
module CHIP ( clk, rst_n, mem_read_D, mem_write_D, mem_addr_D, mem_wdata_D, 
        mem_rdata_D, mem_ready_D, mem_read_I, mem_write_I, mem_addr_I, 
        mem_wdata_I, mem_rdata_I, mem_ready_I, DCACHE_addr, DCACHE_wdata, 
        DCACHE_wen );
  output [31:4] mem_addr_D;
  output [127:0] mem_wdata_D;
  input [127:0] mem_rdata_D;
  output [31:4] mem_addr_I;
  output [127:0] mem_wdata_I;
  input [127:0] mem_rdata_I;
  output [29:0] DCACHE_addr;
  output [31:0] DCACHE_wdata;
  input clk, rst_n, mem_ready_D, mem_ready_I;
  output mem_read_D, mem_write_D, mem_read_I, mem_write_I, DCACHE_wen;
  wire   n10165, n10166, n10167, n10168, n10169, n10170, n10171, n10172,
         n10173, n10174, n10175, n10176, n10177, n10178, n10179, n10180,
         n10181, n10182, n10183, n10184, n10185, n10186, n10187, n10188,
         n10189, n10190, n10191, n10192, n10193, n10194, n10195, n10196,
         n10197, n10198, n10199, n10200, n10201, n10202, n10203, n10204,
         n10205, n10206, n10207, n10208, n10209, n10210, n10211, n10212,
         n10213, n10214, n10215, n10216, n10217, n10218, n10219, n10220,
         n10221, n10222, n10223, n10224, n10225, n10226, n10227, n10228,
         n10229, n10230, n10231, n10232, n10233, n10234, n10235, n10236,
         n10237, n10238, n10239, n10240, n10241, n10242, n10243, n10244,
         n10245, n10246, n10247, n10248, n10249, n10250, n10251, n10252,
         n10253, n10254, n10255, n10256, n10257, n10258, n10259, n10260,
         n10261, n10262, n10263, n10264, n10265, n10266, n10267, n10268,
         n10269, n10270, n10271, n10272, n10273, n10274, n10275, n10276,
         n10277, n10278, n10279, n10280, n10281, n10282, n10283, n10284,
         n10285, n10286, n10287, n10288, n10289, n10290, n10291, n10292,
         n10293, n10294, n10295, n10296, n10297, n10298, n10299, n10300,
         n10301, n10302, n10303, n10304, n10305, n10306, n10307, n10308,
         n10309, n10310, n10311, n10312, n10313, n10314, n10315, n10316,
         n10317, n10318, n10319, n10320, n10321, n10322, n10323, n10324,
         n10325, n10326, n10327, n10328, n10329, n10330, n10331, n10332,
         n10333, n10334, n10335, n10336, n10337, n10338, n10339, n10340,
         n10341, n10342, n10343, n10344, n10345, n10346, n10347, n10348,
         n10349, n10350, n10351, n10352, n10353, n10354, n10355, n10356,
         DCACHE_ren, \i_MIPS/n563 , \i_MIPS/n562 , \i_MIPS/n561 ,
         \i_MIPS/n560 , \i_MIPS/n559 , \i_MIPS/n558 , \i_MIPS/n557 ,
         \i_MIPS/n556 , \i_MIPS/n555 , \i_MIPS/n554 , \i_MIPS/n553 ,
         \i_MIPS/n552 , \i_MIPS/n551 , \i_MIPS/n550 , \i_MIPS/n549 ,
         \i_MIPS/n548 , \i_MIPS/n547 , \i_MIPS/n546 , \i_MIPS/n545 ,
         \i_MIPS/n544 , \i_MIPS/n543 , \i_MIPS/n542 , \i_MIPS/n541 ,
         \i_MIPS/n540 , \i_MIPS/n539 , \i_MIPS/n538 , \i_MIPS/n537 ,
         \i_MIPS/n536 , \i_MIPS/n535 , \i_MIPS/n534 , \i_MIPS/n533 ,
         \i_MIPS/n532 , \i_MIPS/n531 , \i_MIPS/n530 , \i_MIPS/n529 ,
         \i_MIPS/n528 , \i_MIPS/n527 , \i_MIPS/n526 , \i_MIPS/n525 ,
         \i_MIPS/n524 , \i_MIPS/n523 , \i_MIPS/n522 , \i_MIPS/n521 ,
         \i_MIPS/n520 , \i_MIPS/n519 , \i_MIPS/n518 , \i_MIPS/n517 ,
         \i_MIPS/n516 , \i_MIPS/n515 , \i_MIPS/n514 , \i_MIPS/n513 ,
         \i_MIPS/n512 , \i_MIPS/n511 , \i_MIPS/n510 , \i_MIPS/n509 ,
         \i_MIPS/n508 , \i_MIPS/n507 , \i_MIPS/n506 , \i_MIPS/n505 ,
         \i_MIPS/n504 , \i_MIPS/n503 , \i_MIPS/n502 , \i_MIPS/n501 ,
         \i_MIPS/n500 , \i_MIPS/n499 , \i_MIPS/n498 , \i_MIPS/n497 ,
         \i_MIPS/n496 , \i_MIPS/n495 , \i_MIPS/n494 , \i_MIPS/n493 ,
         \i_MIPS/n492 , \i_MIPS/n491 , \i_MIPS/n490 , \i_MIPS/n489 ,
         \i_MIPS/n488 , \i_MIPS/n487 , \i_MIPS/n486 , \i_MIPS/n485 ,
         \i_MIPS/n484 , \i_MIPS/n483 , \i_MIPS/n482 , \i_MIPS/n481 ,
         \i_MIPS/n480 , \i_MIPS/n479 , \i_MIPS/n478 , \i_MIPS/n477 ,
         \i_MIPS/n476 , \i_MIPS/n475 , \i_MIPS/n474 , \i_MIPS/n473 ,
         \i_MIPS/n472 , \i_MIPS/n471 , \i_MIPS/n470 , \i_MIPS/n469 ,
         \i_MIPS/n468 , \i_MIPS/n467 , \i_MIPS/n466 , \i_MIPS/n465 ,
         \i_MIPS/n464 , \i_MIPS/n463 , \i_MIPS/n462 , \i_MIPS/n461 ,
         \i_MIPS/n460 , \i_MIPS/n459 , \i_MIPS/n458 , \i_MIPS/n457 ,
         \i_MIPS/n456 , \i_MIPS/n455 , \i_MIPS/n454 , \i_MIPS/n453 ,
         \i_MIPS/n452 , \i_MIPS/n451 , \i_MIPS/n450 , \i_MIPS/n449 ,
         \i_MIPS/n448 , \i_MIPS/n447 , \i_MIPS/n446 , \i_MIPS/n445 ,
         \i_MIPS/n444 , \i_MIPS/n443 , \i_MIPS/n442 , \i_MIPS/n441 ,
         \i_MIPS/n440 , \i_MIPS/n439 , \i_MIPS/n438 , \i_MIPS/n437 ,
         \i_MIPS/n436 , \i_MIPS/n435 , \i_MIPS/n434 , \i_MIPS/n433 ,
         \i_MIPS/n432 , \i_MIPS/n431 , \i_MIPS/n430 , \i_MIPS/n429 ,
         \i_MIPS/n428 , \i_MIPS/n427 , \i_MIPS/n426 , \i_MIPS/n425 ,
         \i_MIPS/n424 , \i_MIPS/n423 , \i_MIPS/n422 , \i_MIPS/n421 ,
         \i_MIPS/n420 , \i_MIPS/n419 , \i_MIPS/n418 , \i_MIPS/n417 ,
         \i_MIPS/n416 , \i_MIPS/n415 , \i_MIPS/n414 , \i_MIPS/n413 ,
         \i_MIPS/n412 , \i_MIPS/n411 , \i_MIPS/n410 , \i_MIPS/n409 ,
         \i_MIPS/n408 , \i_MIPS/n407 , \i_MIPS/n406 , \i_MIPS/n405 ,
         \i_MIPS/n404 , \i_MIPS/n403 , \i_MIPS/n402 , \i_MIPS/n401 ,
         \i_MIPS/n400 , \i_MIPS/n399 , \i_MIPS/n398 , \i_MIPS/n397 ,
         \i_MIPS/n396 , \i_MIPS/n395 , \i_MIPS/n394 , \i_MIPS/n393 ,
         \i_MIPS/n392 , \i_MIPS/n391 , \i_MIPS/n390 , \i_MIPS/n389 ,
         \i_MIPS/n388 , \i_MIPS/n387 , \i_MIPS/n386 , \i_MIPS/n385 ,
         \i_MIPS/n384 , \i_MIPS/n383 , \i_MIPS/n382 , \i_MIPS/n381 ,
         \i_MIPS/n380 , \i_MIPS/n379 , \i_MIPS/n378 , \i_MIPS/n377 ,
         \i_MIPS/n376 , \i_MIPS/n375 , \i_MIPS/n374 , \i_MIPS/n373 ,
         \i_MIPS/n372 , \i_MIPS/n371 , \i_MIPS/n370 , \i_MIPS/n369 ,
         \i_MIPS/n368 , \i_MIPS/n367 , \i_MIPS/n366 , \i_MIPS/n365 ,
         \i_MIPS/n364 , \i_MIPS/n363 , \i_MIPS/n362 , \i_MIPS/n361 ,
         \i_MIPS/n360 , \i_MIPS/n359 , \i_MIPS/n358 , \i_MIPS/n357 ,
         \i_MIPS/n356 , \i_MIPS/n355 , \i_MIPS/n354 , \i_MIPS/n353 ,
         \i_MIPS/n352 , \i_MIPS/n351 , \i_MIPS/n350 , \i_MIPS/n349 ,
         \i_MIPS/n348 , \i_MIPS/n347 , \i_MIPS/n346 , \i_MIPS/n345 ,
         \i_MIPS/n344 , \i_MIPS/n343 , \i_MIPS/n342 , \i_MIPS/n341 ,
         \i_MIPS/n340 , \i_MIPS/n339 , \i_MIPS/n338 , \i_MIPS/n337 ,
         \i_MIPS/n336 , \i_MIPS/n335 , \i_MIPS/n334 , \i_MIPS/n333 ,
         \i_MIPS/n332 , \i_MIPS/n331 , \i_MIPS/n330 , \i_MIPS/n329 ,
         \i_MIPS/n328 , \i_MIPS/n327 , \i_MIPS/n326 , \i_MIPS/n325 ,
         \i_MIPS/n324 , \i_MIPS/n323 , \i_MIPS/n322 , \i_MIPS/n321 ,
         \i_MIPS/n320 , \i_MIPS/n319 , \i_MIPS/n318 , \i_MIPS/n317 ,
         \i_MIPS/n316 , \i_MIPS/n315 , \i_MIPS/n314 , \i_MIPS/n313 ,
         \i_MIPS/n312 , \i_MIPS/n311 , \i_MIPS/n310 , \i_MIPS/n309 ,
         \i_MIPS/n308 , \i_MIPS/n307 , \i_MIPS/n306 , \i_MIPS/n305 ,
         \i_MIPS/n304 , \i_MIPS/n303 , \i_MIPS/n302 , \i_MIPS/n301 ,
         \i_MIPS/n300 , \i_MIPS/n299 , \i_MIPS/n298 , \i_MIPS/n297 ,
         \i_MIPS/n296 , \i_MIPS/n295 , \i_MIPS/n294 , \i_MIPS/n293 ,
         \i_MIPS/n292 , \i_MIPS/n291 , \i_MIPS/n290 , \i_MIPS/n289 ,
         \i_MIPS/n288 , \i_MIPS/n287 , \i_MIPS/n286 , \i_MIPS/n285 ,
         \i_MIPS/n284 , \i_MIPS/n283 , \i_MIPS/n282 , \i_MIPS/n281 ,
         \i_MIPS/n280 , \i_MIPS/n279 , \i_MIPS/n278 , \i_MIPS/n277 ,
         \i_MIPS/n276 , \i_MIPS/n275 , \i_MIPS/n274 , \i_MIPS/n273 ,
         \i_MIPS/n272 , \i_MIPS/n271 , \i_MIPS/n270 , \i_MIPS/n269 ,
         \i_MIPS/n268 , \i_MIPS/n267 , \i_MIPS/n266 , \i_MIPS/n265 ,
         \i_MIPS/n264 , \i_MIPS/n263 , \i_MIPS/n262 , \i_MIPS/n261 ,
         \i_MIPS/n260 , \i_MIPS/n259 , \i_MIPS/n258 , \i_MIPS/n257 ,
         \i_MIPS/n256 , \i_MIPS/n255 , \i_MIPS/n254 , \i_MIPS/n253 ,
         \i_MIPS/n252 , \i_MIPS/n251 , \i_MIPS/n250 , \i_MIPS/n249 ,
         \i_MIPS/n248 , \i_MIPS/n247 , \i_MIPS/n246 , \i_MIPS/n245 ,
         \i_MIPS/n244 , \i_MIPS/n243 , \i_MIPS/n242 , \i_MIPS/n241 ,
         \i_MIPS/n240 , \i_MIPS/n239 , \i_MIPS/n238 , \i_MIPS/n237 ,
         \i_MIPS/n236 , \i_MIPS/n235 , \i_MIPS/n234 , \i_MIPS/n233 ,
         \i_MIPS/n232 , \i_MIPS/n231 , \i_MIPS/n230 , \i_MIPS/n229 ,
         \i_MIPS/n228 , \i_MIPS/n227 , \i_MIPS/n226 , \i_MIPS/n225 ,
         \i_MIPS/n224 , \i_MIPS/n223 , \i_MIPS/n222 , \i_MIPS/n221 ,
         \i_MIPS/n220 , \i_MIPS/n219 , \i_MIPS/n218 , \i_MIPS/n217 ,
         \i_MIPS/n216 , \i_MIPS/n215 , \i_MIPS/n214 , \i_MIPS/n213 ,
         \i_MIPS/n212 , \i_MIPS/n211 , \i_MIPS/n210 , \i_MIPS/n209 ,
         \i_MIPS/n208 , \i_MIPS/n207 , \i_MIPS/n206 , \i_MIPS/n205 ,
         \i_MIPS/n204 , \i_MIPS/n203 , \i_MIPS/n202 , \i_MIPS/n201 ,
         \i_MIPS/n200 , \i_MIPS/n199 , \i_MIPS/n198 , \i_MIPS/n197 ,
         \i_MIPS/n196 , \i_MIPS/n195 , \i_MIPS/n194 , \i_MIPS/n193 ,
         \i_MIPS/n192 , \i_MIPS/n191 , \i_MIPS/n190 , \i_MIPS/n189 ,
         \i_MIPS/n188 , \i_MIPS/n187 , \i_MIPS/n186 , \i_MIPS/n185 ,
         \i_MIPS/n184 , \i_MIPS/n183 , \i_MIPS/n182 , \i_MIPS/n181 ,
         \i_MIPS/n180 , \i_MIPS/n178 , \i_MIPS/n177 , \i_MIPS/n176 ,
         \i_MIPS/n175 , \i_MIPS/n174 , \i_MIPS/n173 , \i_MIPS/n172 ,
         \i_MIPS/n171 , \i_MIPS/n170 , \i_MIPS/n169 , \i_MIPS/n168 ,
         \i_MIPS/n167 , \i_MIPS/n166 , \i_MIPS/n165 , \i_MIPS/n164 ,
         \i_MIPS/n163 , \i_MIPS/n162 , \i_MIPS/n161 , \i_MIPS/n160 ,
         \i_MIPS/n159 , \i_MIPS/N120 , \i_MIPS/N119 , \i_MIPS/N118 ,
         \i_MIPS/N117 , \i_MIPS/N116 , \i_MIPS/N115 , \i_MIPS/N114 ,
         \i_MIPS/N113 , \i_MIPS/N112 , \i_MIPS/N111 , \i_MIPS/N110 ,
         \i_MIPS/N109 , \i_MIPS/N108 , \i_MIPS/N107 , \i_MIPS/N106 ,
         \i_MIPS/N105 , \i_MIPS/N104 , \i_MIPS/N103 , \i_MIPS/N102 ,
         \i_MIPS/N101 , \i_MIPS/N100 , \i_MIPS/N99 , \i_MIPS/N98 ,
         \i_MIPS/N97 , \i_MIPS/N96 , \i_MIPS/N95 , \i_MIPS/N94 , \i_MIPS/N93 ,
         \i_MIPS/N92 , \i_MIPS/N91 , \i_MIPS/N90 , \i_MIPS/N89 , \i_MIPS/N88 ,
         \i_MIPS/N87 , \i_MIPS/N86 , \i_MIPS/N85 , \i_MIPS/N84 , \i_MIPS/N83 ,
         \i_MIPS/N82 , \i_MIPS/N81 , \i_MIPS/N80 , \i_MIPS/N79 , \i_MIPS/N78 ,
         \i_MIPS/N77 , \i_MIPS/N76 , \i_MIPS/N75 , \i_MIPS/N74 , \i_MIPS/N73 ,
         \i_MIPS/N72 , \i_MIPS/N71 , \i_MIPS/N70 , \i_MIPS/N69 , \i_MIPS/N68 ,
         \i_MIPS/N67 , \i_MIPS/N66 , \i_MIPS/N65 , \i_MIPS/N64 , \i_MIPS/N63 ,
         \i_MIPS/N62 , \i_MIPS/N61 , \i_MIPS/N60 , \i_MIPS/N59 , \i_MIPS/N58 ,
         \i_MIPS/N57 , \i_MIPS/N56 , \i_MIPS/N55 , \i_MIPS/N54 , \i_MIPS/N53 ,
         \i_MIPS/N52 , \i_MIPS/N51 , \i_MIPS/N50 , \i_MIPS/N49 , \i_MIPS/N48 ,
         \i_MIPS/N47 , \i_MIPS/N46 , \i_MIPS/N45 , \i_MIPS/N44 , \i_MIPS/N43 ,
         \i_MIPS/N42 , \i_MIPS/N41 , \i_MIPS/N40 , \i_MIPS/N39 , \i_MIPS/N38 ,
         \i_MIPS/N37 , \i_MIPS/N36 , \i_MIPS/N35 , \i_MIPS/N34 , \i_MIPS/N33 ,
         \i_MIPS/N32 , \i_MIPS/N31 , \i_MIPS/N30 , \i_MIPS/N29 , \i_MIPS/N28 ,
         \i_MIPS/N27 , \i_MIPS/N26 , \i_MIPS/N25 , \i_MIPS/N24 , \i_MIPS/N23 ,
         \i_MIPS/ALUin1[30] , \i_MIPS/ALUin1[29] , \i_MIPS/ALUin1[28] ,
         \i_MIPS/ALUin1[27] , \i_MIPS/ALUin1[26] , \i_MIPS/ALUin1[25] ,
         \i_MIPS/ALUin1[24] , \i_MIPS/ALUin1[23] , \i_MIPS/ALUin1[22] ,
         \i_MIPS/ALUin1[21] , \i_MIPS/ALUin1[20] , \i_MIPS/ALUin1[19] ,
         \i_MIPS/ALUin1[18] , \i_MIPS/ALUin1[17] , \i_MIPS/ALUin1[16] ,
         \i_MIPS/ALUin1[15] , \i_MIPS/ALUin1[14] , \i_MIPS/ALUin1[13] ,
         \i_MIPS/ALUin1[12] , \i_MIPS/ALUin1[11] , \i_MIPS/ALUin1[10] ,
         \i_MIPS/ALUin1[9] , \i_MIPS/ALUin1[8] , \i_MIPS/ALUin1[7] ,
         \i_MIPS/ALUin1[6] , \i_MIPS/ALUin1[5] , \i_MIPS/ALUin1[4] ,
         \i_MIPS/ALUin1[3] , \i_MIPS/ALUin1[2] , \i_MIPS/ALUin1[1] ,
         \i_MIPS/ALUin1[0] , \i_MIPS/ALUOp[0] , \i_MIPS/ALUOp[1] ,
         \i_MIPS/EX_MEM_0 , \i_MIPS/EX_MEM_1 , \i_MIPS/EX_MEM[5] ,
         \i_MIPS/EX_MEM[6] , \i_MIPS/EX_MEM_74 , \i_MIPS/EX_MEM_next[69] ,
         \i_MIPS/EX_MEM_next[70] , \i_MIPS/EX_MEM_next[71] ,
         \i_MIPS/Sign_Extend_ID[31] , \i_MIPS/Sign_Extend_ID[8] ,
         \i_MIPS/Sign_Extend_ID[6] , \i_MIPS/Sign_Extend_ID[5] ,
         \i_MIPS/Sign_Extend_ID[4] , \i_MIPS/Sign_Extend_ID[3] ,
         \i_MIPS/Sign_Extend_ID[2] , \i_MIPS/Sign_Extend_ID[1] ,
         \i_MIPS/Sign_Extend_ID[0] , \i_MIPS/ID_EX_0 , \i_MIPS/ID_EX_3 ,
         \i_MIPS/ID_EX_5 , \i_MIPS/ID_EX[47] , \i_MIPS/ID_EX[49] ,
         \i_MIPS/ID_EX[50] , \i_MIPS/ID_EX[52] , \i_MIPS/ID_EX[57] ,
         \i_MIPS/ID_EX[58] , \i_MIPS/ID_EX[59] , \i_MIPS/ID_EX[60] ,
         \i_MIPS/ID_EX[61] , \i_MIPS/ID_EX[62] , \i_MIPS/ID_EX[63] ,
         \i_MIPS/ID_EX[64] , \i_MIPS/ID_EX[65] , \i_MIPS/ID_EX[66] ,
         \i_MIPS/ID_EX[67] , \i_MIPS/ID_EX[68] , \i_MIPS/ID_EX[69] ,
         \i_MIPS/ID_EX[70] , \i_MIPS/ID_EX[71] , \i_MIPS/ID_EX[73] ,
         \i_MIPS/ID_EX[74] , \i_MIPS/ID_EX[75] , \i_MIPS/ID_EX[76] ,
         \i_MIPS/ID_EX[77] , \i_MIPS/ID_EX[78] , \i_MIPS/ID_EX[79] ,
         \i_MIPS/ID_EX[80] , \i_MIPS/ID_EX[82] , \i_MIPS/ID_EX[83] ,
         \i_MIPS/ID_EX[84] , \i_MIPS/ID_EX[85] , \i_MIPS/ID_EX[86] ,
         \i_MIPS/ID_EX[87] , \i_MIPS/ID_EX[88] , \i_MIPS/ID_EX[89] ,
         \i_MIPS/ID_EX[90] , \i_MIPS/ID_EX[91] , \i_MIPS/ID_EX[92] ,
         \i_MIPS/ID_EX[93] , \i_MIPS/ID_EX[94] , \i_MIPS/ID_EX[95] ,
         \i_MIPS/ID_EX[96] , \i_MIPS/ID_EX[97] , \i_MIPS/ID_EX[98] ,
         \i_MIPS/ID_EX[99] , \i_MIPS/ID_EX[100] , \i_MIPS/ID_EX[101] ,
         \i_MIPS/ID_EX[102] , \i_MIPS/ID_EX[103] , \i_MIPS/ID_EX[104] ,
         \i_MIPS/ID_EX[105] , \i_MIPS/ID_EX[106] , \i_MIPS/ID_EX[107] ,
         \i_MIPS/ID_EX[109] , \i_MIPS/ID_EX[110] , \i_MIPS/ID_EX[111] ,
         \i_MIPS/ID_EX[112] , \i_MIPS/ID_EX[113] , \i_MIPS/ID_EX[114] ,
         \i_MIPS/ID_EX[115] , \i_MIPS/control_out[7] , \i_MIPS/control_out[0] ,
         \i_MIPS/Reg_W[0] , \i_MIPS/Reg_W[1] , \i_MIPS/Reg_W[2] ,
         \i_MIPS/Reg_W[3] , \i_MIPS/Reg_W[4] , \i_MIPS/IR_ID[16] ,
         \i_MIPS/IR_ID[17] , \i_MIPS/IR_ID[18] , \i_MIPS/IR_ID[19] ,
         \i_MIPS/IR_ID[20] , \i_MIPS/IR_ID[21] , \i_MIPS/IR_ID[22] ,
         \i_MIPS/IR_ID[23] , \i_MIPS/IR_ID[24] , \i_MIPS/IR_ID[25] ,
         \i_MIPS/IR_ID[26] , \i_MIPS/IR_ID[27] , \i_MIPS/IR_ID[28] ,
         \i_MIPS/IR_ID[29] , \i_MIPS/IR_ID[30] , \i_MIPS/IR_ID[31] ,
         \i_MIPS/IF_ID_0 , \i_MIPS/IF_ID_1 , \i_MIPS/IF_ID_28 ,
         \i_MIPS/IF_ID_29 , \i_MIPS/IF_ID_30 , \i_MIPS/IF_ID_31 ,
         \i_MIPS/IF_ID[97] , \i_MIPS/IF_ID[96] , \i_MIPS/IF_ID[95] ,
         \i_MIPS/IF_ID[94] , \i_MIPS/IF_ID[93] , \i_MIPS/IF_ID[92] ,
         \i_MIPS/IF_ID[91] , \i_MIPS/IF_ID[90] , \i_MIPS/IF_ID[89] ,
         \i_MIPS/IF_ID[88] , \i_MIPS/IF_ID[87] , \i_MIPS/IF_ID[86] ,
         \i_MIPS/IF_ID[85] , \i_MIPS/IF_ID[84] , \i_MIPS/IF_ID[83] ,
         \i_MIPS/IF_ID[82] , \i_MIPS/IF_ID[81] , \i_MIPS/IF_ID[80] ,
         \i_MIPS/IF_ID[79] , \i_MIPS/IF_ID[78] , \i_MIPS/IF_ID[77] ,
         \i_MIPS/IF_ID[76] , \i_MIPS/IF_ID[75] , \i_MIPS/IF_ID[74] ,
         \i_MIPS/IF_ID[73] , \i_MIPS/IF_ID[72] , \i_MIPS/IF_ID[71] ,
         \i_MIPS/IF_ID[70] , \i_MIPS/IF_ID[69] , \i_MIPS/IF_ID[68] ,
         \i_MIPS/IF_ID[67] , \i_MIPS/IF_ID[66] , \i_MIPS/IF_ID[65] ,
         \i_MIPS/IF_ID[64] , \i_MIPS/PC_o[1] , \i_MIPS/BranchAddr[0] ,
         \D_cache/n2106 , \D_cache/n2105 , \D_cache/n2104 , \D_cache/n2103 ,
         \D_cache/n2102 , \D_cache/n2101 , \D_cache/n2100 , \D_cache/n2099 ,
         \D_cache/n2098 , \D_cache/n2097 , \D_cache/n2096 , \D_cache/n2095 ,
         \D_cache/n2094 , \D_cache/n2093 , \D_cache/n2092 , \D_cache/n2091 ,
         \D_cache/n2090 , \D_cache/n2089 , \D_cache/n2088 , \D_cache/n2087 ,
         \D_cache/n2086 , \D_cache/n2085 , \D_cache/n2084 , \D_cache/n2083 ,
         \D_cache/n2082 , \D_cache/n2081 , \D_cache/n2080 , \D_cache/n2079 ,
         \D_cache/n2078 , \D_cache/n2077 , \D_cache/n2076 , \D_cache/n2075 ,
         \D_cache/n2074 , \D_cache/n2073 , \D_cache/n2072 , \D_cache/n2071 ,
         \D_cache/n2070 , \D_cache/n2069 , \D_cache/n2068 , \D_cache/n2067 ,
         \D_cache/n2066 , \D_cache/n2065 , \D_cache/n2064 , \D_cache/n2063 ,
         \D_cache/n2062 , \D_cache/n2061 , \D_cache/n2060 , \D_cache/n2059 ,
         \D_cache/n2058 , \D_cache/n2057 , \D_cache/n2056 , \D_cache/n2055 ,
         \D_cache/n2054 , \D_cache/n2053 , \D_cache/n2052 , \D_cache/n2051 ,
         \D_cache/n2050 , \D_cache/n2049 , \D_cache/n2048 , \D_cache/n2047 ,
         \D_cache/n2046 , \D_cache/n2045 , \D_cache/n2044 , \D_cache/n2043 ,
         \D_cache/n2042 , \D_cache/n2041 , \D_cache/n2040 , \D_cache/n2039 ,
         \D_cache/n2038 , \D_cache/n2037 , \D_cache/n2036 , \D_cache/n2035 ,
         \D_cache/n2034 , \D_cache/n2033 , \D_cache/n2032 , \D_cache/n2031 ,
         \D_cache/n2030 , \D_cache/n2029 , \D_cache/n2028 , \D_cache/n2027 ,
         \D_cache/n2026 , \D_cache/n2025 , \D_cache/n2024 , \D_cache/n2023 ,
         \D_cache/n2022 , \D_cache/n2021 , \D_cache/n2020 , \D_cache/n2019 ,
         \D_cache/n2018 , \D_cache/n2017 , \D_cache/n2016 , \D_cache/n2015 ,
         \D_cache/n2014 , \D_cache/n2013 , \D_cache/n2012 , \D_cache/n2011 ,
         \D_cache/n2010 , \D_cache/n2009 , \D_cache/n2008 , \D_cache/n2007 ,
         \D_cache/n2006 , \D_cache/n2005 , \D_cache/n2004 , \D_cache/n2003 ,
         \D_cache/n2002 , \D_cache/n2001 , \D_cache/n2000 , \D_cache/n1999 ,
         \D_cache/n1998 , \D_cache/n1997 , \D_cache/n1996 , \D_cache/n1995 ,
         \D_cache/n1994 , \D_cache/n1993 , \D_cache/n1992 , \D_cache/n1991 ,
         \D_cache/n1990 , \D_cache/n1989 , \D_cache/n1988 , \D_cache/n1987 ,
         \D_cache/n1986 , \D_cache/n1985 , \D_cache/n1984 , \D_cache/n1983 ,
         \D_cache/n1982 , \D_cache/n1981 , \D_cache/n1980 , \D_cache/n1979 ,
         \D_cache/n1978 , \D_cache/n1977 , \D_cache/n1976 , \D_cache/n1975 ,
         \D_cache/n1974 , \D_cache/n1973 , \D_cache/n1972 , \D_cache/n1971 ,
         \D_cache/n1970 , \D_cache/n1969 , \D_cache/n1968 , \D_cache/n1967 ,
         \D_cache/n1966 , \D_cache/n1965 , \D_cache/n1964 , \D_cache/n1963 ,
         \D_cache/n1962 , \D_cache/n1961 , \D_cache/n1960 , \D_cache/n1959 ,
         \D_cache/n1958 , \D_cache/n1957 , \D_cache/n1956 , \D_cache/n1955 ,
         \D_cache/n1954 , \D_cache/n1953 , \D_cache/n1952 , \D_cache/n1951 ,
         \D_cache/n1950 , \D_cache/n1949 , \D_cache/n1948 , \D_cache/n1947 ,
         \D_cache/n1946 , \D_cache/n1945 , \D_cache/n1944 , \D_cache/n1943 ,
         \D_cache/n1942 , \D_cache/n1941 , \D_cache/n1940 , \D_cache/n1939 ,
         \D_cache/n1938 , \D_cache/n1937 , \D_cache/n1936 , \D_cache/n1935 ,
         \D_cache/n1934 , \D_cache/n1933 , \D_cache/n1932 , \D_cache/n1931 ,
         \D_cache/n1930 , \D_cache/n1929 , \D_cache/n1928 , \D_cache/n1927 ,
         \D_cache/n1926 , \D_cache/n1925 , \D_cache/n1860 , \D_cache/n1859 ,
         \D_cache/n1858 , \D_cache/n1857 , \D_cache/n1856 , \D_cache/n1855 ,
         \D_cache/n1854 , \D_cache/n1853 , \D_cache/n1852 , \D_cache/n1851 ,
         \D_cache/n1850 , \D_cache/n1849 , \D_cache/n1848 , \D_cache/n1847 ,
         \D_cache/n1846 , \D_cache/n1845 , \D_cache/n1844 , \D_cache/n1843 ,
         \D_cache/n1842 , \D_cache/n1841 , \D_cache/n1840 , \D_cache/n1839 ,
         \D_cache/n1838 , \D_cache/n1837 , \D_cache/n1836 , \D_cache/n1835 ,
         \D_cache/n1834 , \D_cache/n1833 , \D_cache/n1832 , \D_cache/n1831 ,
         \D_cache/n1830 , \D_cache/n1829 , \D_cache/n1828 , \D_cache/n1827 ,
         \D_cache/n1826 , \D_cache/n1825 , \D_cache/n1824 , \D_cache/n1823 ,
         \D_cache/n1822 , \D_cache/n1821 , \D_cache/n1820 , \D_cache/n1819 ,
         \D_cache/n1818 , \D_cache/n1817 , \D_cache/n1816 , \D_cache/n1815 ,
         \D_cache/n1814 , \D_cache/n1813 , \D_cache/n1812 , \D_cache/n1811 ,
         \D_cache/n1810 , \D_cache/n1809 , \D_cache/n1808 , \D_cache/n1807 ,
         \D_cache/n1806 , \D_cache/n1805 , \D_cache/n1804 , \D_cache/n1803 ,
         \D_cache/n1802 , \D_cache/n1801 , \D_cache/n1800 , \D_cache/n1799 ,
         \D_cache/n1798 , \D_cache/n1797 , \D_cache/n1796 , \D_cache/n1795 ,
         \D_cache/n1794 , \D_cache/n1793 , \D_cache/n1792 , \D_cache/n1791 ,
         \D_cache/n1790 , \D_cache/n1789 , \D_cache/n1788 , \D_cache/n1787 ,
         \D_cache/n1786 , \D_cache/n1785 , \D_cache/n1784 , \D_cache/n1783 ,
         \D_cache/n1782 , \D_cache/n1781 , \D_cache/n1780 , \D_cache/n1779 ,
         \D_cache/n1778 , \D_cache/n1777 , \D_cache/n1776 , \D_cache/n1775 ,
         \D_cache/n1774 , \D_cache/n1773 , \D_cache/n1772 , \D_cache/n1771 ,
         \D_cache/n1770 , \D_cache/n1769 , \D_cache/n1768 , \D_cache/n1767 ,
         \D_cache/n1766 , \D_cache/n1765 , \D_cache/n1764 , \D_cache/n1763 ,
         \D_cache/n1762 , \D_cache/n1761 , \D_cache/n1760 , \D_cache/n1759 ,
         \D_cache/n1758 , \D_cache/n1757 , \D_cache/n1756 , \D_cache/n1755 ,
         \D_cache/n1754 , \D_cache/n1753 , \D_cache/n1752 , \D_cache/n1751 ,
         \D_cache/n1750 , \D_cache/n1749 , \D_cache/n1748 , \D_cache/n1747 ,
         \D_cache/n1746 , \D_cache/n1745 , \D_cache/n1744 , \D_cache/n1743 ,
         \D_cache/n1742 , \D_cache/n1741 , \D_cache/n1740 , \D_cache/n1739 ,
         \D_cache/n1738 , \D_cache/n1737 , \D_cache/n1736 , \D_cache/n1735 ,
         \D_cache/n1734 , \D_cache/n1733 , \D_cache/n1732 , \D_cache/n1731 ,
         \D_cache/n1730 , \D_cache/n1729 , \D_cache/n1728 , \D_cache/n1727 ,
         \D_cache/n1726 , \D_cache/n1725 , \D_cache/n1724 , \D_cache/n1723 ,
         \D_cache/n1722 , \D_cache/n1721 , \D_cache/n1720 , \D_cache/n1719 ,
         \D_cache/n1718 , \D_cache/n1717 , \D_cache/n1716 , \D_cache/n1715 ,
         \D_cache/n1714 , \D_cache/n1713 , \D_cache/n1712 , \D_cache/n1711 ,
         \D_cache/n1710 , \D_cache/n1709 , \D_cache/n1708 , \D_cache/n1707 ,
         \D_cache/n1706 , \D_cache/n1705 , \D_cache/n1704 , \D_cache/n1703 ,
         \D_cache/n1702 , \D_cache/n1701 , \D_cache/n1700 , \D_cache/n1699 ,
         \D_cache/n1698 , \D_cache/n1697 , \D_cache/n1696 , \D_cache/n1695 ,
         \D_cache/n1694 , \D_cache/n1693 , \D_cache/n1692 , \D_cache/n1691 ,
         \D_cache/n1690 , \D_cache/n1689 , \D_cache/n1688 , \D_cache/n1687 ,
         \D_cache/n1686 , \D_cache/n1685 , \D_cache/n1684 , \D_cache/n1683 ,
         \D_cache/n1682 , \D_cache/n1681 , \D_cache/n1680 , \D_cache/n1679 ,
         \D_cache/n1678 , \D_cache/n1677 , \D_cache/n1676 , \D_cache/n1675 ,
         \D_cache/n1674 , \D_cache/n1673 , \D_cache/n1672 , \D_cache/n1671 ,
         \D_cache/n1670 , \D_cache/n1669 , \D_cache/n1668 , \D_cache/n1667 ,
         \D_cache/n1666 , \D_cache/n1665 , \D_cache/n1664 , \D_cache/n1663 ,
         \D_cache/n1662 , \D_cache/n1661 , \D_cache/n1660 , \D_cache/n1659 ,
         \D_cache/n1658 , \D_cache/n1657 , \D_cache/n1656 , \D_cache/n1655 ,
         \D_cache/n1654 , \D_cache/n1653 , \D_cache/n1652 , \D_cache/n1651 ,
         \D_cache/n1650 , \D_cache/n1649 , \D_cache/n1648 , \D_cache/n1647 ,
         \D_cache/n1646 , \D_cache/n1645 , \D_cache/n1644 , \D_cache/n1643 ,
         \D_cache/n1642 , \D_cache/n1641 , \D_cache/n1640 , \D_cache/n1639 ,
         \D_cache/n1638 , \D_cache/n1637 , \D_cache/n1636 , \D_cache/n1635 ,
         \D_cache/n1634 , \D_cache/n1633 , \D_cache/n1632 , \D_cache/n1631 ,
         \D_cache/n1630 , \D_cache/n1629 , \D_cache/n1628 , \D_cache/n1627 ,
         \D_cache/n1626 , \D_cache/n1625 , \D_cache/n1624 , \D_cache/n1623 ,
         \D_cache/n1622 , \D_cache/n1621 , \D_cache/n1620 , \D_cache/n1619 ,
         \D_cache/n1618 , \D_cache/n1617 , \D_cache/n1616 , \D_cache/n1615 ,
         \D_cache/n1614 , \D_cache/n1613 , \D_cache/n1612 , \D_cache/n1611 ,
         \D_cache/n1610 , \D_cache/n1609 , \D_cache/n1608 , \D_cache/n1607 ,
         \D_cache/n1606 , \D_cache/n1605 , \D_cache/n1604 , \D_cache/n1603 ,
         \D_cache/n1602 , \D_cache/n1601 , \D_cache/n1600 , \D_cache/n1599 ,
         \D_cache/n1598 , \D_cache/n1597 , \D_cache/n1596 , \D_cache/n1595 ,
         \D_cache/n1594 , \D_cache/n1593 , \D_cache/n1592 , \D_cache/n1591 ,
         \D_cache/n1590 , \D_cache/n1589 , \D_cache/n1588 , \D_cache/n1587 ,
         \D_cache/n1586 , \D_cache/n1585 , \D_cache/n1584 , \D_cache/n1583 ,
         \D_cache/n1582 , \D_cache/n1581 , \D_cache/n1580 , \D_cache/n1579 ,
         \D_cache/n1578 , \D_cache/n1577 , \D_cache/n1576 , \D_cache/n1575 ,
         \D_cache/n1574 , \D_cache/n1573 , \D_cache/n1572 , \D_cache/n1571 ,
         \D_cache/n1570 , \D_cache/n1569 , \D_cache/n1568 , \D_cache/n1567 ,
         \D_cache/n1566 , \D_cache/n1565 , \D_cache/n1564 , \D_cache/n1563 ,
         \D_cache/n1562 , \D_cache/n1561 , \D_cache/n1560 , \D_cache/n1559 ,
         \D_cache/n1558 , \D_cache/n1557 , \D_cache/n1556 , \D_cache/n1555 ,
         \D_cache/n1554 , \D_cache/n1553 , \D_cache/n1552 , \D_cache/n1551 ,
         \D_cache/n1550 , \D_cache/n1549 , \D_cache/n1548 , \D_cache/n1547 ,
         \D_cache/n1546 , \D_cache/n1545 , \D_cache/n1544 , \D_cache/n1543 ,
         \D_cache/n1542 , \D_cache/n1541 , \D_cache/n1540 , \D_cache/n1539 ,
         \D_cache/n1538 , \D_cache/n1537 , \D_cache/n1536 , \D_cache/n1535 ,
         \D_cache/n1534 , \D_cache/n1533 , \D_cache/n1532 , \D_cache/n1531 ,
         \D_cache/n1530 , \D_cache/n1529 , \D_cache/n1528 , \D_cache/n1527 ,
         \D_cache/n1526 , \D_cache/n1525 , \D_cache/n1524 , \D_cache/n1523 ,
         \D_cache/n1522 , \D_cache/n1521 , \D_cache/n1520 , \D_cache/n1519 ,
         \D_cache/n1518 , \D_cache/n1517 , \D_cache/n1516 , \D_cache/n1515 ,
         \D_cache/n1514 , \D_cache/n1513 , \D_cache/n1512 , \D_cache/n1511 ,
         \D_cache/n1510 , \D_cache/n1509 , \D_cache/n1508 , \D_cache/n1507 ,
         \D_cache/n1506 , \D_cache/n1505 , \D_cache/n1504 , \D_cache/n1503 ,
         \D_cache/n1502 , \D_cache/n1501 , \D_cache/n1500 , \D_cache/n1499 ,
         \D_cache/n1498 , \D_cache/n1497 , \D_cache/n1496 , \D_cache/n1495 ,
         \D_cache/n1494 , \D_cache/n1493 , \D_cache/n1492 , \D_cache/n1491 ,
         \D_cache/n1490 , \D_cache/n1489 , \D_cache/n1488 , \D_cache/n1487 ,
         \D_cache/n1486 , \D_cache/n1485 , \D_cache/n1484 , \D_cache/n1483 ,
         \D_cache/n1482 , \D_cache/n1481 , \D_cache/n1480 , \D_cache/n1479 ,
         \D_cache/n1478 , \D_cache/n1477 , \D_cache/n1476 , \D_cache/n1475 ,
         \D_cache/n1474 , \D_cache/n1473 , \D_cache/n1472 , \D_cache/n1471 ,
         \D_cache/n1470 , \D_cache/n1469 , \D_cache/n1468 , \D_cache/n1467 ,
         \D_cache/n1466 , \D_cache/n1465 , \D_cache/n1464 , \D_cache/n1463 ,
         \D_cache/n1462 , \D_cache/n1461 , \D_cache/n1460 , \D_cache/n1459 ,
         \D_cache/n1458 , \D_cache/n1457 , \D_cache/n1456 , \D_cache/n1455 ,
         \D_cache/n1454 , \D_cache/n1453 , \D_cache/n1452 , \D_cache/n1451 ,
         \D_cache/n1450 , \D_cache/n1449 , \D_cache/n1448 , \D_cache/n1447 ,
         \D_cache/n1446 , \D_cache/n1445 , \D_cache/n1444 , \D_cache/n1443 ,
         \D_cache/n1442 , \D_cache/n1441 , \D_cache/n1440 , \D_cache/n1439 ,
         \D_cache/n1438 , \D_cache/n1437 , \D_cache/n1436 , \D_cache/n1435 ,
         \D_cache/n1434 , \D_cache/n1433 , \D_cache/n1432 , \D_cache/n1431 ,
         \D_cache/n1430 , \D_cache/n1429 , \D_cache/n1428 , \D_cache/n1427 ,
         \D_cache/n1426 , \D_cache/n1425 , \D_cache/n1424 , \D_cache/n1423 ,
         \D_cache/n1422 , \D_cache/n1421 , \D_cache/n1420 , \D_cache/n1419 ,
         \D_cache/n1418 , \D_cache/n1417 , \D_cache/n1416 , \D_cache/n1415 ,
         \D_cache/n1414 , \D_cache/n1413 , \D_cache/n1412 , \D_cache/n1411 ,
         \D_cache/n1410 , \D_cache/n1409 , \D_cache/n1408 , \D_cache/n1407 ,
         \D_cache/n1406 , \D_cache/n1405 , \D_cache/n1404 , \D_cache/n1403 ,
         \D_cache/n1402 , \D_cache/n1401 , \D_cache/n1400 , \D_cache/n1399 ,
         \D_cache/n1398 , \D_cache/n1397 , \D_cache/n1396 , \D_cache/n1395 ,
         \D_cache/n1394 , \D_cache/n1393 , \D_cache/n1392 , \D_cache/n1391 ,
         \D_cache/n1390 , \D_cache/n1389 , \D_cache/n1388 , \D_cache/n1387 ,
         \D_cache/n1386 , \D_cache/n1385 , \D_cache/n1384 , \D_cache/n1383 ,
         \D_cache/n1382 , \D_cache/n1381 , \D_cache/n1380 , \D_cache/n1379 ,
         \D_cache/n1378 , \D_cache/n1377 , \D_cache/n1376 , \D_cache/n1375 ,
         \D_cache/n1374 , \D_cache/n1373 , \D_cache/n1372 , \D_cache/n1371 ,
         \D_cache/n1370 , \D_cache/n1369 , \D_cache/n1368 , \D_cache/n1367 ,
         \D_cache/n1366 , \D_cache/n1365 , \D_cache/n1364 , \D_cache/n1363 ,
         \D_cache/n1362 , \D_cache/n1361 , \D_cache/n1360 , \D_cache/n1359 ,
         \D_cache/n1358 , \D_cache/n1357 , \D_cache/n1356 , \D_cache/n1355 ,
         \D_cache/n1354 , \D_cache/n1353 , \D_cache/n1352 , \D_cache/n1351 ,
         \D_cache/n1350 , \D_cache/n1349 , \D_cache/n1348 , \D_cache/n1347 ,
         \D_cache/n1346 , \D_cache/n1345 , \D_cache/n1344 , \D_cache/n1343 ,
         \D_cache/n1342 , \D_cache/n1341 , \D_cache/n1340 , \D_cache/n1339 ,
         \D_cache/n1338 , \D_cache/n1337 , \D_cache/n1336 , \D_cache/n1335 ,
         \D_cache/n1334 , \D_cache/n1333 , \D_cache/n1332 , \D_cache/n1331 ,
         \D_cache/n1330 , \D_cache/n1329 , \D_cache/n1328 , \D_cache/n1327 ,
         \D_cache/n1326 , \D_cache/n1325 , \D_cache/n1324 , \D_cache/n1323 ,
         \D_cache/n1322 , \D_cache/n1321 , \D_cache/n1320 , \D_cache/n1319 ,
         \D_cache/n1318 , \D_cache/n1317 , \D_cache/n1316 , \D_cache/n1315 ,
         \D_cache/n1314 , \D_cache/n1313 , \D_cache/n1312 , \D_cache/n1311 ,
         \D_cache/n1310 , \D_cache/n1309 , \D_cache/n1308 , \D_cache/n1307 ,
         \D_cache/n1306 , \D_cache/n1305 , \D_cache/n1304 , \D_cache/n1303 ,
         \D_cache/n1302 , \D_cache/n1301 , \D_cache/n1300 , \D_cache/n1299 ,
         \D_cache/n1298 , \D_cache/n1297 , \D_cache/n1296 , \D_cache/n1295 ,
         \D_cache/n1294 , \D_cache/n1293 , \D_cache/n1292 , \D_cache/n1291 ,
         \D_cache/n1290 , \D_cache/n1289 , \D_cache/n1288 , \D_cache/n1287 ,
         \D_cache/n1286 , \D_cache/n1285 , \D_cache/n1284 , \D_cache/n1283 ,
         \D_cache/n1282 , \D_cache/n1281 , \D_cache/n1280 , \D_cache/n1279 ,
         \D_cache/n1278 , \D_cache/n1277 , \D_cache/n1276 , \D_cache/n1275 ,
         \D_cache/n1274 , \D_cache/n1273 , \D_cache/n1272 , \D_cache/n1271 ,
         \D_cache/n1270 , \D_cache/n1269 , \D_cache/n1268 , \D_cache/n1267 ,
         \D_cache/n1266 , \D_cache/n1265 , \D_cache/n1264 , \D_cache/n1263 ,
         \D_cache/n1262 , \D_cache/n1261 , \D_cache/n1260 , \D_cache/n1259 ,
         \D_cache/n1258 , \D_cache/n1257 , \D_cache/n1256 , \D_cache/n1255 ,
         \D_cache/n1254 , \D_cache/n1253 , \D_cache/n1252 , \D_cache/n1251 ,
         \D_cache/n1250 , \D_cache/n1249 , \D_cache/n1248 , \D_cache/n1247 ,
         \D_cache/n1246 , \D_cache/n1245 , \D_cache/n1244 , \D_cache/n1243 ,
         \D_cache/n1242 , \D_cache/n1241 , \D_cache/n1240 , \D_cache/n1239 ,
         \D_cache/n1238 , \D_cache/n1237 , \D_cache/n1236 , \D_cache/n1235 ,
         \D_cache/n1234 , \D_cache/n1233 , \D_cache/n1232 , \D_cache/n1231 ,
         \D_cache/n1230 , \D_cache/n1229 , \D_cache/n1228 , \D_cache/n1227 ,
         \D_cache/n1226 , \D_cache/n1225 , \D_cache/n1224 , \D_cache/n1223 ,
         \D_cache/n1222 , \D_cache/n1221 , \D_cache/n1220 , \D_cache/n1219 ,
         \D_cache/n1218 , \D_cache/n1217 , \D_cache/n1216 , \D_cache/n1215 ,
         \D_cache/n1214 , \D_cache/n1213 , \D_cache/n1212 , \D_cache/n1211 ,
         \D_cache/n1210 , \D_cache/n1209 , \D_cache/n1208 , \D_cache/n1207 ,
         \D_cache/n1206 , \D_cache/n1205 , \D_cache/n1204 , \D_cache/n1203 ,
         \D_cache/n1202 , \D_cache/n1201 , \D_cache/n1200 , \D_cache/n1199 ,
         \D_cache/n1198 , \D_cache/n1197 , \D_cache/n1196 , \D_cache/n1195 ,
         \D_cache/n1194 , \D_cache/n1193 , \D_cache/n1192 , \D_cache/n1191 ,
         \D_cache/n1190 , \D_cache/n1189 , \D_cache/n1188 , \D_cache/n1187 ,
         \D_cache/n1186 , \D_cache/n1185 , \D_cache/n1184 , \D_cache/n1183 ,
         \D_cache/n1182 , \D_cache/n1181 , \D_cache/n1180 , \D_cache/n1179 ,
         \D_cache/n1178 , \D_cache/n1177 , \D_cache/n1176 , \D_cache/n1175 ,
         \D_cache/n1174 , \D_cache/n1173 , \D_cache/n1172 , \D_cache/n1171 ,
         \D_cache/n1170 , \D_cache/n1169 , \D_cache/n1168 , \D_cache/n1167 ,
         \D_cache/n1166 , \D_cache/n1165 , \D_cache/n1164 , \D_cache/n1163 ,
         \D_cache/n1162 , \D_cache/n1161 , \D_cache/n1160 , \D_cache/n1159 ,
         \D_cache/n1158 , \D_cache/n1157 , \D_cache/n1156 , \D_cache/n1155 ,
         \D_cache/n1154 , \D_cache/n1153 , \D_cache/n1152 , \D_cache/n1151 ,
         \D_cache/n1150 , \D_cache/n1149 , \D_cache/n1148 , \D_cache/n1147 ,
         \D_cache/n1146 , \D_cache/n1145 , \D_cache/n1144 , \D_cache/n1143 ,
         \D_cache/n1142 , \D_cache/n1141 , \D_cache/n1140 , \D_cache/n1139 ,
         \D_cache/n1138 , \D_cache/n1137 , \D_cache/n1136 , \D_cache/n1135 ,
         \D_cache/n1134 , \D_cache/n1133 , \D_cache/n1132 , \D_cache/n1131 ,
         \D_cache/n1130 , \D_cache/n1129 , \D_cache/n1128 , \D_cache/n1127 ,
         \D_cache/n1126 , \D_cache/n1125 , \D_cache/n1124 , \D_cache/n1123 ,
         \D_cache/n1122 , \D_cache/n1121 , \D_cache/n1120 , \D_cache/n1119 ,
         \D_cache/n1118 , \D_cache/n1117 , \D_cache/n1116 , \D_cache/n1115 ,
         \D_cache/n1114 , \D_cache/n1113 , \D_cache/n1112 , \D_cache/n1111 ,
         \D_cache/n1110 , \D_cache/n1109 , \D_cache/n1108 , \D_cache/n1107 ,
         \D_cache/n1106 , \D_cache/n1105 , \D_cache/n1104 , \D_cache/n1103 ,
         \D_cache/n1102 , \D_cache/n1101 , \D_cache/n1100 , \D_cache/n1099 ,
         \D_cache/n1098 , \D_cache/n1097 , \D_cache/n1096 , \D_cache/n1095 ,
         \D_cache/n1094 , \D_cache/n1093 , \D_cache/n1092 , \D_cache/n1091 ,
         \D_cache/n1090 , \D_cache/n1089 , \D_cache/n1088 , \D_cache/n1087 ,
         \D_cache/n1086 , \D_cache/n1085 , \D_cache/n1084 , \D_cache/n1083 ,
         \D_cache/n1082 , \D_cache/n1081 , \D_cache/n1080 , \D_cache/n1079 ,
         \D_cache/n1078 , \D_cache/n1077 , \D_cache/n1076 , \D_cache/n1075 ,
         \D_cache/n1074 , \D_cache/n1073 , \D_cache/n1072 , \D_cache/n1071 ,
         \D_cache/n1070 , \D_cache/n1069 , \D_cache/n1068 , \D_cache/n1067 ,
         \D_cache/n1066 , \D_cache/n1065 , \D_cache/n1064 , \D_cache/n1063 ,
         \D_cache/n1062 , \D_cache/n1061 , \D_cache/n1060 , \D_cache/n1059 ,
         \D_cache/n1058 , \D_cache/n1057 , \D_cache/n1056 , \D_cache/n1055 ,
         \D_cache/n1054 , \D_cache/n1053 , \D_cache/n1052 , \D_cache/n1051 ,
         \D_cache/n1050 , \D_cache/n1049 , \D_cache/n1048 , \D_cache/n1047 ,
         \D_cache/n1046 , \D_cache/n1045 , \D_cache/n1044 , \D_cache/n1043 ,
         \D_cache/n1042 , \D_cache/n1041 , \D_cache/n1040 , \D_cache/n1039 ,
         \D_cache/n1038 , \D_cache/n1037 , \D_cache/n1036 , \D_cache/n1035 ,
         \D_cache/n1034 , \D_cache/n1033 , \D_cache/n1032 , \D_cache/n1031 ,
         \D_cache/n1030 , \D_cache/n1029 , \D_cache/n1028 , \D_cache/n1027 ,
         \D_cache/n1026 , \D_cache/n1025 , \D_cache/n1024 , \D_cache/n1023 ,
         \D_cache/n1022 , \D_cache/n1021 , \D_cache/n1020 , \D_cache/n1019 ,
         \D_cache/n1018 , \D_cache/n1017 , \D_cache/n1016 , \D_cache/n1015 ,
         \D_cache/n1014 , \D_cache/n1013 , \D_cache/n1012 , \D_cache/n1011 ,
         \D_cache/n1010 , \D_cache/n1009 , \D_cache/n1008 , \D_cache/n1007 ,
         \D_cache/n1006 , \D_cache/n1005 , \D_cache/n1004 , \D_cache/n1003 ,
         \D_cache/n1002 , \D_cache/n1001 , \D_cache/n1000 , \D_cache/n999 ,
         \D_cache/n998 , \D_cache/n997 , \D_cache/n996 , \D_cache/n995 ,
         \D_cache/n994 , \D_cache/n993 , \D_cache/n992 , \D_cache/n991 ,
         \D_cache/n990 , \D_cache/n989 , \D_cache/n988 , \D_cache/n987 ,
         \D_cache/n986 , \D_cache/n985 , \D_cache/n984 , \D_cache/n983 ,
         \D_cache/n982 , \D_cache/n981 , \D_cache/n980 , \D_cache/n979 ,
         \D_cache/n978 , \D_cache/n977 , \D_cache/n976 , \D_cache/n975 ,
         \D_cache/n974 , \D_cache/n973 , \D_cache/n972 , \D_cache/n971 ,
         \D_cache/n970 , \D_cache/n969 , \D_cache/n968 , \D_cache/n967 ,
         \D_cache/n966 , \D_cache/n965 , \D_cache/n964 , \D_cache/n963 ,
         \D_cache/n962 , \D_cache/n961 , \D_cache/n960 , \D_cache/n959 ,
         \D_cache/n958 , \D_cache/n957 , \D_cache/n956 , \D_cache/n955 ,
         \D_cache/n954 , \D_cache/n953 , \D_cache/n952 , \D_cache/n951 ,
         \D_cache/n950 , \D_cache/n949 , \D_cache/n948 , \D_cache/n947 ,
         \D_cache/n946 , \D_cache/n945 , \D_cache/n944 , \D_cache/n943 ,
         \D_cache/n942 , \D_cache/n941 , \D_cache/n940 , \D_cache/n939 ,
         \D_cache/n938 , \D_cache/n937 , \D_cache/n936 , \D_cache/n935 ,
         \D_cache/n934 , \D_cache/n933 , \D_cache/n932 , \D_cache/n931 ,
         \D_cache/n930 , \D_cache/n929 , \D_cache/n928 , \D_cache/n927 ,
         \D_cache/n926 , \D_cache/n925 , \D_cache/n924 , \D_cache/n923 ,
         \D_cache/n922 , \D_cache/n921 , \D_cache/n920 , \D_cache/n919 ,
         \D_cache/n918 , \D_cache/n917 , \D_cache/n916 , \D_cache/n915 ,
         \D_cache/n914 , \D_cache/n913 , \D_cache/n912 , \D_cache/n911 ,
         \D_cache/n910 , \D_cache/n909 , \D_cache/n908 , \D_cache/n907 ,
         \D_cache/n906 , \D_cache/n905 , \D_cache/n904 , \D_cache/n903 ,
         \D_cache/n902 , \D_cache/n901 , \D_cache/n900 , \D_cache/n899 ,
         \D_cache/n898 , \D_cache/n897 , \D_cache/n896 , \D_cache/n895 ,
         \D_cache/n894 , \D_cache/n893 , \D_cache/n892 , \D_cache/n891 ,
         \D_cache/n890 , \D_cache/n889 , \D_cache/n888 , \D_cache/n887 ,
         \D_cache/n886 , \D_cache/n885 , \D_cache/n884 , \D_cache/n883 ,
         \D_cache/n882 , \D_cache/n881 , \D_cache/n880 , \D_cache/n879 ,
         \D_cache/n878 , \D_cache/n877 , \D_cache/n876 , \D_cache/n875 ,
         \D_cache/n874 , \D_cache/n873 , \D_cache/n872 , \D_cache/n871 ,
         \D_cache/n870 , \D_cache/n869 , \D_cache/n868 , \D_cache/n867 ,
         \D_cache/n866 , \D_cache/n865 , \D_cache/n864 , \D_cache/n863 ,
         \D_cache/n862 , \D_cache/n861 , \D_cache/n860 , \D_cache/n859 ,
         \D_cache/n858 , \D_cache/n857 , \D_cache/n856 , \D_cache/n855 ,
         \D_cache/n854 , \D_cache/n853 , \D_cache/n852 , \D_cache/n851 ,
         \D_cache/n850 , \D_cache/n849 , \D_cache/n848 , \D_cache/n847 ,
         \D_cache/n846 , \D_cache/n845 , \D_cache/n844 , \D_cache/n843 ,
         \D_cache/n842 , \D_cache/n841 , \D_cache/n840 , \D_cache/n839 ,
         \D_cache/n838 , \D_cache/n837 , \D_cache/n836 , \D_cache/n835 ,
         \D_cache/n834 , \D_cache/n833 , \D_cache/n832 , \D_cache/n831 ,
         \D_cache/n830 , \D_cache/n829 , \D_cache/n828 , \D_cache/n827 ,
         \D_cache/n826 , \D_cache/n825 , \D_cache/n824 , \D_cache/n823 ,
         \D_cache/n822 , \D_cache/n821 , \D_cache/n820 , \D_cache/n819 ,
         \D_cache/n818 , \D_cache/n817 , \D_cache/n816 , \D_cache/n815 ,
         \D_cache/n814 , \D_cache/n813 , \D_cache/n812 , \D_cache/n811 ,
         \D_cache/n810 , \D_cache/n809 , \D_cache/n808 , \D_cache/n807 ,
         \D_cache/n806 , \D_cache/n805 , \D_cache/n804 , \D_cache/n803 ,
         \D_cache/n802 , \D_cache/n801 , \D_cache/n800 , \D_cache/n799 ,
         \D_cache/n798 , \D_cache/n797 , \D_cache/n796 , \D_cache/n795 ,
         \D_cache/n794 , \D_cache/n793 , \D_cache/n792 , \D_cache/n791 ,
         \D_cache/n790 , \D_cache/n789 , \D_cache/n788 , \D_cache/n787 ,
         \D_cache/n786 , \D_cache/n785 , \D_cache/n784 , \D_cache/n783 ,
         \D_cache/n782 , \D_cache/n781 , \D_cache/n780 , \D_cache/n779 ,
         \D_cache/n778 , \D_cache/n777 , \D_cache/n776 , \D_cache/n775 ,
         \D_cache/n774 , \D_cache/n773 , \D_cache/n772 , \D_cache/n771 ,
         \D_cache/n770 , \D_cache/n769 , \D_cache/n768 , \D_cache/n767 ,
         \D_cache/n766 , \D_cache/n765 , \D_cache/n764 , \D_cache/n763 ,
         \D_cache/n762 , \D_cache/n761 , \D_cache/n760 , \D_cache/n759 ,
         \D_cache/n758 , \D_cache/n757 , \D_cache/n756 , \D_cache/n755 ,
         \D_cache/n754 , \D_cache/n753 , \D_cache/n752 , \D_cache/n751 ,
         \D_cache/n750 , \D_cache/n749 , \D_cache/n748 , \D_cache/n747 ,
         \D_cache/n746 , \D_cache/n745 , \D_cache/n744 , \D_cache/n743 ,
         \D_cache/n742 , \D_cache/n741 , \D_cache/n740 , \D_cache/n739 ,
         \D_cache/n738 , \D_cache/n737 , \D_cache/n736 , \D_cache/n735 ,
         \D_cache/n734 , \D_cache/n733 , \D_cache/n732 , \D_cache/n731 ,
         \D_cache/n730 , \D_cache/n729 , \D_cache/n728 , \D_cache/n727 ,
         \D_cache/n726 , \D_cache/n725 , \D_cache/n724 , \D_cache/n723 ,
         \D_cache/n722 , \D_cache/n721 , \D_cache/n720 , \D_cache/n719 ,
         \D_cache/n718 , \D_cache/n717 , \D_cache/n716 , \D_cache/n715 ,
         \D_cache/n714 , \D_cache/n713 , \D_cache/n712 , \D_cache/n711 ,
         \D_cache/n710 , \D_cache/n709 , \D_cache/n708 , \D_cache/n707 ,
         \D_cache/n706 , \D_cache/n705 , \D_cache/n704 , \D_cache/n703 ,
         \D_cache/n702 , \D_cache/n701 , \D_cache/n700 , \D_cache/n699 ,
         \D_cache/n698 , \D_cache/n697 , \D_cache/n696 , \D_cache/n695 ,
         \D_cache/n694 , \D_cache/n693 , \D_cache/n692 , \D_cache/n691 ,
         \D_cache/n690 , \D_cache/n689 , \D_cache/n688 , \D_cache/n687 ,
         \D_cache/n686 , \D_cache/n685 , \D_cache/n684 , \D_cache/n683 ,
         \D_cache/n682 , \D_cache/n681 , \D_cache/n680 , \D_cache/n679 ,
         \D_cache/n678 , \D_cache/n677 , \D_cache/n676 , \D_cache/n675 ,
         \D_cache/n674 , \D_cache/n673 , \D_cache/n672 , \D_cache/n671 ,
         \D_cache/n670 , \D_cache/n669 , \D_cache/n668 , \D_cache/n667 ,
         \D_cache/n666 , \D_cache/n665 , \D_cache/n664 , \D_cache/n663 ,
         \D_cache/n662 , \D_cache/n661 , \D_cache/n660 , \D_cache/n659 ,
         \D_cache/n658 , \D_cache/n657 , \D_cache/n656 , \D_cache/n655 ,
         \D_cache/n654 , \D_cache/n653 , \D_cache/n652 , \D_cache/n651 ,
         \D_cache/n650 , \D_cache/n649 , \D_cache/n648 , \D_cache/n647 ,
         \D_cache/n646 , \D_cache/n645 , \D_cache/n644 , \D_cache/n643 ,
         \D_cache/n642 , \D_cache/n641 , \D_cache/n640 , \D_cache/n639 ,
         \D_cache/n638 , \D_cache/n637 , \D_cache/n636 , \D_cache/n635 ,
         \D_cache/n634 , \D_cache/n633 , \D_cache/n632 , \D_cache/n631 ,
         \D_cache/n630 , \D_cache/n629 , \D_cache/n628 , \D_cache/n627 ,
         \D_cache/n626 , \D_cache/n625 , \D_cache/n624 , \D_cache/n623 ,
         \D_cache/n622 , \D_cache/n621 , \D_cache/n620 , \D_cache/n619 ,
         \D_cache/n618 , \D_cache/n617 , \D_cache/n616 , \D_cache/n615 ,
         \D_cache/n614 , \D_cache/n613 , \D_cache/n612 , \D_cache/n611 ,
         \D_cache/n610 , \D_cache/n609 , \D_cache/n608 , \D_cache/n607 ,
         \D_cache/n606 , \D_cache/n605 , \D_cache/n604 , \D_cache/n603 ,
         \D_cache/n602 , \D_cache/n601 , \D_cache/n600 , \D_cache/n599 ,
         \D_cache/n598 , \D_cache/n597 , \D_cache/n596 , \D_cache/n595 ,
         \D_cache/n594 , \D_cache/n593 , \D_cache/n592 , \D_cache/n591 ,
         \D_cache/n590 , \D_cache/n589 , \D_cache/n588 , \D_cache/n587 ,
         \D_cache/n586 , \D_cache/n585 , \D_cache/n584 , \D_cache/n583 ,
         \D_cache/n582 , \D_cache/n581 , \D_cache/n580 , \D_cache/n579 ,
         \D_cache/n578 , \D_cache/n577 , \D_cache/n576 , \D_cache/n575 ,
         \D_cache/n574 , \D_cache/n573 , \D_cache/n572 , \D_cache/n571 ,
         \D_cache/n570 , \D_cache/n569 , \D_cache/n568 , \D_cache/n567 ,
         \D_cache/n566 , \D_cache/n565 , \D_cache/n564 , \D_cache/n563 ,
         \D_cache/n562 , \D_cache/n561 , \D_cache/n560 , \D_cache/n559 ,
         \D_cache/n558 , \D_cache/n557 , \D_cache/n556 , \D_cache/n555 ,
         \D_cache/n554 , \D_cache/n553 , \D_cache/n552 , \D_cache/n551 ,
         \D_cache/n550 , \D_cache/n542 , \D_cache/n541 , \D_cache/n540 ,
         \D_cache/n539 , \D_cache/n538 , \D_cache/n537 , \D_cache/n536 ,
         \D_cache/n535 , \D_cache/n534 , \D_cache/n533 , \D_cache/n532 ,
         \D_cache/n531 , \D_cache/n530 , \D_cache/n529 , \D_cache/n528 ,
         \D_cache/n527 , \D_cache/n526 , \D_cache/n525 , \D_cache/n523 ,
         \D_cache/n522 , \D_cache/n520 , \D_cache/n519 , \D_cache/n518 ,
         \D_cache/n517 , \D_cache/n516 , \D_cache/n515 , \D_cache/n514 ,
         \D_cache/n513 , \D_cache/n512 , \D_cache/n511 , \D_cache/n510 ,
         \D_cache/n509 , \D_cache/n508 , \D_cache/n507 , \D_cache/n506 ,
         \D_cache/n505 , \D_cache/n504 , \D_cache/n503 , \D_cache/n502 ,
         \D_cache/n501 , \D_cache/n500 , \D_cache/n499 , \D_cache/n498 ,
         \D_cache/n497 , \D_cache/n496 , \D_cache/n495 , \D_cache/n494 ,
         \D_cache/n493 , \D_cache/n492 , \D_cache/n491 , \D_cache/n490 ,
         \D_cache/n489 , \D_cache/n488 , \D_cache/n487 , \D_cache/n486 ,
         \D_cache/n485 , \D_cache/n484 , \D_cache/n483 , \D_cache/n482 ,
         \D_cache/n481 , \D_cache/n480 , \D_cache/n479 , \D_cache/n478 ,
         \D_cache/n477 , \D_cache/n476 , \D_cache/n475 , \D_cache/n474 ,
         \D_cache/n473 , \D_cache/n472 , \D_cache/n471 , \D_cache/n470 ,
         \D_cache/n469 , \D_cache/n468 , \D_cache/n467 , \D_cache/n466 ,
         \D_cache/n465 , \D_cache/n464 , \D_cache/n463 , \D_cache/n462 ,
         \D_cache/n461 , \D_cache/n460 , \D_cache/n459 , \D_cache/n458 ,
         \D_cache/n457 , \D_cache/n456 , \D_cache/n455 , \D_cache/n454 ,
         \D_cache/n453 , \D_cache/n452 , \D_cache/n451 , \D_cache/n450 ,
         \D_cache/n449 , \D_cache/n448 , \D_cache/n447 , \D_cache/n446 ,
         \D_cache/n445 , \D_cache/n444 , \D_cache/n443 , \D_cache/n442 ,
         \D_cache/n441 , \D_cache/n440 , \D_cache/n439 , \D_cache/n438 ,
         \D_cache/n437 , \D_cache/n436 , \D_cache/n435 , \D_cache/n434 ,
         \D_cache/n433 , \D_cache/n432 , \D_cache/n431 , \D_cache/n430 ,
         \D_cache/n429 , \D_cache/n428 , \D_cache/n427 , \D_cache/n426 ,
         \D_cache/n425 , \D_cache/n424 , \D_cache/n423 , \D_cache/n422 ,
         \D_cache/n421 , \D_cache/n420 , \D_cache/n419 , \D_cache/n418 ,
         \D_cache/n417 , \D_cache/n416 , \D_cache/n415 , \D_cache/n414 ,
         \D_cache/n413 , \D_cache/n412 , \D_cache/n411 , \D_cache/n410 ,
         \D_cache/n409 , \D_cache/n408 , \D_cache/n407 , \D_cache/n406 ,
         \D_cache/n405 , \D_cache/n404 , \D_cache/n403 , \D_cache/n402 ,
         \D_cache/n401 , \D_cache/n400 , \D_cache/n399 , \D_cache/n398 ,
         \D_cache/n397 , \D_cache/n396 , \D_cache/n395 , \D_cache/n394 ,
         \D_cache/n393 , \D_cache/n392 , \D_cache/n391 , \D_cache/n390 ,
         \D_cache/n389 , \D_cache/n388 , \D_cache/n387 , \D_cache/n386 ,
         \D_cache/n385 , \D_cache/n384 , \D_cache/n383 , \D_cache/n382 ,
         \D_cache/n381 , \D_cache/n380 , \D_cache/n379 , \D_cache/n378 ,
         \D_cache/n377 , \D_cache/n376 , \D_cache/n375 , \D_cache/n374 ,
         \D_cache/n373 , \D_cache/n372 , \D_cache/n371 , \D_cache/n370 ,
         \D_cache/n369 , \D_cache/n368 , \D_cache/n367 , \D_cache/n366 ,
         \D_cache/n365 , \D_cache/n364 , \D_cache/n363 , \D_cache/n362 ,
         \D_cache/n361 , \D_cache/n360 , \D_cache/n359 , \D_cache/n358 ,
         \D_cache/n357 , \D_cache/n356 , \D_cache/n355 , \D_cache/n354 ,
         \D_cache/n353 , \D_cache/n352 , \D_cache/n351 , \D_cache/n350 ,
         \D_cache/n349 , \D_cache/n348 , \D_cache/n347 , \D_cache/n346 ,
         \D_cache/n345 , \D_cache/n344 , \D_cache/n343 , \D_cache/n342 ,
         \D_cache/n341 , \D_cache/n340 , \D_cache/n339 , \D_cache/n338 ,
         \D_cache/n337 , \D_cache/n336 , \D_cache/n335 , \D_cache/n334 ,
         \D_cache/n333 , \D_cache/n332 , \D_cache/n331 , \D_cache/n330 ,
         \D_cache/n329 , \D_cache/n328 , \D_cache/n327 , \D_cache/n326 ,
         \D_cache/n325 , \D_cache/n324 , \D_cache/n323 , \D_cache/n322 ,
         \D_cache/n321 , \D_cache/n320 , \D_cache/n319 , \D_cache/n318 ,
         \D_cache/n317 , \D_cache/n316 , \D_cache/n315 , \D_cache/n314 ,
         \D_cache/n313 , \D_cache/n312 , \D_cache/n311 , \D_cache/n310 ,
         \D_cache/n309 , \D_cache/n308 , \D_cache/n307 , \D_cache/n306 ,
         \D_cache/n305 , \D_cache/n304 , \D_cache/n303 , \D_cache/n302 ,
         \D_cache/n301 , \D_cache/n300 , \D_cache/n299 , \D_cache/n298 ,
         \D_cache/n297 , \D_cache/n296 , \D_cache/n295 , \D_cache/n294 ,
         \D_cache/n293 , \D_cache/n292 , \D_cache/n291 , \D_cache/n290 ,
         \D_cache/n289 , \D_cache/n288 , \D_cache/n287 , \D_cache/n286 ,
         \D_cache/n285 , \D_cache/n284 , \D_cache/n283 , \D_cache/n282 ,
         \D_cache/n281 , \D_cache/n280 , \D_cache/n279 , \D_cache/n278 ,
         \D_cache/n277 , \D_cache/n276 , \D_cache/n275 , \D_cache/n274 ,
         \D_cache/n273 , \D_cache/n272 , \D_cache/n271 , \D_cache/n270 ,
         \D_cache/n269 , \D_cache/n268 , \D_cache/n267 , \D_cache/n266 ,
         \D_cache/n265 , \D_cache/n264 , \D_cache/n263 , \D_cache/n262 ,
         \D_cache/n261 , \D_cache/n260 , \D_cache/n259 , \D_cache/n258 ,
         \D_cache/n257 , \D_cache/n256 , \D_cache/n255 , \D_cache/n254 ,
         \D_cache/n253 , \D_cache/n252 , \D_cache/n251 , \D_cache/n250 ,
         \D_cache/n249 , \D_cache/n248 , \D_cache/n247 , \D_cache/n246 ,
         \D_cache/n245 , \D_cache/n244 , \D_cache/n243 , \D_cache/n242 ,
         \D_cache/n241 , \D_cache/n240 , \D_cache/n239 , \D_cache/n238 ,
         \D_cache/n237 , \D_cache/n236 , \D_cache/n235 , \D_cache/n234 ,
         \D_cache/n233 , \D_cache/n232 , \D_cache/n231 , \D_cache/n230 ,
         \D_cache/n229 , \D_cache/n228 , \D_cache/n227 , \D_cache/n226 ,
         \D_cache/n225 , \D_cache/n224 , \D_cache/n223 , \D_cache/n222 ,
         \D_cache/n218 , \D_cache/n217 , \D_cache/n216 , \D_cache/n215 ,
         \D_cache/n214 , \D_cache/n213 , \D_cache/n212 , \D_cache/n211 ,
         \D_cache/n210 , \D_cache/n209 , \D_cache/n208 , \D_cache/n207 ,
         \D_cache/n206 , \D_cache/n205 , \D_cache/n204 , \D_cache/n203 ,
         \D_cache/n202 , \D_cache/n201 , \D_cache/n200 , \D_cache/n199 ,
         \D_cache/n198 , \D_cache/n197 , \D_cache/n196 , \D_cache/n195 ,
         \D_cache/n194 , \D_cache/n193 , \D_cache/n192 , \D_cache/n191 ,
         \D_cache/n190 , \D_cache/n189 , \D_cache/n188 , \D_cache/n187 ,
         \D_cache/n186 , \D_cache/n185 , \D_cache/n184 , \D_cache/n183 ,
         \D_cache/n182 , \D_cache/n181 , \D_cache/n180 , \D_cache/n179 ,
         \D_cache/n178 , \D_cache/n177 , \D_cache/n176 , \D_cache/n175 ,
         \D_cache/n174 , \D_cache/n173 , \D_cache/n172 , \D_cache/n171 ,
         \D_cache/n170 , \D_cache/n169 , \D_cache/n166 , \D_cache/n165 ,
         \D_cache/n164 , \D_cache/N184 , \D_cache/N183 , \D_cache/N182 ,
         \D_cache/N181 , \D_cache/N180 , \D_cache/N179 , \D_cache/N178 ,
         \D_cache/N177 , \D_cache/N176 , \D_cache/N175 , \D_cache/N174 ,
         \D_cache/N173 , \D_cache/N172 , \D_cache/N171 , \D_cache/N170 ,
         \D_cache/N169 , \D_cache/N168 , \D_cache/N167 , \D_cache/N166 ,
         \D_cache/N165 , \D_cache/N164 , \D_cache/N163 , \D_cache/N162 ,
         \D_cache/N161 , \D_cache/N160 , \D_cache/N159 , \D_cache/N158 ,
         \D_cache/N157 , \D_cache/N156 , \D_cache/N155 , \D_cache/N154 ,
         \D_cache/N153 , \D_cache/N152 , \D_cache/N151 , \D_cache/N150 ,
         \D_cache/N149 , \D_cache/N148 , \D_cache/N147 , \D_cache/N146 ,
         \D_cache/N145 , \D_cache/N144 , \D_cache/N143 , \D_cache/N142 ,
         \D_cache/N141 , \D_cache/N140 , \D_cache/N139 , \D_cache/N138 ,
         \D_cache/N137 , \D_cache/N136 , \D_cache/N135 , \D_cache/N134 ,
         \D_cache/N133 , \D_cache/N132 , \D_cache/N131 , \D_cache/N130 ,
         \D_cache/N129 , \D_cache/N128 , \D_cache/N127 , \D_cache/N126 ,
         \D_cache/N125 , \D_cache/N124 , \D_cache/N123 , \D_cache/N122 ,
         \D_cache/N121 , \D_cache/N120 , \D_cache/N119 , \D_cache/N118 ,
         \D_cache/N117 , \D_cache/N116 , \D_cache/N115 , \D_cache/N114 ,
         \D_cache/N113 , \D_cache/N112 , \D_cache/N111 , \D_cache/N110 ,
         \D_cache/N109 , \D_cache/N108 , \D_cache/N107 , \D_cache/N106 ,
         \D_cache/N105 , \D_cache/N104 , \D_cache/N103 , \D_cache/N102 ,
         \D_cache/N101 , \D_cache/N100 , \D_cache/N99 , \D_cache/N98 ,
         \D_cache/N97 , \D_cache/N96 , \D_cache/N95 , \D_cache/N94 ,
         \D_cache/N93 , \D_cache/N92 , \D_cache/N91 , \D_cache/N90 ,
         \D_cache/N89 , \D_cache/N88 , \D_cache/N87 , \D_cache/N86 ,
         \D_cache/N85 , \D_cache/N84 , \D_cache/N83 , \D_cache/N82 ,
         \D_cache/N81 , \D_cache/N80 , \D_cache/N79 , \D_cache/N78 ,
         \D_cache/N77 , \D_cache/N76 , \D_cache/N75 , \D_cache/N74 ,
         \D_cache/N73 , \D_cache/N72 , \D_cache/N71 , \D_cache/N70 ,
         \D_cache/N69 , \D_cache/N68 , \D_cache/N67 , \D_cache/N66 ,
         \D_cache/N65 , \D_cache/N64 , \D_cache/N63 , \D_cache/N62 ,
         \D_cache/N61 , \D_cache/N60 , \D_cache/N59 , \D_cache/N58 ,
         \D_cache/N57 , \D_cache/N56 , \D_cache/N55 , \D_cache/N54 ,
         \D_cache/N53 , \D_cache/N52 , \D_cache/N51 , \D_cache/N50 ,
         \D_cache/N49 , \D_cache/N48 , \D_cache/N47 , \D_cache/N46 ,
         \D_cache/N45 , \D_cache/N44 , \D_cache/N43 , \D_cache/N42 ,
         \D_cache/N41 , \D_cache/N40 , \D_cache/N39 , \D_cache/N38 ,
         \D_cache/N37 , \D_cache/N36 , \D_cache/N35 , \D_cache/N34 ,
         \D_cache/N33 , \D_cache/N32 , \D_cache/N31 , \D_cache/N30 ,
         \D_cache/cache[7][0] , \D_cache/cache[7][1] , \D_cache/cache[7][2] ,
         \D_cache/cache[7][3] , \D_cache/cache[7][4] , \D_cache/cache[7][5] ,
         \D_cache/cache[7][6] , \D_cache/cache[7][7] , \D_cache/cache[7][8] ,
         \D_cache/cache[7][9] , \D_cache/cache[7][10] , \D_cache/cache[7][11] ,
         \D_cache/cache[7][12] , \D_cache/cache[7][13] ,
         \D_cache/cache[7][14] , \D_cache/cache[7][15] ,
         \D_cache/cache[7][16] , \D_cache/cache[7][17] ,
         \D_cache/cache[7][18] , \D_cache/cache[7][19] ,
         \D_cache/cache[7][20] , \D_cache/cache[7][21] ,
         \D_cache/cache[7][22] , \D_cache/cache[7][23] ,
         \D_cache/cache[7][24] , \D_cache/cache[7][25] ,
         \D_cache/cache[7][26] , \D_cache/cache[7][27] ,
         \D_cache/cache[7][28] , \D_cache/cache[7][29] ,
         \D_cache/cache[7][30] , \D_cache/cache[7][31] ,
         \D_cache/cache[7][32] , \D_cache/cache[7][33] ,
         \D_cache/cache[7][34] , \D_cache/cache[7][35] ,
         \D_cache/cache[7][36] , \D_cache/cache[7][37] ,
         \D_cache/cache[7][38] , \D_cache/cache[7][39] ,
         \D_cache/cache[7][40] , \D_cache/cache[7][41] ,
         \D_cache/cache[7][42] , \D_cache/cache[7][43] ,
         \D_cache/cache[7][44] , \D_cache/cache[7][45] ,
         \D_cache/cache[7][46] , \D_cache/cache[7][47] ,
         \D_cache/cache[7][48] , \D_cache/cache[7][49] ,
         \D_cache/cache[7][50] , \D_cache/cache[7][51] ,
         \D_cache/cache[7][52] , \D_cache/cache[7][53] ,
         \D_cache/cache[7][54] , \D_cache/cache[7][55] ,
         \D_cache/cache[7][56] , \D_cache/cache[7][57] ,
         \D_cache/cache[7][58] , \D_cache/cache[7][59] ,
         \D_cache/cache[7][60] , \D_cache/cache[7][61] ,
         \D_cache/cache[7][62] , \D_cache/cache[7][63] ,
         \D_cache/cache[7][64] , \D_cache/cache[7][65] ,
         \D_cache/cache[7][66] , \D_cache/cache[7][67] ,
         \D_cache/cache[7][68] , \D_cache/cache[7][69] ,
         \D_cache/cache[7][70] , \D_cache/cache[7][71] ,
         \D_cache/cache[7][72] , \D_cache/cache[7][73] ,
         \D_cache/cache[7][74] , \D_cache/cache[7][75] ,
         \D_cache/cache[7][76] , \D_cache/cache[7][77] ,
         \D_cache/cache[7][78] , \D_cache/cache[7][79] ,
         \D_cache/cache[7][80] , \D_cache/cache[7][81] ,
         \D_cache/cache[7][82] , \D_cache/cache[7][83] ,
         \D_cache/cache[7][84] , \D_cache/cache[7][85] ,
         \D_cache/cache[7][86] , \D_cache/cache[7][87] ,
         \D_cache/cache[7][88] , \D_cache/cache[7][89] ,
         \D_cache/cache[7][90] , \D_cache/cache[7][91] ,
         \D_cache/cache[7][92] , \D_cache/cache[7][93] ,
         \D_cache/cache[7][94] , \D_cache/cache[7][95] ,
         \D_cache/cache[7][96] , \D_cache/cache[7][97] ,
         \D_cache/cache[7][98] , \D_cache/cache[7][99] ,
         \D_cache/cache[7][100] , \D_cache/cache[7][101] ,
         \D_cache/cache[7][102] , \D_cache/cache[7][103] ,
         \D_cache/cache[7][104] , \D_cache/cache[7][105] ,
         \D_cache/cache[7][106] , \D_cache/cache[7][107] ,
         \D_cache/cache[7][108] , \D_cache/cache[7][109] ,
         \D_cache/cache[7][110] , \D_cache/cache[7][111] ,
         \D_cache/cache[7][112] , \D_cache/cache[7][113] ,
         \D_cache/cache[7][114] , \D_cache/cache[7][115] ,
         \D_cache/cache[7][116] , \D_cache/cache[7][117] ,
         \D_cache/cache[7][118] , \D_cache/cache[7][119] ,
         \D_cache/cache[7][120] , \D_cache/cache[7][121] ,
         \D_cache/cache[7][122] , \D_cache/cache[7][123] ,
         \D_cache/cache[7][124] , \D_cache/cache[7][125] ,
         \D_cache/cache[7][126] , \D_cache/cache[7][127] ,
         \D_cache/cache[7][128] , \D_cache/cache[7][129] ,
         \D_cache/cache[7][130] , \D_cache/cache[7][131] ,
         \D_cache/cache[7][132] , \D_cache/cache[7][133] ,
         \D_cache/cache[7][134] , \D_cache/cache[7][135] ,
         \D_cache/cache[7][136] , \D_cache/cache[7][137] ,
         \D_cache/cache[7][138] , \D_cache/cache[7][139] ,
         \D_cache/cache[7][140] , \D_cache/cache[7][141] ,
         \D_cache/cache[7][142] , \D_cache/cache[7][143] ,
         \D_cache/cache[7][144] , \D_cache/cache[7][145] ,
         \D_cache/cache[7][146] , \D_cache/cache[7][147] ,
         \D_cache/cache[7][148] , \D_cache/cache[7][149] ,
         \D_cache/cache[7][150] , \D_cache/cache[7][151] ,
         \D_cache/cache[7][152] , \D_cache/cache[7][153] ,
         \D_cache/cache[7][154] , \D_cache/cache[6][0] , \D_cache/cache[6][1] ,
         \D_cache/cache[6][2] , \D_cache/cache[6][3] , \D_cache/cache[6][4] ,
         \D_cache/cache[6][5] , \D_cache/cache[6][6] , \D_cache/cache[6][7] ,
         \D_cache/cache[6][8] , \D_cache/cache[6][9] , \D_cache/cache[6][10] ,
         \D_cache/cache[6][11] , \D_cache/cache[6][12] ,
         \D_cache/cache[6][13] , \D_cache/cache[6][14] ,
         \D_cache/cache[6][15] , \D_cache/cache[6][16] ,
         \D_cache/cache[6][17] , \D_cache/cache[6][18] ,
         \D_cache/cache[6][19] , \D_cache/cache[6][20] ,
         \D_cache/cache[6][21] , \D_cache/cache[6][22] ,
         \D_cache/cache[6][23] , \D_cache/cache[6][24] ,
         \D_cache/cache[6][25] , \D_cache/cache[6][26] ,
         \D_cache/cache[6][27] , \D_cache/cache[6][28] ,
         \D_cache/cache[6][29] , \D_cache/cache[6][30] ,
         \D_cache/cache[6][31] , \D_cache/cache[6][32] ,
         \D_cache/cache[6][33] , \D_cache/cache[6][34] ,
         \D_cache/cache[6][35] , \D_cache/cache[6][36] ,
         \D_cache/cache[6][37] , \D_cache/cache[6][38] ,
         \D_cache/cache[6][39] , \D_cache/cache[6][40] ,
         \D_cache/cache[6][41] , \D_cache/cache[6][42] ,
         \D_cache/cache[6][43] , \D_cache/cache[6][44] ,
         \D_cache/cache[6][45] , \D_cache/cache[6][46] ,
         \D_cache/cache[6][47] , \D_cache/cache[6][48] ,
         \D_cache/cache[6][49] , \D_cache/cache[6][50] ,
         \D_cache/cache[6][51] , \D_cache/cache[6][52] ,
         \D_cache/cache[6][53] , \D_cache/cache[6][54] ,
         \D_cache/cache[6][55] , \D_cache/cache[6][56] ,
         \D_cache/cache[6][57] , \D_cache/cache[6][58] ,
         \D_cache/cache[6][59] , \D_cache/cache[6][60] ,
         \D_cache/cache[6][61] , \D_cache/cache[6][62] ,
         \D_cache/cache[6][63] , \D_cache/cache[6][64] ,
         \D_cache/cache[6][65] , \D_cache/cache[6][66] ,
         \D_cache/cache[6][67] , \D_cache/cache[6][68] ,
         \D_cache/cache[6][69] , \D_cache/cache[6][70] ,
         \D_cache/cache[6][71] , \D_cache/cache[6][72] ,
         \D_cache/cache[6][73] , \D_cache/cache[6][74] ,
         \D_cache/cache[6][75] , \D_cache/cache[6][76] ,
         \D_cache/cache[6][77] , \D_cache/cache[6][78] ,
         \D_cache/cache[6][79] , \D_cache/cache[6][80] ,
         \D_cache/cache[6][81] , \D_cache/cache[6][82] ,
         \D_cache/cache[6][83] , \D_cache/cache[6][84] ,
         \D_cache/cache[6][85] , \D_cache/cache[6][86] ,
         \D_cache/cache[6][87] , \D_cache/cache[6][88] ,
         \D_cache/cache[6][89] , \D_cache/cache[6][90] ,
         \D_cache/cache[6][91] , \D_cache/cache[6][92] ,
         \D_cache/cache[6][93] , \D_cache/cache[6][94] ,
         \D_cache/cache[6][95] , \D_cache/cache[6][96] ,
         \D_cache/cache[6][97] , \D_cache/cache[6][98] ,
         \D_cache/cache[6][99] , \D_cache/cache[6][100] ,
         \D_cache/cache[6][101] , \D_cache/cache[6][102] ,
         \D_cache/cache[6][103] , \D_cache/cache[6][104] ,
         \D_cache/cache[6][105] , \D_cache/cache[6][106] ,
         \D_cache/cache[6][107] , \D_cache/cache[6][108] ,
         \D_cache/cache[6][109] , \D_cache/cache[6][110] ,
         \D_cache/cache[6][111] , \D_cache/cache[6][112] ,
         \D_cache/cache[6][113] , \D_cache/cache[6][114] ,
         \D_cache/cache[6][115] , \D_cache/cache[6][116] ,
         \D_cache/cache[6][117] , \D_cache/cache[6][118] ,
         \D_cache/cache[6][119] , \D_cache/cache[6][120] ,
         \D_cache/cache[6][121] , \D_cache/cache[6][122] ,
         \D_cache/cache[6][123] , \D_cache/cache[6][124] ,
         \D_cache/cache[6][125] , \D_cache/cache[6][126] ,
         \D_cache/cache[6][127] , \D_cache/cache[6][128] ,
         \D_cache/cache[6][129] , \D_cache/cache[6][130] ,
         \D_cache/cache[6][131] , \D_cache/cache[6][132] ,
         \D_cache/cache[6][133] , \D_cache/cache[6][134] ,
         \D_cache/cache[6][135] , \D_cache/cache[6][136] ,
         \D_cache/cache[6][137] , \D_cache/cache[6][138] ,
         \D_cache/cache[6][139] , \D_cache/cache[6][140] ,
         \D_cache/cache[6][141] , \D_cache/cache[6][142] ,
         \D_cache/cache[6][143] , \D_cache/cache[6][144] ,
         \D_cache/cache[6][145] , \D_cache/cache[6][146] ,
         \D_cache/cache[6][147] , \D_cache/cache[6][148] ,
         \D_cache/cache[6][149] , \D_cache/cache[6][150] ,
         \D_cache/cache[6][151] , \D_cache/cache[6][152] ,
         \D_cache/cache[6][153] , \D_cache/cache[6][154] ,
         \D_cache/cache[5][0] , \D_cache/cache[5][1] , \D_cache/cache[5][2] ,
         \D_cache/cache[5][3] , \D_cache/cache[5][4] , \D_cache/cache[5][5] ,
         \D_cache/cache[5][6] , \D_cache/cache[5][7] , \D_cache/cache[5][8] ,
         \D_cache/cache[5][9] , \D_cache/cache[5][10] , \D_cache/cache[5][11] ,
         \D_cache/cache[5][12] , \D_cache/cache[5][13] ,
         \D_cache/cache[5][14] , \D_cache/cache[5][15] ,
         \D_cache/cache[5][16] , \D_cache/cache[5][17] ,
         \D_cache/cache[5][18] , \D_cache/cache[5][19] ,
         \D_cache/cache[5][20] , \D_cache/cache[5][21] ,
         \D_cache/cache[5][22] , \D_cache/cache[5][23] ,
         \D_cache/cache[5][24] , \D_cache/cache[5][25] ,
         \D_cache/cache[5][26] , \D_cache/cache[5][27] ,
         \D_cache/cache[5][28] , \D_cache/cache[5][29] ,
         \D_cache/cache[5][30] , \D_cache/cache[5][31] ,
         \D_cache/cache[5][32] , \D_cache/cache[5][33] ,
         \D_cache/cache[5][34] , \D_cache/cache[5][35] ,
         \D_cache/cache[5][36] , \D_cache/cache[5][37] ,
         \D_cache/cache[5][38] , \D_cache/cache[5][39] ,
         \D_cache/cache[5][40] , \D_cache/cache[5][41] ,
         \D_cache/cache[5][42] , \D_cache/cache[5][43] ,
         \D_cache/cache[5][44] , \D_cache/cache[5][45] ,
         \D_cache/cache[5][46] , \D_cache/cache[5][47] ,
         \D_cache/cache[5][48] , \D_cache/cache[5][49] ,
         \D_cache/cache[5][50] , \D_cache/cache[5][51] ,
         \D_cache/cache[5][52] , \D_cache/cache[5][53] ,
         \D_cache/cache[5][54] , \D_cache/cache[5][55] ,
         \D_cache/cache[5][56] , \D_cache/cache[5][57] ,
         \D_cache/cache[5][58] , \D_cache/cache[5][59] ,
         \D_cache/cache[5][60] , \D_cache/cache[5][61] ,
         \D_cache/cache[5][62] , \D_cache/cache[5][63] ,
         \D_cache/cache[5][64] , \D_cache/cache[5][65] ,
         \D_cache/cache[5][66] , \D_cache/cache[5][67] ,
         \D_cache/cache[5][68] , \D_cache/cache[5][69] ,
         \D_cache/cache[5][70] , \D_cache/cache[5][71] ,
         \D_cache/cache[5][72] , \D_cache/cache[5][73] ,
         \D_cache/cache[5][74] , \D_cache/cache[5][75] ,
         \D_cache/cache[5][76] , \D_cache/cache[5][77] ,
         \D_cache/cache[5][78] , \D_cache/cache[5][79] ,
         \D_cache/cache[5][80] , \D_cache/cache[5][81] ,
         \D_cache/cache[5][82] , \D_cache/cache[5][83] ,
         \D_cache/cache[5][84] , \D_cache/cache[5][85] ,
         \D_cache/cache[5][86] , \D_cache/cache[5][87] ,
         \D_cache/cache[5][88] , \D_cache/cache[5][89] ,
         \D_cache/cache[5][90] , \D_cache/cache[5][91] ,
         \D_cache/cache[5][92] , \D_cache/cache[5][93] ,
         \D_cache/cache[5][94] , \D_cache/cache[5][95] ,
         \D_cache/cache[5][96] , \D_cache/cache[5][97] ,
         \D_cache/cache[5][98] , \D_cache/cache[5][99] ,
         \D_cache/cache[5][100] , \D_cache/cache[5][101] ,
         \D_cache/cache[5][102] , \D_cache/cache[5][103] ,
         \D_cache/cache[5][104] , \D_cache/cache[5][105] ,
         \D_cache/cache[5][106] , \D_cache/cache[5][107] ,
         \D_cache/cache[5][108] , \D_cache/cache[5][109] ,
         \D_cache/cache[5][110] , \D_cache/cache[5][111] ,
         \D_cache/cache[5][112] , \D_cache/cache[5][113] ,
         \D_cache/cache[5][114] , \D_cache/cache[5][115] ,
         \D_cache/cache[5][116] , \D_cache/cache[5][117] ,
         \D_cache/cache[5][118] , \D_cache/cache[5][119] ,
         \D_cache/cache[5][120] , \D_cache/cache[5][121] ,
         \D_cache/cache[5][122] , \D_cache/cache[5][123] ,
         \D_cache/cache[5][124] , \D_cache/cache[5][125] ,
         \D_cache/cache[5][126] , \D_cache/cache[5][127] ,
         \D_cache/cache[5][128] , \D_cache/cache[5][129] ,
         \D_cache/cache[5][130] , \D_cache/cache[5][131] ,
         \D_cache/cache[5][132] , \D_cache/cache[5][133] ,
         \D_cache/cache[5][134] , \D_cache/cache[5][135] ,
         \D_cache/cache[5][136] , \D_cache/cache[5][137] ,
         \D_cache/cache[5][138] , \D_cache/cache[5][139] ,
         \D_cache/cache[5][140] , \D_cache/cache[5][141] ,
         \D_cache/cache[5][142] , \D_cache/cache[5][143] ,
         \D_cache/cache[5][144] , \D_cache/cache[5][145] ,
         \D_cache/cache[5][146] , \D_cache/cache[5][147] ,
         \D_cache/cache[5][148] , \D_cache/cache[5][149] ,
         \D_cache/cache[5][150] , \D_cache/cache[5][151] ,
         \D_cache/cache[5][152] , \D_cache/cache[5][153] ,
         \D_cache/cache[5][154] , \D_cache/cache[4][0] , \D_cache/cache[4][1] ,
         \D_cache/cache[4][2] , \D_cache/cache[4][3] , \D_cache/cache[4][4] ,
         \D_cache/cache[4][5] , \D_cache/cache[4][6] , \D_cache/cache[4][7] ,
         \D_cache/cache[4][8] , \D_cache/cache[4][9] , \D_cache/cache[4][10] ,
         \D_cache/cache[4][11] , \D_cache/cache[4][12] ,
         \D_cache/cache[4][13] , \D_cache/cache[4][14] ,
         \D_cache/cache[4][15] , \D_cache/cache[4][16] ,
         \D_cache/cache[4][17] , \D_cache/cache[4][18] ,
         \D_cache/cache[4][19] , \D_cache/cache[4][20] ,
         \D_cache/cache[4][21] , \D_cache/cache[4][22] ,
         \D_cache/cache[4][23] , \D_cache/cache[4][24] ,
         \D_cache/cache[4][25] , \D_cache/cache[4][26] ,
         \D_cache/cache[4][27] , \D_cache/cache[4][28] ,
         \D_cache/cache[4][29] , \D_cache/cache[4][30] ,
         \D_cache/cache[4][31] , \D_cache/cache[4][32] ,
         \D_cache/cache[4][33] , \D_cache/cache[4][34] ,
         \D_cache/cache[4][35] , \D_cache/cache[4][36] ,
         \D_cache/cache[4][37] , \D_cache/cache[4][38] ,
         \D_cache/cache[4][39] , \D_cache/cache[4][40] ,
         \D_cache/cache[4][41] , \D_cache/cache[4][42] ,
         \D_cache/cache[4][43] , \D_cache/cache[4][44] ,
         \D_cache/cache[4][45] , \D_cache/cache[4][46] ,
         \D_cache/cache[4][47] , \D_cache/cache[4][48] ,
         \D_cache/cache[4][49] , \D_cache/cache[4][50] ,
         \D_cache/cache[4][51] , \D_cache/cache[4][52] ,
         \D_cache/cache[4][53] , \D_cache/cache[4][54] ,
         \D_cache/cache[4][55] , \D_cache/cache[4][56] ,
         \D_cache/cache[4][57] , \D_cache/cache[4][58] ,
         \D_cache/cache[4][59] , \D_cache/cache[4][60] ,
         \D_cache/cache[4][61] , \D_cache/cache[4][62] ,
         \D_cache/cache[4][63] , \D_cache/cache[4][64] ,
         \D_cache/cache[4][65] , \D_cache/cache[4][66] ,
         \D_cache/cache[4][67] , \D_cache/cache[4][68] ,
         \D_cache/cache[4][69] , \D_cache/cache[4][70] ,
         \D_cache/cache[4][71] , \D_cache/cache[4][72] ,
         \D_cache/cache[4][73] , \D_cache/cache[4][74] ,
         \D_cache/cache[4][75] , \D_cache/cache[4][76] ,
         \D_cache/cache[4][77] , \D_cache/cache[4][78] ,
         \D_cache/cache[4][79] , \D_cache/cache[4][80] ,
         \D_cache/cache[4][81] , \D_cache/cache[4][82] ,
         \D_cache/cache[4][83] , \D_cache/cache[4][84] ,
         \D_cache/cache[4][85] , \D_cache/cache[4][86] ,
         \D_cache/cache[4][87] , \D_cache/cache[4][88] ,
         \D_cache/cache[4][89] , \D_cache/cache[4][90] ,
         \D_cache/cache[4][91] , \D_cache/cache[4][92] ,
         \D_cache/cache[4][93] , \D_cache/cache[4][94] ,
         \D_cache/cache[4][95] , \D_cache/cache[4][96] ,
         \D_cache/cache[4][97] , \D_cache/cache[4][98] ,
         \D_cache/cache[4][99] , \D_cache/cache[4][100] ,
         \D_cache/cache[4][101] , \D_cache/cache[4][102] ,
         \D_cache/cache[4][103] , \D_cache/cache[4][104] ,
         \D_cache/cache[4][105] , \D_cache/cache[4][106] ,
         \D_cache/cache[4][107] , \D_cache/cache[4][108] ,
         \D_cache/cache[4][109] , \D_cache/cache[4][110] ,
         \D_cache/cache[4][111] , \D_cache/cache[4][112] ,
         \D_cache/cache[4][113] , \D_cache/cache[4][114] ,
         \D_cache/cache[4][115] , \D_cache/cache[4][116] ,
         \D_cache/cache[4][117] , \D_cache/cache[4][118] ,
         \D_cache/cache[4][119] , \D_cache/cache[4][120] ,
         \D_cache/cache[4][121] , \D_cache/cache[4][122] ,
         \D_cache/cache[4][123] , \D_cache/cache[4][124] ,
         \D_cache/cache[4][125] , \D_cache/cache[4][126] ,
         \D_cache/cache[4][127] , \D_cache/cache[4][128] ,
         \D_cache/cache[4][129] , \D_cache/cache[4][130] ,
         \D_cache/cache[4][131] , \D_cache/cache[4][132] ,
         \D_cache/cache[4][133] , \D_cache/cache[4][134] ,
         \D_cache/cache[4][135] , \D_cache/cache[4][136] ,
         \D_cache/cache[4][137] , \D_cache/cache[4][138] ,
         \D_cache/cache[4][139] , \D_cache/cache[4][140] ,
         \D_cache/cache[4][141] , \D_cache/cache[4][142] ,
         \D_cache/cache[4][143] , \D_cache/cache[4][144] ,
         \D_cache/cache[4][145] , \D_cache/cache[4][146] ,
         \D_cache/cache[4][147] , \D_cache/cache[4][148] ,
         \D_cache/cache[4][149] , \D_cache/cache[4][150] ,
         \D_cache/cache[4][151] , \D_cache/cache[4][152] ,
         \D_cache/cache[4][153] , \D_cache/cache[4][154] ,
         \D_cache/cache[3][0] , \D_cache/cache[3][1] , \D_cache/cache[3][2] ,
         \D_cache/cache[3][3] , \D_cache/cache[3][4] , \D_cache/cache[3][5] ,
         \D_cache/cache[3][6] , \D_cache/cache[3][7] , \D_cache/cache[3][8] ,
         \D_cache/cache[3][9] , \D_cache/cache[3][10] , \D_cache/cache[3][11] ,
         \D_cache/cache[3][12] , \D_cache/cache[3][13] ,
         \D_cache/cache[3][14] , \D_cache/cache[3][15] ,
         \D_cache/cache[3][16] , \D_cache/cache[3][17] ,
         \D_cache/cache[3][18] , \D_cache/cache[3][19] ,
         \D_cache/cache[3][20] , \D_cache/cache[3][21] ,
         \D_cache/cache[3][22] , \D_cache/cache[3][23] ,
         \D_cache/cache[3][24] , \D_cache/cache[3][25] ,
         \D_cache/cache[3][26] , \D_cache/cache[3][27] ,
         \D_cache/cache[3][28] , \D_cache/cache[3][29] ,
         \D_cache/cache[3][30] , \D_cache/cache[3][31] ,
         \D_cache/cache[3][32] , \D_cache/cache[3][33] ,
         \D_cache/cache[3][34] , \D_cache/cache[3][35] ,
         \D_cache/cache[3][36] , \D_cache/cache[3][37] ,
         \D_cache/cache[3][38] , \D_cache/cache[3][39] ,
         \D_cache/cache[3][40] , \D_cache/cache[3][41] ,
         \D_cache/cache[3][42] , \D_cache/cache[3][43] ,
         \D_cache/cache[3][44] , \D_cache/cache[3][45] ,
         \D_cache/cache[3][46] , \D_cache/cache[3][47] ,
         \D_cache/cache[3][48] , \D_cache/cache[3][49] ,
         \D_cache/cache[3][50] , \D_cache/cache[3][51] ,
         \D_cache/cache[3][52] , \D_cache/cache[3][53] ,
         \D_cache/cache[3][54] , \D_cache/cache[3][55] ,
         \D_cache/cache[3][56] , \D_cache/cache[3][57] ,
         \D_cache/cache[3][58] , \D_cache/cache[3][59] ,
         \D_cache/cache[3][60] , \D_cache/cache[3][61] ,
         \D_cache/cache[3][62] , \D_cache/cache[3][63] ,
         \D_cache/cache[3][64] , \D_cache/cache[3][65] ,
         \D_cache/cache[3][66] , \D_cache/cache[3][67] ,
         \D_cache/cache[3][68] , \D_cache/cache[3][69] ,
         \D_cache/cache[3][70] , \D_cache/cache[3][71] ,
         \D_cache/cache[3][72] , \D_cache/cache[3][73] ,
         \D_cache/cache[3][74] , \D_cache/cache[3][75] ,
         \D_cache/cache[3][76] , \D_cache/cache[3][77] ,
         \D_cache/cache[3][78] , \D_cache/cache[3][79] ,
         \D_cache/cache[3][80] , \D_cache/cache[3][81] ,
         \D_cache/cache[3][82] , \D_cache/cache[3][83] ,
         \D_cache/cache[3][84] , \D_cache/cache[3][85] ,
         \D_cache/cache[3][86] , \D_cache/cache[3][87] ,
         \D_cache/cache[3][88] , \D_cache/cache[3][89] ,
         \D_cache/cache[3][90] , \D_cache/cache[3][91] ,
         \D_cache/cache[3][92] , \D_cache/cache[3][93] ,
         \D_cache/cache[3][94] , \D_cache/cache[3][95] ,
         \D_cache/cache[3][96] , \D_cache/cache[3][97] ,
         \D_cache/cache[3][98] , \D_cache/cache[3][99] ,
         \D_cache/cache[3][100] , \D_cache/cache[3][101] ,
         \D_cache/cache[3][102] , \D_cache/cache[3][103] ,
         \D_cache/cache[3][104] , \D_cache/cache[3][105] ,
         \D_cache/cache[3][106] , \D_cache/cache[3][107] ,
         \D_cache/cache[3][108] , \D_cache/cache[3][109] ,
         \D_cache/cache[3][110] , \D_cache/cache[3][111] ,
         \D_cache/cache[3][112] , \D_cache/cache[3][113] ,
         \D_cache/cache[3][114] , \D_cache/cache[3][115] ,
         \D_cache/cache[3][116] , \D_cache/cache[3][117] ,
         \D_cache/cache[3][118] , \D_cache/cache[3][119] ,
         \D_cache/cache[3][120] , \D_cache/cache[3][121] ,
         \D_cache/cache[3][122] , \D_cache/cache[3][123] ,
         \D_cache/cache[3][124] , \D_cache/cache[3][125] ,
         \D_cache/cache[3][126] , \D_cache/cache[3][127] ,
         \D_cache/cache[3][128] , \D_cache/cache[3][129] ,
         \D_cache/cache[3][130] , \D_cache/cache[3][131] ,
         \D_cache/cache[3][132] , \D_cache/cache[3][133] ,
         \D_cache/cache[3][134] , \D_cache/cache[3][135] ,
         \D_cache/cache[3][136] , \D_cache/cache[3][137] ,
         \D_cache/cache[3][138] , \D_cache/cache[3][139] ,
         \D_cache/cache[3][140] , \D_cache/cache[3][141] ,
         \D_cache/cache[3][142] , \D_cache/cache[3][143] ,
         \D_cache/cache[3][144] , \D_cache/cache[3][145] ,
         \D_cache/cache[3][146] , \D_cache/cache[3][147] ,
         \D_cache/cache[3][148] , \D_cache/cache[3][149] ,
         \D_cache/cache[3][150] , \D_cache/cache[3][151] ,
         \D_cache/cache[3][152] , \D_cache/cache[3][153] ,
         \D_cache/cache[3][154] , \D_cache/cache[2][0] , \D_cache/cache[2][1] ,
         \D_cache/cache[2][2] , \D_cache/cache[2][3] , \D_cache/cache[2][4] ,
         \D_cache/cache[2][5] , \D_cache/cache[2][6] , \D_cache/cache[2][7] ,
         \D_cache/cache[2][8] , \D_cache/cache[2][9] , \D_cache/cache[2][10] ,
         \D_cache/cache[2][11] , \D_cache/cache[2][12] ,
         \D_cache/cache[2][13] , \D_cache/cache[2][14] ,
         \D_cache/cache[2][15] , \D_cache/cache[2][16] ,
         \D_cache/cache[2][17] , \D_cache/cache[2][18] ,
         \D_cache/cache[2][19] , \D_cache/cache[2][20] ,
         \D_cache/cache[2][21] , \D_cache/cache[2][22] ,
         \D_cache/cache[2][23] , \D_cache/cache[2][24] ,
         \D_cache/cache[2][25] , \D_cache/cache[2][26] ,
         \D_cache/cache[2][27] , \D_cache/cache[2][28] ,
         \D_cache/cache[2][29] , \D_cache/cache[2][30] ,
         \D_cache/cache[2][31] , \D_cache/cache[2][32] ,
         \D_cache/cache[2][33] , \D_cache/cache[2][34] ,
         \D_cache/cache[2][35] , \D_cache/cache[2][36] ,
         \D_cache/cache[2][37] , \D_cache/cache[2][38] ,
         \D_cache/cache[2][39] , \D_cache/cache[2][40] ,
         \D_cache/cache[2][41] , \D_cache/cache[2][42] ,
         \D_cache/cache[2][43] , \D_cache/cache[2][44] ,
         \D_cache/cache[2][45] , \D_cache/cache[2][46] ,
         \D_cache/cache[2][47] , \D_cache/cache[2][48] ,
         \D_cache/cache[2][49] , \D_cache/cache[2][50] ,
         \D_cache/cache[2][51] , \D_cache/cache[2][52] ,
         \D_cache/cache[2][53] , \D_cache/cache[2][54] ,
         \D_cache/cache[2][55] , \D_cache/cache[2][56] ,
         \D_cache/cache[2][57] , \D_cache/cache[2][58] ,
         \D_cache/cache[2][59] , \D_cache/cache[2][60] ,
         \D_cache/cache[2][61] , \D_cache/cache[2][62] ,
         \D_cache/cache[2][63] , \D_cache/cache[2][64] ,
         \D_cache/cache[2][65] , \D_cache/cache[2][66] ,
         \D_cache/cache[2][67] , \D_cache/cache[2][68] ,
         \D_cache/cache[2][69] , \D_cache/cache[2][70] ,
         \D_cache/cache[2][71] , \D_cache/cache[2][72] ,
         \D_cache/cache[2][73] , \D_cache/cache[2][74] ,
         \D_cache/cache[2][75] , \D_cache/cache[2][76] ,
         \D_cache/cache[2][77] , \D_cache/cache[2][78] ,
         \D_cache/cache[2][79] , \D_cache/cache[2][80] ,
         \D_cache/cache[2][81] , \D_cache/cache[2][82] ,
         \D_cache/cache[2][83] , \D_cache/cache[2][84] ,
         \D_cache/cache[2][85] , \D_cache/cache[2][86] ,
         \D_cache/cache[2][87] , \D_cache/cache[2][88] ,
         \D_cache/cache[2][89] , \D_cache/cache[2][90] ,
         \D_cache/cache[2][91] , \D_cache/cache[2][92] ,
         \D_cache/cache[2][93] , \D_cache/cache[2][94] ,
         \D_cache/cache[2][95] , \D_cache/cache[2][96] ,
         \D_cache/cache[2][97] , \D_cache/cache[2][98] ,
         \D_cache/cache[2][99] , \D_cache/cache[2][100] ,
         \D_cache/cache[2][101] , \D_cache/cache[2][102] ,
         \D_cache/cache[2][103] , \D_cache/cache[2][104] ,
         \D_cache/cache[2][105] , \D_cache/cache[2][106] ,
         \D_cache/cache[2][107] , \D_cache/cache[2][108] ,
         \D_cache/cache[2][109] , \D_cache/cache[2][110] ,
         \D_cache/cache[2][111] , \D_cache/cache[2][112] ,
         \D_cache/cache[2][113] , \D_cache/cache[2][114] ,
         \D_cache/cache[2][115] , \D_cache/cache[2][116] ,
         \D_cache/cache[2][117] , \D_cache/cache[2][118] ,
         \D_cache/cache[2][119] , \D_cache/cache[2][120] ,
         \D_cache/cache[2][121] , \D_cache/cache[2][122] ,
         \D_cache/cache[2][123] , \D_cache/cache[2][124] ,
         \D_cache/cache[2][125] , \D_cache/cache[2][126] ,
         \D_cache/cache[2][127] , \D_cache/cache[2][128] ,
         \D_cache/cache[2][129] , \D_cache/cache[2][130] ,
         \D_cache/cache[2][131] , \D_cache/cache[2][132] ,
         \D_cache/cache[2][133] , \D_cache/cache[2][134] ,
         \D_cache/cache[2][135] , \D_cache/cache[2][136] ,
         \D_cache/cache[2][137] , \D_cache/cache[2][138] ,
         \D_cache/cache[2][139] , \D_cache/cache[2][140] ,
         \D_cache/cache[2][141] , \D_cache/cache[2][142] ,
         \D_cache/cache[2][143] , \D_cache/cache[2][144] ,
         \D_cache/cache[2][145] , \D_cache/cache[2][146] ,
         \D_cache/cache[2][147] , \D_cache/cache[2][148] ,
         \D_cache/cache[2][149] , \D_cache/cache[2][150] ,
         \D_cache/cache[2][151] , \D_cache/cache[2][152] ,
         \D_cache/cache[2][153] , \D_cache/cache[2][154] ,
         \D_cache/cache[1][0] , \D_cache/cache[1][1] , \D_cache/cache[1][2] ,
         \D_cache/cache[1][3] , \D_cache/cache[1][4] , \D_cache/cache[1][5] ,
         \D_cache/cache[1][6] , \D_cache/cache[1][7] , \D_cache/cache[1][8] ,
         \D_cache/cache[1][9] , \D_cache/cache[1][10] , \D_cache/cache[1][11] ,
         \D_cache/cache[1][12] , \D_cache/cache[1][13] ,
         \D_cache/cache[1][14] , \D_cache/cache[1][15] ,
         \D_cache/cache[1][16] , \D_cache/cache[1][17] ,
         \D_cache/cache[1][18] , \D_cache/cache[1][19] ,
         \D_cache/cache[1][20] , \D_cache/cache[1][21] ,
         \D_cache/cache[1][22] , \D_cache/cache[1][23] ,
         \D_cache/cache[1][24] , \D_cache/cache[1][25] ,
         \D_cache/cache[1][26] , \D_cache/cache[1][27] ,
         \D_cache/cache[1][28] , \D_cache/cache[1][29] ,
         \D_cache/cache[1][30] , \D_cache/cache[1][31] ,
         \D_cache/cache[1][32] , \D_cache/cache[1][33] ,
         \D_cache/cache[1][34] , \D_cache/cache[1][35] ,
         \D_cache/cache[1][36] , \D_cache/cache[1][37] ,
         \D_cache/cache[1][38] , \D_cache/cache[1][39] ,
         \D_cache/cache[1][40] , \D_cache/cache[1][41] ,
         \D_cache/cache[1][42] , \D_cache/cache[1][43] ,
         \D_cache/cache[1][44] , \D_cache/cache[1][45] ,
         \D_cache/cache[1][46] , \D_cache/cache[1][47] ,
         \D_cache/cache[1][48] , \D_cache/cache[1][49] ,
         \D_cache/cache[1][50] , \D_cache/cache[1][51] ,
         \D_cache/cache[1][52] , \D_cache/cache[1][53] ,
         \D_cache/cache[1][54] , \D_cache/cache[1][55] ,
         \D_cache/cache[1][56] , \D_cache/cache[1][57] ,
         \D_cache/cache[1][58] , \D_cache/cache[1][59] ,
         \D_cache/cache[1][60] , \D_cache/cache[1][61] ,
         \D_cache/cache[1][62] , \D_cache/cache[1][63] ,
         \D_cache/cache[1][64] , \D_cache/cache[1][65] ,
         \D_cache/cache[1][66] , \D_cache/cache[1][67] ,
         \D_cache/cache[1][68] , \D_cache/cache[1][69] ,
         \D_cache/cache[1][70] , \D_cache/cache[1][71] ,
         \D_cache/cache[1][72] , \D_cache/cache[1][73] ,
         \D_cache/cache[1][74] , \D_cache/cache[1][75] ,
         \D_cache/cache[1][76] , \D_cache/cache[1][77] ,
         \D_cache/cache[1][78] , \D_cache/cache[1][79] ,
         \D_cache/cache[1][80] , \D_cache/cache[1][81] ,
         \D_cache/cache[1][82] , \D_cache/cache[1][83] ,
         \D_cache/cache[1][84] , \D_cache/cache[1][85] ,
         \D_cache/cache[1][86] , \D_cache/cache[1][87] ,
         \D_cache/cache[1][88] , \D_cache/cache[1][89] ,
         \D_cache/cache[1][90] , \D_cache/cache[1][91] ,
         \D_cache/cache[1][92] , \D_cache/cache[1][93] ,
         \D_cache/cache[1][94] , \D_cache/cache[1][95] ,
         \D_cache/cache[1][96] , \D_cache/cache[1][97] ,
         \D_cache/cache[1][98] , \D_cache/cache[1][99] ,
         \D_cache/cache[1][100] , \D_cache/cache[1][101] ,
         \D_cache/cache[1][102] , \D_cache/cache[1][103] ,
         \D_cache/cache[1][104] , \D_cache/cache[1][105] ,
         \D_cache/cache[1][106] , \D_cache/cache[1][107] ,
         \D_cache/cache[1][108] , \D_cache/cache[1][109] ,
         \D_cache/cache[1][110] , \D_cache/cache[1][111] ,
         \D_cache/cache[1][112] , \D_cache/cache[1][113] ,
         \D_cache/cache[1][114] , \D_cache/cache[1][115] ,
         \D_cache/cache[1][116] , \D_cache/cache[1][117] ,
         \D_cache/cache[1][118] , \D_cache/cache[1][119] ,
         \D_cache/cache[1][120] , \D_cache/cache[1][121] ,
         \D_cache/cache[1][122] , \D_cache/cache[1][123] ,
         \D_cache/cache[1][124] , \D_cache/cache[1][125] ,
         \D_cache/cache[1][126] , \D_cache/cache[1][127] ,
         \D_cache/cache[1][128] , \D_cache/cache[1][129] ,
         \D_cache/cache[1][130] , \D_cache/cache[1][131] ,
         \D_cache/cache[1][132] , \D_cache/cache[1][133] ,
         \D_cache/cache[1][134] , \D_cache/cache[1][135] ,
         \D_cache/cache[1][136] , \D_cache/cache[1][137] ,
         \D_cache/cache[1][138] , \D_cache/cache[1][139] ,
         \D_cache/cache[1][140] , \D_cache/cache[1][141] ,
         \D_cache/cache[1][142] , \D_cache/cache[1][143] ,
         \D_cache/cache[1][144] , \D_cache/cache[1][145] ,
         \D_cache/cache[1][146] , \D_cache/cache[1][147] ,
         \D_cache/cache[1][148] , \D_cache/cache[1][149] ,
         \D_cache/cache[1][150] , \D_cache/cache[1][151] ,
         \D_cache/cache[1][152] , \D_cache/cache[1][153] ,
         \D_cache/cache[1][154] , \D_cache/cache[0][0] , \D_cache/cache[0][1] ,
         \D_cache/cache[0][2] , \D_cache/cache[0][3] , \D_cache/cache[0][4] ,
         \D_cache/cache[0][5] , \D_cache/cache[0][6] , \D_cache/cache[0][7] ,
         \D_cache/cache[0][8] , \D_cache/cache[0][9] , \D_cache/cache[0][10] ,
         \D_cache/cache[0][11] , \D_cache/cache[0][12] ,
         \D_cache/cache[0][13] , \D_cache/cache[0][14] ,
         \D_cache/cache[0][15] , \D_cache/cache[0][16] ,
         \D_cache/cache[0][17] , \D_cache/cache[0][18] ,
         \D_cache/cache[0][19] , \D_cache/cache[0][20] ,
         \D_cache/cache[0][21] , \D_cache/cache[0][22] ,
         \D_cache/cache[0][23] , \D_cache/cache[0][24] ,
         \D_cache/cache[0][25] , \D_cache/cache[0][26] ,
         \D_cache/cache[0][27] , \D_cache/cache[0][28] ,
         \D_cache/cache[0][29] , \D_cache/cache[0][30] ,
         \D_cache/cache[0][31] , \D_cache/cache[0][32] ,
         \D_cache/cache[0][33] , \D_cache/cache[0][34] ,
         \D_cache/cache[0][35] , \D_cache/cache[0][36] ,
         \D_cache/cache[0][37] , \D_cache/cache[0][38] ,
         \D_cache/cache[0][39] , \D_cache/cache[0][40] ,
         \D_cache/cache[0][41] , \D_cache/cache[0][42] ,
         \D_cache/cache[0][43] , \D_cache/cache[0][44] ,
         \D_cache/cache[0][45] , \D_cache/cache[0][46] ,
         \D_cache/cache[0][47] , \D_cache/cache[0][48] ,
         \D_cache/cache[0][49] , \D_cache/cache[0][50] ,
         \D_cache/cache[0][51] , \D_cache/cache[0][52] ,
         \D_cache/cache[0][53] , \D_cache/cache[0][54] ,
         \D_cache/cache[0][55] , \D_cache/cache[0][56] ,
         \D_cache/cache[0][57] , \D_cache/cache[0][58] ,
         \D_cache/cache[0][59] , \D_cache/cache[0][60] ,
         \D_cache/cache[0][61] , \D_cache/cache[0][62] ,
         \D_cache/cache[0][63] , \D_cache/cache[0][64] ,
         \D_cache/cache[0][65] , \D_cache/cache[0][66] ,
         \D_cache/cache[0][67] , \D_cache/cache[0][68] ,
         \D_cache/cache[0][69] , \D_cache/cache[0][70] ,
         \D_cache/cache[0][71] , \D_cache/cache[0][72] ,
         \D_cache/cache[0][73] , \D_cache/cache[0][74] ,
         \D_cache/cache[0][75] , \D_cache/cache[0][76] ,
         \D_cache/cache[0][77] , \D_cache/cache[0][78] ,
         \D_cache/cache[0][79] , \D_cache/cache[0][80] ,
         \D_cache/cache[0][81] , \D_cache/cache[0][82] ,
         \D_cache/cache[0][83] , \D_cache/cache[0][84] ,
         \D_cache/cache[0][85] , \D_cache/cache[0][86] ,
         \D_cache/cache[0][87] , \D_cache/cache[0][88] ,
         \D_cache/cache[0][89] , \D_cache/cache[0][90] ,
         \D_cache/cache[0][91] , \D_cache/cache[0][92] ,
         \D_cache/cache[0][93] , \D_cache/cache[0][94] ,
         \D_cache/cache[0][95] , \D_cache/cache[0][96] ,
         \D_cache/cache[0][97] , \D_cache/cache[0][98] ,
         \D_cache/cache[0][99] , \D_cache/cache[0][100] ,
         \D_cache/cache[0][101] , \D_cache/cache[0][102] ,
         \D_cache/cache[0][103] , \D_cache/cache[0][104] ,
         \D_cache/cache[0][105] , \D_cache/cache[0][106] ,
         \D_cache/cache[0][107] , \D_cache/cache[0][108] ,
         \D_cache/cache[0][109] , \D_cache/cache[0][110] ,
         \D_cache/cache[0][111] , \D_cache/cache[0][112] ,
         \D_cache/cache[0][113] , \D_cache/cache[0][114] ,
         \D_cache/cache[0][115] , \D_cache/cache[0][116] ,
         \D_cache/cache[0][117] , \D_cache/cache[0][118] ,
         \D_cache/cache[0][119] , \D_cache/cache[0][120] ,
         \D_cache/cache[0][121] , \D_cache/cache[0][122] ,
         \D_cache/cache[0][123] , \D_cache/cache[0][124] ,
         \D_cache/cache[0][125] , \D_cache/cache[0][126] ,
         \D_cache/cache[0][127] , \D_cache/cache[0][128] ,
         \D_cache/cache[0][129] , \D_cache/cache[0][130] ,
         \D_cache/cache[0][131] , \D_cache/cache[0][132] ,
         \D_cache/cache[0][133] , \D_cache/cache[0][134] ,
         \D_cache/cache[0][135] , \D_cache/cache[0][136] ,
         \D_cache/cache[0][137] , \D_cache/cache[0][138] ,
         \D_cache/cache[0][139] , \D_cache/cache[0][140] ,
         \D_cache/cache[0][141] , \D_cache/cache[0][142] ,
         \D_cache/cache[0][143] , \D_cache/cache[0][144] ,
         \D_cache/cache[0][145] , \D_cache/cache[0][146] ,
         \D_cache/cache[0][147] , \D_cache/cache[0][148] ,
         \D_cache/cache[0][149] , \D_cache/cache[0][150] ,
         \D_cache/cache[0][151] , \D_cache/cache[0][152] ,
         \D_cache/cache[0][153] , \D_cache/cache[0][154] ,
         \i_MIPS/Pred_1bit/n2 , \i_MIPS/Pred_1bit/current_state ,
         \i_MIPS/PC/n65 , \i_MIPS/PC/n64 , \i_MIPS/PC/n63 , \i_MIPS/PC/n62 ,
         \i_MIPS/PC/n61 , \i_MIPS/PC/n60 , \i_MIPS/PC/n59 , \i_MIPS/PC/n58 ,
         \i_MIPS/PC/n57 , \i_MIPS/PC/n56 , \i_MIPS/PC/n55 , \i_MIPS/PC/n54 ,
         \i_MIPS/PC/n53 , \i_MIPS/PC/n52 , \i_MIPS/PC/n51 , \i_MIPS/PC/n50 ,
         \i_MIPS/PC/n49 , \i_MIPS/PC/n48 , \i_MIPS/PC/n47 , \i_MIPS/PC/n46 ,
         \i_MIPS/PC/n45 , \i_MIPS/PC/n44 , \i_MIPS/PC/n43 , \i_MIPS/PC/n42 ,
         \i_MIPS/PC/n41 , \i_MIPS/PC/n40 , \i_MIPS/PC/n39 , \i_MIPS/PC/n38 ,
         \i_MIPS/PC/n37 , \i_MIPS/PC/n36 , \i_MIPS/PC/n35 , \i_MIPS/PC/n34 ,
         \i_MIPS/PC/n33 , \i_MIPS/PC/n32 , \i_MIPS/PC/n31 , \i_MIPS/PC/n30 ,
         \i_MIPS/PC/n29 , \i_MIPS/PC/n28 , \i_MIPS/PC/n27 , \i_MIPS/PC/n26 ,
         \i_MIPS/PC/n25 , \i_MIPS/PC/n24 , \i_MIPS/PC/n23 , \i_MIPS/PC/n22 ,
         \i_MIPS/PC/n21 , \i_MIPS/PC/n20 , \i_MIPS/PC/n19 , \i_MIPS/PC/n18 ,
         \i_MIPS/PC/n17 , \i_MIPS/PC/n16 , \i_MIPS/PC/n15 , \i_MIPS/PC/n14 ,
         \i_MIPS/PC/n13 , \i_MIPS/PC/n12 , \i_MIPS/PC/n11 , \i_MIPS/PC/n10 ,
         \i_MIPS/PC/n9 , \i_MIPS/PC/n8 , \i_MIPS/PC/n7 , \i_MIPS/PC/n6 ,
         \i_MIPS/PC/n5 , \i_MIPS/PC/n4 , \i_MIPS/PC/n3 , \i_MIPS/PC/n2 ,
         \i_MIPS/Register/n1139 , \i_MIPS/Register/n1138 ,
         \i_MIPS/Register/n1137 , \i_MIPS/Register/n1136 ,
         \i_MIPS/Register/n1135 , \i_MIPS/Register/n1134 ,
         \i_MIPS/Register/n1133 , \i_MIPS/Register/n1132 ,
         \i_MIPS/Register/n1131 , \i_MIPS/Register/n1130 ,
         \i_MIPS/Register/n1129 , \i_MIPS/Register/n1128 ,
         \i_MIPS/Register/n1127 , \i_MIPS/Register/n1126 ,
         \i_MIPS/Register/n1125 , \i_MIPS/Register/n1124 ,
         \i_MIPS/Register/n1123 , \i_MIPS/Register/n1122 ,
         \i_MIPS/Register/n1121 , \i_MIPS/Register/n1120 ,
         \i_MIPS/Register/n1119 , \i_MIPS/Register/n1118 ,
         \i_MIPS/Register/n1117 , \i_MIPS/Register/n1116 ,
         \i_MIPS/Register/n1115 , \i_MIPS/Register/n1114 ,
         \i_MIPS/Register/n1113 , \i_MIPS/Register/n1112 ,
         \i_MIPS/Register/n1111 , \i_MIPS/Register/n1110 ,
         \i_MIPS/Register/n1109 , \i_MIPS/Register/n1108 ,
         \i_MIPS/Register/n1107 , \i_MIPS/Register/n1106 ,
         \i_MIPS/Register/n1105 , \i_MIPS/Register/n1104 ,
         \i_MIPS/Register/n1103 , \i_MIPS/Register/n1102 ,
         \i_MIPS/Register/n1101 , \i_MIPS/Register/n1100 ,
         \i_MIPS/Register/n1099 , \i_MIPS/Register/n1098 ,
         \i_MIPS/Register/n1097 , \i_MIPS/Register/n1096 ,
         \i_MIPS/Register/n1095 , \i_MIPS/Register/n1094 ,
         \i_MIPS/Register/n1093 , \i_MIPS/Register/n1092 ,
         \i_MIPS/Register/n1091 , \i_MIPS/Register/n1090 ,
         \i_MIPS/Register/n1089 , \i_MIPS/Register/n1088 ,
         \i_MIPS/Register/n1087 , \i_MIPS/Register/n1086 ,
         \i_MIPS/Register/n1085 , \i_MIPS/Register/n1084 ,
         \i_MIPS/Register/n1083 , \i_MIPS/Register/n1082 ,
         \i_MIPS/Register/n1081 , \i_MIPS/Register/n1080 ,
         \i_MIPS/Register/n1079 , \i_MIPS/Register/n1078 ,
         \i_MIPS/Register/n1077 , \i_MIPS/Register/n1076 ,
         \i_MIPS/Register/n1075 , \i_MIPS/Register/n1074 ,
         \i_MIPS/Register/n1073 , \i_MIPS/Register/n1072 ,
         \i_MIPS/Register/n1071 , \i_MIPS/Register/n1070 ,
         \i_MIPS/Register/n1069 , \i_MIPS/Register/n1068 ,
         \i_MIPS/Register/n1067 , \i_MIPS/Register/n1066 ,
         \i_MIPS/Register/n1065 , \i_MIPS/Register/n1064 ,
         \i_MIPS/Register/n1063 , \i_MIPS/Register/n1062 ,
         \i_MIPS/Register/n1061 , \i_MIPS/Register/n1060 ,
         \i_MIPS/Register/n1059 , \i_MIPS/Register/n1058 ,
         \i_MIPS/Register/n1057 , \i_MIPS/Register/n1056 ,
         \i_MIPS/Register/n1055 , \i_MIPS/Register/n1054 ,
         \i_MIPS/Register/n1053 , \i_MIPS/Register/n1052 ,
         \i_MIPS/Register/n1051 , \i_MIPS/Register/n1050 ,
         \i_MIPS/Register/n1049 , \i_MIPS/Register/n1048 ,
         \i_MIPS/Register/n1047 , \i_MIPS/Register/n1046 ,
         \i_MIPS/Register/n1045 , \i_MIPS/Register/n1044 ,
         \i_MIPS/Register/n1043 , \i_MIPS/Register/n1042 ,
         \i_MIPS/Register/n1041 , \i_MIPS/Register/n1040 ,
         \i_MIPS/Register/n1039 , \i_MIPS/Register/n1038 ,
         \i_MIPS/Register/n1037 , \i_MIPS/Register/n1036 ,
         \i_MIPS/Register/n1035 , \i_MIPS/Register/n1034 ,
         \i_MIPS/Register/n1033 , \i_MIPS/Register/n1032 ,
         \i_MIPS/Register/n1031 , \i_MIPS/Register/n1030 ,
         \i_MIPS/Register/n1029 , \i_MIPS/Register/n1028 ,
         \i_MIPS/Register/n1027 , \i_MIPS/Register/n1026 ,
         \i_MIPS/Register/n1025 , \i_MIPS/Register/n1024 ,
         \i_MIPS/Register/n1023 , \i_MIPS/Register/n1022 ,
         \i_MIPS/Register/n1021 , \i_MIPS/Register/n1020 ,
         \i_MIPS/Register/n1019 , \i_MIPS/Register/n1018 ,
         \i_MIPS/Register/n1017 , \i_MIPS/Register/n1016 ,
         \i_MIPS/Register/n1015 , \i_MIPS/Register/n1014 ,
         \i_MIPS/Register/n1013 , \i_MIPS/Register/n1012 ,
         \i_MIPS/Register/n1011 , \i_MIPS/Register/n1010 ,
         \i_MIPS/Register/n1009 , \i_MIPS/Register/n1008 ,
         \i_MIPS/Register/n1007 , \i_MIPS/Register/n1006 ,
         \i_MIPS/Register/n1005 , \i_MIPS/Register/n1004 ,
         \i_MIPS/Register/n1003 , \i_MIPS/Register/n1002 ,
         \i_MIPS/Register/n1001 , \i_MIPS/Register/n1000 ,
         \i_MIPS/Register/n999 , \i_MIPS/Register/n998 ,
         \i_MIPS/Register/n997 , \i_MIPS/Register/n996 ,
         \i_MIPS/Register/n995 , \i_MIPS/Register/n994 ,
         \i_MIPS/Register/n993 , \i_MIPS/Register/n992 ,
         \i_MIPS/Register/n991 , \i_MIPS/Register/n990 ,
         \i_MIPS/Register/n989 , \i_MIPS/Register/n988 ,
         \i_MIPS/Register/n987 , \i_MIPS/Register/n986 ,
         \i_MIPS/Register/n985 , \i_MIPS/Register/n984 ,
         \i_MIPS/Register/n983 , \i_MIPS/Register/n982 ,
         \i_MIPS/Register/n981 , \i_MIPS/Register/n980 ,
         \i_MIPS/Register/n979 , \i_MIPS/Register/n978 ,
         \i_MIPS/Register/n977 , \i_MIPS/Register/n976 ,
         \i_MIPS/Register/n975 , \i_MIPS/Register/n974 ,
         \i_MIPS/Register/n973 , \i_MIPS/Register/n972 ,
         \i_MIPS/Register/n971 , \i_MIPS/Register/n970 ,
         \i_MIPS/Register/n969 , \i_MIPS/Register/n968 ,
         \i_MIPS/Register/n967 , \i_MIPS/Register/n966 ,
         \i_MIPS/Register/n965 , \i_MIPS/Register/n964 ,
         \i_MIPS/Register/n963 , \i_MIPS/Register/n962 ,
         \i_MIPS/Register/n961 , \i_MIPS/Register/n960 ,
         \i_MIPS/Register/n959 , \i_MIPS/Register/n958 ,
         \i_MIPS/Register/n957 , \i_MIPS/Register/n956 ,
         \i_MIPS/Register/n955 , \i_MIPS/Register/n954 ,
         \i_MIPS/Register/n953 , \i_MIPS/Register/n952 ,
         \i_MIPS/Register/n951 , \i_MIPS/Register/n950 ,
         \i_MIPS/Register/n949 , \i_MIPS/Register/n948 ,
         \i_MIPS/Register/n947 , \i_MIPS/Register/n946 ,
         \i_MIPS/Register/n945 , \i_MIPS/Register/n944 ,
         \i_MIPS/Register/n943 , \i_MIPS/Register/n942 ,
         \i_MIPS/Register/n941 , \i_MIPS/Register/n940 ,
         \i_MIPS/Register/n939 , \i_MIPS/Register/n938 ,
         \i_MIPS/Register/n937 , \i_MIPS/Register/n936 ,
         \i_MIPS/Register/n935 , \i_MIPS/Register/n934 ,
         \i_MIPS/Register/n933 , \i_MIPS/Register/n932 ,
         \i_MIPS/Register/n931 , \i_MIPS/Register/n930 ,
         \i_MIPS/Register/n929 , \i_MIPS/Register/n928 ,
         \i_MIPS/Register/n927 , \i_MIPS/Register/n926 ,
         \i_MIPS/Register/n925 , \i_MIPS/Register/n924 ,
         \i_MIPS/Register/n923 , \i_MIPS/Register/n922 ,
         \i_MIPS/Register/n921 , \i_MIPS/Register/n920 ,
         \i_MIPS/Register/n919 , \i_MIPS/Register/n918 ,
         \i_MIPS/Register/n917 , \i_MIPS/Register/n916 ,
         \i_MIPS/Register/n915 , \i_MIPS/Register/n914 ,
         \i_MIPS/Register/n913 , \i_MIPS/Register/n912 ,
         \i_MIPS/Register/n911 , \i_MIPS/Register/n910 ,
         \i_MIPS/Register/n909 , \i_MIPS/Register/n908 ,
         \i_MIPS/Register/n907 , \i_MIPS/Register/n906 ,
         \i_MIPS/Register/n905 , \i_MIPS/Register/n904 ,
         \i_MIPS/Register/n903 , \i_MIPS/Register/n902 ,
         \i_MIPS/Register/n901 , \i_MIPS/Register/n900 ,
         \i_MIPS/Register/n899 , \i_MIPS/Register/n898 ,
         \i_MIPS/Register/n897 , \i_MIPS/Register/n896 ,
         \i_MIPS/Register/n895 , \i_MIPS/Register/n894 ,
         \i_MIPS/Register/n893 , \i_MIPS/Register/n892 ,
         \i_MIPS/Register/n891 , \i_MIPS/Register/n890 ,
         \i_MIPS/Register/n889 , \i_MIPS/Register/n888 ,
         \i_MIPS/Register/n887 , \i_MIPS/Register/n886 ,
         \i_MIPS/Register/n885 , \i_MIPS/Register/n884 ,
         \i_MIPS/Register/n883 , \i_MIPS/Register/n882 ,
         \i_MIPS/Register/n881 , \i_MIPS/Register/n880 ,
         \i_MIPS/Register/n879 , \i_MIPS/Register/n878 ,
         \i_MIPS/Register/n877 , \i_MIPS/Register/n876 ,
         \i_MIPS/Register/n875 , \i_MIPS/Register/n874 ,
         \i_MIPS/Register/n873 , \i_MIPS/Register/n872 ,
         \i_MIPS/Register/n871 , \i_MIPS/Register/n870 ,
         \i_MIPS/Register/n869 , \i_MIPS/Register/n868 ,
         \i_MIPS/Register/n867 , \i_MIPS/Register/n866 ,
         \i_MIPS/Register/n865 , \i_MIPS/Register/n864 ,
         \i_MIPS/Register/n863 , \i_MIPS/Register/n862 ,
         \i_MIPS/Register/n861 , \i_MIPS/Register/n860 ,
         \i_MIPS/Register/n859 , \i_MIPS/Register/n858 ,
         \i_MIPS/Register/n857 , \i_MIPS/Register/n856 ,
         \i_MIPS/Register/n855 , \i_MIPS/Register/n854 ,
         \i_MIPS/Register/n853 , \i_MIPS/Register/n852 ,
         \i_MIPS/Register/n851 , \i_MIPS/Register/n850 ,
         \i_MIPS/Register/n849 , \i_MIPS/Register/n848 ,
         \i_MIPS/Register/n847 , \i_MIPS/Register/n846 ,
         \i_MIPS/Register/n845 , \i_MIPS/Register/n844 ,
         \i_MIPS/Register/n843 , \i_MIPS/Register/n842 ,
         \i_MIPS/Register/n841 , \i_MIPS/Register/n840 ,
         \i_MIPS/Register/n839 , \i_MIPS/Register/n838 ,
         \i_MIPS/Register/n837 , \i_MIPS/Register/n836 ,
         \i_MIPS/Register/n835 , \i_MIPS/Register/n834 ,
         \i_MIPS/Register/n833 , \i_MIPS/Register/n832 ,
         \i_MIPS/Register/n831 , \i_MIPS/Register/n830 ,
         \i_MIPS/Register/n829 , \i_MIPS/Register/n828 ,
         \i_MIPS/Register/n827 , \i_MIPS/Register/n826 ,
         \i_MIPS/Register/n825 , \i_MIPS/Register/n824 ,
         \i_MIPS/Register/n823 , \i_MIPS/Register/n822 ,
         \i_MIPS/Register/n821 , \i_MIPS/Register/n820 ,
         \i_MIPS/Register/n819 , \i_MIPS/Register/n818 ,
         \i_MIPS/Register/n817 , \i_MIPS/Register/n816 ,
         \i_MIPS/Register/n815 , \i_MIPS/Register/n814 ,
         \i_MIPS/Register/n813 , \i_MIPS/Register/n812 ,
         \i_MIPS/Register/n811 , \i_MIPS/Register/n810 ,
         \i_MIPS/Register/n809 , \i_MIPS/Register/n808 ,
         \i_MIPS/Register/n807 , \i_MIPS/Register/n806 ,
         \i_MIPS/Register/n805 , \i_MIPS/Register/n804 ,
         \i_MIPS/Register/n803 , \i_MIPS/Register/n802 ,
         \i_MIPS/Register/n801 , \i_MIPS/Register/n800 ,
         \i_MIPS/Register/n799 , \i_MIPS/Register/n798 ,
         \i_MIPS/Register/n797 , \i_MIPS/Register/n796 ,
         \i_MIPS/Register/n795 , \i_MIPS/Register/n794 ,
         \i_MIPS/Register/n793 , \i_MIPS/Register/n792 ,
         \i_MIPS/Register/n791 , \i_MIPS/Register/n790 ,
         \i_MIPS/Register/n789 , \i_MIPS/Register/n788 ,
         \i_MIPS/Register/n787 , \i_MIPS/Register/n786 ,
         \i_MIPS/Register/n785 , \i_MIPS/Register/n784 ,
         \i_MIPS/Register/n783 , \i_MIPS/Register/n782 ,
         \i_MIPS/Register/n781 , \i_MIPS/Register/n780 ,
         \i_MIPS/Register/n779 , \i_MIPS/Register/n778 ,
         \i_MIPS/Register/n777 , \i_MIPS/Register/n776 ,
         \i_MIPS/Register/n775 , \i_MIPS/Register/n774 ,
         \i_MIPS/Register/n773 , \i_MIPS/Register/n772 ,
         \i_MIPS/Register/n771 , \i_MIPS/Register/n770 ,
         \i_MIPS/Register/n769 , \i_MIPS/Register/n768 ,
         \i_MIPS/Register/n767 , \i_MIPS/Register/n766 ,
         \i_MIPS/Register/n765 , \i_MIPS/Register/n764 ,
         \i_MIPS/Register/n763 , \i_MIPS/Register/n762 ,
         \i_MIPS/Register/n761 , \i_MIPS/Register/n760 ,
         \i_MIPS/Register/n759 , \i_MIPS/Register/n758 ,
         \i_MIPS/Register/n757 , \i_MIPS/Register/n756 ,
         \i_MIPS/Register/n755 , \i_MIPS/Register/n754 ,
         \i_MIPS/Register/n753 , \i_MIPS/Register/n752 ,
         \i_MIPS/Register/n751 , \i_MIPS/Register/n750 ,
         \i_MIPS/Register/n749 , \i_MIPS/Register/n748 ,
         \i_MIPS/Register/n747 , \i_MIPS/Register/n746 ,
         \i_MIPS/Register/n745 , \i_MIPS/Register/n744 ,
         \i_MIPS/Register/n743 , \i_MIPS/Register/n742 ,
         \i_MIPS/Register/n741 , \i_MIPS/Register/n740 ,
         \i_MIPS/Register/n739 , \i_MIPS/Register/n738 ,
         \i_MIPS/Register/n737 , \i_MIPS/Register/n736 ,
         \i_MIPS/Register/n735 , \i_MIPS/Register/n734 ,
         \i_MIPS/Register/n733 , \i_MIPS/Register/n732 ,
         \i_MIPS/Register/n731 , \i_MIPS/Register/n730 ,
         \i_MIPS/Register/n729 , \i_MIPS/Register/n728 ,
         \i_MIPS/Register/n727 , \i_MIPS/Register/n726 ,
         \i_MIPS/Register/n725 , \i_MIPS/Register/n724 ,
         \i_MIPS/Register/n723 , \i_MIPS/Register/n722 ,
         \i_MIPS/Register/n721 , \i_MIPS/Register/n720 ,
         \i_MIPS/Register/n719 , \i_MIPS/Register/n718 ,
         \i_MIPS/Register/n717 , \i_MIPS/Register/n716 ,
         \i_MIPS/Register/n715 , \i_MIPS/Register/n714 ,
         \i_MIPS/Register/n713 , \i_MIPS/Register/n712 ,
         \i_MIPS/Register/n711 , \i_MIPS/Register/n710 ,
         \i_MIPS/Register/n709 , \i_MIPS/Register/n708 ,
         \i_MIPS/Register/n707 , \i_MIPS/Register/n706 ,
         \i_MIPS/Register/n705 , \i_MIPS/Register/n704 ,
         \i_MIPS/Register/n703 , \i_MIPS/Register/n702 ,
         \i_MIPS/Register/n701 , \i_MIPS/Register/n700 ,
         \i_MIPS/Register/n699 , \i_MIPS/Register/n698 ,
         \i_MIPS/Register/n697 , \i_MIPS/Register/n696 ,
         \i_MIPS/Register/n695 , \i_MIPS/Register/n694 ,
         \i_MIPS/Register/n693 , \i_MIPS/Register/n692 ,
         \i_MIPS/Register/n691 , \i_MIPS/Register/n690 ,
         \i_MIPS/Register/n689 , \i_MIPS/Register/n688 ,
         \i_MIPS/Register/n687 , \i_MIPS/Register/n686 ,
         \i_MIPS/Register/n685 , \i_MIPS/Register/n684 ,
         \i_MIPS/Register/n683 , \i_MIPS/Register/n682 ,
         \i_MIPS/Register/n681 , \i_MIPS/Register/n680 ,
         \i_MIPS/Register/n679 , \i_MIPS/Register/n678 ,
         \i_MIPS/Register/n677 , \i_MIPS/Register/n676 ,
         \i_MIPS/Register/n675 , \i_MIPS/Register/n674 ,
         \i_MIPS/Register/n673 , \i_MIPS/Register/n672 ,
         \i_MIPS/Register/n671 , \i_MIPS/Register/n670 ,
         \i_MIPS/Register/n669 , \i_MIPS/Register/n668 ,
         \i_MIPS/Register/n667 , \i_MIPS/Register/n666 ,
         \i_MIPS/Register/n665 , \i_MIPS/Register/n664 ,
         \i_MIPS/Register/n663 , \i_MIPS/Register/n662 ,
         \i_MIPS/Register/n661 , \i_MIPS/Register/n660 ,
         \i_MIPS/Register/n659 , \i_MIPS/Register/n658 ,
         \i_MIPS/Register/n657 , \i_MIPS/Register/n656 ,
         \i_MIPS/Register/n655 , \i_MIPS/Register/n654 ,
         \i_MIPS/Register/n653 , \i_MIPS/Register/n652 ,
         \i_MIPS/Register/n651 , \i_MIPS/Register/n650 ,
         \i_MIPS/Register/n649 , \i_MIPS/Register/n648 ,
         \i_MIPS/Register/n647 , \i_MIPS/Register/n646 ,
         \i_MIPS/Register/n645 , \i_MIPS/Register/n644 ,
         \i_MIPS/Register/n643 , \i_MIPS/Register/n642 ,
         \i_MIPS/Register/n641 , \i_MIPS/Register/n640 ,
         \i_MIPS/Register/n639 , \i_MIPS/Register/n638 ,
         \i_MIPS/Register/n637 , \i_MIPS/Register/n636 ,
         \i_MIPS/Register/n635 , \i_MIPS/Register/n634 ,
         \i_MIPS/Register/n633 , \i_MIPS/Register/n632 ,
         \i_MIPS/Register/n631 , \i_MIPS/Register/n630 ,
         \i_MIPS/Register/n629 , \i_MIPS/Register/n628 ,
         \i_MIPS/Register/n627 , \i_MIPS/Register/n626 ,
         \i_MIPS/Register/n625 , \i_MIPS/Register/n624 ,
         \i_MIPS/Register/n623 , \i_MIPS/Register/n622 ,
         \i_MIPS/Register/n621 , \i_MIPS/Register/n620 ,
         \i_MIPS/Register/n619 , \i_MIPS/Register/n618 ,
         \i_MIPS/Register/n617 , \i_MIPS/Register/n616 ,
         \i_MIPS/Register/n615 , \i_MIPS/Register/n614 ,
         \i_MIPS/Register/n613 , \i_MIPS/Register/n612 ,
         \i_MIPS/Register/n611 , \i_MIPS/Register/n610 ,
         \i_MIPS/Register/n609 , \i_MIPS/Register/n608 ,
         \i_MIPS/Register/n607 , \i_MIPS/Register/n606 ,
         \i_MIPS/Register/n605 , \i_MIPS/Register/n604 ,
         \i_MIPS/Register/n603 , \i_MIPS/Register/n602 ,
         \i_MIPS/Register/n601 , \i_MIPS/Register/n600 ,
         \i_MIPS/Register/n599 , \i_MIPS/Register/n598 ,
         \i_MIPS/Register/n597 , \i_MIPS/Register/n596 ,
         \i_MIPS/Register/n595 , \i_MIPS/Register/n594 ,
         \i_MIPS/Register/n593 , \i_MIPS/Register/n592 ,
         \i_MIPS/Register/n591 , \i_MIPS/Register/n590 ,
         \i_MIPS/Register/n589 , \i_MIPS/Register/n588 ,
         \i_MIPS/Register/n587 , \i_MIPS/Register/n586 ,
         \i_MIPS/Register/n585 , \i_MIPS/Register/n584 ,
         \i_MIPS/Register/n583 , \i_MIPS/Register/n582 ,
         \i_MIPS/Register/n581 , \i_MIPS/Register/n580 ,
         \i_MIPS/Register/n579 , \i_MIPS/Register/n578 ,
         \i_MIPS/Register/n577 , \i_MIPS/Register/n576 ,
         \i_MIPS/Register/n575 , \i_MIPS/Register/n574 ,
         \i_MIPS/Register/n573 , \i_MIPS/Register/n572 ,
         \i_MIPS/Register/n571 , \i_MIPS/Register/n570 ,
         \i_MIPS/Register/n569 , \i_MIPS/Register/n568 ,
         \i_MIPS/Register/n567 , \i_MIPS/Register/n566 ,
         \i_MIPS/Register/n565 , \i_MIPS/Register/n564 ,
         \i_MIPS/Register/n563 , \i_MIPS/Register/n562 ,
         \i_MIPS/Register/n561 , \i_MIPS/Register/n560 ,
         \i_MIPS/Register/n559 , \i_MIPS/Register/n558 ,
         \i_MIPS/Register/n557 , \i_MIPS/Register/n556 ,
         \i_MIPS/Register/n555 , \i_MIPS/Register/n554 ,
         \i_MIPS/Register/n553 , \i_MIPS/Register/n552 ,
         \i_MIPS/Register/n551 , \i_MIPS/Register/n550 ,
         \i_MIPS/Register/n549 , \i_MIPS/Register/n548 ,
         \i_MIPS/Register/n547 , \i_MIPS/Register/n546 ,
         \i_MIPS/Register/n545 , \i_MIPS/Register/n544 ,
         \i_MIPS/Register/n543 , \i_MIPS/Register/n542 ,
         \i_MIPS/Register/n541 , \i_MIPS/Register/n540 ,
         \i_MIPS/Register/n539 , \i_MIPS/Register/n538 ,
         \i_MIPS/Register/n537 , \i_MIPS/Register/n536 ,
         \i_MIPS/Register/n535 , \i_MIPS/Register/n534 ,
         \i_MIPS/Register/n533 , \i_MIPS/Register/n532 ,
         \i_MIPS/Register/n531 , \i_MIPS/Register/n530 ,
         \i_MIPS/Register/n529 , \i_MIPS/Register/n528 ,
         \i_MIPS/Register/n527 , \i_MIPS/Register/n526 ,
         \i_MIPS/Register/n525 , \i_MIPS/Register/n524 ,
         \i_MIPS/Register/n523 , \i_MIPS/Register/n522 ,
         \i_MIPS/Register/n521 , \i_MIPS/Register/n520 ,
         \i_MIPS/Register/n519 , \i_MIPS/Register/n518 ,
         \i_MIPS/Register/n517 , \i_MIPS/Register/n516 ,
         \i_MIPS/Register/n515 , \i_MIPS/Register/n514 ,
         \i_MIPS/Register/n513 , \i_MIPS/Register/n512 ,
         \i_MIPS/Register/n511 , \i_MIPS/Register/n510 ,
         \i_MIPS/Register/n509 , \i_MIPS/Register/n508 ,
         \i_MIPS/Register/n507 , \i_MIPS/Register/n506 ,
         \i_MIPS/Register/n505 , \i_MIPS/Register/n504 ,
         \i_MIPS/Register/n503 , \i_MIPS/Register/n502 ,
         \i_MIPS/Register/n501 , \i_MIPS/Register/n500 ,
         \i_MIPS/Register/n499 , \i_MIPS/Register/n498 ,
         \i_MIPS/Register/n497 , \i_MIPS/Register/n496 ,
         \i_MIPS/Register/n495 , \i_MIPS/Register/n494 ,
         \i_MIPS/Register/n493 , \i_MIPS/Register/n492 ,
         \i_MIPS/Register/n491 , \i_MIPS/Register/n490 ,
         \i_MIPS/Register/n489 , \i_MIPS/Register/n488 ,
         \i_MIPS/Register/n487 , \i_MIPS/Register/n486 ,
         \i_MIPS/Register/n485 , \i_MIPS/Register/n484 ,
         \i_MIPS/Register/n483 , \i_MIPS/Register/n482 ,
         \i_MIPS/Register/n481 , \i_MIPS/Register/n480 ,
         \i_MIPS/Register/n479 , \i_MIPS/Register/n478 ,
         \i_MIPS/Register/n477 , \i_MIPS/Register/n476 ,
         \i_MIPS/Register/n475 , \i_MIPS/Register/n474 ,
         \i_MIPS/Register/n473 , \i_MIPS/Register/n472 ,
         \i_MIPS/Register/n471 , \i_MIPS/Register/n470 ,
         \i_MIPS/Register/n469 , \i_MIPS/Register/n468 ,
         \i_MIPS/Register/n467 , \i_MIPS/Register/n466 ,
         \i_MIPS/Register/n465 , \i_MIPS/Register/n464 ,
         \i_MIPS/Register/n463 , \i_MIPS/Register/n462 ,
         \i_MIPS/Register/n461 , \i_MIPS/Register/n460 ,
         \i_MIPS/Register/n459 , \i_MIPS/Register/n458 ,
         \i_MIPS/Register/n457 , \i_MIPS/Register/n456 ,
         \i_MIPS/Register/n455 , \i_MIPS/Register/n454 ,
         \i_MIPS/Register/n453 , \i_MIPS/Register/n452 ,
         \i_MIPS/Register/n451 , \i_MIPS/Register/n450 ,
         \i_MIPS/Register/n449 , \i_MIPS/Register/n448 ,
         \i_MIPS/Register/n447 , \i_MIPS/Register/n446 ,
         \i_MIPS/Register/n445 , \i_MIPS/Register/n444 ,
         \i_MIPS/Register/n443 , \i_MIPS/Register/n442 ,
         \i_MIPS/Register/n441 , \i_MIPS/Register/n440 ,
         \i_MIPS/Register/n439 , \i_MIPS/Register/n438 ,
         \i_MIPS/Register/n437 , \i_MIPS/Register/n436 ,
         \i_MIPS/Register/n435 , \i_MIPS/Register/n434 ,
         \i_MIPS/Register/n433 , \i_MIPS/Register/n432 ,
         \i_MIPS/Register/n431 , \i_MIPS/Register/n430 ,
         \i_MIPS/Register/n429 , \i_MIPS/Register/n428 ,
         \i_MIPS/Register/n427 , \i_MIPS/Register/n426 ,
         \i_MIPS/Register/n425 , \i_MIPS/Register/n424 ,
         \i_MIPS/Register/n423 , \i_MIPS/Register/n422 ,
         \i_MIPS/Register/n421 , \i_MIPS/Register/n420 ,
         \i_MIPS/Register/n419 , \i_MIPS/Register/n418 ,
         \i_MIPS/Register/n417 , \i_MIPS/Register/n416 ,
         \i_MIPS/Register/n415 , \i_MIPS/Register/n414 ,
         \i_MIPS/Register/n413 , \i_MIPS/Register/n412 ,
         \i_MIPS/Register/n411 , \i_MIPS/Register/n410 ,
         \i_MIPS/Register/n409 , \i_MIPS/Register/n408 ,
         \i_MIPS/Register/n407 , \i_MIPS/Register/n406 ,
         \i_MIPS/Register/n405 , \i_MIPS/Register/n404 ,
         \i_MIPS/Register/n403 , \i_MIPS/Register/n402 ,
         \i_MIPS/Register/n401 , \i_MIPS/Register/n400 ,
         \i_MIPS/Register/n399 , \i_MIPS/Register/n398 ,
         \i_MIPS/Register/n397 , \i_MIPS/Register/n396 ,
         \i_MIPS/Register/n395 , \i_MIPS/Register/n394 ,
         \i_MIPS/Register/n393 , \i_MIPS/Register/n392 ,
         \i_MIPS/Register/n391 , \i_MIPS/Register/n390 ,
         \i_MIPS/Register/n389 , \i_MIPS/Register/n388 ,
         \i_MIPS/Register/n387 , \i_MIPS/Register/n386 ,
         \i_MIPS/Register/n385 , \i_MIPS/Register/n384 ,
         \i_MIPS/Register/n383 , \i_MIPS/Register/n382 ,
         \i_MIPS/Register/n381 , \i_MIPS/Register/n380 ,
         \i_MIPS/Register/n379 , \i_MIPS/Register/n378 ,
         \i_MIPS/Register/n377 , \i_MIPS/Register/n376 ,
         \i_MIPS/Register/n375 , \i_MIPS/Register/n374 ,
         \i_MIPS/Register/n373 , \i_MIPS/Register/n372 ,
         \i_MIPS/Register/n371 , \i_MIPS/Register/n370 ,
         \i_MIPS/Register/n369 , \i_MIPS/Register/n368 ,
         \i_MIPS/Register/n367 , \i_MIPS/Register/n366 ,
         \i_MIPS/Register/n365 , \i_MIPS/Register/n364 ,
         \i_MIPS/Register/n363 , \i_MIPS/Register/n362 ,
         \i_MIPS/Register/n361 , \i_MIPS/Register/n360 ,
         \i_MIPS/Register/n359 , \i_MIPS/Register/n358 ,
         \i_MIPS/Register/n357 , \i_MIPS/Register/n356 ,
         \i_MIPS/Register/n355 , \i_MIPS/Register/n354 ,
         \i_MIPS/Register/n353 , \i_MIPS/Register/n352 ,
         \i_MIPS/Register/n351 , \i_MIPS/Register/n350 ,
         \i_MIPS/Register/n349 , \i_MIPS/Register/n348 ,
         \i_MIPS/Register/n347 , \i_MIPS/Register/n346 ,
         \i_MIPS/Register/n345 , \i_MIPS/Register/n344 ,
         \i_MIPS/Register/n343 , \i_MIPS/Register/n342 ,
         \i_MIPS/Register/n341 , \i_MIPS/Register/n340 ,
         \i_MIPS/Register/n339 , \i_MIPS/Register/n338 ,
         \i_MIPS/Register/n337 , \i_MIPS/Register/n336 ,
         \i_MIPS/Register/n335 , \i_MIPS/Register/n334 ,
         \i_MIPS/Register/n333 , \i_MIPS/Register/n332 ,
         \i_MIPS/Register/n331 , \i_MIPS/Register/n330 ,
         \i_MIPS/Register/n329 , \i_MIPS/Register/n328 ,
         \i_MIPS/Register/n327 , \i_MIPS/Register/n326 ,
         \i_MIPS/Register/n325 , \i_MIPS/Register/n324 ,
         \i_MIPS/Register/n323 , \i_MIPS/Register/n322 ,
         \i_MIPS/Register/n321 , \i_MIPS/Register/n320 ,
         \i_MIPS/Register/n319 , \i_MIPS/Register/n318 ,
         \i_MIPS/Register/n317 , \i_MIPS/Register/n316 ,
         \i_MIPS/Register/n315 , \i_MIPS/Register/n314 ,
         \i_MIPS/Register/n313 , \i_MIPS/Register/n312 ,
         \i_MIPS/Register/n311 , \i_MIPS/Register/n310 ,
         \i_MIPS/Register/n309 , \i_MIPS/Register/n308 ,
         \i_MIPS/Register/n307 , \i_MIPS/Register/n306 ,
         \i_MIPS/Register/n305 , \i_MIPS/Register/n304 ,
         \i_MIPS/Register/n303 , \i_MIPS/Register/n302 ,
         \i_MIPS/Register/n301 , \i_MIPS/Register/n300 ,
         \i_MIPS/Register/n299 , \i_MIPS/Register/n298 ,
         \i_MIPS/Register/n297 , \i_MIPS/Register/n296 ,
         \i_MIPS/Register/n295 , \i_MIPS/Register/n294 ,
         \i_MIPS/Register/n293 , \i_MIPS/Register/n292 ,
         \i_MIPS/Register/n291 , \i_MIPS/Register/n290 ,
         \i_MIPS/Register/n289 , \i_MIPS/Register/n288 ,
         \i_MIPS/Register/n287 , \i_MIPS/Register/n286 ,
         \i_MIPS/Register/n285 , \i_MIPS/Register/n284 ,
         \i_MIPS/Register/n283 , \i_MIPS/Register/n282 ,
         \i_MIPS/Register/n281 , \i_MIPS/Register/n280 ,
         \i_MIPS/Register/n279 , \i_MIPS/Register/n278 ,
         \i_MIPS/Register/n277 , \i_MIPS/Register/n276 ,
         \i_MIPS/Register/n275 , \i_MIPS/Register/n274 ,
         \i_MIPS/Register/n273 , \i_MIPS/Register/n272 ,
         \i_MIPS/Register/n271 , \i_MIPS/Register/n270 ,
         \i_MIPS/Register/n269 , \i_MIPS/Register/n268 ,
         \i_MIPS/Register/n267 , \i_MIPS/Register/n266 ,
         \i_MIPS/Register/n265 , \i_MIPS/Register/n264 ,
         \i_MIPS/Register/n263 , \i_MIPS/Register/n262 ,
         \i_MIPS/Register/n261 , \i_MIPS/Register/n260 ,
         \i_MIPS/Register/n259 , \i_MIPS/Register/n258 ,
         \i_MIPS/Register/n257 , \i_MIPS/Register/n256 ,
         \i_MIPS/Register/n255 , \i_MIPS/Register/n254 ,
         \i_MIPS/Register/n253 , \i_MIPS/Register/n252 ,
         \i_MIPS/Register/n251 , \i_MIPS/Register/n250 ,
         \i_MIPS/Register/n249 , \i_MIPS/Register/n248 ,
         \i_MIPS/Register/n247 , \i_MIPS/Register/n246 ,
         \i_MIPS/Register/n245 , \i_MIPS/Register/n244 ,
         \i_MIPS/Register/n243 , \i_MIPS/Register/n242 ,
         \i_MIPS/Register/n241 , \i_MIPS/Register/n240 ,
         \i_MIPS/Register/n239 , \i_MIPS/Register/n238 ,
         \i_MIPS/Register/n237 , \i_MIPS/Register/n236 ,
         \i_MIPS/Register/n235 , \i_MIPS/Register/n234 ,
         \i_MIPS/Register/n233 , \i_MIPS/Register/n232 ,
         \i_MIPS/Register/n231 , \i_MIPS/Register/n230 ,
         \i_MIPS/Register/n229 , \i_MIPS/Register/n228 ,
         \i_MIPS/Register/n227 , \i_MIPS/Register/n226 ,
         \i_MIPS/Register/n225 , \i_MIPS/Register/n224 ,
         \i_MIPS/Register/n223 , \i_MIPS/Register/n222 ,
         \i_MIPS/Register/n221 , \i_MIPS/Register/n220 ,
         \i_MIPS/Register/n219 , \i_MIPS/Register/n218 ,
         \i_MIPS/Register/n217 , \i_MIPS/Register/n216 ,
         \i_MIPS/Register/n215 , \i_MIPS/Register/n214 ,
         \i_MIPS/Register/n213 , \i_MIPS/Register/n212 ,
         \i_MIPS/Register/n211 , \i_MIPS/Register/n210 ,
         \i_MIPS/Register/n209 , \i_MIPS/Register/n208 ,
         \i_MIPS/Register/n207 , \i_MIPS/Register/n206 ,
         \i_MIPS/Register/n205 , \i_MIPS/Register/n204 ,
         \i_MIPS/Register/n203 , \i_MIPS/Register/n202 ,
         \i_MIPS/Register/n201 , \i_MIPS/Register/n200 ,
         \i_MIPS/Register/n199 , \i_MIPS/Register/n198 ,
         \i_MIPS/Register/n197 , \i_MIPS/Register/n196 ,
         \i_MIPS/Register/n195 , \i_MIPS/Register/n194 ,
         \i_MIPS/Register/n193 , \i_MIPS/Register/n192 ,
         \i_MIPS/Register/n191 , \i_MIPS/Register/n190 ,
         \i_MIPS/Register/n189 , \i_MIPS/Register/n188 ,
         \i_MIPS/Register/n187 , \i_MIPS/Register/n186 ,
         \i_MIPS/Register/n185 , \i_MIPS/Register/n184 ,
         \i_MIPS/Register/n183 , \i_MIPS/Register/n182 ,
         \i_MIPS/Register/n181 , \i_MIPS/Register/n180 ,
         \i_MIPS/Register/n179 , \i_MIPS/Register/n178 ,
         \i_MIPS/Register/n177 , \i_MIPS/Register/n176 ,
         \i_MIPS/Register/n175 , \i_MIPS/Register/n174 ,
         \i_MIPS/Register/n173 , \i_MIPS/Register/n172 ,
         \i_MIPS/Register/n171 , \i_MIPS/Register/n170 ,
         \i_MIPS/Register/n169 , \i_MIPS/Register/n168 ,
         \i_MIPS/Register/n167 , \i_MIPS/Register/n166 ,
         \i_MIPS/Register/n165 , \i_MIPS/Register/n164 ,
         \i_MIPS/Register/n163 , \i_MIPS/Register/n162 ,
         \i_MIPS/Register/n161 , \i_MIPS/Register/n160 ,
         \i_MIPS/Register/n159 , \i_MIPS/Register/n158 ,
         \i_MIPS/Register/n157 , \i_MIPS/Register/n156 ,
         \i_MIPS/Register/n155 , \i_MIPS/Register/n154 ,
         \i_MIPS/Register/n153 , \i_MIPS/Register/n152 ,
         \i_MIPS/Register/n151 , \i_MIPS/Register/n150 ,
         \i_MIPS/Register/n149 , \i_MIPS/Register/n148 ,
         \i_MIPS/Register/n140 , \i_MIPS/Register/n131 ,
         \i_MIPS/Register/n122 , \i_MIPS/Register/n120 ,
         \i_MIPS/Register/n119 , \i_MIPS/Register/n118 ,
         \i_MIPS/Register/n117 , \i_MIPS/Register/n116 ,
         \i_MIPS/Register/n115 , \i_MIPS/Register/n114 ,
         \i_MIPS/Register/n113 , \i_MIPS/Register/n112 ,
         \i_MIPS/Register/n111 , \i_MIPS/Register/n110 ,
         \i_MIPS/Register/n109 , \i_MIPS/Register/n108 ,
         \i_MIPS/Register/n107 , \i_MIPS/Register/n106 ,
         \i_MIPS/Register/n105 , \i_MIPS/Register/n104 ,
         \i_MIPS/Register/register[30][0] , \i_MIPS/Register/register[30][1] ,
         \i_MIPS/Register/register[30][2] , \i_MIPS/Register/register[30][3] ,
         \i_MIPS/Register/register[30][4] , \i_MIPS/Register/register[30][5] ,
         \i_MIPS/Register/register[30][6] , \i_MIPS/Register/register[30][7] ,
         \i_MIPS/Register/register[30][8] , \i_MIPS/Register/register[30][9] ,
         \i_MIPS/Register/register[30][10] ,
         \i_MIPS/Register/register[30][11] ,
         \i_MIPS/Register/register[30][12] ,
         \i_MIPS/Register/register[30][13] ,
         \i_MIPS/Register/register[30][14] ,
         \i_MIPS/Register/register[30][15] ,
         \i_MIPS/Register/register[30][16] ,
         \i_MIPS/Register/register[30][17] ,
         \i_MIPS/Register/register[30][18] ,
         \i_MIPS/Register/register[30][19] ,
         \i_MIPS/Register/register[30][20] ,
         \i_MIPS/Register/register[30][21] ,
         \i_MIPS/Register/register[30][22] ,
         \i_MIPS/Register/register[30][23] ,
         \i_MIPS/Register/register[30][24] ,
         \i_MIPS/Register/register[30][25] ,
         \i_MIPS/Register/register[30][26] ,
         \i_MIPS/Register/register[30][27] ,
         \i_MIPS/Register/register[30][28] ,
         \i_MIPS/Register/register[30][29] ,
         \i_MIPS/Register/register[30][30] ,
         \i_MIPS/Register/register[30][31] , \i_MIPS/Register/register[29][0] ,
         \i_MIPS/Register/register[29][1] , \i_MIPS/Register/register[29][2] ,
         \i_MIPS/Register/register[29][3] , \i_MIPS/Register/register[29][4] ,
         \i_MIPS/Register/register[29][5] , \i_MIPS/Register/register[29][6] ,
         \i_MIPS/Register/register[29][7] , \i_MIPS/Register/register[29][8] ,
         \i_MIPS/Register/register[29][9] , \i_MIPS/Register/register[29][10] ,
         \i_MIPS/Register/register[29][11] ,
         \i_MIPS/Register/register[29][12] ,
         \i_MIPS/Register/register[29][13] ,
         \i_MIPS/Register/register[29][14] ,
         \i_MIPS/Register/register[29][15] ,
         \i_MIPS/Register/register[29][16] ,
         \i_MIPS/Register/register[29][17] ,
         \i_MIPS/Register/register[29][18] ,
         \i_MIPS/Register/register[29][19] ,
         \i_MIPS/Register/register[29][20] ,
         \i_MIPS/Register/register[29][21] ,
         \i_MIPS/Register/register[29][22] ,
         \i_MIPS/Register/register[29][23] ,
         \i_MIPS/Register/register[29][24] ,
         \i_MIPS/Register/register[29][25] ,
         \i_MIPS/Register/register[29][26] ,
         \i_MIPS/Register/register[29][27] ,
         \i_MIPS/Register/register[29][28] ,
         \i_MIPS/Register/register[29][29] ,
         \i_MIPS/Register/register[29][30] ,
         \i_MIPS/Register/register[29][31] , \i_MIPS/Register/register[28][0] ,
         \i_MIPS/Register/register[28][1] , \i_MIPS/Register/register[28][2] ,
         \i_MIPS/Register/register[28][3] , \i_MIPS/Register/register[28][4] ,
         \i_MIPS/Register/register[28][5] , \i_MIPS/Register/register[28][6] ,
         \i_MIPS/Register/register[28][7] , \i_MIPS/Register/register[28][8] ,
         \i_MIPS/Register/register[28][9] , \i_MIPS/Register/register[28][10] ,
         \i_MIPS/Register/register[28][11] ,
         \i_MIPS/Register/register[28][12] ,
         \i_MIPS/Register/register[28][13] ,
         \i_MIPS/Register/register[28][14] ,
         \i_MIPS/Register/register[28][15] ,
         \i_MIPS/Register/register[28][16] ,
         \i_MIPS/Register/register[28][17] ,
         \i_MIPS/Register/register[28][18] ,
         \i_MIPS/Register/register[28][19] ,
         \i_MIPS/Register/register[28][20] ,
         \i_MIPS/Register/register[28][21] ,
         \i_MIPS/Register/register[28][22] ,
         \i_MIPS/Register/register[28][23] ,
         \i_MIPS/Register/register[28][24] ,
         \i_MIPS/Register/register[28][25] ,
         \i_MIPS/Register/register[28][26] ,
         \i_MIPS/Register/register[28][27] ,
         \i_MIPS/Register/register[28][28] ,
         \i_MIPS/Register/register[28][29] ,
         \i_MIPS/Register/register[28][30] ,
         \i_MIPS/Register/register[28][31] , \i_MIPS/Register/register[27][0] ,
         \i_MIPS/Register/register[27][1] , \i_MIPS/Register/register[27][2] ,
         \i_MIPS/Register/register[27][3] , \i_MIPS/Register/register[27][4] ,
         \i_MIPS/Register/register[27][5] , \i_MIPS/Register/register[27][6] ,
         \i_MIPS/Register/register[27][7] , \i_MIPS/Register/register[27][8] ,
         \i_MIPS/Register/register[27][9] , \i_MIPS/Register/register[27][10] ,
         \i_MIPS/Register/register[27][11] ,
         \i_MIPS/Register/register[27][12] ,
         \i_MIPS/Register/register[27][13] ,
         \i_MIPS/Register/register[27][14] ,
         \i_MIPS/Register/register[27][15] ,
         \i_MIPS/Register/register[27][16] ,
         \i_MIPS/Register/register[27][17] ,
         \i_MIPS/Register/register[27][18] ,
         \i_MIPS/Register/register[27][19] ,
         \i_MIPS/Register/register[27][20] ,
         \i_MIPS/Register/register[27][21] ,
         \i_MIPS/Register/register[27][22] ,
         \i_MIPS/Register/register[27][23] ,
         \i_MIPS/Register/register[27][24] ,
         \i_MIPS/Register/register[27][25] ,
         \i_MIPS/Register/register[27][26] ,
         \i_MIPS/Register/register[27][27] ,
         \i_MIPS/Register/register[27][28] ,
         \i_MIPS/Register/register[27][29] ,
         \i_MIPS/Register/register[27][30] ,
         \i_MIPS/Register/register[27][31] , \i_MIPS/Register/register[26][0] ,
         \i_MIPS/Register/register[26][1] , \i_MIPS/Register/register[26][2] ,
         \i_MIPS/Register/register[26][3] , \i_MIPS/Register/register[26][4] ,
         \i_MIPS/Register/register[26][5] , \i_MIPS/Register/register[26][6] ,
         \i_MIPS/Register/register[26][7] , \i_MIPS/Register/register[26][8] ,
         \i_MIPS/Register/register[26][9] , \i_MIPS/Register/register[26][10] ,
         \i_MIPS/Register/register[26][11] ,
         \i_MIPS/Register/register[26][12] ,
         \i_MIPS/Register/register[26][13] ,
         \i_MIPS/Register/register[26][14] ,
         \i_MIPS/Register/register[26][15] ,
         \i_MIPS/Register/register[26][16] ,
         \i_MIPS/Register/register[26][17] ,
         \i_MIPS/Register/register[26][18] ,
         \i_MIPS/Register/register[26][19] ,
         \i_MIPS/Register/register[26][20] ,
         \i_MIPS/Register/register[26][21] ,
         \i_MIPS/Register/register[26][22] ,
         \i_MIPS/Register/register[26][23] ,
         \i_MIPS/Register/register[26][24] ,
         \i_MIPS/Register/register[26][25] ,
         \i_MIPS/Register/register[26][26] ,
         \i_MIPS/Register/register[26][27] ,
         \i_MIPS/Register/register[26][28] ,
         \i_MIPS/Register/register[26][29] ,
         \i_MIPS/Register/register[26][30] ,
         \i_MIPS/Register/register[26][31] , \i_MIPS/Register/register[25][0] ,
         \i_MIPS/Register/register[25][1] , \i_MIPS/Register/register[25][2] ,
         \i_MIPS/Register/register[25][3] , \i_MIPS/Register/register[25][4] ,
         \i_MIPS/Register/register[25][5] , \i_MIPS/Register/register[25][6] ,
         \i_MIPS/Register/register[25][7] , \i_MIPS/Register/register[25][8] ,
         \i_MIPS/Register/register[25][9] , \i_MIPS/Register/register[25][10] ,
         \i_MIPS/Register/register[25][11] ,
         \i_MIPS/Register/register[25][12] ,
         \i_MIPS/Register/register[25][13] ,
         \i_MIPS/Register/register[25][14] ,
         \i_MIPS/Register/register[25][15] ,
         \i_MIPS/Register/register[25][16] ,
         \i_MIPS/Register/register[25][17] ,
         \i_MIPS/Register/register[25][18] ,
         \i_MIPS/Register/register[25][19] ,
         \i_MIPS/Register/register[25][20] ,
         \i_MIPS/Register/register[25][21] ,
         \i_MIPS/Register/register[25][22] ,
         \i_MIPS/Register/register[25][23] ,
         \i_MIPS/Register/register[25][24] ,
         \i_MIPS/Register/register[25][25] ,
         \i_MIPS/Register/register[25][26] ,
         \i_MIPS/Register/register[25][27] ,
         \i_MIPS/Register/register[25][28] ,
         \i_MIPS/Register/register[25][29] ,
         \i_MIPS/Register/register[25][30] ,
         \i_MIPS/Register/register[25][31] , \i_MIPS/Register/register[24][0] ,
         \i_MIPS/Register/register[24][1] , \i_MIPS/Register/register[24][2] ,
         \i_MIPS/Register/register[24][3] , \i_MIPS/Register/register[24][4] ,
         \i_MIPS/Register/register[24][5] , \i_MIPS/Register/register[24][6] ,
         \i_MIPS/Register/register[24][7] , \i_MIPS/Register/register[24][8] ,
         \i_MIPS/Register/register[24][9] , \i_MIPS/Register/register[24][10] ,
         \i_MIPS/Register/register[24][11] ,
         \i_MIPS/Register/register[24][12] ,
         \i_MIPS/Register/register[24][13] ,
         \i_MIPS/Register/register[24][14] ,
         \i_MIPS/Register/register[24][15] ,
         \i_MIPS/Register/register[24][16] ,
         \i_MIPS/Register/register[24][17] ,
         \i_MIPS/Register/register[24][18] ,
         \i_MIPS/Register/register[24][19] ,
         \i_MIPS/Register/register[24][20] ,
         \i_MIPS/Register/register[24][21] ,
         \i_MIPS/Register/register[24][22] ,
         \i_MIPS/Register/register[24][23] ,
         \i_MIPS/Register/register[24][24] ,
         \i_MIPS/Register/register[24][25] ,
         \i_MIPS/Register/register[24][26] ,
         \i_MIPS/Register/register[24][27] ,
         \i_MIPS/Register/register[24][28] ,
         \i_MIPS/Register/register[24][29] ,
         \i_MIPS/Register/register[24][30] ,
         \i_MIPS/Register/register[24][31] , \i_MIPS/Register/register[23][0] ,
         \i_MIPS/Register/register[23][1] , \i_MIPS/Register/register[23][2] ,
         \i_MIPS/Register/register[23][3] , \i_MIPS/Register/register[23][4] ,
         \i_MIPS/Register/register[23][5] , \i_MIPS/Register/register[23][6] ,
         \i_MIPS/Register/register[23][7] , \i_MIPS/Register/register[23][8] ,
         \i_MIPS/Register/register[23][9] , \i_MIPS/Register/register[23][10] ,
         \i_MIPS/Register/register[23][11] ,
         \i_MIPS/Register/register[23][12] ,
         \i_MIPS/Register/register[23][13] ,
         \i_MIPS/Register/register[23][14] ,
         \i_MIPS/Register/register[23][15] ,
         \i_MIPS/Register/register[23][16] ,
         \i_MIPS/Register/register[23][17] ,
         \i_MIPS/Register/register[23][18] ,
         \i_MIPS/Register/register[23][19] ,
         \i_MIPS/Register/register[23][20] ,
         \i_MIPS/Register/register[23][21] ,
         \i_MIPS/Register/register[23][22] ,
         \i_MIPS/Register/register[23][23] ,
         \i_MIPS/Register/register[23][24] ,
         \i_MIPS/Register/register[23][25] ,
         \i_MIPS/Register/register[23][26] ,
         \i_MIPS/Register/register[23][27] ,
         \i_MIPS/Register/register[23][28] ,
         \i_MIPS/Register/register[23][29] ,
         \i_MIPS/Register/register[23][30] ,
         \i_MIPS/Register/register[23][31] , \i_MIPS/Register/register[22][0] ,
         \i_MIPS/Register/register[22][1] , \i_MIPS/Register/register[22][2] ,
         \i_MIPS/Register/register[22][3] , \i_MIPS/Register/register[22][4] ,
         \i_MIPS/Register/register[22][5] , \i_MIPS/Register/register[22][6] ,
         \i_MIPS/Register/register[22][7] , \i_MIPS/Register/register[22][8] ,
         \i_MIPS/Register/register[22][9] , \i_MIPS/Register/register[22][10] ,
         \i_MIPS/Register/register[22][11] ,
         \i_MIPS/Register/register[22][12] ,
         \i_MIPS/Register/register[22][13] ,
         \i_MIPS/Register/register[22][14] ,
         \i_MIPS/Register/register[22][15] ,
         \i_MIPS/Register/register[22][16] ,
         \i_MIPS/Register/register[22][17] ,
         \i_MIPS/Register/register[22][18] ,
         \i_MIPS/Register/register[22][19] ,
         \i_MIPS/Register/register[22][20] ,
         \i_MIPS/Register/register[22][21] ,
         \i_MIPS/Register/register[22][22] ,
         \i_MIPS/Register/register[22][23] ,
         \i_MIPS/Register/register[22][24] ,
         \i_MIPS/Register/register[22][25] ,
         \i_MIPS/Register/register[22][26] ,
         \i_MIPS/Register/register[22][27] ,
         \i_MIPS/Register/register[22][28] ,
         \i_MIPS/Register/register[22][29] ,
         \i_MIPS/Register/register[22][30] ,
         \i_MIPS/Register/register[22][31] , \i_MIPS/Register/register[21][0] ,
         \i_MIPS/Register/register[21][1] , \i_MIPS/Register/register[21][2] ,
         \i_MIPS/Register/register[21][3] , \i_MIPS/Register/register[21][4] ,
         \i_MIPS/Register/register[21][5] , \i_MIPS/Register/register[21][6] ,
         \i_MIPS/Register/register[21][7] , \i_MIPS/Register/register[21][8] ,
         \i_MIPS/Register/register[21][9] , \i_MIPS/Register/register[21][10] ,
         \i_MIPS/Register/register[21][11] ,
         \i_MIPS/Register/register[21][12] ,
         \i_MIPS/Register/register[21][13] ,
         \i_MIPS/Register/register[21][14] ,
         \i_MIPS/Register/register[21][15] ,
         \i_MIPS/Register/register[21][16] ,
         \i_MIPS/Register/register[21][17] ,
         \i_MIPS/Register/register[21][18] ,
         \i_MIPS/Register/register[21][19] ,
         \i_MIPS/Register/register[21][20] ,
         \i_MIPS/Register/register[21][21] ,
         \i_MIPS/Register/register[21][22] ,
         \i_MIPS/Register/register[21][23] ,
         \i_MIPS/Register/register[21][24] ,
         \i_MIPS/Register/register[21][25] ,
         \i_MIPS/Register/register[21][26] ,
         \i_MIPS/Register/register[21][27] ,
         \i_MIPS/Register/register[21][28] ,
         \i_MIPS/Register/register[21][29] ,
         \i_MIPS/Register/register[21][30] ,
         \i_MIPS/Register/register[21][31] , \i_MIPS/Register/register[20][0] ,
         \i_MIPS/Register/register[20][1] , \i_MIPS/Register/register[20][2] ,
         \i_MIPS/Register/register[20][3] , \i_MIPS/Register/register[20][4] ,
         \i_MIPS/Register/register[20][5] , \i_MIPS/Register/register[20][6] ,
         \i_MIPS/Register/register[20][7] , \i_MIPS/Register/register[20][8] ,
         \i_MIPS/Register/register[20][9] , \i_MIPS/Register/register[20][10] ,
         \i_MIPS/Register/register[20][11] ,
         \i_MIPS/Register/register[20][12] ,
         \i_MIPS/Register/register[20][13] ,
         \i_MIPS/Register/register[20][14] ,
         \i_MIPS/Register/register[20][15] ,
         \i_MIPS/Register/register[20][16] ,
         \i_MIPS/Register/register[20][17] ,
         \i_MIPS/Register/register[20][18] ,
         \i_MIPS/Register/register[20][19] ,
         \i_MIPS/Register/register[20][20] ,
         \i_MIPS/Register/register[20][21] ,
         \i_MIPS/Register/register[20][22] ,
         \i_MIPS/Register/register[20][23] ,
         \i_MIPS/Register/register[20][24] ,
         \i_MIPS/Register/register[20][25] ,
         \i_MIPS/Register/register[20][26] ,
         \i_MIPS/Register/register[20][27] ,
         \i_MIPS/Register/register[20][28] ,
         \i_MIPS/Register/register[20][29] ,
         \i_MIPS/Register/register[20][30] ,
         \i_MIPS/Register/register[20][31] , \i_MIPS/Register/register[19][0] ,
         \i_MIPS/Register/register[19][1] , \i_MIPS/Register/register[19][2] ,
         \i_MIPS/Register/register[19][3] , \i_MIPS/Register/register[19][4] ,
         \i_MIPS/Register/register[19][5] , \i_MIPS/Register/register[19][6] ,
         \i_MIPS/Register/register[19][7] , \i_MIPS/Register/register[19][8] ,
         \i_MIPS/Register/register[19][9] , \i_MIPS/Register/register[19][10] ,
         \i_MIPS/Register/register[19][11] ,
         \i_MIPS/Register/register[19][12] ,
         \i_MIPS/Register/register[19][13] ,
         \i_MIPS/Register/register[19][14] ,
         \i_MIPS/Register/register[19][15] ,
         \i_MIPS/Register/register[19][16] ,
         \i_MIPS/Register/register[19][17] ,
         \i_MIPS/Register/register[19][18] ,
         \i_MIPS/Register/register[19][19] ,
         \i_MIPS/Register/register[19][20] ,
         \i_MIPS/Register/register[19][21] ,
         \i_MIPS/Register/register[19][22] ,
         \i_MIPS/Register/register[19][23] ,
         \i_MIPS/Register/register[19][24] ,
         \i_MIPS/Register/register[19][25] ,
         \i_MIPS/Register/register[19][26] ,
         \i_MIPS/Register/register[19][27] ,
         \i_MIPS/Register/register[19][28] ,
         \i_MIPS/Register/register[19][29] ,
         \i_MIPS/Register/register[19][30] ,
         \i_MIPS/Register/register[19][31] , \i_MIPS/Register/register[18][0] ,
         \i_MIPS/Register/register[18][1] , \i_MIPS/Register/register[18][2] ,
         \i_MIPS/Register/register[18][3] , \i_MIPS/Register/register[18][4] ,
         \i_MIPS/Register/register[18][5] , \i_MIPS/Register/register[18][6] ,
         \i_MIPS/Register/register[18][7] , \i_MIPS/Register/register[18][8] ,
         \i_MIPS/Register/register[18][9] , \i_MIPS/Register/register[18][10] ,
         \i_MIPS/Register/register[18][11] ,
         \i_MIPS/Register/register[18][12] ,
         \i_MIPS/Register/register[18][13] ,
         \i_MIPS/Register/register[18][14] ,
         \i_MIPS/Register/register[18][15] ,
         \i_MIPS/Register/register[18][16] ,
         \i_MIPS/Register/register[18][17] ,
         \i_MIPS/Register/register[18][18] ,
         \i_MIPS/Register/register[18][19] ,
         \i_MIPS/Register/register[18][20] ,
         \i_MIPS/Register/register[18][21] ,
         \i_MIPS/Register/register[18][22] ,
         \i_MIPS/Register/register[18][23] ,
         \i_MIPS/Register/register[18][24] ,
         \i_MIPS/Register/register[18][25] ,
         \i_MIPS/Register/register[18][26] ,
         \i_MIPS/Register/register[18][27] ,
         \i_MIPS/Register/register[18][28] ,
         \i_MIPS/Register/register[18][29] ,
         \i_MIPS/Register/register[18][30] ,
         \i_MIPS/Register/register[18][31] , \i_MIPS/Register/register[17][0] ,
         \i_MIPS/Register/register[17][1] , \i_MIPS/Register/register[17][2] ,
         \i_MIPS/Register/register[17][3] , \i_MIPS/Register/register[17][4] ,
         \i_MIPS/Register/register[17][5] , \i_MIPS/Register/register[17][6] ,
         \i_MIPS/Register/register[17][7] , \i_MIPS/Register/register[17][8] ,
         \i_MIPS/Register/register[17][9] , \i_MIPS/Register/register[17][10] ,
         \i_MIPS/Register/register[17][11] ,
         \i_MIPS/Register/register[17][12] ,
         \i_MIPS/Register/register[17][13] ,
         \i_MIPS/Register/register[17][14] ,
         \i_MIPS/Register/register[17][15] ,
         \i_MIPS/Register/register[17][16] ,
         \i_MIPS/Register/register[17][17] ,
         \i_MIPS/Register/register[17][18] ,
         \i_MIPS/Register/register[17][19] ,
         \i_MIPS/Register/register[17][20] ,
         \i_MIPS/Register/register[17][21] ,
         \i_MIPS/Register/register[17][22] ,
         \i_MIPS/Register/register[17][23] ,
         \i_MIPS/Register/register[17][24] ,
         \i_MIPS/Register/register[17][25] ,
         \i_MIPS/Register/register[17][26] ,
         \i_MIPS/Register/register[17][27] ,
         \i_MIPS/Register/register[17][28] ,
         \i_MIPS/Register/register[17][29] ,
         \i_MIPS/Register/register[17][30] ,
         \i_MIPS/Register/register[17][31] , \i_MIPS/Register/register[16][0] ,
         \i_MIPS/Register/register[16][1] , \i_MIPS/Register/register[16][2] ,
         \i_MIPS/Register/register[16][3] , \i_MIPS/Register/register[16][4] ,
         \i_MIPS/Register/register[16][5] , \i_MIPS/Register/register[16][6] ,
         \i_MIPS/Register/register[16][7] , \i_MIPS/Register/register[16][8] ,
         \i_MIPS/Register/register[16][9] , \i_MIPS/Register/register[16][10] ,
         \i_MIPS/Register/register[16][11] ,
         \i_MIPS/Register/register[16][12] ,
         \i_MIPS/Register/register[16][13] ,
         \i_MIPS/Register/register[16][14] ,
         \i_MIPS/Register/register[16][15] ,
         \i_MIPS/Register/register[16][16] ,
         \i_MIPS/Register/register[16][17] ,
         \i_MIPS/Register/register[16][18] ,
         \i_MIPS/Register/register[16][19] ,
         \i_MIPS/Register/register[16][20] ,
         \i_MIPS/Register/register[16][21] ,
         \i_MIPS/Register/register[16][22] ,
         \i_MIPS/Register/register[16][23] ,
         \i_MIPS/Register/register[16][24] ,
         \i_MIPS/Register/register[16][25] ,
         \i_MIPS/Register/register[16][26] ,
         \i_MIPS/Register/register[16][27] ,
         \i_MIPS/Register/register[16][28] ,
         \i_MIPS/Register/register[16][29] ,
         \i_MIPS/Register/register[16][30] ,
         \i_MIPS/Register/register[16][31] , \i_MIPS/Register/register[15][0] ,
         \i_MIPS/Register/register[15][1] , \i_MIPS/Register/register[15][2] ,
         \i_MIPS/Register/register[15][3] , \i_MIPS/Register/register[15][4] ,
         \i_MIPS/Register/register[15][5] , \i_MIPS/Register/register[15][6] ,
         \i_MIPS/Register/register[15][7] , \i_MIPS/Register/register[15][8] ,
         \i_MIPS/Register/register[15][9] , \i_MIPS/Register/register[15][10] ,
         \i_MIPS/Register/register[15][11] ,
         \i_MIPS/Register/register[15][12] ,
         \i_MIPS/Register/register[15][13] ,
         \i_MIPS/Register/register[15][14] ,
         \i_MIPS/Register/register[15][15] ,
         \i_MIPS/Register/register[15][16] ,
         \i_MIPS/Register/register[15][17] ,
         \i_MIPS/Register/register[15][18] ,
         \i_MIPS/Register/register[15][19] ,
         \i_MIPS/Register/register[15][20] ,
         \i_MIPS/Register/register[15][21] ,
         \i_MIPS/Register/register[15][22] ,
         \i_MIPS/Register/register[15][23] ,
         \i_MIPS/Register/register[15][24] ,
         \i_MIPS/Register/register[15][25] ,
         \i_MIPS/Register/register[15][26] ,
         \i_MIPS/Register/register[15][27] ,
         \i_MIPS/Register/register[15][28] ,
         \i_MIPS/Register/register[15][29] ,
         \i_MIPS/Register/register[15][30] ,
         \i_MIPS/Register/register[15][31] , \i_MIPS/Register/register[14][0] ,
         \i_MIPS/Register/register[14][1] , \i_MIPS/Register/register[14][2] ,
         \i_MIPS/Register/register[14][3] , \i_MIPS/Register/register[14][4] ,
         \i_MIPS/Register/register[14][5] , \i_MIPS/Register/register[14][6] ,
         \i_MIPS/Register/register[14][7] , \i_MIPS/Register/register[14][8] ,
         \i_MIPS/Register/register[14][9] , \i_MIPS/Register/register[14][10] ,
         \i_MIPS/Register/register[14][11] ,
         \i_MIPS/Register/register[14][12] ,
         \i_MIPS/Register/register[14][13] ,
         \i_MIPS/Register/register[14][14] ,
         \i_MIPS/Register/register[14][15] ,
         \i_MIPS/Register/register[14][16] ,
         \i_MIPS/Register/register[14][17] ,
         \i_MIPS/Register/register[14][18] ,
         \i_MIPS/Register/register[14][19] ,
         \i_MIPS/Register/register[14][20] ,
         \i_MIPS/Register/register[14][21] ,
         \i_MIPS/Register/register[14][22] ,
         \i_MIPS/Register/register[14][23] ,
         \i_MIPS/Register/register[14][24] ,
         \i_MIPS/Register/register[14][25] ,
         \i_MIPS/Register/register[14][26] ,
         \i_MIPS/Register/register[14][27] ,
         \i_MIPS/Register/register[14][28] ,
         \i_MIPS/Register/register[14][29] ,
         \i_MIPS/Register/register[14][30] ,
         \i_MIPS/Register/register[14][31] , \i_MIPS/Register/register[13][0] ,
         \i_MIPS/Register/register[13][1] , \i_MIPS/Register/register[13][2] ,
         \i_MIPS/Register/register[13][3] , \i_MIPS/Register/register[13][4] ,
         \i_MIPS/Register/register[13][5] , \i_MIPS/Register/register[13][6] ,
         \i_MIPS/Register/register[13][7] , \i_MIPS/Register/register[13][8] ,
         \i_MIPS/Register/register[13][9] , \i_MIPS/Register/register[13][10] ,
         \i_MIPS/Register/register[13][11] ,
         \i_MIPS/Register/register[13][12] ,
         \i_MIPS/Register/register[13][13] ,
         \i_MIPS/Register/register[13][14] ,
         \i_MIPS/Register/register[13][15] ,
         \i_MIPS/Register/register[13][16] ,
         \i_MIPS/Register/register[13][17] ,
         \i_MIPS/Register/register[13][18] ,
         \i_MIPS/Register/register[13][19] ,
         \i_MIPS/Register/register[13][20] ,
         \i_MIPS/Register/register[13][21] ,
         \i_MIPS/Register/register[13][22] ,
         \i_MIPS/Register/register[13][23] ,
         \i_MIPS/Register/register[13][24] ,
         \i_MIPS/Register/register[13][25] ,
         \i_MIPS/Register/register[13][26] ,
         \i_MIPS/Register/register[13][27] ,
         \i_MIPS/Register/register[13][28] ,
         \i_MIPS/Register/register[13][29] ,
         \i_MIPS/Register/register[13][30] ,
         \i_MIPS/Register/register[13][31] , \i_MIPS/Register/register[12][0] ,
         \i_MIPS/Register/register[12][1] , \i_MIPS/Register/register[12][2] ,
         \i_MIPS/Register/register[12][3] , \i_MIPS/Register/register[12][4] ,
         \i_MIPS/Register/register[12][5] , \i_MIPS/Register/register[12][6] ,
         \i_MIPS/Register/register[12][7] , \i_MIPS/Register/register[12][8] ,
         \i_MIPS/Register/register[12][9] , \i_MIPS/Register/register[12][10] ,
         \i_MIPS/Register/register[12][11] ,
         \i_MIPS/Register/register[12][12] ,
         \i_MIPS/Register/register[12][13] ,
         \i_MIPS/Register/register[12][14] ,
         \i_MIPS/Register/register[12][15] ,
         \i_MIPS/Register/register[12][16] ,
         \i_MIPS/Register/register[12][17] ,
         \i_MIPS/Register/register[12][18] ,
         \i_MIPS/Register/register[12][19] ,
         \i_MIPS/Register/register[12][20] ,
         \i_MIPS/Register/register[12][21] ,
         \i_MIPS/Register/register[12][22] ,
         \i_MIPS/Register/register[12][23] ,
         \i_MIPS/Register/register[12][24] ,
         \i_MIPS/Register/register[12][25] ,
         \i_MIPS/Register/register[12][26] ,
         \i_MIPS/Register/register[12][27] ,
         \i_MIPS/Register/register[12][28] ,
         \i_MIPS/Register/register[12][29] ,
         \i_MIPS/Register/register[12][30] ,
         \i_MIPS/Register/register[12][31] , \i_MIPS/Register/register[11][0] ,
         \i_MIPS/Register/register[11][1] , \i_MIPS/Register/register[11][2] ,
         \i_MIPS/Register/register[11][3] , \i_MIPS/Register/register[11][4] ,
         \i_MIPS/Register/register[11][5] , \i_MIPS/Register/register[11][6] ,
         \i_MIPS/Register/register[11][7] , \i_MIPS/Register/register[11][8] ,
         \i_MIPS/Register/register[11][9] , \i_MIPS/Register/register[11][10] ,
         \i_MIPS/Register/register[11][11] ,
         \i_MIPS/Register/register[11][12] ,
         \i_MIPS/Register/register[11][13] ,
         \i_MIPS/Register/register[11][14] ,
         \i_MIPS/Register/register[11][15] ,
         \i_MIPS/Register/register[11][16] ,
         \i_MIPS/Register/register[11][17] ,
         \i_MIPS/Register/register[11][18] ,
         \i_MIPS/Register/register[11][19] ,
         \i_MIPS/Register/register[11][20] ,
         \i_MIPS/Register/register[11][21] ,
         \i_MIPS/Register/register[11][22] ,
         \i_MIPS/Register/register[11][23] ,
         \i_MIPS/Register/register[11][24] ,
         \i_MIPS/Register/register[11][25] ,
         \i_MIPS/Register/register[11][26] ,
         \i_MIPS/Register/register[11][27] ,
         \i_MIPS/Register/register[11][28] ,
         \i_MIPS/Register/register[11][29] ,
         \i_MIPS/Register/register[11][30] ,
         \i_MIPS/Register/register[11][31] , \i_MIPS/Register/register[10][0] ,
         \i_MIPS/Register/register[10][1] , \i_MIPS/Register/register[10][2] ,
         \i_MIPS/Register/register[10][3] , \i_MIPS/Register/register[10][4] ,
         \i_MIPS/Register/register[10][5] , \i_MIPS/Register/register[10][6] ,
         \i_MIPS/Register/register[10][7] , \i_MIPS/Register/register[10][8] ,
         \i_MIPS/Register/register[10][9] , \i_MIPS/Register/register[10][10] ,
         \i_MIPS/Register/register[10][11] ,
         \i_MIPS/Register/register[10][12] ,
         \i_MIPS/Register/register[10][13] ,
         \i_MIPS/Register/register[10][14] ,
         \i_MIPS/Register/register[10][15] ,
         \i_MIPS/Register/register[10][16] ,
         \i_MIPS/Register/register[10][17] ,
         \i_MIPS/Register/register[10][18] ,
         \i_MIPS/Register/register[10][19] ,
         \i_MIPS/Register/register[10][20] ,
         \i_MIPS/Register/register[10][21] ,
         \i_MIPS/Register/register[10][22] ,
         \i_MIPS/Register/register[10][23] ,
         \i_MIPS/Register/register[10][24] ,
         \i_MIPS/Register/register[10][25] ,
         \i_MIPS/Register/register[10][26] ,
         \i_MIPS/Register/register[10][27] ,
         \i_MIPS/Register/register[10][28] ,
         \i_MIPS/Register/register[10][29] ,
         \i_MIPS/Register/register[10][30] ,
         \i_MIPS/Register/register[10][31] , \i_MIPS/Register/register[9][0] ,
         \i_MIPS/Register/register[9][1] , \i_MIPS/Register/register[9][2] ,
         \i_MIPS/Register/register[9][3] , \i_MIPS/Register/register[9][4] ,
         \i_MIPS/Register/register[9][5] , \i_MIPS/Register/register[9][6] ,
         \i_MIPS/Register/register[9][7] , \i_MIPS/Register/register[9][8] ,
         \i_MIPS/Register/register[9][9] , \i_MIPS/Register/register[9][10] ,
         \i_MIPS/Register/register[9][11] , \i_MIPS/Register/register[9][12] ,
         \i_MIPS/Register/register[9][13] , \i_MIPS/Register/register[9][14] ,
         \i_MIPS/Register/register[9][15] , \i_MIPS/Register/register[9][16] ,
         \i_MIPS/Register/register[9][17] , \i_MIPS/Register/register[9][18] ,
         \i_MIPS/Register/register[9][19] , \i_MIPS/Register/register[9][20] ,
         \i_MIPS/Register/register[9][21] , \i_MIPS/Register/register[9][22] ,
         \i_MIPS/Register/register[9][23] , \i_MIPS/Register/register[9][24] ,
         \i_MIPS/Register/register[9][25] , \i_MIPS/Register/register[9][26] ,
         \i_MIPS/Register/register[9][27] , \i_MIPS/Register/register[9][28] ,
         \i_MIPS/Register/register[9][29] , \i_MIPS/Register/register[9][30] ,
         \i_MIPS/Register/register[9][31] , \i_MIPS/Register/register[8][0] ,
         \i_MIPS/Register/register[8][1] , \i_MIPS/Register/register[8][2] ,
         \i_MIPS/Register/register[8][3] , \i_MIPS/Register/register[8][4] ,
         \i_MIPS/Register/register[8][5] , \i_MIPS/Register/register[8][6] ,
         \i_MIPS/Register/register[8][7] , \i_MIPS/Register/register[8][8] ,
         \i_MIPS/Register/register[8][9] , \i_MIPS/Register/register[8][10] ,
         \i_MIPS/Register/register[8][11] , \i_MIPS/Register/register[8][12] ,
         \i_MIPS/Register/register[8][13] , \i_MIPS/Register/register[8][14] ,
         \i_MIPS/Register/register[8][15] , \i_MIPS/Register/register[8][16] ,
         \i_MIPS/Register/register[8][17] , \i_MIPS/Register/register[8][18] ,
         \i_MIPS/Register/register[8][19] , \i_MIPS/Register/register[8][20] ,
         \i_MIPS/Register/register[8][21] , \i_MIPS/Register/register[8][22] ,
         \i_MIPS/Register/register[8][23] , \i_MIPS/Register/register[8][24] ,
         \i_MIPS/Register/register[8][25] , \i_MIPS/Register/register[8][26] ,
         \i_MIPS/Register/register[8][27] , \i_MIPS/Register/register[8][28] ,
         \i_MIPS/Register/register[8][29] , \i_MIPS/Register/register[8][30] ,
         \i_MIPS/Register/register[8][31] , \i_MIPS/Register/register[7][0] ,
         \i_MIPS/Register/register[7][1] , \i_MIPS/Register/register[7][2] ,
         \i_MIPS/Register/register[7][3] , \i_MIPS/Register/register[7][4] ,
         \i_MIPS/Register/register[7][5] , \i_MIPS/Register/register[7][6] ,
         \i_MIPS/Register/register[7][7] , \i_MIPS/Register/register[7][8] ,
         \i_MIPS/Register/register[7][9] , \i_MIPS/Register/register[7][10] ,
         \i_MIPS/Register/register[7][11] , \i_MIPS/Register/register[7][12] ,
         \i_MIPS/Register/register[7][13] , \i_MIPS/Register/register[7][14] ,
         \i_MIPS/Register/register[7][15] , \i_MIPS/Register/register[7][16] ,
         \i_MIPS/Register/register[7][17] , \i_MIPS/Register/register[7][18] ,
         \i_MIPS/Register/register[7][19] , \i_MIPS/Register/register[7][20] ,
         \i_MIPS/Register/register[7][21] , \i_MIPS/Register/register[7][22] ,
         \i_MIPS/Register/register[7][23] , \i_MIPS/Register/register[7][24] ,
         \i_MIPS/Register/register[7][25] , \i_MIPS/Register/register[7][26] ,
         \i_MIPS/Register/register[7][27] , \i_MIPS/Register/register[7][28] ,
         \i_MIPS/Register/register[7][29] , \i_MIPS/Register/register[7][30] ,
         \i_MIPS/Register/register[7][31] , \i_MIPS/Register/register[6][0] ,
         \i_MIPS/Register/register[6][1] , \i_MIPS/Register/register[6][2] ,
         \i_MIPS/Register/register[6][3] , \i_MIPS/Register/register[6][4] ,
         \i_MIPS/Register/register[6][5] , \i_MIPS/Register/register[6][6] ,
         \i_MIPS/Register/register[6][7] , \i_MIPS/Register/register[6][8] ,
         \i_MIPS/Register/register[6][9] , \i_MIPS/Register/register[6][10] ,
         \i_MIPS/Register/register[6][11] , \i_MIPS/Register/register[6][12] ,
         \i_MIPS/Register/register[6][13] , \i_MIPS/Register/register[6][14] ,
         \i_MIPS/Register/register[6][15] , \i_MIPS/Register/register[6][16] ,
         \i_MIPS/Register/register[6][17] , \i_MIPS/Register/register[6][18] ,
         \i_MIPS/Register/register[6][19] , \i_MIPS/Register/register[6][20] ,
         \i_MIPS/Register/register[6][21] , \i_MIPS/Register/register[6][22] ,
         \i_MIPS/Register/register[6][23] , \i_MIPS/Register/register[6][24] ,
         \i_MIPS/Register/register[6][25] , \i_MIPS/Register/register[6][26] ,
         \i_MIPS/Register/register[6][27] , \i_MIPS/Register/register[6][28] ,
         \i_MIPS/Register/register[6][29] , \i_MIPS/Register/register[6][30] ,
         \i_MIPS/Register/register[6][31] , \i_MIPS/Register/register[5][0] ,
         \i_MIPS/Register/register[5][1] , \i_MIPS/Register/register[5][2] ,
         \i_MIPS/Register/register[5][3] , \i_MIPS/Register/register[5][4] ,
         \i_MIPS/Register/register[5][5] , \i_MIPS/Register/register[5][6] ,
         \i_MIPS/Register/register[5][7] , \i_MIPS/Register/register[5][8] ,
         \i_MIPS/Register/register[5][9] , \i_MIPS/Register/register[5][10] ,
         \i_MIPS/Register/register[5][11] , \i_MIPS/Register/register[5][12] ,
         \i_MIPS/Register/register[5][13] , \i_MIPS/Register/register[5][14] ,
         \i_MIPS/Register/register[5][15] , \i_MIPS/Register/register[5][16] ,
         \i_MIPS/Register/register[5][17] , \i_MIPS/Register/register[5][18] ,
         \i_MIPS/Register/register[5][19] , \i_MIPS/Register/register[5][20] ,
         \i_MIPS/Register/register[5][21] , \i_MIPS/Register/register[5][22] ,
         \i_MIPS/Register/register[5][23] , \i_MIPS/Register/register[5][24] ,
         \i_MIPS/Register/register[5][25] , \i_MIPS/Register/register[5][26] ,
         \i_MIPS/Register/register[5][27] , \i_MIPS/Register/register[5][28] ,
         \i_MIPS/Register/register[5][29] , \i_MIPS/Register/register[5][30] ,
         \i_MIPS/Register/register[5][31] , \i_MIPS/Register/register[4][0] ,
         \i_MIPS/Register/register[4][1] , \i_MIPS/Register/register[4][2] ,
         \i_MIPS/Register/register[4][3] , \i_MIPS/Register/register[4][4] ,
         \i_MIPS/Register/register[4][5] , \i_MIPS/Register/register[4][6] ,
         \i_MIPS/Register/register[4][7] , \i_MIPS/Register/register[4][8] ,
         \i_MIPS/Register/register[4][9] , \i_MIPS/Register/register[4][10] ,
         \i_MIPS/Register/register[4][11] , \i_MIPS/Register/register[4][12] ,
         \i_MIPS/Register/register[4][13] , \i_MIPS/Register/register[4][14] ,
         \i_MIPS/Register/register[4][15] , \i_MIPS/Register/register[4][16] ,
         \i_MIPS/Register/register[4][17] , \i_MIPS/Register/register[4][18] ,
         \i_MIPS/Register/register[4][19] , \i_MIPS/Register/register[4][20] ,
         \i_MIPS/Register/register[4][21] , \i_MIPS/Register/register[4][22] ,
         \i_MIPS/Register/register[4][23] , \i_MIPS/Register/register[4][24] ,
         \i_MIPS/Register/register[4][25] , \i_MIPS/Register/register[4][26] ,
         \i_MIPS/Register/register[4][27] , \i_MIPS/Register/register[4][28] ,
         \i_MIPS/Register/register[4][29] , \i_MIPS/Register/register[4][30] ,
         \i_MIPS/Register/register[4][31] , \i_MIPS/Register/register[3][0] ,
         \i_MIPS/Register/register[3][1] , \i_MIPS/Register/register[3][2] ,
         \i_MIPS/Register/register[3][3] , \i_MIPS/Register/register[3][4] ,
         \i_MIPS/Register/register[3][5] , \i_MIPS/Register/register[3][6] ,
         \i_MIPS/Register/register[3][7] , \i_MIPS/Register/register[3][8] ,
         \i_MIPS/Register/register[3][9] , \i_MIPS/Register/register[3][10] ,
         \i_MIPS/Register/register[3][11] , \i_MIPS/Register/register[3][12] ,
         \i_MIPS/Register/register[3][13] , \i_MIPS/Register/register[3][14] ,
         \i_MIPS/Register/register[3][15] , \i_MIPS/Register/register[3][16] ,
         \i_MIPS/Register/register[3][17] , \i_MIPS/Register/register[3][18] ,
         \i_MIPS/Register/register[3][19] , \i_MIPS/Register/register[3][20] ,
         \i_MIPS/Register/register[3][21] , \i_MIPS/Register/register[3][22] ,
         \i_MIPS/Register/register[3][23] , \i_MIPS/Register/register[3][24] ,
         \i_MIPS/Register/register[3][25] , \i_MIPS/Register/register[3][26] ,
         \i_MIPS/Register/register[3][27] , \i_MIPS/Register/register[3][28] ,
         \i_MIPS/Register/register[3][29] , \i_MIPS/Register/register[3][30] ,
         \i_MIPS/Register/register[3][31] , \i_MIPS/Register/register[2][0] ,
         \i_MIPS/Register/register[2][1] , \i_MIPS/Register/register[2][2] ,
         \i_MIPS/Register/register[2][3] , \i_MIPS/Register/register[2][4] ,
         \i_MIPS/Register/register[2][5] , \i_MIPS/Register/register[2][6] ,
         \i_MIPS/Register/register[2][7] , \i_MIPS/Register/register[2][8] ,
         \i_MIPS/Register/register[2][9] , \i_MIPS/Register/register[2][10] ,
         \i_MIPS/Register/register[2][11] , \i_MIPS/Register/register[2][12] ,
         \i_MIPS/Register/register[2][13] , \i_MIPS/Register/register[2][14] ,
         \i_MIPS/Register/register[2][15] , \i_MIPS/Register/register[2][16] ,
         \i_MIPS/Register/register[2][17] , \i_MIPS/Register/register[2][18] ,
         \i_MIPS/Register/register[2][19] , \i_MIPS/Register/register[2][20] ,
         \i_MIPS/Register/register[2][21] , \i_MIPS/Register/register[2][22] ,
         \i_MIPS/Register/register[2][23] , \i_MIPS/Register/register[2][24] ,
         \i_MIPS/Register/register[2][25] , \i_MIPS/Register/register[2][26] ,
         \i_MIPS/Register/register[2][27] , \i_MIPS/Register/register[2][28] ,
         \i_MIPS/Register/register[2][29] , \i_MIPS/Register/register[2][30] ,
         \i_MIPS/Register/register[2][31] , \i_MIPS/Register/register[1][0] ,
         \i_MIPS/Register/register[1][1] , \i_MIPS/Register/register[1][2] ,
         \i_MIPS/Register/register[1][3] , \i_MIPS/Register/register[1][4] ,
         \i_MIPS/Register/register[1][5] , \i_MIPS/Register/register[1][6] ,
         \i_MIPS/Register/register[1][7] , \i_MIPS/Register/register[1][8] ,
         \i_MIPS/Register/register[1][9] , \i_MIPS/Register/register[1][10] ,
         \i_MIPS/Register/register[1][11] , \i_MIPS/Register/register[1][12] ,
         \i_MIPS/Register/register[1][13] , \i_MIPS/Register/register[1][14] ,
         \i_MIPS/Register/register[1][15] , \i_MIPS/Register/register[1][16] ,
         \i_MIPS/Register/register[1][17] , \i_MIPS/Register/register[1][18] ,
         \i_MIPS/Register/register[1][19] , \i_MIPS/Register/register[1][20] ,
         \i_MIPS/Register/register[1][21] , \i_MIPS/Register/register[1][22] ,
         \i_MIPS/Register/register[1][23] , \i_MIPS/Register/register[1][24] ,
         \i_MIPS/Register/register[1][25] , \i_MIPS/Register/register[1][26] ,
         \i_MIPS/Register/register[1][27] , \i_MIPS/Register/register[1][28] ,
         \i_MIPS/Register/register[1][29] , \i_MIPS/Register/register[1][30] ,
         \i_MIPS/Register/register[1][31] , \i_MIPS/Register/register[0][0] ,
         \i_MIPS/Register/register[0][1] , \i_MIPS/Register/register[0][2] ,
         \i_MIPS/Register/register[0][3] , \i_MIPS/Register/register[0][4] ,
         \i_MIPS/Register/register[0][5] , \i_MIPS/Register/register[0][6] ,
         \i_MIPS/Register/register[0][7] , \i_MIPS/Register/register[0][8] ,
         \i_MIPS/Register/register[0][9] , \i_MIPS/Register/register[0][10] ,
         \i_MIPS/Register/register[0][11] , \i_MIPS/Register/register[0][12] ,
         \i_MIPS/Register/register[0][13] , \i_MIPS/Register/register[0][14] ,
         \i_MIPS/Register/register[0][15] , \i_MIPS/Register/register[0][16] ,
         \i_MIPS/Register/register[0][17] , \i_MIPS/Register/register[0][18] ,
         \i_MIPS/Register/register[0][19] , \i_MIPS/Register/register[0][20] ,
         \i_MIPS/Register/register[0][21] , \i_MIPS/Register/register[0][22] ,
         \i_MIPS/Register/register[0][23] , \i_MIPS/Register/register[0][24] ,
         \i_MIPS/Register/register[0][25] , \i_MIPS/Register/register[0][26] ,
         \i_MIPS/Register/register[0][27] , \i_MIPS/Register/register[0][28] ,
         \i_MIPS/Register/register[0][29] , \i_MIPS/Register/register[0][30] ,
         \i_MIPS/Register/register[0][31] , \i_MIPS/Control_ID/n15 ,
         \i_MIPS/Control_ID/n12 , \i_MIPS/Control_ID/n10 ,
         \i_MIPS/Hazard_detection/n13 , \i_MIPS/Hazard_detection/n12 ,
         \i_MIPS/Hazard_detection/n11 , \i_MIPS/Hazard_detection/n10 ,
         \i_MIPS/Hazard_detection/n9 , \i_MIPS/Hazard_detection/n8 ,
         \i_MIPS/Hazard_detection/n7 , \i_MIPS/Hazard_detection/n4 ,
         \i_MIPS/forward_unit/n32 , \i_MIPS/forward_unit/n25 ,
         \i_MIPS/forward_unit/n15 , \i_MIPS/forward_unit/n10 ,
         \i_MIPS/ALU_Control/n20 , \i_MIPS/ALU_Control/n18 ,
         \i_MIPS/ALU_Control/n15 , \i_MIPS/ALU_Control/n11 ,
         \i_MIPS/ALU_Control/n10 , \i_MIPS/ALU/N303 , \I_cache/cache[7][0] ,
         \I_cache/cache[7][1] , \I_cache/cache[7][2] , \I_cache/cache[7][3] ,
         \I_cache/cache[7][4] , \I_cache/cache[7][5] , \I_cache/cache[7][6] ,
         \I_cache/cache[7][7] , \I_cache/cache[7][8] , \I_cache/cache[7][9] ,
         \I_cache/cache[7][10] , \I_cache/cache[7][11] ,
         \I_cache/cache[7][12] , \I_cache/cache[7][13] ,
         \I_cache/cache[7][14] , \I_cache/cache[7][15] ,
         \I_cache/cache[7][16] , \I_cache/cache[7][17] ,
         \I_cache/cache[7][18] , \I_cache/cache[7][19] ,
         \I_cache/cache[7][20] , \I_cache/cache[7][21] ,
         \I_cache/cache[7][22] , \I_cache/cache[7][23] ,
         \I_cache/cache[7][24] , \I_cache/cache[7][25] ,
         \I_cache/cache[7][26] , \I_cache/cache[7][27] ,
         \I_cache/cache[7][28] , \I_cache/cache[7][29] ,
         \I_cache/cache[7][30] , \I_cache/cache[7][31] ,
         \I_cache/cache[7][32] , \I_cache/cache[7][33] ,
         \I_cache/cache[7][34] , \I_cache/cache[7][35] ,
         \I_cache/cache[7][36] , \I_cache/cache[7][37] ,
         \I_cache/cache[7][38] , \I_cache/cache[7][39] ,
         \I_cache/cache[7][40] , \I_cache/cache[7][41] ,
         \I_cache/cache[7][42] , \I_cache/cache[7][43] ,
         \I_cache/cache[7][44] , \I_cache/cache[7][45] ,
         \I_cache/cache[7][46] , \I_cache/cache[7][47] ,
         \I_cache/cache[7][48] , \I_cache/cache[7][49] ,
         \I_cache/cache[7][50] , \I_cache/cache[7][51] ,
         \I_cache/cache[7][52] , \I_cache/cache[7][53] ,
         \I_cache/cache[7][54] , \I_cache/cache[7][55] ,
         \I_cache/cache[7][56] , \I_cache/cache[7][57] ,
         \I_cache/cache[7][58] , \I_cache/cache[7][59] ,
         \I_cache/cache[7][60] , \I_cache/cache[7][61] ,
         \I_cache/cache[7][62] , \I_cache/cache[7][63] ,
         \I_cache/cache[7][64] , \I_cache/cache[7][65] ,
         \I_cache/cache[7][66] , \I_cache/cache[7][67] ,
         \I_cache/cache[7][68] , \I_cache/cache[7][69] ,
         \I_cache/cache[7][70] , \I_cache/cache[7][71] ,
         \I_cache/cache[7][72] , \I_cache/cache[7][73] ,
         \I_cache/cache[7][74] , \I_cache/cache[7][75] ,
         \I_cache/cache[7][76] , \I_cache/cache[7][77] ,
         \I_cache/cache[7][78] , \I_cache/cache[7][79] ,
         \I_cache/cache[7][80] , \I_cache/cache[7][81] ,
         \I_cache/cache[7][82] , \I_cache/cache[7][83] ,
         \I_cache/cache[7][84] , \I_cache/cache[7][85] ,
         \I_cache/cache[7][86] , \I_cache/cache[7][87] ,
         \I_cache/cache[7][88] , \I_cache/cache[7][89] ,
         \I_cache/cache[7][90] , \I_cache/cache[7][91] ,
         \I_cache/cache[7][92] , \I_cache/cache[7][93] ,
         \I_cache/cache[7][94] , \I_cache/cache[7][95] ,
         \I_cache/cache[7][96] , \I_cache/cache[7][97] ,
         \I_cache/cache[7][98] , \I_cache/cache[7][99] ,
         \I_cache/cache[7][100] , \I_cache/cache[7][101] ,
         \I_cache/cache[7][102] , \I_cache/cache[7][103] ,
         \I_cache/cache[7][104] , \I_cache/cache[7][105] ,
         \I_cache/cache[7][106] , \I_cache/cache[7][107] ,
         \I_cache/cache[7][108] , \I_cache/cache[7][109] ,
         \I_cache/cache[7][110] , \I_cache/cache[7][111] ,
         \I_cache/cache[7][112] , \I_cache/cache[7][113] ,
         \I_cache/cache[7][114] , \I_cache/cache[7][115] ,
         \I_cache/cache[7][116] , \I_cache/cache[7][117] ,
         \I_cache/cache[7][118] , \I_cache/cache[7][119] ,
         \I_cache/cache[7][120] , \I_cache/cache[7][121] ,
         \I_cache/cache[7][122] , \I_cache/cache[7][123] ,
         \I_cache/cache[7][124] , \I_cache/cache[7][125] ,
         \I_cache/cache[7][126] , \I_cache/cache[7][127] ,
         \I_cache/cache[7][128] , \I_cache/cache[7][129] ,
         \I_cache/cache[7][130] , \I_cache/cache[7][131] ,
         \I_cache/cache[7][132] , \I_cache/cache[7][133] ,
         \I_cache/cache[7][134] , \I_cache/cache[7][135] ,
         \I_cache/cache[7][136] , \I_cache/cache[7][137] ,
         \I_cache/cache[7][138] , \I_cache/cache[7][139] ,
         \I_cache/cache[7][140] , \I_cache/cache[7][141] ,
         \I_cache/cache[7][142] , \I_cache/cache[7][143] ,
         \I_cache/cache[7][144] , \I_cache/cache[7][145] ,
         \I_cache/cache[7][146] , \I_cache/cache[7][147] ,
         \I_cache/cache[7][148] , \I_cache/cache[7][149] ,
         \I_cache/cache[7][150] , \I_cache/cache[7][151] ,
         \I_cache/cache[7][152] , \I_cache/cache[7][153] ,
         \I_cache/cache[7][154] , \I_cache/cache[6][0] , \I_cache/cache[6][1] ,
         \I_cache/cache[6][2] , \I_cache/cache[6][3] , \I_cache/cache[6][4] ,
         \I_cache/cache[6][5] , \I_cache/cache[6][6] , \I_cache/cache[6][7] ,
         \I_cache/cache[6][8] , \I_cache/cache[6][9] , \I_cache/cache[6][10] ,
         \I_cache/cache[6][11] , \I_cache/cache[6][12] ,
         \I_cache/cache[6][13] , \I_cache/cache[6][14] ,
         \I_cache/cache[6][15] , \I_cache/cache[6][16] ,
         \I_cache/cache[6][17] , \I_cache/cache[6][18] ,
         \I_cache/cache[6][19] , \I_cache/cache[6][20] ,
         \I_cache/cache[6][21] , \I_cache/cache[6][22] ,
         \I_cache/cache[6][23] , \I_cache/cache[6][24] ,
         \I_cache/cache[6][25] , \I_cache/cache[6][26] ,
         \I_cache/cache[6][27] , \I_cache/cache[6][28] ,
         \I_cache/cache[6][29] , \I_cache/cache[6][30] ,
         \I_cache/cache[6][31] , \I_cache/cache[6][32] ,
         \I_cache/cache[6][33] , \I_cache/cache[6][34] ,
         \I_cache/cache[6][35] , \I_cache/cache[6][36] ,
         \I_cache/cache[6][37] , \I_cache/cache[6][38] ,
         \I_cache/cache[6][39] , \I_cache/cache[6][40] ,
         \I_cache/cache[6][41] , \I_cache/cache[6][42] ,
         \I_cache/cache[6][43] , \I_cache/cache[6][44] ,
         \I_cache/cache[6][45] , \I_cache/cache[6][46] ,
         \I_cache/cache[6][47] , \I_cache/cache[6][48] ,
         \I_cache/cache[6][49] , \I_cache/cache[6][50] ,
         \I_cache/cache[6][51] , \I_cache/cache[6][52] ,
         \I_cache/cache[6][53] , \I_cache/cache[6][54] ,
         \I_cache/cache[6][55] , \I_cache/cache[6][56] ,
         \I_cache/cache[6][57] , \I_cache/cache[6][58] ,
         \I_cache/cache[6][59] , \I_cache/cache[6][60] ,
         \I_cache/cache[6][61] , \I_cache/cache[6][62] ,
         \I_cache/cache[6][63] , \I_cache/cache[6][64] ,
         \I_cache/cache[6][65] , \I_cache/cache[6][66] ,
         \I_cache/cache[6][67] , \I_cache/cache[6][68] ,
         \I_cache/cache[6][69] , \I_cache/cache[6][70] ,
         \I_cache/cache[6][71] , \I_cache/cache[6][72] ,
         \I_cache/cache[6][73] , \I_cache/cache[6][74] ,
         \I_cache/cache[6][75] , \I_cache/cache[6][76] ,
         \I_cache/cache[6][77] , \I_cache/cache[6][78] ,
         \I_cache/cache[6][79] , \I_cache/cache[6][80] ,
         \I_cache/cache[6][81] , \I_cache/cache[6][82] ,
         \I_cache/cache[6][83] , \I_cache/cache[6][84] ,
         \I_cache/cache[6][85] , \I_cache/cache[6][86] ,
         \I_cache/cache[6][87] , \I_cache/cache[6][88] ,
         \I_cache/cache[6][89] , \I_cache/cache[6][90] ,
         \I_cache/cache[6][91] , \I_cache/cache[6][92] ,
         \I_cache/cache[6][93] , \I_cache/cache[6][94] ,
         \I_cache/cache[6][95] , \I_cache/cache[6][96] ,
         \I_cache/cache[6][97] , \I_cache/cache[6][98] ,
         \I_cache/cache[6][99] , \I_cache/cache[6][100] ,
         \I_cache/cache[6][101] , \I_cache/cache[6][102] ,
         \I_cache/cache[6][103] , \I_cache/cache[6][104] ,
         \I_cache/cache[6][105] , \I_cache/cache[6][106] ,
         \I_cache/cache[6][107] , \I_cache/cache[6][108] ,
         \I_cache/cache[6][109] , \I_cache/cache[6][110] ,
         \I_cache/cache[6][111] , \I_cache/cache[6][112] ,
         \I_cache/cache[6][113] , \I_cache/cache[6][114] ,
         \I_cache/cache[6][115] , \I_cache/cache[6][116] ,
         \I_cache/cache[6][117] , \I_cache/cache[6][118] ,
         \I_cache/cache[6][119] , \I_cache/cache[6][120] ,
         \I_cache/cache[6][121] , \I_cache/cache[6][122] ,
         \I_cache/cache[6][123] , \I_cache/cache[6][124] ,
         \I_cache/cache[6][125] , \I_cache/cache[6][126] ,
         \I_cache/cache[6][127] , \I_cache/cache[6][128] ,
         \I_cache/cache[6][129] , \I_cache/cache[6][130] ,
         \I_cache/cache[6][131] , \I_cache/cache[6][132] ,
         \I_cache/cache[6][133] , \I_cache/cache[6][134] ,
         \I_cache/cache[6][135] , \I_cache/cache[6][136] ,
         \I_cache/cache[6][137] , \I_cache/cache[6][138] ,
         \I_cache/cache[6][139] , \I_cache/cache[6][140] ,
         \I_cache/cache[6][141] , \I_cache/cache[6][142] ,
         \I_cache/cache[6][143] , \I_cache/cache[6][144] ,
         \I_cache/cache[6][145] , \I_cache/cache[6][146] ,
         \I_cache/cache[6][147] , \I_cache/cache[6][148] ,
         \I_cache/cache[6][149] , \I_cache/cache[6][150] ,
         \I_cache/cache[6][151] , \I_cache/cache[6][152] ,
         \I_cache/cache[6][153] , \I_cache/cache[6][154] ,
         \I_cache/cache[5][0] , \I_cache/cache[5][1] , \I_cache/cache[5][2] ,
         \I_cache/cache[5][3] , \I_cache/cache[5][4] , \I_cache/cache[5][5] ,
         \I_cache/cache[5][6] , \I_cache/cache[5][7] , \I_cache/cache[5][8] ,
         \I_cache/cache[5][9] , \I_cache/cache[5][10] , \I_cache/cache[5][11] ,
         \I_cache/cache[5][12] , \I_cache/cache[5][13] ,
         \I_cache/cache[5][14] , \I_cache/cache[5][15] ,
         \I_cache/cache[5][16] , \I_cache/cache[5][17] ,
         \I_cache/cache[5][18] , \I_cache/cache[5][19] ,
         \I_cache/cache[5][20] , \I_cache/cache[5][21] ,
         \I_cache/cache[5][22] , \I_cache/cache[5][23] ,
         \I_cache/cache[5][24] , \I_cache/cache[5][25] ,
         \I_cache/cache[5][26] , \I_cache/cache[5][27] ,
         \I_cache/cache[5][28] , \I_cache/cache[5][29] ,
         \I_cache/cache[5][30] , \I_cache/cache[5][31] ,
         \I_cache/cache[5][32] , \I_cache/cache[5][33] ,
         \I_cache/cache[5][34] , \I_cache/cache[5][35] ,
         \I_cache/cache[5][36] , \I_cache/cache[5][37] ,
         \I_cache/cache[5][38] , \I_cache/cache[5][39] ,
         \I_cache/cache[5][40] , \I_cache/cache[5][41] ,
         \I_cache/cache[5][42] , \I_cache/cache[5][43] ,
         \I_cache/cache[5][44] , \I_cache/cache[5][45] ,
         \I_cache/cache[5][46] , \I_cache/cache[5][47] ,
         \I_cache/cache[5][48] , \I_cache/cache[5][49] ,
         \I_cache/cache[5][50] , \I_cache/cache[5][51] ,
         \I_cache/cache[5][52] , \I_cache/cache[5][53] ,
         \I_cache/cache[5][54] , \I_cache/cache[5][55] ,
         \I_cache/cache[5][56] , \I_cache/cache[5][57] ,
         \I_cache/cache[5][58] , \I_cache/cache[5][59] ,
         \I_cache/cache[5][60] , \I_cache/cache[5][61] ,
         \I_cache/cache[5][62] , \I_cache/cache[5][63] ,
         \I_cache/cache[5][64] , \I_cache/cache[5][65] ,
         \I_cache/cache[5][66] , \I_cache/cache[5][67] ,
         \I_cache/cache[5][68] , \I_cache/cache[5][69] ,
         \I_cache/cache[5][70] , \I_cache/cache[5][71] ,
         \I_cache/cache[5][72] , \I_cache/cache[5][73] ,
         \I_cache/cache[5][74] , \I_cache/cache[5][75] ,
         \I_cache/cache[5][76] , \I_cache/cache[5][77] ,
         \I_cache/cache[5][78] , \I_cache/cache[5][79] ,
         \I_cache/cache[5][80] , \I_cache/cache[5][81] ,
         \I_cache/cache[5][82] , \I_cache/cache[5][83] ,
         \I_cache/cache[5][84] , \I_cache/cache[5][85] ,
         \I_cache/cache[5][86] , \I_cache/cache[5][87] ,
         \I_cache/cache[5][88] , \I_cache/cache[5][89] ,
         \I_cache/cache[5][90] , \I_cache/cache[5][91] ,
         \I_cache/cache[5][92] , \I_cache/cache[5][93] ,
         \I_cache/cache[5][94] , \I_cache/cache[5][95] ,
         \I_cache/cache[5][96] , \I_cache/cache[5][97] ,
         \I_cache/cache[5][98] , \I_cache/cache[5][99] ,
         \I_cache/cache[5][100] , \I_cache/cache[5][101] ,
         \I_cache/cache[5][102] , \I_cache/cache[5][103] ,
         \I_cache/cache[5][104] , \I_cache/cache[5][105] ,
         \I_cache/cache[5][106] , \I_cache/cache[5][107] ,
         \I_cache/cache[5][108] , \I_cache/cache[5][109] ,
         \I_cache/cache[5][110] , \I_cache/cache[5][111] ,
         \I_cache/cache[5][112] , \I_cache/cache[5][113] ,
         \I_cache/cache[5][114] , \I_cache/cache[5][115] ,
         \I_cache/cache[5][116] , \I_cache/cache[5][117] ,
         \I_cache/cache[5][118] , \I_cache/cache[5][119] ,
         \I_cache/cache[5][120] , \I_cache/cache[5][121] ,
         \I_cache/cache[5][122] , \I_cache/cache[5][123] ,
         \I_cache/cache[5][124] , \I_cache/cache[5][125] ,
         \I_cache/cache[5][126] , \I_cache/cache[5][127] ,
         \I_cache/cache[5][128] , \I_cache/cache[5][129] ,
         \I_cache/cache[5][130] , \I_cache/cache[5][131] ,
         \I_cache/cache[5][132] , \I_cache/cache[5][133] ,
         \I_cache/cache[5][134] , \I_cache/cache[5][135] ,
         \I_cache/cache[5][136] , \I_cache/cache[5][137] ,
         \I_cache/cache[5][138] , \I_cache/cache[5][139] ,
         \I_cache/cache[5][140] , \I_cache/cache[5][141] ,
         \I_cache/cache[5][142] , \I_cache/cache[5][143] ,
         \I_cache/cache[5][144] , \I_cache/cache[5][145] ,
         \I_cache/cache[5][146] , \I_cache/cache[5][147] ,
         \I_cache/cache[5][148] , \I_cache/cache[5][149] ,
         \I_cache/cache[5][150] , \I_cache/cache[5][151] ,
         \I_cache/cache[5][152] , \I_cache/cache[5][153] ,
         \I_cache/cache[5][154] , \I_cache/cache[4][0] , \I_cache/cache[4][1] ,
         \I_cache/cache[4][2] , \I_cache/cache[4][3] , \I_cache/cache[4][4] ,
         \I_cache/cache[4][5] , \I_cache/cache[4][6] , \I_cache/cache[4][7] ,
         \I_cache/cache[4][8] , \I_cache/cache[4][9] , \I_cache/cache[4][10] ,
         \I_cache/cache[4][11] , \I_cache/cache[4][12] ,
         \I_cache/cache[4][13] , \I_cache/cache[4][14] ,
         \I_cache/cache[4][15] , \I_cache/cache[4][16] ,
         \I_cache/cache[4][17] , \I_cache/cache[4][18] ,
         \I_cache/cache[4][19] , \I_cache/cache[4][20] ,
         \I_cache/cache[4][21] , \I_cache/cache[4][22] ,
         \I_cache/cache[4][23] , \I_cache/cache[4][24] ,
         \I_cache/cache[4][25] , \I_cache/cache[4][26] ,
         \I_cache/cache[4][27] , \I_cache/cache[4][28] ,
         \I_cache/cache[4][29] , \I_cache/cache[4][30] ,
         \I_cache/cache[4][31] , \I_cache/cache[4][32] ,
         \I_cache/cache[4][33] , \I_cache/cache[4][34] ,
         \I_cache/cache[4][35] , \I_cache/cache[4][36] ,
         \I_cache/cache[4][37] , \I_cache/cache[4][38] ,
         \I_cache/cache[4][39] , \I_cache/cache[4][40] ,
         \I_cache/cache[4][41] , \I_cache/cache[4][42] ,
         \I_cache/cache[4][43] , \I_cache/cache[4][44] ,
         \I_cache/cache[4][45] , \I_cache/cache[4][46] ,
         \I_cache/cache[4][47] , \I_cache/cache[4][48] ,
         \I_cache/cache[4][49] , \I_cache/cache[4][50] ,
         \I_cache/cache[4][51] , \I_cache/cache[4][52] ,
         \I_cache/cache[4][53] , \I_cache/cache[4][54] ,
         \I_cache/cache[4][55] , \I_cache/cache[4][56] ,
         \I_cache/cache[4][57] , \I_cache/cache[4][58] ,
         \I_cache/cache[4][59] , \I_cache/cache[4][60] ,
         \I_cache/cache[4][61] , \I_cache/cache[4][62] ,
         \I_cache/cache[4][63] , \I_cache/cache[4][64] ,
         \I_cache/cache[4][65] , \I_cache/cache[4][66] ,
         \I_cache/cache[4][67] , \I_cache/cache[4][68] ,
         \I_cache/cache[4][69] , \I_cache/cache[4][70] ,
         \I_cache/cache[4][71] , \I_cache/cache[4][72] ,
         \I_cache/cache[4][73] , \I_cache/cache[4][74] ,
         \I_cache/cache[4][75] , \I_cache/cache[4][76] ,
         \I_cache/cache[4][77] , \I_cache/cache[4][78] ,
         \I_cache/cache[4][79] , \I_cache/cache[4][80] ,
         \I_cache/cache[4][81] , \I_cache/cache[4][82] ,
         \I_cache/cache[4][83] , \I_cache/cache[4][84] ,
         \I_cache/cache[4][85] , \I_cache/cache[4][86] ,
         \I_cache/cache[4][87] , \I_cache/cache[4][88] ,
         \I_cache/cache[4][89] , \I_cache/cache[4][90] ,
         \I_cache/cache[4][91] , \I_cache/cache[4][92] ,
         \I_cache/cache[4][93] , \I_cache/cache[4][94] ,
         \I_cache/cache[4][95] , \I_cache/cache[4][96] ,
         \I_cache/cache[4][97] , \I_cache/cache[4][98] ,
         \I_cache/cache[4][99] , \I_cache/cache[4][100] ,
         \I_cache/cache[4][101] , \I_cache/cache[4][102] ,
         \I_cache/cache[4][103] , \I_cache/cache[4][104] ,
         \I_cache/cache[4][105] , \I_cache/cache[4][106] ,
         \I_cache/cache[4][107] , \I_cache/cache[4][108] ,
         \I_cache/cache[4][109] , \I_cache/cache[4][110] ,
         \I_cache/cache[4][111] , \I_cache/cache[4][112] ,
         \I_cache/cache[4][113] , \I_cache/cache[4][114] ,
         \I_cache/cache[4][115] , \I_cache/cache[4][116] ,
         \I_cache/cache[4][117] , \I_cache/cache[4][118] ,
         \I_cache/cache[4][119] , \I_cache/cache[4][120] ,
         \I_cache/cache[4][121] , \I_cache/cache[4][122] ,
         \I_cache/cache[4][123] , \I_cache/cache[4][124] ,
         \I_cache/cache[4][125] , \I_cache/cache[4][126] ,
         \I_cache/cache[4][127] , \I_cache/cache[4][128] ,
         \I_cache/cache[4][129] , \I_cache/cache[4][130] ,
         \I_cache/cache[4][131] , \I_cache/cache[4][132] ,
         \I_cache/cache[4][133] , \I_cache/cache[4][134] ,
         \I_cache/cache[4][135] , \I_cache/cache[4][136] ,
         \I_cache/cache[4][137] , \I_cache/cache[4][138] ,
         \I_cache/cache[4][139] , \I_cache/cache[4][140] ,
         \I_cache/cache[4][141] , \I_cache/cache[4][142] ,
         \I_cache/cache[4][143] , \I_cache/cache[4][144] ,
         \I_cache/cache[4][145] , \I_cache/cache[4][146] ,
         \I_cache/cache[4][147] , \I_cache/cache[4][148] ,
         \I_cache/cache[4][149] , \I_cache/cache[4][150] ,
         \I_cache/cache[4][151] , \I_cache/cache[4][152] ,
         \I_cache/cache[4][153] , \I_cache/cache[4][154] ,
         \I_cache/cache[3][0] , \I_cache/cache[3][1] , \I_cache/cache[3][2] ,
         \I_cache/cache[3][3] , \I_cache/cache[3][4] , \I_cache/cache[3][5] ,
         \I_cache/cache[3][6] , \I_cache/cache[3][7] , \I_cache/cache[3][8] ,
         \I_cache/cache[3][9] , \I_cache/cache[3][10] , \I_cache/cache[3][11] ,
         \I_cache/cache[3][12] , \I_cache/cache[3][13] ,
         \I_cache/cache[3][14] , \I_cache/cache[3][15] ,
         \I_cache/cache[3][16] , \I_cache/cache[3][17] ,
         \I_cache/cache[3][18] , \I_cache/cache[3][19] ,
         \I_cache/cache[3][20] , \I_cache/cache[3][21] ,
         \I_cache/cache[3][22] , \I_cache/cache[3][23] ,
         \I_cache/cache[3][24] , \I_cache/cache[3][25] ,
         \I_cache/cache[3][26] , \I_cache/cache[3][27] ,
         \I_cache/cache[3][28] , \I_cache/cache[3][29] ,
         \I_cache/cache[3][30] , \I_cache/cache[3][31] ,
         \I_cache/cache[3][32] , \I_cache/cache[3][33] ,
         \I_cache/cache[3][34] , \I_cache/cache[3][35] ,
         \I_cache/cache[3][36] , \I_cache/cache[3][37] ,
         \I_cache/cache[3][38] , \I_cache/cache[3][39] ,
         \I_cache/cache[3][40] , \I_cache/cache[3][41] ,
         \I_cache/cache[3][42] , \I_cache/cache[3][43] ,
         \I_cache/cache[3][44] , \I_cache/cache[3][45] ,
         \I_cache/cache[3][46] , \I_cache/cache[3][47] ,
         \I_cache/cache[3][48] , \I_cache/cache[3][49] ,
         \I_cache/cache[3][50] , \I_cache/cache[3][51] ,
         \I_cache/cache[3][52] , \I_cache/cache[3][53] ,
         \I_cache/cache[3][54] , \I_cache/cache[3][55] ,
         \I_cache/cache[3][56] , \I_cache/cache[3][57] ,
         \I_cache/cache[3][58] , \I_cache/cache[3][59] ,
         \I_cache/cache[3][60] , \I_cache/cache[3][61] ,
         \I_cache/cache[3][62] , \I_cache/cache[3][63] ,
         \I_cache/cache[3][64] , \I_cache/cache[3][65] ,
         \I_cache/cache[3][66] , \I_cache/cache[3][67] ,
         \I_cache/cache[3][68] , \I_cache/cache[3][69] ,
         \I_cache/cache[3][70] , \I_cache/cache[3][71] ,
         \I_cache/cache[3][72] , \I_cache/cache[3][73] ,
         \I_cache/cache[3][74] , \I_cache/cache[3][75] ,
         \I_cache/cache[3][76] , \I_cache/cache[3][77] ,
         \I_cache/cache[3][78] , \I_cache/cache[3][79] ,
         \I_cache/cache[3][80] , \I_cache/cache[3][81] ,
         \I_cache/cache[3][82] , \I_cache/cache[3][83] ,
         \I_cache/cache[3][84] , \I_cache/cache[3][85] ,
         \I_cache/cache[3][86] , \I_cache/cache[3][87] ,
         \I_cache/cache[3][88] , \I_cache/cache[3][89] ,
         \I_cache/cache[3][90] , \I_cache/cache[3][91] ,
         \I_cache/cache[3][92] , \I_cache/cache[3][93] ,
         \I_cache/cache[3][94] , \I_cache/cache[3][95] ,
         \I_cache/cache[3][96] , \I_cache/cache[3][97] ,
         \I_cache/cache[3][98] , \I_cache/cache[3][99] ,
         \I_cache/cache[3][100] , \I_cache/cache[3][101] ,
         \I_cache/cache[3][102] , \I_cache/cache[3][103] ,
         \I_cache/cache[3][104] , \I_cache/cache[3][105] ,
         \I_cache/cache[3][106] , \I_cache/cache[3][107] ,
         \I_cache/cache[3][108] , \I_cache/cache[3][109] ,
         \I_cache/cache[3][110] , \I_cache/cache[3][111] ,
         \I_cache/cache[3][112] , \I_cache/cache[3][113] ,
         \I_cache/cache[3][114] , \I_cache/cache[3][115] ,
         \I_cache/cache[3][116] , \I_cache/cache[3][117] ,
         \I_cache/cache[3][118] , \I_cache/cache[3][119] ,
         \I_cache/cache[3][120] , \I_cache/cache[3][121] ,
         \I_cache/cache[3][122] , \I_cache/cache[3][123] ,
         \I_cache/cache[3][124] , \I_cache/cache[3][125] ,
         \I_cache/cache[3][126] , \I_cache/cache[3][127] ,
         \I_cache/cache[3][128] , \I_cache/cache[3][129] ,
         \I_cache/cache[3][130] , \I_cache/cache[3][131] ,
         \I_cache/cache[3][132] , \I_cache/cache[3][133] ,
         \I_cache/cache[3][134] , \I_cache/cache[3][135] ,
         \I_cache/cache[3][136] , \I_cache/cache[3][137] ,
         \I_cache/cache[3][138] , \I_cache/cache[3][139] ,
         \I_cache/cache[3][140] , \I_cache/cache[3][141] ,
         \I_cache/cache[3][142] , \I_cache/cache[3][143] ,
         \I_cache/cache[3][144] , \I_cache/cache[3][145] ,
         \I_cache/cache[3][146] , \I_cache/cache[3][147] ,
         \I_cache/cache[3][148] , \I_cache/cache[3][149] ,
         \I_cache/cache[3][150] , \I_cache/cache[3][151] ,
         \I_cache/cache[3][152] , \I_cache/cache[3][153] ,
         \I_cache/cache[3][154] , \I_cache/cache[2][0] , \I_cache/cache[2][1] ,
         \I_cache/cache[2][2] , \I_cache/cache[2][3] , \I_cache/cache[2][4] ,
         \I_cache/cache[2][5] , \I_cache/cache[2][6] , \I_cache/cache[2][7] ,
         \I_cache/cache[2][8] , \I_cache/cache[2][9] , \I_cache/cache[2][10] ,
         \I_cache/cache[2][11] , \I_cache/cache[2][12] ,
         \I_cache/cache[2][13] , \I_cache/cache[2][14] ,
         \I_cache/cache[2][15] , \I_cache/cache[2][16] ,
         \I_cache/cache[2][17] , \I_cache/cache[2][18] ,
         \I_cache/cache[2][19] , \I_cache/cache[2][20] ,
         \I_cache/cache[2][21] , \I_cache/cache[2][22] ,
         \I_cache/cache[2][23] , \I_cache/cache[2][24] ,
         \I_cache/cache[2][25] , \I_cache/cache[2][26] ,
         \I_cache/cache[2][27] , \I_cache/cache[2][28] ,
         \I_cache/cache[2][29] , \I_cache/cache[2][30] ,
         \I_cache/cache[2][31] , \I_cache/cache[2][32] ,
         \I_cache/cache[2][33] , \I_cache/cache[2][34] ,
         \I_cache/cache[2][35] , \I_cache/cache[2][36] ,
         \I_cache/cache[2][37] , \I_cache/cache[2][38] ,
         \I_cache/cache[2][39] , \I_cache/cache[2][40] ,
         \I_cache/cache[2][41] , \I_cache/cache[2][42] ,
         \I_cache/cache[2][43] , \I_cache/cache[2][44] ,
         \I_cache/cache[2][45] , \I_cache/cache[2][46] ,
         \I_cache/cache[2][47] , \I_cache/cache[2][48] ,
         \I_cache/cache[2][49] , \I_cache/cache[2][50] ,
         \I_cache/cache[2][51] , \I_cache/cache[2][52] ,
         \I_cache/cache[2][53] , \I_cache/cache[2][54] ,
         \I_cache/cache[2][55] , \I_cache/cache[2][56] ,
         \I_cache/cache[2][57] , \I_cache/cache[2][58] ,
         \I_cache/cache[2][59] , \I_cache/cache[2][60] ,
         \I_cache/cache[2][61] , \I_cache/cache[2][62] ,
         \I_cache/cache[2][63] , \I_cache/cache[2][64] ,
         \I_cache/cache[2][65] , \I_cache/cache[2][66] ,
         \I_cache/cache[2][67] , \I_cache/cache[2][68] ,
         \I_cache/cache[2][69] , \I_cache/cache[2][70] ,
         \I_cache/cache[2][71] , \I_cache/cache[2][72] ,
         \I_cache/cache[2][73] , \I_cache/cache[2][74] ,
         \I_cache/cache[2][75] , \I_cache/cache[2][76] ,
         \I_cache/cache[2][77] , \I_cache/cache[2][78] ,
         \I_cache/cache[2][79] , \I_cache/cache[2][80] ,
         \I_cache/cache[2][81] , \I_cache/cache[2][82] ,
         \I_cache/cache[2][83] , \I_cache/cache[2][84] ,
         \I_cache/cache[2][85] , \I_cache/cache[2][86] ,
         \I_cache/cache[2][87] , \I_cache/cache[2][88] ,
         \I_cache/cache[2][89] , \I_cache/cache[2][90] ,
         \I_cache/cache[2][91] , \I_cache/cache[2][92] ,
         \I_cache/cache[2][93] , \I_cache/cache[2][94] ,
         \I_cache/cache[2][95] , \I_cache/cache[2][96] ,
         \I_cache/cache[2][97] , \I_cache/cache[2][98] ,
         \I_cache/cache[2][99] , \I_cache/cache[2][100] ,
         \I_cache/cache[2][101] , \I_cache/cache[2][102] ,
         \I_cache/cache[2][103] , \I_cache/cache[2][104] ,
         \I_cache/cache[2][105] , \I_cache/cache[2][106] ,
         \I_cache/cache[2][107] , \I_cache/cache[2][108] ,
         \I_cache/cache[2][109] , \I_cache/cache[2][110] ,
         \I_cache/cache[2][111] , \I_cache/cache[2][112] ,
         \I_cache/cache[2][113] , \I_cache/cache[2][114] ,
         \I_cache/cache[2][115] , \I_cache/cache[2][116] ,
         \I_cache/cache[2][117] , \I_cache/cache[2][118] ,
         \I_cache/cache[2][119] , \I_cache/cache[2][120] ,
         \I_cache/cache[2][121] , \I_cache/cache[2][122] ,
         \I_cache/cache[2][123] , \I_cache/cache[2][124] ,
         \I_cache/cache[2][125] , \I_cache/cache[2][126] ,
         \I_cache/cache[2][127] , \I_cache/cache[2][128] ,
         \I_cache/cache[2][129] , \I_cache/cache[2][130] ,
         \I_cache/cache[2][131] , \I_cache/cache[2][132] ,
         \I_cache/cache[2][133] , \I_cache/cache[2][134] ,
         \I_cache/cache[2][135] , \I_cache/cache[2][136] ,
         \I_cache/cache[2][137] , \I_cache/cache[2][138] ,
         \I_cache/cache[2][139] , \I_cache/cache[2][140] ,
         \I_cache/cache[2][141] , \I_cache/cache[2][142] ,
         \I_cache/cache[2][143] , \I_cache/cache[2][144] ,
         \I_cache/cache[2][145] , \I_cache/cache[2][146] ,
         \I_cache/cache[2][147] , \I_cache/cache[2][148] ,
         \I_cache/cache[2][149] , \I_cache/cache[2][150] ,
         \I_cache/cache[2][151] , \I_cache/cache[2][152] ,
         \I_cache/cache[2][153] , \I_cache/cache[2][154] ,
         \I_cache/cache[1][0] , \I_cache/cache[1][1] , \I_cache/cache[1][2] ,
         \I_cache/cache[1][3] , \I_cache/cache[1][4] , \I_cache/cache[1][5] ,
         \I_cache/cache[1][6] , \I_cache/cache[1][7] , \I_cache/cache[1][8] ,
         \I_cache/cache[1][9] , \I_cache/cache[1][10] , \I_cache/cache[1][11] ,
         \I_cache/cache[1][12] , \I_cache/cache[1][13] ,
         \I_cache/cache[1][14] , \I_cache/cache[1][15] ,
         \I_cache/cache[1][16] , \I_cache/cache[1][17] ,
         \I_cache/cache[1][18] , \I_cache/cache[1][19] ,
         \I_cache/cache[1][20] , \I_cache/cache[1][21] ,
         \I_cache/cache[1][22] , \I_cache/cache[1][23] ,
         \I_cache/cache[1][24] , \I_cache/cache[1][25] ,
         \I_cache/cache[1][26] , \I_cache/cache[1][27] ,
         \I_cache/cache[1][28] , \I_cache/cache[1][29] ,
         \I_cache/cache[1][30] , \I_cache/cache[1][31] ,
         \I_cache/cache[1][32] , \I_cache/cache[1][33] ,
         \I_cache/cache[1][34] , \I_cache/cache[1][35] ,
         \I_cache/cache[1][36] , \I_cache/cache[1][37] ,
         \I_cache/cache[1][38] , \I_cache/cache[1][39] ,
         \I_cache/cache[1][40] , \I_cache/cache[1][41] ,
         \I_cache/cache[1][42] , \I_cache/cache[1][43] ,
         \I_cache/cache[1][44] , \I_cache/cache[1][45] ,
         \I_cache/cache[1][46] , \I_cache/cache[1][47] ,
         \I_cache/cache[1][48] , \I_cache/cache[1][49] ,
         \I_cache/cache[1][50] , \I_cache/cache[1][51] ,
         \I_cache/cache[1][52] , \I_cache/cache[1][53] ,
         \I_cache/cache[1][54] , \I_cache/cache[1][55] ,
         \I_cache/cache[1][56] , \I_cache/cache[1][57] ,
         \I_cache/cache[1][58] , \I_cache/cache[1][59] ,
         \I_cache/cache[1][60] , \I_cache/cache[1][61] ,
         \I_cache/cache[1][62] , \I_cache/cache[1][63] ,
         \I_cache/cache[1][64] , \I_cache/cache[1][65] ,
         \I_cache/cache[1][66] , \I_cache/cache[1][67] ,
         \I_cache/cache[1][68] , \I_cache/cache[1][69] ,
         \I_cache/cache[1][70] , \I_cache/cache[1][71] ,
         \I_cache/cache[1][72] , \I_cache/cache[1][73] ,
         \I_cache/cache[1][74] , \I_cache/cache[1][75] ,
         \I_cache/cache[1][76] , \I_cache/cache[1][77] ,
         \I_cache/cache[1][78] , \I_cache/cache[1][79] ,
         \I_cache/cache[1][80] , \I_cache/cache[1][81] ,
         \I_cache/cache[1][82] , \I_cache/cache[1][83] ,
         \I_cache/cache[1][84] , \I_cache/cache[1][85] ,
         \I_cache/cache[1][86] , \I_cache/cache[1][87] ,
         \I_cache/cache[1][88] , \I_cache/cache[1][89] ,
         \I_cache/cache[1][90] , \I_cache/cache[1][91] ,
         \I_cache/cache[1][92] , \I_cache/cache[1][93] ,
         \I_cache/cache[1][94] , \I_cache/cache[1][95] ,
         \I_cache/cache[1][96] , \I_cache/cache[1][97] ,
         \I_cache/cache[1][98] , \I_cache/cache[1][99] ,
         \I_cache/cache[1][100] , \I_cache/cache[1][101] ,
         \I_cache/cache[1][102] , \I_cache/cache[1][103] ,
         \I_cache/cache[1][104] , \I_cache/cache[1][105] ,
         \I_cache/cache[1][106] , \I_cache/cache[1][107] ,
         \I_cache/cache[1][108] , \I_cache/cache[1][109] ,
         \I_cache/cache[1][110] , \I_cache/cache[1][111] ,
         \I_cache/cache[1][112] , \I_cache/cache[1][113] ,
         \I_cache/cache[1][114] , \I_cache/cache[1][115] ,
         \I_cache/cache[1][116] , \I_cache/cache[1][117] ,
         \I_cache/cache[1][118] , \I_cache/cache[1][119] ,
         \I_cache/cache[1][120] , \I_cache/cache[1][121] ,
         \I_cache/cache[1][122] , \I_cache/cache[1][123] ,
         \I_cache/cache[1][124] , \I_cache/cache[1][125] ,
         \I_cache/cache[1][126] , \I_cache/cache[1][127] ,
         \I_cache/cache[1][128] , \I_cache/cache[1][129] ,
         \I_cache/cache[1][130] , \I_cache/cache[1][131] ,
         \I_cache/cache[1][132] , \I_cache/cache[1][133] ,
         \I_cache/cache[1][134] , \I_cache/cache[1][135] ,
         \I_cache/cache[1][136] , \I_cache/cache[1][137] ,
         \I_cache/cache[1][138] , \I_cache/cache[1][139] ,
         \I_cache/cache[1][140] , \I_cache/cache[1][141] ,
         \I_cache/cache[1][142] , \I_cache/cache[1][143] ,
         \I_cache/cache[1][144] , \I_cache/cache[1][145] ,
         \I_cache/cache[1][146] , \I_cache/cache[1][147] ,
         \I_cache/cache[1][148] , \I_cache/cache[1][149] ,
         \I_cache/cache[1][150] , \I_cache/cache[1][151] ,
         \I_cache/cache[1][152] , \I_cache/cache[1][153] ,
         \I_cache/cache[1][154] , \I_cache/cache[0][0] , \I_cache/cache[0][1] ,
         \I_cache/cache[0][2] , \I_cache/cache[0][3] , \I_cache/cache[0][4] ,
         \I_cache/cache[0][5] , \I_cache/cache[0][6] , \I_cache/cache[0][7] ,
         \I_cache/cache[0][8] , \I_cache/cache[0][9] , \I_cache/cache[0][10] ,
         \I_cache/cache[0][11] , \I_cache/cache[0][12] ,
         \I_cache/cache[0][13] , \I_cache/cache[0][14] ,
         \I_cache/cache[0][15] , \I_cache/cache[0][16] ,
         \I_cache/cache[0][17] , \I_cache/cache[0][18] ,
         \I_cache/cache[0][19] , \I_cache/cache[0][20] ,
         \I_cache/cache[0][21] , \I_cache/cache[0][22] ,
         \I_cache/cache[0][23] , \I_cache/cache[0][24] ,
         \I_cache/cache[0][25] , \I_cache/cache[0][26] ,
         \I_cache/cache[0][27] , \I_cache/cache[0][28] ,
         \I_cache/cache[0][29] , \I_cache/cache[0][30] ,
         \I_cache/cache[0][31] , \I_cache/cache[0][32] ,
         \I_cache/cache[0][33] , \I_cache/cache[0][34] ,
         \I_cache/cache[0][35] , \I_cache/cache[0][36] ,
         \I_cache/cache[0][37] , \I_cache/cache[0][38] ,
         \I_cache/cache[0][39] , \I_cache/cache[0][40] ,
         \I_cache/cache[0][41] , \I_cache/cache[0][42] ,
         \I_cache/cache[0][43] , \I_cache/cache[0][44] ,
         \I_cache/cache[0][45] , \I_cache/cache[0][46] ,
         \I_cache/cache[0][47] , \I_cache/cache[0][48] ,
         \I_cache/cache[0][49] , \I_cache/cache[0][50] ,
         \I_cache/cache[0][51] , \I_cache/cache[0][52] ,
         \I_cache/cache[0][53] , \I_cache/cache[0][54] ,
         \I_cache/cache[0][55] , \I_cache/cache[0][56] ,
         \I_cache/cache[0][57] , \I_cache/cache[0][58] ,
         \I_cache/cache[0][59] , \I_cache/cache[0][60] ,
         \I_cache/cache[0][61] , \I_cache/cache[0][62] ,
         \I_cache/cache[0][63] , \I_cache/cache[0][64] ,
         \I_cache/cache[0][65] , \I_cache/cache[0][66] ,
         \I_cache/cache[0][67] , \I_cache/cache[0][68] ,
         \I_cache/cache[0][69] , \I_cache/cache[0][70] ,
         \I_cache/cache[0][71] , \I_cache/cache[0][72] ,
         \I_cache/cache[0][73] , \I_cache/cache[0][74] ,
         \I_cache/cache[0][75] , \I_cache/cache[0][76] ,
         \I_cache/cache[0][77] , \I_cache/cache[0][78] ,
         \I_cache/cache[0][79] , \I_cache/cache[0][80] ,
         \I_cache/cache[0][81] , \I_cache/cache[0][82] ,
         \I_cache/cache[0][83] , \I_cache/cache[0][84] ,
         \I_cache/cache[0][85] , \I_cache/cache[0][86] ,
         \I_cache/cache[0][87] , \I_cache/cache[0][88] ,
         \I_cache/cache[0][89] , \I_cache/cache[0][90] ,
         \I_cache/cache[0][91] , \I_cache/cache[0][92] ,
         \I_cache/cache[0][93] , \I_cache/cache[0][94] ,
         \I_cache/cache[0][95] , \I_cache/cache[0][96] ,
         \I_cache/cache[0][97] , \I_cache/cache[0][98] ,
         \I_cache/cache[0][99] , \I_cache/cache[0][100] ,
         \I_cache/cache[0][101] , \I_cache/cache[0][102] ,
         \I_cache/cache[0][103] , \I_cache/cache[0][104] ,
         \I_cache/cache[0][105] , \I_cache/cache[0][106] ,
         \I_cache/cache[0][107] , \I_cache/cache[0][108] ,
         \I_cache/cache[0][109] , \I_cache/cache[0][110] ,
         \I_cache/cache[0][111] , \I_cache/cache[0][112] ,
         \I_cache/cache[0][113] , \I_cache/cache[0][114] ,
         \I_cache/cache[0][115] , \I_cache/cache[0][116] ,
         \I_cache/cache[0][117] , \I_cache/cache[0][118] ,
         \I_cache/cache[0][119] , \I_cache/cache[0][120] ,
         \I_cache/cache[0][121] , \I_cache/cache[0][122] ,
         \I_cache/cache[0][123] , \I_cache/cache[0][124] ,
         \I_cache/cache[0][125] , \I_cache/cache[0][126] ,
         \I_cache/cache[0][127] , \I_cache/cache[0][128] ,
         \I_cache/cache[0][129] , \I_cache/cache[0][130] ,
         \I_cache/cache[0][131] , \I_cache/cache[0][132] ,
         \I_cache/cache[0][133] , \I_cache/cache[0][134] ,
         \I_cache/cache[0][135] , \I_cache/cache[0][136] ,
         \I_cache/cache[0][137] , \I_cache/cache[0][138] ,
         \I_cache/cache[0][139] , \I_cache/cache[0][140] ,
         \I_cache/cache[0][141] , \I_cache/cache[0][142] ,
         \I_cache/cache[0][143] , \I_cache/cache[0][144] ,
         \I_cache/cache[0][145] , \I_cache/cache[0][146] ,
         \I_cache/cache[0][147] , \I_cache/cache[0][148] ,
         \I_cache/cache[0][149] , \I_cache/cache[0][150] ,
         \I_cache/cache[0][151] , \I_cache/cache[0][152] ,
         \I_cache/cache[0][153] , \I_cache/cache[0][154] , n2, n3, n4, n5, n6,
         n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n139, n140, n141, n142, n143, n144, n145, n146, n147,
         n148, n149, n150, n151, n152, n153, n154, n155, n156, n157, n158,
         n159, n160, n161, n162, n163, n164, n165, n166, n167, n168, n169,
         n170, n171, n172, n173, n174, n175, n176, n177, n178, n179, n180,
         n181, n182, n183, n184, n185, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n305, n306, n307, n308, n309, n310, n311, n312,
         n313, n314, n315, n316, n317, n318, n319, n320, n321, n322, n323,
         n324, n325, n326, n327, n328, n329, n330, n331, n332, n333, n334,
         n335, n336, n337, n338, n339, n340, n341, n342, n343, n344, n345,
         n346, n347, n348, n349, n350, n351, n352, n353, n354, n355, n356,
         n357, n358, n359, n360, n361, n362, n363, n364, n365, n366, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694, n695, n696, n697,
         n698, n699, n700, n701, n702, n703, n704, n705, n706, n707, n708,
         n709, n710, n711, n712, n713, n714, n715, n716, n717, n718, n719,
         n720, n721, n722, n723, n724, n725, n726, n727, n728, n729, n730,
         n731, n732, n733, n734, n735, n736, n737, n738, n739, n740, n741,
         n742, n743, n744, n745, n746, n747, n748, n749, n750, n751, n752,
         n753, n754, n755, n756, n757, n758, n759, n760, n761, n762, n763,
         n764, n765, n766, n767, n768, n769, n770, n771, n772, n773, n774,
         n775, n776, n777, n778, n779, n780, n781, n782, n783, n784, n785,
         n786, n787, n788, n789, n790, n791, n792, n793, n794, n795, n796,
         n797, n798, n799, n800, n801, n802, n803, n804, n805, n806, n807,
         n808, n809, n810, n811, n812, n813, n814, n815, n816, n817, n818,
         n819, n820, n821, n822, n823, n824, n825, n826, n827, n828, n829,
         n830, n831, n832, n833, n834, n835, n836, n837, n838, n839, n840,
         n841, n842, n843, n844, n845, n846, n847, n848, n849, n850, n851,
         n852, n853, n854, n855, n856, n857, n858, n859, n860, n861, n862,
         n863, n864, n865, n866, n867, n868, n869, n870, n871, n872, n873,
         n874, n875, n876, n877, n878, n879, n880, n881, n882, n883, n884,
         n885, n886, n887, n888, n889, n890, n891, n892, n893, n894, n895,
         n896, n897, n898, n899, n900, n901, n902, n903, n904, n905, n906,
         n907, n908, n909, n910, n911, n912, n913, n914, n915, n916, n917,
         n918, n919, n920, n921, n922, n923, n924, n925, n926, n927, n928,
         n929, n930, n931, n932, n933, n934, n935, n936, n937, n938, n939,
         n940, n941, n942, n943, n944, n945, n946, n947, n948, n949, n950,
         n951, n952, n953, n954, n955, n956, n957, n958, n959, n960, n961,
         n962, n963, n964, n965, n966, n967, n968, n969, n970, n971, n972,
         n973, n974, n975, n976, n977, n978, n979, n980, n981, n982, n983,
         n984, n985, n986, n987, n988, n989, n990, n991, n992, n993, n994,
         n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004,
         n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014,
         n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024,
         n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034,
         n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044,
         n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054,
         n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064,
         n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074,
         n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084,
         n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094,
         n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104,
         n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114,
         n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123, n1124,
         n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134,
         n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144,
         n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154,
         n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164,
         n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174,
         n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184,
         n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1194,
         n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203, n1204,
         n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213, n1214,
         n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223, n1224,
         n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233, n1234,
         n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243, n1244,
         n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253, n1254,
         n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263, n1264,
         n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273, n1274,
         n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283, n1284,
         n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293, n1294,
         n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303, n1304,
         n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313, n1314,
         n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323, n1324,
         n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333, n1334,
         n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343, n1344,
         n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353, n1354,
         n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363, n1364,
         n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373, n1374,
         n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383, n1384,
         n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393, n1394,
         n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403, n1404,
         n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413, n1414,
         n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423, n1424,
         n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433, n1434,
         n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443, n1444,
         n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453, n1454,
         n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463, n1464,
         n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474,
         n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484,
         n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494,
         n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504,
         n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514,
         n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524,
         n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534,
         n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544,
         n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554,
         n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564,
         n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574,
         n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583, n1584,
         n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593, n1594,
         n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603, n1604,
         n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613, n1614,
         n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623, n1624,
         n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633, n1634,
         n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643, n1644,
         n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653, n1654,
         n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663, n1664,
         n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673, n1674,
         n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683, n1684,
         n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693, n1694,
         n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703, n1704,
         n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713, n1714,
         n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723, n1724,
         n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733, n1734,
         n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743, n1744,
         n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753, n1754,
         n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763, n1764,
         n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773, n1774,
         n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783, n1784,
         n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793, n1794,
         n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803, n1804,
         n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813, n1814,
         n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823, n1824,
         n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833, n1834,
         n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843, n1844,
         n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853, n1854,
         n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863, n1864,
         n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873, n1874,
         n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883, n1884,
         n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893, n1894,
         n1915, n1917, n1919, n1921, n1923, n1925, n1927, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2223, n2224,
         n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233, n2234,
         n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243, n2244,
         n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253, n2254,
         n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263, n2264,
         n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273, n2274,
         n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283, n2284,
         n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293, n2294,
         n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303, n2304,
         n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313, n2314,
         n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323, n2324,
         n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333, n2334,
         n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343, n2344,
         n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353, n2354,
         n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363, n2364,
         n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373, n2374,
         n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383, n2384,
         n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393, n2394,
         n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403, n2404,
         n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413, n2414,
         n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423, n2424,
         n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433, n2434,
         n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2448, n2449, n2450,
         n2451, n2452, n2453, n2464, n2465, n2466, n2467, n2468, n2469, n2485,
         n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2508,
         n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518,
         n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575,
         n2576, n2577, n2578, n2579, n2596, n2597, n2598, n2599, n2600, n2601,
         n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2623, n2624,
         n2625, n2626, n2627, n2628, n2630, n2631, n2632, n2633, n2650, n2651,
         n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661,
         n2701, n2703, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2724,
         n2725, n2726, n2727, n2728, n2730, n2731, n2732, n2733, n2734, n2735,
         n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745,
         n2746, n2747, n2748, n2750, n2751, n2752, n2753, n2754, n2755, n2756,
         n2757, n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766,
         n2767, n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776,
         n2777, n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786,
         n2787, n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796,
         n2797, n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806,
         n2807, n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816,
         n2817, n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826,
         n2827, n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836,
         n2837, n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846,
         n2847, n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856,
         n2857, n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866,
         n2867, n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876,
         n2877, n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886,
         n2887, n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896,
         n2897, n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906,
         n2907, n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916,
         n2917, n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926,
         n2927, n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936,
         n2937, n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946,
         n2947, n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956,
         n2957, n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966,
         n2967, n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976,
         n2977, n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986,
         n2987, n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996,
         n2997, n3000, n3001, n3002, n3010, n3015, n3016, n3017, n3019, n3020,
         n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030,
         n3031, n3032, n3033, n3034, n3036, n3037, n3038, n3039, n3040, n3041,
         n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
         n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
         n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
         n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
         n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
         n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
         n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
         n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
         n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
         n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
         n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
         n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
         n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
         n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
         n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
         n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
         n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
         n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
         n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
         n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
         n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
         n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
         n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
         n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
         n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953,
         n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963,
         n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973,
         n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983,
         n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993,
         n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
         n4004, n4005, n4006, n4007, n4010, n4011, n4012, n4013, n4014, n4015,
         n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023, n4024, n4025,
         n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033, n4034, n4035,
         n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043, n4044, n4045,
         n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053, n4054, n4055,
         n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063, n4064, n4065,
         n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075,
         n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085,
         n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095,
         n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105,
         n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115,
         n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125,
         n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135,
         n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145,
         n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155,
         n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165,
         n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175,
         n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185,
         n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195,
         n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205,
         n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215,
         n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225,
         n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235,
         n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245,
         n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253, n4254, n4255,
         n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263, n4264, n4265,
         n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273, n4274, n4275,
         n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283, n4284, n4285,
         n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293, n4294, n4295,
         n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305,
         n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315,
         n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325,
         n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335,
         n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345,
         n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355,
         n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365,
         n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375,
         n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385,
         n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395,
         n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405,
         n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415,
         n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425,
         n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435,
         n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445,
         n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455,
         n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465,
         n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475,
         n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485,
         n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495,
         n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505,
         n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515,
         n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525,
         n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535,
         n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4545,
         n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553, n4554, n4555,
         n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563, n4564, n4565,
         n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573, n4574, n4575,
         n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583, n4584, n4585,
         n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593, n4594, n4595,
         n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603, n4604, n4605,
         n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614, n4615,
         n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625,
         n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635,
         n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645,
         n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655,
         n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665,
         n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
         n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
         n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
         n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
         n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
         n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
         n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
         n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
         n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
         n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
         n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
         n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
         n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,
         n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,
         n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
         n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
         n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
         n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,
         n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125,
         n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,
         n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145,
         n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155,
         n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165,
         n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175,
         n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185,
         n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195,
         n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205,
         n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215,
         n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225,
         n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235,
         n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245,
         n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255,
         n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265,
         n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275,
         n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285,
         n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295,
         n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305,
         n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315,
         n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325,
         n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335,
         n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345,
         n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355,
         n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365,
         n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
         n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,
         n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395,
         n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405,
         n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415,
         n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425,
         n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435,
         n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445,
         n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455,
         n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465,
         n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475,
         n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485,
         n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495,
         n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505,
         n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515,
         n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525,
         n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535,
         n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545,
         n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553, n5554, n5555,
         n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563, n5564, n5565,
         n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573, n5574, n5575,
         n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583, n5584, n5585,
         n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593, n5594, n5595,
         n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603, n5604, n5605,
         n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613, n5614, n5615,
         n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623, n5624, n5625,
         n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633, n5634, n5635,
         n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643, n5644, n5645,
         n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653, n5654, n5655,
         n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663, n5664, n5665,
         n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673, n5674, n5675,
         n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683, n5684, n5685,
         n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693, n5694, n5695,
         n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703, n5704, n5705,
         n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713, n5714, n5715,
         n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723, n5724, n5725,
         n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733, n5734, n5735,
         n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743, n5744, n5745,
         n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753, n5754, n5755,
         n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763, n5764, n5765,
         n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773, n5774, n5775,
         n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783, n5784, n5785,
         n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793, n5794, n5795,
         n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803, n5804, n5805,
         n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813, n5814, n5815,
         n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823, n5824, n5825,
         n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833, n5834, n5835,
         n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843, n5844, n5845,
         n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853, n5854, n5855,
         n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863, n5864, n5865,
         n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873, n5874, n5875,
         n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883, n5884, n5885,
         n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893, n5894, n5895,
         n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903, n5904, n5905,
         n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913, n5914, n5915,
         n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923, n5924, n5925,
         n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933, n5934, n5935,
         n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943, n5944, n5945,
         n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953, n5954, n5955,
         n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963, n5964, n5965,
         n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973, n5974, n5975,
         n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983, n5984, n5985,
         n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993, n5994, n5995,
         n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003, n6004, n6005,
         n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013, n6014, n6015,
         n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023, n6024, n6025,
         n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033, n6034, n6035,
         n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043, n6044, n6045,
         n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053, n6054, n6055,
         n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063, n6064, n6065,
         n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073, n6074, n6075,
         n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083, n6084, n6085,
         n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093, n6094, n6095,
         n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103, n6104, n6105,
         n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113, n6114, n6115,
         n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123, n6124, n6125,
         n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133, n6134, n6135,
         n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143, n6144, n6145,
         n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153, n6154, n6155,
         n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163, n6164, n6165,
         n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173, n6174, n6175,
         n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183, n6184, n6185,
         n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193, n6194, n6195,
         n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203, n6204, n6205,
         n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213, n6214, n6215,
         n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223, n6224, n6225,
         n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233, n6234, n6235,
         n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243, n6244, n6245,
         n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253, n6254, n6255,
         n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263, n6264, n6265,
         n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273, n6274, n6275,
         n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283, n6284, n6285,
         n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293, n6294, n6295,
         n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303, n6304, n6305,
         n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313, n6314, n6315,
         n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323, n6324, n6325,
         n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333, n6334, n6335,
         n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343, n6344, n6345,
         n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353, n6354, n6355,
         n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363, n6364, n6365,
         n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373, n6374, n6375,
         n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383, n6384, n6385,
         n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393, n6394, n6395,
         n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403, n6404, n6405,
         n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413, n6414, n6415,
         n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423, n6424, n6425,
         n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433, n6434, n6435,
         n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443, n6444, n6445,
         n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453, n6454, n6455,
         n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463, n6464, n6465,
         n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473, n6474, n6475,
         n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483, n6484, n6485,
         n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493, n6494, n6495,
         n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503, n6504, n6505,
         n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513, n6514, n6515,
         n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523, n6524, n6525,
         n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533, n6534, n6535,
         n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543, n6544, n6545,
         n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553, n6554, n6555,
         n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563, n6564, n6565,
         n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573, n6574, n6575,
         n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583, n6584, n6585,
         n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593, n6594, n6595,
         n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603, n6604, n6605,
         n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613, n6614, n6615,
         n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623, n6624, n6625,
         n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633, n6634, n6635,
         n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643, n6644, n6645,
         n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653, n6654, n6655,
         n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663, n6664, n6665,
         n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673, n6674, n6675,
         n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683, n6684, n6685,
         n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693, n6694, n6695,
         n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703, n6704, n6705,
         n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713, n6714, n6715,
         n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723, n6724, n6725,
         n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733, n6734, n6735,
         n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743, n6744, n6745,
         n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753, n6754, n6755,
         n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763, n6764, n6765,
         n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773, n6774, n6775,
         n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783, n6784, n6785,
         n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793, n6794, n6795,
         n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803, n6804, n6805,
         n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813, n6814, n6815,
         n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823, n6824, n6825,
         n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833, n6834, n6835,
         n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843, n6844, n6845,
         n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853, n6854, n6855,
         n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863, n6864, n6865,
         n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873, n6874, n6875,
         n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883, n6884, n6885,
         n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893, n6894, n6895,
         n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903, n6904, n6905,
         n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913, n6914, n6915,
         n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923, n6924, n6925,
         n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933, n6934, n6935,
         n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943, n6944, n6945,
         n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953, n6954, n6955,
         n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963, n6964, n6965,
         n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973, n6974, n6975,
         n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983, n6984, n6985,
         n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993, n6994, n6995,
         n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003, n7004, n7005,
         n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013, n7014, n7015,
         n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023, n7024, n7025,
         n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033, n7034, n7035,
         n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043, n7044, n7045,
         n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053, n7054, n7055,
         n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063, n7064, n7065,
         n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073, n7074, n7075,
         n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083, n7084, n7085,
         n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093, n7094, n7095,
         n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103, n7104, n7105,
         n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113, n7114, n7115,
         n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123, n7124, n7125,
         n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133, n7134, n7135,
         n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143, n7144, n7145,
         n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153, n7154, n7155,
         n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163, n7164, n7165,
         n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173, n7174, n7175,
         n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183, n7184, n7185,
         n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193, n7194, n7195,
         n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203, n7204, n7205,
         n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213, n7214, n7215,
         n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223, n7224, n7225,
         n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233, n7234, n7235,
         n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243, n7244, n7245,
         n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253, n7254, n7255,
         n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263, n7264, n7265,
         n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273, n7274, n7275,
         n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283, n7284, n7285,
         n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293, n7294, n7295,
         n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303, n7304, n7305,
         n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313, n7314, n7315,
         n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323, n7324, n7325,
         n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333, n7334, n7335,
         n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343, n7344, n7345,
         n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353, n7354, n7355,
         n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363, n7364, n7365,
         n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373, n7374, n7375,
         n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383, n7384, n7385,
         n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393, n7394, n7395,
         n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403, n7404, n7405,
         n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413, n7414, n7415,
         n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423, n7424, n7425,
         n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433, n7434, n7435,
         n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443, n7444, n7445,
         n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453, n7454, n7455,
         n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463, n7464, n7465,
         n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473, n7474, n7475,
         n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483, n7484, n7485,
         n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493, n7494, n7495,
         n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503, n7504, n7505,
         n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513, n7514, n7515,
         n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523, n7524, n7525,
         n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533, n7534, n7535,
         n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543, n7544, n7545,
         n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553, n7554, n7555,
         n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563, n7564, n7565,
         n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573, n7574, n7575,
         n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583, n7584, n7585,
         n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593, n7594, n7595,
         n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603, n7604, n7605,
         n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613, n7614, n7615,
         n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623, n7624, n7625,
         n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633, n7634, n7635,
         n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643, n7644, n7645,
         n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653, n7654, n7655,
         n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663, n7664, n7665,
         n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673, n7674, n7675,
         n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683, n7684, n7685,
         n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693, n7694, n7695,
         n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703, n7704, n7705,
         n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713, n7714, n7715,
         n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723, n7724, n7725,
         n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733, n7734, n7735,
         n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743, n7744, n7745,
         n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753, n7754, n7755,
         n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763, n7764, n7765,
         n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773, n7774, n7775,
         n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783, n7784, n7785,
         n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793, n7794, n7795,
         n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803, n7804, n7805,
         n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813, n7814, n7815,
         n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823, n7824, n7825,
         n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833, n7834, n7835,
         n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843, n7844, n7845,
         n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853, n7854, n7855,
         n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863, n7864, n7865,
         n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873, n7874, n7875,
         n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883, n7884, n7885,
         n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893, n7894, n7895,
         n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903, n7904, n7905,
         n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913, n7914, n7915,
         n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923, n7924, n7925,
         n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933, n7934, n7935,
         n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943, n7944, n7945,
         n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953, n7954, n7955,
         n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963, n7964, n7965,
         n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973, n7974, n7975,
         n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983, n7984, n7985,
         n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993, n7994, n7995,
         n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003, n8004, n8005,
         n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013, n8014, n8015,
         n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023, n8024, n8025,
         n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033, n8034, n8035,
         n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043, n8044, n8045,
         n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053, n8054, n8055,
         n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063, n8064, n8065,
         n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073, n8074, n8075,
         n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083, n8084, n8085,
         n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093, n8094, n8095,
         n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103, n8104, n8105,
         n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113, n8114, n8115,
         n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123, n8124, n8125,
         n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133, n8134, n8135,
         n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143, n8144, n8145,
         n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153, n8154, n8155,
         n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163, n8164, n8165,
         n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173, n8174, n8175,
         n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183, n8184, n8185,
         n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193, n8194, n8195,
         n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203, n8204, n8205,
         n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213, n8214, n8215,
         n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223, n8224, n8225,
         n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233, n8234, n8235,
         n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243, n8244, n8245,
         n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253, n8254, n8255,
         n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263, n8264, n8265,
         n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273, n8274, n8275,
         n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283, n8284, n8285,
         n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293, n8294, n8295,
         n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303, n8304, n8305,
         n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313, n8314, n8315,
         n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323, n8324, n8325,
         n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333, n8334, n8335,
         n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343, n8344, n8345,
         n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353, n8354, n8355,
         n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363, n8364, n8365,
         n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373, n8374, n8375,
         n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383, n8384, n8385,
         n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393, n8394, n8395,
         n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403, n8404, n8405,
         n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413, n8414, n8415,
         n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423, n8424, n8425,
         n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433, n8434, n8435,
         n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443, n8444, n8445,
         n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453, n8454, n8455,
         n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463, n8464, n8465,
         n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473, n8474, n8475,
         n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483, n8484, n8485,
         n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493, n8494, n8495,
         n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503, n8504, n8505,
         n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513, n8514, n8515,
         n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523, n8524, n8525,
         n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533, n8534, n8535,
         n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543, n8544, n8545,
         n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553, n8554, n8555,
         n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563, n8564, n8565,
         n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573, n8574, n8575,
         n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583, n8584, n8585,
         n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593, n8594, n8595,
         n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603, n8604, n8605,
         n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613, n8614, n8615,
         n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623, n8624, n8625,
         n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633, n8634, n8635,
         n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643, n8644, n8645,
         n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653, n8654, n8655,
         n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663, n8664, n8665,
         n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673, n8674, n8675,
         n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683, n8684, n8685,
         n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693, n8694, n8695,
         n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703, n8704, n8705,
         n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713, n8714, n8715,
         n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723, n8724, n8725,
         n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733, n8734, n8735,
         n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743, n8744, n8745,
         n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753, n8754, n8755,
         n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763, n8764, n8765,
         n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773, n8774, n8775,
         n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783, n8784, n8785,
         n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793, n8794, n8795,
         n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803, n8804, n8805,
         n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813, n8814, n8815,
         n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823, n8824, n8825,
         n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833, n8834, n8835,
         n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843, n8844, n8845,
         n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853, n8854, n8855,
         n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863, n8864, n8865,
         n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873, n8874, n8875,
         n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883, n8884, n8885,
         n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893, n8894, n8895,
         n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903, n8904, n8905,
         n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913, n8914, n8915,
         n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923, n8924, n8925,
         n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933, n8934, n8935,
         n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943, n8944, n8945,
         n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953, n8954, n8955,
         n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963, n8964, n8965,
         n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973, n8974, n8975,
         n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983, n8984, n8985,
         n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993, n8994, n8995,
         n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003, n9004, n9005,
         n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013, n9014, n9015,
         n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023, n9024, n9025,
         n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033, n9034, n9035,
         n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043, n9044, n9045,
         n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053, n9054, n9055,
         n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063, n9064, n9065,
         n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073, n9074, n9075,
         n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083, n9084, n9085,
         n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093, n9094, n9095,
         n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103, n9104, n9105,
         n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113, n9114, n9115,
         n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123, n9124, n9125,
         n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133, n9134, n9135,
         n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143, n9144, n9145,
         n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153, n9154, n9155,
         n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163, n9164, n9165,
         n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173, n9174, n9175,
         n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183, n9184, n9185,
         n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193, n9194, n9195,
         n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203, n9204, n9205,
         n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213, n9214, n9215,
         n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223, n9224, n9225,
         n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233, n9234, n9235,
         n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243, n9244, n9245,
         n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253, n9254, n9255,
         n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263, n9264, n9265,
         n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273, n9274, n9275,
         n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283, n9284, n9285,
         n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293, n9294, n9295,
         n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303, n9304, n9305,
         n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313, n9314, n9315,
         n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323, n9324, n9325,
         n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333, n9334, n9335,
         n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343, n9344, n9345,
         n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353, n9354, n9355,
         n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363, n9364, n9365,
         n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373, n9374, n9375,
         n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383, n9384, n9385,
         n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393, n9394, n9395,
         n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403, n9404, n9405,
         n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413, n9414, n9415,
         n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423, n9424, n9425,
         n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433, n9434, n9435,
         n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443, n9444, n9445,
         n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453, n9454, n9455,
         n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463, n9464, n9465,
         n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473, n9474, n9475,
         n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483, n9484, n9485,
         n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493, n9494, n9495,
         n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503, n9504, n9505,
         n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513, n9514, n9515,
         n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523, n9524, n9525,
         n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533, n9534, n9535,
         n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543, n9544, n9545,
         n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553, n9554, n9555,
         n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563, n9564, n9565,
         n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573, n9574, n9575,
         n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583, n9584, n9585,
         n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593, n9594, n9595,
         n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603, n9604, n9605,
         n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613, n9614, n9615,
         n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623, n9624, n9625,
         n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633, n9634, n9635,
         n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643, n9644, n9645,
         n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653, n9654, n9655,
         n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663, n9664, n9665,
         n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673, n9674, n9675,
         n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683, n9684, n9685,
         n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693, n9694, n9695,
         n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703, n9704, n9705,
         n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713, n9714, n9715,
         n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723, n9724, n9725,
         n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733, n9734, n9735,
         n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743, n9744, n9745,
         n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753, n9754, n9755,
         n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763, n9764, n9765,
         n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773, n9774, n9775,
         n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783, n9784, n9785,
         n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793, n9794, n9795,
         n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803, n9804, n9805,
         n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813, n9814, n9815,
         n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823, n9824, n9825,
         n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833, n9834, n9835,
         n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843, n9844, n9845,
         n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853, n9854, n9855,
         n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863, n9864, n9865,
         n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873, n9874, n9875,
         n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883, n9884, n9885,
         n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893, n9894, n9895,
         n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903, n9904, n9905,
         n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913, n9914, n9915,
         n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923, n9924, n9925,
         n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933, n9934, n9935,
         n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943, n9944, n9945,
         n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953, n9954, n9955,
         n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963, n9964, n9965,
         n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973, n9974, n9975,
         n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983, n9984, n9985,
         n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993, n9994, n9995,
         n9996, n9997, n9998, n9999, n10000, n10001, n10002, n10003, n10004,
         n10005, n10006, n10007, n10008, n10009, n10010, n10011, n10012,
         n10013, n10014, n10015, n10016, n10017, n10018, n10019, n10020,
         n10021, n10022, n10023, n10024, n10025, n10026, n10027, n10028,
         n10029, n10030, n10031, n10032, n10033, n10034, n10035, n10036,
         n10037, n10038, n10039, n10040, n10041, n10042, n10043, n10044,
         n10045, n10046, n10047, n10048, n10049, n10050, n10051, n10052,
         n10053, n10054, n10055, n10056, n10057, n10058, n10059, n10060,
         n10061, n10062, n10063, n10064, n10065, n10066, n10067, n10068,
         n10069, n10070, n10071, n10072, n10073, n10074, n10075, n10076,
         n10077, n10078, n10079, n10080, n10081, n10082, n10083, n10084,
         n10085, n10086, n10087, n10088, n10089, n10090, n10091, n10092,
         n10093, n10094, n10095, n10096, n10097, n10098, n10099, n10100,
         n10101, n10102, n10103, n10104, n10105, n10106, n10107, n10108,
         n10109, n10110, n10111, n10112, n10113, n10114, n10115, n10116,
         n10117, n10118, n10119, n10120, n10121, n10122, n10123, n10124,
         n10125, n10126, n10127, n10128, n10129, n10130, n10131, n10132,
         n10133, n10134, n10135, n10136, n10137, n10138, n10139, n10140,
         n10141, n10142, n10143, n10144, n10145, n10146, n10147, n10148,
         n10149, n10150, n10151, n10152, n10153, n10154, n10155, n10156,
         n10157, n10158, n10159, n10160, n10161, n10162, n10163, n10164;
  wire   [29:0] ICACHE_addr;
  wire   [31:0] DCACHE_rdata;

  NOR4X6 \D_cache/U1793  ( .A(\D_cache/n528 ), .B(\D_cache/n529 ), .C(
        \D_cache/n530 ), .D(\D_cache/n531 ), .Y(\D_cache/n527 ) );
  DFFRX4 \i_MIPS/PC/PC_o_reg[4]  ( .D(\i_MIPS/PC/n38 ), .CK(clk), .RN(n4066), 
        .Q(ICACHE_addr[2]), .QN(\i_MIPS/PC/n6 ) );
  DFFRX4 \i_MIPS/PC/PC_o_reg[5]  ( .D(\i_MIPS/PC/n39 ), .CK(clk), .RN(n4066), 
        .Q(ICACHE_addr[3]), .QN(\i_MIPS/PC/n7 ) );
  DFFRX4 \i_MIPS/PC/PC_o_reg[6]  ( .D(\i_MIPS/PC/n40 ), .CK(clk), .RN(n4066), 
        .Q(ICACHE_addr[4]), .QN(\i_MIPS/PC/n8 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[1]  ( .D(\i_MIPS/n526 ), .CK(clk), .RN(n4062), .Q(
        \i_MIPS/EX_MEM_1 ), .QN(\i_MIPS/n336 ) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[21]  ( .D(\i_MIPS/PC/n55 ), .CK(clk), .RN(n4067), 
        .Q(ICACHE_addr[19]), .QN(\i_MIPS/PC/n23 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[50]  ( .D(\i_MIPS/n419 ), .CK(clk), .RN(n4051), .Q(
        \i_MIPS/ID_EX[50] ), .QN(\i_MIPS/n291 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[22]  ( .D(\i_MIPS/n452 ), .CK(clk), .RN(n4054), 
        .Q(n10311), .QN(n1625) );
  DFFRX1 \i_MIPS/EX_MEM_reg[16]  ( .D(\i_MIPS/n458 ), .CK(clk), .RN(n4054), 
        .Q(n10317), .QN(n1622) );
  DFFRX1 \i_MIPS/EX_MEM_reg[30]  ( .D(\i_MIPS/n444 ), .CK(clk), .RN(n4053), 
        .Q(n10303), .QN(n1089) );
  DFFRX1 \i_MIPS/EX_MEM_reg[15]  ( .D(\i_MIPS/n459 ), .CK(clk), .RN(n4054), 
        .Q(n10318), .QN(n1626) );
  DFFRX1 \i_MIPS/EX_MEM_reg[26]  ( .D(\i_MIPS/n448 ), .CK(clk), .RN(n4053), 
        .Q(n10307), .QN(n1088) );
  DFFRX1 \i_MIPS/EX_MEM_reg[34]  ( .D(\i_MIPS/n440 ), .CK(clk), .RN(n4053), 
        .Q(n10299), .QN(n1092) );
  DFFRX1 \i_MIPS/EX_MEM_reg[13]  ( .D(\i_MIPS/n461 ), .CK(clk), .RN(n4054), 
        .Q(n10320), .QN(n1623) );
  DFFRX1 \i_MIPS/EX_MEM_reg[25]  ( .D(\i_MIPS/n449 ), .CK(clk), .RN(n4053), 
        .Q(n10308), .QN(n1087) );
  DFFRX1 \i_MIPS/EX_MEM_reg[29]  ( .D(\i_MIPS/n445 ), .CK(clk), .RN(n4053), 
        .Q(n10304), .QN(n1090) );
  DFFRX1 \i_MIPS/EX_MEM_reg[14]  ( .D(\i_MIPS/n460 ), .CK(clk), .RN(n4054), 
        .Q(n10319), .QN(n1624) );
  DFFRX1 \i_MIPS/EX_MEM_reg[27]  ( .D(\i_MIPS/n447 ), .CK(clk), .RN(n4053), 
        .Q(n10306), .QN(n1091) );
  DFFRX1 \i_MIPS/EX_MEM_reg[19]  ( .D(\i_MIPS/n455 ), .CK(clk), .RN(n4054), 
        .Q(n10314), .QN(n1071) );
  DFFRX1 \i_MIPS/EX_MEM_reg[21]  ( .D(\i_MIPS/n453 ), .CK(clk), .RN(n4054), 
        .Q(n10312), .QN(n1070) );
  DFFRX1 \i_MIPS/IF_ID_reg[38]  ( .D(\i_MIPS/N61 ), .CK(clk), .RN(n4059), .Q(
        \i_MIPS/Sign_Extend_ID[6] ), .QN(\i_MIPS/n218 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[39]  ( .D(\i_MIPS/N62 ), .CK(clk), .RN(n4059), .QN(
        \i_MIPS/n219 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[40]  ( .D(\i_MIPS/N63 ), .CK(clk), .RN(n4059), .Q(
        \i_MIPS/Sign_Extend_ID[8] ), .QN(\i_MIPS/n220 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[41]  ( .D(\i_MIPS/N64 ), .CK(clk), .RN(n4059), .QN(
        \i_MIPS/n221 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[42]  ( .D(\i_MIPS/N65 ), .CK(clk), .RN(n4059), .QN(
        \i_MIPS/n222 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[43]  ( .D(\i_MIPS/N66 ), .CK(clk), .RN(n4059), .QN(
        \i_MIPS/n223 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[44]  ( .D(\i_MIPS/N67 ), .CK(clk), .RN(n4060), .QN(
        \i_MIPS/n224 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[45]  ( .D(\i_MIPS/N68 ), .CK(clk), .RN(n4060), .QN(
        \i_MIPS/n225 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[46]  ( .D(\i_MIPS/N69 ), .CK(clk), .RN(n4060), .QN(
        \i_MIPS/n226 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[47]  ( .D(\i_MIPS/N70 ), .CK(clk), .RN(n4060), .Q(
        \i_MIPS/Sign_Extend_ID[31] ), .QN(\i_MIPS/n227 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[27]  ( .D(\i_MIPS/N50 ), .CK(clk), .RN(n4045), .QN(
        \i_MIPS/n207 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[26]  ( .D(\i_MIPS/N49 ), .CK(clk), .RN(n4045), .QN(
        \i_MIPS/n206 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[25]  ( .D(\i_MIPS/N48 ), .CK(clk), .RN(n4045), .QN(
        \i_MIPS/n205 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[24]  ( .D(\i_MIPS/N47 ), .CK(clk), .RN(n4045), .QN(
        \i_MIPS/n204 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[23]  ( .D(\i_MIPS/N46 ), .CK(clk), .RN(n4045), .QN(
        \i_MIPS/n203 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[22]  ( .D(\i_MIPS/N45 ), .CK(clk), .RN(n4045), .QN(
        \i_MIPS/n202 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[21]  ( .D(\i_MIPS/N44 ), .CK(clk), .RN(n4045), .QN(
        \i_MIPS/n201 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[20]  ( .D(\i_MIPS/N43 ), .CK(clk), .RN(n4045), .QN(
        \i_MIPS/n200 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[19]  ( .D(\i_MIPS/N42 ), .CK(clk), .RN(n4045), .QN(
        \i_MIPS/n199 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[18]  ( .D(\i_MIPS/N41 ), .CK(clk), .RN(n4045), .QN(
        \i_MIPS/n198 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[17]  ( .D(\i_MIPS/N40 ), .CK(clk), .RN(n4045), .QN(
        \i_MIPS/n197 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[16]  ( .D(\i_MIPS/N39 ), .CK(clk), .RN(n4045), .QN(
        \i_MIPS/n196 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[15]  ( .D(\i_MIPS/N38 ), .CK(clk), .RN(n4046), .QN(
        \i_MIPS/n195 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[14]  ( .D(\i_MIPS/N37 ), .CK(clk), .RN(n4046), .QN(
        \i_MIPS/n194 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[13]  ( .D(\i_MIPS/N36 ), .CK(clk), .RN(n4046), .QN(
        \i_MIPS/n193 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[12]  ( .D(\i_MIPS/N35 ), .CK(clk), .RN(n4046), .QN(
        \i_MIPS/n192 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[11]  ( .D(\i_MIPS/N34 ), .CK(clk), .RN(n4046), .QN(
        \i_MIPS/n191 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[10]  ( .D(\i_MIPS/N33 ), .CK(clk), .RN(n4046), .QN(
        \i_MIPS/n190 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[9]  ( .D(\i_MIPS/N32 ), .CK(clk), .RN(n4046), .QN(
        \i_MIPS/n189 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[8]  ( .D(\i_MIPS/N31 ), .CK(clk), .RN(n4046), .QN(
        \i_MIPS/n188 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[7]  ( .D(\i_MIPS/N30 ), .CK(clk), .RN(n4046), .QN(
        \i_MIPS/n187 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[6]  ( .D(\i_MIPS/N29 ), .CK(clk), .RN(n4046), .QN(
        \i_MIPS/n186 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[5]  ( .D(\i_MIPS/N28 ), .CK(clk), .RN(n4046), .QN(
        \i_MIPS/n185 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[4]  ( .D(\i_MIPS/N27 ), .CK(clk), .RN(n4046), .QN(
        \i_MIPS/n184 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[3]  ( .D(\i_MIPS/N26 ), .CK(clk), .RN(n4047), .QN(
        \i_MIPS/n183 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[2]  ( .D(\i_MIPS/N25 ), .CK(clk), .RN(n4047), .QN(
        \i_MIPS/n182 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[92]  ( .D(\i_MIPS/N115 ), .CK(clk), .RN(n4042), .Q(
        \i_MIPS/IF_ID[92] ), .QN(\i_MIPS/n174 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[91]  ( .D(\i_MIPS/N114 ), .CK(clk), .RN(n4042), .Q(
        \i_MIPS/IF_ID[91] ), .QN(\i_MIPS/n173 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[90]  ( .D(\i_MIPS/N113 ), .CK(clk), .RN(n4042), .Q(
        \i_MIPS/IF_ID[90] ), .QN(\i_MIPS/n172 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[89]  ( .D(\i_MIPS/N112 ), .CK(clk), .RN(n4042), .Q(
        \i_MIPS/IF_ID[89] ), .QN(\i_MIPS/n171 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[88]  ( .D(\i_MIPS/N111 ), .CK(clk), .RN(n4042), .Q(
        \i_MIPS/IF_ID[88] ), .QN(\i_MIPS/n170 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[87]  ( .D(\i_MIPS/N110 ), .CK(clk), .RN(n4042), .Q(
        \i_MIPS/IF_ID[87] ), .QN(\i_MIPS/n169 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[86]  ( .D(\i_MIPS/N109 ), .CK(clk), .RN(n4042), .Q(
        \i_MIPS/IF_ID[86] ), .QN(\i_MIPS/n168 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[84]  ( .D(\i_MIPS/N107 ), .CK(clk), .RN(n4043), .Q(
        \i_MIPS/IF_ID[84] ), .QN(\i_MIPS/n166 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[83]  ( .D(\i_MIPS/N106 ), .CK(clk), .RN(n4043), .Q(
        \i_MIPS/IF_ID[83] ), .QN(\i_MIPS/n165 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[82]  ( .D(\i_MIPS/N105 ), .CK(clk), .RN(n4043), .Q(
        \i_MIPS/IF_ID[82] ), .QN(\i_MIPS/n164 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[81]  ( .D(\i_MIPS/N104 ), .CK(clk), .RN(n4043), .Q(
        \i_MIPS/IF_ID[81] ), .QN(\i_MIPS/n163 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[80]  ( .D(\i_MIPS/N103 ), .CK(clk), .RN(n4043), .Q(
        \i_MIPS/IF_ID[80] ), .QN(\i_MIPS/n162 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[79]  ( .D(\i_MIPS/N102 ), .CK(clk), .RN(n4043), .Q(
        \i_MIPS/IF_ID[79] ), .QN(\i_MIPS/n161 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[78]  ( .D(\i_MIPS/N101 ), .CK(clk), .RN(n4043), .Q(
        \i_MIPS/IF_ID[78] ), .QN(\i_MIPS/n160 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[77]  ( .D(\i_MIPS/N100 ), .CK(clk), .RN(n4043), .Q(
        \i_MIPS/IF_ID[77] ), .QN(\i_MIPS/n159 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[76]  ( .D(\i_MIPS/N99 ), .CK(clk), .RN(n4043), .Q(
        \i_MIPS/IF_ID[76] ), .QN(\i_MIPS/n245 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[75]  ( .D(\i_MIPS/N98 ), .CK(clk), .RN(n4043), .Q(
        \i_MIPS/IF_ID[75] ), .QN(\i_MIPS/n244 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[74]  ( .D(\i_MIPS/N97 ), .CK(clk), .RN(n4043), .Q(
        \i_MIPS/IF_ID[74] ), .QN(\i_MIPS/n243 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[73]  ( .D(\i_MIPS/N96 ), .CK(clk), .RN(n4044), .Q(
        \i_MIPS/IF_ID[73] ), .QN(\i_MIPS/n242 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[72]  ( .D(\i_MIPS/N95 ), .CK(clk), .RN(n4044), .Q(
        \i_MIPS/IF_ID[72] ), .QN(\i_MIPS/n241 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[71]  ( .D(\i_MIPS/N94 ), .CK(clk), .RN(n4044), .Q(
        \i_MIPS/IF_ID[71] ), .QN(\i_MIPS/n240 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[70]  ( .D(\i_MIPS/N93 ), .CK(clk), .RN(n4044), .Q(
        \i_MIPS/IF_ID[70] ), .QN(\i_MIPS/n239 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[69]  ( .D(\i_MIPS/N92 ), .CK(clk), .RN(n4044), .Q(
        \i_MIPS/IF_ID[69] ), .QN(\i_MIPS/n238 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[68]  ( .D(\i_MIPS/N91 ), .CK(clk), .RN(n4044), .Q(
        \i_MIPS/IF_ID[68] ), .QN(\i_MIPS/n237 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[67]  ( .D(\i_MIPS/N90 ), .CK(clk), .RN(n4044), .Q(
        \i_MIPS/IF_ID[67] ), .QN(\i_MIPS/n236 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[96]  ( .D(\i_MIPS/N119 ), .CK(clk), .RN(n4042), .Q(
        \i_MIPS/IF_ID[96] ), .QN(\i_MIPS/n178 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[94]  ( .D(\i_MIPS/N117 ), .CK(clk), .RN(n4042), .Q(
        \i_MIPS/IF_ID[94] ), .QN(\i_MIPS/n176 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[93]  ( .D(\i_MIPS/N116 ), .CK(clk), .RN(n4042), .Q(
        \i_MIPS/IF_ID[93] ), .QN(\i_MIPS/n175 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[65]  ( .D(\i_MIPS/N88 ), .CK(clk), .RN(n4044), .Q(
        \i_MIPS/IF_ID[65] ), .QN(\i_MIPS/n234 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[31]  ( .D(\i_MIPS/N54 ), .CK(clk), .RN(n4042), .Q(
        \i_MIPS/IF_ID_31 ), .QN(\i_MIPS/n211 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[29]  ( .D(\i_MIPS/N52 ), .CK(clk), .RN(n4044), .Q(
        \i_MIPS/IF_ID_29 ), .QN(\i_MIPS/n209 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[28]  ( .D(\i_MIPS/N51 ), .CK(clk), .RN(n4044), .Q(
        \i_MIPS/IF_ID_28 ), .QN(\i_MIPS/n208 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[0]  ( .D(\i_MIPS/N23 ), .CK(clk), .RN(n4047), .Q(
        \i_MIPS/IF_ID_0 ), .QN(\i_MIPS/n180 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[4]  ( .D(\i_MIPS/n480 ), .CK(clk), .RN(n4056), .Q(
        n1894), .QN(\i_MIPS/n311 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[1]  ( .D(\i_MIPS/n527 ), .CK(clk), .RN(n4062), .Q(
        n1893), .QN(\i_MIPS/n337 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[116]  ( .D(\i_MIPS/n530 ), .CK(clk), .RN(n4063), 
        .Q(n1892), .QN(\i_MIPS/n339 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[3]  ( .D(\i_MIPS/n525 ), .CK(clk), .RN(n4062), .Q(
        \i_MIPS/ID_EX_3 ), .QN(\i_MIPS/n335 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[36]  ( .D(\i_MIPS/N59 ), .CK(clk), .RN(n4059), .Q(
        \i_MIPS/Sign_Extend_ID[4] ), .QN(\i_MIPS/n216 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[34]  ( .D(\i_MIPS/N57 ), .CK(clk), .RN(n4059), .Q(
        \i_MIPS/Sign_Extend_ID[2] ), .QN(\i_MIPS/n214 ) );
  DFFSX1 \i_MIPS/Pred_1bit/current_state_reg  ( .D(\i_MIPS/Pred_1bit/n2 ), 
        .CK(clk), .SN(n4360), .Q(\i_MIPS/Pred_1bit/current_state ) );
  DFFRX1 \i_MIPS/IF_ID_reg[33]  ( .D(\i_MIPS/N56 ), .CK(clk), .RN(n4059), .Q(
        \i_MIPS/Sign_Extend_ID[1] ), .QN(\i_MIPS/n213 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[35]  ( .D(\i_MIPS/N58 ), .CK(clk), .RN(n4059), .Q(
        \i_MIPS/Sign_Extend_ID[3] ), .QN(\i_MIPS/n215 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[37]  ( .D(\i_MIPS/N60 ), .CK(clk), .RN(n4059), .Q(
        \i_MIPS/Sign_Extend_ID[5] ), .QN(\i_MIPS/n217 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[32]  ( .D(\i_MIPS/N55 ), .CK(clk), .RN(n4063), .Q(
        \i_MIPS/Sign_Extend_ID[0] ), .QN(\i_MIPS/n212 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[64]  ( .D(\i_MIPS/N87 ), .CK(clk), .RN(n4047), .Q(
        \i_MIPS/IF_ID[64] ), .QN(\i_MIPS/n233 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[97]  ( .D(\i_MIPS/N120 ), .CK(clk), .RN(n4047), .Q(
        \i_MIPS/IF_ID[97] ), .QN(n1627) );
  DFFRX1 \i_MIPS/Register/register_reg[31][0]  ( .D(n8804), .CK(clk), .RN(
        n4068), .QN(n70) );
  DFFRX1 \i_MIPS/Register/register_reg[31][1]  ( .D(n8803), .CK(clk), .RN(
        n4068), .QN(n206) );
  DFFRX1 \i_MIPS/Register/register_reg[31][2]  ( .D(n8802), .CK(clk), .RN(
        n4068), .QN(n200) );
  DFFRX1 \i_MIPS/Register/register_reg[31][3]  ( .D(n8801), .CK(clk), .RN(
        n4068), .QN(n201) );
  DFFRX1 \i_MIPS/Register/register_reg[31][4]  ( .D(n8800), .CK(clk), .RN(
        n4069), .QN(n197) );
  DFFRX1 \i_MIPS/Register/register_reg[31][5]  ( .D(n8799), .CK(clk), .RN(
        n4069), .QN(n207) );
  DFFRX1 \i_MIPS/Register/register_reg[31][6]  ( .D(n8798), .CK(clk), .RN(
        n4069), .QN(n199) );
  DFFRX1 \i_MIPS/Register/register_reg[31][7]  ( .D(n8797), .CK(clk), .RN(
        n4069), .QN(n61) );
  DFFRX1 \i_MIPS/Register/register_reg[31][9]  ( .D(n8795), .CK(clk), .RN(
        n4069), .QN(n57) );
  DFFRX1 \i_MIPS/Register/register_reg[31][10]  ( .D(n8794), .CK(clk), .RN(
        n4069), .QN(n198) );
  DFFRX1 \i_MIPS/Register/register_reg[31][11]  ( .D(n8793), .CK(clk), .RN(
        n4069), .QN(n60) );
  DFFRX1 \i_MIPS/Register/register_reg[31][12]  ( .D(n8792), .CK(clk), .RN(
        n4069), .QN(n209) );
  DFFRX1 \i_MIPS/Register/register_reg[31][13]  ( .D(n8791), .CK(clk), .RN(
        n4069), .QN(n58) );
  DFFRX1 \i_MIPS/Register/register_reg[31][14]  ( .D(n8790), .CK(clk), .RN(
        n4069), .QN(n59) );
  DFFRX1 \i_MIPS/Register/register_reg[31][15]  ( .D(n8789), .CK(clk), .RN(
        n4069), .QN(n62) );
  DFFRX1 \i_MIPS/Register/register_reg[31][16]  ( .D(n8788), .CK(clk), .RN(
        n4070), .QN(n63) );
  DFFRX1 \i_MIPS/Register/register_reg[31][17]  ( .D(n8787), .CK(clk), .RN(
        n4070), .QN(n65) );
  DFFRX1 \i_MIPS/Register/register_reg[31][18]  ( .D(n8786), .CK(clk), .RN(
        n4070), .QN(n64) );
  DFFRX1 \i_MIPS/Register/register_reg[31][19]  ( .D(n8785), .CK(clk), .RN(
        n4070), .QN(n194) );
  DFFRX1 \i_MIPS/Register/register_reg[31][20]  ( .D(n8784), .CK(clk), .RN(
        n4070), .QN(n204) );
  DFFRX1 \i_MIPS/Register/register_reg[31][21]  ( .D(n8783), .CK(clk), .RN(
        n4070), .QN(n205) );
  DFFRX1 \i_MIPS/Register/register_reg[31][22]  ( .D(n8782), .CK(clk), .RN(
        n4070), .QN(n202) );
  DFFRX1 \i_MIPS/Register/register_reg[31][23]  ( .D(n8781), .CK(clk), .RN(
        n4070), .QN(n203) );
  DFFRX1 \i_MIPS/Register/register_reg[31][24]  ( .D(n8780), .CK(clk), .RN(
        n4070), .QN(n208) );
  DFFRX1 \i_MIPS/Register/register_reg[31][25]  ( .D(n8779), .CK(clk), .RN(
        n4070), .QN(n193) );
  DFFRX1 \i_MIPS/Register/register_reg[31][26]  ( .D(n8778), .CK(clk), .RN(
        n4070), .QN(n71) );
  DFFRX1 \i_MIPS/Register/register_reg[31][27]  ( .D(n8777), .CK(clk), .RN(
        n4070), .QN(n195) );
  DFFRX1 \i_MIPS/Register/register_reg[31][28]  ( .D(n8776), .CK(clk), .RN(
        n4071), .QN(n67) );
  DFFRX1 \i_MIPS/Register/register_reg[31][29]  ( .D(n8775), .CK(clk), .RN(
        n4071), .QN(n69) );
  DFFRX1 \i_MIPS/Register/register_reg[31][30]  ( .D(n8774), .CK(clk), .RN(
        n4071), .QN(n68) );
  DFFRX1 \i_MIPS/Register/register_reg[31][31]  ( .D(n8773), .CK(clk), .RN(
        n4071), .QN(n66) );
  DFFRX1 \i_MIPS/EX_MEM_reg[74]  ( .D(\i_MIPS/n529 ), .CK(clk), .RN(n4063), 
        .Q(\i_MIPS/EX_MEM_74 ), .QN(\i_MIPS/n338 ) );
  DFFRX1 \i_MIPS/Register/register_reg[29][0]  ( .D(\i_MIPS/Register/n180 ), 
        .CK(clk), .RN(n4074), .Q(\i_MIPS/Register/register[29][0] ), .QN(n278)
         );
  DFFRX1 \i_MIPS/Register/register_reg[27][0]  ( .D(\i_MIPS/Register/n244 ), 
        .CK(clk), .RN(n4079), .Q(\i_MIPS/Register/register[27][0] ), .QN(n277)
         );
  DFFRX1 \i_MIPS/Register/register_reg[27][1]  ( .D(\i_MIPS/Register/n245 ), 
        .CK(clk), .RN(n4079), .Q(\i_MIPS/Register/register[27][1] ), .QN(n272)
         );
  DFFRX1 \i_MIPS/Register/register_reg[25][0]  ( .D(\i_MIPS/Register/n308 ), 
        .CK(clk), .RN(n4084), .Q(\i_MIPS/Register/register[25][0] ), .QN(n228)
         );
  DFFRX1 \i_MIPS/Register/register_reg[23][0]  ( .D(\i_MIPS/Register/n372 ), 
        .CK(clk), .RN(n4090), .Q(\i_MIPS/Register/register[23][0] ), .QN(n1171) );
  DFFRX1 \i_MIPS/Register/register_reg[23][1]  ( .D(\i_MIPS/Register/n373 ), 
        .CK(clk), .RN(n4090), .Q(\i_MIPS/Register/register[23][1] ), .QN(n1165) );
  DFFRX1 \i_MIPS/Register/register_reg[21][0]  ( .D(\i_MIPS/Register/n436 ), 
        .CK(clk), .RN(n4095), .Q(\i_MIPS/Register/register[21][0] ), .QN(n1173) );
  DFFRX1 \i_MIPS/Register/register_reg[19][0]  ( .D(\i_MIPS/Register/n500 ), 
        .CK(clk), .RN(n4100), .Q(\i_MIPS/Register/register[19][0] ), .QN(n1172) );
  DFFRX1 \i_MIPS/Register/register_reg[17][0]  ( .D(\i_MIPS/Register/n564 ), 
        .CK(clk), .RN(n4106), .Q(\i_MIPS/Register/register[17][0] ), .QN(n1348) );
  DFFRX1 \i_MIPS/Register/register_reg[15][0]  ( .D(\i_MIPS/Register/n628 ), 
        .CK(clk), .RN(n4111), .Q(\i_MIPS/Register/register[15][0] ), .QN(n279)
         );
  DFFRX1 \i_MIPS/Register/register_reg[15][1]  ( .D(\i_MIPS/Register/n629 ), 
        .CK(clk), .RN(n4111), .Q(\i_MIPS/Register/register[15][1] ), .QN(n274)
         );
  DFFRX1 \i_MIPS/Register/register_reg[13][0]  ( .D(\i_MIPS/Register/n692 ), 
        .CK(clk), .RN(n4116), .Q(\i_MIPS/Register/register[13][0] ), .QN(n281)
         );
  DFFRX1 \i_MIPS/Register/register_reg[11][0]  ( .D(\i_MIPS/Register/n756 ), 
        .CK(clk), .RN(n4122), .Q(\i_MIPS/Register/register[11][0] ), .QN(n280)
         );
  DFFRX1 \i_MIPS/Register/register_reg[11][1]  ( .D(\i_MIPS/Register/n757 ), 
        .CK(clk), .RN(n4122), .Q(\i_MIPS/Register/register[11][1] ), .QN(n275)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][0]  ( .D(\i_MIPS/Register/n820 ), 
        .CK(clk), .RN(n4127), .Q(\i_MIPS/Register/register[9][0] ), .QN(n395)
         );
  DFFRX1 \i_MIPS/Register/register_reg[7][0]  ( .D(\i_MIPS/Register/n884 ), 
        .CK(clk), .RN(n4132), .Q(\i_MIPS/Register/register[7][0] ), .QN(n1174)
         );
  DFFRX1 \i_MIPS/Register/register_reg[7][1]  ( .D(\i_MIPS/Register/n885 ), 
        .CK(clk), .RN(n4132), .Q(\i_MIPS/Register/register[7][1] ), .QN(n1168)
         );
  DFFRX1 \i_MIPS/Register/register_reg[5][0]  ( .D(\i_MIPS/Register/n948 ), 
        .CK(clk), .RN(n4138), .Q(\i_MIPS/Register/register[5][0] ), .QN(n1176)
         );
  DFFRX1 \i_MIPS/Register/register_reg[5][24]  ( .D(\i_MIPS/Register/n972 ), 
        .CK(clk), .RN(n4140), .Q(\i_MIPS/Register/register[5][24] ), .QN(n1212) );
  DFFRX1 \i_MIPS/Register/register_reg[5][26]  ( .D(\i_MIPS/Register/n974 ), 
        .CK(clk), .RN(n4140), .Q(\i_MIPS/Register/register[5][26] ), .QN(n1218) );
  DFFRX1 \i_MIPS/Register/register_reg[3][0]  ( .D(\i_MIPS/Register/n1012 ), 
        .CK(clk), .RN(n4143), .Q(\i_MIPS/Register/register[3][0] ), .QN(n1175)
         );
  DFFRX1 \i_MIPS/Register/register_reg[3][12]  ( .D(\i_MIPS/Register/n1024 ), 
        .CK(clk), .RN(n4144), .Q(\i_MIPS/Register/register[3][12] ), .QN(n1117) );
  DFFRX1 \i_MIPS/Register/register_reg[3][24]  ( .D(\i_MIPS/Register/n1036 ), 
        .CK(clk), .RN(n4145), .Q(\i_MIPS/Register/register[3][24] ), .QN(n1211) );
  DFFRX1 \i_MIPS/Register/register_reg[3][26]  ( .D(\i_MIPS/Register/n1038 ), 
        .CK(clk), .RN(n4145), .Q(\i_MIPS/Register/register[3][26] ), .QN(n1217) );
  DFFRX1 \i_MIPS/Register/register_reg[1][0]  ( .D(\i_MIPS/Register/n1076 ), 
        .CK(clk), .RN(n4148), .Q(\i_MIPS/Register/register[1][0] ), .QN(n1309)
         );
  DFFRX1 \i_MIPS/Register/register_reg[1][24]  ( .D(\i_MIPS/Register/n1100 ), 
        .CK(clk), .RN(n4150), .Q(\i_MIPS/Register/register[1][24] ), .QN(n1321) );
  DFFRX1 \i_MIPS/Register/register_reg[1][26]  ( .D(\i_MIPS/Register/n1102 ), 
        .CK(clk), .RN(n4150), .Q(\i_MIPS/Register/register[1][26] ), .QN(n1323) );
  DFFRX1 \D_cache/cache_reg[3][15]  ( .D(\D_cache/n1673 ), .CK(clk), .RN(n4164), .Q(\D_cache/cache[3][15] ) );
  DFFRX1 \D_cache/cache_reg[3][16]  ( .D(\D_cache/n1665 ), .CK(clk), .RN(n4164), .Q(\D_cache/cache[3][16] ) );
  DFFRX1 \D_cache/cache_reg[7][16]  ( .D(\D_cache/n1661 ), .CK(clk), .RN(n4165), .Q(\D_cache/cache[7][16] ) );
  DFFRX1 \D_cache/cache_reg[3][29]  ( .D(\D_cache/n1561 ), .CK(clk), .RN(n4173), .Q(\D_cache/cache[3][29] ) );
  DFFRX1 \D_cache/cache_reg[7][29]  ( .D(\D_cache/n1557 ), .CK(clk), .RN(n4173), .Q(\D_cache/cache[7][29] ) );
  DFFRX1 \D_cache/cache_reg[3][30]  ( .D(\D_cache/n1553 ), .CK(clk), .RN(n4174), .Q(\D_cache/cache[3][30] ) );
  DFFRX1 \D_cache/cache_reg[7][30]  ( .D(\D_cache/n1549 ), .CK(clk), .RN(n4174), .Q(\D_cache/cache[7][30] ) );
  DFFRX1 \D_cache/cache_reg[3][32]  ( .D(\D_cache/n1537 ), .CK(clk), .RN(n4175), .Q(\D_cache/cache[3][32] ) );
  DFFRX1 \D_cache/cache_reg[7][32]  ( .D(\D_cache/n1533 ), .CK(clk), .RN(n4175), .Q(\D_cache/cache[7][32] ) );
  DFFRX1 \D_cache/cache_reg[3][33]  ( .D(\D_cache/n1529 ), .CK(clk), .RN(n4176), .Q(\D_cache/cache[3][33] ) );
  DFFRX1 \D_cache/cache_reg[7][33]  ( .D(\D_cache/n1525 ), .CK(clk), .RN(n4176), .Q(\D_cache/cache[7][33] ) );
  DFFRX1 \D_cache/cache_reg[3][34]  ( .D(\D_cache/n1521 ), .CK(clk), .RN(n4176), .Q(\D_cache/cache[3][34] ) );
  DFFRX1 \D_cache/cache_reg[7][34]  ( .D(\D_cache/n1517 ), .CK(clk), .RN(n4177), .Q(\D_cache/cache[7][34] ) );
  DFFRX1 \D_cache/cache_reg[3][35]  ( .D(\D_cache/n1513 ), .CK(clk), .RN(n4177), .Q(\D_cache/cache[3][35] ) );
  DFFRX1 \D_cache/cache_reg[7][35]  ( .D(\D_cache/n1509 ), .CK(clk), .RN(n4177), .Q(\D_cache/cache[7][35] ) );
  DFFRX1 \D_cache/cache_reg[3][36]  ( .D(\D_cache/n1505 ), .CK(clk), .RN(n4178), .Q(\D_cache/cache[3][36] ) );
  DFFRX1 \D_cache/cache_reg[7][36]  ( .D(\D_cache/n1501 ), .CK(clk), .RN(n4178), .Q(\D_cache/cache[7][36] ) );
  DFFRX1 \D_cache/cache_reg[3][37]  ( .D(\D_cache/n1497 ), .CK(clk), .RN(n4178), .Q(\D_cache/cache[3][37] ) );
  DFFRX1 \D_cache/cache_reg[7][37]  ( .D(\D_cache/n1493 ), .CK(clk), .RN(n4179), .Q(\D_cache/cache[7][37] ) );
  DFFRX1 \D_cache/cache_reg[3][38]  ( .D(\D_cache/n1489 ), .CK(clk), .RN(n4179), .Q(\D_cache/cache[3][38] ) );
  DFFRX1 \D_cache/cache_reg[7][38]  ( .D(\D_cache/n1485 ), .CK(clk), .RN(n4179), .Q(\D_cache/cache[7][38] ) );
  DFFRX1 \D_cache/cache_reg[3][40]  ( .D(\D_cache/n1473 ), .CK(clk), .RN(n4180), .Q(\D_cache/cache[3][40] ) );
  DFFRX1 \D_cache/cache_reg[7][40]  ( .D(\D_cache/n1469 ), .CK(clk), .RN(n4181), .Q(\D_cache/cache[7][40] ) );
  DFFRX1 \D_cache/cache_reg[3][42]  ( .D(\D_cache/n1457 ), .CK(clk), .RN(n4182), .Q(\D_cache/cache[3][42] ) );
  DFFRX1 \D_cache/cache_reg[7][42]  ( .D(\D_cache/n1453 ), .CK(clk), .RN(n4182), .Q(\D_cache/cache[7][42] ) );
  DFFRX1 \D_cache/cache_reg[3][44]  ( .D(\D_cache/n1441 ), .CK(clk), .RN(n4183), .Q(\D_cache/cache[3][44] ) );
  DFFRX1 \D_cache/cache_reg[7][44]  ( .D(\D_cache/n1437 ), .CK(clk), .RN(n4183), .Q(\D_cache/cache[7][44] ) );
  DFFRX1 \D_cache/cache_reg[3][46]  ( .D(\D_cache/n1425 ), .CK(clk), .RN(n4184), .Q(\D_cache/cache[3][46] ) );
  DFFRX1 \D_cache/cache_reg[7][46]  ( .D(\D_cache/n1421 ), .CK(clk), .RN(n4185), .Q(\D_cache/cache[7][46] ) );
  DFFRX1 \D_cache/cache_reg[3][47]  ( .D(\D_cache/n1417 ), .CK(clk), .RN(n4185), .Q(\D_cache/cache[3][47] ) );
  DFFRX1 \D_cache/cache_reg[7][47]  ( .D(\D_cache/n1413 ), .CK(clk), .RN(n4185), .Q(\D_cache/cache[7][47] ) );
  DFFRX1 \D_cache/cache_reg[3][48]  ( .D(\D_cache/n1409 ), .CK(clk), .RN(n4186), .Q(\D_cache/cache[3][48] ) );
  DFFRX1 \D_cache/cache_reg[7][48]  ( .D(\D_cache/n1405 ), .CK(clk), .RN(n4186), .Q(\D_cache/cache[7][48] ) );
  DFFRX1 \D_cache/cache_reg[3][49]  ( .D(\D_cache/n1401 ), .CK(clk), .RN(n4186), .Q(\D_cache/cache[3][49] ) );
  DFFRX1 \D_cache/cache_reg[7][49]  ( .D(\D_cache/n1397 ), .CK(clk), .RN(n4187), .Q(\D_cache/cache[7][49] ) );
  DFFRX1 \D_cache/cache_reg[3][50]  ( .D(\D_cache/n1393 ), .CK(clk), .RN(n4187), .Q(\D_cache/cache[3][50] ) );
  DFFRX1 \D_cache/cache_reg[7][50]  ( .D(\D_cache/n1389 ), .CK(clk), .RN(n4187), .Q(\D_cache/cache[7][50] ) );
  DFFRX1 \D_cache/cache_reg[3][51]  ( .D(\D_cache/n1385 ), .CK(clk), .RN(n4188), .Q(\D_cache/cache[3][51] ) );
  DFFRX1 \D_cache/cache_reg[7][51]  ( .D(\D_cache/n1381 ), .CK(clk), .RN(n4188), .Q(\D_cache/cache[7][51] ) );
  DFFRX1 \D_cache/cache_reg[3][52]  ( .D(\D_cache/n1377 ), .CK(clk), .RN(n4188), .Q(\D_cache/cache[3][52] ) );
  DFFRX1 \D_cache/cache_reg[7][52]  ( .D(\D_cache/n1373 ), .CK(clk), .RN(n4189), .Q(\D_cache/cache[7][52] ) );
  DFFRX1 \D_cache/cache_reg[7][53]  ( .D(\D_cache/n1365 ), .CK(clk), .RN(n4189), .Q(\D_cache/cache[7][53] ) );
  DFFRX1 \D_cache/cache_reg[3][55]  ( .D(\D_cache/n1353 ), .CK(clk), .RN(n4190), .Q(\D_cache/cache[3][55] ) );
  DFFRX1 \D_cache/cache_reg[7][55]  ( .D(\D_cache/n1349 ), .CK(clk), .RN(n4191), .Q(\D_cache/cache[7][55] ) );
  DFFRX1 \D_cache/cache_reg[3][56]  ( .D(\D_cache/n1345 ), .CK(clk), .RN(n4191), .Q(\D_cache/cache[3][56] ) );
  DFFRX1 \D_cache/cache_reg[7][56]  ( .D(\D_cache/n1341 ), .CK(clk), .RN(n4191), .Q(\D_cache/cache[7][56] ) );
  DFFRX1 \D_cache/cache_reg[3][57]  ( .D(\D_cache/n1337 ), .CK(clk), .RN(n4192), .Q(\D_cache/cache[3][57] ) );
  DFFRX1 \D_cache/cache_reg[7][57]  ( .D(\D_cache/n1333 ), .CK(clk), .RN(n4192), .Q(\D_cache/cache[7][57] ) );
  DFFRX1 \D_cache/cache_reg[3][58]  ( .D(\D_cache/n1329 ), .CK(clk), .RN(n4192), .Q(\D_cache/cache[3][58] ) );
  DFFRX1 \D_cache/cache_reg[7][58]  ( .D(\D_cache/n1325 ), .CK(clk), .RN(n4193), .Q(\D_cache/cache[7][58] ) );
  DFFRX1 \D_cache/cache_reg[3][59]  ( .D(\D_cache/n1321 ), .CK(clk), .RN(n4193), .Q(\D_cache/cache[3][59] ) );
  DFFRX1 \D_cache/cache_reg[7][59]  ( .D(\D_cache/n1317 ), .CK(clk), .RN(n4193), .Q(\D_cache/cache[7][59] ) );
  DFFRX1 \D_cache/cache_reg[3][60]  ( .D(\D_cache/n1313 ), .CK(clk), .RN(n4194), .Q(\D_cache/cache[3][60] ) );
  DFFRX1 \D_cache/cache_reg[7][60]  ( .D(\D_cache/n1309 ), .CK(clk), .RN(n4194), .Q(\D_cache/cache[7][60] ) );
  DFFRX1 \D_cache/cache_reg[3][61]  ( .D(\D_cache/n1305 ), .CK(clk), .RN(n4194), .Q(\D_cache/cache[3][61] ) );
  DFFRX1 \D_cache/cache_reg[7][61]  ( .D(\D_cache/n1301 ), .CK(clk), .RN(n4195), .Q(\D_cache/cache[7][61] ) );
  DFFRX1 \D_cache/cache_reg[3][62]  ( .D(\D_cache/n1297 ), .CK(clk), .RN(n4195), .Q(\D_cache/cache[3][62] ) );
  DFFRX1 \D_cache/cache_reg[7][62]  ( .D(\D_cache/n1293 ), .CK(clk), .RN(n4195), .Q(\D_cache/cache[7][62] ) );
  DFFRX1 \D_cache/cache_reg[3][63]  ( .D(\D_cache/n1289 ), .CK(clk), .RN(n4196), .Q(\D_cache/cache[3][63] ) );
  DFFRX1 \D_cache/cache_reg[7][63]  ( .D(\D_cache/n1285 ), .CK(clk), .RN(n4196), .Q(\D_cache/cache[7][63] ) );
  DFFRX1 \D_cache/cache_reg[3][64]  ( .D(\D_cache/n1281 ), .CK(clk), .RN(n4196), .Q(\D_cache/cache[3][64] ) );
  DFFRX1 \D_cache/cache_reg[7][64]  ( .D(\D_cache/n1277 ), .CK(clk), .RN(n4197), .Q(\D_cache/cache[7][64] ) );
  DFFRX1 \D_cache/cache_reg[3][65]  ( .D(\D_cache/n1273 ), .CK(clk), .RN(n4197), .Q(\D_cache/cache[3][65] ) );
  DFFRX1 \D_cache/cache_reg[7][65]  ( .D(\D_cache/n1269 ), .CK(clk), .RN(n4197), .Q(\D_cache/cache[7][65] ) );
  DFFRX1 \D_cache/cache_reg[3][66]  ( .D(\D_cache/n1265 ), .CK(clk), .RN(n4198), .Q(\D_cache/cache[3][66] ) );
  DFFRX1 \D_cache/cache_reg[7][66]  ( .D(\D_cache/n1261 ), .CK(clk), .RN(n4198), .Q(\D_cache/cache[7][66] ) );
  DFFRX1 \D_cache/cache_reg[3][67]  ( .D(\D_cache/n1257 ), .CK(clk), .RN(n4198), .Q(\D_cache/cache[3][67] ) );
  DFFRX1 \D_cache/cache_reg[7][67]  ( .D(\D_cache/n1253 ), .CK(clk), .RN(n4199), .Q(\D_cache/cache[7][67] ) );
  DFFRX1 \D_cache/cache_reg[3][68]  ( .D(\D_cache/n1249 ), .CK(clk), .RN(n4199), .Q(\D_cache/cache[3][68] ) );
  DFFRX1 \D_cache/cache_reg[7][68]  ( .D(\D_cache/n1245 ), .CK(clk), .RN(n4199), .Q(\D_cache/cache[7][68] ) );
  DFFRX1 \D_cache/cache_reg[3][74]  ( .D(\D_cache/n1201 ), .CK(clk), .RN(n4203), .Q(\D_cache/cache[3][74] ) );
  DFFRX1 \D_cache/cache_reg[3][78]  ( .D(\D_cache/n1169 ), .CK(clk), .RN(n4206), .Q(\D_cache/cache[3][78] ) );
  DFFRX1 \D_cache/cache_reg[7][78]  ( .D(\D_cache/n1165 ), .CK(clk), .RN(n4206), .Q(\D_cache/cache[7][78] ) );
  DFFRX1 \D_cache/cache_reg[3][79]  ( .D(\D_cache/n1161 ), .CK(clk), .RN(n4206), .Q(\D_cache/cache[3][79] ) );
  DFFRX1 \D_cache/cache_reg[7][79]  ( .D(\D_cache/n1157 ), .CK(clk), .RN(n4207), .Q(\D_cache/cache[7][79] ) );
  DFFRX1 \D_cache/cache_reg[3][80]  ( .D(\D_cache/n1153 ), .CK(clk), .RN(n4207), .Q(\D_cache/cache[3][80] ) );
  DFFRX1 \D_cache/cache_reg[7][80]  ( .D(\D_cache/n1149 ), .CK(clk), .RN(n4207), .Q(\D_cache/cache[7][80] ) );
  DFFRX1 \D_cache/cache_reg[3][81]  ( .D(\D_cache/n1145 ), .CK(clk), .RN(n4208), .Q(\D_cache/cache[3][81] ) );
  DFFRX1 \D_cache/cache_reg[7][81]  ( .D(\D_cache/n1141 ), .CK(clk), .RN(n4208), .Q(\D_cache/cache[7][81] ) );
  DFFRX1 \D_cache/cache_reg[3][82]  ( .D(\D_cache/n1137 ), .CK(clk), .RN(n4208), .Q(\D_cache/cache[3][82] ) );
  DFFRX1 \D_cache/cache_reg[7][82]  ( .D(\D_cache/n1133 ), .CK(clk), .RN(n4209), .Q(\D_cache/cache[7][82] ) );
  DFFRX1 \D_cache/cache_reg[3][83]  ( .D(\D_cache/n1129 ), .CK(clk), .RN(n4209), .Q(\D_cache/cache[3][83] ) );
  DFFRX1 \D_cache/cache_reg[7][83]  ( .D(\D_cache/n1125 ), .CK(clk), .RN(n4209), .Q(\D_cache/cache[7][83] ) );
  DFFRX1 \D_cache/cache_reg[3][84]  ( .D(\D_cache/n1121 ), .CK(clk), .RN(n4210), .Q(\D_cache/cache[3][84] ) );
  DFFRX1 \D_cache/cache_reg[7][84]  ( .D(\D_cache/n1117 ), .CK(clk), .RN(n4210), .Q(\D_cache/cache[7][84] ) );
  DFFRX1 \D_cache/cache_reg[3][85]  ( .D(\D_cache/n1113 ), .CK(clk), .RN(n4210), .Q(\D_cache/cache[3][85] ) );
  DFFRX1 \D_cache/cache_reg[7][85]  ( .D(\D_cache/n1109 ), .CK(clk), .RN(n4211), .Q(\D_cache/cache[7][85] ) );
  DFFRX1 \D_cache/cache_reg[3][86]  ( .D(\D_cache/n1105 ), .CK(clk), .RN(n4211), .Q(\D_cache/cache[3][86] ) );
  DFFRX1 \D_cache/cache_reg[7][86]  ( .D(\D_cache/n1101 ), .CK(clk), .RN(n4211), .Q(\D_cache/cache[7][86] ) );
  DFFRX1 \D_cache/cache_reg[3][87]  ( .D(\D_cache/n1097 ), .CK(clk), .RN(n4212), .Q(\D_cache/cache[3][87] ) );
  DFFRX1 \D_cache/cache_reg[7][87]  ( .D(\D_cache/n1093 ), .CK(clk), .RN(n4212), .Q(\D_cache/cache[7][87] ) );
  DFFRX1 \D_cache/cache_reg[3][88]  ( .D(\D_cache/n1089 ), .CK(clk), .RN(n4212), .Q(\D_cache/cache[3][88] ) );
  DFFRX1 \D_cache/cache_reg[7][88]  ( .D(\D_cache/n1085 ), .CK(clk), .RN(n4213), .Q(\D_cache/cache[7][88] ) );
  DFFRX1 \D_cache/cache_reg[3][89]  ( .D(\D_cache/n1081 ), .CK(clk), .RN(n4213), .Q(\D_cache/cache[3][89] ) );
  DFFRX1 \D_cache/cache_reg[7][89]  ( .D(\D_cache/n1077 ), .CK(clk), .RN(n4213), .Q(\D_cache/cache[7][89] ) );
  DFFRX1 \D_cache/cache_reg[3][90]  ( .D(\D_cache/n1073 ), .CK(clk), .RN(n4214), .Q(\D_cache/cache[3][90] ) );
  DFFRX1 \D_cache/cache_reg[7][90]  ( .D(\D_cache/n1069 ), .CK(clk), .RN(n4214), .Q(\D_cache/cache[7][90] ) );
  DFFRX1 \D_cache/cache_reg[3][91]  ( .D(\D_cache/n1065 ), .CK(clk), .RN(n4214), .Q(\D_cache/cache[3][91] ) );
  DFFRX1 \D_cache/cache_reg[7][91]  ( .D(\D_cache/n1061 ), .CK(clk), .RN(n4215), .Q(\D_cache/cache[7][91] ) );
  DFFRX1 \D_cache/cache_reg[3][92]  ( .D(\D_cache/n1057 ), .CK(clk), .RN(n4215), .Q(\D_cache/cache[3][92] ) );
  DFFRX1 \D_cache/cache_reg[7][92]  ( .D(\D_cache/n1053 ), .CK(clk), .RN(n4215), .Q(\D_cache/cache[7][92] ) );
  DFFRX1 \D_cache/cache_reg[3][93]  ( .D(\D_cache/n1049 ), .CK(clk), .RN(n4216), .Q(\D_cache/cache[3][93] ) );
  DFFRX1 \D_cache/cache_reg[7][93]  ( .D(\D_cache/n1045 ), .CK(clk), .RN(n4216), .Q(\D_cache/cache[7][93] ) );
  DFFRX1 \D_cache/cache_reg[3][94]  ( .D(\D_cache/n1041 ), .CK(clk), .RN(n4216), .Q(\D_cache/cache[3][94] ) );
  DFFRX1 \D_cache/cache_reg[7][94]  ( .D(\D_cache/n1037 ), .CK(clk), .RN(n4217), .Q(\D_cache/cache[7][94] ) );
  DFFRX1 \D_cache/cache_reg[3][95]  ( .D(\D_cache/n1033 ), .CK(clk), .RN(n4217), .Q(\D_cache/cache[3][95] ) );
  DFFRX1 \D_cache/cache_reg[7][95]  ( .D(\D_cache/n1029 ), .CK(clk), .RN(n4217), .Q(\D_cache/cache[7][95] ) );
  DFFRX1 \D_cache/cache_reg[3][97]  ( .D(\D_cache/n1017 ), .CK(clk), .RN(n4218), .Q(\D_cache/cache[3][97] ) );
  DFFRX1 \D_cache/cache_reg[7][97]  ( .D(\D_cache/n1013 ), .CK(clk), .RN(n4219), .Q(\D_cache/cache[7][97] ) );
  DFFRX1 \D_cache/cache_reg[3][99]  ( .D(\D_cache/n1001 ), .CK(clk), .RN(n4220), .Q(\D_cache/cache[3][99] ) );
  DFFRX1 \D_cache/cache_reg[7][99]  ( .D(\D_cache/n997 ), .CK(clk), .RN(n4220), 
        .Q(\D_cache/cache[7][99] ) );
  DFFRX1 \D_cache/cache_reg[3][111]  ( .D(\D_cache/n905 ), .CK(clk), .RN(n4228), .Q(\D_cache/cache[3][111] ) );
  DFFRX1 \D_cache/cache_reg[7][111]  ( .D(\D_cache/n901 ), .CK(clk), .RN(n4228), .Q(\D_cache/cache[7][111] ) );
  DFFRX1 \D_cache/cache_reg[3][112]  ( .D(\D_cache/n897 ), .CK(clk), .RN(n4228), .Q(\D_cache/cache[3][112] ) );
  DFFRX1 \D_cache/cache_reg[7][112]  ( .D(\D_cache/n893 ), .CK(clk), .RN(n4229), .Q(\D_cache/cache[7][112] ) );
  DFFRX1 \D_cache/cache_reg[3][113]  ( .D(\D_cache/n889 ), .CK(clk), .RN(n4229), .Q(\D_cache/cache[3][113] ) );
  DFFRX1 \D_cache/cache_reg[7][113]  ( .D(\D_cache/n885 ), .CK(clk), .RN(n4229), .Q(\D_cache/cache[7][113] ) );
  DFFRX1 \D_cache/cache_reg[3][114]  ( .D(\D_cache/n881 ), .CK(clk), .RN(n4230), .Q(\D_cache/cache[3][114] ) );
  DFFRX1 \D_cache/cache_reg[7][114]  ( .D(\D_cache/n877 ), .CK(clk), .RN(n4230), .Q(\D_cache/cache[7][114] ) );
  DFFRX1 \D_cache/cache_reg[3][115]  ( .D(\D_cache/n873 ), .CK(clk), .RN(n4230), .Q(\D_cache/cache[3][115] ) );
  DFFRX1 \D_cache/cache_reg[7][115]  ( .D(\D_cache/n869 ), .CK(clk), .RN(n4231), .Q(\D_cache/cache[7][115] ) );
  DFFRX1 \D_cache/cache_reg[3][116]  ( .D(\D_cache/n865 ), .CK(clk), .RN(n4231), .Q(\D_cache/cache[3][116] ) );
  DFFRX1 \D_cache/cache_reg[7][116]  ( .D(\D_cache/n861 ), .CK(clk), .RN(n4231), .Q(\D_cache/cache[7][116] ) );
  DFFRX1 \D_cache/cache_reg[3][117]  ( .D(\D_cache/n857 ), .CK(clk), .RN(n4232), .Q(\D_cache/cache[3][117] ) );
  DFFRX1 \D_cache/cache_reg[7][117]  ( .D(\D_cache/n853 ), .CK(clk), .RN(n4232), .Q(\D_cache/cache[7][117] ) );
  DFFRX1 \D_cache/cache_reg[3][119]  ( .D(\D_cache/n841 ), .CK(clk), .RN(n4233), .Q(\D_cache/cache[3][119] ) );
  DFFRX1 \D_cache/cache_reg[7][119]  ( .D(\D_cache/n837 ), .CK(clk), .RN(n4233), .Q(\D_cache/cache[7][119] ) );
  DFFRX1 \D_cache/cache_reg[3][120]  ( .D(\D_cache/n833 ), .CK(clk), .RN(n4234), .Q(\D_cache/cache[3][120] ) );
  DFFRX1 \D_cache/cache_reg[7][120]  ( .D(\D_cache/n829 ), .CK(clk), .RN(n4234), .Q(\D_cache/cache[7][120] ) );
  DFFRX1 \D_cache/cache_reg[3][121]  ( .D(\D_cache/n825 ), .CK(clk), .RN(n4234), .Q(\D_cache/cache[3][121] ) );
  DFFRX1 \D_cache/cache_reg[7][121]  ( .D(\D_cache/n821 ), .CK(clk), .RN(n4235), .Q(\D_cache/cache[7][121] ) );
  DFFRX1 \D_cache/cache_reg[3][122]  ( .D(\D_cache/n817 ), .CK(clk), .RN(n4235), .Q(\D_cache/cache[3][122] ) );
  DFFRX1 \D_cache/cache_reg[7][122]  ( .D(\D_cache/n813 ), .CK(clk), .RN(n4235), .Q(\D_cache/cache[7][122] ) );
  DFFRX1 \D_cache/cache_reg[3][123]  ( .D(\D_cache/n809 ), .CK(clk), .RN(n4236), .Q(\D_cache/cache[3][123] ) );
  DFFRX1 \D_cache/cache_reg[7][123]  ( .D(\D_cache/n805 ), .CK(clk), .RN(n4236), .Q(\D_cache/cache[7][123] ) );
  DFFRX1 \D_cache/cache_reg[3][124]  ( .D(\D_cache/n801 ), .CK(clk), .RN(n4236), .Q(\D_cache/cache[3][124] ) );
  DFFRX1 \D_cache/cache_reg[7][124]  ( .D(\D_cache/n797 ), .CK(clk), .RN(n4237), .Q(\D_cache/cache[7][124] ) );
  DFFRX1 \D_cache/cache_reg[3][125]  ( .D(\D_cache/n793 ), .CK(clk), .RN(n4237), .Q(\D_cache/cache[3][125] ) );
  DFFRX1 \D_cache/cache_reg[7][125]  ( .D(\D_cache/n789 ), .CK(clk), .RN(n4237), .Q(\D_cache/cache[7][125] ) );
  DFFRX1 \D_cache/cache_reg[3][126]  ( .D(\D_cache/n785 ), .CK(clk), .RN(n4238), .Q(\D_cache/cache[3][126] ) );
  DFFRX1 \D_cache/cache_reg[7][126]  ( .D(\D_cache/n781 ), .CK(clk), .RN(n4238), .Q(\D_cache/cache[7][126] ) );
  DFFRX1 \D_cache/cache_reg[3][127]  ( .D(\D_cache/n777 ), .CK(clk), .RN(n4238), .Q(\D_cache/cache[3][127] ) );
  DFFRX1 \D_cache/cache_reg[7][127]  ( .D(\D_cache/n773 ), .CK(clk), .RN(n4239), .Q(\D_cache/cache[7][127] ) );
  DFFRX1 \D_cache/cache_reg[1][16]  ( .D(\D_cache/n1667 ), .CK(clk), .RN(n4164), .Q(\D_cache/cache[1][16] ) );
  DFFRX1 \D_cache/cache_reg[5][16]  ( .D(\D_cache/n1663 ), .CK(clk), .RN(n4165), .Q(\D_cache/cache[5][16] ) );
  DFFRX1 \D_cache/cache_reg[1][29]  ( .D(\D_cache/n1563 ), .CK(clk), .RN(n4173), .Q(\D_cache/cache[1][29] ) );
  DFFRX1 \D_cache/cache_reg[5][29]  ( .D(\D_cache/n1559 ), .CK(clk), .RN(n4173), .Q(\D_cache/cache[5][29] ) );
  DFFRX1 \D_cache/cache_reg[1][30]  ( .D(\D_cache/n1555 ), .CK(clk), .RN(n4174), .Q(\D_cache/cache[1][30] ) );
  DFFRX1 \D_cache/cache_reg[5][30]  ( .D(\D_cache/n1551 ), .CK(clk), .RN(n4174), .Q(\D_cache/cache[5][30] ) );
  DFFRX1 \D_cache/cache_reg[1][33]  ( .D(\D_cache/n1531 ), .CK(clk), .RN(n4176), .Q(\D_cache/cache[1][33] ) );
  DFFRX1 \D_cache/cache_reg[5][33]  ( .D(\D_cache/n1527 ), .CK(clk), .RN(n4176), .Q(\D_cache/cache[5][33] ) );
  DFFRX1 \D_cache/cache_reg[1][34]  ( .D(\D_cache/n1523 ), .CK(clk), .RN(n4176), .Q(\D_cache/cache[1][34] ) );
  DFFRX1 \D_cache/cache_reg[5][34]  ( .D(\D_cache/n1519 ), .CK(clk), .RN(n4177), .Q(\D_cache/cache[5][34] ) );
  DFFRX1 \D_cache/cache_reg[1][35]  ( .D(\D_cache/n1515 ), .CK(clk), .RN(n4177), .Q(\D_cache/cache[1][35] ) );
  DFFRX1 \D_cache/cache_reg[5][35]  ( .D(\D_cache/n1511 ), .CK(clk), .RN(n4177), .Q(\D_cache/cache[5][35] ) );
  DFFRX1 \D_cache/cache_reg[1][37]  ( .D(\D_cache/n1499 ), .CK(clk), .RN(n4178), .Q(\D_cache/cache[1][37] ) );
  DFFRX1 \D_cache/cache_reg[5][37]  ( .D(\D_cache/n1495 ), .CK(clk), .RN(n4179), .Q(\D_cache/cache[5][37] ) );
  DFFRX1 \D_cache/cache_reg[1][38]  ( .D(\D_cache/n1491 ), .CK(clk), .RN(n4179), .Q(\D_cache/cache[1][38] ) );
  DFFRX1 \D_cache/cache_reg[5][38]  ( .D(\D_cache/n1487 ), .CK(clk), .RN(n4179), .Q(\D_cache/cache[5][38] ) );
  DFFRX1 \D_cache/cache_reg[1][42]  ( .D(\D_cache/n1459 ), .CK(clk), .RN(n4182), .Q(\D_cache/cache[1][42] ) );
  DFFRX1 \D_cache/cache_reg[5][42]  ( .D(\D_cache/n1455 ), .CK(clk), .RN(n4182), .Q(\D_cache/cache[5][42] ) );
  DFFRX1 \D_cache/cache_reg[1][46]  ( .D(\D_cache/n1427 ), .CK(clk), .RN(n4184), .Q(\D_cache/cache[1][46] ) );
  DFFRX1 \D_cache/cache_reg[5][46]  ( .D(\D_cache/n1423 ), .CK(clk), .RN(n4185), .Q(\D_cache/cache[5][46] ) );
  DFFRX1 \D_cache/cache_reg[1][47]  ( .D(\D_cache/n1419 ), .CK(clk), .RN(n4185), .Q(\D_cache/cache[1][47] ) );
  DFFRX1 \D_cache/cache_reg[5][47]  ( .D(\D_cache/n1415 ), .CK(clk), .RN(n4185), .Q(\D_cache/cache[5][47] ) );
  DFFRX1 \D_cache/cache_reg[1][48]  ( .D(\D_cache/n1411 ), .CK(clk), .RN(n4186), .Q(\D_cache/cache[1][48] ) );
  DFFRX1 \D_cache/cache_reg[5][48]  ( .D(\D_cache/n1407 ), .CK(clk), .RN(n4186), .Q(\D_cache/cache[5][48] ) );
  DFFRX1 \D_cache/cache_reg[1][49]  ( .D(\D_cache/n1403 ), .CK(clk), .RN(n4186), .Q(\D_cache/cache[1][49] ) );
  DFFRX1 \D_cache/cache_reg[5][49]  ( .D(\D_cache/n1399 ), .CK(clk), .RN(n4187), .Q(\D_cache/cache[5][49] ) );
  DFFRX1 \D_cache/cache_reg[1][50]  ( .D(\D_cache/n1395 ), .CK(clk), .RN(n4187), .Q(\D_cache/cache[1][50] ) );
  DFFRX1 \D_cache/cache_reg[5][50]  ( .D(\D_cache/n1391 ), .CK(clk), .RN(n4187), .Q(\D_cache/cache[5][50] ) );
  DFFRX1 \D_cache/cache_reg[1][51]  ( .D(\D_cache/n1387 ), .CK(clk), .RN(n4188), .Q(\D_cache/cache[1][51] ) );
  DFFRX1 \D_cache/cache_reg[5][51]  ( .D(\D_cache/n1383 ), .CK(clk), .RN(n4188), .Q(\D_cache/cache[5][51] ) );
  DFFRX1 \D_cache/cache_reg[1][52]  ( .D(\D_cache/n1379 ), .CK(clk), .RN(n4188), .Q(\D_cache/cache[1][52] ) );
  DFFRX1 \D_cache/cache_reg[5][52]  ( .D(\D_cache/n1375 ), .CK(clk), .RN(n4189), .Q(\D_cache/cache[5][52] ) );
  DFFRX1 \D_cache/cache_reg[1][55]  ( .D(\D_cache/n1355 ), .CK(clk), .RN(n4190), .Q(\D_cache/cache[1][55] ) );
  DFFRX1 \D_cache/cache_reg[5][55]  ( .D(\D_cache/n1351 ), .CK(clk), .RN(n4191), .Q(\D_cache/cache[5][55] ) );
  DFFRX1 \D_cache/cache_reg[1][56]  ( .D(\D_cache/n1347 ), .CK(clk), .RN(n4191), .Q(\D_cache/cache[1][56] ) );
  DFFRX1 \D_cache/cache_reg[5][56]  ( .D(\D_cache/n1343 ), .CK(clk), .RN(n4191), .Q(\D_cache/cache[5][56] ) );
  DFFRX1 \D_cache/cache_reg[1][57]  ( .D(\D_cache/n1339 ), .CK(clk), .RN(n4192), .Q(\D_cache/cache[1][57] ) );
  DFFRX1 \D_cache/cache_reg[5][57]  ( .D(\D_cache/n1335 ), .CK(clk), .RN(n4192), .Q(\D_cache/cache[5][57] ) );
  DFFRX1 \D_cache/cache_reg[1][58]  ( .D(\D_cache/n1331 ), .CK(clk), .RN(n4192), .Q(\D_cache/cache[1][58] ) );
  DFFRX1 \D_cache/cache_reg[5][58]  ( .D(\D_cache/n1327 ), .CK(clk), .RN(n4193), .Q(\D_cache/cache[5][58] ) );
  DFFRX1 \D_cache/cache_reg[1][59]  ( .D(\D_cache/n1323 ), .CK(clk), .RN(n4193), .Q(\D_cache/cache[1][59] ) );
  DFFRX1 \D_cache/cache_reg[5][59]  ( .D(\D_cache/n1319 ), .CK(clk), .RN(n4193), .Q(\D_cache/cache[5][59] ) );
  DFFRX1 \D_cache/cache_reg[1][61]  ( .D(\D_cache/n1307 ), .CK(clk), .RN(n4194), .Q(\D_cache/cache[1][61] ) );
  DFFRX1 \D_cache/cache_reg[5][61]  ( .D(\D_cache/n1303 ), .CK(clk), .RN(n4195), .Q(\D_cache/cache[5][61] ) );
  DFFRX1 \D_cache/cache_reg[1][62]  ( .D(\D_cache/n1299 ), .CK(clk), .RN(n4195), .Q(\D_cache/cache[1][62] ) );
  DFFRX1 \D_cache/cache_reg[5][62]  ( .D(\D_cache/n1295 ), .CK(clk), .RN(n4195), .Q(\D_cache/cache[5][62] ) );
  DFFRX1 \D_cache/cache_reg[1][63]  ( .D(\D_cache/n1291 ), .CK(clk), .RN(n4196), .Q(\D_cache/cache[1][63] ) );
  DFFRX1 \D_cache/cache_reg[5][63]  ( .D(\D_cache/n1287 ), .CK(clk), .RN(n4196), .Q(\D_cache/cache[5][63] ) );
  DFFRX1 \D_cache/cache_reg[1][64]  ( .D(\D_cache/n1283 ), .CK(clk), .RN(n4196), .Q(\D_cache/cache[1][64] ) );
  DFFRX1 \D_cache/cache_reg[1][65]  ( .D(\D_cache/n1275 ), .CK(clk), .RN(n4197), .Q(\D_cache/cache[1][65] ) );
  DFFRX1 \D_cache/cache_reg[5][65]  ( .D(\D_cache/n1271 ), .CK(clk), .RN(n4197), .Q(\D_cache/cache[5][65] ) );
  DFFRX1 \D_cache/cache_reg[1][66]  ( .D(\D_cache/n1267 ), .CK(clk), .RN(n4198), .Q(\D_cache/cache[1][66] ) );
  DFFRX1 \D_cache/cache_reg[1][67]  ( .D(\D_cache/n1259 ), .CK(clk), .RN(n4198), .Q(\D_cache/cache[1][67] ) );
  DFFRX1 \D_cache/cache_reg[5][67]  ( .D(\D_cache/n1255 ), .CK(clk), .RN(n4199), .Q(\D_cache/cache[5][67] ) );
  DFFRX1 \D_cache/cache_reg[1][68]  ( .D(\D_cache/n1251 ), .CK(clk), .RN(n4199), .Q(\D_cache/cache[1][68] ) );
  DFFRX1 \D_cache/cache_reg[5][68]  ( .D(\D_cache/n1247 ), .CK(clk), .RN(n4199), .Q(\D_cache/cache[5][68] ) );
  DFFRX1 \D_cache/cache_reg[1][78]  ( .D(\D_cache/n1171 ), .CK(clk), .RN(n4206), .Q(\D_cache/cache[1][78] ) );
  DFFRX1 \D_cache/cache_reg[5][78]  ( .D(\D_cache/n1167 ), .CK(clk), .RN(n4206), .Q(\D_cache/cache[5][78] ) );
  DFFRX1 \D_cache/cache_reg[1][79]  ( .D(\D_cache/n1163 ), .CK(clk), .RN(n4206), .Q(\D_cache/cache[1][79] ) );
  DFFRX1 \D_cache/cache_reg[5][79]  ( .D(\D_cache/n1159 ), .CK(clk), .RN(n4207), .Q(\D_cache/cache[5][79] ) );
  DFFRX1 \D_cache/cache_reg[1][80]  ( .D(\D_cache/n1155 ), .CK(clk), .RN(n4207), .Q(\D_cache/cache[1][80] ) );
  DFFRX1 \D_cache/cache_reg[5][80]  ( .D(\D_cache/n1151 ), .CK(clk), .RN(n4207), .Q(\D_cache/cache[5][80] ) );
  DFFRX1 \D_cache/cache_reg[1][81]  ( .D(\D_cache/n1147 ), .CK(clk), .RN(n4208), .Q(\D_cache/cache[1][81] ) );
  DFFRX1 \D_cache/cache_reg[5][81]  ( .D(\D_cache/n1143 ), .CK(clk), .RN(n4208), .Q(\D_cache/cache[5][81] ) );
  DFFRX1 \D_cache/cache_reg[1][82]  ( .D(\D_cache/n1139 ), .CK(clk), .RN(n4208), .Q(\D_cache/cache[1][82] ) );
  DFFRX1 \D_cache/cache_reg[5][82]  ( .D(\D_cache/n1135 ), .CK(clk), .RN(n4209), .Q(\D_cache/cache[5][82] ) );
  DFFRX1 \D_cache/cache_reg[1][83]  ( .D(\D_cache/n1131 ), .CK(clk), .RN(n4209), .Q(\D_cache/cache[1][83] ) );
  DFFRX1 \D_cache/cache_reg[5][83]  ( .D(\D_cache/n1127 ), .CK(clk), .RN(n4209), .Q(\D_cache/cache[5][83] ) );
  DFFRX1 \D_cache/cache_reg[1][84]  ( .D(\D_cache/n1123 ), .CK(clk), .RN(n4210), .Q(\D_cache/cache[1][84] ) );
  DFFRX1 \D_cache/cache_reg[5][84]  ( .D(\D_cache/n1119 ), .CK(clk), .RN(n4210), .Q(\D_cache/cache[5][84] ) );
  DFFRX1 \D_cache/cache_reg[1][85]  ( .D(\D_cache/n1115 ), .CK(clk), .RN(n4210), .Q(\D_cache/cache[1][85] ) );
  DFFRX1 \D_cache/cache_reg[5][85]  ( .D(\D_cache/n1111 ), .CK(clk), .RN(n4211), .Q(\D_cache/cache[5][85] ) );
  DFFRX1 \D_cache/cache_reg[1][86]  ( .D(\D_cache/n1107 ), .CK(clk), .RN(n4211), .Q(\D_cache/cache[1][86] ) );
  DFFRX1 \D_cache/cache_reg[5][86]  ( .D(\D_cache/n1103 ), .CK(clk), .RN(n4211), .Q(\D_cache/cache[5][86] ) );
  DFFRX1 \D_cache/cache_reg[1][87]  ( .D(\D_cache/n1099 ), .CK(clk), .RN(n4212), .Q(\D_cache/cache[1][87] ) );
  DFFRX1 \D_cache/cache_reg[5][87]  ( .D(\D_cache/n1095 ), .CK(clk), .RN(n4212), .Q(\D_cache/cache[5][87] ) );
  DFFRX1 \D_cache/cache_reg[1][88]  ( .D(\D_cache/n1091 ), .CK(clk), .RN(n4212), .Q(\D_cache/cache[1][88] ) );
  DFFRX1 \D_cache/cache_reg[5][88]  ( .D(\D_cache/n1087 ), .CK(clk), .RN(n4213), .Q(\D_cache/cache[5][88] ) );
  DFFRX1 \D_cache/cache_reg[1][89]  ( .D(\D_cache/n1083 ), .CK(clk), .RN(n4213), .Q(\D_cache/cache[1][89] ) );
  DFFRX1 \D_cache/cache_reg[5][89]  ( .D(\D_cache/n1079 ), .CK(clk), .RN(n4213), .Q(\D_cache/cache[5][89] ) );
  DFFRX1 \D_cache/cache_reg[1][90]  ( .D(\D_cache/n1075 ), .CK(clk), .RN(n4214), .Q(\D_cache/cache[1][90] ) );
  DFFRX1 \D_cache/cache_reg[5][90]  ( .D(\D_cache/n1071 ), .CK(clk), .RN(n4214), .Q(\D_cache/cache[5][90] ) );
  DFFRX1 \D_cache/cache_reg[1][91]  ( .D(\D_cache/n1067 ), .CK(clk), .RN(n4214), .Q(\D_cache/cache[1][91] ) );
  DFFRX1 \D_cache/cache_reg[5][91]  ( .D(\D_cache/n1063 ), .CK(clk), .RN(n4215), .Q(\D_cache/cache[5][91] ) );
  DFFRX1 \D_cache/cache_reg[1][92]  ( .D(\D_cache/n1059 ), .CK(clk), .RN(n4215), .Q(\D_cache/cache[1][92] ) );
  DFFRX1 \D_cache/cache_reg[5][92]  ( .D(\D_cache/n1055 ), .CK(clk), .RN(n4215), .Q(\D_cache/cache[5][92] ) );
  DFFRX1 \D_cache/cache_reg[1][93]  ( .D(\D_cache/n1051 ), .CK(clk), .RN(n4216), .Q(\D_cache/cache[1][93] ) );
  DFFRX1 \D_cache/cache_reg[5][93]  ( .D(\D_cache/n1047 ), .CK(clk), .RN(n4216), .Q(\D_cache/cache[5][93] ) );
  DFFRX1 \D_cache/cache_reg[1][94]  ( .D(\D_cache/n1043 ), .CK(clk), .RN(n4216), .Q(\D_cache/cache[1][94] ) );
  DFFRX1 \D_cache/cache_reg[5][94]  ( .D(\D_cache/n1039 ), .CK(clk), .RN(n4217), .Q(\D_cache/cache[5][94] ) );
  DFFRX1 \D_cache/cache_reg[1][95]  ( .D(\D_cache/n1035 ), .CK(clk), .RN(n4217), .Q(\D_cache/cache[1][95] ) );
  DFFRX1 \D_cache/cache_reg[5][95]  ( .D(\D_cache/n1031 ), .CK(clk), .RN(n4217), .Q(\D_cache/cache[5][95] ) );
  DFFRX1 \D_cache/cache_reg[1][97]  ( .D(\D_cache/n1019 ), .CK(clk), .RN(n4218), .Q(\D_cache/cache[1][97] ) );
  DFFRX1 \D_cache/cache_reg[5][97]  ( .D(\D_cache/n1015 ), .CK(clk), .RN(n4219), .Q(\D_cache/cache[5][97] ) );
  DFFRX1 \D_cache/cache_reg[1][111]  ( .D(\D_cache/n907 ), .CK(clk), .RN(n4228), .Q(\D_cache/cache[1][111] ) );
  DFFRX1 \D_cache/cache_reg[5][111]  ( .D(\D_cache/n903 ), .CK(clk), .RN(n4228), .Q(\D_cache/cache[5][111] ) );
  DFFRX1 \D_cache/cache_reg[1][112]  ( .D(\D_cache/n899 ), .CK(clk), .RN(n4228), .Q(\D_cache/cache[1][112] ) );
  DFFRX1 \D_cache/cache_reg[5][112]  ( .D(\D_cache/n895 ), .CK(clk), .RN(n4229), .Q(\D_cache/cache[5][112] ) );
  DFFRX1 \D_cache/cache_reg[1][113]  ( .D(\D_cache/n891 ), .CK(clk), .RN(n4229), .Q(\D_cache/cache[1][113] ) );
  DFFRX1 \D_cache/cache_reg[5][113]  ( .D(\D_cache/n887 ), .CK(clk), .RN(n4229), .Q(\D_cache/cache[5][113] ) );
  DFFRX1 \D_cache/cache_reg[1][114]  ( .D(\D_cache/n883 ), .CK(clk), .RN(n4230), .Q(\D_cache/cache[1][114] ) );
  DFFRX1 \D_cache/cache_reg[5][114]  ( .D(\D_cache/n879 ), .CK(clk), .RN(n4230), .Q(\D_cache/cache[5][114] ) );
  DFFRX1 \D_cache/cache_reg[1][115]  ( .D(\D_cache/n875 ), .CK(clk), .RN(n4230), .Q(\D_cache/cache[1][115] ) );
  DFFRX1 \D_cache/cache_reg[5][115]  ( .D(\D_cache/n871 ), .CK(clk), .RN(n4231), .Q(\D_cache/cache[5][115] ) );
  DFFRX1 \D_cache/cache_reg[1][116]  ( .D(\D_cache/n867 ), .CK(clk), .RN(n4231), .Q(\D_cache/cache[1][116] ) );
  DFFRX1 \D_cache/cache_reg[5][116]  ( .D(\D_cache/n863 ), .CK(clk), .RN(n4231), .Q(\D_cache/cache[5][116] ) );
  DFFRX1 \D_cache/cache_reg[1][117]  ( .D(\D_cache/n859 ), .CK(clk), .RN(n4232), .Q(\D_cache/cache[1][117] ) );
  DFFRX1 \D_cache/cache_reg[5][117]  ( .D(\D_cache/n855 ), .CK(clk), .RN(n4232), .Q(\D_cache/cache[5][117] ) );
  DFFRX1 \D_cache/cache_reg[1][119]  ( .D(\D_cache/n843 ), .CK(clk), .RN(n4233), .Q(\D_cache/cache[1][119] ) );
  DFFRX1 \D_cache/cache_reg[5][119]  ( .D(\D_cache/n839 ), .CK(clk), .RN(n4233), .Q(\D_cache/cache[5][119] ) );
  DFFRX1 \D_cache/cache_reg[1][120]  ( .D(\D_cache/n835 ), .CK(clk), .RN(n4234), .Q(\D_cache/cache[1][120] ) );
  DFFRX1 \D_cache/cache_reg[5][120]  ( .D(\D_cache/n831 ), .CK(clk), .RN(n4234), .Q(\D_cache/cache[5][120] ) );
  DFFRX1 \D_cache/cache_reg[1][121]  ( .D(\D_cache/n827 ), .CK(clk), .RN(n4234), .Q(\D_cache/cache[1][121] ) );
  DFFRX1 \D_cache/cache_reg[5][121]  ( .D(\D_cache/n823 ), .CK(clk), .RN(n4235), .Q(\D_cache/cache[5][121] ) );
  DFFRX1 \D_cache/cache_reg[1][122]  ( .D(\D_cache/n819 ), .CK(clk), .RN(n4235), .Q(\D_cache/cache[1][122] ) );
  DFFRX1 \D_cache/cache_reg[5][122]  ( .D(\D_cache/n815 ), .CK(clk), .RN(n4235), .Q(\D_cache/cache[5][122] ) );
  DFFRX1 \D_cache/cache_reg[1][123]  ( .D(\D_cache/n811 ), .CK(clk), .RN(n4236), .Q(\D_cache/cache[1][123] ) );
  DFFRX1 \D_cache/cache_reg[5][123]  ( .D(\D_cache/n807 ), .CK(clk), .RN(n4236), .Q(\D_cache/cache[5][123] ) );
  DFFRX1 \D_cache/cache_reg[1][124]  ( .D(\D_cache/n803 ), .CK(clk), .RN(n4236), .Q(\D_cache/cache[1][124] ) );
  DFFRX1 \D_cache/cache_reg[5][124]  ( .D(\D_cache/n799 ), .CK(clk), .RN(n4237), .Q(\D_cache/cache[5][124] ) );
  DFFRX1 \D_cache/cache_reg[1][125]  ( .D(\D_cache/n795 ), .CK(clk), .RN(n4237), .Q(\D_cache/cache[1][125] ) );
  DFFRX1 \D_cache/cache_reg[5][125]  ( .D(\D_cache/n791 ), .CK(clk), .RN(n4237), .Q(\D_cache/cache[5][125] ) );
  DFFRX1 \D_cache/cache_reg[1][126]  ( .D(\D_cache/n787 ), .CK(clk), .RN(n4238), .Q(\D_cache/cache[1][126] ) );
  DFFRX1 \D_cache/cache_reg[5][126]  ( .D(\D_cache/n783 ), .CK(clk), .RN(n4238), .Q(\D_cache/cache[5][126] ) );
  DFFRX1 \D_cache/cache_reg[1][127]  ( .D(\D_cache/n779 ), .CK(clk), .RN(n4238), .Q(\D_cache/cache[1][127] ) );
  DFFRX1 \D_cache/cache_reg[5][127]  ( .D(\D_cache/n775 ), .CK(clk), .RN(n4239), .Q(\D_cache/cache[5][127] ) );
  DFFRX1 \D_cache/cache_reg[0][16]  ( .D(\D_cache/n1668 ), .CK(clk), .RN(n4164), .Q(\D_cache/cache[0][16] ) );
  DFFRX1 \D_cache/cache_reg[4][16]  ( .D(\D_cache/n1664 ), .CK(clk), .RN(n4165), .Q(\D_cache/cache[4][16] ) );
  DFFRX1 \D_cache/cache_reg[0][29]  ( .D(\D_cache/n1564 ), .CK(clk), .RN(n4173), .Q(\D_cache/cache[0][29] ) );
  DFFRX1 \D_cache/cache_reg[4][29]  ( .D(\D_cache/n1560 ), .CK(clk), .RN(n4173), .Q(\D_cache/cache[4][29] ) );
  DFFRX1 \D_cache/cache_reg[0][30]  ( .D(\D_cache/n1556 ), .CK(clk), .RN(n4174), .Q(\D_cache/cache[0][30] ) );
  DFFRX1 \D_cache/cache_reg[4][30]  ( .D(\D_cache/n1552 ), .CK(clk), .RN(n4174), .Q(\D_cache/cache[4][30] ) );
  DFFRX1 \D_cache/cache_reg[0][33]  ( .D(\D_cache/n1532 ), .CK(clk), .RN(n4176), .Q(\D_cache/cache[0][33] ) );
  DFFRX1 \D_cache/cache_reg[4][33]  ( .D(\D_cache/n1528 ), .CK(clk), .RN(n4176), .Q(\D_cache/cache[4][33] ) );
  DFFRX1 \D_cache/cache_reg[0][34]  ( .D(\D_cache/n1524 ), .CK(clk), .RN(n4176), .Q(\D_cache/cache[0][34] ) );
  DFFRX1 \D_cache/cache_reg[4][34]  ( .D(\D_cache/n1520 ), .CK(clk), .RN(n4177), .Q(\D_cache/cache[4][34] ) );
  DFFRX1 \D_cache/cache_reg[0][35]  ( .D(\D_cache/n1516 ), .CK(clk), .RN(n4177), .Q(\D_cache/cache[0][35] ) );
  DFFRX1 \D_cache/cache_reg[4][35]  ( .D(\D_cache/n1512 ), .CK(clk), .RN(n4177), .Q(\D_cache/cache[4][35] ) );
  DFFRX1 \D_cache/cache_reg[0][37]  ( .D(\D_cache/n1500 ), .CK(clk), .RN(n4178), .Q(\D_cache/cache[0][37] ) );
  DFFRX1 \D_cache/cache_reg[4][37]  ( .D(\D_cache/n1496 ), .CK(clk), .RN(n4179), .Q(\D_cache/cache[4][37] ) );
  DFFRX1 \D_cache/cache_reg[0][38]  ( .D(\D_cache/n1492 ), .CK(clk), .RN(n4179), .Q(\D_cache/cache[0][38] ) );
  DFFRX1 \D_cache/cache_reg[4][38]  ( .D(\D_cache/n1488 ), .CK(clk), .RN(n4179), .Q(\D_cache/cache[4][38] ) );
  DFFRX1 \D_cache/cache_reg[0][42]  ( .D(\D_cache/n1460 ), .CK(clk), .RN(n4182), .Q(\D_cache/cache[0][42] ) );
  DFFRX1 \D_cache/cache_reg[4][42]  ( .D(\D_cache/n1456 ), .CK(clk), .RN(n4182), .Q(\D_cache/cache[4][42] ) );
  DFFRX1 \D_cache/cache_reg[0][46]  ( .D(\D_cache/n1428 ), .CK(clk), .RN(n4184), .Q(\D_cache/cache[0][46] ) );
  DFFRX1 \D_cache/cache_reg[4][46]  ( .D(\D_cache/n1424 ), .CK(clk), .RN(n4185), .Q(\D_cache/cache[4][46] ) );
  DFFRX1 \D_cache/cache_reg[0][47]  ( .D(\D_cache/n1420 ), .CK(clk), .RN(n4185), .Q(\D_cache/cache[0][47] ) );
  DFFRX1 \D_cache/cache_reg[4][47]  ( .D(\D_cache/n1416 ), .CK(clk), .RN(n4185), .Q(\D_cache/cache[4][47] ) );
  DFFRX1 \D_cache/cache_reg[0][48]  ( .D(\D_cache/n1412 ), .CK(clk), .RN(n4186), .Q(\D_cache/cache[0][48] ) );
  DFFRX1 \D_cache/cache_reg[4][48]  ( .D(\D_cache/n1408 ), .CK(clk), .RN(n4186), .Q(\D_cache/cache[4][48] ) );
  DFFRX1 \D_cache/cache_reg[0][49]  ( .D(\D_cache/n1404 ), .CK(clk), .RN(n4186), .Q(\D_cache/cache[0][49] ) );
  DFFRX1 \D_cache/cache_reg[4][49]  ( .D(\D_cache/n1400 ), .CK(clk), .RN(n4187), .Q(\D_cache/cache[4][49] ) );
  DFFRX1 \D_cache/cache_reg[0][50]  ( .D(\D_cache/n1396 ), .CK(clk), .RN(n4187), .Q(\D_cache/cache[0][50] ) );
  DFFRX1 \D_cache/cache_reg[4][50]  ( .D(\D_cache/n1392 ), .CK(clk), .RN(n4187), .Q(\D_cache/cache[4][50] ) );
  DFFRX1 \D_cache/cache_reg[0][51]  ( .D(\D_cache/n1388 ), .CK(clk), .RN(n4188), .Q(\D_cache/cache[0][51] ) );
  DFFRX1 \D_cache/cache_reg[4][51]  ( .D(\D_cache/n1384 ), .CK(clk), .RN(n4188), .Q(\D_cache/cache[4][51] ) );
  DFFRX1 \D_cache/cache_reg[0][52]  ( .D(\D_cache/n1380 ), .CK(clk), .RN(n4188), .Q(\D_cache/cache[0][52] ) );
  DFFRX1 \D_cache/cache_reg[4][52]  ( .D(\D_cache/n1376 ), .CK(clk), .RN(n4189), .Q(\D_cache/cache[4][52] ) );
  DFFRX1 \D_cache/cache_reg[0][55]  ( .D(\D_cache/n1356 ), .CK(clk), .RN(n4190), .Q(\D_cache/cache[0][55] ) );
  DFFRX1 \D_cache/cache_reg[4][55]  ( .D(\D_cache/n1352 ), .CK(clk), .RN(n4191), .Q(\D_cache/cache[4][55] ) );
  DFFRX1 \D_cache/cache_reg[0][56]  ( .D(\D_cache/n1348 ), .CK(clk), .RN(n4191), .Q(\D_cache/cache[0][56] ) );
  DFFRX1 \D_cache/cache_reg[4][56]  ( .D(\D_cache/n1344 ), .CK(clk), .RN(n4191), .Q(\D_cache/cache[4][56] ) );
  DFFRX1 \D_cache/cache_reg[0][57]  ( .D(\D_cache/n1340 ), .CK(clk), .RN(n4192), .Q(\D_cache/cache[0][57] ) );
  DFFRX1 \D_cache/cache_reg[4][57]  ( .D(\D_cache/n1336 ), .CK(clk), .RN(n4192), .Q(\D_cache/cache[4][57] ) );
  DFFRX1 \D_cache/cache_reg[0][58]  ( .D(\D_cache/n1332 ), .CK(clk), .RN(n4192), .Q(\D_cache/cache[0][58] ) );
  DFFRX1 \D_cache/cache_reg[4][58]  ( .D(\D_cache/n1328 ), .CK(clk), .RN(n4193), .Q(\D_cache/cache[4][58] ) );
  DFFRX1 \D_cache/cache_reg[0][59]  ( .D(\D_cache/n1324 ), .CK(clk), .RN(n4193), .Q(\D_cache/cache[0][59] ) );
  DFFRX1 \D_cache/cache_reg[4][59]  ( .D(\D_cache/n1320 ), .CK(clk), .RN(n4193), .Q(\D_cache/cache[4][59] ) );
  DFFRX1 \D_cache/cache_reg[0][61]  ( .D(\D_cache/n1308 ), .CK(clk), .RN(n4194), .Q(\D_cache/cache[0][61] ) );
  DFFRX1 \D_cache/cache_reg[4][61]  ( .D(\D_cache/n1304 ), .CK(clk), .RN(n4195), .Q(\D_cache/cache[4][61] ) );
  DFFRX1 \D_cache/cache_reg[0][62]  ( .D(\D_cache/n1300 ), .CK(clk), .RN(n4195), .Q(\D_cache/cache[0][62] ) );
  DFFRX1 \D_cache/cache_reg[4][62]  ( .D(\D_cache/n1296 ), .CK(clk), .RN(n4195), .Q(\D_cache/cache[4][62] ) );
  DFFRX1 \D_cache/cache_reg[0][63]  ( .D(\D_cache/n1292 ), .CK(clk), .RN(n4196), .Q(\D_cache/cache[0][63] ) );
  DFFRX1 \D_cache/cache_reg[4][63]  ( .D(\D_cache/n1288 ), .CK(clk), .RN(n4196), .Q(\D_cache/cache[4][63] ) );
  DFFRX1 \D_cache/cache_reg[0][64]  ( .D(\D_cache/n1284 ), .CK(clk), .RN(n4196), .Q(\D_cache/cache[0][64] ) );
  DFFRX1 \D_cache/cache_reg[0][65]  ( .D(\D_cache/n1276 ), .CK(clk), .RN(n4197), .Q(\D_cache/cache[0][65] ) );
  DFFRX1 \D_cache/cache_reg[4][65]  ( .D(\D_cache/n1272 ), .CK(clk), .RN(n4197), .Q(\D_cache/cache[4][65] ) );
  DFFRX1 \D_cache/cache_reg[0][67]  ( .D(\D_cache/n1260 ), .CK(clk), .RN(n4198), .Q(\D_cache/cache[0][67] ) );
  DFFRX1 \D_cache/cache_reg[4][67]  ( .D(\D_cache/n1256 ), .CK(clk), .RN(n4199), .Q(\D_cache/cache[4][67] ) );
  DFFRX1 \D_cache/cache_reg[0][68]  ( .D(\D_cache/n1252 ), .CK(clk), .RN(n4199), .Q(\D_cache/cache[0][68] ) );
  DFFRX1 \D_cache/cache_reg[4][68]  ( .D(\D_cache/n1248 ), .CK(clk), .RN(n4199), .Q(\D_cache/cache[4][68] ) );
  DFFRX1 \D_cache/cache_reg[0][78]  ( .D(\D_cache/n1172 ), .CK(clk), .RN(n4206), .Q(\D_cache/cache[0][78] ) );
  DFFRX1 \D_cache/cache_reg[4][78]  ( .D(\D_cache/n1168 ), .CK(clk), .RN(n4206), .Q(\D_cache/cache[4][78] ) );
  DFFRX1 \D_cache/cache_reg[0][79]  ( .D(\D_cache/n1164 ), .CK(clk), .RN(n4206), .Q(\D_cache/cache[0][79] ) );
  DFFRX1 \D_cache/cache_reg[4][79]  ( .D(\D_cache/n1160 ), .CK(clk), .RN(n4207), .Q(\D_cache/cache[4][79] ) );
  DFFRX1 \D_cache/cache_reg[0][80]  ( .D(\D_cache/n1156 ), .CK(clk), .RN(n4207), .Q(\D_cache/cache[0][80] ) );
  DFFRX1 \D_cache/cache_reg[4][80]  ( .D(\D_cache/n1152 ), .CK(clk), .RN(n4207), .Q(\D_cache/cache[4][80] ) );
  DFFRX1 \D_cache/cache_reg[0][81]  ( .D(\D_cache/n1148 ), .CK(clk), .RN(n4208), .Q(\D_cache/cache[0][81] ) );
  DFFRX1 \D_cache/cache_reg[4][81]  ( .D(\D_cache/n1144 ), .CK(clk), .RN(n4208), .Q(\D_cache/cache[4][81] ) );
  DFFRX1 \D_cache/cache_reg[0][82]  ( .D(\D_cache/n1140 ), .CK(clk), .RN(n4208), .Q(\D_cache/cache[0][82] ) );
  DFFRX1 \D_cache/cache_reg[4][82]  ( .D(\D_cache/n1136 ), .CK(clk), .RN(n4209), .Q(\D_cache/cache[4][82] ) );
  DFFRX1 \D_cache/cache_reg[0][83]  ( .D(\D_cache/n1132 ), .CK(clk), .RN(n4209), .Q(\D_cache/cache[0][83] ) );
  DFFRX1 \D_cache/cache_reg[4][83]  ( .D(\D_cache/n1128 ), .CK(clk), .RN(n4209), .Q(\D_cache/cache[4][83] ) );
  DFFRX1 \D_cache/cache_reg[0][84]  ( .D(\D_cache/n1124 ), .CK(clk), .RN(n4210), .Q(\D_cache/cache[0][84] ) );
  DFFRX1 \D_cache/cache_reg[4][84]  ( .D(\D_cache/n1120 ), .CK(clk), .RN(n4210), .Q(\D_cache/cache[4][84] ) );
  DFFRX1 \D_cache/cache_reg[0][85]  ( .D(\D_cache/n1116 ), .CK(clk), .RN(n4210), .Q(\D_cache/cache[0][85] ) );
  DFFRX1 \D_cache/cache_reg[4][85]  ( .D(\D_cache/n1112 ), .CK(clk), .RN(n4211), .Q(\D_cache/cache[4][85] ) );
  DFFRX1 \D_cache/cache_reg[0][86]  ( .D(\D_cache/n1108 ), .CK(clk), .RN(n4211), .Q(\D_cache/cache[0][86] ) );
  DFFRX1 \D_cache/cache_reg[4][86]  ( .D(\D_cache/n1104 ), .CK(clk), .RN(n4211), .Q(\D_cache/cache[4][86] ) );
  DFFRX1 \D_cache/cache_reg[0][87]  ( .D(\D_cache/n1100 ), .CK(clk), .RN(n4212), .Q(\D_cache/cache[0][87] ) );
  DFFRX1 \D_cache/cache_reg[4][87]  ( .D(\D_cache/n1096 ), .CK(clk), .RN(n4212), .Q(\D_cache/cache[4][87] ) );
  DFFRX1 \D_cache/cache_reg[0][88]  ( .D(\D_cache/n1092 ), .CK(clk), .RN(n4212), .Q(\D_cache/cache[0][88] ) );
  DFFRX1 \D_cache/cache_reg[4][88]  ( .D(\D_cache/n1088 ), .CK(clk), .RN(n4213), .Q(\D_cache/cache[4][88] ) );
  DFFRX1 \D_cache/cache_reg[0][89]  ( .D(\D_cache/n1084 ), .CK(clk), .RN(n4213), .Q(\D_cache/cache[0][89] ) );
  DFFRX1 \D_cache/cache_reg[4][89]  ( .D(\D_cache/n1080 ), .CK(clk), .RN(n4213), .Q(\D_cache/cache[4][89] ) );
  DFFRX1 \D_cache/cache_reg[0][90]  ( .D(\D_cache/n1076 ), .CK(clk), .RN(n4214), .Q(\D_cache/cache[0][90] ) );
  DFFRX1 \D_cache/cache_reg[4][90]  ( .D(\D_cache/n1072 ), .CK(clk), .RN(n4214), .Q(\D_cache/cache[4][90] ) );
  DFFRX1 \D_cache/cache_reg[0][91]  ( .D(\D_cache/n1068 ), .CK(clk), .RN(n4214), .Q(\D_cache/cache[0][91] ) );
  DFFRX1 \D_cache/cache_reg[4][91]  ( .D(\D_cache/n1064 ), .CK(clk), .RN(n4215), .Q(\D_cache/cache[4][91] ) );
  DFFRX1 \D_cache/cache_reg[0][92]  ( .D(\D_cache/n1060 ), .CK(clk), .RN(n4215), .Q(\D_cache/cache[0][92] ) );
  DFFRX1 \D_cache/cache_reg[4][92]  ( .D(\D_cache/n1056 ), .CK(clk), .RN(n4215), .Q(\D_cache/cache[4][92] ) );
  DFFRX1 \D_cache/cache_reg[0][93]  ( .D(\D_cache/n1052 ), .CK(clk), .RN(n4216), .Q(\D_cache/cache[0][93] ) );
  DFFRX1 \D_cache/cache_reg[4][93]  ( .D(\D_cache/n1048 ), .CK(clk), .RN(n4216), .Q(\D_cache/cache[4][93] ) );
  DFFRX1 \D_cache/cache_reg[0][94]  ( .D(\D_cache/n1044 ), .CK(clk), .RN(n4216), .Q(\D_cache/cache[0][94] ) );
  DFFRX1 \D_cache/cache_reg[4][94]  ( .D(\D_cache/n1040 ), .CK(clk), .RN(n4217), .Q(\D_cache/cache[4][94] ) );
  DFFRX1 \D_cache/cache_reg[0][95]  ( .D(\D_cache/n1036 ), .CK(clk), .RN(n4217), .Q(\D_cache/cache[0][95] ) );
  DFFRX1 \D_cache/cache_reg[4][95]  ( .D(\D_cache/n1032 ), .CK(clk), .RN(n4217), .Q(\D_cache/cache[4][95] ) );
  DFFRX1 \D_cache/cache_reg[0][97]  ( .D(\D_cache/n1020 ), .CK(clk), .RN(n4218), .Q(\D_cache/cache[0][97] ) );
  DFFRX1 \D_cache/cache_reg[4][97]  ( .D(\D_cache/n1016 ), .CK(clk), .RN(n4219), .Q(\D_cache/cache[4][97] ) );
  DFFRX1 \D_cache/cache_reg[0][111]  ( .D(\D_cache/n908 ), .CK(clk), .RN(n4228), .Q(\D_cache/cache[0][111] ) );
  DFFRX1 \D_cache/cache_reg[4][111]  ( .D(\D_cache/n904 ), .CK(clk), .RN(n4228), .Q(\D_cache/cache[4][111] ) );
  DFFRX1 \D_cache/cache_reg[0][112]  ( .D(\D_cache/n900 ), .CK(clk), .RN(n4228), .Q(\D_cache/cache[0][112] ) );
  DFFRX1 \D_cache/cache_reg[4][112]  ( .D(\D_cache/n896 ), .CK(clk), .RN(n4229), .Q(\D_cache/cache[4][112] ) );
  DFFRX1 \D_cache/cache_reg[0][113]  ( .D(\D_cache/n892 ), .CK(clk), .RN(n4229), .Q(\D_cache/cache[0][113] ) );
  DFFRX1 \D_cache/cache_reg[4][113]  ( .D(\D_cache/n888 ), .CK(clk), .RN(n4229), .Q(\D_cache/cache[4][113] ) );
  DFFRX1 \D_cache/cache_reg[0][114]  ( .D(\D_cache/n884 ), .CK(clk), .RN(n4230), .Q(\D_cache/cache[0][114] ) );
  DFFRX1 \D_cache/cache_reg[4][114]  ( .D(\D_cache/n880 ), .CK(clk), .RN(n4230), .Q(\D_cache/cache[4][114] ) );
  DFFRX1 \D_cache/cache_reg[0][115]  ( .D(\D_cache/n876 ), .CK(clk), .RN(n4230), .Q(\D_cache/cache[0][115] ) );
  DFFRX1 \D_cache/cache_reg[4][115]  ( .D(\D_cache/n872 ), .CK(clk), .RN(n4231), .Q(\D_cache/cache[4][115] ) );
  DFFRX1 \D_cache/cache_reg[0][116]  ( .D(\D_cache/n868 ), .CK(clk), .RN(n4231), .Q(\D_cache/cache[0][116] ) );
  DFFRX1 \D_cache/cache_reg[4][116]  ( .D(\D_cache/n864 ), .CK(clk), .RN(n4231), .Q(\D_cache/cache[4][116] ) );
  DFFRX1 \D_cache/cache_reg[0][117]  ( .D(\D_cache/n860 ), .CK(clk), .RN(n4232), .Q(\D_cache/cache[0][117] ) );
  DFFRX1 \D_cache/cache_reg[4][117]  ( .D(\D_cache/n856 ), .CK(clk), .RN(n4232), .Q(\D_cache/cache[4][117] ) );
  DFFRX1 \D_cache/cache_reg[0][119]  ( .D(\D_cache/n844 ), .CK(clk), .RN(n4233), .Q(\D_cache/cache[0][119] ) );
  DFFRX1 \D_cache/cache_reg[4][119]  ( .D(\D_cache/n840 ), .CK(clk), .RN(n4233), .Q(\D_cache/cache[4][119] ) );
  DFFRX1 \D_cache/cache_reg[0][120]  ( .D(\D_cache/n836 ), .CK(clk), .RN(n4234), .Q(\D_cache/cache[0][120] ) );
  DFFRX1 \D_cache/cache_reg[4][120]  ( .D(\D_cache/n832 ), .CK(clk), .RN(n4234), .Q(\D_cache/cache[4][120] ) );
  DFFRX1 \D_cache/cache_reg[0][121]  ( .D(\D_cache/n828 ), .CK(clk), .RN(n4234), .Q(\D_cache/cache[0][121] ) );
  DFFRX1 \D_cache/cache_reg[4][121]  ( .D(\D_cache/n824 ), .CK(clk), .RN(n4235), .Q(\D_cache/cache[4][121] ) );
  DFFRX1 \D_cache/cache_reg[0][122]  ( .D(\D_cache/n820 ), .CK(clk), .RN(n4235), .Q(\D_cache/cache[0][122] ) );
  DFFRX1 \D_cache/cache_reg[4][122]  ( .D(\D_cache/n816 ), .CK(clk), .RN(n4235), .Q(\D_cache/cache[4][122] ) );
  DFFRX1 \D_cache/cache_reg[0][123]  ( .D(\D_cache/n812 ), .CK(clk), .RN(n4236), .Q(\D_cache/cache[0][123] ) );
  DFFRX1 \D_cache/cache_reg[4][123]  ( .D(\D_cache/n808 ), .CK(clk), .RN(n4236), .Q(\D_cache/cache[4][123] ) );
  DFFRX1 \D_cache/cache_reg[0][124]  ( .D(\D_cache/n804 ), .CK(clk), .RN(n4236), .Q(\D_cache/cache[0][124] ) );
  DFFRX1 \D_cache/cache_reg[4][124]  ( .D(\D_cache/n800 ), .CK(clk), .RN(n4237), .Q(\D_cache/cache[4][124] ) );
  DFFRX1 \D_cache/cache_reg[0][125]  ( .D(\D_cache/n796 ), .CK(clk), .RN(n4237), .Q(\D_cache/cache[0][125] ) );
  DFFRX1 \D_cache/cache_reg[4][125]  ( .D(\D_cache/n792 ), .CK(clk), .RN(n4237), .Q(\D_cache/cache[4][125] ) );
  DFFRX1 \D_cache/cache_reg[0][126]  ( .D(\D_cache/n788 ), .CK(clk), .RN(n4238), .Q(\D_cache/cache[0][126] ) );
  DFFRX1 \D_cache/cache_reg[4][126]  ( .D(\D_cache/n784 ), .CK(clk), .RN(n4238), .Q(\D_cache/cache[4][126] ) );
  DFFRX1 \D_cache/cache_reg[0][127]  ( .D(\D_cache/n780 ), .CK(clk), .RN(n4238), .Q(\D_cache/cache[0][127] ) );
  DFFRX1 \D_cache/cache_reg[4][127]  ( .D(\D_cache/n776 ), .CK(clk), .RN(n4239), .Q(\D_cache/cache[4][127] ) );
  DFFRX1 \D_cache/cache_reg[2][15]  ( .D(\D_cache/n1674 ), .CK(clk), .RN(n4164), .Q(\D_cache/cache[2][15] ) );
  DFFRX1 \D_cache/cache_reg[2][16]  ( .D(\D_cache/n1666 ), .CK(clk), .RN(n4164), .Q(\D_cache/cache[2][16] ) );
  DFFRX1 \D_cache/cache_reg[6][16]  ( .D(\D_cache/n1662 ), .CK(clk), .RN(n4165), .Q(\D_cache/cache[6][16] ) );
  DFFRX1 \D_cache/cache_reg[2][29]  ( .D(\D_cache/n1562 ), .CK(clk), .RN(n4173), .Q(\D_cache/cache[2][29] ) );
  DFFRX1 \D_cache/cache_reg[6][29]  ( .D(\D_cache/n1558 ), .CK(clk), .RN(n4173), .Q(\D_cache/cache[6][29] ) );
  DFFRX1 \D_cache/cache_reg[2][30]  ( .D(\D_cache/n1554 ), .CK(clk), .RN(n4174), .Q(\D_cache/cache[2][30] ) );
  DFFRX1 \D_cache/cache_reg[6][30]  ( .D(\D_cache/n1550 ), .CK(clk), .RN(n4174), .Q(\D_cache/cache[6][30] ) );
  DFFRX1 \D_cache/cache_reg[2][32]  ( .D(\D_cache/n1538 ), .CK(clk), .RN(n4175), .Q(\D_cache/cache[2][32] ) );
  DFFRX1 \D_cache/cache_reg[6][32]  ( .D(\D_cache/n1534 ), .CK(clk), .RN(n4175), .Q(\D_cache/cache[6][32] ) );
  DFFRX1 \D_cache/cache_reg[2][33]  ( .D(\D_cache/n1530 ), .CK(clk), .RN(n4176), .Q(\D_cache/cache[2][33] ) );
  DFFRX1 \D_cache/cache_reg[6][33]  ( .D(\D_cache/n1526 ), .CK(clk), .RN(n4176), .Q(\D_cache/cache[6][33] ) );
  DFFRX1 \D_cache/cache_reg[2][34]  ( .D(\D_cache/n1522 ), .CK(clk), .RN(n4176), .Q(\D_cache/cache[2][34] ) );
  DFFRX1 \D_cache/cache_reg[6][34]  ( .D(\D_cache/n1518 ), .CK(clk), .RN(n4177), .Q(\D_cache/cache[6][34] ) );
  DFFRX1 \D_cache/cache_reg[2][35]  ( .D(\D_cache/n1514 ), .CK(clk), .RN(n4177), .Q(\D_cache/cache[2][35] ) );
  DFFRX1 \D_cache/cache_reg[6][35]  ( .D(\D_cache/n1510 ), .CK(clk), .RN(n4177), .Q(\D_cache/cache[6][35] ) );
  DFFRX1 \D_cache/cache_reg[2][36]  ( .D(\D_cache/n1506 ), .CK(clk), .RN(n4178), .Q(\D_cache/cache[2][36] ) );
  DFFRX1 \D_cache/cache_reg[6][36]  ( .D(\D_cache/n1502 ), .CK(clk), .RN(n4178), .Q(\D_cache/cache[6][36] ) );
  DFFRX1 \D_cache/cache_reg[2][37]  ( .D(\D_cache/n1498 ), .CK(clk), .RN(n4178), .Q(\D_cache/cache[2][37] ) );
  DFFRX1 \D_cache/cache_reg[6][37]  ( .D(\D_cache/n1494 ), .CK(clk), .RN(n4179), .Q(\D_cache/cache[6][37] ) );
  DFFRX1 \D_cache/cache_reg[2][38]  ( .D(\D_cache/n1490 ), .CK(clk), .RN(n4179), .Q(\D_cache/cache[2][38] ) );
  DFFRX1 \D_cache/cache_reg[6][38]  ( .D(\D_cache/n1486 ), .CK(clk), .RN(n4179), .Q(\D_cache/cache[6][38] ) );
  DFFRX1 \D_cache/cache_reg[2][40]  ( .D(\D_cache/n1474 ), .CK(clk), .RN(n4180), .Q(\D_cache/cache[2][40] ) );
  DFFRX1 \D_cache/cache_reg[6][40]  ( .D(\D_cache/n1470 ), .CK(clk), .RN(n4181), .Q(\D_cache/cache[6][40] ) );
  DFFRX1 \D_cache/cache_reg[2][42]  ( .D(\D_cache/n1458 ), .CK(clk), .RN(n4182), .Q(\D_cache/cache[2][42] ) );
  DFFRX1 \D_cache/cache_reg[6][42]  ( .D(\D_cache/n1454 ), .CK(clk), .RN(n4182), .Q(\D_cache/cache[6][42] ) );
  DFFRX1 \D_cache/cache_reg[2][44]  ( .D(\D_cache/n1442 ), .CK(clk), .RN(n4183), .Q(\D_cache/cache[2][44] ) );
  DFFRX1 \D_cache/cache_reg[6][44]  ( .D(\D_cache/n1438 ), .CK(clk), .RN(n4183), .Q(\D_cache/cache[6][44] ) );
  DFFRX1 \D_cache/cache_reg[2][46]  ( .D(\D_cache/n1426 ), .CK(clk), .RN(n4184), .Q(\D_cache/cache[2][46] ) );
  DFFRX1 \D_cache/cache_reg[6][46]  ( .D(\D_cache/n1422 ), .CK(clk), .RN(n4185), .Q(\D_cache/cache[6][46] ) );
  DFFRX1 \D_cache/cache_reg[2][47]  ( .D(\D_cache/n1418 ), .CK(clk), .RN(n4185), .Q(\D_cache/cache[2][47] ) );
  DFFRX1 \D_cache/cache_reg[6][47]  ( .D(\D_cache/n1414 ), .CK(clk), .RN(n4185), .Q(\D_cache/cache[6][47] ) );
  DFFRX1 \D_cache/cache_reg[2][48]  ( .D(\D_cache/n1410 ), .CK(clk), .RN(n4186), .Q(\D_cache/cache[2][48] ) );
  DFFRX1 \D_cache/cache_reg[6][48]  ( .D(\D_cache/n1406 ), .CK(clk), .RN(n4186), .Q(\D_cache/cache[6][48] ) );
  DFFRX1 \D_cache/cache_reg[2][49]  ( .D(\D_cache/n1402 ), .CK(clk), .RN(n4186), .Q(\D_cache/cache[2][49] ) );
  DFFRX1 \D_cache/cache_reg[6][49]  ( .D(\D_cache/n1398 ), .CK(clk), .RN(n4187), .Q(\D_cache/cache[6][49] ) );
  DFFRX1 \D_cache/cache_reg[2][50]  ( .D(\D_cache/n1394 ), .CK(clk), .RN(n4187), .Q(\D_cache/cache[2][50] ) );
  DFFRX1 \D_cache/cache_reg[6][50]  ( .D(\D_cache/n1390 ), .CK(clk), .RN(n4187), .Q(\D_cache/cache[6][50] ) );
  DFFRX1 \D_cache/cache_reg[2][51]  ( .D(\D_cache/n1386 ), .CK(clk), .RN(n4188), .Q(\D_cache/cache[2][51] ) );
  DFFRX1 \D_cache/cache_reg[6][51]  ( .D(\D_cache/n1382 ), .CK(clk), .RN(n4188), .Q(\D_cache/cache[6][51] ) );
  DFFRX1 \D_cache/cache_reg[2][52]  ( .D(\D_cache/n1378 ), .CK(clk), .RN(n4188), .Q(\D_cache/cache[2][52] ) );
  DFFRX1 \D_cache/cache_reg[6][52]  ( .D(\D_cache/n1374 ), .CK(clk), .RN(n4189), .Q(\D_cache/cache[6][52] ) );
  DFFRX1 \D_cache/cache_reg[6][53]  ( .D(\D_cache/n1366 ), .CK(clk), .RN(n4189), .Q(\D_cache/cache[6][53] ) );
  DFFRX1 \D_cache/cache_reg[2][55]  ( .D(\D_cache/n1354 ), .CK(clk), .RN(n4190), .Q(\D_cache/cache[2][55] ) );
  DFFRX1 \D_cache/cache_reg[6][55]  ( .D(\D_cache/n1350 ), .CK(clk), .RN(n4191), .Q(\D_cache/cache[6][55] ) );
  DFFRX1 \D_cache/cache_reg[2][56]  ( .D(\D_cache/n1346 ), .CK(clk), .RN(n4191), .Q(\D_cache/cache[2][56] ) );
  DFFRX1 \D_cache/cache_reg[6][56]  ( .D(\D_cache/n1342 ), .CK(clk), .RN(n4191), .Q(\D_cache/cache[6][56] ) );
  DFFRX1 \D_cache/cache_reg[2][57]  ( .D(\D_cache/n1338 ), .CK(clk), .RN(n4192), .Q(\D_cache/cache[2][57] ) );
  DFFRX1 \D_cache/cache_reg[6][57]  ( .D(\D_cache/n1334 ), .CK(clk), .RN(n4192), .Q(\D_cache/cache[6][57] ) );
  DFFRX1 \D_cache/cache_reg[2][58]  ( .D(\D_cache/n1330 ), .CK(clk), .RN(n4192), .Q(\D_cache/cache[2][58] ) );
  DFFRX1 \D_cache/cache_reg[6][58]  ( .D(\D_cache/n1326 ), .CK(clk), .RN(n4193), .Q(\D_cache/cache[6][58] ) );
  DFFRX1 \D_cache/cache_reg[2][59]  ( .D(\D_cache/n1322 ), .CK(clk), .RN(n4193), .Q(\D_cache/cache[2][59] ) );
  DFFRX1 \D_cache/cache_reg[6][59]  ( .D(\D_cache/n1318 ), .CK(clk), .RN(n4193), .Q(\D_cache/cache[6][59] ) );
  DFFRX1 \D_cache/cache_reg[2][60]  ( .D(\D_cache/n1314 ), .CK(clk), .RN(n4194), .Q(\D_cache/cache[2][60] ) );
  DFFRX1 \D_cache/cache_reg[6][60]  ( .D(\D_cache/n1310 ), .CK(clk), .RN(n4194), .Q(\D_cache/cache[6][60] ) );
  DFFRX1 \D_cache/cache_reg[2][61]  ( .D(\D_cache/n1306 ), .CK(clk), .RN(n4194), .Q(\D_cache/cache[2][61] ) );
  DFFRX1 \D_cache/cache_reg[6][61]  ( .D(\D_cache/n1302 ), .CK(clk), .RN(n4195), .Q(\D_cache/cache[6][61] ) );
  DFFRX1 \D_cache/cache_reg[2][62]  ( .D(\D_cache/n1298 ), .CK(clk), .RN(n4195), .Q(\D_cache/cache[2][62] ) );
  DFFRX1 \D_cache/cache_reg[6][62]  ( .D(\D_cache/n1294 ), .CK(clk), .RN(n4195), .Q(\D_cache/cache[6][62] ) );
  DFFRX1 \D_cache/cache_reg[2][63]  ( .D(\D_cache/n1290 ), .CK(clk), .RN(n4196), .Q(\D_cache/cache[2][63] ) );
  DFFRX1 \D_cache/cache_reg[6][63]  ( .D(\D_cache/n1286 ), .CK(clk), .RN(n4196), .Q(\D_cache/cache[6][63] ) );
  DFFRX1 \D_cache/cache_reg[2][64]  ( .D(\D_cache/n1282 ), .CK(clk), .RN(n4196), .Q(\D_cache/cache[2][64] ) );
  DFFRX1 \D_cache/cache_reg[6][64]  ( .D(\D_cache/n1278 ), .CK(clk), .RN(n4197), .Q(\D_cache/cache[6][64] ) );
  DFFRX1 \D_cache/cache_reg[2][65]  ( .D(\D_cache/n1274 ), .CK(clk), .RN(n4197), .Q(\D_cache/cache[2][65] ) );
  DFFRX1 \D_cache/cache_reg[6][65]  ( .D(\D_cache/n1270 ), .CK(clk), .RN(n4197), .Q(\D_cache/cache[6][65] ) );
  DFFRX1 \D_cache/cache_reg[2][66]  ( .D(\D_cache/n1266 ), .CK(clk), .RN(n4198), .Q(\D_cache/cache[2][66] ) );
  DFFRX1 \D_cache/cache_reg[6][66]  ( .D(\D_cache/n1262 ), .CK(clk), .RN(n4198), .Q(\D_cache/cache[6][66] ) );
  DFFRX1 \D_cache/cache_reg[2][67]  ( .D(\D_cache/n1258 ), .CK(clk), .RN(n4198), .Q(\D_cache/cache[2][67] ) );
  DFFRX1 \D_cache/cache_reg[6][67]  ( .D(\D_cache/n1254 ), .CK(clk), .RN(n4199), .Q(\D_cache/cache[6][67] ) );
  DFFRX1 \D_cache/cache_reg[2][68]  ( .D(\D_cache/n1250 ), .CK(clk), .RN(n4199), .Q(\D_cache/cache[2][68] ) );
  DFFRX1 \D_cache/cache_reg[6][68]  ( .D(\D_cache/n1246 ), .CK(clk), .RN(n4199), .Q(\D_cache/cache[6][68] ) );
  DFFRX1 \D_cache/cache_reg[2][78]  ( .D(\D_cache/n1170 ), .CK(clk), .RN(n4206), .Q(\D_cache/cache[2][78] ) );
  DFFRX1 \D_cache/cache_reg[6][78]  ( .D(\D_cache/n1166 ), .CK(clk), .RN(n4206), .Q(\D_cache/cache[6][78] ) );
  DFFRX1 \D_cache/cache_reg[2][79]  ( .D(\D_cache/n1162 ), .CK(clk), .RN(n4206), .Q(\D_cache/cache[2][79] ) );
  DFFRX1 \D_cache/cache_reg[6][79]  ( .D(\D_cache/n1158 ), .CK(clk), .RN(n4207), .Q(\D_cache/cache[6][79] ) );
  DFFRX1 \D_cache/cache_reg[2][80]  ( .D(\D_cache/n1154 ), .CK(clk), .RN(n4207), .Q(\D_cache/cache[2][80] ) );
  DFFRX1 \D_cache/cache_reg[6][80]  ( .D(\D_cache/n1150 ), .CK(clk), .RN(n4207), .Q(\D_cache/cache[6][80] ) );
  DFFRX1 \D_cache/cache_reg[2][81]  ( .D(\D_cache/n1146 ), .CK(clk), .RN(n4208), .Q(\D_cache/cache[2][81] ) );
  DFFRX1 \D_cache/cache_reg[6][81]  ( .D(\D_cache/n1142 ), .CK(clk), .RN(n4208), .Q(\D_cache/cache[6][81] ) );
  DFFRX1 \D_cache/cache_reg[2][82]  ( .D(\D_cache/n1138 ), .CK(clk), .RN(n4208), .Q(\D_cache/cache[2][82] ) );
  DFFRX1 \D_cache/cache_reg[6][82]  ( .D(\D_cache/n1134 ), .CK(clk), .RN(n4209), .Q(\D_cache/cache[6][82] ) );
  DFFRX1 \D_cache/cache_reg[2][83]  ( .D(\D_cache/n1130 ), .CK(clk), .RN(n4209), .Q(\D_cache/cache[2][83] ) );
  DFFRX1 \D_cache/cache_reg[6][83]  ( .D(\D_cache/n1126 ), .CK(clk), .RN(n4209), .Q(\D_cache/cache[6][83] ) );
  DFFRX1 \D_cache/cache_reg[2][84]  ( .D(\D_cache/n1122 ), .CK(clk), .RN(n4210), .Q(\D_cache/cache[2][84] ) );
  DFFRX1 \D_cache/cache_reg[6][84]  ( .D(\D_cache/n1118 ), .CK(clk), .RN(n4210), .Q(\D_cache/cache[6][84] ) );
  DFFRX1 \D_cache/cache_reg[2][85]  ( .D(\D_cache/n1114 ), .CK(clk), .RN(n4210), .Q(\D_cache/cache[2][85] ) );
  DFFRX1 \D_cache/cache_reg[6][85]  ( .D(\D_cache/n1110 ), .CK(clk), .RN(n4211), .Q(\D_cache/cache[6][85] ) );
  DFFRX1 \D_cache/cache_reg[2][86]  ( .D(\D_cache/n1106 ), .CK(clk), .RN(n4211), .Q(\D_cache/cache[2][86] ) );
  DFFRX1 \D_cache/cache_reg[6][86]  ( .D(\D_cache/n1102 ), .CK(clk), .RN(n4211), .Q(\D_cache/cache[6][86] ) );
  DFFRX1 \D_cache/cache_reg[2][87]  ( .D(\D_cache/n1098 ), .CK(clk), .RN(n4212), .Q(\D_cache/cache[2][87] ) );
  DFFRX1 \D_cache/cache_reg[6][87]  ( .D(\D_cache/n1094 ), .CK(clk), .RN(n4212), .Q(\D_cache/cache[6][87] ) );
  DFFRX1 \D_cache/cache_reg[2][88]  ( .D(\D_cache/n1090 ), .CK(clk), .RN(n4212), .Q(\D_cache/cache[2][88] ) );
  DFFRX1 \D_cache/cache_reg[6][88]  ( .D(\D_cache/n1086 ), .CK(clk), .RN(n4213), .Q(\D_cache/cache[6][88] ) );
  DFFRX1 \D_cache/cache_reg[2][89]  ( .D(\D_cache/n1082 ), .CK(clk), .RN(n4213), .Q(\D_cache/cache[2][89] ) );
  DFFRX1 \D_cache/cache_reg[6][89]  ( .D(\D_cache/n1078 ), .CK(clk), .RN(n4213), .Q(\D_cache/cache[6][89] ) );
  DFFRX1 \D_cache/cache_reg[2][90]  ( .D(\D_cache/n1074 ), .CK(clk), .RN(n4214), .Q(\D_cache/cache[2][90] ) );
  DFFRX1 \D_cache/cache_reg[6][90]  ( .D(\D_cache/n1070 ), .CK(clk), .RN(n4214), .Q(\D_cache/cache[6][90] ) );
  DFFRX1 \D_cache/cache_reg[2][91]  ( .D(\D_cache/n1066 ), .CK(clk), .RN(n4214), .Q(\D_cache/cache[2][91] ) );
  DFFRX1 \D_cache/cache_reg[6][91]  ( .D(\D_cache/n1062 ), .CK(clk), .RN(n4215), .Q(\D_cache/cache[6][91] ) );
  DFFRX1 \D_cache/cache_reg[2][92]  ( .D(\D_cache/n1058 ), .CK(clk), .RN(n4215), .Q(\D_cache/cache[2][92] ) );
  DFFRX1 \D_cache/cache_reg[6][92]  ( .D(\D_cache/n1054 ), .CK(clk), .RN(n4215), .Q(\D_cache/cache[6][92] ) );
  DFFRX1 \D_cache/cache_reg[2][93]  ( .D(\D_cache/n1050 ), .CK(clk), .RN(n4216), .Q(\D_cache/cache[2][93] ) );
  DFFRX1 \D_cache/cache_reg[6][93]  ( .D(\D_cache/n1046 ), .CK(clk), .RN(n4216), .Q(\D_cache/cache[6][93] ) );
  DFFRX1 \D_cache/cache_reg[2][94]  ( .D(\D_cache/n1042 ), .CK(clk), .RN(n4216), .Q(\D_cache/cache[2][94] ) );
  DFFRX1 \D_cache/cache_reg[6][94]  ( .D(\D_cache/n1038 ), .CK(clk), .RN(n4217), .Q(\D_cache/cache[6][94] ) );
  DFFRX1 \D_cache/cache_reg[2][95]  ( .D(\D_cache/n1034 ), .CK(clk), .RN(n4217), .Q(\D_cache/cache[2][95] ) );
  DFFRX1 \D_cache/cache_reg[6][95]  ( .D(\D_cache/n1030 ), .CK(clk), .RN(n4217), .Q(\D_cache/cache[6][95] ) );
  DFFRX1 \D_cache/cache_reg[2][97]  ( .D(\D_cache/n1018 ), .CK(clk), .RN(n4218), .Q(\D_cache/cache[2][97] ) );
  DFFRX1 \D_cache/cache_reg[6][97]  ( .D(\D_cache/n1014 ), .CK(clk), .RN(n4219), .Q(\D_cache/cache[6][97] ) );
  DFFRX1 \D_cache/cache_reg[2][99]  ( .D(\D_cache/n1002 ), .CK(clk), .RN(n4220), .Q(\D_cache/cache[2][99] ) );
  DFFRX1 \D_cache/cache_reg[2][111]  ( .D(\D_cache/n906 ), .CK(clk), .RN(n4228), .Q(\D_cache/cache[2][111] ) );
  DFFRX1 \D_cache/cache_reg[6][111]  ( .D(\D_cache/n902 ), .CK(clk), .RN(n4228), .Q(\D_cache/cache[6][111] ) );
  DFFRX1 \D_cache/cache_reg[2][112]  ( .D(\D_cache/n898 ), .CK(clk), .RN(n4228), .Q(\D_cache/cache[2][112] ) );
  DFFRX1 \D_cache/cache_reg[6][112]  ( .D(\D_cache/n894 ), .CK(clk), .RN(n4229), .Q(\D_cache/cache[6][112] ) );
  DFFRX1 \D_cache/cache_reg[2][113]  ( .D(\D_cache/n890 ), .CK(clk), .RN(n4229), .Q(\D_cache/cache[2][113] ) );
  DFFRX1 \D_cache/cache_reg[6][113]  ( .D(\D_cache/n886 ), .CK(clk), .RN(n4229), .Q(\D_cache/cache[6][113] ) );
  DFFRX1 \D_cache/cache_reg[2][114]  ( .D(\D_cache/n882 ), .CK(clk), .RN(n4230), .Q(\D_cache/cache[2][114] ) );
  DFFRX1 \D_cache/cache_reg[6][114]  ( .D(\D_cache/n878 ), .CK(clk), .RN(n4230), .Q(\D_cache/cache[6][114] ) );
  DFFRX1 \D_cache/cache_reg[2][115]  ( .D(\D_cache/n874 ), .CK(clk), .RN(n4230), .Q(\D_cache/cache[2][115] ) );
  DFFRX1 \D_cache/cache_reg[6][115]  ( .D(\D_cache/n870 ), .CK(clk), .RN(n4231), .Q(\D_cache/cache[6][115] ) );
  DFFRX1 \D_cache/cache_reg[2][116]  ( .D(\D_cache/n866 ), .CK(clk), .RN(n4231), .Q(\D_cache/cache[2][116] ) );
  DFFRX1 \D_cache/cache_reg[6][116]  ( .D(\D_cache/n862 ), .CK(clk), .RN(n4231), .Q(\D_cache/cache[6][116] ) );
  DFFRX1 \D_cache/cache_reg[2][117]  ( .D(\D_cache/n858 ), .CK(clk), .RN(n4232), .Q(\D_cache/cache[2][117] ) );
  DFFRX1 \D_cache/cache_reg[6][117]  ( .D(\D_cache/n854 ), .CK(clk), .RN(n4232), .Q(\D_cache/cache[6][117] ) );
  DFFRX1 \D_cache/cache_reg[2][119]  ( .D(\D_cache/n842 ), .CK(clk), .RN(n4233), .Q(\D_cache/cache[2][119] ) );
  DFFRX1 \D_cache/cache_reg[6][119]  ( .D(\D_cache/n838 ), .CK(clk), .RN(n4233), .Q(\D_cache/cache[6][119] ) );
  DFFRX1 \D_cache/cache_reg[2][120]  ( .D(\D_cache/n834 ), .CK(clk), .RN(n4234), .Q(\D_cache/cache[2][120] ) );
  DFFRX1 \D_cache/cache_reg[6][120]  ( .D(\D_cache/n830 ), .CK(clk), .RN(n4234), .Q(\D_cache/cache[6][120] ) );
  DFFRX1 \D_cache/cache_reg[2][121]  ( .D(\D_cache/n826 ), .CK(clk), .RN(n4234), .Q(\D_cache/cache[2][121] ) );
  DFFRX1 \D_cache/cache_reg[6][121]  ( .D(\D_cache/n822 ), .CK(clk), .RN(n4235), .Q(\D_cache/cache[6][121] ) );
  DFFRX1 \D_cache/cache_reg[2][122]  ( .D(\D_cache/n818 ), .CK(clk), .RN(n4235), .Q(\D_cache/cache[2][122] ) );
  DFFRX1 \D_cache/cache_reg[6][122]  ( .D(\D_cache/n814 ), .CK(clk), .RN(n4235), .Q(\D_cache/cache[6][122] ) );
  DFFRX1 \D_cache/cache_reg[2][123]  ( .D(\D_cache/n810 ), .CK(clk), .RN(n4236), .Q(\D_cache/cache[2][123] ) );
  DFFRX1 \D_cache/cache_reg[6][123]  ( .D(\D_cache/n806 ), .CK(clk), .RN(n4236), .Q(\D_cache/cache[6][123] ) );
  DFFRX1 \D_cache/cache_reg[2][124]  ( .D(\D_cache/n802 ), .CK(clk), .RN(n4236), .Q(\D_cache/cache[2][124] ) );
  DFFRX1 \D_cache/cache_reg[6][124]  ( .D(\D_cache/n798 ), .CK(clk), .RN(n4237), .Q(\D_cache/cache[6][124] ) );
  DFFRX1 \D_cache/cache_reg[2][125]  ( .D(\D_cache/n794 ), .CK(clk), .RN(n4237), .Q(\D_cache/cache[2][125] ) );
  DFFRX1 \D_cache/cache_reg[6][125]  ( .D(\D_cache/n790 ), .CK(clk), .RN(n4237), .Q(\D_cache/cache[6][125] ) );
  DFFRX1 \D_cache/cache_reg[2][126]  ( .D(\D_cache/n786 ), .CK(clk), .RN(n4238), .Q(\D_cache/cache[2][126] ) );
  DFFRX1 \D_cache/cache_reg[6][126]  ( .D(\D_cache/n782 ), .CK(clk), .RN(n4238), .Q(\D_cache/cache[6][126] ) );
  DFFRX1 \D_cache/cache_reg[2][127]  ( .D(\D_cache/n778 ), .CK(clk), .RN(n4238), .Q(\D_cache/cache[2][127] ) );
  DFFRX1 \D_cache/cache_reg[6][127]  ( .D(\D_cache/n774 ), .CK(clk), .RN(n4239), .Q(\D_cache/cache[6][127] ) );
  DFFRX1 \i_MIPS/Register/register_reg[29][2]  ( .D(\i_MIPS/Register/n182 ), 
        .CK(clk), .RN(n4074), .Q(\i_MIPS/Register/register[29][2] ), .QN(n283)
         );
  DFFRX1 \i_MIPS/Register/register_reg[29][3]  ( .D(\i_MIPS/Register/n183 ), 
        .CK(clk), .RN(n4074), .Q(\i_MIPS/Register/register[29][3] ), .QN(n288)
         );
  DFFRX1 \i_MIPS/Register/register_reg[29][4]  ( .D(\i_MIPS/Register/n184 ), 
        .CK(clk), .RN(n4074), .Q(\i_MIPS/Register/register[29][4] ), .QN(n245)
         );
  DFFRX1 \i_MIPS/Register/register_reg[29][7]  ( .D(\i_MIPS/Register/n187 ), 
        .CK(clk), .RN(n4074), .Q(\i_MIPS/Register/register[29][7] ), .QN(n263)
         );
  DFFRX1 \i_MIPS/Register/register_reg[29][11]  ( .D(\i_MIPS/Register/n191 ), 
        .CK(clk), .RN(n4074), .Q(\i_MIPS/Register/register[29][11] ), .QN(
        n1109) );
  DFFRX1 \i_MIPS/Register/register_reg[29][12]  ( .D(\i_MIPS/Register/n192 ), 
        .CK(clk), .RN(n4075), .Q(\i_MIPS/Register/register[29][12] ), .QN(n230) );
  DFFRX1 \i_MIPS/Register/register_reg[29][13]  ( .D(\i_MIPS/Register/n193 ), 
        .CK(clk), .RN(n4075), .Q(\i_MIPS/Register/register[29][13] ), .QN(n215) );
  DFFRX1 \i_MIPS/Register/register_reg[29][15]  ( .D(\i_MIPS/Register/n195 ), 
        .CK(clk), .RN(n4075), .Q(\i_MIPS/Register/register[29][15] ), .QN(n298) );
  DFFRX1 \i_MIPS/Register/register_reg[29][16]  ( .D(\i_MIPS/Register/n196 ), 
        .CK(clk), .RN(n4075), .Q(\i_MIPS/Register/register[29][16] ), .QN(n318) );
  DFFRX1 \i_MIPS/Register/register_reg[29][17]  ( .D(\i_MIPS/Register/n197 ), 
        .CK(clk), .RN(n4075), .Q(\i_MIPS/Register/register[29][17] ), .QN(n373) );
  DFFRX1 \i_MIPS/Register/register_reg[29][18]  ( .D(\i_MIPS/Register/n198 ), 
        .CK(clk), .RN(n4075), .Q(\i_MIPS/Register/register[29][18] ), .QN(n368) );
  DFFRX1 \i_MIPS/Register/register_reg[29][19]  ( .D(\i_MIPS/Register/n199 ), 
        .CK(clk), .RN(n4075), .Q(\i_MIPS/Register/register[29][19] ), .QN(n323) );
  DFFRX1 \i_MIPS/Register/register_reg[29][20]  ( .D(\i_MIPS/Register/n200 ), 
        .CK(clk), .RN(n4075), .Q(\i_MIPS/Register/register[29][20] ), .QN(n363) );
  DFFRX1 \i_MIPS/Register/register_reg[29][21]  ( .D(\i_MIPS/Register/n201 ), 
        .CK(clk), .RN(n4075), .Q(\i_MIPS/Register/register[29][21] ), .QN(n303) );
  DFFRX1 \i_MIPS/Register/register_reg[29][22]  ( .D(\i_MIPS/Register/n202 ), 
        .CK(clk), .RN(n4075), .Q(\i_MIPS/Register/register[29][22] ), .QN(n353) );
  DFFRX1 \i_MIPS/Register/register_reg[29][23]  ( .D(\i_MIPS/Register/n203 ), 
        .CK(clk), .RN(n4075), .Q(\i_MIPS/Register/register[29][23] ), .QN(n358) );
  DFFRX1 \i_MIPS/Register/register_reg[29][24]  ( .D(\i_MIPS/Register/n204 ), 
        .CK(clk), .RN(n4076), .Q(\i_MIPS/Register/register[29][24] ), .QN(n308) );
  DFFRX1 \i_MIPS/Register/register_reg[29][25]  ( .D(\i_MIPS/Register/n205 ), 
        .CK(clk), .RN(n4076), .Q(\i_MIPS/Register/register[29][25] ), .QN(n293) );
  DFFRX1 \i_MIPS/Register/register_reg[29][26]  ( .D(\i_MIPS/Register/n206 ), 
        .CK(clk), .RN(n4076), .Q(\i_MIPS/Register/register[29][26] ), .QN(n313) );
  DFFRX1 \i_MIPS/Register/register_reg[29][27]  ( .D(\i_MIPS/Register/n207 ), 
        .CK(clk), .RN(n4076), .Q(\i_MIPS/Register/register[29][27] ), .QN(n328) );
  DFFRX1 \i_MIPS/Register/register_reg[29][28]  ( .D(\i_MIPS/Register/n208 ), 
        .CK(clk), .RN(n4076), .Q(\i_MIPS/Register/register[29][28] ), .QN(n338) );
  DFFRX1 \i_MIPS/Register/register_reg[29][29]  ( .D(\i_MIPS/Register/n209 ), 
        .CK(clk), .RN(n4076), .Q(\i_MIPS/Register/register[29][29] ), .QN(n333) );
  DFFRX1 \i_MIPS/Register/register_reg[29][30]  ( .D(\i_MIPS/Register/n210 ), 
        .CK(clk), .RN(n4076), .Q(\i_MIPS/Register/register[29][30] ), .QN(n348) );
  DFFRX1 \i_MIPS/Register/register_reg[29][31]  ( .D(\i_MIPS/Register/n211 ), 
        .CK(clk), .RN(n4076), .Q(\i_MIPS/Register/register[29][31] ), .QN(n343) );
  DFFRX1 \i_MIPS/Register/register_reg[27][2]  ( .D(\i_MIPS/Register/n246 ), 
        .CK(clk), .RN(n4079), .Q(\i_MIPS/Register/register[27][2] ), .QN(n282)
         );
  DFFRX1 \i_MIPS/Register/register_reg[27][3]  ( .D(\i_MIPS/Register/n247 ), 
        .CK(clk), .RN(n4079), .Q(\i_MIPS/Register/register[27][3] ), .QN(n287)
         );
  DFFRX1 \i_MIPS/Register/register_reg[27][4]  ( .D(\i_MIPS/Register/n248 ), 
        .CK(clk), .RN(n4079), .Q(\i_MIPS/Register/register[27][4] ), .QN(n244)
         );
  DFFRX1 \i_MIPS/Register/register_reg[27][5]  ( .D(\i_MIPS/Register/n249 ), 
        .CK(clk), .RN(n4079), .Q(\i_MIPS/Register/register[27][5] ), .QN(n257)
         );
  DFFRX1 \i_MIPS/Register/register_reg[27][6]  ( .D(\i_MIPS/Register/n250 ), 
        .CK(clk), .RN(n4079), .Q(\i_MIPS/Register/register[27][6] ), .QN(n267)
         );
  DFFRX1 \i_MIPS/Register/register_reg[27][7]  ( .D(\i_MIPS/Register/n251 ), 
        .CK(clk), .RN(n4079), .Q(\i_MIPS/Register/register[27][7] ), .QN(n262)
         );
  DFFRX1 \i_MIPS/Register/register_reg[27][10]  ( .D(\i_MIPS/Register/n254 ), 
        .CK(clk), .RN(n4080), .Q(\i_MIPS/Register/register[27][10] ), .QN(n252) );
  DFFRX1 \i_MIPS/Register/register_reg[27][11]  ( .D(\i_MIPS/Register/n255 ), 
        .CK(clk), .RN(n4080), .Q(\i_MIPS/Register/register[27][11] ), .QN(n249) );
  DFFRX1 \i_MIPS/Register/register_reg[27][12]  ( .D(\i_MIPS/Register/n256 ), 
        .CK(clk), .RN(n4080), .Q(\i_MIPS/Register/register[27][12] ), .QN(n229) );
  DFFRX1 \i_MIPS/Register/register_reg[27][13]  ( .D(\i_MIPS/Register/n257 ), 
        .CK(clk), .RN(n4080), .Q(\i_MIPS/Register/register[27][13] ), .QN(n214) );
  DFFRX1 \i_MIPS/Register/register_reg[27][15]  ( .D(\i_MIPS/Register/n259 ), 
        .CK(clk), .RN(n4080), .Q(\i_MIPS/Register/register[27][15] ), .QN(n297) );
  DFFRX1 \i_MIPS/Register/register_reg[27][16]  ( .D(\i_MIPS/Register/n260 ), 
        .CK(clk), .RN(n4080), .Q(\i_MIPS/Register/register[27][16] ), .QN(n317) );
  DFFRX1 \i_MIPS/Register/register_reg[27][17]  ( .D(\i_MIPS/Register/n261 ), 
        .CK(clk), .RN(n4080), .Q(\i_MIPS/Register/register[27][17] ), .QN(n372) );
  DFFRX1 \i_MIPS/Register/register_reg[27][18]  ( .D(\i_MIPS/Register/n262 ), 
        .CK(clk), .RN(n4080), .Q(\i_MIPS/Register/register[27][18] ), .QN(n367) );
  DFFRX1 \i_MIPS/Register/register_reg[27][19]  ( .D(\i_MIPS/Register/n263 ), 
        .CK(clk), .RN(n4080), .Q(\i_MIPS/Register/register[27][19] ), .QN(n322) );
  DFFRX1 \i_MIPS/Register/register_reg[27][20]  ( .D(\i_MIPS/Register/n264 ), 
        .CK(clk), .RN(n4081), .Q(\i_MIPS/Register/register[27][20] ), .QN(n362) );
  DFFRX1 \i_MIPS/Register/register_reg[27][21]  ( .D(\i_MIPS/Register/n265 ), 
        .CK(clk), .RN(n4081), .Q(\i_MIPS/Register/register[27][21] ), .QN(n302) );
  DFFRX1 \i_MIPS/Register/register_reg[27][22]  ( .D(\i_MIPS/Register/n266 ), 
        .CK(clk), .RN(n4081), .Q(\i_MIPS/Register/register[27][22] ), .QN(n352) );
  DFFRX1 \i_MIPS/Register/register_reg[27][23]  ( .D(\i_MIPS/Register/n267 ), 
        .CK(clk), .RN(n4081), .Q(\i_MIPS/Register/register[27][23] ), .QN(n357) );
  DFFRX1 \i_MIPS/Register/register_reg[27][24]  ( .D(\i_MIPS/Register/n268 ), 
        .CK(clk), .RN(n4081), .Q(\i_MIPS/Register/register[27][24] ), .QN(n307) );
  DFFRX1 \i_MIPS/Register/register_reg[27][25]  ( .D(\i_MIPS/Register/n269 ), 
        .CK(clk), .RN(n4081), .Q(\i_MIPS/Register/register[27][25] ), .QN(n292) );
  DFFRX1 \i_MIPS/Register/register_reg[27][26]  ( .D(\i_MIPS/Register/n270 ), 
        .CK(clk), .RN(n4081), .Q(\i_MIPS/Register/register[27][26] ), .QN(n312) );
  DFFRX1 \i_MIPS/Register/register_reg[27][27]  ( .D(\i_MIPS/Register/n271 ), 
        .CK(clk), .RN(n4081), .Q(\i_MIPS/Register/register[27][27] ), .QN(n327) );
  DFFRX1 \i_MIPS/Register/register_reg[27][28]  ( .D(\i_MIPS/Register/n272 ), 
        .CK(clk), .RN(n4081), .Q(\i_MIPS/Register/register[27][28] ), .QN(n337) );
  DFFRX1 \i_MIPS/Register/register_reg[27][29]  ( .D(\i_MIPS/Register/n273 ), 
        .CK(clk), .RN(n4081), .Q(\i_MIPS/Register/register[27][29] ), .QN(n332) );
  DFFRX1 \i_MIPS/Register/register_reg[27][30]  ( .D(\i_MIPS/Register/n274 ), 
        .CK(clk), .RN(n4081), .Q(\i_MIPS/Register/register[27][30] ), .QN(n347) );
  DFFRX1 \i_MIPS/Register/register_reg[27][31]  ( .D(\i_MIPS/Register/n275 ), 
        .CK(clk), .RN(n4081), .Q(\i_MIPS/Register/register[27][31] ), .QN(n342) );
  DFFRX1 \i_MIPS/Register/register_reg[25][2]  ( .D(\i_MIPS/Register/n310 ), 
        .CK(clk), .RN(n4084), .Q(\i_MIPS/Register/register[25][2] ), .QN(n396)
         );
  DFFRX1 \i_MIPS/Register/register_reg[25][3]  ( .D(\i_MIPS/Register/n311 ), 
        .CK(clk), .RN(n4084), .Q(\i_MIPS/Register/register[25][3] ), .QN(n398)
         );
  DFFRX1 \i_MIPS/Register/register_reg[25][4]  ( .D(\i_MIPS/Register/n312 ), 
        .CK(clk), .RN(n4085), .Q(\i_MIPS/Register/register[25][4] ), .QN(n383)
         );
  DFFRX1 \i_MIPS/Register/register_reg[25][11]  ( .D(\i_MIPS/Register/n319 ), 
        .CK(clk), .RN(n4085), .Q(\i_MIPS/Register/register[25][11] ), .QN(
        n1111) );
  DFFRX1 \i_MIPS/Register/register_reg[25][13]  ( .D(\i_MIPS/Register/n321 ), 
        .CK(clk), .RN(n4085), .Q(\i_MIPS/Register/register[25][13] ), .QN(n220) );
  DFFRX1 \i_MIPS/Register/register_reg[25][15]  ( .D(\i_MIPS/Register/n323 ), 
        .CK(clk), .RN(n4085), .Q(\i_MIPS/Register/register[25][15] ), .QN(n402) );
  DFFRX1 \i_MIPS/Register/register_reg[25][16]  ( .D(\i_MIPS/Register/n324 ), 
        .CK(clk), .RN(n4086), .Q(\i_MIPS/Register/register[25][16] ), .QN(n410) );
  DFFRX1 \i_MIPS/Register/register_reg[25][17]  ( .D(\i_MIPS/Register/n325 ), 
        .CK(clk), .RN(n4086), .Q(\i_MIPS/Register/register[25][17] ), .QN(n432) );
  DFFRX1 \i_MIPS/Register/register_reg[25][18]  ( .D(\i_MIPS/Register/n326 ), 
        .CK(clk), .RN(n4086), .Q(\i_MIPS/Register/register[25][18] ), .QN(n430) );
  DFFRX1 \i_MIPS/Register/register_reg[25][19]  ( .D(\i_MIPS/Register/n327 ), 
        .CK(clk), .RN(n4086), .Q(\i_MIPS/Register/register[25][19] ), .QN(n412) );
  DFFRX1 \i_MIPS/Register/register_reg[25][20]  ( .D(\i_MIPS/Register/n328 ), 
        .CK(clk), .RN(n4086), .Q(\i_MIPS/Register/register[25][20] ), .QN(n428) );
  DFFRX1 \i_MIPS/Register/register_reg[25][21]  ( .D(\i_MIPS/Register/n329 ), 
        .CK(clk), .RN(n4086), .Q(\i_MIPS/Register/register[25][21] ), .QN(n404) );
  DFFRX1 \i_MIPS/Register/register_reg[25][22]  ( .D(\i_MIPS/Register/n330 ), 
        .CK(clk), .RN(n4086), .Q(\i_MIPS/Register/register[25][22] ), .QN(n424) );
  DFFRX1 \i_MIPS/Register/register_reg[25][23]  ( .D(\i_MIPS/Register/n331 ), 
        .CK(clk), .RN(n4086), .Q(\i_MIPS/Register/register[25][23] ), .QN(n426) );
  DFFRX1 \i_MIPS/Register/register_reg[25][24]  ( .D(\i_MIPS/Register/n332 ), 
        .CK(clk), .RN(n4086), .Q(\i_MIPS/Register/register[25][24] ), .QN(n406) );
  DFFRX1 \i_MIPS/Register/register_reg[25][25]  ( .D(\i_MIPS/Register/n333 ), 
        .CK(clk), .RN(n4086), .Q(\i_MIPS/Register/register[25][25] ), .QN(n400) );
  DFFRX1 \i_MIPS/Register/register_reg[25][26]  ( .D(\i_MIPS/Register/n334 ), 
        .CK(clk), .RN(n4086), .Q(\i_MIPS/Register/register[25][26] ), .QN(n408) );
  DFFRX1 \i_MIPS/Register/register_reg[25][27]  ( .D(\i_MIPS/Register/n335 ), 
        .CK(clk), .RN(n4086), .Q(\i_MIPS/Register/register[25][27] ), .QN(n414) );
  DFFRX1 \i_MIPS/Register/register_reg[25][28]  ( .D(\i_MIPS/Register/n336 ), 
        .CK(clk), .RN(n4087), .Q(\i_MIPS/Register/register[25][28] ), .QN(n418) );
  DFFRX1 \i_MIPS/Register/register_reg[25][29]  ( .D(\i_MIPS/Register/n337 ), 
        .CK(clk), .RN(n4087), .Q(\i_MIPS/Register/register[25][29] ), .QN(n416) );
  DFFRX1 \i_MIPS/Register/register_reg[25][30]  ( .D(\i_MIPS/Register/n338 ), 
        .CK(clk), .RN(n4087), .Q(\i_MIPS/Register/register[25][30] ), .QN(n422) );
  DFFRX1 \i_MIPS/Register/register_reg[25][31]  ( .D(\i_MIPS/Register/n339 ), 
        .CK(clk), .RN(n4087), .Q(\i_MIPS/Register/register[25][31] ), .QN(n420) );
  DFFRX1 \i_MIPS/Register/register_reg[23][2]  ( .D(\i_MIPS/Register/n374 ), 
        .CK(clk), .RN(n4090), .Q(\i_MIPS/Register/register[23][2] ), .QN(n1177) );
  DFFRX1 \i_MIPS/Register/register_reg[23][3]  ( .D(\i_MIPS/Register/n375 ), 
        .CK(clk), .RN(n4090), .Q(\i_MIPS/Register/register[23][3] ), .QN(n1183) );
  DFFRX1 \i_MIPS/Register/register_reg[23][4]  ( .D(\i_MIPS/Register/n376 ), 
        .CK(clk), .RN(n4090), .Q(\i_MIPS/Register/register[23][4] ), .QN(n1131) );
  DFFRX1 \i_MIPS/Register/register_reg[23][5]  ( .D(\i_MIPS/Register/n377 ), 
        .CK(clk), .RN(n4090), .Q(\i_MIPS/Register/register[23][5] ), .QN(n1147) );
  DFFRX1 \i_MIPS/Register/register_reg[23][6]  ( .D(\i_MIPS/Register/n378 ), 
        .CK(clk), .RN(n4090), .Q(\i_MIPS/Register/register[23][6] ), .QN(n1159) );
  DFFRX1 \i_MIPS/Register/register_reg[23][7]  ( .D(\i_MIPS/Register/n379 ), 
        .CK(clk), .RN(n4090), .Q(\i_MIPS/Register/register[23][7] ), .QN(n1153) );
  DFFRX1 \i_MIPS/Register/register_reg[23][9]  ( .D(\i_MIPS/Register/n381 ), 
        .CK(clk), .RN(n4090), .Q(\i_MIPS/Register/register[23][9] ), .QN(n1119) );
  DFFRX1 \i_MIPS/Register/register_reg[23][10]  ( .D(\i_MIPS/Register/n382 ), 
        .CK(clk), .RN(n4090), .Q(\i_MIPS/Register/register[23][10] ), .QN(
        n1141) );
  DFFRX1 \i_MIPS/Register/register_reg[23][11]  ( .D(\i_MIPS/Register/n383 ), 
        .CK(clk), .RN(n4090), .Q(\i_MIPS/Register/register[23][11] ), .QN(
        n1137) );
  DFFRX1 \i_MIPS/Register/register_reg[23][12]  ( .D(\i_MIPS/Register/n384 ), 
        .CK(clk), .RN(n4091), .Q(\i_MIPS/Register/register[23][12] ), .QN(
        n1113) );
  DFFRX1 \i_MIPS/Register/register_reg[23][13]  ( .D(\i_MIPS/Register/n385 ), 
        .CK(clk), .RN(n4091), .Q(\i_MIPS/Register/register[23][13] ), .QN(
        n1098) );
  DFFRX1 \i_MIPS/Register/register_reg[23][14]  ( .D(\i_MIPS/Register/n386 ), 
        .CK(clk), .RN(n4091), .Q(\i_MIPS/Register/register[23][14] ), .QN(
        n1125) );
  DFFRX1 \i_MIPS/Register/register_reg[23][15]  ( .D(\i_MIPS/Register/n387 ), 
        .CK(clk), .RN(n4091), .Q(\i_MIPS/Register/register[23][15] ), .QN(
        n1195) );
  DFFRX1 \i_MIPS/Register/register_reg[23][16]  ( .D(\i_MIPS/Register/n388 ), 
        .CK(clk), .RN(n4091), .Q(\i_MIPS/Register/register[23][16] ), .QN(
        n1219) );
  DFFRX1 \i_MIPS/Register/register_reg[23][17]  ( .D(\i_MIPS/Register/n389 ), 
        .CK(clk), .RN(n4091), .Q(\i_MIPS/Register/register[23][17] ), .QN(
        n1285) );
  DFFRX1 \i_MIPS/Register/register_reg[23][18]  ( .D(\i_MIPS/Register/n390 ), 
        .CK(clk), .RN(n4091), .Q(\i_MIPS/Register/register[23][18] ), .QN(
        n1279) );
  DFFRX1 \i_MIPS/Register/register_reg[23][19]  ( .D(\i_MIPS/Register/n391 ), 
        .CK(clk), .RN(n4091), .Q(\i_MIPS/Register/register[23][19] ), .QN(
        n1225) );
  DFFRX1 \i_MIPS/Register/register_reg[23][20]  ( .D(\i_MIPS/Register/n392 ), 
        .CK(clk), .RN(n4091), .Q(\i_MIPS/Register/register[23][20] ), .QN(
        n1273) );
  DFFRX1 \i_MIPS/Register/register_reg[23][21]  ( .D(\i_MIPS/Register/n393 ), 
        .CK(clk), .RN(n4091), .Q(\i_MIPS/Register/register[23][21] ), .QN(
        n1201) );
  DFFRX1 \i_MIPS/Register/register_reg[23][22]  ( .D(\i_MIPS/Register/n394 ), 
        .CK(clk), .RN(n4091), .Q(\i_MIPS/Register/register[23][22] ), .QN(
        n1261) );
  DFFRX1 \i_MIPS/Register/register_reg[23][23]  ( .D(\i_MIPS/Register/n395 ), 
        .CK(clk), .RN(n4091), .Q(\i_MIPS/Register/register[23][23] ), .QN(
        n1267) );
  DFFRX1 \i_MIPS/Register/register_reg[23][24]  ( .D(\i_MIPS/Register/n396 ), 
        .CK(clk), .RN(n4092), .Q(\i_MIPS/Register/register[23][24] ), .QN(
        n1207) );
  DFFRX1 \i_MIPS/Register/register_reg[23][25]  ( .D(\i_MIPS/Register/n397 ), 
        .CK(clk), .RN(n4092), .Q(\i_MIPS/Register/register[23][25] ), .QN(
        n1189) );
  DFFRX1 \i_MIPS/Register/register_reg[23][26]  ( .D(\i_MIPS/Register/n398 ), 
        .CK(clk), .RN(n4092), .Q(\i_MIPS/Register/register[23][26] ), .QN(
        n1213) );
  DFFRX1 \i_MIPS/Register/register_reg[23][27]  ( .D(\i_MIPS/Register/n399 ), 
        .CK(clk), .RN(n4092), .Q(\i_MIPS/Register/register[23][27] ), .QN(
        n1231) );
  DFFRX1 \i_MIPS/Register/register_reg[23][28]  ( .D(\i_MIPS/Register/n400 ), 
        .CK(clk), .RN(n4092), .Q(\i_MIPS/Register/register[23][28] ), .QN(
        n1243) );
  DFFRX1 \i_MIPS/Register/register_reg[23][29]  ( .D(\i_MIPS/Register/n401 ), 
        .CK(clk), .RN(n4092), .Q(\i_MIPS/Register/register[23][29] ), .QN(
        n1237) );
  DFFRX1 \i_MIPS/Register/register_reg[23][30]  ( .D(\i_MIPS/Register/n402 ), 
        .CK(clk), .RN(n4092), .Q(\i_MIPS/Register/register[23][30] ), .QN(
        n1255) );
  DFFRX1 \i_MIPS/Register/register_reg[23][31]  ( .D(\i_MIPS/Register/n403 ), 
        .CK(clk), .RN(n4092), .Q(\i_MIPS/Register/register[23][31] ), .QN(
        n1249) );
  DFFRX1 \i_MIPS/Register/register_reg[21][2]  ( .D(\i_MIPS/Register/n438 ), 
        .CK(clk), .RN(n4095), .Q(\i_MIPS/Register/register[21][2] ), .QN(n1179) );
  DFFRX1 \i_MIPS/Register/register_reg[21][3]  ( .D(\i_MIPS/Register/n439 ), 
        .CK(clk), .RN(n4095), .Q(\i_MIPS/Register/register[21][3] ), .QN(n1185) );
  DFFRX1 \i_MIPS/Register/register_reg[21][4]  ( .D(\i_MIPS/Register/n440 ), 
        .CK(clk), .RN(n4095), .Q(\i_MIPS/Register/register[21][4] ), .QN(n1133) );
  DFFRX1 \i_MIPS/Register/register_reg[21][15]  ( .D(\i_MIPS/Register/n451 ), 
        .CK(clk), .RN(n4096), .Q(\i_MIPS/Register/register[21][15] ), .QN(
        n1197) );
  DFFRX1 \i_MIPS/Register/register_reg[21][16]  ( .D(\i_MIPS/Register/n452 ), 
        .CK(clk), .RN(n4096), .Q(\i_MIPS/Register/register[21][16] ), .QN(
        n1221) );
  DFFRX1 \i_MIPS/Register/register_reg[21][17]  ( .D(\i_MIPS/Register/n453 ), 
        .CK(clk), .RN(n4096), .Q(\i_MIPS/Register/register[21][17] ), .QN(
        n1287) );
  DFFRX1 \i_MIPS/Register/register_reg[21][18]  ( .D(\i_MIPS/Register/n454 ), 
        .CK(clk), .RN(n4096), .Q(\i_MIPS/Register/register[21][18] ), .QN(
        n1281) );
  DFFRX1 \i_MIPS/Register/register_reg[21][19]  ( .D(\i_MIPS/Register/n455 ), 
        .CK(clk), .RN(n4096), .Q(\i_MIPS/Register/register[21][19] ), .QN(
        n1227) );
  DFFRX1 \i_MIPS/Register/register_reg[21][20]  ( .D(\i_MIPS/Register/n456 ), 
        .CK(clk), .RN(n4097), .Q(\i_MIPS/Register/register[21][20] ), .QN(
        n1275) );
  DFFRX1 \i_MIPS/Register/register_reg[21][21]  ( .D(\i_MIPS/Register/n457 ), 
        .CK(clk), .RN(n4097), .Q(\i_MIPS/Register/register[21][21] ), .QN(
        n1203) );
  DFFRX1 \i_MIPS/Register/register_reg[21][22]  ( .D(\i_MIPS/Register/n458 ), 
        .CK(clk), .RN(n4097), .Q(\i_MIPS/Register/register[21][22] ), .QN(
        n1263) );
  DFFRX1 \i_MIPS/Register/register_reg[21][23]  ( .D(\i_MIPS/Register/n459 ), 
        .CK(clk), .RN(n4097), .Q(\i_MIPS/Register/register[21][23] ), .QN(
        n1269) );
  DFFRX1 \i_MIPS/Register/register_reg[21][24]  ( .D(\i_MIPS/Register/n460 ), 
        .CK(clk), .RN(n4097), .Q(\i_MIPS/Register/register[21][24] ), .QN(
        n1209) );
  DFFRX1 \i_MIPS/Register/register_reg[21][25]  ( .D(\i_MIPS/Register/n461 ), 
        .CK(clk), .RN(n4097), .Q(\i_MIPS/Register/register[21][25] ), .QN(
        n1191) );
  DFFRX1 \i_MIPS/Register/register_reg[21][26]  ( .D(\i_MIPS/Register/n462 ), 
        .CK(clk), .RN(n4097), .Q(\i_MIPS/Register/register[21][26] ), .QN(
        n1215) );
  DFFRX1 \i_MIPS/Register/register_reg[21][27]  ( .D(\i_MIPS/Register/n463 ), 
        .CK(clk), .RN(n4097), .Q(\i_MIPS/Register/register[21][27] ), .QN(
        n1233) );
  DFFRX1 \i_MIPS/Register/register_reg[21][28]  ( .D(\i_MIPS/Register/n464 ), 
        .CK(clk), .RN(n4097), .Q(\i_MIPS/Register/register[21][28] ), .QN(
        n1245) );
  DFFRX1 \i_MIPS/Register/register_reg[21][29]  ( .D(\i_MIPS/Register/n465 ), 
        .CK(clk), .RN(n4097), .Q(\i_MIPS/Register/register[21][29] ), .QN(
        n1239) );
  DFFRX1 \i_MIPS/Register/register_reg[21][30]  ( .D(\i_MIPS/Register/n466 ), 
        .CK(clk), .RN(n4097), .Q(\i_MIPS/Register/register[21][30] ), .QN(
        n1257) );
  DFFRX1 \i_MIPS/Register/register_reg[21][31]  ( .D(\i_MIPS/Register/n467 ), 
        .CK(clk), .RN(n4097), .Q(\i_MIPS/Register/register[21][31] ), .QN(
        n1251) );
  DFFRX1 \i_MIPS/Register/register_reg[19][2]  ( .D(\i_MIPS/Register/n502 ), 
        .CK(clk), .RN(n4100), .Q(\i_MIPS/Register/register[19][2] ), .QN(n1178) );
  DFFRX1 \i_MIPS/Register/register_reg[19][3]  ( .D(\i_MIPS/Register/n503 ), 
        .CK(clk), .RN(n4100), .Q(\i_MIPS/Register/register[19][3] ), .QN(n1184) );
  DFFRX1 \i_MIPS/Register/register_reg[19][4]  ( .D(\i_MIPS/Register/n504 ), 
        .CK(clk), .RN(n4101), .Q(\i_MIPS/Register/register[19][4] ), .QN(n1132) );
  DFFRX1 \i_MIPS/Register/register_reg[19][7]  ( .D(\i_MIPS/Register/n507 ), 
        .CK(clk), .RN(n4101), .Q(\i_MIPS/Register/register[19][7] ), .QN(n1154) );
  DFFRX1 \i_MIPS/Register/register_reg[19][11]  ( .D(\i_MIPS/Register/n511 ), 
        .CK(clk), .RN(n4101), .Q(\i_MIPS/Register/register[19][11] ), .QN(
        n1138) );
  DFFRX1 \i_MIPS/Register/register_reg[19][12]  ( .D(\i_MIPS/Register/n512 ), 
        .CK(clk), .RN(n4101), .Q(\i_MIPS/Register/register[19][12] ), .QN(
        n1114) );
  DFFRX1 \i_MIPS/Register/register_reg[19][13]  ( .D(\i_MIPS/Register/n513 ), 
        .CK(clk), .RN(n4101), .Q(\i_MIPS/Register/register[19][13] ), .QN(
        n1099) );
  DFFRX1 \i_MIPS/Register/register_reg[19][15]  ( .D(\i_MIPS/Register/n515 ), 
        .CK(clk), .RN(n4101), .Q(\i_MIPS/Register/register[19][15] ), .QN(
        n1196) );
  DFFRX1 \i_MIPS/Register/register_reg[19][16]  ( .D(\i_MIPS/Register/n516 ), 
        .CK(clk), .RN(n4102), .Q(\i_MIPS/Register/register[19][16] ), .QN(
        n1220) );
  DFFRX1 \i_MIPS/Register/register_reg[19][17]  ( .D(\i_MIPS/Register/n517 ), 
        .CK(clk), .RN(n4102), .Q(\i_MIPS/Register/register[19][17] ), .QN(
        n1286) );
  DFFRX1 \i_MIPS/Register/register_reg[19][18]  ( .D(\i_MIPS/Register/n518 ), 
        .CK(clk), .RN(n4102), .Q(\i_MIPS/Register/register[19][18] ), .QN(
        n1280) );
  DFFRX1 \i_MIPS/Register/register_reg[19][19]  ( .D(\i_MIPS/Register/n519 ), 
        .CK(clk), .RN(n4102), .Q(\i_MIPS/Register/register[19][19] ), .QN(
        n1226) );
  DFFRX1 \i_MIPS/Register/register_reg[19][20]  ( .D(\i_MIPS/Register/n520 ), 
        .CK(clk), .RN(n4102), .Q(\i_MIPS/Register/register[19][20] ), .QN(
        n1274) );
  DFFRX1 \i_MIPS/Register/register_reg[19][21]  ( .D(\i_MIPS/Register/n521 ), 
        .CK(clk), .RN(n4102), .Q(\i_MIPS/Register/register[19][21] ), .QN(
        n1202) );
  DFFRX1 \i_MIPS/Register/register_reg[19][22]  ( .D(\i_MIPS/Register/n522 ), 
        .CK(clk), .RN(n4102), .Q(\i_MIPS/Register/register[19][22] ), .QN(
        n1262) );
  DFFRX1 \i_MIPS/Register/register_reg[19][23]  ( .D(\i_MIPS/Register/n523 ), 
        .CK(clk), .RN(n4102), .Q(\i_MIPS/Register/register[19][23] ), .QN(
        n1268) );
  DFFRX1 \i_MIPS/Register/register_reg[19][24]  ( .D(\i_MIPS/Register/n524 ), 
        .CK(clk), .RN(n4102), .Q(\i_MIPS/Register/register[19][24] ), .QN(
        n1208) );
  DFFRX1 \i_MIPS/Register/register_reg[19][25]  ( .D(\i_MIPS/Register/n525 ), 
        .CK(clk), .RN(n4102), .Q(\i_MIPS/Register/register[19][25] ), .QN(
        n1190) );
  DFFRX1 \i_MIPS/Register/register_reg[19][26]  ( .D(\i_MIPS/Register/n526 ), 
        .CK(clk), .RN(n4102), .Q(\i_MIPS/Register/register[19][26] ), .QN(
        n1214) );
  DFFRX1 \i_MIPS/Register/register_reg[19][27]  ( .D(\i_MIPS/Register/n527 ), 
        .CK(clk), .RN(n4102), .Q(\i_MIPS/Register/register[19][27] ), .QN(
        n1232) );
  DFFRX1 \i_MIPS/Register/register_reg[19][28]  ( .D(\i_MIPS/Register/n528 ), 
        .CK(clk), .RN(n4103), .Q(\i_MIPS/Register/register[19][28] ), .QN(
        n1244) );
  DFFRX1 \i_MIPS/Register/register_reg[19][29]  ( .D(\i_MIPS/Register/n529 ), 
        .CK(clk), .RN(n4103), .Q(\i_MIPS/Register/register[19][29] ), .QN(
        n1238) );
  DFFRX1 \i_MIPS/Register/register_reg[19][30]  ( .D(\i_MIPS/Register/n530 ), 
        .CK(clk), .RN(n4103), .Q(\i_MIPS/Register/register[19][30] ), .QN(
        n1256) );
  DFFRX1 \i_MIPS/Register/register_reg[19][31]  ( .D(\i_MIPS/Register/n531 ), 
        .CK(clk), .RN(n4103), .Q(\i_MIPS/Register/register[19][31] ), .QN(
        n1250) );
  DFFRX1 \i_MIPS/Register/register_reg[17][15]  ( .D(\i_MIPS/Register/n579 ), 
        .CK(clk), .RN(n4107), .Q(\i_MIPS/Register/register[17][15] ), .QN(
        n1316) );
  DFFRX1 \i_MIPS/Register/register_reg[17][16]  ( .D(\i_MIPS/Register/n580 ), 
        .CK(clk), .RN(n4107), .Q(\i_MIPS/Register/register[17][16] ), .QN(
        n1324) );
  DFFRX1 \i_MIPS/Register/register_reg[17][17]  ( .D(\i_MIPS/Register/n581 ), 
        .CK(clk), .RN(n4107), .Q(\i_MIPS/Register/register[17][17] ), .QN(
        n1346) );
  DFFRX1 \i_MIPS/Register/register_reg[17][18]  ( .D(\i_MIPS/Register/n582 ), 
        .CK(clk), .RN(n4107), .Q(\i_MIPS/Register/register[17][18] ), .QN(
        n1344) );
  DFFRX1 \i_MIPS/Register/register_reg[17][19]  ( .D(\i_MIPS/Register/n583 ), 
        .CK(clk), .RN(n4107), .Q(\i_MIPS/Register/register[17][19] ), .QN(
        n1326) );
  DFFRX1 \i_MIPS/Register/register_reg[17][20]  ( .D(\i_MIPS/Register/n584 ), 
        .CK(clk), .RN(n4107), .Q(\i_MIPS/Register/register[17][20] ), .QN(
        n1342) );
  DFFRX1 \i_MIPS/Register/register_reg[17][21]  ( .D(\i_MIPS/Register/n585 ), 
        .CK(clk), .RN(n4107), .Q(\i_MIPS/Register/register[17][21] ), .QN(
        n1318) );
  DFFRX1 \i_MIPS/Register/register_reg[17][22]  ( .D(\i_MIPS/Register/n586 ), 
        .CK(clk), .RN(n4107), .Q(\i_MIPS/Register/register[17][22] ), .QN(
        n1338) );
  DFFRX1 \i_MIPS/Register/register_reg[17][23]  ( .D(\i_MIPS/Register/n587 ), 
        .CK(clk), .RN(n4107), .Q(\i_MIPS/Register/register[17][23] ), .QN(
        n1340) );
  DFFRX1 \i_MIPS/Register/register_reg[17][24]  ( .D(\i_MIPS/Register/n588 ), 
        .CK(clk), .RN(n4108), .Q(\i_MIPS/Register/register[17][24] ), .QN(
        n1320) );
  DFFRX1 \i_MIPS/Register/register_reg[17][25]  ( .D(\i_MIPS/Register/n589 ), 
        .CK(clk), .RN(n4108), .Q(\i_MIPS/Register/register[17][25] ), .QN(
        n1314) );
  DFFRX1 \i_MIPS/Register/register_reg[17][26]  ( .D(\i_MIPS/Register/n590 ), 
        .CK(clk), .RN(n4108), .Q(\i_MIPS/Register/register[17][26] ), .QN(
        n1322) );
  DFFRX1 \i_MIPS/Register/register_reg[17][27]  ( .D(\i_MIPS/Register/n591 ), 
        .CK(clk), .RN(n4108), .Q(\i_MIPS/Register/register[17][27] ), .QN(
        n1328) );
  DFFRX1 \i_MIPS/Register/register_reg[17][28]  ( .D(\i_MIPS/Register/n592 ), 
        .CK(clk), .RN(n4108), .Q(\i_MIPS/Register/register[17][28] ), .QN(
        n1332) );
  DFFRX1 \i_MIPS/Register/register_reg[17][29]  ( .D(\i_MIPS/Register/n593 ), 
        .CK(clk), .RN(n4108), .Q(\i_MIPS/Register/register[17][29] ), .QN(
        n1330) );
  DFFRX1 \i_MIPS/Register/register_reg[17][30]  ( .D(\i_MIPS/Register/n594 ), 
        .CK(clk), .RN(n4108), .Q(\i_MIPS/Register/register[17][30] ), .QN(
        n1336) );
  DFFRX1 \i_MIPS/Register/register_reg[17][31]  ( .D(\i_MIPS/Register/n595 ), 
        .CK(clk), .RN(n4108), .Q(\i_MIPS/Register/register[17][31] ), .QN(
        n1334) );
  DFFRX1 \i_MIPS/Register/register_reg[15][2]  ( .D(\i_MIPS/Register/n630 ), 
        .CK(clk), .RN(n4111), .Q(\i_MIPS/Register/register[15][2] ), .QN(n284)
         );
  DFFRX1 \i_MIPS/Register/register_reg[15][3]  ( .D(\i_MIPS/Register/n631 ), 
        .CK(clk), .RN(n4111), .Q(\i_MIPS/Register/register[15][3] ), .QN(n289)
         );
  DFFRX1 \i_MIPS/Register/register_reg[15][4]  ( .D(\i_MIPS/Register/n632 ), 
        .CK(clk), .RN(n4111), .Q(\i_MIPS/Register/register[15][4] ), .QN(n246)
         );
  DFFRX1 \i_MIPS/Register/register_reg[15][5]  ( .D(\i_MIPS/Register/n633 ), 
        .CK(clk), .RN(n4111), .Q(\i_MIPS/Register/register[15][5] ), .QN(n259)
         );
  DFFRX1 \i_MIPS/Register/register_reg[15][6]  ( .D(\i_MIPS/Register/n634 ), 
        .CK(clk), .RN(n4111), .Q(\i_MIPS/Register/register[15][6] ), .QN(n269)
         );
  DFFRX1 \i_MIPS/Register/register_reg[15][7]  ( .D(\i_MIPS/Register/n635 ), 
        .CK(clk), .RN(n4111), .Q(\i_MIPS/Register/register[15][7] ), .QN(n264)
         );
  DFFRX1 \i_MIPS/Register/register_reg[15][8]  ( .D(\i_MIPS/Register/n636 ), 
        .CK(clk), .RN(n4112), .Q(\i_MIPS/Register/register[15][8] ), .QN(n1107) );
  DFFRX1 \i_MIPS/Register/register_reg[15][9]  ( .D(\i_MIPS/Register/n637 ), 
        .CK(clk), .RN(n4112), .Q(\i_MIPS/Register/register[15][9] ), .QN(n236)
         );
  DFFRX1 \i_MIPS/Register/register_reg[15][10]  ( .D(\i_MIPS/Register/n638 ), 
        .CK(clk), .RN(n4112), .Q(\i_MIPS/Register/register[15][10] ), .QN(n254) );
  DFFRX1 \i_MIPS/Register/register_reg[15][11]  ( .D(\i_MIPS/Register/n639 ), 
        .CK(clk), .RN(n4112), .Q(\i_MIPS/Register/register[15][11] ), .QN(n250) );
  DFFRX1 \i_MIPS/Register/register_reg[15][12]  ( .D(\i_MIPS/Register/n640 ), 
        .CK(clk), .RN(n4112), .Q(\i_MIPS/Register/register[15][12] ), .QN(n231) );
  DFFRX1 \i_MIPS/Register/register_reg[15][13]  ( .D(\i_MIPS/Register/n641 ), 
        .CK(clk), .RN(n4112), .Q(\i_MIPS/Register/register[15][13] ), .QN(
        n1108) );
  DFFRX1 \i_MIPS/Register/register_reg[15][14]  ( .D(\i_MIPS/Register/n642 ), 
        .CK(clk), .RN(n4112), .Q(\i_MIPS/Register/register[15][14] ), .QN(n241) );
  DFFRX1 \i_MIPS/Register/register_reg[15][15]  ( .D(\i_MIPS/Register/n643 ), 
        .CK(clk), .RN(n4112), .Q(\i_MIPS/Register/register[15][15] ), .QN(n299) );
  DFFRX1 \i_MIPS/Register/register_reg[15][16]  ( .D(\i_MIPS/Register/n644 ), 
        .CK(clk), .RN(n4112), .Q(\i_MIPS/Register/register[15][16] ), .QN(n319) );
  DFFRX1 \i_MIPS/Register/register_reg[15][17]  ( .D(\i_MIPS/Register/n645 ), 
        .CK(clk), .RN(n4112), .Q(\i_MIPS/Register/register[15][17] ), .QN(n374) );
  DFFRX1 \i_MIPS/Register/register_reg[15][18]  ( .D(\i_MIPS/Register/n646 ), 
        .CK(clk), .RN(n4112), .Q(\i_MIPS/Register/register[15][18] ), .QN(n369) );
  DFFRX1 \i_MIPS/Register/register_reg[15][19]  ( .D(\i_MIPS/Register/n647 ), 
        .CK(clk), .RN(n4112), .Q(\i_MIPS/Register/register[15][19] ), .QN(n324) );
  DFFRX1 \i_MIPS/Register/register_reg[15][20]  ( .D(\i_MIPS/Register/n648 ), 
        .CK(clk), .RN(n4113), .Q(\i_MIPS/Register/register[15][20] ), .QN(n364) );
  DFFRX1 \i_MIPS/Register/register_reg[15][21]  ( .D(\i_MIPS/Register/n649 ), 
        .CK(clk), .RN(n4113), .Q(\i_MIPS/Register/register[15][21] ), .QN(n304) );
  DFFRX1 \i_MIPS/Register/register_reg[15][22]  ( .D(\i_MIPS/Register/n650 ), 
        .CK(clk), .RN(n4113), .Q(\i_MIPS/Register/register[15][22] ), .QN(n354) );
  DFFRX1 \i_MIPS/Register/register_reg[15][23]  ( .D(\i_MIPS/Register/n651 ), 
        .CK(clk), .RN(n4113), .Q(\i_MIPS/Register/register[15][23] ), .QN(n359) );
  DFFRX1 \i_MIPS/Register/register_reg[15][24]  ( .D(\i_MIPS/Register/n652 ), 
        .CK(clk), .RN(n4113), .Q(\i_MIPS/Register/register[15][24] ), .QN(n309) );
  DFFRX1 \i_MIPS/Register/register_reg[15][25]  ( .D(\i_MIPS/Register/n653 ), 
        .CK(clk), .RN(n4113), .Q(\i_MIPS/Register/register[15][25] ), .QN(n294) );
  DFFRX1 \i_MIPS/Register/register_reg[15][26]  ( .D(\i_MIPS/Register/n654 ), 
        .CK(clk), .RN(n4113), .Q(\i_MIPS/Register/register[15][26] ), .QN(n314) );
  DFFRX1 \i_MIPS/Register/register_reg[15][27]  ( .D(\i_MIPS/Register/n655 ), 
        .CK(clk), .RN(n4113), .Q(\i_MIPS/Register/register[15][27] ), .QN(n329) );
  DFFRX1 \i_MIPS/Register/register_reg[15][28]  ( .D(\i_MIPS/Register/n656 ), 
        .CK(clk), .RN(n4113), .Q(\i_MIPS/Register/register[15][28] ), .QN(n339) );
  DFFRX1 \i_MIPS/Register/register_reg[15][29]  ( .D(\i_MIPS/Register/n657 ), 
        .CK(clk), .RN(n4113), .Q(\i_MIPS/Register/register[15][29] ), .QN(n334) );
  DFFRX1 \i_MIPS/Register/register_reg[15][30]  ( .D(\i_MIPS/Register/n658 ), 
        .CK(clk), .RN(n4113), .Q(\i_MIPS/Register/register[15][30] ), .QN(n349) );
  DFFRX1 \i_MIPS/Register/register_reg[15][31]  ( .D(\i_MIPS/Register/n659 ), 
        .CK(clk), .RN(n4113), .Q(\i_MIPS/Register/register[15][31] ), .QN(n344) );
  DFFRX1 \i_MIPS/Register/register_reg[13][2]  ( .D(\i_MIPS/Register/n694 ), 
        .CK(clk), .RN(n4116), .Q(\i_MIPS/Register/register[13][2] ), .QN(n286)
         );
  DFFRX1 \i_MIPS/Register/register_reg[13][3]  ( .D(\i_MIPS/Register/n695 ), 
        .CK(clk), .RN(n4116), .Q(\i_MIPS/Register/register[13][3] ), .QN(n291)
         );
  DFFRX1 \i_MIPS/Register/register_reg[13][4]  ( .D(\i_MIPS/Register/n696 ), 
        .CK(clk), .RN(n4117), .Q(\i_MIPS/Register/register[13][4] ), .QN(n248)
         );
  DFFRX1 \i_MIPS/Register/register_reg[13][7]  ( .D(\i_MIPS/Register/n699 ), 
        .CK(clk), .RN(n4117), .Q(\i_MIPS/Register/register[13][7] ), .QN(n266)
         );
  DFFRX1 \i_MIPS/Register/register_reg[13][11]  ( .D(\i_MIPS/Register/n703 ), 
        .CK(clk), .RN(n4117), .Q(\i_MIPS/Register/register[13][11] ), .QN(
        n1110) );
  DFFRX1 \i_MIPS/Register/register_reg[13][12]  ( .D(\i_MIPS/Register/n704 ), 
        .CK(clk), .RN(n4117), .Q(\i_MIPS/Register/register[13][12] ), .QN(n233) );
  DFFRX1 \i_MIPS/Register/register_reg[13][13]  ( .D(\i_MIPS/Register/n705 ), 
        .CK(clk), .RN(n4117), .Q(\i_MIPS/Register/register[13][13] ), .QN(n217) );
  DFFRX1 \i_MIPS/Register/register_reg[13][15]  ( .D(\i_MIPS/Register/n707 ), 
        .CK(clk), .RN(n4117), .Q(\i_MIPS/Register/register[13][15] ), .QN(n301) );
  DFFRX1 \i_MIPS/Register/register_reg[13][16]  ( .D(\i_MIPS/Register/n708 ), 
        .CK(clk), .RN(n4118), .Q(\i_MIPS/Register/register[13][16] ), .QN(n321) );
  DFFRX1 \i_MIPS/Register/register_reg[13][17]  ( .D(\i_MIPS/Register/n709 ), 
        .CK(clk), .RN(n4118), .Q(\i_MIPS/Register/register[13][17] ), .QN(n376) );
  DFFRX1 \i_MIPS/Register/register_reg[13][18]  ( .D(\i_MIPS/Register/n710 ), 
        .CK(clk), .RN(n4118), .Q(\i_MIPS/Register/register[13][18] ), .QN(n371) );
  DFFRX1 \i_MIPS/Register/register_reg[13][19]  ( .D(\i_MIPS/Register/n711 ), 
        .CK(clk), .RN(n4118), .Q(\i_MIPS/Register/register[13][19] ), .QN(n326) );
  DFFRX1 \i_MIPS/Register/register_reg[13][20]  ( .D(\i_MIPS/Register/n712 ), 
        .CK(clk), .RN(n4118), .Q(\i_MIPS/Register/register[13][20] ), .QN(n366) );
  DFFRX1 \i_MIPS/Register/register_reg[13][21]  ( .D(\i_MIPS/Register/n713 ), 
        .CK(clk), .RN(n4118), .Q(\i_MIPS/Register/register[13][21] ), .QN(n306) );
  DFFRX1 \i_MIPS/Register/register_reg[13][22]  ( .D(\i_MIPS/Register/n714 ), 
        .CK(clk), .RN(n4118), .Q(\i_MIPS/Register/register[13][22] ), .QN(n356) );
  DFFRX1 \i_MIPS/Register/register_reg[13][23]  ( .D(\i_MIPS/Register/n715 ), 
        .CK(clk), .RN(n4118), .Q(\i_MIPS/Register/register[13][23] ), .QN(n361) );
  DFFRX1 \i_MIPS/Register/register_reg[13][24]  ( .D(\i_MIPS/Register/n716 ), 
        .CK(clk), .RN(n4118), .Q(\i_MIPS/Register/register[13][24] ), .QN(n311) );
  DFFRX1 \i_MIPS/Register/register_reg[13][25]  ( .D(\i_MIPS/Register/n717 ), 
        .CK(clk), .RN(n4118), .Q(\i_MIPS/Register/register[13][25] ), .QN(n296) );
  DFFRX1 \i_MIPS/Register/register_reg[13][26]  ( .D(\i_MIPS/Register/n718 ), 
        .CK(clk), .RN(n4118), .Q(\i_MIPS/Register/register[13][26] ), .QN(n316) );
  DFFRX1 \i_MIPS/Register/register_reg[13][27]  ( .D(\i_MIPS/Register/n719 ), 
        .CK(clk), .RN(n4118), .Q(\i_MIPS/Register/register[13][27] ), .QN(n331) );
  DFFRX1 \i_MIPS/Register/register_reg[13][28]  ( .D(\i_MIPS/Register/n720 ), 
        .CK(clk), .RN(n4119), .Q(\i_MIPS/Register/register[13][28] ), .QN(n341) );
  DFFRX1 \i_MIPS/Register/register_reg[13][29]  ( .D(\i_MIPS/Register/n721 ), 
        .CK(clk), .RN(n4119), .Q(\i_MIPS/Register/register[13][29] ), .QN(n336) );
  DFFRX1 \i_MIPS/Register/register_reg[13][30]  ( .D(\i_MIPS/Register/n722 ), 
        .CK(clk), .RN(n4119), .Q(\i_MIPS/Register/register[13][30] ), .QN(n351) );
  DFFRX1 \i_MIPS/Register/register_reg[13][31]  ( .D(\i_MIPS/Register/n723 ), 
        .CK(clk), .RN(n4119), .Q(\i_MIPS/Register/register[13][31] ), .QN(n346) );
  DFFRX1 \i_MIPS/Register/register_reg[11][2]  ( .D(\i_MIPS/Register/n758 ), 
        .CK(clk), .RN(n4122), .Q(\i_MIPS/Register/register[11][2] ), .QN(n285)
         );
  DFFRX1 \i_MIPS/Register/register_reg[11][3]  ( .D(\i_MIPS/Register/n759 ), 
        .CK(clk), .RN(n4122), .Q(\i_MIPS/Register/register[11][3] ), .QN(n290)
         );
  DFFRX1 \i_MIPS/Register/register_reg[11][4]  ( .D(\i_MIPS/Register/n760 ), 
        .CK(clk), .RN(n4122), .Q(\i_MIPS/Register/register[11][4] ), .QN(n247)
         );
  DFFRX1 \i_MIPS/Register/register_reg[11][5]  ( .D(\i_MIPS/Register/n761 ), 
        .CK(clk), .RN(n4122), .Q(\i_MIPS/Register/register[11][5] ), .QN(n260)
         );
  DFFRX1 \i_MIPS/Register/register_reg[11][6]  ( .D(\i_MIPS/Register/n762 ), 
        .CK(clk), .RN(n4122), .Q(\i_MIPS/Register/register[11][6] ), .QN(n270)
         );
  DFFRX1 \i_MIPS/Register/register_reg[11][7]  ( .D(\i_MIPS/Register/n763 ), 
        .CK(clk), .RN(n4122), .Q(\i_MIPS/Register/register[11][7] ), .QN(n265)
         );
  DFFRX1 \i_MIPS/Register/register_reg[11][10]  ( .D(\i_MIPS/Register/n766 ), 
        .CK(clk), .RN(n4122), .Q(\i_MIPS/Register/register[11][10] ), .QN(n255) );
  DFFRX1 \i_MIPS/Register/register_reg[11][11]  ( .D(\i_MIPS/Register/n767 ), 
        .CK(clk), .RN(n4122), .Q(\i_MIPS/Register/register[11][11] ), .QN(n251) );
  DFFRX1 \i_MIPS/Register/register_reg[11][12]  ( .D(\i_MIPS/Register/n768 ), 
        .CK(clk), .RN(n4123), .Q(\i_MIPS/Register/register[11][12] ), .QN(n232) );
  DFFRX1 \i_MIPS/Register/register_reg[11][13]  ( .D(\i_MIPS/Register/n769 ), 
        .CK(clk), .RN(n4123), .Q(\i_MIPS/Register/register[11][13] ), .QN(n216) );
  DFFRX1 \i_MIPS/Register/register_reg[11][14]  ( .D(\i_MIPS/Register/n770 ), 
        .CK(clk), .RN(n4123), .Q(\i_MIPS/Register/register[11][14] ), .QN(n242) );
  DFFRX1 \i_MIPS/Register/register_reg[11][15]  ( .D(\i_MIPS/Register/n771 ), 
        .CK(clk), .RN(n4123), .Q(\i_MIPS/Register/register[11][15] ), .QN(n300) );
  DFFRX1 \i_MIPS/Register/register_reg[11][16]  ( .D(\i_MIPS/Register/n772 ), 
        .CK(clk), .RN(n4123), .Q(\i_MIPS/Register/register[11][16] ), .QN(n320) );
  DFFRX1 \i_MIPS/Register/register_reg[11][17]  ( .D(\i_MIPS/Register/n773 ), 
        .CK(clk), .RN(n4123), .Q(\i_MIPS/Register/register[11][17] ), .QN(n375) );
  DFFRX1 \i_MIPS/Register/register_reg[11][18]  ( .D(\i_MIPS/Register/n774 ), 
        .CK(clk), .RN(n4123), .Q(\i_MIPS/Register/register[11][18] ), .QN(n370) );
  DFFRX1 \i_MIPS/Register/register_reg[11][19]  ( .D(\i_MIPS/Register/n775 ), 
        .CK(clk), .RN(n4123), .Q(\i_MIPS/Register/register[11][19] ), .QN(n325) );
  DFFRX1 \i_MIPS/Register/register_reg[11][20]  ( .D(\i_MIPS/Register/n776 ), 
        .CK(clk), .RN(n4123), .Q(\i_MIPS/Register/register[11][20] ), .QN(n365) );
  DFFRX1 \i_MIPS/Register/register_reg[11][21]  ( .D(\i_MIPS/Register/n777 ), 
        .CK(clk), .RN(n4123), .Q(\i_MIPS/Register/register[11][21] ), .QN(n305) );
  DFFRX1 \i_MIPS/Register/register_reg[11][22]  ( .D(\i_MIPS/Register/n778 ), 
        .CK(clk), .RN(n4123), .Q(\i_MIPS/Register/register[11][22] ), .QN(n355) );
  DFFRX1 \i_MIPS/Register/register_reg[11][23]  ( .D(\i_MIPS/Register/n779 ), 
        .CK(clk), .RN(n4123), .Q(\i_MIPS/Register/register[11][23] ), .QN(n360) );
  DFFRX1 \i_MIPS/Register/register_reg[11][24]  ( .D(\i_MIPS/Register/n780 ), 
        .CK(clk), .RN(n4124), .Q(\i_MIPS/Register/register[11][24] ), .QN(n310) );
  DFFRX1 \i_MIPS/Register/register_reg[11][25]  ( .D(\i_MIPS/Register/n781 ), 
        .CK(clk), .RN(n4124), .Q(\i_MIPS/Register/register[11][25] ), .QN(n295) );
  DFFRX1 \i_MIPS/Register/register_reg[11][26]  ( .D(\i_MIPS/Register/n782 ), 
        .CK(clk), .RN(n4124), .Q(\i_MIPS/Register/register[11][26] ), .QN(n315) );
  DFFRX1 \i_MIPS/Register/register_reg[11][27]  ( .D(\i_MIPS/Register/n783 ), 
        .CK(clk), .RN(n4124), .Q(\i_MIPS/Register/register[11][27] ), .QN(n330) );
  DFFRX1 \i_MIPS/Register/register_reg[11][28]  ( .D(\i_MIPS/Register/n784 ), 
        .CK(clk), .RN(n4124), .Q(\i_MIPS/Register/register[11][28] ), .QN(n340) );
  DFFRX1 \i_MIPS/Register/register_reg[11][29]  ( .D(\i_MIPS/Register/n785 ), 
        .CK(clk), .RN(n4124), .Q(\i_MIPS/Register/register[11][29] ), .QN(n335) );
  DFFRX1 \i_MIPS/Register/register_reg[11][30]  ( .D(\i_MIPS/Register/n786 ), 
        .CK(clk), .RN(n4124), .Q(\i_MIPS/Register/register[11][30] ), .QN(n350) );
  DFFRX1 \i_MIPS/Register/register_reg[11][31]  ( .D(\i_MIPS/Register/n787 ), 
        .CK(clk), .RN(n4124), .Q(\i_MIPS/Register/register[11][31] ), .QN(n345) );
  DFFRX1 \i_MIPS/Register/register_reg[9][2]  ( .D(\i_MIPS/Register/n822 ), 
        .CK(clk), .RN(n4127), .Q(\i_MIPS/Register/register[9][2] ), .QN(n397)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][3]  ( .D(\i_MIPS/Register/n823 ), 
        .CK(clk), .RN(n4127), .Q(\i_MIPS/Register/register[9][3] ), .QN(n399)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][4]  ( .D(\i_MIPS/Register/n824 ), 
        .CK(clk), .RN(n4127), .Q(\i_MIPS/Register/register[9][4] ), .QN(n384)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][11]  ( .D(\i_MIPS/Register/n831 ), 
        .CK(clk), .RN(n4128), .Q(\i_MIPS/Register/register[9][11] ), .QN(n1112) );
  DFFRX1 \i_MIPS/Register/register_reg[9][13]  ( .D(\i_MIPS/Register/n833 ), 
        .CK(clk), .RN(n4128), .Q(\i_MIPS/Register/register[9][13] ), .QN(n221)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][15]  ( .D(\i_MIPS/Register/n835 ), 
        .CK(clk), .RN(n4128), .Q(\i_MIPS/Register/register[9][15] ), .QN(n403)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][16]  ( .D(\i_MIPS/Register/n836 ), 
        .CK(clk), .RN(n4128), .Q(\i_MIPS/Register/register[9][16] ), .QN(n411)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][17]  ( .D(\i_MIPS/Register/n837 ), 
        .CK(clk), .RN(n4128), .Q(\i_MIPS/Register/register[9][17] ), .QN(n433)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][18]  ( .D(\i_MIPS/Register/n838 ), 
        .CK(clk), .RN(n4128), .Q(\i_MIPS/Register/register[9][18] ), .QN(n431)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][19]  ( .D(\i_MIPS/Register/n839 ), 
        .CK(clk), .RN(n4128), .Q(\i_MIPS/Register/register[9][19] ), .QN(n413)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][20]  ( .D(\i_MIPS/Register/n840 ), 
        .CK(clk), .RN(n4129), .Q(\i_MIPS/Register/register[9][20] ), .QN(n429)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][21]  ( .D(\i_MIPS/Register/n841 ), 
        .CK(clk), .RN(n4129), .Q(\i_MIPS/Register/register[9][21] ), .QN(n405)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][22]  ( .D(\i_MIPS/Register/n842 ), 
        .CK(clk), .RN(n4129), .Q(\i_MIPS/Register/register[9][22] ), .QN(n425)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][23]  ( .D(\i_MIPS/Register/n843 ), 
        .CK(clk), .RN(n4129), .Q(\i_MIPS/Register/register[9][23] ), .QN(n427)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][24]  ( .D(\i_MIPS/Register/n844 ), 
        .CK(clk), .RN(n4129), .Q(\i_MIPS/Register/register[9][24] ), .QN(n407)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][25]  ( .D(\i_MIPS/Register/n845 ), 
        .CK(clk), .RN(n4129), .Q(\i_MIPS/Register/register[9][25] ), .QN(n401)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][26]  ( .D(\i_MIPS/Register/n846 ), 
        .CK(clk), .RN(n4129), .Q(\i_MIPS/Register/register[9][26] ), .QN(n409)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][27]  ( .D(\i_MIPS/Register/n847 ), 
        .CK(clk), .RN(n4129), .Q(\i_MIPS/Register/register[9][27] ), .QN(n415)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][28]  ( .D(\i_MIPS/Register/n848 ), 
        .CK(clk), .RN(n4129), .Q(\i_MIPS/Register/register[9][28] ), .QN(n419)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][29]  ( .D(\i_MIPS/Register/n849 ), 
        .CK(clk), .RN(n4129), .Q(\i_MIPS/Register/register[9][29] ), .QN(n417)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][30]  ( .D(\i_MIPS/Register/n850 ), 
        .CK(clk), .RN(n4129), .Q(\i_MIPS/Register/register[9][30] ), .QN(n423)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][31]  ( .D(\i_MIPS/Register/n851 ), 
        .CK(clk), .RN(n4129), .Q(\i_MIPS/Register/register[9][31] ), .QN(n421)
         );
  DFFRX1 \i_MIPS/Register/register_reg[7][2]  ( .D(\i_MIPS/Register/n886 ), 
        .CK(clk), .RN(n4132), .Q(\i_MIPS/Register/register[7][2] ), .QN(n1180)
         );
  DFFRX1 \i_MIPS/Register/register_reg[7][3]  ( .D(\i_MIPS/Register/n887 ), 
        .CK(clk), .RN(n4132), .Q(\i_MIPS/Register/register[7][3] ), .QN(n1186)
         );
  DFFRX1 \i_MIPS/Register/register_reg[7][4]  ( .D(\i_MIPS/Register/n888 ), 
        .CK(clk), .RN(n4133), .Q(\i_MIPS/Register/register[7][4] ), .QN(n1134)
         );
  DFFRX1 \i_MIPS/Register/register_reg[7][5]  ( .D(\i_MIPS/Register/n889 ), 
        .CK(clk), .RN(n4133), .Q(\i_MIPS/Register/register[7][5] ), .QN(n1150)
         );
  DFFRX1 \i_MIPS/Register/register_reg[7][6]  ( .D(\i_MIPS/Register/n890 ), 
        .CK(clk), .RN(n4133), .Q(\i_MIPS/Register/register[7][6] ), .QN(n1162)
         );
  DFFRX1 \i_MIPS/Register/register_reg[7][7]  ( .D(\i_MIPS/Register/n891 ), 
        .CK(clk), .RN(n4133), .Q(\i_MIPS/Register/register[7][7] ), .QN(n1156)
         );
  DFFRX1 \i_MIPS/Register/register_reg[7][9]  ( .D(\i_MIPS/Register/n893 ), 
        .CK(clk), .RN(n4133), .Q(\i_MIPS/Register/register[7][9] ), .QN(n1122)
         );
  DFFRX1 \i_MIPS/Register/register_reg[7][10]  ( .D(\i_MIPS/Register/n894 ), 
        .CK(clk), .RN(n4133), .Q(\i_MIPS/Register/register[7][10] ), .QN(n1144) );
  DFFRX1 \i_MIPS/Register/register_reg[7][11]  ( .D(\i_MIPS/Register/n895 ), 
        .CK(clk), .RN(n4133), .Q(\i_MIPS/Register/register[7][11] ), .QN(n1139) );
  DFFRX1 \i_MIPS/Register/register_reg[7][12]  ( .D(\i_MIPS/Register/n896 ), 
        .CK(clk), .RN(n4133), .Q(\i_MIPS/Register/register[7][12] ), .QN(n1116) );
  DFFRX1 \i_MIPS/Register/register_reg[7][13]  ( .D(\i_MIPS/Register/n897 ), 
        .CK(clk), .RN(n4133), .Q(\i_MIPS/Register/register[7][13] ), .QN(n223)
         );
  DFFRX1 \i_MIPS/Register/register_reg[7][14]  ( .D(\i_MIPS/Register/n898 ), 
        .CK(clk), .RN(n4133), .Q(\i_MIPS/Register/register[7][14] ), .QN(n1128) );
  DFFRX1 \i_MIPS/Register/register_reg[7][15]  ( .D(\i_MIPS/Register/n899 ), 
        .CK(clk), .RN(n4133), .Q(\i_MIPS/Register/register[7][15] ), .QN(n1198) );
  DFFRX1 \i_MIPS/Register/register_reg[7][16]  ( .D(\i_MIPS/Register/n900 ), 
        .CK(clk), .RN(n4134), .Q(\i_MIPS/Register/register[7][16] ), .QN(n1222) );
  DFFRX1 \i_MIPS/Register/register_reg[7][17]  ( .D(\i_MIPS/Register/n901 ), 
        .CK(clk), .RN(n4134), .Q(\i_MIPS/Register/register[7][17] ), .QN(n1288) );
  DFFRX1 \i_MIPS/Register/register_reg[7][18]  ( .D(\i_MIPS/Register/n902 ), 
        .CK(clk), .RN(n4134), .Q(\i_MIPS/Register/register[7][18] ), .QN(n1282) );
  DFFRX1 \i_MIPS/Register/register_reg[7][19]  ( .D(\i_MIPS/Register/n903 ), 
        .CK(clk), .RN(n4134), .Q(\i_MIPS/Register/register[7][19] ), .QN(n1228) );
  DFFRX1 \i_MIPS/Register/register_reg[7][20]  ( .D(\i_MIPS/Register/n904 ), 
        .CK(clk), .RN(n4134), .Q(\i_MIPS/Register/register[7][20] ), .QN(n1276) );
  DFFRX1 \i_MIPS/Register/register_reg[7][21]  ( .D(\i_MIPS/Register/n905 ), 
        .CK(clk), .RN(n4134), .Q(\i_MIPS/Register/register[7][21] ), .QN(n1204) );
  DFFRX1 \i_MIPS/Register/register_reg[7][22]  ( .D(\i_MIPS/Register/n906 ), 
        .CK(clk), .RN(n4134), .Q(\i_MIPS/Register/register[7][22] ), .QN(n1264) );
  DFFRX1 \i_MIPS/Register/register_reg[7][23]  ( .D(\i_MIPS/Register/n907 ), 
        .CK(clk), .RN(n4134), .Q(\i_MIPS/Register/register[7][23] ), .QN(n1270) );
  DFFRX1 \i_MIPS/Register/register_reg[7][24]  ( .D(\i_MIPS/Register/n908 ), 
        .CK(clk), .RN(n4134), .Q(\i_MIPS/Register/register[7][24] ), .QN(n1210) );
  DFFRX1 \i_MIPS/Register/register_reg[7][25]  ( .D(\i_MIPS/Register/n909 ), 
        .CK(clk), .RN(n4134), .Q(\i_MIPS/Register/register[7][25] ), .QN(n1192) );
  DFFRX1 \i_MIPS/Register/register_reg[7][26]  ( .D(\i_MIPS/Register/n910 ), 
        .CK(clk), .RN(n4134), .Q(\i_MIPS/Register/register[7][26] ), .QN(n1216) );
  DFFRX1 \i_MIPS/Register/register_reg[7][27]  ( .D(\i_MIPS/Register/n911 ), 
        .CK(clk), .RN(n4134), .Q(\i_MIPS/Register/register[7][27] ), .QN(n1234) );
  DFFRX1 \i_MIPS/Register/register_reg[7][28]  ( .D(\i_MIPS/Register/n912 ), 
        .CK(clk), .RN(n4135), .Q(\i_MIPS/Register/register[7][28] ), .QN(n1246) );
  DFFRX1 \i_MIPS/Register/register_reg[7][29]  ( .D(\i_MIPS/Register/n913 ), 
        .CK(clk), .RN(n4135), .Q(\i_MIPS/Register/register[7][29] ), .QN(n1240) );
  DFFRX1 \i_MIPS/Register/register_reg[7][30]  ( .D(\i_MIPS/Register/n914 ), 
        .CK(clk), .RN(n4135), .Q(\i_MIPS/Register/register[7][30] ), .QN(n1258) );
  DFFRX1 \i_MIPS/Register/register_reg[7][31]  ( .D(\i_MIPS/Register/n915 ), 
        .CK(clk), .RN(n4135), .Q(\i_MIPS/Register/register[7][31] ), .QN(n1252) );
  DFFRX1 \i_MIPS/Register/register_reg[5][2]  ( .D(\i_MIPS/Register/n950 ), 
        .CK(clk), .RN(n4138), .Q(\i_MIPS/Register/register[5][2] ), .QN(n1182)
         );
  DFFRX1 \i_MIPS/Register/register_reg[5][3]  ( .D(\i_MIPS/Register/n951 ), 
        .CK(clk), .RN(n4138), .Q(\i_MIPS/Register/register[5][3] ), .QN(n1188)
         );
  DFFRX1 \i_MIPS/Register/register_reg[5][4]  ( .D(\i_MIPS/Register/n952 ), 
        .CK(clk), .RN(n4138), .Q(\i_MIPS/Register/register[5][4] ), .QN(n1136)
         );
  DFFRX1 \i_MIPS/Register/register_reg[5][15]  ( .D(\i_MIPS/Register/n963 ), 
        .CK(clk), .RN(n4139), .Q(\i_MIPS/Register/register[5][15] ), .QN(n1200) );
  DFFRX1 \i_MIPS/Register/register_reg[5][16]  ( .D(\i_MIPS/Register/n964 ), 
        .CK(clk), .RN(n4139), .Q(\i_MIPS/Register/register[5][16] ), .QN(n1224) );
  DFFRX1 \i_MIPS/Register/register_reg[5][17]  ( .D(\i_MIPS/Register/n965 ), 
        .CK(clk), .RN(n4139), .Q(\i_MIPS/Register/register[5][17] ), .QN(n1290) );
  DFFRX1 \i_MIPS/Register/register_reg[5][18]  ( .D(\i_MIPS/Register/n966 ), 
        .CK(clk), .RN(n4139), .Q(\i_MIPS/Register/register[5][18] ), .QN(n1284) );
  DFFRX1 \i_MIPS/Register/register_reg[5][19]  ( .D(\i_MIPS/Register/n967 ), 
        .CK(clk), .RN(n4139), .Q(\i_MIPS/Register/register[5][19] ), .QN(n1230) );
  DFFRX1 \i_MIPS/Register/register_reg[5][20]  ( .D(\i_MIPS/Register/n968 ), 
        .CK(clk), .RN(n4139), .Q(\i_MIPS/Register/register[5][20] ), .QN(n1278) );
  DFFRX1 \i_MIPS/Register/register_reg[5][21]  ( .D(\i_MIPS/Register/n969 ), 
        .CK(clk), .RN(n4139), .Q(\i_MIPS/Register/register[5][21] ), .QN(n1206) );
  DFFRX1 \i_MIPS/Register/register_reg[5][22]  ( .D(\i_MIPS/Register/n970 ), 
        .CK(clk), .RN(n4139), .Q(\i_MIPS/Register/register[5][22] ), .QN(n1266) );
  DFFRX1 \i_MIPS/Register/register_reg[5][23]  ( .D(\i_MIPS/Register/n971 ), 
        .CK(clk), .RN(n4139), .Q(\i_MIPS/Register/register[5][23] ), .QN(n1272) );
  DFFRX1 \i_MIPS/Register/register_reg[5][25]  ( .D(\i_MIPS/Register/n973 ), 
        .CK(clk), .RN(n4140), .Q(\i_MIPS/Register/register[5][25] ), .QN(n1194) );
  DFFRX1 \i_MIPS/Register/register_reg[5][27]  ( .D(\i_MIPS/Register/n975 ), 
        .CK(clk), .RN(n4140), .Q(\i_MIPS/Register/register[5][27] ), .QN(n1236) );
  DFFRX1 \i_MIPS/Register/register_reg[5][28]  ( .D(\i_MIPS/Register/n976 ), 
        .CK(clk), .RN(n4140), .Q(\i_MIPS/Register/register[5][28] ), .QN(n1248) );
  DFFRX1 \i_MIPS/Register/register_reg[5][29]  ( .D(\i_MIPS/Register/n977 ), 
        .CK(clk), .RN(n4140), .Q(\i_MIPS/Register/register[5][29] ), .QN(n1242) );
  DFFRX1 \i_MIPS/Register/register_reg[5][30]  ( .D(\i_MIPS/Register/n978 ), 
        .CK(clk), .RN(n4140), .Q(\i_MIPS/Register/register[5][30] ), .QN(n1260) );
  DFFRX1 \i_MIPS/Register/register_reg[5][31]  ( .D(\i_MIPS/Register/n979 ), 
        .CK(clk), .RN(n4140), .Q(\i_MIPS/Register/register[5][31] ), .QN(n1254) );
  DFFRX1 \i_MIPS/Register/register_reg[3][2]  ( .D(\i_MIPS/Register/n1014 ), 
        .CK(clk), .RN(n4143), .Q(\i_MIPS/Register/register[3][2] ), .QN(n1181)
         );
  DFFRX1 \i_MIPS/Register/register_reg[3][3]  ( .D(\i_MIPS/Register/n1015 ), 
        .CK(clk), .RN(n4143), .Q(\i_MIPS/Register/register[3][3] ), .QN(n1187)
         );
  DFFRX1 \i_MIPS/Register/register_reg[3][4]  ( .D(\i_MIPS/Register/n1016 ), 
        .CK(clk), .RN(n4143), .Q(\i_MIPS/Register/register[3][4] ), .QN(n1135)
         );
  DFFRX1 \i_MIPS/Register/register_reg[3][7]  ( .D(\i_MIPS/Register/n1019 ), 
        .CK(clk), .RN(n4143), .Q(\i_MIPS/Register/register[3][7] ), .QN(n1157)
         );
  DFFRX1 \i_MIPS/Register/register_reg[3][11]  ( .D(\i_MIPS/Register/n1023 ), 
        .CK(clk), .RN(n4144), .Q(\i_MIPS/Register/register[3][11] ), .QN(n1140) );
  DFFRX1 \i_MIPS/Register/register_reg[3][13]  ( .D(\i_MIPS/Register/n1025 ), 
        .CK(clk), .RN(n4144), .Q(\i_MIPS/Register/register[3][13] ), .QN(n1101) );
  DFFRX1 \i_MIPS/Register/register_reg[3][15]  ( .D(\i_MIPS/Register/n1027 ), 
        .CK(clk), .RN(n4144), .Q(\i_MIPS/Register/register[3][15] ), .QN(n1199) );
  DFFRX1 \i_MIPS/Register/register_reg[3][16]  ( .D(\i_MIPS/Register/n1028 ), 
        .CK(clk), .RN(n4144), .Q(\i_MIPS/Register/register[3][16] ), .QN(n1223) );
  DFFRX1 \i_MIPS/Register/register_reg[3][17]  ( .D(\i_MIPS/Register/n1029 ), 
        .CK(clk), .RN(n4144), .Q(\i_MIPS/Register/register[3][17] ), .QN(n1289) );
  DFFRX1 \i_MIPS/Register/register_reg[3][18]  ( .D(\i_MIPS/Register/n1030 ), 
        .CK(clk), .RN(n4144), .Q(\i_MIPS/Register/register[3][18] ), .QN(n1283) );
  DFFRX1 \i_MIPS/Register/register_reg[3][19]  ( .D(\i_MIPS/Register/n1031 ), 
        .CK(clk), .RN(n4144), .Q(\i_MIPS/Register/register[3][19] ), .QN(n1229) );
  DFFRX1 \i_MIPS/Register/register_reg[3][20]  ( .D(\i_MIPS/Register/n1032 ), 
        .CK(clk), .RN(n4145), .Q(\i_MIPS/Register/register[3][20] ), .QN(n1277) );
  DFFRX1 \i_MIPS/Register/register_reg[3][21]  ( .D(\i_MIPS/Register/n1033 ), 
        .CK(clk), .RN(n4145), .Q(\i_MIPS/Register/register[3][21] ), .QN(n1205) );
  DFFRX1 \i_MIPS/Register/register_reg[3][22]  ( .D(\i_MIPS/Register/n1034 ), 
        .CK(clk), .RN(n4145), .Q(\i_MIPS/Register/register[3][22] ), .QN(n1265) );
  DFFRX1 \i_MIPS/Register/register_reg[3][23]  ( .D(\i_MIPS/Register/n1035 ), 
        .CK(clk), .RN(n4145), .Q(\i_MIPS/Register/register[3][23] ), .QN(n1271) );
  DFFRX1 \i_MIPS/Register/register_reg[3][25]  ( .D(\i_MIPS/Register/n1037 ), 
        .CK(clk), .RN(n4145), .Q(\i_MIPS/Register/register[3][25] ), .QN(n1193) );
  DFFRX1 \i_MIPS/Register/register_reg[3][27]  ( .D(\i_MIPS/Register/n1039 ), 
        .CK(clk), .RN(n4145), .Q(\i_MIPS/Register/register[3][27] ), .QN(n1235) );
  DFFRX1 \i_MIPS/Register/register_reg[3][28]  ( .D(\i_MIPS/Register/n1040 ), 
        .CK(clk), .RN(n4145), .Q(\i_MIPS/Register/register[3][28] ), .QN(n1247) );
  DFFRX1 \i_MIPS/Register/register_reg[3][29]  ( .D(\i_MIPS/Register/n1041 ), 
        .CK(clk), .RN(n4145), .Q(\i_MIPS/Register/register[3][29] ), .QN(n1241) );
  DFFRX1 \i_MIPS/Register/register_reg[3][30]  ( .D(\i_MIPS/Register/n1042 ), 
        .CK(clk), .RN(n4145), .Q(\i_MIPS/Register/register[3][30] ), .QN(n1259) );
  DFFRX1 \i_MIPS/Register/register_reg[3][31]  ( .D(\i_MIPS/Register/n1043 ), 
        .CK(clk), .RN(n4145), .Q(\i_MIPS/Register/register[3][31] ), .QN(n1253) );
  DFFRX1 \i_MIPS/Register/register_reg[1][4]  ( .D(\i_MIPS/Register/n1080 ), 
        .CK(clk), .RN(n4149), .Q(\i_MIPS/Register/register[1][4] ), .QN(n1298)
         );
  DFFRX1 \i_MIPS/Register/register_reg[1][15]  ( .D(\i_MIPS/Register/n1091 ), 
        .CK(clk), .RN(n4149), .Q(\i_MIPS/Register/register[1][15] ), .QN(n1317) );
  DFFRX1 \i_MIPS/Register/register_reg[1][16]  ( .D(\i_MIPS/Register/n1092 ), 
        .CK(clk), .RN(n4150), .Q(\i_MIPS/Register/register[1][16] ), .QN(n1325) );
  DFFRX1 \i_MIPS/Register/register_reg[1][17]  ( .D(\i_MIPS/Register/n1093 ), 
        .CK(clk), .RN(n4150), .Q(\i_MIPS/Register/register[1][17] ), .QN(n1347) );
  DFFRX1 \i_MIPS/Register/register_reg[1][18]  ( .D(\i_MIPS/Register/n1094 ), 
        .CK(clk), .RN(n4150), .Q(\i_MIPS/Register/register[1][18] ), .QN(n1345) );
  DFFRX1 \i_MIPS/Register/register_reg[1][19]  ( .D(\i_MIPS/Register/n1095 ), 
        .CK(clk), .RN(n4150), .Q(\i_MIPS/Register/register[1][19] ), .QN(n1327) );
  DFFRX1 \i_MIPS/Register/register_reg[1][20]  ( .D(\i_MIPS/Register/n1096 ), 
        .CK(clk), .RN(n4150), .Q(\i_MIPS/Register/register[1][20] ), .QN(n1343) );
  DFFRX1 \i_MIPS/Register/register_reg[1][21]  ( .D(\i_MIPS/Register/n1097 ), 
        .CK(clk), .RN(n4150), .Q(\i_MIPS/Register/register[1][21] ), .QN(n1319) );
  DFFRX1 \i_MIPS/Register/register_reg[1][22]  ( .D(\i_MIPS/Register/n1098 ), 
        .CK(clk), .RN(n4150), .Q(\i_MIPS/Register/register[1][22] ), .QN(n1339) );
  DFFRX1 \i_MIPS/Register/register_reg[1][23]  ( .D(\i_MIPS/Register/n1099 ), 
        .CK(clk), .RN(n4150), .Q(\i_MIPS/Register/register[1][23] ), .QN(n1341) );
  DFFRX1 \i_MIPS/Register/register_reg[1][25]  ( .D(\i_MIPS/Register/n1101 ), 
        .CK(clk), .RN(n4150), .Q(\i_MIPS/Register/register[1][25] ), .QN(n1315) );
  DFFRX1 \i_MIPS/Register/register_reg[1][27]  ( .D(\i_MIPS/Register/n1103 ), 
        .CK(clk), .RN(n4150), .Q(\i_MIPS/Register/register[1][27] ), .QN(n1329) );
  DFFRX1 \i_MIPS/Register/register_reg[1][28]  ( .D(\i_MIPS/Register/n1104 ), 
        .CK(clk), .RN(n4151), .Q(\i_MIPS/Register/register[1][28] ), .QN(n1333) );
  DFFRX1 \i_MIPS/Register/register_reg[1][29]  ( .D(\i_MIPS/Register/n1105 ), 
        .CK(clk), .RN(n4151), .Q(\i_MIPS/Register/register[1][29] ), .QN(n1331) );
  DFFRX1 \i_MIPS/Register/register_reg[1][30]  ( .D(\i_MIPS/Register/n1106 ), 
        .CK(clk), .RN(n4151), .Q(\i_MIPS/Register/register[1][30] ), .QN(n1337) );
  DFFRX1 \i_MIPS/Register/register_reg[1][31]  ( .D(\i_MIPS/Register/n1107 ), 
        .CK(clk), .RN(n4151), .Q(\i_MIPS/Register/register[1][31] ), .QN(n1335) );
  DFFRX1 \I_cache/cache_reg[0][10]  ( .D(n10084), .CK(clk), .RN(n4264), .Q(
        \I_cache/cache[0][10] ), .QN(n632) );
  DFFRX1 \I_cache/cache_reg[1][10]  ( .D(n10083), .CK(clk), .RN(n4264), .Q(
        \I_cache/cache[1][10] ), .QN(n1551) );
  DFFRX1 \I_cache/cache_reg[2][10]  ( .D(n10082), .CK(clk), .RN(n4264), .Q(
        \I_cache/cache[2][10] ), .QN(n631) );
  DFFRX1 \I_cache/cache_reg[4][10]  ( .D(n10080), .CK(clk), .RN(n4264), .Q(
        \I_cache/cache[4][10] ), .QN(n670) );
  DFFRX1 \I_cache/cache_reg[6][10]  ( .D(n10078), .CK(clk), .RN(n4264), .Q(
        \I_cache/cache[6][10] ), .QN(n630) );
  DFFRX1 \I_cache/cache_reg[0][14]  ( .D(n10052), .CK(clk), .RN(n4266), .Q(
        \I_cache/cache[0][14] ), .QN(n520) );
  DFFRX1 \I_cache/cache_reg[2][14]  ( .D(n10050), .CK(clk), .RN(n4266), .Q(
        \I_cache/cache[2][14] ), .QN(n519) );
  DFFRX1 \I_cache/cache_reg[0][16]  ( .D(n10036), .CK(clk), .RN(n4268), .Q(
        \I_cache/cache[0][16] ), .QN(n1856) );
  DFFRX1 \I_cache/cache_reg[1][16]  ( .D(n10035), .CK(clk), .RN(n4268), .Q(
        \I_cache/cache[1][16] ), .QN(n922) );
  DFFRX1 \I_cache/cache_reg[2][16]  ( .D(n10034), .CK(clk), .RN(n4268), .Q(
        \I_cache/cache[2][16] ), .QN(n1857) );
  DFFRX1 \I_cache/cache_reg[3][16]  ( .D(n10033), .CK(clk), .RN(n4268), .Q(
        \I_cache/cache[3][16] ), .QN(n923) );
  DFFRX1 \I_cache/cache_reg[4][16]  ( .D(n10032), .CK(clk), .RN(n4268), .Q(
        \I_cache/cache[4][16] ), .QN(n810) );
  DFFRX1 \I_cache/cache_reg[5][16]  ( .D(n10031), .CK(clk), .RN(n4268), .Q(
        \I_cache/cache[5][16] ), .QN(n1743) );
  DFFRX1 \I_cache/cache_reg[6][16]  ( .D(n10030), .CK(clk), .RN(n4268), .Q(
        \I_cache/cache[6][16] ), .QN(n852) );
  DFFRX1 \I_cache/cache_reg[7][16]  ( .D(n10029), .CK(clk), .RN(n4268), .Q(
        \I_cache/cache[7][16] ), .QN(n1785) );
  DFFRX1 \I_cache/cache_reg[0][17]  ( .D(n10028), .CK(clk), .RN(n4268), .Q(
        \I_cache/cache[0][17] ), .QN(n888) );
  DFFRX1 \I_cache/cache_reg[1][17]  ( .D(n10027), .CK(clk), .RN(n4268), .Q(
        \I_cache/cache[1][17] ), .QN(n1821) );
  DFFRX1 \I_cache/cache_reg[2][17]  ( .D(n10026), .CK(clk), .RN(n4268), .Q(
        \I_cache/cache[2][17] ), .QN(n890) );
  DFFRX1 \I_cache/cache_reg[3][17]  ( .D(n10025), .CK(clk), .RN(n4268), .Q(
        \I_cache/cache[3][17] ), .QN(n1823) );
  DFFRX1 \I_cache/cache_reg[4][17]  ( .D(n10024), .CK(clk), .RN(n4269), .Q(
        \I_cache/cache[4][17] ), .QN(n889) );
  DFFRX1 \I_cache/cache_reg[5][17]  ( .D(n10023), .CK(clk), .RN(n4269), .Q(
        \I_cache/cache[5][17] ), .QN(n1822) );
  DFFRX1 \I_cache/cache_reg[6][17]  ( .D(n10022), .CK(clk), .RN(n4269), .Q(
        \I_cache/cache[6][17] ), .QN(n908) );
  DFFRX1 \I_cache/cache_reg[7][17]  ( .D(n10021), .CK(clk), .RN(n4269), .Q(
        \I_cache/cache[7][17] ), .QN(n1841) );
  DFFRX1 \I_cache/cache_reg[0][18]  ( .D(n10020), .CK(clk), .RN(n4269), .Q(
        \I_cache/cache[0][18] ), .QN(n1854) );
  DFFRX1 \I_cache/cache_reg[1][18]  ( .D(n10019), .CK(clk), .RN(n4269), .Q(
        \I_cache/cache[1][18] ), .QN(n920) );
  DFFRX1 \I_cache/cache_reg[2][18]  ( .D(n10018), .CK(clk), .RN(n4269), .Q(
        \I_cache/cache[2][18] ), .QN(n1855) );
  DFFRX1 \I_cache/cache_reg[3][18]  ( .D(n10017), .CK(clk), .RN(n4269), .Q(
        \I_cache/cache[3][18] ), .QN(n921) );
  DFFRX1 \I_cache/cache_reg[4][18]  ( .D(n10016), .CK(clk), .RN(n4269), .Q(
        \I_cache/cache[4][18] ), .QN(n797) );
  DFFRX1 \I_cache/cache_reg[5][18]  ( .D(n10015), .CK(clk), .RN(n4269), .Q(
        \I_cache/cache[5][18] ), .QN(n1730) );
  DFFRX1 \I_cache/cache_reg[6][18]  ( .D(n10014), .CK(clk), .RN(n4269), .Q(
        \I_cache/cache[6][18] ), .QN(n847) );
  DFFRX1 \I_cache/cache_reg[7][18]  ( .D(n10013), .CK(clk), .RN(n4269), .Q(
        \I_cache/cache[7][18] ), .QN(n1780) );
  DFFRX1 \I_cache/cache_reg[0][19]  ( .D(n10012), .CK(clk), .RN(n4270), .Q(
        \I_cache/cache[0][19] ), .QN(n1848) );
  DFFRX1 \I_cache/cache_reg[1][19]  ( .D(n10011), .CK(clk), .RN(n4270), .Q(
        \I_cache/cache[1][19] ), .QN(n914) );
  DFFRX1 \I_cache/cache_reg[2][19]  ( .D(n10010), .CK(clk), .RN(n4270), .Q(
        \I_cache/cache[2][19] ), .QN(n1849) );
  DFFRX1 \I_cache/cache_reg[3][19]  ( .D(n10009), .CK(clk), .RN(n4270), .Q(
        \I_cache/cache[3][19] ), .QN(n915) );
  DFFRX1 \I_cache/cache_reg[4][19]  ( .D(n10008), .CK(clk), .RN(n4270), .Q(
        \I_cache/cache[4][19] ), .QN(n773) );
  DFFRX1 \I_cache/cache_reg[5][19]  ( .D(n10007), .CK(clk), .RN(n4270), .Q(
        \I_cache/cache[5][19] ), .QN(n1706) );
  DFFRX1 \I_cache/cache_reg[6][19]  ( .D(n10006), .CK(clk), .RN(n4270), .Q(
        \I_cache/cache[6][19] ), .QN(n837) );
  DFFRX1 \I_cache/cache_reg[7][19]  ( .D(n10005), .CK(clk), .RN(n4270), .Q(
        \I_cache/cache[7][19] ), .QN(n1770) );
  DFFRX1 \I_cache/cache_reg[0][20]  ( .D(n10004), .CK(clk), .RN(n4270), .Q(
        \I_cache/cache[0][20] ), .QN(n1864) );
  DFFRX1 \I_cache/cache_reg[1][20]  ( .D(n10003), .CK(clk), .RN(n4270), .Q(
        \I_cache/cache[1][20] ), .QN(n930) );
  DFFRX1 \I_cache/cache_reg[2][20]  ( .D(n10002), .CK(clk), .RN(n4270), .Q(
        \I_cache/cache[2][20] ), .QN(n1866) );
  DFFRX1 \I_cache/cache_reg[3][20]  ( .D(n10001), .CK(clk), .RN(n4270), .Q(
        \I_cache/cache[3][20] ), .QN(n932) );
  DFFRX1 \I_cache/cache_reg[4][20]  ( .D(n10000), .CK(clk), .RN(n4271), .Q(
        \I_cache/cache[4][20] ), .QN(n1865) );
  DFFRX1 \I_cache/cache_reg[5][20]  ( .D(n9999), .CK(clk), .RN(n4271), .Q(
        \I_cache/cache[5][20] ), .QN(n931) );
  DFFRX1 \I_cache/cache_reg[6][20]  ( .D(n9998), .CK(clk), .RN(n4271), .Q(
        \I_cache/cache[6][20] ), .QN(n898) );
  DFFRX1 \I_cache/cache_reg[7][20]  ( .D(n9997), .CK(clk), .RN(n4271), .Q(
        \I_cache/cache[7][20] ), .QN(n1831) );
  DFFRX1 \I_cache/cache_reg[0][21]  ( .D(n9996), .CK(clk), .RN(n4271), .Q(
        \I_cache/cache[0][21] ), .QN(n1851) );
  DFFRX1 \I_cache/cache_reg[1][21]  ( .D(n9995), .CK(clk), .RN(n4271), .Q(
        \I_cache/cache[1][21] ), .QN(n917) );
  DFFRX1 \I_cache/cache_reg[2][21]  ( .D(n9994), .CK(clk), .RN(n4271), .Q(
        \I_cache/cache[2][21] ), .QN(n1852) );
  DFFRX1 \I_cache/cache_reg[3][21]  ( .D(n9993), .CK(clk), .RN(n4271), .Q(
        \I_cache/cache[3][21] ), .QN(n918) );
  DFFRX1 \I_cache/cache_reg[4][21]  ( .D(n9992), .CK(clk), .RN(n4271), .Q(
        \I_cache/cache[4][21] ), .QN(n785) );
  DFFRX1 \I_cache/cache_reg[5][21]  ( .D(n9991), .CK(clk), .RN(n4271), .Q(
        \I_cache/cache[5][21] ), .QN(n1718) );
  DFFRX1 \I_cache/cache_reg[6][21]  ( .D(n9990), .CK(clk), .RN(n4271), .Q(
        \I_cache/cache[6][21] ), .QN(n842) );
  DFFRX1 \I_cache/cache_reg[7][21]  ( .D(n9989), .CK(clk), .RN(n4271), .Q(
        \I_cache/cache[7][21] ), .QN(n1775) );
  DFFRX1 \I_cache/cache_reg[0][22]  ( .D(n9988), .CK(clk), .RN(n4272), .Q(
        \I_cache/cache[0][22] ), .QN(n1869) );
  DFFRX1 \I_cache/cache_reg[1][22]  ( .D(n9987), .CK(clk), .RN(n4272), .Q(
        \I_cache/cache[1][22] ), .QN(n935) );
  DFFRX1 \I_cache/cache_reg[2][22]  ( .D(n9986), .CK(clk), .RN(n4272), .Q(
        \I_cache/cache[2][22] ), .QN(n1871) );
  DFFRX1 \I_cache/cache_reg[3][22]  ( .D(n9985), .CK(clk), .RN(n4272), .Q(
        \I_cache/cache[3][22] ), .QN(n937) );
  DFFRX1 \I_cache/cache_reg[4][22]  ( .D(n9984), .CK(clk), .RN(n4272), .Q(
        \I_cache/cache[4][22] ), .QN(n1870) );
  DFFRX1 \I_cache/cache_reg[5][22]  ( .D(n9983), .CK(clk), .RN(n4272), .Q(
        \I_cache/cache[5][22] ), .QN(n936) );
  DFFRX1 \I_cache/cache_reg[6][22]  ( .D(n9982), .CK(clk), .RN(n4272), .Q(
        \I_cache/cache[6][22] ), .QN(n910) );
  DFFRX1 \I_cache/cache_reg[7][22]  ( .D(n9981), .CK(clk), .RN(n4272), .Q(
        \I_cache/cache[7][22] ), .QN(n1843) );
  DFFRX1 \I_cache/cache_reg[0][23]  ( .D(n9980), .CK(clk), .RN(n4272), .Q(
        \I_cache/cache[0][23] ), .QN(n1879) );
  DFFRX1 \I_cache/cache_reg[1][23]  ( .D(n9979), .CK(clk), .RN(n4272), .Q(
        \I_cache/cache[1][23] ), .QN(n945) );
  DFFRX1 \I_cache/cache_reg[2][23]  ( .D(n9978), .CK(clk), .RN(n4272), .Q(
        \I_cache/cache[2][23] ), .QN(n881) );
  DFFRX1 \I_cache/cache_reg[3][23]  ( .D(n9977), .CK(clk), .RN(n4272), .Q(
        \I_cache/cache[3][23] ), .QN(n1814) );
  DFFRX1 \I_cache/cache_reg[4][23]  ( .D(n9976), .CK(clk), .RN(n4273), .Q(
        \I_cache/cache[4][23] ), .QN(n880) );
  DFFRX1 \I_cache/cache_reg[5][23]  ( .D(n9975), .CK(clk), .RN(n4273), .Q(
        \I_cache/cache[5][23] ), .QN(n1813) );
  DFFRX1 \I_cache/cache_reg[6][23]  ( .D(n9974), .CK(clk), .RN(n4273), .Q(
        \I_cache/cache[6][23] ), .QN(n905) );
  DFFRX1 \I_cache/cache_reg[7][23]  ( .D(n9973), .CK(clk), .RN(n4273), .Q(
        \I_cache/cache[7][23] ), .QN(n1838) );
  DFFRX1 \I_cache/cache_reg[0][24]  ( .D(n9972), .CK(clk), .RN(n4273), .Q(
        \I_cache/cache[0][24] ), .QN(n1858) );
  DFFRX1 \I_cache/cache_reg[1][24]  ( .D(n9971), .CK(clk), .RN(n4273), .Q(
        \I_cache/cache[1][24] ), .QN(n924) );
  DFFRX1 \I_cache/cache_reg[2][24]  ( .D(n9970), .CK(clk), .RN(n4273), .Q(
        \I_cache/cache[2][24] ), .QN(n1860) );
  DFFRX1 \I_cache/cache_reg[3][24]  ( .D(n9969), .CK(clk), .RN(n4273), .Q(
        \I_cache/cache[3][24] ), .QN(n926) );
  DFFRX1 \I_cache/cache_reg[4][24]  ( .D(n9968), .CK(clk), .RN(n4273), .Q(
        \I_cache/cache[4][24] ), .QN(n1859) );
  DFFRX1 \I_cache/cache_reg[5][24]  ( .D(n9967), .CK(clk), .RN(n4273), .Q(
        \I_cache/cache[5][24] ), .QN(n925) );
  DFFRX1 \I_cache/cache_reg[6][24]  ( .D(n9966), .CK(clk), .RN(n4273), .Q(
        \I_cache/cache[6][24] ), .QN(n1880) );
  DFFRX1 \I_cache/cache_reg[7][24]  ( .D(n9965), .CK(clk), .RN(n4273), .Q(
        \I_cache/cache[7][24] ), .QN(n946) );
  DFFRX1 \I_cache/cache_reg[0][25]  ( .D(n9964), .CK(clk), .RN(n4274), .Q(
        \I_cache/cache[0][25] ), .QN(n1874) );
  DFFRX1 \I_cache/cache_reg[1][25]  ( .D(n9963), .CK(clk), .RN(n4274), .Q(
        \I_cache/cache[1][25] ), .QN(n940) );
  DFFRX1 \I_cache/cache_reg[2][25]  ( .D(n9962), .CK(clk), .RN(n4274), .Q(
        \I_cache/cache[2][25] ), .QN(n1876) );
  DFFRX1 \I_cache/cache_reg[3][25]  ( .D(n9961), .CK(clk), .RN(n4274), .Q(
        \I_cache/cache[3][25] ), .QN(n942) );
  DFFRX1 \I_cache/cache_reg[4][25]  ( .D(n9960), .CK(clk), .RN(n4274), .Q(
        \I_cache/cache[4][25] ), .QN(n1875) );
  DFFRX1 \I_cache/cache_reg[5][25]  ( .D(n9959), .CK(clk), .RN(n4274), .Q(
        \I_cache/cache[5][25] ), .QN(n941) );
  DFFRX1 \I_cache/cache_reg[6][25]  ( .D(n9958), .CK(clk), .RN(n4274), .Q(
        \I_cache/cache[6][25] ), .QN(n902) );
  DFFRX1 \I_cache/cache_reg[7][25]  ( .D(n9957), .CK(clk), .RN(n4274), .Q(
        \I_cache/cache[7][25] ), .QN(n1835) );
  DFFRX1 \I_cache/cache_reg[0][26]  ( .D(n9956), .CK(clk), .RN(n4274), .Q(
        \I_cache/cache[0][26] ), .QN(n695) );
  DFFRX1 \I_cache/cache_reg[1][26]  ( .D(n9955), .CK(clk), .RN(n4274), .Q(
        \I_cache/cache[1][26] ), .QN(n1628) );
  DFFRX1 \I_cache/cache_reg[2][26]  ( .D(n9954), .CK(clk), .RN(n4274), .Q(
        \I_cache/cache[2][26] ), .QN(n697) );
  DFFRX1 \I_cache/cache_reg[3][26]  ( .D(n9953), .CK(clk), .RN(n4274), .Q(
        \I_cache/cache[3][26] ), .QN(n1630) );
  DFFRX1 \I_cache/cache_reg[4][26]  ( .D(n9952), .CK(clk), .RN(n4275), .Q(
        \I_cache/cache[4][26] ), .QN(n696) );
  DFFRX1 \I_cache/cache_reg[5][26]  ( .D(n9951), .CK(clk), .RN(n4275), .Q(
        \I_cache/cache[5][26] ), .QN(n1629) );
  DFFRX1 \I_cache/cache_reg[6][26]  ( .D(n9950), .CK(clk), .RN(n4275), .Q(
        \I_cache/cache[6][26] ), .QN(n811) );
  DFFRX1 \I_cache/cache_reg[7][26]  ( .D(n9949), .CK(clk), .RN(n4275), .Q(
        \I_cache/cache[7][26] ), .QN(n1744) );
  DFFRX1 \I_cache/cache_reg[0][27]  ( .D(n9948), .CK(clk), .RN(n4275), .Q(
        \I_cache/cache[0][27] ), .QN(n752) );
  DFFRX1 \I_cache/cache_reg[1][27]  ( .D(n9947), .CK(clk), .RN(n4275), .Q(
        \I_cache/cache[1][27] ), .QN(n1685) );
  DFFRX1 \I_cache/cache_reg[2][27]  ( .D(n9946), .CK(clk), .RN(n4275), .Q(
        \I_cache/cache[2][27] ), .QN(n754) );
  DFFRX1 \I_cache/cache_reg[3][27]  ( .D(n9945), .CK(clk), .RN(n4275), .Q(
        \I_cache/cache[3][27] ), .QN(n1687) );
  DFFRX1 \I_cache/cache_reg[4][27]  ( .D(n9944), .CK(clk), .RN(n4275), .Q(
        \I_cache/cache[4][27] ), .QN(n753) );
  DFFRX1 \I_cache/cache_reg[5][27]  ( .D(n9943), .CK(clk), .RN(n4275), .Q(
        \I_cache/cache[5][27] ), .QN(n1686) );
  DFFRX1 \I_cache/cache_reg[6][27]  ( .D(n9942), .CK(clk), .RN(n4275), .Q(
        \I_cache/cache[6][27] ), .QN(n830) );
  DFFRX1 \I_cache/cache_reg[7][27]  ( .D(n9941), .CK(clk), .RN(n4275), .Q(
        \I_cache/cache[7][27] ), .QN(n1763) );
  DFFRX1 \I_cache/cache_reg[0][28]  ( .D(n9940), .CK(clk), .RN(n4276), .Q(
        \I_cache/cache[0][28] ), .QN(n740) );
  DFFRX1 \I_cache/cache_reg[1][28]  ( .D(n9939), .CK(clk), .RN(n4276), .Q(
        \I_cache/cache[1][28] ), .QN(n1673) );
  DFFRX1 \I_cache/cache_reg[2][28]  ( .D(n9938), .CK(clk), .RN(n4276), .Q(
        \I_cache/cache[2][28] ), .QN(n742) );
  DFFRX1 \I_cache/cache_reg[3][28]  ( .D(n9937), .CK(clk), .RN(n4276), .Q(
        \I_cache/cache[3][28] ), .QN(n1675) );
  DFFRX1 \I_cache/cache_reg[4][28]  ( .D(n9936), .CK(clk), .RN(n4276), .Q(
        \I_cache/cache[4][28] ), .QN(n741) );
  DFFRX1 \I_cache/cache_reg[5][28]  ( .D(n9935), .CK(clk), .RN(n4276), .Q(
        \I_cache/cache[5][28] ), .QN(n1674) );
  DFFRX1 \I_cache/cache_reg[6][28]  ( .D(n9934), .CK(clk), .RN(n4276), .Q(
        \I_cache/cache[6][28] ), .QN(n826) );
  DFFRX1 \I_cache/cache_reg[7][28]  ( .D(n9933), .CK(clk), .RN(n4276), .Q(
        \I_cache/cache[7][28] ), .QN(n1759) );
  DFFRX1 \I_cache/cache_reg[0][29]  ( .D(n9932), .CK(clk), .RN(n4276), .Q(
        \I_cache/cache[0][29] ), .QN(n707) );
  DFFRX1 \I_cache/cache_reg[1][29]  ( .D(n9931), .CK(clk), .RN(n4276), .Q(
        \I_cache/cache[1][29] ), .QN(n1640) );
  DFFRX1 \I_cache/cache_reg[2][29]  ( .D(n9930), .CK(clk), .RN(n4276), .Q(
        \I_cache/cache[2][29] ), .QN(n709) );
  DFFRX1 \I_cache/cache_reg[3][29]  ( .D(n9929), .CK(clk), .RN(n4276), .Q(
        \I_cache/cache[3][29] ), .QN(n1642) );
  DFFRX1 \I_cache/cache_reg[4][29]  ( .D(n9928), .CK(clk), .RN(n4277), .Q(
        \I_cache/cache[4][29] ), .QN(n708) );
  DFFRX1 \I_cache/cache_reg[5][29]  ( .D(n9927), .CK(clk), .RN(n4277), .Q(
        \I_cache/cache[5][29] ), .QN(n1641) );
  DFFRX1 \I_cache/cache_reg[6][29]  ( .D(n9926), .CK(clk), .RN(n4277), .Q(
        \I_cache/cache[6][29] ), .QN(n815) );
  DFFRX1 \I_cache/cache_reg[7][29]  ( .D(n9925), .CK(clk), .RN(n4277), .Q(
        \I_cache/cache[7][29] ), .QN(n1748) );
  DFFRX1 \I_cache/cache_reg[0][30]  ( .D(n9924), .CK(clk), .RN(n4277), .Q(
        \I_cache/cache[0][30] ), .QN(n728) );
  DFFRX1 \I_cache/cache_reg[1][30]  ( .D(n9923), .CK(clk), .RN(n4277), .Q(
        \I_cache/cache[1][30] ), .QN(n1661) );
  DFFRX1 \I_cache/cache_reg[2][30]  ( .D(n9922), .CK(clk), .RN(n4277), .Q(
        \I_cache/cache[2][30] ), .QN(n730) );
  DFFRX1 \I_cache/cache_reg[3][30]  ( .D(n9921), .CK(clk), .RN(n4277), .Q(
        \I_cache/cache[3][30] ), .QN(n1663) );
  DFFRX1 \I_cache/cache_reg[4][30]  ( .D(n9920), .CK(clk), .RN(n4277), .Q(
        \I_cache/cache[4][30] ), .QN(n729) );
  DFFRX1 \I_cache/cache_reg[5][30]  ( .D(n9919), .CK(clk), .RN(n4277), .Q(
        \I_cache/cache[5][30] ), .QN(n1662) );
  DFFRX1 \I_cache/cache_reg[6][30]  ( .D(n9918), .CK(clk), .RN(n4277), .Q(
        \I_cache/cache[6][30] ), .QN(n822) );
  DFFRX1 \I_cache/cache_reg[7][30]  ( .D(n9917), .CK(clk), .RN(n4277), .Q(
        \I_cache/cache[7][30] ), .QN(n1755) );
  DFFRX1 \I_cache/cache_reg[0][31]  ( .D(n9916), .CK(clk), .RN(n4278), .Q(
        \I_cache/cache[0][31] ), .QN(n719) );
  DFFRX1 \I_cache/cache_reg[1][31]  ( .D(n9915), .CK(clk), .RN(n4278), .Q(
        \I_cache/cache[1][31] ), .QN(n1652) );
  DFFRX1 \I_cache/cache_reg[2][31]  ( .D(n9914), .CK(clk), .RN(n4278), .Q(
        \I_cache/cache[2][31] ), .QN(n721) );
  DFFRX1 \I_cache/cache_reg[3][31]  ( .D(n9913), .CK(clk), .RN(n4278), .Q(
        \I_cache/cache[3][31] ), .QN(n1654) );
  DFFRX1 \I_cache/cache_reg[4][31]  ( .D(n9912), .CK(clk), .RN(n4278), .Q(
        \I_cache/cache[4][31] ), .QN(n720) );
  DFFRX1 \I_cache/cache_reg[5][31]  ( .D(n9911), .CK(clk), .RN(n4278), .Q(
        \I_cache/cache[5][31] ), .QN(n1653) );
  DFFRX1 \I_cache/cache_reg[6][31]  ( .D(n9910), .CK(clk), .RN(n4278), .Q(
        \I_cache/cache[6][31] ), .QN(n819) );
  DFFRX1 \I_cache/cache_reg[7][31]  ( .D(n9909), .CK(clk), .RN(n4278), .Q(
        \I_cache/cache[7][31] ), .QN(n1752) );
  DFFRX1 \I_cache/cache_reg[0][42]  ( .D(n9828), .CK(clk), .RN(n4285), .Q(
        \I_cache/cache[0][42] ), .QN(n629) );
  DFFRX1 \I_cache/cache_reg[2][42]  ( .D(n9826), .CK(clk), .RN(n4285), .Q(
        \I_cache/cache[2][42] ), .QN(n628) );
  DFFRX1 \I_cache/cache_reg[4][42]  ( .D(n9824), .CK(clk), .RN(n4285), .Q(
        \I_cache/cache[4][42] ), .QN(n669) );
  DFFRX1 \I_cache/cache_reg[0][46]  ( .D(n9796), .CK(clk), .RN(n4288), .Q(
        \I_cache/cache[0][46] ), .QN(n596) );
  DFFRX1 \I_cache/cache_reg[0][48]  ( .D(n9780), .CK(clk), .RN(n4289), .Q(
        \I_cache/cache[0][48] ), .QN(n804) );
  DFFRX1 \I_cache/cache_reg[1][48]  ( .D(n9779), .CK(clk), .RN(n4289), .Q(
        \I_cache/cache[1][48] ), .QN(n1737) );
  DFFRX1 \I_cache/cache_reg[2][48]  ( .D(n9778), .CK(clk), .RN(n4289), .Q(
        \I_cache/cache[2][48] ), .QN(n806) );
  DFFRX1 \I_cache/cache_reg[3][48]  ( .D(n9777), .CK(clk), .RN(n4289), .Q(
        \I_cache/cache[3][48] ), .QN(n1739) );
  DFFRX1 \I_cache/cache_reg[4][48]  ( .D(n9776), .CK(clk), .RN(n4289), .Q(
        \I_cache/cache[4][48] ), .QN(n805) );
  DFFRX1 \I_cache/cache_reg[5][48]  ( .D(n9775), .CK(clk), .RN(n4289), .Q(
        \I_cache/cache[5][48] ), .QN(n1738) );
  DFFRX1 \I_cache/cache_reg[6][48]  ( .D(n9774), .CK(clk), .RN(n4289), .Q(
        \I_cache/cache[6][48] ), .QN(n850) );
  DFFRX1 \I_cache/cache_reg[7][48]  ( .D(n9773), .CK(clk), .RN(n4289), .Q(
        \I_cache/cache[7][48] ), .QN(n1783) );
  DFFRX1 \I_cache/cache_reg[0][49]  ( .D(n9772), .CK(clk), .RN(n4290), .Q(
        \I_cache/cache[0][49] ), .QN(n891) );
  DFFRX1 \I_cache/cache_reg[1][49]  ( .D(n9771), .CK(clk), .RN(n4290), .Q(
        \I_cache/cache[1][49] ), .QN(n1824) );
  DFFRX1 \I_cache/cache_reg[2][49]  ( .D(n9770), .CK(clk), .RN(n4290), .Q(
        \I_cache/cache[2][49] ), .QN(n893) );
  DFFRX1 \I_cache/cache_reg[3][49]  ( .D(n9769), .CK(clk), .RN(n4290), .Q(
        \I_cache/cache[3][49] ), .QN(n1826) );
  DFFRX1 \I_cache/cache_reg[4][49]  ( .D(n9768), .CK(clk), .RN(n4290), .Q(
        \I_cache/cache[4][49] ), .QN(n892) );
  DFFRX1 \I_cache/cache_reg[5][49]  ( .D(n9767), .CK(clk), .RN(n4290), .Q(
        \I_cache/cache[5][49] ), .QN(n1825) );
  DFFRX1 \I_cache/cache_reg[6][49]  ( .D(n9766), .CK(clk), .RN(n4290), .Q(
        \I_cache/cache[6][49] ), .QN(n909) );
  DFFRX1 \I_cache/cache_reg[7][49]  ( .D(n9765), .CK(clk), .RN(n4290), .Q(
        \I_cache/cache[7][49] ), .QN(n1842) );
  DFFRX1 \I_cache/cache_reg[0][50]  ( .D(n9764), .CK(clk), .RN(n4290), .Q(
        \I_cache/cache[0][50] ), .QN(n791) );
  DFFRX1 \I_cache/cache_reg[1][50]  ( .D(n9763), .CK(clk), .RN(n4290), .Q(
        \I_cache/cache[1][50] ), .QN(n1724) );
  DFFRX1 \I_cache/cache_reg[2][50]  ( .D(n9762), .CK(clk), .RN(n4290), .Q(
        \I_cache/cache[2][50] ), .QN(n793) );
  DFFRX1 \I_cache/cache_reg[3][50]  ( .D(n9761), .CK(clk), .RN(n4290), .Q(
        \I_cache/cache[3][50] ), .QN(n1726) );
  DFFRX1 \I_cache/cache_reg[4][50]  ( .D(n9760), .CK(clk), .RN(n4291), .Q(
        \I_cache/cache[4][50] ), .QN(n792) );
  DFFRX1 \I_cache/cache_reg[5][50]  ( .D(n9759), .CK(clk), .RN(n4291), .Q(
        \I_cache/cache[5][50] ), .QN(n1725) );
  DFFRX1 \I_cache/cache_reg[6][50]  ( .D(n9758), .CK(clk), .RN(n4291), .Q(
        \I_cache/cache[6][50] ), .QN(n845) );
  DFFRX1 \I_cache/cache_reg[7][50]  ( .D(n9757), .CK(clk), .RN(n4291), .Q(
        \I_cache/cache[7][50] ), .QN(n1778) );
  DFFRX1 \I_cache/cache_reg[0][51]  ( .D(n9756), .CK(clk), .RN(n4291), .Q(
        \I_cache/cache[0][51] ), .QN(n767) );
  DFFRX1 \I_cache/cache_reg[1][51]  ( .D(n9755), .CK(clk), .RN(n4291), .Q(
        \I_cache/cache[1][51] ), .QN(n1700) );
  DFFRX1 \I_cache/cache_reg[2][51]  ( .D(n9754), .CK(clk), .RN(n4291), .Q(
        \I_cache/cache[2][51] ), .QN(n769) );
  DFFRX1 \I_cache/cache_reg[3][51]  ( .D(n9753), .CK(clk), .RN(n4291), .Q(
        \I_cache/cache[3][51] ), .QN(n1702) );
  DFFRX1 \I_cache/cache_reg[4][51]  ( .D(n9752), .CK(clk), .RN(n4291), .Q(
        \I_cache/cache[4][51] ), .QN(n768) );
  DFFRX1 \I_cache/cache_reg[5][51]  ( .D(n9751), .CK(clk), .RN(n4291), .Q(
        \I_cache/cache[5][51] ), .QN(n1701) );
  DFFRX1 \I_cache/cache_reg[6][51]  ( .D(n9750), .CK(clk), .RN(n4291), .Q(
        \I_cache/cache[6][51] ), .QN(n835) );
  DFFRX1 \I_cache/cache_reg[7][51]  ( .D(n9749), .CK(clk), .RN(n4291), .Q(
        \I_cache/cache[7][51] ), .QN(n1768) );
  DFFRX1 \I_cache/cache_reg[0][52]  ( .D(n9748), .CK(clk), .RN(n4292), .Q(
        \I_cache/cache[0][52] ), .QN(n1867) );
  DFFRX1 \I_cache/cache_reg[1][52]  ( .D(n9747), .CK(clk), .RN(n4292), .Q(
        \I_cache/cache[1][52] ), .QN(n933) );
  DFFRX1 \I_cache/cache_reg[2][52]  ( .D(n9746), .CK(clk), .RN(n4292), .Q(
        \I_cache/cache[2][52] ), .QN(n1868) );
  DFFRX1 \I_cache/cache_reg[3][52]  ( .D(n9745), .CK(clk), .RN(n4292), .Q(
        \I_cache/cache[3][52] ), .QN(n934) );
  DFFRX1 \I_cache/cache_reg[4][52]  ( .D(n9744), .CK(clk), .RN(n4292), .Q(
        \I_cache/cache[4][52] ), .QN(n865) );
  DFFRX1 \I_cache/cache_reg[5][52]  ( .D(n9743), .CK(clk), .RN(n4292), .Q(
        \I_cache/cache[5][52] ), .QN(n1798) );
  DFFRX1 \I_cache/cache_reg[6][52]  ( .D(n9742), .CK(clk), .RN(n4292), .Q(
        \I_cache/cache[6][52] ), .QN(n900) );
  DFFRX1 \I_cache/cache_reg[7][52]  ( .D(n9741), .CK(clk), .RN(n4292), .Q(
        \I_cache/cache[7][52] ), .QN(n1833) );
  DFFRX1 \I_cache/cache_reg[0][53]  ( .D(n9740), .CK(clk), .RN(n4292), .Q(
        \I_cache/cache[0][53] ), .QN(n1853) );
  DFFRX1 \I_cache/cache_reg[1][53]  ( .D(n9739), .CK(clk), .RN(n4292), .Q(
        \I_cache/cache[1][53] ), .QN(n919) );
  DFFRX1 \I_cache/cache_reg[2][53]  ( .D(n9738), .CK(clk), .RN(n4292), .Q(
        \I_cache/cache[2][53] ), .QN(n787) );
  DFFRX1 \I_cache/cache_reg[3][53]  ( .D(n9737), .CK(clk), .RN(n4292), .Q(
        \I_cache/cache[3][53] ), .QN(n1720) );
  DFFRX1 \I_cache/cache_reg[4][53]  ( .D(n9736), .CK(clk), .RN(n4293), .Q(
        \I_cache/cache[4][53] ), .QN(n786) );
  DFFRX1 \I_cache/cache_reg[5][53]  ( .D(n9735), .CK(clk), .RN(n4293), .Q(
        \I_cache/cache[5][53] ), .QN(n1719) );
  DFFRX1 \I_cache/cache_reg[6][53]  ( .D(n9734), .CK(clk), .RN(n4293), .Q(
        \I_cache/cache[6][53] ), .QN(n843) );
  DFFRX1 \I_cache/cache_reg[7][53]  ( .D(n9733), .CK(clk), .RN(n4293), .Q(
        \I_cache/cache[7][53] ), .QN(n1776) );
  DFFRX1 \I_cache/cache_reg[0][54]  ( .D(n9732), .CK(clk), .RN(n4293), .Q(
        \I_cache/cache[0][54] ), .QN(n1872) );
  DFFRX1 \I_cache/cache_reg[1][54]  ( .D(n9731), .CK(clk), .RN(n4293), .Q(
        \I_cache/cache[1][54] ), .QN(n938) );
  DFFRX1 \I_cache/cache_reg[2][54]  ( .D(n9730), .CK(clk), .RN(n4293), .Q(
        \I_cache/cache[2][54] ), .QN(n1873) );
  DFFRX1 \I_cache/cache_reg[3][54]  ( .D(n9729), .CK(clk), .RN(n4293), .Q(
        \I_cache/cache[3][54] ), .QN(n939) );
  DFFRX1 \I_cache/cache_reg[4][54]  ( .D(n9728), .CK(clk), .RN(n4293), .Q(
        \I_cache/cache[4][54] ), .QN(n872) );
  DFFRX1 \I_cache/cache_reg[5][54]  ( .D(n9727), .CK(clk), .RN(n4293), .Q(
        \I_cache/cache[5][54] ), .QN(n1805) );
  DFFRX1 \I_cache/cache_reg[6][54]  ( .D(n9726), .CK(clk), .RN(n4293), .Q(
        \I_cache/cache[6][54] ), .QN(n913) );
  DFFRX1 \I_cache/cache_reg[7][54]  ( .D(n9725), .CK(clk), .RN(n4293), .Q(
        \I_cache/cache[7][54] ), .QN(n1846) );
  DFFRX1 \I_cache/cache_reg[0][55]  ( .D(n9724), .CK(clk), .RN(n4294), .Q(
        \I_cache/cache[0][55] ), .QN(n1850) );
  DFFRX1 \I_cache/cache_reg[1][55]  ( .D(n9723), .CK(clk), .RN(n4294), .Q(
        \I_cache/cache[1][55] ), .QN(n916) );
  DFFRX1 \I_cache/cache_reg[2][55]  ( .D(n9722), .CK(clk), .RN(n4294), .Q(
        \I_cache/cache[2][55] ), .QN(n781) );
  DFFRX1 \I_cache/cache_reg[3][55]  ( .D(n9721), .CK(clk), .RN(n4294), .Q(
        \I_cache/cache[3][55] ), .QN(n1714) );
  DFFRX1 \I_cache/cache_reg[4][55]  ( .D(n9720), .CK(clk), .RN(n4294), .Q(
        \I_cache/cache[4][55] ), .QN(n780) );
  DFFRX1 \I_cache/cache_reg[5][55]  ( .D(n9719), .CK(clk), .RN(n4294), .Q(
        \I_cache/cache[5][55] ), .QN(n1713) );
  DFFRX1 \I_cache/cache_reg[6][55]  ( .D(n9718), .CK(clk), .RN(n4294), .Q(
        \I_cache/cache[6][55] ), .QN(n840) );
  DFFRX1 \I_cache/cache_reg[7][55]  ( .D(n9717), .CK(clk), .RN(n4294), .Q(
        \I_cache/cache[7][55] ), .QN(n1773) );
  DFFRX1 \I_cache/cache_reg[0][56]  ( .D(n9716), .CK(clk), .RN(n4294), .Q(
        \I_cache/cache[0][56] ), .QN(n1861) );
  DFFRX1 \I_cache/cache_reg[1][56]  ( .D(n9715), .CK(clk), .RN(n4294), .Q(
        \I_cache/cache[1][56] ), .QN(n927) );
  DFFRX1 \I_cache/cache_reg[2][56]  ( .D(n9714), .CK(clk), .RN(n4294), .Q(
        \I_cache/cache[2][56] ), .QN(n1863) );
  DFFRX1 \I_cache/cache_reg[3][56]  ( .D(n9713), .CK(clk), .RN(n4294), .Q(
        \I_cache/cache[3][56] ), .QN(n929) );
  DFFRX1 \I_cache/cache_reg[4][56]  ( .D(n9712), .CK(clk), .RN(n4295), .Q(
        \I_cache/cache[4][56] ), .QN(n1862) );
  DFFRX1 \I_cache/cache_reg[5][56]  ( .D(n9711), .CK(clk), .RN(n4295), .Q(
        \I_cache/cache[5][56] ), .QN(n928) );
  DFFRX1 \I_cache/cache_reg[6][56]  ( .D(n9710), .CK(clk), .RN(n4295), .Q(
        \I_cache/cache[6][56] ), .QN(n896) );
  DFFRX1 \I_cache/cache_reg[7][56]  ( .D(n9709), .CK(clk), .RN(n4295), .Q(
        \I_cache/cache[7][56] ), .QN(n1829) );
  DFFRX1 \I_cache/cache_reg[0][57]  ( .D(n9708), .CK(clk), .RN(n4295), .Q(
        \I_cache/cache[0][57] ), .QN(n1877) );
  DFFRX1 \I_cache/cache_reg[1][57]  ( .D(n9707), .CK(clk), .RN(n4295), .Q(
        \I_cache/cache[1][57] ), .QN(n943) );
  DFFRX1 \I_cache/cache_reg[2][57]  ( .D(n9706), .CK(clk), .RN(n4295), .Q(
        \I_cache/cache[2][57] ), .QN(n1878) );
  DFFRX1 \I_cache/cache_reg[3][57]  ( .D(n9705), .CK(clk), .RN(n4295), .Q(
        \I_cache/cache[3][57] ), .QN(n944) );
  DFFRX1 \I_cache/cache_reg[4][57]  ( .D(n9704), .CK(clk), .RN(n4295), .Q(
        \I_cache/cache[4][57] ), .QN(n879) );
  DFFRX1 \I_cache/cache_reg[5][57]  ( .D(n9703), .CK(clk), .RN(n4295), .Q(
        \I_cache/cache[5][57] ), .QN(n1812) );
  DFFRX1 \I_cache/cache_reg[6][57]  ( .D(n9702), .CK(clk), .RN(n4295), .Q(
        \I_cache/cache[6][57] ), .QN(n904) );
  DFFRX1 \I_cache/cache_reg[7][57]  ( .D(n9701), .CK(clk), .RN(n4295), .Q(
        \I_cache/cache[7][57] ), .QN(n1837) );
  DFFRX1 \I_cache/cache_reg[0][58]  ( .D(n9700), .CK(clk), .RN(n4296), .Q(
        \I_cache/cache[0][58] ), .QN(n701) );
  DFFRX1 \I_cache/cache_reg[1][58]  ( .D(n9699), .CK(clk), .RN(n4296), .Q(
        \I_cache/cache[1][58] ), .QN(n1634) );
  DFFRX1 \I_cache/cache_reg[2][58]  ( .D(n9698), .CK(clk), .RN(n4296), .Q(
        \I_cache/cache[2][58] ), .QN(n703) );
  DFFRX1 \I_cache/cache_reg[3][58]  ( .D(n9697), .CK(clk), .RN(n4296), .Q(
        \I_cache/cache[3][58] ), .QN(n1636) );
  DFFRX1 \I_cache/cache_reg[4][58]  ( .D(n9696), .CK(clk), .RN(n4296), .Q(
        \I_cache/cache[4][58] ), .QN(n702) );
  DFFRX1 \I_cache/cache_reg[5][58]  ( .D(n9695), .CK(clk), .RN(n4296), .Q(
        \I_cache/cache[5][58] ), .QN(n1635) );
  DFFRX1 \I_cache/cache_reg[6][58]  ( .D(n9694), .CK(clk), .RN(n4296), .Q(
        \I_cache/cache[6][58] ), .QN(n813) );
  DFFRX1 \I_cache/cache_reg[7][58]  ( .D(n9693), .CK(clk), .RN(n4296), .Q(
        \I_cache/cache[7][58] ), .QN(n1746) );
  DFFRX1 \I_cache/cache_reg[0][59]  ( .D(n9692), .CK(clk), .RN(n4296), .Q(
        \I_cache/cache[0][59] ), .QN(n758) );
  DFFRX1 \I_cache/cache_reg[1][59]  ( .D(n9691), .CK(clk), .RN(n4296), .Q(
        \I_cache/cache[1][59] ), .QN(n1691) );
  DFFRX1 \I_cache/cache_reg[2][59]  ( .D(n9690), .CK(clk), .RN(n4296), .Q(
        \I_cache/cache[2][59] ), .QN(n760) );
  DFFRX1 \I_cache/cache_reg[3][59]  ( .D(n9689), .CK(clk), .RN(n4296), .Q(
        \I_cache/cache[3][59] ), .QN(n1693) );
  DFFRX1 \I_cache/cache_reg[4][59]  ( .D(n9688), .CK(clk), .RN(n4297), .Q(
        \I_cache/cache[4][59] ), .QN(n759) );
  DFFRX1 \I_cache/cache_reg[5][59]  ( .D(n9687), .CK(clk), .RN(n4297), .Q(
        \I_cache/cache[5][59] ), .QN(n1692) );
  DFFRX1 \I_cache/cache_reg[6][59]  ( .D(n9686), .CK(clk), .RN(n4297), .Q(
        \I_cache/cache[6][59] ), .QN(n832) );
  DFFRX1 \I_cache/cache_reg[7][59]  ( .D(n9685), .CK(clk), .RN(n4297), .Q(
        \I_cache/cache[7][59] ), .QN(n1765) );
  DFFRX1 \I_cache/cache_reg[0][60]  ( .D(n9684), .CK(clk), .RN(n4297), .Q(
        \I_cache/cache[0][60] ), .QN(n746) );
  DFFRX1 \I_cache/cache_reg[1][60]  ( .D(n9683), .CK(clk), .RN(n4297), .Q(
        \I_cache/cache[1][60] ), .QN(n1679) );
  DFFRX1 \I_cache/cache_reg[2][60]  ( .D(n9682), .CK(clk), .RN(n4297), .Q(
        \I_cache/cache[2][60] ), .QN(n748) );
  DFFRX1 \I_cache/cache_reg[3][60]  ( .D(n9681), .CK(clk), .RN(n4297), .Q(
        \I_cache/cache[3][60] ), .QN(n1681) );
  DFFRX1 \I_cache/cache_reg[4][60]  ( .D(n9680), .CK(clk), .RN(n4297), .Q(
        \I_cache/cache[4][60] ), .QN(n747) );
  DFFRX1 \I_cache/cache_reg[5][60]  ( .D(n9679), .CK(clk), .RN(n4297), .Q(
        \I_cache/cache[5][60] ), .QN(n1680) );
  DFFRX1 \I_cache/cache_reg[6][60]  ( .D(n9678), .CK(clk), .RN(n4297), .Q(
        \I_cache/cache[6][60] ), .QN(n828) );
  DFFRX1 \I_cache/cache_reg[7][60]  ( .D(n9677), .CK(clk), .RN(n4297), .Q(
        \I_cache/cache[7][60] ), .QN(n1761) );
  DFFRX1 \I_cache/cache_reg[0][61]  ( .D(n9676), .CK(clk), .RN(n4298), .Q(
        \I_cache/cache[0][61] ), .QN(n716) );
  DFFRX1 \I_cache/cache_reg[1][61]  ( .D(n9675), .CK(clk), .RN(n4298), .Q(
        \I_cache/cache[1][61] ), .QN(n1649) );
  DFFRX1 \I_cache/cache_reg[2][61]  ( .D(n9674), .CK(clk), .RN(n4298), .Q(
        \I_cache/cache[2][61] ), .QN(n718) );
  DFFRX1 \I_cache/cache_reg[3][61]  ( .D(n9673), .CK(clk), .RN(n4298), .Q(
        \I_cache/cache[3][61] ), .QN(n1651) );
  DFFRX1 \I_cache/cache_reg[4][61]  ( .D(n9672), .CK(clk), .RN(n4298), .Q(
        \I_cache/cache[4][61] ), .QN(n717) );
  DFFRX1 \I_cache/cache_reg[5][61]  ( .D(n9671), .CK(clk), .RN(n4298), .Q(
        \I_cache/cache[5][61] ), .QN(n1650) );
  DFFRX1 \I_cache/cache_reg[6][61]  ( .D(n9670), .CK(clk), .RN(n4298), .Q(
        \I_cache/cache[6][61] ), .QN(n818) );
  DFFRX1 \I_cache/cache_reg[7][61]  ( .D(n9669), .CK(clk), .RN(n4298), .Q(
        \I_cache/cache[7][61] ), .QN(n1751) );
  DFFRX1 \I_cache/cache_reg[0][62]  ( .D(n9668), .CK(clk), .RN(n4298), .Q(
        \I_cache/cache[0][62] ), .QN(n737) );
  DFFRX1 \I_cache/cache_reg[1][62]  ( .D(n9667), .CK(clk), .RN(n4298), .Q(
        \I_cache/cache[1][62] ), .QN(n1670) );
  DFFRX1 \I_cache/cache_reg[2][62]  ( .D(n9666), .CK(clk), .RN(n4298), .Q(
        \I_cache/cache[2][62] ), .QN(n739) );
  DFFRX1 \I_cache/cache_reg[3][62]  ( .D(n9665), .CK(clk), .RN(n4298), .Q(
        \I_cache/cache[3][62] ), .QN(n1672) );
  DFFRX1 \I_cache/cache_reg[4][62]  ( .D(n9664), .CK(clk), .RN(n4299), .Q(
        \I_cache/cache[4][62] ), .QN(n738) );
  DFFRX1 \I_cache/cache_reg[5][62]  ( .D(n9663), .CK(clk), .RN(n4299), .Q(
        \I_cache/cache[5][62] ), .QN(n1671) );
  DFFRX1 \I_cache/cache_reg[6][62]  ( .D(n9662), .CK(clk), .RN(n4299), .Q(
        \I_cache/cache[6][62] ), .QN(n825) );
  DFFRX1 \I_cache/cache_reg[7][62]  ( .D(n9661), .CK(clk), .RN(n4299), .Q(
        \I_cache/cache[7][62] ), .QN(n1758) );
  DFFRX1 \I_cache/cache_reg[0][63]  ( .D(n9660), .CK(clk), .RN(n4299), .Q(
        \I_cache/cache[0][63] ), .QN(n725) );
  DFFRX1 \I_cache/cache_reg[1][63]  ( .D(n9659), .CK(clk), .RN(n4299), .Q(
        \I_cache/cache[1][63] ), .QN(n1658) );
  DFFRX1 \I_cache/cache_reg[2][63]  ( .D(n9658), .CK(clk), .RN(n4299), .Q(
        \I_cache/cache[2][63] ), .QN(n727) );
  DFFRX1 \I_cache/cache_reg[3][63]  ( .D(n9657), .CK(clk), .RN(n4299), .Q(
        \I_cache/cache[3][63] ), .QN(n1660) );
  DFFRX1 \I_cache/cache_reg[4][63]  ( .D(n9656), .CK(clk), .RN(n4299), .Q(
        \I_cache/cache[4][63] ), .QN(n726) );
  DFFRX1 \I_cache/cache_reg[5][63]  ( .D(n9655), .CK(clk), .RN(n4299), .Q(
        \I_cache/cache[5][63] ), .QN(n1659) );
  DFFRX1 \I_cache/cache_reg[6][63]  ( .D(n9654), .CK(clk), .RN(n4299), .Q(
        \I_cache/cache[6][63] ), .QN(n821) );
  DFFRX1 \I_cache/cache_reg[7][63]  ( .D(n9653), .CK(clk), .RN(n4299), .Q(
        \I_cache/cache[7][63] ), .QN(n1754) );
  DFFRX1 \I_cache/cache_reg[0][74]  ( .D(n9572), .CK(clk), .RN(n4306), .Q(
        \I_cache/cache[0][74] ), .QN(n623) );
  DFFRX1 \I_cache/cache_reg[0][80]  ( .D(n9524), .CK(clk), .RN(n4310), .Q(
        \I_cache/cache[0][80] ), .QN(n801) );
  DFFRX1 \I_cache/cache_reg[1][80]  ( .D(n9523), .CK(clk), .RN(n4310), .Q(
        \I_cache/cache[1][80] ), .QN(n1734) );
  DFFRX1 \I_cache/cache_reg[2][80]  ( .D(n9522), .CK(clk), .RN(n4310), .Q(
        \I_cache/cache[2][80] ), .QN(n803) );
  DFFRX1 \I_cache/cache_reg[3][80]  ( .D(n9521), .CK(clk), .RN(n4310), .Q(
        \I_cache/cache[3][80] ), .QN(n1736) );
  DFFRX1 \I_cache/cache_reg[4][80]  ( .D(n9520), .CK(clk), .RN(n4311), .Q(
        \I_cache/cache[4][80] ), .QN(n802) );
  DFFRX1 \I_cache/cache_reg[5][80]  ( .D(n9519), .CK(clk), .RN(n4311), .Q(
        \I_cache/cache[5][80] ), .QN(n1735) );
  DFFRX1 \I_cache/cache_reg[6][80]  ( .D(n9518), .CK(clk), .RN(n4311), .Q(
        \I_cache/cache[6][80] ), .QN(n849) );
  DFFRX1 \I_cache/cache_reg[7][80]  ( .D(n9517), .CK(clk), .RN(n4311), .Q(
        \I_cache/cache[7][80] ), .QN(n1782) );
  DFFRX1 \I_cache/cache_reg[0][81]  ( .D(n9516), .CK(clk), .RN(n4311), .Q(
        \I_cache/cache[0][81] ), .QN(n798) );
  DFFRX1 \I_cache/cache_reg[1][81]  ( .D(n9515), .CK(clk), .RN(n4311), .Q(
        \I_cache/cache[1][81] ), .QN(n1731) );
  DFFRX1 \I_cache/cache_reg[2][81]  ( .D(n9514), .CK(clk), .RN(n4311), .Q(
        \I_cache/cache[2][81] ), .QN(n800) );
  DFFRX1 \I_cache/cache_reg[3][81]  ( .D(n9513), .CK(clk), .RN(n4311), .Q(
        \I_cache/cache[3][81] ), .QN(n1733) );
  DFFRX1 \I_cache/cache_reg[4][81]  ( .D(n9512), .CK(clk), .RN(n4311), .Q(
        \I_cache/cache[4][81] ), .QN(n799) );
  DFFRX1 \I_cache/cache_reg[5][81]  ( .D(n9511), .CK(clk), .RN(n4311), .Q(
        \I_cache/cache[5][81] ), .QN(n1732) );
  DFFRX1 \I_cache/cache_reg[6][81]  ( .D(n9510), .CK(clk), .RN(n4311), .Q(
        \I_cache/cache[6][81] ), .QN(n848) );
  DFFRX1 \I_cache/cache_reg[7][81]  ( .D(n9509), .CK(clk), .RN(n4311), .Q(
        \I_cache/cache[7][81] ), .QN(n1781) );
  DFFRX1 \I_cache/cache_reg[0][82]  ( .D(n9508), .CK(clk), .RN(n4312), .Q(
        \I_cache/cache[0][82] ), .QN(n788) );
  DFFRX1 \I_cache/cache_reg[1][82]  ( .D(n9507), .CK(clk), .RN(n4312), .Q(
        \I_cache/cache[1][82] ), .QN(n1721) );
  DFFRX1 \I_cache/cache_reg[2][82]  ( .D(n9506), .CK(clk), .RN(n4312), .Q(
        \I_cache/cache[2][82] ), .QN(n790) );
  DFFRX1 \I_cache/cache_reg[3][82]  ( .D(n9505), .CK(clk), .RN(n4312), .Q(
        \I_cache/cache[3][82] ), .QN(n1723) );
  DFFRX1 \I_cache/cache_reg[4][82]  ( .D(n9504), .CK(clk), .RN(n4312), .Q(
        \I_cache/cache[4][82] ), .QN(n789) );
  DFFRX1 \I_cache/cache_reg[5][82]  ( .D(n9503), .CK(clk), .RN(n4312), .Q(
        \I_cache/cache[5][82] ), .QN(n1722) );
  DFFRX1 \I_cache/cache_reg[6][82]  ( .D(n9502), .CK(clk), .RN(n4312), .Q(
        \I_cache/cache[6][82] ), .QN(n844) );
  DFFRX1 \I_cache/cache_reg[7][82]  ( .D(n9501), .CK(clk), .RN(n4312), .Q(
        \I_cache/cache[7][82] ), .QN(n1777) );
  DFFRX1 \I_cache/cache_reg[0][83]  ( .D(n9500), .CK(clk), .RN(n4312), .Q(
        \I_cache/cache[0][83] ), .QN(n764) );
  DFFRX1 \I_cache/cache_reg[1][83]  ( .D(n9499), .CK(clk), .RN(n4312), .Q(
        \I_cache/cache[1][83] ), .QN(n1697) );
  DFFRX1 \I_cache/cache_reg[2][83]  ( .D(n9498), .CK(clk), .RN(n4312), .Q(
        \I_cache/cache[2][83] ), .QN(n766) );
  DFFRX1 \I_cache/cache_reg[3][83]  ( .D(n9497), .CK(clk), .RN(n4312), .Q(
        \I_cache/cache[3][83] ), .QN(n1699) );
  DFFRX1 \I_cache/cache_reg[4][83]  ( .D(n9496), .CK(clk), .RN(n4313), .Q(
        \I_cache/cache[4][83] ), .QN(n765) );
  DFFRX1 \I_cache/cache_reg[5][83]  ( .D(n9495), .CK(clk), .RN(n4313), .Q(
        \I_cache/cache[5][83] ), .QN(n1698) );
  DFFRX1 \I_cache/cache_reg[6][83]  ( .D(n9494), .CK(clk), .RN(n4313), .Q(
        \I_cache/cache[6][83] ), .QN(n834) );
  DFFRX1 \I_cache/cache_reg[7][83]  ( .D(n9493), .CK(clk), .RN(n4313), .Q(
        \I_cache/cache[7][83] ), .QN(n1767) );
  DFFRX1 \I_cache/cache_reg[0][84]  ( .D(n9492), .CK(clk), .RN(n4313), .Q(
        \I_cache/cache[0][84] ), .QN(n862) );
  DFFRX1 \I_cache/cache_reg[1][84]  ( .D(n9491), .CK(clk), .RN(n4313), .Q(
        \I_cache/cache[1][84] ), .QN(n1795) );
  DFFRX1 \I_cache/cache_reg[2][84]  ( .D(n9490), .CK(clk), .RN(n4313), .Q(
        \I_cache/cache[2][84] ), .QN(n864) );
  DFFRX1 \I_cache/cache_reg[3][84]  ( .D(n9489), .CK(clk), .RN(n4313), .Q(
        \I_cache/cache[3][84] ), .QN(n1797) );
  DFFRX1 \I_cache/cache_reg[4][84]  ( .D(n9488), .CK(clk), .RN(n4313), .Q(
        \I_cache/cache[4][84] ), .QN(n863) );
  DFFRX1 \I_cache/cache_reg[5][84]  ( .D(n9487), .CK(clk), .RN(n4313), .Q(
        \I_cache/cache[5][84] ), .QN(n1796) );
  DFFRX1 \I_cache/cache_reg[6][84]  ( .D(n9486), .CK(clk), .RN(n4313), .Q(
        \I_cache/cache[6][84] ), .QN(n899) );
  DFFRX1 \I_cache/cache_reg[7][84]  ( .D(n9485), .CK(clk), .RN(n4313), .Q(
        \I_cache/cache[7][84] ), .QN(n1832) );
  DFFRX1 \I_cache/cache_reg[0][85]  ( .D(n9484), .CK(clk), .RN(n4314), .Q(
        \I_cache/cache[0][85] ), .QN(n882) );
  DFFRX1 \I_cache/cache_reg[1][85]  ( .D(n9483), .CK(clk), .RN(n4314), .Q(
        \I_cache/cache[1][85] ), .QN(n1815) );
  DFFRX1 \I_cache/cache_reg[2][85]  ( .D(n9482), .CK(clk), .RN(n4314), .Q(
        \I_cache/cache[2][85] ), .QN(n884) );
  DFFRX1 \I_cache/cache_reg[3][85]  ( .D(n9481), .CK(clk), .RN(n4314), .Q(
        \I_cache/cache[3][85] ), .QN(n1817) );
  DFFRX1 \I_cache/cache_reg[4][85]  ( .D(n9480), .CK(clk), .RN(n4314), .Q(
        \I_cache/cache[4][85] ), .QN(n883) );
  DFFRX1 \I_cache/cache_reg[5][85]  ( .D(n9479), .CK(clk), .RN(n4314), .Q(
        \I_cache/cache[5][85] ), .QN(n1816) );
  DFFRX1 \I_cache/cache_reg[6][85]  ( .D(n9478), .CK(clk), .RN(n4314), .Q(
        \I_cache/cache[6][85] ), .QN(n906) );
  DFFRX1 \I_cache/cache_reg[7][85]  ( .D(n9477), .CK(clk), .RN(n4314), .Q(
        \I_cache/cache[7][85] ), .QN(n1839) );
  DFFRX1 \I_cache/cache_reg[0][86]  ( .D(n9476), .CK(clk), .RN(n4314), .Q(
        \I_cache/cache[0][86] ), .QN(n869) );
  DFFRX1 \I_cache/cache_reg[1][86]  ( .D(n9475), .CK(clk), .RN(n4314), .Q(
        \I_cache/cache[1][86] ), .QN(n1802) );
  DFFRX1 \I_cache/cache_reg[2][86]  ( .D(n9474), .CK(clk), .RN(n4314), .Q(
        \I_cache/cache[2][86] ), .QN(n871) );
  DFFRX1 \I_cache/cache_reg[3][86]  ( .D(n9473), .CK(clk), .RN(n4314), .Q(
        \I_cache/cache[3][86] ), .QN(n1804) );
  DFFRX1 \I_cache/cache_reg[4][86]  ( .D(n9472), .CK(clk), .RN(n4315), .Q(
        \I_cache/cache[4][86] ), .QN(n870) );
  DFFRX1 \I_cache/cache_reg[5][86]  ( .D(n9471), .CK(clk), .RN(n4315), .Q(
        \I_cache/cache[5][86] ), .QN(n1803) );
  DFFRX1 \I_cache/cache_reg[6][86]  ( .D(n9470), .CK(clk), .RN(n4315), .Q(
        \I_cache/cache[6][86] ), .QN(n912) );
  DFFRX1 \I_cache/cache_reg[7][86]  ( .D(n9469), .CK(clk), .RN(n4315), .Q(
        \I_cache/cache[7][86] ), .QN(n1845) );
  DFFRX1 \I_cache/cache_reg[0][87]  ( .D(n9468), .CK(clk), .RN(n4315), .Q(
        \I_cache/cache[0][87] ), .QN(n777) );
  DFFRX1 \I_cache/cache_reg[1][87]  ( .D(n9467), .CK(clk), .RN(n4315), .Q(
        \I_cache/cache[1][87] ), .QN(n1710) );
  DFFRX1 \I_cache/cache_reg[2][87]  ( .D(n9466), .CK(clk), .RN(n4315), .Q(
        \I_cache/cache[2][87] ), .QN(n779) );
  DFFRX1 \I_cache/cache_reg[3][87]  ( .D(n9465), .CK(clk), .RN(n4315), .Q(
        \I_cache/cache[3][87] ), .QN(n1712) );
  DFFRX1 \I_cache/cache_reg[4][87]  ( .D(n9464), .CK(clk), .RN(n4315), .Q(
        \I_cache/cache[4][87] ), .QN(n778) );
  DFFRX1 \I_cache/cache_reg[5][87]  ( .D(n9463), .CK(clk), .RN(n4315), .Q(
        \I_cache/cache[5][87] ), .QN(n1711) );
  DFFRX1 \I_cache/cache_reg[6][87]  ( .D(n9462), .CK(clk), .RN(n4315), .Q(
        \I_cache/cache[6][87] ), .QN(n839) );
  DFFRX1 \I_cache/cache_reg[7][87]  ( .D(n9461), .CK(clk), .RN(n4315), .Q(
        \I_cache/cache[7][87] ), .QN(n1772) );
  DFFRX1 \I_cache/cache_reg[0][88]  ( .D(n9460), .CK(clk), .RN(n4316), .Q(
        \I_cache/cache[0][88] ), .QN(n856) );
  DFFRX1 \I_cache/cache_reg[1][88]  ( .D(n9459), .CK(clk), .RN(n4316), .Q(
        \I_cache/cache[1][88] ), .QN(n1789) );
  DFFRX1 \I_cache/cache_reg[2][88]  ( .D(n9458), .CK(clk), .RN(n4316), .Q(
        \I_cache/cache[2][88] ), .QN(n858) );
  DFFRX1 \I_cache/cache_reg[3][88]  ( .D(n9457), .CK(clk), .RN(n4316), .Q(
        \I_cache/cache[3][88] ), .QN(n1791) );
  DFFRX1 \I_cache/cache_reg[4][88]  ( .D(n9456), .CK(clk), .RN(n4316), .Q(
        \I_cache/cache[4][88] ), .QN(n857) );
  DFFRX1 \I_cache/cache_reg[5][88]  ( .D(n9455), .CK(clk), .RN(n4316), .Q(
        \I_cache/cache[5][88] ), .QN(n1790) );
  DFFRX1 \I_cache/cache_reg[6][88]  ( .D(n9454), .CK(clk), .RN(n4316), .Q(
        \I_cache/cache[6][88] ), .QN(n895) );
  DFFRX1 \I_cache/cache_reg[7][88]  ( .D(n9453), .CK(clk), .RN(n4316), .Q(
        \I_cache/cache[7][88] ), .QN(n1828) );
  DFFRX1 \I_cache/cache_reg[0][89]  ( .D(n9452), .CK(clk), .RN(n4316), .Q(
        \I_cache/cache[0][89] ), .QN(n876) );
  DFFRX1 \I_cache/cache_reg[1][89]  ( .D(n9451), .CK(clk), .RN(n4316), .Q(
        \I_cache/cache[1][89] ), .QN(n1809) );
  DFFRX1 \I_cache/cache_reg[2][89]  ( .D(n9450), .CK(clk), .RN(n4316), .Q(
        \I_cache/cache[2][89] ), .QN(n878) );
  DFFRX1 \I_cache/cache_reg[3][89]  ( .D(n9449), .CK(clk), .RN(n4316), .Q(
        \I_cache/cache[3][89] ), .QN(n1811) );
  DFFRX1 \I_cache/cache_reg[4][89]  ( .D(n9448), .CK(clk), .RN(n4317), .Q(
        \I_cache/cache[4][89] ), .QN(n877) );
  DFFRX1 \I_cache/cache_reg[5][89]  ( .D(n9447), .CK(clk), .RN(n4317), .Q(
        \I_cache/cache[5][89] ), .QN(n1810) );
  DFFRX1 \I_cache/cache_reg[6][89]  ( .D(n9446), .CK(clk), .RN(n4317), .Q(
        \I_cache/cache[6][89] ), .QN(n903) );
  DFFRX1 \I_cache/cache_reg[7][89]  ( .D(n9445), .CK(clk), .RN(n4317), .Q(
        \I_cache/cache[7][89] ), .QN(n1836) );
  DFFRX1 \I_cache/cache_reg[0][90]  ( .D(n9444), .CK(clk), .RN(n4317), .Q(
        \I_cache/cache[0][90] ), .QN(n698) );
  DFFRX1 \I_cache/cache_reg[1][90]  ( .D(n9443), .CK(clk), .RN(n4317), .Q(
        \I_cache/cache[1][90] ), .QN(n1631) );
  DFFRX1 \I_cache/cache_reg[2][90]  ( .D(n9442), .CK(clk), .RN(n4317), .Q(
        \I_cache/cache[2][90] ), .QN(n700) );
  DFFRX1 \I_cache/cache_reg[3][90]  ( .D(n9441), .CK(clk), .RN(n4317), .Q(
        \I_cache/cache[3][90] ), .QN(n1633) );
  DFFRX1 \I_cache/cache_reg[4][90]  ( .D(n9440), .CK(clk), .RN(n4317), .Q(
        \I_cache/cache[4][90] ), .QN(n699) );
  DFFRX1 \I_cache/cache_reg[5][90]  ( .D(n9439), .CK(clk), .RN(n4317), .Q(
        \I_cache/cache[5][90] ), .QN(n1632) );
  DFFRX1 \I_cache/cache_reg[6][90]  ( .D(n9438), .CK(clk), .RN(n4317), .Q(
        \I_cache/cache[6][90] ), .QN(n812) );
  DFFRX1 \I_cache/cache_reg[7][90]  ( .D(n9437), .CK(clk), .RN(n4317), .Q(
        \I_cache/cache[7][90] ), .QN(n1745) );
  DFFRX1 \I_cache/cache_reg[0][91]  ( .D(n9436), .CK(clk), .RN(n4318), .Q(
        \I_cache/cache[0][91] ), .QN(n755) );
  DFFRX1 \I_cache/cache_reg[1][91]  ( .D(n9435), .CK(clk), .RN(n4318), .Q(
        \I_cache/cache[1][91] ), .QN(n1688) );
  DFFRX1 \I_cache/cache_reg[2][91]  ( .D(n9434), .CK(clk), .RN(n4318), .Q(
        \I_cache/cache[2][91] ), .QN(n757) );
  DFFRX1 \I_cache/cache_reg[3][91]  ( .D(n9433), .CK(clk), .RN(n4318), .Q(
        \I_cache/cache[3][91] ), .QN(n1690) );
  DFFRX1 \I_cache/cache_reg[4][91]  ( .D(n9432), .CK(clk), .RN(n4318), .Q(
        \I_cache/cache[4][91] ), .QN(n756) );
  DFFRX1 \I_cache/cache_reg[5][91]  ( .D(n9431), .CK(clk), .RN(n4318), .Q(
        \I_cache/cache[5][91] ), .QN(n1689) );
  DFFRX1 \I_cache/cache_reg[6][91]  ( .D(n9430), .CK(clk), .RN(n4318), .Q(
        \I_cache/cache[6][91] ), .QN(n831) );
  DFFRX1 \I_cache/cache_reg[7][91]  ( .D(n9429), .CK(clk), .RN(n4318), .Q(
        \I_cache/cache[7][91] ), .QN(n1764) );
  DFFRX1 \I_cache/cache_reg[0][92]  ( .D(n9428), .CK(clk), .RN(n4318), .Q(
        \I_cache/cache[0][92] ), .QN(n743) );
  DFFRX1 \I_cache/cache_reg[1][92]  ( .D(n9427), .CK(clk), .RN(n4318), .Q(
        \I_cache/cache[1][92] ), .QN(n1676) );
  DFFRX1 \I_cache/cache_reg[2][92]  ( .D(n9426), .CK(clk), .RN(n4318), .Q(
        \I_cache/cache[2][92] ), .QN(n745) );
  DFFRX1 \I_cache/cache_reg[3][92]  ( .D(n9425), .CK(clk), .RN(n4318), .Q(
        \I_cache/cache[3][92] ), .QN(n1678) );
  DFFRX1 \I_cache/cache_reg[4][92]  ( .D(n9424), .CK(clk), .RN(n4319), .Q(
        \I_cache/cache[4][92] ), .QN(n744) );
  DFFRX1 \I_cache/cache_reg[5][92]  ( .D(n9423), .CK(clk), .RN(n4319), .Q(
        \I_cache/cache[5][92] ), .QN(n1677) );
  DFFRX1 \I_cache/cache_reg[6][92]  ( .D(n9422), .CK(clk), .RN(n4319), .Q(
        \I_cache/cache[6][92] ), .QN(n827) );
  DFFRX1 \I_cache/cache_reg[7][92]  ( .D(n9421), .CK(clk), .RN(n4319), .Q(
        \I_cache/cache[7][92] ), .QN(n1760) );
  DFFRX1 \I_cache/cache_reg[0][93]  ( .D(n9420), .CK(clk), .RN(n4319), .Q(
        \I_cache/cache[0][93] ), .QN(n713) );
  DFFRX1 \I_cache/cache_reg[1][93]  ( .D(n9419), .CK(clk), .RN(n4319), .Q(
        \I_cache/cache[1][93] ), .QN(n1646) );
  DFFRX1 \I_cache/cache_reg[2][93]  ( .D(n9418), .CK(clk), .RN(n4319), .Q(
        \I_cache/cache[2][93] ), .QN(n715) );
  DFFRX1 \I_cache/cache_reg[3][93]  ( .D(n9417), .CK(clk), .RN(n4319), .Q(
        \I_cache/cache[3][93] ), .QN(n1648) );
  DFFRX1 \I_cache/cache_reg[4][93]  ( .D(n9416), .CK(clk), .RN(n4319), .Q(
        \I_cache/cache[4][93] ), .QN(n714) );
  DFFRX1 \I_cache/cache_reg[5][93]  ( .D(n9415), .CK(clk), .RN(n4319), .Q(
        \I_cache/cache[5][93] ), .QN(n1647) );
  DFFRX1 \I_cache/cache_reg[6][93]  ( .D(n9414), .CK(clk), .RN(n4319), .Q(
        \I_cache/cache[6][93] ), .QN(n817) );
  DFFRX1 \I_cache/cache_reg[7][93]  ( .D(n9413), .CK(clk), .RN(n4319), .Q(
        \I_cache/cache[7][93] ), .QN(n1750) );
  DFFRX1 \I_cache/cache_reg[0][94]  ( .D(n9412), .CK(clk), .RN(n4320), .Q(
        \I_cache/cache[0][94] ), .QN(n734) );
  DFFRX1 \I_cache/cache_reg[1][94]  ( .D(n9411), .CK(clk), .RN(n4320), .Q(
        \I_cache/cache[1][94] ), .QN(n1667) );
  DFFRX1 \I_cache/cache_reg[2][94]  ( .D(n9410), .CK(clk), .RN(n4320), .Q(
        \I_cache/cache[2][94] ), .QN(n736) );
  DFFRX1 \I_cache/cache_reg[3][94]  ( .D(n9409), .CK(clk), .RN(n4320), .Q(
        \I_cache/cache[3][94] ), .QN(n1669) );
  DFFRX1 \I_cache/cache_reg[4][94]  ( .D(n9408), .CK(clk), .RN(n4320), .Q(
        \I_cache/cache[4][94] ), .QN(n735) );
  DFFRX1 \I_cache/cache_reg[5][94]  ( .D(n9407), .CK(clk), .RN(n4320), .Q(
        \I_cache/cache[5][94] ), .QN(n1668) );
  DFFRX1 \I_cache/cache_reg[6][94]  ( .D(n9406), .CK(clk), .RN(n4320), .Q(
        \I_cache/cache[6][94] ), .QN(n824) );
  DFFRX1 \I_cache/cache_reg[7][94]  ( .D(n9405), .CK(clk), .RN(n4320), .Q(
        \I_cache/cache[7][94] ), .QN(n1757) );
  DFFRX1 \I_cache/cache_reg[0][95]  ( .D(n9404), .CK(clk), .RN(n4320), .Q(
        \I_cache/cache[0][95] ), .QN(n637) );
  DFFRX1 \I_cache/cache_reg[1][95]  ( .D(n9403), .CK(clk), .RN(n4320), .Q(
        \I_cache/cache[1][95] ), .QN(n1556) );
  DFFRX1 \I_cache/cache_reg[2][95]  ( .D(n9402), .CK(clk), .RN(n4320), .Q(
        \I_cache/cache[2][95] ), .QN(n639) );
  DFFRX1 \I_cache/cache_reg[3][95]  ( .D(n9401), .CK(clk), .RN(n4320), .Q(
        \I_cache/cache[3][95] ), .QN(n1558) );
  DFFRX1 \I_cache/cache_reg[4][95]  ( .D(n9400), .CK(clk), .RN(n4321), .Q(
        \I_cache/cache[4][95] ), .QN(n638) );
  DFFRX1 \I_cache/cache_reg[5][95]  ( .D(n9399), .CK(clk), .RN(n4321), .Q(
        \I_cache/cache[5][95] ), .QN(n1557) );
  DFFRX1 \I_cache/cache_reg[6][95]  ( .D(n9398), .CK(clk), .RN(n4321), .Q(
        \I_cache/cache[6][95] ), .QN(n678) );
  DFFRX1 \I_cache/cache_reg[7][95]  ( .D(n9397), .CK(clk), .RN(n4321), .Q(
        \I_cache/cache[7][95] ), .QN(n1597) );
  DFFRX1 \I_cache/cache_reg[0][106]  ( .D(n9316), .CK(clk), .RN(n4328), .Q(
        \I_cache/cache[0][106] ), .QN(n626) );
  DFFRX1 \I_cache/cache_reg[2][106]  ( .D(n9314), .CK(clk), .RN(n4328), .Q(
        \I_cache/cache[2][106] ), .QN(n625) );
  DFFRX1 \I_cache/cache_reg[0][112]  ( .D(n9268), .CK(clk), .RN(n4332), .Q(
        \I_cache/cache[0][112] ), .QN(n807) );
  DFFRX1 \I_cache/cache_reg[1][112]  ( .D(n9267), .CK(clk), .RN(n4332), .Q(
        \I_cache/cache[1][112] ), .QN(n1740) );
  DFFRX1 \I_cache/cache_reg[2][112]  ( .D(n9266), .CK(clk), .RN(n4332), .Q(
        \I_cache/cache[2][112] ), .QN(n809) );
  DFFRX1 \I_cache/cache_reg[3][112]  ( .D(n9265), .CK(clk), .RN(n4332), .Q(
        \I_cache/cache[3][112] ), .QN(n1742) );
  DFFRX1 \I_cache/cache_reg[4][112]  ( .D(n9264), .CK(clk), .RN(n4332), .Q(
        \I_cache/cache[4][112] ), .QN(n808) );
  DFFRX1 \I_cache/cache_reg[5][112]  ( .D(n9263), .CK(clk), .RN(n4332), .Q(
        \I_cache/cache[5][112] ), .QN(n1741) );
  DFFRX1 \I_cache/cache_reg[6][112]  ( .D(n9262), .CK(clk), .RN(n4332), .Q(
        \I_cache/cache[6][112] ), .QN(n851) );
  DFFRX1 \I_cache/cache_reg[7][112]  ( .D(n9261), .CK(clk), .RN(n4332), .Q(
        \I_cache/cache[7][112] ), .QN(n1784) );
  DFFRX1 \I_cache/cache_reg[0][113]  ( .D(n9260), .CK(clk), .RN(n4332), .Q(
        \I_cache/cache[0][113] ), .QN(n885) );
  DFFRX1 \I_cache/cache_reg[1][113]  ( .D(n9259), .CK(clk), .RN(n4332), .Q(
        \I_cache/cache[1][113] ), .QN(n1818) );
  DFFRX1 \I_cache/cache_reg[2][113]  ( .D(n9258), .CK(clk), .RN(n4332), .Q(
        \I_cache/cache[2][113] ), .QN(n887) );
  DFFRX1 \I_cache/cache_reg[3][113]  ( .D(n9257), .CK(clk), .RN(n4332), .Q(
        \I_cache/cache[3][113] ), .QN(n1820) );
  DFFRX1 \I_cache/cache_reg[4][113]  ( .D(n9256), .CK(clk), .RN(n4333), .Q(
        \I_cache/cache[4][113] ), .QN(n886) );
  DFFRX1 \I_cache/cache_reg[5][113]  ( .D(n9255), .CK(clk), .RN(n4333), .Q(
        \I_cache/cache[5][113] ), .QN(n1819) );
  DFFRX1 \I_cache/cache_reg[6][113]  ( .D(n9254), .CK(clk), .RN(n4333), .Q(
        \I_cache/cache[6][113] ), .QN(n907) );
  DFFRX1 \I_cache/cache_reg[7][113]  ( .D(n9253), .CK(clk), .RN(n4333), .Q(
        \I_cache/cache[7][113] ), .QN(n1840) );
  DFFRX1 \I_cache/cache_reg[0][114]  ( .D(n9252), .CK(clk), .RN(n4333), .Q(
        \I_cache/cache[0][114] ), .QN(n794) );
  DFFRX1 \I_cache/cache_reg[1][114]  ( .D(n9251), .CK(clk), .RN(n4333), .Q(
        \I_cache/cache[1][114] ), .QN(n1727) );
  DFFRX1 \I_cache/cache_reg[2][114]  ( .D(n9250), .CK(clk), .RN(n4333), .Q(
        \I_cache/cache[2][114] ), .QN(n796) );
  DFFRX1 \I_cache/cache_reg[3][114]  ( .D(n9249), .CK(clk), .RN(n4333), .Q(
        \I_cache/cache[3][114] ), .QN(n1729) );
  DFFRX1 \I_cache/cache_reg[4][114]  ( .D(n9248), .CK(clk), .RN(n4333), .Q(
        \I_cache/cache[4][114] ), .QN(n795) );
  DFFRX1 \I_cache/cache_reg[5][114]  ( .D(n9247), .CK(clk), .RN(n4333), .Q(
        \I_cache/cache[5][114] ), .QN(n1728) );
  DFFRX1 \I_cache/cache_reg[6][114]  ( .D(n9246), .CK(clk), .RN(n4333), .Q(
        \I_cache/cache[6][114] ), .QN(n846) );
  DFFRX1 \I_cache/cache_reg[7][114]  ( .D(n9245), .CK(clk), .RN(n4333), .Q(
        \I_cache/cache[7][114] ), .QN(n1779) );
  DFFRX1 \I_cache/cache_reg[0][115]  ( .D(n9244), .CK(clk), .RN(n4334), .Q(
        \I_cache/cache[0][115] ), .QN(n770) );
  DFFRX1 \I_cache/cache_reg[1][115]  ( .D(n9243), .CK(clk), .RN(n4334), .Q(
        \I_cache/cache[1][115] ), .QN(n1703) );
  DFFRX1 \I_cache/cache_reg[2][115]  ( .D(n9242), .CK(clk), .RN(n4334), .Q(
        \I_cache/cache[2][115] ), .QN(n772) );
  DFFRX1 \I_cache/cache_reg[3][115]  ( .D(n9241), .CK(clk), .RN(n4334), .Q(
        \I_cache/cache[3][115] ), .QN(n1705) );
  DFFRX1 \I_cache/cache_reg[4][115]  ( .D(n9240), .CK(clk), .RN(n4334), .Q(
        \I_cache/cache[4][115] ), .QN(n771) );
  DFFRX1 \I_cache/cache_reg[5][115]  ( .D(n9239), .CK(clk), .RN(n4334), .Q(
        \I_cache/cache[5][115] ), .QN(n1704) );
  DFFRX1 \I_cache/cache_reg[6][115]  ( .D(n9238), .CK(clk), .RN(n4334), .Q(
        \I_cache/cache[6][115] ), .QN(n836) );
  DFFRX1 \I_cache/cache_reg[7][115]  ( .D(n9237), .CK(clk), .RN(n4334), .Q(
        \I_cache/cache[7][115] ), .QN(n1769) );
  DFFRX1 \I_cache/cache_reg[0][116]  ( .D(n9236), .CK(clk), .RN(n4334), .Q(
        \I_cache/cache[0][116] ), .QN(n859) );
  DFFRX1 \I_cache/cache_reg[1][116]  ( .D(n9235), .CK(clk), .RN(n4334), .Q(
        \I_cache/cache[1][116] ), .QN(n1792) );
  DFFRX1 \I_cache/cache_reg[2][116]  ( .D(n9234), .CK(clk), .RN(n4334), .Q(
        \I_cache/cache[2][116] ), .QN(n861) );
  DFFRX1 \I_cache/cache_reg[3][116]  ( .D(n9233), .CK(clk), .RN(n4334), .Q(
        \I_cache/cache[3][116] ), .QN(n1794) );
  DFFRX1 \I_cache/cache_reg[4][116]  ( .D(n9232), .CK(clk), .RN(n4335), .Q(
        \I_cache/cache[4][116] ), .QN(n860) );
  DFFRX1 \I_cache/cache_reg[5][116]  ( .D(n9231), .CK(clk), .RN(n4335), .Q(
        \I_cache/cache[5][116] ), .QN(n1793) );
  DFFRX1 \I_cache/cache_reg[6][116]  ( .D(n9230), .CK(clk), .RN(n4335), .Q(
        \I_cache/cache[6][116] ), .QN(n897) );
  DFFRX1 \I_cache/cache_reg[7][116]  ( .D(n9229), .CK(clk), .RN(n4335), .Q(
        \I_cache/cache[7][116] ), .QN(n1830) );
  DFFRX1 \I_cache/cache_reg[0][117]  ( .D(n9228), .CK(clk), .RN(n4335), .Q(
        \I_cache/cache[0][117] ), .QN(n782) );
  DFFRX1 \I_cache/cache_reg[1][117]  ( .D(n9227), .CK(clk), .RN(n4335), .Q(
        \I_cache/cache[1][117] ), .QN(n1715) );
  DFFRX1 \I_cache/cache_reg[2][117]  ( .D(n9226), .CK(clk), .RN(n4335), .Q(
        \I_cache/cache[2][117] ), .QN(n784) );
  DFFRX1 \I_cache/cache_reg[3][117]  ( .D(n9225), .CK(clk), .RN(n4335), .Q(
        \I_cache/cache[3][117] ), .QN(n1717) );
  DFFRX1 \I_cache/cache_reg[4][117]  ( .D(n9224), .CK(clk), .RN(n4335), .Q(
        \I_cache/cache[4][117] ), .QN(n783) );
  DFFRX1 \I_cache/cache_reg[5][117]  ( .D(n9223), .CK(clk), .RN(n4335), .Q(
        \I_cache/cache[5][117] ), .QN(n1716) );
  DFFRX1 \I_cache/cache_reg[6][117]  ( .D(n9222), .CK(clk), .RN(n4335), .Q(
        \I_cache/cache[6][117] ), .QN(n841) );
  DFFRX1 \I_cache/cache_reg[7][117]  ( .D(n9221), .CK(clk), .RN(n4335), .Q(
        \I_cache/cache[7][117] ), .QN(n1774) );
  DFFRX1 \I_cache/cache_reg[0][118]  ( .D(n9220), .CK(clk), .RN(n4336), .Q(
        \I_cache/cache[0][118] ), .QN(n866) );
  DFFRX1 \I_cache/cache_reg[1][118]  ( .D(n9219), .CK(clk), .RN(n4336), .Q(
        \I_cache/cache[1][118] ), .QN(n1799) );
  DFFRX1 \I_cache/cache_reg[2][118]  ( .D(n9218), .CK(clk), .RN(n4336), .Q(
        \I_cache/cache[2][118] ), .QN(n868) );
  DFFRX1 \I_cache/cache_reg[3][118]  ( .D(n9217), .CK(clk), .RN(n4336), .Q(
        \I_cache/cache[3][118] ), .QN(n1801) );
  DFFRX1 \I_cache/cache_reg[4][118]  ( .D(n9216), .CK(clk), .RN(n4336), .Q(
        \I_cache/cache[4][118] ), .QN(n867) );
  DFFRX1 \I_cache/cache_reg[5][118]  ( .D(n9215), .CK(clk), .RN(n4336), .Q(
        \I_cache/cache[5][118] ), .QN(n1800) );
  DFFRX1 \I_cache/cache_reg[6][118]  ( .D(n9214), .CK(clk), .RN(n4336), .Q(
        \I_cache/cache[6][118] ), .QN(n911) );
  DFFRX1 \I_cache/cache_reg[7][118]  ( .D(n9213), .CK(clk), .RN(n4336), .Q(
        \I_cache/cache[7][118] ), .QN(n1844) );
  DFFRX1 \I_cache/cache_reg[0][119]  ( .D(n9212), .CK(clk), .RN(n4336), .Q(
        \I_cache/cache[0][119] ), .QN(n774) );
  DFFRX1 \I_cache/cache_reg[1][119]  ( .D(n9211), .CK(clk), .RN(n4336), .Q(
        \I_cache/cache[1][119] ), .QN(n1707) );
  DFFRX1 \I_cache/cache_reg[2][119]  ( .D(n9210), .CK(clk), .RN(n4336), .Q(
        \I_cache/cache[2][119] ), .QN(n776) );
  DFFRX1 \I_cache/cache_reg[3][119]  ( .D(n9209), .CK(clk), .RN(n4336), .Q(
        \I_cache/cache[3][119] ), .QN(n1709) );
  DFFRX1 \I_cache/cache_reg[4][119]  ( .D(n9208), .CK(clk), .RN(n4337), .Q(
        \I_cache/cache[4][119] ), .QN(n775) );
  DFFRX1 \I_cache/cache_reg[5][119]  ( .D(n9207), .CK(clk), .RN(n4337), .Q(
        \I_cache/cache[5][119] ), .QN(n1708) );
  DFFRX1 \I_cache/cache_reg[6][119]  ( .D(n9206), .CK(clk), .RN(n4337), .Q(
        \I_cache/cache[6][119] ), .QN(n838) );
  DFFRX1 \I_cache/cache_reg[7][119]  ( .D(n9205), .CK(clk), .RN(n4337), .Q(
        \I_cache/cache[7][119] ), .QN(n1771) );
  DFFRX1 \I_cache/cache_reg[0][120]  ( .D(n9204), .CK(clk), .RN(n4337), .Q(
        \I_cache/cache[0][120] ), .QN(n853) );
  DFFRX1 \I_cache/cache_reg[1][120]  ( .D(n9203), .CK(clk), .RN(n4337), .Q(
        \I_cache/cache[1][120] ), .QN(n1786) );
  DFFRX1 \I_cache/cache_reg[2][120]  ( .D(n9202), .CK(clk), .RN(n4337), .Q(
        \I_cache/cache[2][120] ), .QN(n855) );
  DFFRX1 \I_cache/cache_reg[3][120]  ( .D(n9201), .CK(clk), .RN(n4337), .Q(
        \I_cache/cache[3][120] ), .QN(n1788) );
  DFFRX1 \I_cache/cache_reg[4][120]  ( .D(n9200), .CK(clk), .RN(n4337), .Q(
        \I_cache/cache[4][120] ), .QN(n854) );
  DFFRX1 \I_cache/cache_reg[5][120]  ( .D(n9199), .CK(clk), .RN(n4337), .Q(
        \I_cache/cache[5][120] ), .QN(n1787) );
  DFFRX1 \I_cache/cache_reg[6][120]  ( .D(n9198), .CK(clk), .RN(n4337), .Q(
        \I_cache/cache[6][120] ), .QN(n894) );
  DFFRX1 \I_cache/cache_reg[7][120]  ( .D(n9197), .CK(clk), .RN(n4337), .Q(
        \I_cache/cache[7][120] ), .QN(n1827) );
  DFFRX1 \I_cache/cache_reg[0][121]  ( .D(n9196), .CK(clk), .RN(n4338), .Q(
        \I_cache/cache[0][121] ), .QN(n873) );
  DFFRX1 \I_cache/cache_reg[1][121]  ( .D(n9195), .CK(clk), .RN(n4338), .Q(
        \I_cache/cache[1][121] ), .QN(n1806) );
  DFFRX1 \I_cache/cache_reg[2][121]  ( .D(n9194), .CK(clk), .RN(n4338), .Q(
        \I_cache/cache[2][121] ), .QN(n875) );
  DFFRX1 \I_cache/cache_reg[3][121]  ( .D(n9193), .CK(clk), .RN(n4338), .Q(
        \I_cache/cache[3][121] ), .QN(n1808) );
  DFFRX1 \I_cache/cache_reg[4][121]  ( .D(n9192), .CK(clk), .RN(n4338), .Q(
        \I_cache/cache[4][121] ), .QN(n874) );
  DFFRX1 \I_cache/cache_reg[5][121]  ( .D(n9191), .CK(clk), .RN(n4338), .Q(
        \I_cache/cache[5][121] ), .QN(n1807) );
  DFFRX1 \I_cache/cache_reg[6][121]  ( .D(n9190), .CK(clk), .RN(n4338), .Q(
        \I_cache/cache[6][121] ), .QN(n901) );
  DFFRX1 \I_cache/cache_reg[7][121]  ( .D(n9189), .CK(clk), .RN(n4338), .Q(
        \I_cache/cache[7][121] ), .QN(n1834) );
  DFFRX1 \I_cache/cache_reg[0][122]  ( .D(n9188), .CK(clk), .RN(n4338), .Q(
        \I_cache/cache[0][122] ), .QN(n704) );
  DFFRX1 \I_cache/cache_reg[1][122]  ( .D(n9187), .CK(clk), .RN(n4338), .Q(
        \I_cache/cache[1][122] ), .QN(n1637) );
  DFFRX1 \I_cache/cache_reg[2][122]  ( .D(n9186), .CK(clk), .RN(n4338), .Q(
        \I_cache/cache[2][122] ), .QN(n706) );
  DFFRX1 \I_cache/cache_reg[3][122]  ( .D(n9185), .CK(clk), .RN(n4338), .Q(
        \I_cache/cache[3][122] ), .QN(n1639) );
  DFFRX1 \I_cache/cache_reg[4][122]  ( .D(n9184), .CK(clk), .RN(n4339), .Q(
        \I_cache/cache[4][122] ), .QN(n705) );
  DFFRX1 \I_cache/cache_reg[5][122]  ( .D(n9183), .CK(clk), .RN(n4339), .Q(
        \I_cache/cache[5][122] ), .QN(n1638) );
  DFFRX1 \I_cache/cache_reg[6][122]  ( .D(n9182), .CK(clk), .RN(n4339), .Q(
        \I_cache/cache[6][122] ), .QN(n814) );
  DFFRX1 \I_cache/cache_reg[7][122]  ( .D(n9181), .CK(clk), .RN(n4339), .Q(
        \I_cache/cache[7][122] ), .QN(n1747) );
  DFFRX1 \I_cache/cache_reg[0][123]  ( .D(n9180), .CK(clk), .RN(n4339), .Q(
        \I_cache/cache[0][123] ), .QN(n761) );
  DFFRX1 \I_cache/cache_reg[1][123]  ( .D(n9179), .CK(clk), .RN(n4339), .Q(
        \I_cache/cache[1][123] ), .QN(n1694) );
  DFFRX1 \I_cache/cache_reg[2][123]  ( .D(n9178), .CK(clk), .RN(n4339), .Q(
        \I_cache/cache[2][123] ), .QN(n763) );
  DFFRX1 \I_cache/cache_reg[3][123]  ( .D(n9177), .CK(clk), .RN(n4339), .Q(
        \I_cache/cache[3][123] ), .QN(n1696) );
  DFFRX1 \I_cache/cache_reg[4][123]  ( .D(n9176), .CK(clk), .RN(n4339), .Q(
        \I_cache/cache[4][123] ), .QN(n762) );
  DFFRX1 \I_cache/cache_reg[5][123]  ( .D(n9175), .CK(clk), .RN(n4339), .Q(
        \I_cache/cache[5][123] ), .QN(n1695) );
  DFFRX1 \I_cache/cache_reg[6][123]  ( .D(n9174), .CK(clk), .RN(n4339), .Q(
        \I_cache/cache[6][123] ), .QN(n833) );
  DFFRX1 \I_cache/cache_reg[7][123]  ( .D(n9173), .CK(clk), .RN(n4339), .Q(
        \I_cache/cache[7][123] ), .QN(n1766) );
  DFFRX1 \I_cache/cache_reg[0][124]  ( .D(n9172), .CK(clk), .RN(n4340), .Q(
        \I_cache/cache[0][124] ), .QN(n749) );
  DFFRX1 \I_cache/cache_reg[1][124]  ( .D(n9171), .CK(clk), .RN(n4340), .Q(
        \I_cache/cache[1][124] ), .QN(n1682) );
  DFFRX1 \I_cache/cache_reg[2][124]  ( .D(n9170), .CK(clk), .RN(n4340), .Q(
        \I_cache/cache[2][124] ), .QN(n751) );
  DFFRX1 \I_cache/cache_reg[3][124]  ( .D(n9169), .CK(clk), .RN(n4340), .Q(
        \I_cache/cache[3][124] ), .QN(n1684) );
  DFFRX1 \I_cache/cache_reg[4][124]  ( .D(n9168), .CK(clk), .RN(n4340), .Q(
        \I_cache/cache[4][124] ), .QN(n750) );
  DFFRX1 \I_cache/cache_reg[5][124]  ( .D(n9167), .CK(clk), .RN(n4340), .Q(
        \I_cache/cache[5][124] ), .QN(n1683) );
  DFFRX1 \I_cache/cache_reg[6][124]  ( .D(n9166), .CK(clk), .RN(n4340), .Q(
        \I_cache/cache[6][124] ), .QN(n829) );
  DFFRX1 \I_cache/cache_reg[7][124]  ( .D(n9165), .CK(clk), .RN(n4340), .Q(
        \I_cache/cache[7][124] ), .QN(n1762) );
  DFFRX1 \I_cache/cache_reg[0][125]  ( .D(n9164), .CK(clk), .RN(n4340), .Q(
        \I_cache/cache[0][125] ), .QN(n710) );
  DFFRX1 \I_cache/cache_reg[1][125]  ( .D(n9163), .CK(clk), .RN(n4340), .Q(
        \I_cache/cache[1][125] ), .QN(n1643) );
  DFFRX1 \I_cache/cache_reg[2][125]  ( .D(n9162), .CK(clk), .RN(n4340), .Q(
        \I_cache/cache[2][125] ), .QN(n712) );
  DFFRX1 \I_cache/cache_reg[3][125]  ( .D(n9161), .CK(clk), .RN(n4340), .Q(
        \I_cache/cache[3][125] ), .QN(n1645) );
  DFFRX1 \I_cache/cache_reg[4][125]  ( .D(n9160), .CK(clk), .RN(n4341), .Q(
        \I_cache/cache[4][125] ), .QN(n711) );
  DFFRX1 \I_cache/cache_reg[5][125]  ( .D(n9159), .CK(clk), .RN(n4341), .Q(
        \I_cache/cache[5][125] ), .QN(n1644) );
  DFFRX1 \I_cache/cache_reg[6][125]  ( .D(n9158), .CK(clk), .RN(n4341), .Q(
        \I_cache/cache[6][125] ), .QN(n816) );
  DFFRX1 \I_cache/cache_reg[7][125]  ( .D(n9157), .CK(clk), .RN(n4341), .Q(
        \I_cache/cache[7][125] ), .QN(n1749) );
  DFFRX1 \I_cache/cache_reg[0][126]  ( .D(n9156), .CK(clk), .RN(n4341), .Q(
        \I_cache/cache[0][126] ), .QN(n731) );
  DFFRX1 \I_cache/cache_reg[1][126]  ( .D(n9155), .CK(clk), .RN(n4341), .Q(
        \I_cache/cache[1][126] ), .QN(n1664) );
  DFFRX1 \I_cache/cache_reg[2][126]  ( .D(n9154), .CK(clk), .RN(n4341), .Q(
        \I_cache/cache[2][126] ), .QN(n733) );
  DFFRX1 \I_cache/cache_reg[3][126]  ( .D(n9153), .CK(clk), .RN(n4341), .Q(
        \I_cache/cache[3][126] ), .QN(n1666) );
  DFFRX1 \I_cache/cache_reg[4][126]  ( .D(n9152), .CK(clk), .RN(n4341), .Q(
        \I_cache/cache[4][126] ), .QN(n732) );
  DFFRX1 \I_cache/cache_reg[5][126]  ( .D(n9151), .CK(clk), .RN(n4341), .Q(
        \I_cache/cache[5][126] ), .QN(n1665) );
  DFFRX1 \I_cache/cache_reg[6][126]  ( .D(n9150), .CK(clk), .RN(n4341), .Q(
        \I_cache/cache[6][126] ), .QN(n823) );
  DFFRX1 \I_cache/cache_reg[7][126]  ( .D(n9149), .CK(clk), .RN(n4341), .Q(
        \I_cache/cache[7][126] ), .QN(n1756) );
  DFFRX1 \I_cache/cache_reg[0][127]  ( .D(n9148), .CK(clk), .RN(n4342), .Q(
        \I_cache/cache[0][127] ), .QN(n722) );
  DFFRX1 \I_cache/cache_reg[1][127]  ( .D(n9147), .CK(clk), .RN(n4342), .Q(
        \I_cache/cache[1][127] ), .QN(n1655) );
  DFFRX1 \I_cache/cache_reg[2][127]  ( .D(n9146), .CK(clk), .RN(n4342), .Q(
        \I_cache/cache[2][127] ), .QN(n724) );
  DFFRX1 \I_cache/cache_reg[3][127]  ( .D(n9145), .CK(clk), .RN(n4342), .Q(
        \I_cache/cache[3][127] ), .QN(n1657) );
  DFFRX1 \I_cache/cache_reg[4][127]  ( .D(n9144), .CK(clk), .RN(n4342), .Q(
        \I_cache/cache[4][127] ), .QN(n723) );
  DFFRX1 \I_cache/cache_reg[5][127]  ( .D(n9143), .CK(clk), .RN(n4342), .Q(
        \I_cache/cache[5][127] ), .QN(n1656) );
  DFFRX1 \I_cache/cache_reg[6][127]  ( .D(n9142), .CK(clk), .RN(n4342), .Q(
        \I_cache/cache[6][127] ), .QN(n820) );
  DFFRX1 \I_cache/cache_reg[7][127]  ( .D(n9141), .CK(clk), .RN(n4342), .Q(
        \I_cache/cache[7][127] ), .QN(n1753) );
  DFFRX1 \i_MIPS/IF_ID_reg[58]  ( .D(\i_MIPS/N81 ), .CK(clk), .RN(n4061), .Q(
        \i_MIPS/IR_ID[26] ), .QN(\i_MIPS/n322 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[6]  ( .D(\i_MIPS/n468 ), .CK(clk), .RN(n4055), .Q(
        \i_MIPS/EX_MEM[6] ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[5]  ( .D(\i_MIPS/n469 ), .CK(clk), .RN(n4055), .Q(
        \i_MIPS/EX_MEM[5] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][0]  ( .D(\i_MIPS/Register/n148 ), 
        .CK(clk), .RN(n4071), .Q(\i_MIPS/Register/register[30][0] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][1]  ( .D(\i_MIPS/Register/n149 ), 
        .CK(clk), .RN(n4071), .Q(\i_MIPS/Register/register[30][1] ) );
  DFFRX1 \i_MIPS/Register/register_reg[28][0]  ( .D(\i_MIPS/Register/n212 ), 
        .CK(clk), .RN(n4076), .Q(\i_MIPS/Register/register[28][0] ) );
  DFFRX1 \i_MIPS/Register/register_reg[28][1]  ( .D(\i_MIPS/Register/n213 ), 
        .CK(clk), .RN(n4076), .Q(\i_MIPS/Register/register[28][1] ) );
  DFFRX1 \i_MIPS/Register/register_reg[24][0]  ( .D(\i_MIPS/Register/n340 ), 
        .CK(clk), .RN(n4087), .Q(\i_MIPS/Register/register[24][0] ) );
  DFFRX1 \i_MIPS/Register/register_reg[24][1]  ( .D(\i_MIPS/Register/n341 ), 
        .CK(clk), .RN(n4087), .Q(\i_MIPS/Register/register[24][1] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][0]  ( .D(\i_MIPS/Register/n660 ), 
        .CK(clk), .RN(n4114), .Q(\i_MIPS/Register/register[14][0] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][1]  ( .D(\i_MIPS/Register/n661 ), 
        .CK(clk), .RN(n4114), .Q(\i_MIPS/Register/register[14][1] ) );
  DFFRX1 \i_MIPS/Register/register_reg[12][0]  ( .D(\i_MIPS/Register/n724 ), 
        .CK(clk), .RN(n4119), .Q(\i_MIPS/Register/register[12][0] ) );
  DFFRX1 \i_MIPS/Register/register_reg[12][1]  ( .D(\i_MIPS/Register/n725 ), 
        .CK(clk), .RN(n4119), .Q(\i_MIPS/Register/register[12][1] ) );
  DFFRX1 \i_MIPS/Register/register_reg[8][0]  ( .D(\i_MIPS/Register/n852 ), 
        .CK(clk), .RN(n4130), .Q(\i_MIPS/Register/register[8][0] ) );
  DFFRX1 \i_MIPS/Register/register_reg[8][1]  ( .D(\i_MIPS/Register/n853 ), 
        .CK(clk), .RN(n4130), .Q(\i_MIPS/Register/register[8][1] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][0]  ( .D(\i_MIPS/Register/n404 ), 
        .CK(clk), .RN(n4092), .Q(\i_MIPS/Register/register[22][0] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][1]  ( .D(\i_MIPS/Register/n405 ), 
        .CK(clk), .RN(n4092), .Q(\i_MIPS/Register/register[22][1] ) );
  DFFRX1 \i_MIPS/Register/register_reg[20][0]  ( .D(\i_MIPS/Register/n468 ), 
        .CK(clk), .RN(n4098), .Q(\i_MIPS/Register/register[20][0] ) );
  DFFRX1 \i_MIPS/Register/register_reg[20][1]  ( .D(\i_MIPS/Register/n469 ), 
        .CK(clk), .RN(n4098), .Q(\i_MIPS/Register/register[20][1] ) );
  DFFRX1 \i_MIPS/Register/register_reg[16][0]  ( .D(\i_MIPS/Register/n596 ), 
        .CK(clk), .RN(n4108), .Q(\i_MIPS/Register/register[16][0] ) );
  DFFRX1 \i_MIPS/Register/register_reg[16][1]  ( .D(\i_MIPS/Register/n597 ), 
        .CK(clk), .RN(n4108), .Q(\i_MIPS/Register/register[16][1] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][0]  ( .D(\i_MIPS/Register/n916 ), 
        .CK(clk), .RN(n4135), .Q(\i_MIPS/Register/register[6][0] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][1]  ( .D(\i_MIPS/Register/n917 ), 
        .CK(clk), .RN(n4135), .Q(\i_MIPS/Register/register[6][1] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][5]  ( .D(\i_MIPS/Register/n921 ), 
        .CK(clk), .RN(n4135), .Q(\i_MIPS/Register/register[6][5] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][12]  ( .D(\i_MIPS/Register/n928 ), 
        .CK(clk), .RN(n4136), .Q(\i_MIPS/Register/register[6][12] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][24]  ( .D(\i_MIPS/Register/n940 ), 
        .CK(clk), .RN(n4137), .Q(\i_MIPS/Register/register[6][24] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][26]  ( .D(\i_MIPS/Register/n942 ), 
        .CK(clk), .RN(n4137), .Q(\i_MIPS/Register/register[6][26] ) );
  DFFRX1 \i_MIPS/Register/register_reg[4][0]  ( .D(\i_MIPS/Register/n980 ), 
        .CK(clk), .RN(n4140), .Q(\i_MIPS/Register/register[4][0] ) );
  DFFRX1 \i_MIPS/Register/register_reg[4][1]  ( .D(\i_MIPS/Register/n981 ), 
        .CK(clk), .RN(n4140), .Q(\i_MIPS/Register/register[4][1] ) );
  DFFRX1 \i_MIPS/Register/register_reg[4][5]  ( .D(\i_MIPS/Register/n985 ), 
        .CK(clk), .RN(n4141), .Q(\i_MIPS/Register/register[4][5] ) );
  DFFRX1 \i_MIPS/Register/register_reg[4][12]  ( .D(\i_MIPS/Register/n992 ), 
        .CK(clk), .RN(n4141), .Q(\i_MIPS/Register/register[4][12] ) );
  DFFRX1 \i_MIPS/Register/register_reg[4][24]  ( .D(\i_MIPS/Register/n1004 ), 
        .CK(clk), .RN(n4142), .Q(\i_MIPS/Register/register[4][24] ) );
  DFFRX1 \i_MIPS/Register/register_reg[4][26]  ( .D(\i_MIPS/Register/n1006 ), 
        .CK(clk), .RN(n4142), .Q(\i_MIPS/Register/register[4][26] ) );
  DFFRX1 \i_MIPS/Register/register_reg[0][0]  ( .D(\i_MIPS/Register/n1108 ), 
        .CK(clk), .RN(n4151), .Q(\i_MIPS/Register/register[0][0] ) );
  DFFRX1 \i_MIPS/Register/register_reg[0][1]  ( .D(\i_MIPS/Register/n1109 ), 
        .CK(clk), .RN(n4151), .Q(\i_MIPS/Register/register[0][1] ) );
  DFFRX1 \i_MIPS/Register/register_reg[0][5]  ( .D(\i_MIPS/Register/n1113 ), 
        .CK(clk), .RN(n4151), .Q(\i_MIPS/Register/register[0][5] ) );
  DFFRX1 \i_MIPS/Register/register_reg[0][12]  ( .D(\i_MIPS/Register/n1120 ), 
        .CK(clk), .RN(n4152), .Q(\i_MIPS/Register/register[0][12] ) );
  DFFRX1 \i_MIPS/Register/register_reg[0][24]  ( .D(\i_MIPS/Register/n1132 ), 
        .CK(clk), .RN(n4153), .Q(\i_MIPS/Register/register[0][24] ) );
  DFFRX1 \i_MIPS/Register/register_reg[0][26]  ( .D(\i_MIPS/Register/n1134 ), 
        .CK(clk), .RN(n4153), .Q(\i_MIPS/Register/register[0][26] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][2]  ( .D(\i_MIPS/Register/n150 ), 
        .CK(clk), .RN(n4071), .Q(\i_MIPS/Register/register[30][2] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][3]  ( .D(\i_MIPS/Register/n151 ), 
        .CK(clk), .RN(n4071), .Q(\i_MIPS/Register/register[30][3] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][4]  ( .D(\i_MIPS/Register/n152 ), 
        .CK(clk), .RN(n4071), .Q(\i_MIPS/Register/register[30][4] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][5]  ( .D(\i_MIPS/Register/n153 ), 
        .CK(clk), .RN(n4071), .Q(\i_MIPS/Register/register[30][5] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][6]  ( .D(\i_MIPS/Register/n154 ), 
        .CK(clk), .RN(n4071), .Q(\i_MIPS/Register/register[30][6] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][7]  ( .D(\i_MIPS/Register/n155 ), 
        .CK(clk), .RN(n4071), .Q(\i_MIPS/Register/register[30][7] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][8]  ( .D(\i_MIPS/Register/n156 ), 
        .CK(clk), .RN(n4072), .Q(\i_MIPS/Register/register[30][8] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][9]  ( .D(\i_MIPS/Register/n157 ), 
        .CK(clk), .RN(n4072), .Q(\i_MIPS/Register/register[30][9] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][10]  ( .D(\i_MIPS/Register/n158 ), 
        .CK(clk), .RN(n4072), .Q(\i_MIPS/Register/register[30][10] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][11]  ( .D(\i_MIPS/Register/n159 ), 
        .CK(clk), .RN(n4072), .Q(\i_MIPS/Register/register[30][11] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][12]  ( .D(\i_MIPS/Register/n160 ), 
        .CK(clk), .RN(n4072), .Q(\i_MIPS/Register/register[30][12] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][13]  ( .D(\i_MIPS/Register/n161 ), 
        .CK(clk), .RN(n4072), .Q(\i_MIPS/Register/register[30][13] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][14]  ( .D(\i_MIPS/Register/n162 ), 
        .CK(clk), .RN(n4072), .Q(\i_MIPS/Register/register[30][14] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][15]  ( .D(\i_MIPS/Register/n163 ), 
        .CK(clk), .RN(n4072), .Q(\i_MIPS/Register/register[30][15] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][16]  ( .D(\i_MIPS/Register/n164 ), 
        .CK(clk), .RN(n4072), .Q(\i_MIPS/Register/register[30][16] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][17]  ( .D(\i_MIPS/Register/n165 ), 
        .CK(clk), .RN(n4072), .Q(\i_MIPS/Register/register[30][17] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][18]  ( .D(\i_MIPS/Register/n166 ), 
        .CK(clk), .RN(n4072), .Q(\i_MIPS/Register/register[30][18] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][19]  ( .D(\i_MIPS/Register/n167 ), 
        .CK(clk), .RN(n4072), .Q(\i_MIPS/Register/register[30][19] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][20]  ( .D(\i_MIPS/Register/n168 ), 
        .CK(clk), .RN(n4073), .Q(\i_MIPS/Register/register[30][20] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][21]  ( .D(\i_MIPS/Register/n169 ), 
        .CK(clk), .RN(n4073), .Q(\i_MIPS/Register/register[30][21] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][22]  ( .D(\i_MIPS/Register/n170 ), 
        .CK(clk), .RN(n4073), .Q(\i_MIPS/Register/register[30][22] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][23]  ( .D(\i_MIPS/Register/n171 ), 
        .CK(clk), .RN(n4073), .Q(\i_MIPS/Register/register[30][23] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][24]  ( .D(\i_MIPS/Register/n172 ), 
        .CK(clk), .RN(n4073), .Q(\i_MIPS/Register/register[30][24] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][25]  ( .D(\i_MIPS/Register/n173 ), 
        .CK(clk), .RN(n4073), .Q(\i_MIPS/Register/register[30][25] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][26]  ( .D(\i_MIPS/Register/n174 ), 
        .CK(clk), .RN(n4073), .Q(\i_MIPS/Register/register[30][26] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][27]  ( .D(\i_MIPS/Register/n175 ), 
        .CK(clk), .RN(n4073), .Q(\i_MIPS/Register/register[30][27] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][28]  ( .D(\i_MIPS/Register/n176 ), 
        .CK(clk), .RN(n4073), .Q(\i_MIPS/Register/register[30][28] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][29]  ( .D(\i_MIPS/Register/n177 ), 
        .CK(clk), .RN(n4073), .Q(\i_MIPS/Register/register[30][29] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][30]  ( .D(\i_MIPS/Register/n178 ), 
        .CK(clk), .RN(n4073), .Q(\i_MIPS/Register/register[30][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][31]  ( .D(\i_MIPS/Register/n179 ), 
        .CK(clk), .RN(n4073), .Q(\i_MIPS/Register/register[30][31] ) );
  DFFRX1 \i_MIPS/Register/register_reg[28][2]  ( .D(\i_MIPS/Register/n214 ), 
        .CK(clk), .RN(n4076), .Q(\i_MIPS/Register/register[28][2] ) );
  DFFRX1 \i_MIPS/Register/register_reg[28][3]  ( .D(\i_MIPS/Register/n215 ), 
        .CK(clk), .RN(n4076), .Q(\i_MIPS/Register/register[28][3] ) );
  DFFRX1 \i_MIPS/Register/register_reg[28][4]  ( .D(\i_MIPS/Register/n216 ), 
        .CK(clk), .RN(n4077), .Q(\i_MIPS/Register/register[28][4] ) );
  DFFRX1 \i_MIPS/Register/register_reg[28][5]  ( .D(\i_MIPS/Register/n217 ), 
        .CK(clk), .RN(n4077), .Q(\i_MIPS/Register/register[28][5] ) );
  DFFRX1 \i_MIPS/Register/register_reg[28][6]  ( .D(\i_MIPS/Register/n218 ), 
        .CK(clk), .RN(n4077), .Q(\i_MIPS/Register/register[28][6] ) );
  DFFRX1 \i_MIPS/Register/register_reg[28][7]  ( .D(\i_MIPS/Register/n219 ), 
        .CK(clk), .RN(n4077), .Q(\i_MIPS/Register/register[28][7] ) );
  DFFRX1 \i_MIPS/Register/register_reg[28][8]  ( .D(\i_MIPS/Register/n220 ), 
        .CK(clk), .RN(n4077), .Q(\i_MIPS/Register/register[28][8] ) );
  DFFRX1 \i_MIPS/Register/register_reg[28][9]  ( .D(\i_MIPS/Register/n221 ), 
        .CK(clk), .RN(n4077), .Q(\i_MIPS/Register/register[28][9] ) );
  DFFRX1 \i_MIPS/Register/register_reg[28][10]  ( .D(\i_MIPS/Register/n222 ), 
        .CK(clk), .RN(n4077), .Q(\i_MIPS/Register/register[28][10] ) );
  DFFRX1 \i_MIPS/Register/register_reg[28][11]  ( .D(\i_MIPS/Register/n223 ), 
        .CK(clk), .RN(n4077), .Q(\i_MIPS/Register/register[28][11] ) );
  DFFRX1 \i_MIPS/Register/register_reg[28][12]  ( .D(\i_MIPS/Register/n224 ), 
        .CK(clk), .RN(n4077), .Q(\i_MIPS/Register/register[28][12] ) );
  DFFRX1 \i_MIPS/Register/register_reg[28][13]  ( .D(\i_MIPS/Register/n225 ), 
        .CK(clk), .RN(n4077), .Q(\i_MIPS/Register/register[28][13] ) );
  DFFRX1 \i_MIPS/Register/register_reg[28][14]  ( .D(\i_MIPS/Register/n226 ), 
        .CK(clk), .RN(n4077), .Q(\i_MIPS/Register/register[28][14] ) );
  DFFRX1 \i_MIPS/Register/register_reg[28][15]  ( .D(\i_MIPS/Register/n227 ), 
        .CK(clk), .RN(n4077), .Q(\i_MIPS/Register/register[28][15] ) );
  DFFRX1 \i_MIPS/Register/register_reg[28][16]  ( .D(\i_MIPS/Register/n228 ), 
        .CK(clk), .RN(n4078), .Q(\i_MIPS/Register/register[28][16] ) );
  DFFRX1 \i_MIPS/Register/register_reg[28][17]  ( .D(\i_MIPS/Register/n229 ), 
        .CK(clk), .RN(n4078), .Q(\i_MIPS/Register/register[28][17] ) );
  DFFRX1 \i_MIPS/Register/register_reg[28][18]  ( .D(\i_MIPS/Register/n230 ), 
        .CK(clk), .RN(n4078), .Q(\i_MIPS/Register/register[28][18] ) );
  DFFRX1 \i_MIPS/Register/register_reg[28][19]  ( .D(\i_MIPS/Register/n231 ), 
        .CK(clk), .RN(n4078), .Q(\i_MIPS/Register/register[28][19] ) );
  DFFRX1 \i_MIPS/Register/register_reg[28][20]  ( .D(\i_MIPS/Register/n232 ), 
        .CK(clk), .RN(n4078), .Q(\i_MIPS/Register/register[28][20] ) );
  DFFRX1 \i_MIPS/Register/register_reg[28][21]  ( .D(\i_MIPS/Register/n233 ), 
        .CK(clk), .RN(n4078), .Q(\i_MIPS/Register/register[28][21] ) );
  DFFRX1 \i_MIPS/Register/register_reg[28][22]  ( .D(\i_MIPS/Register/n234 ), 
        .CK(clk), .RN(n4078), .Q(\i_MIPS/Register/register[28][22] ) );
  DFFRX1 \i_MIPS/Register/register_reg[28][23]  ( .D(\i_MIPS/Register/n235 ), 
        .CK(clk), .RN(n4078), .Q(\i_MIPS/Register/register[28][23] ) );
  DFFRX1 \i_MIPS/Register/register_reg[28][24]  ( .D(\i_MIPS/Register/n236 ), 
        .CK(clk), .RN(n4078), .Q(\i_MIPS/Register/register[28][24] ) );
  DFFRX1 \i_MIPS/Register/register_reg[28][25]  ( .D(\i_MIPS/Register/n237 ), 
        .CK(clk), .RN(n4078), .Q(\i_MIPS/Register/register[28][25] ) );
  DFFRX1 \i_MIPS/Register/register_reg[28][26]  ( .D(\i_MIPS/Register/n238 ), 
        .CK(clk), .RN(n4078), .Q(\i_MIPS/Register/register[28][26] ) );
  DFFRX1 \i_MIPS/Register/register_reg[28][27]  ( .D(\i_MIPS/Register/n239 ), 
        .CK(clk), .RN(n4078), .Q(\i_MIPS/Register/register[28][27] ) );
  DFFRX1 \i_MIPS/Register/register_reg[28][28]  ( .D(\i_MIPS/Register/n240 ), 
        .CK(clk), .RN(n4079), .Q(\i_MIPS/Register/register[28][28] ) );
  DFFRX1 \i_MIPS/Register/register_reg[28][29]  ( .D(\i_MIPS/Register/n241 ), 
        .CK(clk), .RN(n4079), .Q(\i_MIPS/Register/register[28][29] ) );
  DFFRX1 \i_MIPS/Register/register_reg[28][30]  ( .D(\i_MIPS/Register/n242 ), 
        .CK(clk), .RN(n4079), .Q(\i_MIPS/Register/register[28][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[28][31]  ( .D(\i_MIPS/Register/n243 ), 
        .CK(clk), .RN(n4079), .Q(\i_MIPS/Register/register[28][31] ) );
  DFFRX1 \i_MIPS/Register/register_reg[24][2]  ( .D(\i_MIPS/Register/n342 ), 
        .CK(clk), .RN(n4087), .Q(\i_MIPS/Register/register[24][2] ) );
  DFFRX1 \i_MIPS/Register/register_reg[24][3]  ( .D(\i_MIPS/Register/n343 ), 
        .CK(clk), .RN(n4087), .Q(\i_MIPS/Register/register[24][3] ) );
  DFFRX1 \i_MIPS/Register/register_reg[24][4]  ( .D(\i_MIPS/Register/n344 ), 
        .CK(clk), .RN(n4087), .Q(\i_MIPS/Register/register[24][4] ) );
  DFFRX1 \i_MIPS/Register/register_reg[24][5]  ( .D(\i_MIPS/Register/n345 ), 
        .CK(clk), .RN(n4087), .Q(\i_MIPS/Register/register[24][5] ) );
  DFFRX1 \i_MIPS/Register/register_reg[24][6]  ( .D(\i_MIPS/Register/n346 ), 
        .CK(clk), .RN(n4087), .Q(\i_MIPS/Register/register[24][6] ) );
  DFFRX1 \i_MIPS/Register/register_reg[24][7]  ( .D(\i_MIPS/Register/n347 ), 
        .CK(clk), .RN(n4087), .Q(\i_MIPS/Register/register[24][7] ) );
  DFFRX1 \i_MIPS/Register/register_reg[24][8]  ( .D(\i_MIPS/Register/n348 ), 
        .CK(clk), .RN(n4088), .Q(\i_MIPS/Register/register[24][8] ) );
  DFFRX1 \i_MIPS/Register/register_reg[24][9]  ( .D(\i_MIPS/Register/n349 ), 
        .CK(clk), .RN(n4088), .Q(\i_MIPS/Register/register[24][9] ) );
  DFFRX1 \i_MIPS/Register/register_reg[24][10]  ( .D(\i_MIPS/Register/n350 ), 
        .CK(clk), .RN(n4088), .Q(\i_MIPS/Register/register[24][10] ) );
  DFFRX1 \i_MIPS/Register/register_reg[24][11]  ( .D(\i_MIPS/Register/n351 ), 
        .CK(clk), .RN(n4088), .Q(\i_MIPS/Register/register[24][11] ) );
  DFFRX1 \i_MIPS/Register/register_reg[24][12]  ( .D(\i_MIPS/Register/n352 ), 
        .CK(clk), .RN(n4088), .Q(\i_MIPS/Register/register[24][12] ) );
  DFFRX1 \i_MIPS/Register/register_reg[24][13]  ( .D(\i_MIPS/Register/n353 ), 
        .CK(clk), .RN(n4088), .Q(\i_MIPS/Register/register[24][13] ) );
  DFFRX1 \i_MIPS/Register/register_reg[24][14]  ( .D(\i_MIPS/Register/n354 ), 
        .CK(clk), .RN(n4088), .Q(\i_MIPS/Register/register[24][14] ) );
  DFFRX1 \i_MIPS/Register/register_reg[24][15]  ( .D(\i_MIPS/Register/n355 ), 
        .CK(clk), .RN(n4088), .Q(\i_MIPS/Register/register[24][15] ) );
  DFFRX1 \i_MIPS/Register/register_reg[24][16]  ( .D(\i_MIPS/Register/n356 ), 
        .CK(clk), .RN(n4088), .Q(\i_MIPS/Register/register[24][16] ) );
  DFFRX1 \i_MIPS/Register/register_reg[24][17]  ( .D(\i_MIPS/Register/n357 ), 
        .CK(clk), .RN(n4088), .Q(\i_MIPS/Register/register[24][17] ) );
  DFFRX1 \i_MIPS/Register/register_reg[24][18]  ( .D(\i_MIPS/Register/n358 ), 
        .CK(clk), .RN(n4088), .Q(\i_MIPS/Register/register[24][18] ) );
  DFFRX1 \i_MIPS/Register/register_reg[24][19]  ( .D(\i_MIPS/Register/n359 ), 
        .CK(clk), .RN(n4088), .Q(\i_MIPS/Register/register[24][19] ) );
  DFFRX1 \i_MIPS/Register/register_reg[24][20]  ( .D(\i_MIPS/Register/n360 ), 
        .CK(clk), .RN(n4089), .Q(\i_MIPS/Register/register[24][20] ) );
  DFFRX1 \i_MIPS/Register/register_reg[24][21]  ( .D(\i_MIPS/Register/n361 ), 
        .CK(clk), .RN(n4089), .Q(\i_MIPS/Register/register[24][21] ) );
  DFFRX1 \i_MIPS/Register/register_reg[24][22]  ( .D(\i_MIPS/Register/n362 ), 
        .CK(clk), .RN(n4089), .Q(\i_MIPS/Register/register[24][22] ) );
  DFFRX1 \i_MIPS/Register/register_reg[24][23]  ( .D(\i_MIPS/Register/n363 ), 
        .CK(clk), .RN(n4089), .Q(\i_MIPS/Register/register[24][23] ) );
  DFFRX1 \i_MIPS/Register/register_reg[24][24]  ( .D(\i_MIPS/Register/n364 ), 
        .CK(clk), .RN(n4089), .Q(\i_MIPS/Register/register[24][24] ) );
  DFFRX1 \i_MIPS/Register/register_reg[24][25]  ( .D(\i_MIPS/Register/n365 ), 
        .CK(clk), .RN(n4089), .Q(\i_MIPS/Register/register[24][25] ) );
  DFFRX1 \i_MIPS/Register/register_reg[24][26]  ( .D(\i_MIPS/Register/n366 ), 
        .CK(clk), .RN(n4089), .Q(\i_MIPS/Register/register[24][26] ) );
  DFFRX1 \i_MIPS/Register/register_reg[24][27]  ( .D(\i_MIPS/Register/n367 ), 
        .CK(clk), .RN(n4089), .Q(\i_MIPS/Register/register[24][27] ) );
  DFFRX1 \i_MIPS/Register/register_reg[24][28]  ( .D(\i_MIPS/Register/n368 ), 
        .CK(clk), .RN(n4089), .Q(\i_MIPS/Register/register[24][28] ) );
  DFFRX1 \i_MIPS/Register/register_reg[24][29]  ( .D(\i_MIPS/Register/n369 ), 
        .CK(clk), .RN(n4089), .Q(\i_MIPS/Register/register[24][29] ) );
  DFFRX1 \i_MIPS/Register/register_reg[24][30]  ( .D(\i_MIPS/Register/n370 ), 
        .CK(clk), .RN(n4089), .Q(\i_MIPS/Register/register[24][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[24][31]  ( .D(\i_MIPS/Register/n371 ), 
        .CK(clk), .RN(n4089), .Q(\i_MIPS/Register/register[24][31] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][2]  ( .D(\i_MIPS/Register/n662 ), 
        .CK(clk), .RN(n4114), .Q(\i_MIPS/Register/register[14][2] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][3]  ( .D(\i_MIPS/Register/n663 ), 
        .CK(clk), .RN(n4114), .Q(\i_MIPS/Register/register[14][3] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][4]  ( .D(\i_MIPS/Register/n664 ), 
        .CK(clk), .RN(n4114), .Q(\i_MIPS/Register/register[14][4] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][5]  ( .D(\i_MIPS/Register/n665 ), 
        .CK(clk), .RN(n4114), .Q(\i_MIPS/Register/register[14][5] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][6]  ( .D(\i_MIPS/Register/n666 ), 
        .CK(clk), .RN(n4114), .Q(\i_MIPS/Register/register[14][6] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][7]  ( .D(\i_MIPS/Register/n667 ), 
        .CK(clk), .RN(n4114), .Q(\i_MIPS/Register/register[14][7] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][8]  ( .D(\i_MIPS/Register/n668 ), 
        .CK(clk), .RN(n4114), .Q(\i_MIPS/Register/register[14][8] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][9]  ( .D(\i_MIPS/Register/n669 ), 
        .CK(clk), .RN(n4114), .Q(\i_MIPS/Register/register[14][9] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][10]  ( .D(\i_MIPS/Register/n670 ), 
        .CK(clk), .RN(n4114), .Q(\i_MIPS/Register/register[14][10] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][11]  ( .D(\i_MIPS/Register/n671 ), 
        .CK(clk), .RN(n4114), .Q(\i_MIPS/Register/register[14][11] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][12]  ( .D(\i_MIPS/Register/n672 ), 
        .CK(clk), .RN(n4115), .Q(\i_MIPS/Register/register[14][12] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][13]  ( .D(\i_MIPS/Register/n673 ), 
        .CK(clk), .RN(n4115), .Q(\i_MIPS/Register/register[14][13] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][14]  ( .D(\i_MIPS/Register/n674 ), 
        .CK(clk), .RN(n4115), .Q(\i_MIPS/Register/register[14][14] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][15]  ( .D(\i_MIPS/Register/n675 ), 
        .CK(clk), .RN(n4115), .Q(\i_MIPS/Register/register[14][15] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][16]  ( .D(\i_MIPS/Register/n676 ), 
        .CK(clk), .RN(n4115), .Q(\i_MIPS/Register/register[14][16] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][17]  ( .D(\i_MIPS/Register/n677 ), 
        .CK(clk), .RN(n4115), .Q(\i_MIPS/Register/register[14][17] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][18]  ( .D(\i_MIPS/Register/n678 ), 
        .CK(clk), .RN(n4115), .Q(\i_MIPS/Register/register[14][18] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][19]  ( .D(\i_MIPS/Register/n679 ), 
        .CK(clk), .RN(n4115), .Q(\i_MIPS/Register/register[14][19] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][20]  ( .D(\i_MIPS/Register/n680 ), 
        .CK(clk), .RN(n4115), .Q(\i_MIPS/Register/register[14][20] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][21]  ( .D(\i_MIPS/Register/n681 ), 
        .CK(clk), .RN(n4115), .Q(\i_MIPS/Register/register[14][21] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][22]  ( .D(\i_MIPS/Register/n682 ), 
        .CK(clk), .RN(n4115), .Q(\i_MIPS/Register/register[14][22] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][23]  ( .D(\i_MIPS/Register/n683 ), 
        .CK(clk), .RN(n4115), .Q(\i_MIPS/Register/register[14][23] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][24]  ( .D(\i_MIPS/Register/n684 ), 
        .CK(clk), .RN(n4116), .Q(\i_MIPS/Register/register[14][24] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][25]  ( .D(\i_MIPS/Register/n685 ), 
        .CK(clk), .RN(n4116), .Q(\i_MIPS/Register/register[14][25] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][26]  ( .D(\i_MIPS/Register/n686 ), 
        .CK(clk), .RN(n4116), .Q(\i_MIPS/Register/register[14][26] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][27]  ( .D(\i_MIPS/Register/n687 ), 
        .CK(clk), .RN(n4116), .Q(\i_MIPS/Register/register[14][27] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][28]  ( .D(\i_MIPS/Register/n688 ), 
        .CK(clk), .RN(n4116), .Q(\i_MIPS/Register/register[14][28] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][29]  ( .D(\i_MIPS/Register/n689 ), 
        .CK(clk), .RN(n4116), .Q(\i_MIPS/Register/register[14][29] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][30]  ( .D(\i_MIPS/Register/n690 ), 
        .CK(clk), .RN(n4116), .Q(\i_MIPS/Register/register[14][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][31]  ( .D(\i_MIPS/Register/n691 ), 
        .CK(clk), .RN(n4116), .Q(\i_MIPS/Register/register[14][31] ) );
  DFFRX1 \i_MIPS/Register/register_reg[12][2]  ( .D(\i_MIPS/Register/n726 ), 
        .CK(clk), .RN(n4119), .Q(\i_MIPS/Register/register[12][2] ) );
  DFFRX1 \i_MIPS/Register/register_reg[12][3]  ( .D(\i_MIPS/Register/n727 ), 
        .CK(clk), .RN(n4119), .Q(\i_MIPS/Register/register[12][3] ) );
  DFFRX1 \i_MIPS/Register/register_reg[12][4]  ( .D(\i_MIPS/Register/n728 ), 
        .CK(clk), .RN(n4119), .Q(\i_MIPS/Register/register[12][4] ) );
  DFFRX1 \i_MIPS/Register/register_reg[12][5]  ( .D(\i_MIPS/Register/n729 ), 
        .CK(clk), .RN(n4119), .Q(\i_MIPS/Register/register[12][5] ) );
  DFFRX1 \i_MIPS/Register/register_reg[12][6]  ( .D(\i_MIPS/Register/n730 ), 
        .CK(clk), .RN(n4119), .Q(\i_MIPS/Register/register[12][6] ) );
  DFFRX1 \i_MIPS/Register/register_reg[12][7]  ( .D(\i_MIPS/Register/n731 ), 
        .CK(clk), .RN(n4119), .Q(\i_MIPS/Register/register[12][7] ) );
  DFFRX1 \i_MIPS/Register/register_reg[12][8]  ( .D(\i_MIPS/Register/n732 ), 
        .CK(clk), .RN(n4120), .Q(\i_MIPS/Register/register[12][8] ) );
  DFFRX1 \i_MIPS/Register/register_reg[12][9]  ( .D(\i_MIPS/Register/n733 ), 
        .CK(clk), .RN(n4120), .Q(\i_MIPS/Register/register[12][9] ) );
  DFFRX1 \i_MIPS/Register/register_reg[12][10]  ( .D(\i_MIPS/Register/n734 ), 
        .CK(clk), .RN(n4120), .Q(\i_MIPS/Register/register[12][10] ) );
  DFFRX1 \i_MIPS/Register/register_reg[12][11]  ( .D(\i_MIPS/Register/n735 ), 
        .CK(clk), .RN(n4120), .Q(\i_MIPS/Register/register[12][11] ) );
  DFFRX1 \i_MIPS/Register/register_reg[12][12]  ( .D(\i_MIPS/Register/n736 ), 
        .CK(clk), .RN(n4120), .Q(\i_MIPS/Register/register[12][12] ) );
  DFFRX1 \i_MIPS/Register/register_reg[12][13]  ( .D(\i_MIPS/Register/n737 ), 
        .CK(clk), .RN(n4120), .Q(\i_MIPS/Register/register[12][13] ) );
  DFFRX1 \i_MIPS/Register/register_reg[12][14]  ( .D(\i_MIPS/Register/n738 ), 
        .CK(clk), .RN(n4120), .Q(\i_MIPS/Register/register[12][14] ) );
  DFFRX1 \i_MIPS/Register/register_reg[12][15]  ( .D(\i_MIPS/Register/n739 ), 
        .CK(clk), .RN(n4120), .Q(\i_MIPS/Register/register[12][15] ) );
  DFFRX1 \i_MIPS/Register/register_reg[12][16]  ( .D(\i_MIPS/Register/n740 ), 
        .CK(clk), .RN(n4120), .Q(\i_MIPS/Register/register[12][16] ) );
  DFFRX1 \i_MIPS/Register/register_reg[12][17]  ( .D(\i_MIPS/Register/n741 ), 
        .CK(clk), .RN(n4120), .Q(\i_MIPS/Register/register[12][17] ) );
  DFFRX1 \i_MIPS/Register/register_reg[12][18]  ( .D(\i_MIPS/Register/n742 ), 
        .CK(clk), .RN(n4120), .Q(\i_MIPS/Register/register[12][18] ) );
  DFFRX1 \i_MIPS/Register/register_reg[12][19]  ( .D(\i_MIPS/Register/n743 ), 
        .CK(clk), .RN(n4120), .Q(\i_MIPS/Register/register[12][19] ) );
  DFFRX1 \i_MIPS/Register/register_reg[12][20]  ( .D(\i_MIPS/Register/n744 ), 
        .CK(clk), .RN(n4121), .Q(\i_MIPS/Register/register[12][20] ) );
  DFFRX1 \i_MIPS/Register/register_reg[12][21]  ( .D(\i_MIPS/Register/n745 ), 
        .CK(clk), .RN(n4121), .Q(\i_MIPS/Register/register[12][21] ) );
  DFFRX1 \i_MIPS/Register/register_reg[12][22]  ( .D(\i_MIPS/Register/n746 ), 
        .CK(clk), .RN(n4121), .Q(\i_MIPS/Register/register[12][22] ) );
  DFFRX1 \i_MIPS/Register/register_reg[12][23]  ( .D(\i_MIPS/Register/n747 ), 
        .CK(clk), .RN(n4121), .Q(\i_MIPS/Register/register[12][23] ) );
  DFFRX1 \i_MIPS/Register/register_reg[12][24]  ( .D(\i_MIPS/Register/n748 ), 
        .CK(clk), .RN(n4121), .Q(\i_MIPS/Register/register[12][24] ) );
  DFFRX1 \i_MIPS/Register/register_reg[12][25]  ( .D(\i_MIPS/Register/n749 ), 
        .CK(clk), .RN(n4121), .Q(\i_MIPS/Register/register[12][25] ) );
  DFFRX1 \i_MIPS/Register/register_reg[12][26]  ( .D(\i_MIPS/Register/n750 ), 
        .CK(clk), .RN(n4121), .Q(\i_MIPS/Register/register[12][26] ) );
  DFFRX1 \i_MIPS/Register/register_reg[12][27]  ( .D(\i_MIPS/Register/n751 ), 
        .CK(clk), .RN(n4121), .Q(\i_MIPS/Register/register[12][27] ) );
  DFFRX1 \i_MIPS/Register/register_reg[12][28]  ( .D(\i_MIPS/Register/n752 ), 
        .CK(clk), .RN(n4121), .Q(\i_MIPS/Register/register[12][28] ) );
  DFFRX1 \i_MIPS/Register/register_reg[12][29]  ( .D(\i_MIPS/Register/n753 ), 
        .CK(clk), .RN(n4121), .Q(\i_MIPS/Register/register[12][29] ) );
  DFFRX1 \i_MIPS/Register/register_reg[12][30]  ( .D(\i_MIPS/Register/n754 ), 
        .CK(clk), .RN(n4121), .Q(\i_MIPS/Register/register[12][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[12][31]  ( .D(\i_MIPS/Register/n755 ), 
        .CK(clk), .RN(n4121), .Q(\i_MIPS/Register/register[12][31] ) );
  DFFRX1 \i_MIPS/Register/register_reg[8][2]  ( .D(\i_MIPS/Register/n854 ), 
        .CK(clk), .RN(n4130), .Q(\i_MIPS/Register/register[8][2] ) );
  DFFRX1 \i_MIPS/Register/register_reg[8][3]  ( .D(\i_MIPS/Register/n855 ), 
        .CK(clk), .RN(n4130), .Q(\i_MIPS/Register/register[8][3] ) );
  DFFRX1 \i_MIPS/Register/register_reg[8][4]  ( .D(\i_MIPS/Register/n856 ), 
        .CK(clk), .RN(n4130), .Q(\i_MIPS/Register/register[8][4] ) );
  DFFRX1 \i_MIPS/Register/register_reg[8][5]  ( .D(\i_MIPS/Register/n857 ), 
        .CK(clk), .RN(n4130), .Q(\i_MIPS/Register/register[8][5] ) );
  DFFRX1 \i_MIPS/Register/register_reg[8][6]  ( .D(\i_MIPS/Register/n858 ), 
        .CK(clk), .RN(n4130), .Q(\i_MIPS/Register/register[8][6] ) );
  DFFRX1 \i_MIPS/Register/register_reg[8][7]  ( .D(\i_MIPS/Register/n859 ), 
        .CK(clk), .RN(n4130), .Q(\i_MIPS/Register/register[8][7] ) );
  DFFRX1 \i_MIPS/Register/register_reg[8][8]  ( .D(\i_MIPS/Register/n860 ), 
        .CK(clk), .RN(n4130), .Q(\i_MIPS/Register/register[8][8] ) );
  DFFRX1 \i_MIPS/Register/register_reg[8][9]  ( .D(\i_MIPS/Register/n861 ), 
        .CK(clk), .RN(n4130), .Q(\i_MIPS/Register/register[8][9] ) );
  DFFRX1 \i_MIPS/Register/register_reg[8][10]  ( .D(\i_MIPS/Register/n862 ), 
        .CK(clk), .RN(n4130), .Q(\i_MIPS/Register/register[8][10] ) );
  DFFRX1 \i_MIPS/Register/register_reg[8][11]  ( .D(\i_MIPS/Register/n863 ), 
        .CK(clk), .RN(n4130), .Q(\i_MIPS/Register/register[8][11] ) );
  DFFRX1 \i_MIPS/Register/register_reg[8][12]  ( .D(\i_MIPS/Register/n864 ), 
        .CK(clk), .RN(n4131), .Q(\i_MIPS/Register/register[8][12] ) );
  DFFRX1 \i_MIPS/Register/register_reg[8][13]  ( .D(\i_MIPS/Register/n865 ), 
        .CK(clk), .RN(n4131), .Q(\i_MIPS/Register/register[8][13] ) );
  DFFRX1 \i_MIPS/Register/register_reg[8][14]  ( .D(\i_MIPS/Register/n866 ), 
        .CK(clk), .RN(n4131), .Q(\i_MIPS/Register/register[8][14] ) );
  DFFRX1 \i_MIPS/Register/register_reg[8][15]  ( .D(\i_MIPS/Register/n867 ), 
        .CK(clk), .RN(n4131), .Q(\i_MIPS/Register/register[8][15] ) );
  DFFRX1 \i_MIPS/Register/register_reg[8][16]  ( .D(\i_MIPS/Register/n868 ), 
        .CK(clk), .RN(n4131), .Q(\i_MIPS/Register/register[8][16] ) );
  DFFRX1 \i_MIPS/Register/register_reg[8][17]  ( .D(\i_MIPS/Register/n869 ), 
        .CK(clk), .RN(n4131), .Q(\i_MIPS/Register/register[8][17] ) );
  DFFRX1 \i_MIPS/Register/register_reg[8][18]  ( .D(\i_MIPS/Register/n870 ), 
        .CK(clk), .RN(n4131), .Q(\i_MIPS/Register/register[8][18] ) );
  DFFRX1 \i_MIPS/Register/register_reg[8][19]  ( .D(\i_MIPS/Register/n871 ), 
        .CK(clk), .RN(n4131), .Q(\i_MIPS/Register/register[8][19] ) );
  DFFRX1 \i_MIPS/Register/register_reg[8][20]  ( .D(\i_MIPS/Register/n872 ), 
        .CK(clk), .RN(n4131), .Q(\i_MIPS/Register/register[8][20] ) );
  DFFRX1 \i_MIPS/Register/register_reg[8][21]  ( .D(\i_MIPS/Register/n873 ), 
        .CK(clk), .RN(n4131), .Q(\i_MIPS/Register/register[8][21] ) );
  DFFRX1 \i_MIPS/Register/register_reg[8][22]  ( .D(\i_MIPS/Register/n874 ), 
        .CK(clk), .RN(n4131), .Q(\i_MIPS/Register/register[8][22] ) );
  DFFRX1 \i_MIPS/Register/register_reg[8][23]  ( .D(\i_MIPS/Register/n875 ), 
        .CK(clk), .RN(n4131), .Q(\i_MIPS/Register/register[8][23] ) );
  DFFRX1 \i_MIPS/Register/register_reg[8][24]  ( .D(\i_MIPS/Register/n876 ), 
        .CK(clk), .RN(n4132), .Q(\i_MIPS/Register/register[8][24] ) );
  DFFRX1 \i_MIPS/Register/register_reg[8][25]  ( .D(\i_MIPS/Register/n877 ), 
        .CK(clk), .RN(n4132), .Q(\i_MIPS/Register/register[8][25] ) );
  DFFRX1 \i_MIPS/Register/register_reg[8][26]  ( .D(\i_MIPS/Register/n878 ), 
        .CK(clk), .RN(n4132), .Q(\i_MIPS/Register/register[8][26] ) );
  DFFRX1 \i_MIPS/Register/register_reg[8][27]  ( .D(\i_MIPS/Register/n879 ), 
        .CK(clk), .RN(n4132), .Q(\i_MIPS/Register/register[8][27] ) );
  DFFRX1 \i_MIPS/Register/register_reg[8][28]  ( .D(\i_MIPS/Register/n880 ), 
        .CK(clk), .RN(n4132), .Q(\i_MIPS/Register/register[8][28] ) );
  DFFRX1 \i_MIPS/Register/register_reg[8][29]  ( .D(\i_MIPS/Register/n881 ), 
        .CK(clk), .RN(n4132), .Q(\i_MIPS/Register/register[8][29] ) );
  DFFRX1 \i_MIPS/Register/register_reg[8][30]  ( .D(\i_MIPS/Register/n882 ), 
        .CK(clk), .RN(n4132), .Q(\i_MIPS/Register/register[8][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[8][31]  ( .D(\i_MIPS/Register/n883 ), 
        .CK(clk), .RN(n4132), .Q(\i_MIPS/Register/register[8][31] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][2]  ( .D(\i_MIPS/Register/n406 ), 
        .CK(clk), .RN(n4092), .Q(\i_MIPS/Register/register[22][2] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][3]  ( .D(\i_MIPS/Register/n407 ), 
        .CK(clk), .RN(n4092), .Q(\i_MIPS/Register/register[22][3] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][4]  ( .D(\i_MIPS/Register/n408 ), 
        .CK(clk), .RN(n4093), .Q(\i_MIPS/Register/register[22][4] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][5]  ( .D(\i_MIPS/Register/n409 ), 
        .CK(clk), .RN(n4093), .Q(\i_MIPS/Register/register[22][5] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][6]  ( .D(\i_MIPS/Register/n410 ), 
        .CK(clk), .RN(n4093), .Q(\i_MIPS/Register/register[22][6] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][7]  ( .D(\i_MIPS/Register/n411 ), 
        .CK(clk), .RN(n4093), .Q(\i_MIPS/Register/register[22][7] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][8]  ( .D(\i_MIPS/Register/n412 ), 
        .CK(clk), .RN(n4093), .Q(\i_MIPS/Register/register[22][8] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][9]  ( .D(\i_MIPS/Register/n413 ), 
        .CK(clk), .RN(n4093), .Q(\i_MIPS/Register/register[22][9] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][10]  ( .D(\i_MIPS/Register/n414 ), 
        .CK(clk), .RN(n4093), .Q(\i_MIPS/Register/register[22][10] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][11]  ( .D(\i_MIPS/Register/n415 ), 
        .CK(clk), .RN(n4093), .Q(\i_MIPS/Register/register[22][11] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][12]  ( .D(\i_MIPS/Register/n416 ), 
        .CK(clk), .RN(n4093), .Q(\i_MIPS/Register/register[22][12] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][13]  ( .D(\i_MIPS/Register/n417 ), 
        .CK(clk), .RN(n4093), .Q(\i_MIPS/Register/register[22][13] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][14]  ( .D(\i_MIPS/Register/n418 ), 
        .CK(clk), .RN(n4093), .Q(\i_MIPS/Register/register[22][14] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][15]  ( .D(\i_MIPS/Register/n419 ), 
        .CK(clk), .RN(n4093), .Q(\i_MIPS/Register/register[22][15] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][16]  ( .D(\i_MIPS/Register/n420 ), 
        .CK(clk), .RN(n4094), .Q(\i_MIPS/Register/register[22][16] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][17]  ( .D(\i_MIPS/Register/n421 ), 
        .CK(clk), .RN(n4094), .Q(\i_MIPS/Register/register[22][17] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][18]  ( .D(\i_MIPS/Register/n422 ), 
        .CK(clk), .RN(n4094), .Q(\i_MIPS/Register/register[22][18] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][19]  ( .D(\i_MIPS/Register/n423 ), 
        .CK(clk), .RN(n4094), .Q(\i_MIPS/Register/register[22][19] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][20]  ( .D(\i_MIPS/Register/n424 ), 
        .CK(clk), .RN(n4094), .Q(\i_MIPS/Register/register[22][20] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][21]  ( .D(\i_MIPS/Register/n425 ), 
        .CK(clk), .RN(n4094), .Q(\i_MIPS/Register/register[22][21] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][22]  ( .D(\i_MIPS/Register/n426 ), 
        .CK(clk), .RN(n4094), .Q(\i_MIPS/Register/register[22][22] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][23]  ( .D(\i_MIPS/Register/n427 ), 
        .CK(clk), .RN(n4094), .Q(\i_MIPS/Register/register[22][23] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][24]  ( .D(\i_MIPS/Register/n428 ), 
        .CK(clk), .RN(n4094), .Q(\i_MIPS/Register/register[22][24] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][25]  ( .D(\i_MIPS/Register/n429 ), 
        .CK(clk), .RN(n4094), .Q(\i_MIPS/Register/register[22][25] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][26]  ( .D(\i_MIPS/Register/n430 ), 
        .CK(clk), .RN(n4094), .Q(\i_MIPS/Register/register[22][26] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][27]  ( .D(\i_MIPS/Register/n431 ), 
        .CK(clk), .RN(n4094), .Q(\i_MIPS/Register/register[22][27] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][28]  ( .D(\i_MIPS/Register/n432 ), 
        .CK(clk), .RN(n4095), .Q(\i_MIPS/Register/register[22][28] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][29]  ( .D(\i_MIPS/Register/n433 ), 
        .CK(clk), .RN(n4095), .Q(\i_MIPS/Register/register[22][29] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][30]  ( .D(\i_MIPS/Register/n434 ), 
        .CK(clk), .RN(n4095), .Q(\i_MIPS/Register/register[22][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][31]  ( .D(\i_MIPS/Register/n435 ), 
        .CK(clk), .RN(n4095), .Q(\i_MIPS/Register/register[22][31] ) );
  DFFRX1 \i_MIPS/Register/register_reg[20][2]  ( .D(\i_MIPS/Register/n470 ), 
        .CK(clk), .RN(n4098), .Q(\i_MIPS/Register/register[20][2] ) );
  DFFRX1 \i_MIPS/Register/register_reg[20][3]  ( .D(\i_MIPS/Register/n471 ), 
        .CK(clk), .RN(n4098), .Q(\i_MIPS/Register/register[20][3] ) );
  DFFRX1 \i_MIPS/Register/register_reg[20][4]  ( .D(\i_MIPS/Register/n472 ), 
        .CK(clk), .RN(n4098), .Q(\i_MIPS/Register/register[20][4] ) );
  DFFRX1 \i_MIPS/Register/register_reg[20][5]  ( .D(\i_MIPS/Register/n473 ), 
        .CK(clk), .RN(n4098), .Q(\i_MIPS/Register/register[20][5] ) );
  DFFRX1 \i_MIPS/Register/register_reg[20][6]  ( .D(\i_MIPS/Register/n474 ), 
        .CK(clk), .RN(n4098), .Q(\i_MIPS/Register/register[20][6] ) );
  DFFRX1 \i_MIPS/Register/register_reg[20][7]  ( .D(\i_MIPS/Register/n475 ), 
        .CK(clk), .RN(n4098), .Q(\i_MIPS/Register/register[20][7] ) );
  DFFRX1 \i_MIPS/Register/register_reg[20][8]  ( .D(\i_MIPS/Register/n476 ), 
        .CK(clk), .RN(n4098), .Q(\i_MIPS/Register/register[20][8] ) );
  DFFRX1 \i_MIPS/Register/register_reg[20][9]  ( .D(\i_MIPS/Register/n477 ), 
        .CK(clk), .RN(n4098), .Q(\i_MIPS/Register/register[20][9] ) );
  DFFRX1 \i_MIPS/Register/register_reg[20][10]  ( .D(\i_MIPS/Register/n478 ), 
        .CK(clk), .RN(n4098), .Q(\i_MIPS/Register/register[20][10] ) );
  DFFRX1 \i_MIPS/Register/register_reg[20][11]  ( .D(\i_MIPS/Register/n479 ), 
        .CK(clk), .RN(n4098), .Q(\i_MIPS/Register/register[20][11] ) );
  DFFRX1 \i_MIPS/Register/register_reg[20][12]  ( .D(\i_MIPS/Register/n480 ), 
        .CK(clk), .RN(n4099), .Q(\i_MIPS/Register/register[20][12] ) );
  DFFRX1 \i_MIPS/Register/register_reg[20][13]  ( .D(\i_MIPS/Register/n481 ), 
        .CK(clk), .RN(n4099), .Q(\i_MIPS/Register/register[20][13] ) );
  DFFRX1 \i_MIPS/Register/register_reg[20][14]  ( .D(\i_MIPS/Register/n482 ), 
        .CK(clk), .RN(n4099), .Q(\i_MIPS/Register/register[20][14] ) );
  DFFRX1 \i_MIPS/Register/register_reg[20][15]  ( .D(\i_MIPS/Register/n483 ), 
        .CK(clk), .RN(n4099), .Q(\i_MIPS/Register/register[20][15] ) );
  DFFRX1 \i_MIPS/Register/register_reg[20][16]  ( .D(\i_MIPS/Register/n484 ), 
        .CK(clk), .RN(n4099), .Q(\i_MIPS/Register/register[20][16] ) );
  DFFRX1 \i_MIPS/Register/register_reg[20][17]  ( .D(\i_MIPS/Register/n485 ), 
        .CK(clk), .RN(n4099), .Q(\i_MIPS/Register/register[20][17] ) );
  DFFRX1 \i_MIPS/Register/register_reg[20][18]  ( .D(\i_MIPS/Register/n486 ), 
        .CK(clk), .RN(n4099), .Q(\i_MIPS/Register/register[20][18] ) );
  DFFRX1 \i_MIPS/Register/register_reg[20][19]  ( .D(\i_MIPS/Register/n487 ), 
        .CK(clk), .RN(n4099), .Q(\i_MIPS/Register/register[20][19] ) );
  DFFRX1 \i_MIPS/Register/register_reg[20][20]  ( .D(\i_MIPS/Register/n488 ), 
        .CK(clk), .RN(n4099), .Q(\i_MIPS/Register/register[20][20] ) );
  DFFRX1 \i_MIPS/Register/register_reg[20][21]  ( .D(\i_MIPS/Register/n489 ), 
        .CK(clk), .RN(n4099), .Q(\i_MIPS/Register/register[20][21] ) );
  DFFRX1 \i_MIPS/Register/register_reg[20][22]  ( .D(\i_MIPS/Register/n490 ), 
        .CK(clk), .RN(n4099), .Q(\i_MIPS/Register/register[20][22] ) );
  DFFRX1 \i_MIPS/Register/register_reg[20][23]  ( .D(\i_MIPS/Register/n491 ), 
        .CK(clk), .RN(n4099), .Q(\i_MIPS/Register/register[20][23] ) );
  DFFRX1 \i_MIPS/Register/register_reg[20][24]  ( .D(\i_MIPS/Register/n492 ), 
        .CK(clk), .RN(n4100), .Q(\i_MIPS/Register/register[20][24] ) );
  DFFRX1 \i_MIPS/Register/register_reg[20][25]  ( .D(\i_MIPS/Register/n493 ), 
        .CK(clk), .RN(n4100), .Q(\i_MIPS/Register/register[20][25] ) );
  DFFRX1 \i_MIPS/Register/register_reg[20][26]  ( .D(\i_MIPS/Register/n494 ), 
        .CK(clk), .RN(n4100), .Q(\i_MIPS/Register/register[20][26] ) );
  DFFRX1 \i_MIPS/Register/register_reg[20][27]  ( .D(\i_MIPS/Register/n495 ), 
        .CK(clk), .RN(n4100), .Q(\i_MIPS/Register/register[20][27] ) );
  DFFRX1 \i_MIPS/Register/register_reg[20][28]  ( .D(\i_MIPS/Register/n496 ), 
        .CK(clk), .RN(n4100), .Q(\i_MIPS/Register/register[20][28] ) );
  DFFRX1 \i_MIPS/Register/register_reg[20][29]  ( .D(\i_MIPS/Register/n497 ), 
        .CK(clk), .RN(n4100), .Q(\i_MIPS/Register/register[20][29] ) );
  DFFRX1 \i_MIPS/Register/register_reg[20][30]  ( .D(\i_MIPS/Register/n498 ), 
        .CK(clk), .RN(n4100), .Q(\i_MIPS/Register/register[20][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[20][31]  ( .D(\i_MIPS/Register/n499 ), 
        .CK(clk), .RN(n4100), .Q(\i_MIPS/Register/register[20][31] ) );
  DFFRX1 \i_MIPS/Register/register_reg[16][2]  ( .D(\i_MIPS/Register/n598 ), 
        .CK(clk), .RN(n4108), .Q(\i_MIPS/Register/register[16][2] ) );
  DFFRX1 \i_MIPS/Register/register_reg[16][3]  ( .D(\i_MIPS/Register/n599 ), 
        .CK(clk), .RN(n4108), .Q(\i_MIPS/Register/register[16][3] ) );
  DFFRX1 \i_MIPS/Register/register_reg[16][4]  ( .D(\i_MIPS/Register/n600 ), 
        .CK(clk), .RN(n4109), .Q(\i_MIPS/Register/register[16][4] ) );
  DFFRX1 \i_MIPS/Register/register_reg[16][5]  ( .D(\i_MIPS/Register/n601 ), 
        .CK(clk), .RN(n4109), .Q(\i_MIPS/Register/register[16][5] ) );
  DFFRX1 \i_MIPS/Register/register_reg[16][6]  ( .D(\i_MIPS/Register/n602 ), 
        .CK(clk), .RN(n4109), .Q(\i_MIPS/Register/register[16][6] ) );
  DFFRX1 \i_MIPS/Register/register_reg[16][7]  ( .D(\i_MIPS/Register/n603 ), 
        .CK(clk), .RN(n4109), .Q(\i_MIPS/Register/register[16][7] ) );
  DFFRX1 \i_MIPS/Register/register_reg[16][8]  ( .D(\i_MIPS/Register/n604 ), 
        .CK(clk), .RN(n4109), .Q(\i_MIPS/Register/register[16][8] ) );
  DFFRX1 \i_MIPS/Register/register_reg[16][9]  ( .D(\i_MIPS/Register/n605 ), 
        .CK(clk), .RN(n4109), .Q(\i_MIPS/Register/register[16][9] ) );
  DFFRX1 \i_MIPS/Register/register_reg[16][10]  ( .D(\i_MIPS/Register/n606 ), 
        .CK(clk), .RN(n4109), .Q(\i_MIPS/Register/register[16][10] ) );
  DFFRX1 \i_MIPS/Register/register_reg[16][11]  ( .D(\i_MIPS/Register/n607 ), 
        .CK(clk), .RN(n4109), .Q(\i_MIPS/Register/register[16][11] ) );
  DFFRX1 \i_MIPS/Register/register_reg[16][12]  ( .D(\i_MIPS/Register/n608 ), 
        .CK(clk), .RN(n4109), .Q(\i_MIPS/Register/register[16][12] ) );
  DFFRX1 \i_MIPS/Register/register_reg[16][13]  ( .D(\i_MIPS/Register/n609 ), 
        .CK(clk), .RN(n4109), .Q(\i_MIPS/Register/register[16][13] ) );
  DFFRX1 \i_MIPS/Register/register_reg[16][14]  ( .D(\i_MIPS/Register/n610 ), 
        .CK(clk), .RN(n4109), .Q(\i_MIPS/Register/register[16][14] ) );
  DFFRX1 \i_MIPS/Register/register_reg[16][15]  ( .D(\i_MIPS/Register/n611 ), 
        .CK(clk), .RN(n4109), .Q(\i_MIPS/Register/register[16][15] ) );
  DFFRX1 \i_MIPS/Register/register_reg[16][16]  ( .D(\i_MIPS/Register/n612 ), 
        .CK(clk), .RN(n4110), .Q(\i_MIPS/Register/register[16][16] ) );
  DFFRX1 \i_MIPS/Register/register_reg[16][17]  ( .D(\i_MIPS/Register/n613 ), 
        .CK(clk), .RN(n4110), .Q(\i_MIPS/Register/register[16][17] ) );
  DFFRX1 \i_MIPS/Register/register_reg[16][18]  ( .D(\i_MIPS/Register/n614 ), 
        .CK(clk), .RN(n4110), .Q(\i_MIPS/Register/register[16][18] ) );
  DFFRX1 \i_MIPS/Register/register_reg[16][19]  ( .D(\i_MIPS/Register/n615 ), 
        .CK(clk), .RN(n4110), .Q(\i_MIPS/Register/register[16][19] ) );
  DFFRX1 \i_MIPS/Register/register_reg[16][20]  ( .D(\i_MIPS/Register/n616 ), 
        .CK(clk), .RN(n4110), .Q(\i_MIPS/Register/register[16][20] ) );
  DFFRX1 \i_MIPS/Register/register_reg[16][21]  ( .D(\i_MIPS/Register/n617 ), 
        .CK(clk), .RN(n4110), .Q(\i_MIPS/Register/register[16][21] ) );
  DFFRX1 \i_MIPS/Register/register_reg[16][22]  ( .D(\i_MIPS/Register/n618 ), 
        .CK(clk), .RN(n4110), .Q(\i_MIPS/Register/register[16][22] ) );
  DFFRX1 \i_MIPS/Register/register_reg[16][23]  ( .D(\i_MIPS/Register/n619 ), 
        .CK(clk), .RN(n4110), .Q(\i_MIPS/Register/register[16][23] ) );
  DFFRX1 \i_MIPS/Register/register_reg[16][24]  ( .D(\i_MIPS/Register/n620 ), 
        .CK(clk), .RN(n4110), .Q(\i_MIPS/Register/register[16][24] ) );
  DFFRX1 \i_MIPS/Register/register_reg[16][25]  ( .D(\i_MIPS/Register/n621 ), 
        .CK(clk), .RN(n4110), .Q(\i_MIPS/Register/register[16][25] ) );
  DFFRX1 \i_MIPS/Register/register_reg[16][26]  ( .D(\i_MIPS/Register/n622 ), 
        .CK(clk), .RN(n4110), .Q(\i_MIPS/Register/register[16][26] ) );
  DFFRX1 \i_MIPS/Register/register_reg[16][27]  ( .D(\i_MIPS/Register/n623 ), 
        .CK(clk), .RN(n4110), .Q(\i_MIPS/Register/register[16][27] ) );
  DFFRX1 \i_MIPS/Register/register_reg[16][28]  ( .D(\i_MIPS/Register/n624 ), 
        .CK(clk), .RN(n4111), .Q(\i_MIPS/Register/register[16][28] ) );
  DFFRX1 \i_MIPS/Register/register_reg[16][29]  ( .D(\i_MIPS/Register/n625 ), 
        .CK(clk), .RN(n4111), .Q(\i_MIPS/Register/register[16][29] ) );
  DFFRX1 \i_MIPS/Register/register_reg[16][30]  ( .D(\i_MIPS/Register/n626 ), 
        .CK(clk), .RN(n4111), .Q(\i_MIPS/Register/register[16][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[16][31]  ( .D(\i_MIPS/Register/n627 ), 
        .CK(clk), .RN(n4111), .Q(\i_MIPS/Register/register[16][31] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][2]  ( .D(\i_MIPS/Register/n918 ), 
        .CK(clk), .RN(n4135), .Q(\i_MIPS/Register/register[6][2] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][3]  ( .D(\i_MIPS/Register/n919 ), 
        .CK(clk), .RN(n4135), .Q(\i_MIPS/Register/register[6][3] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][4]  ( .D(\i_MIPS/Register/n920 ), 
        .CK(clk), .RN(n4135), .Q(\i_MIPS/Register/register[6][4] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][6]  ( .D(\i_MIPS/Register/n922 ), 
        .CK(clk), .RN(n4135), .Q(\i_MIPS/Register/register[6][6] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][7]  ( .D(\i_MIPS/Register/n923 ), 
        .CK(clk), .RN(n4135), .Q(\i_MIPS/Register/register[6][7] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][8]  ( .D(\i_MIPS/Register/n924 ), 
        .CK(clk), .RN(n4136), .Q(\i_MIPS/Register/register[6][8] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][9]  ( .D(\i_MIPS/Register/n925 ), 
        .CK(clk), .RN(n4136), .Q(\i_MIPS/Register/register[6][9] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][10]  ( .D(\i_MIPS/Register/n926 ), 
        .CK(clk), .RN(n4136), .Q(\i_MIPS/Register/register[6][10] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][11]  ( .D(\i_MIPS/Register/n927 ), 
        .CK(clk), .RN(n4136), .Q(\i_MIPS/Register/register[6][11] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][13]  ( .D(\i_MIPS/Register/n929 ), 
        .CK(clk), .RN(n4136), .Q(\i_MIPS/Register/register[6][13] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][14]  ( .D(\i_MIPS/Register/n930 ), 
        .CK(clk), .RN(n4136), .Q(\i_MIPS/Register/register[6][14] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][15]  ( .D(\i_MIPS/Register/n931 ), 
        .CK(clk), .RN(n4136), .Q(\i_MIPS/Register/register[6][15] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][16]  ( .D(\i_MIPS/Register/n932 ), 
        .CK(clk), .RN(n4136), .Q(\i_MIPS/Register/register[6][16] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][17]  ( .D(\i_MIPS/Register/n933 ), 
        .CK(clk), .RN(n4136), .Q(\i_MIPS/Register/register[6][17] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][18]  ( .D(\i_MIPS/Register/n934 ), 
        .CK(clk), .RN(n4136), .Q(\i_MIPS/Register/register[6][18] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][19]  ( .D(\i_MIPS/Register/n935 ), 
        .CK(clk), .RN(n4136), .Q(\i_MIPS/Register/register[6][19] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][20]  ( .D(\i_MIPS/Register/n936 ), 
        .CK(clk), .RN(n4137), .Q(\i_MIPS/Register/register[6][20] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][21]  ( .D(\i_MIPS/Register/n937 ), 
        .CK(clk), .RN(n4137), .Q(\i_MIPS/Register/register[6][21] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][22]  ( .D(\i_MIPS/Register/n938 ), 
        .CK(clk), .RN(n4137), .Q(\i_MIPS/Register/register[6][22] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][23]  ( .D(\i_MIPS/Register/n939 ), 
        .CK(clk), .RN(n4137), .Q(\i_MIPS/Register/register[6][23] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][25]  ( .D(\i_MIPS/Register/n941 ), 
        .CK(clk), .RN(n4137), .Q(\i_MIPS/Register/register[6][25] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][27]  ( .D(\i_MIPS/Register/n943 ), 
        .CK(clk), .RN(n4137), .Q(\i_MIPS/Register/register[6][27] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][28]  ( .D(\i_MIPS/Register/n944 ), 
        .CK(clk), .RN(n4137), .Q(\i_MIPS/Register/register[6][28] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][29]  ( .D(\i_MIPS/Register/n945 ), 
        .CK(clk), .RN(n4137), .Q(\i_MIPS/Register/register[6][29] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][30]  ( .D(\i_MIPS/Register/n946 ), 
        .CK(clk), .RN(n4137), .Q(\i_MIPS/Register/register[6][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][31]  ( .D(\i_MIPS/Register/n947 ), 
        .CK(clk), .RN(n4137), .Q(\i_MIPS/Register/register[6][31] ) );
  DFFRX1 \i_MIPS/Register/register_reg[4][2]  ( .D(\i_MIPS/Register/n982 ), 
        .CK(clk), .RN(n4140), .Q(\i_MIPS/Register/register[4][2] ) );
  DFFRX1 \i_MIPS/Register/register_reg[4][3]  ( .D(\i_MIPS/Register/n983 ), 
        .CK(clk), .RN(n4140), .Q(\i_MIPS/Register/register[4][3] ) );
  DFFRX1 \i_MIPS/Register/register_reg[4][4]  ( .D(\i_MIPS/Register/n984 ), 
        .CK(clk), .RN(n4141), .Q(\i_MIPS/Register/register[4][4] ) );
  DFFRX1 \i_MIPS/Register/register_reg[4][6]  ( .D(\i_MIPS/Register/n986 ), 
        .CK(clk), .RN(n4141), .Q(\i_MIPS/Register/register[4][6] ) );
  DFFRX1 \i_MIPS/Register/register_reg[4][7]  ( .D(\i_MIPS/Register/n987 ), 
        .CK(clk), .RN(n4141), .Q(\i_MIPS/Register/register[4][7] ) );
  DFFRX1 \i_MIPS/Register/register_reg[4][8]  ( .D(\i_MIPS/Register/n988 ), 
        .CK(clk), .RN(n4141), .Q(\i_MIPS/Register/register[4][8] ) );
  DFFRX1 \i_MIPS/Register/register_reg[4][9]  ( .D(\i_MIPS/Register/n989 ), 
        .CK(clk), .RN(n4141), .Q(\i_MIPS/Register/register[4][9] ) );
  DFFRX1 \i_MIPS/Register/register_reg[4][10]  ( .D(\i_MIPS/Register/n990 ), 
        .CK(clk), .RN(n4141), .Q(\i_MIPS/Register/register[4][10] ) );
  DFFRX1 \i_MIPS/Register/register_reg[4][11]  ( .D(\i_MIPS/Register/n991 ), 
        .CK(clk), .RN(n4141), .Q(\i_MIPS/Register/register[4][11] ) );
  DFFRX1 \i_MIPS/Register/register_reg[4][13]  ( .D(\i_MIPS/Register/n993 ), 
        .CK(clk), .RN(n4141), .Q(\i_MIPS/Register/register[4][13] ) );
  DFFRX1 \i_MIPS/Register/register_reg[4][14]  ( .D(\i_MIPS/Register/n994 ), 
        .CK(clk), .RN(n4141), .Q(\i_MIPS/Register/register[4][14] ) );
  DFFRX1 \i_MIPS/Register/register_reg[4][15]  ( .D(\i_MIPS/Register/n995 ), 
        .CK(clk), .RN(n4141), .Q(\i_MIPS/Register/register[4][15] ) );
  DFFRX1 \i_MIPS/Register/register_reg[4][16]  ( .D(\i_MIPS/Register/n996 ), 
        .CK(clk), .RN(n4142), .Q(\i_MIPS/Register/register[4][16] ) );
  DFFRX1 \i_MIPS/Register/register_reg[4][17]  ( .D(\i_MIPS/Register/n997 ), 
        .CK(clk), .RN(n4142), .Q(\i_MIPS/Register/register[4][17] ) );
  DFFRX1 \i_MIPS/Register/register_reg[4][18]  ( .D(\i_MIPS/Register/n998 ), 
        .CK(clk), .RN(n4142), .Q(\i_MIPS/Register/register[4][18] ) );
  DFFRX1 \i_MIPS/Register/register_reg[4][19]  ( .D(\i_MIPS/Register/n999 ), 
        .CK(clk), .RN(n4142), .Q(\i_MIPS/Register/register[4][19] ) );
  DFFRX1 \i_MIPS/Register/register_reg[4][20]  ( .D(\i_MIPS/Register/n1000 ), 
        .CK(clk), .RN(n4142), .Q(\i_MIPS/Register/register[4][20] ) );
  DFFRX1 \i_MIPS/Register/register_reg[4][21]  ( .D(\i_MIPS/Register/n1001 ), 
        .CK(clk), .RN(n4142), .Q(\i_MIPS/Register/register[4][21] ) );
  DFFRX1 \i_MIPS/Register/register_reg[4][22]  ( .D(\i_MIPS/Register/n1002 ), 
        .CK(clk), .RN(n4142), .Q(\i_MIPS/Register/register[4][22] ) );
  DFFRX1 \i_MIPS/Register/register_reg[4][23]  ( .D(\i_MIPS/Register/n1003 ), 
        .CK(clk), .RN(n4142), .Q(\i_MIPS/Register/register[4][23] ) );
  DFFRX1 \i_MIPS/Register/register_reg[4][25]  ( .D(\i_MIPS/Register/n1005 ), 
        .CK(clk), .RN(n4142), .Q(\i_MIPS/Register/register[4][25] ) );
  DFFRX1 \i_MIPS/Register/register_reg[4][27]  ( .D(\i_MIPS/Register/n1007 ), 
        .CK(clk), .RN(n4142), .Q(\i_MIPS/Register/register[4][27] ) );
  DFFRX1 \i_MIPS/Register/register_reg[4][28]  ( .D(\i_MIPS/Register/n1008 ), 
        .CK(clk), .RN(n4143), .Q(\i_MIPS/Register/register[4][28] ) );
  DFFRX1 \i_MIPS/Register/register_reg[4][29]  ( .D(\i_MIPS/Register/n1009 ), 
        .CK(clk), .RN(n4143), .Q(\i_MIPS/Register/register[4][29] ) );
  DFFRX1 \i_MIPS/Register/register_reg[4][30]  ( .D(\i_MIPS/Register/n1010 ), 
        .CK(clk), .RN(n4143), .Q(\i_MIPS/Register/register[4][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[4][31]  ( .D(\i_MIPS/Register/n1011 ), 
        .CK(clk), .RN(n4143), .Q(\i_MIPS/Register/register[4][31] ) );
  DFFRX1 \i_MIPS/Register/register_reg[0][2]  ( .D(\i_MIPS/Register/n1110 ), 
        .CK(clk), .RN(n4151), .Q(\i_MIPS/Register/register[0][2] ) );
  DFFRX1 \i_MIPS/Register/register_reg[0][3]  ( .D(\i_MIPS/Register/n1111 ), 
        .CK(clk), .RN(n4151), .Q(\i_MIPS/Register/register[0][3] ) );
  DFFRX1 \i_MIPS/Register/register_reg[0][4]  ( .D(\i_MIPS/Register/n1112 ), 
        .CK(clk), .RN(n4151), .Q(\i_MIPS/Register/register[0][4] ) );
  DFFRX1 \i_MIPS/Register/register_reg[0][6]  ( .D(\i_MIPS/Register/n1114 ), 
        .CK(clk), .RN(n4151), .Q(\i_MIPS/Register/register[0][6] ) );
  DFFRX1 \i_MIPS/Register/register_reg[0][7]  ( .D(\i_MIPS/Register/n1115 ), 
        .CK(clk), .RN(n4151), .Q(\i_MIPS/Register/register[0][7] ) );
  DFFRX1 \i_MIPS/Register/register_reg[0][8]  ( .D(\i_MIPS/Register/n1116 ), 
        .CK(clk), .RN(n4152), .Q(\i_MIPS/Register/register[0][8] ) );
  DFFRX1 \i_MIPS/Register/register_reg[0][9]  ( .D(\i_MIPS/Register/n1117 ), 
        .CK(clk), .RN(n4152), .Q(\i_MIPS/Register/register[0][9] ) );
  DFFRX1 \i_MIPS/Register/register_reg[0][10]  ( .D(\i_MIPS/Register/n1118 ), 
        .CK(clk), .RN(n4152), .Q(\i_MIPS/Register/register[0][10] ) );
  DFFRX1 \i_MIPS/Register/register_reg[0][11]  ( .D(\i_MIPS/Register/n1119 ), 
        .CK(clk), .RN(n4152), .Q(\i_MIPS/Register/register[0][11] ) );
  DFFRX1 \i_MIPS/Register/register_reg[0][13]  ( .D(\i_MIPS/Register/n1121 ), 
        .CK(clk), .RN(n4152), .Q(\i_MIPS/Register/register[0][13] ) );
  DFFRX1 \i_MIPS/Register/register_reg[0][14]  ( .D(\i_MIPS/Register/n1122 ), 
        .CK(clk), .RN(n4152), .Q(\i_MIPS/Register/register[0][14] ) );
  DFFRX1 \i_MIPS/Register/register_reg[0][15]  ( .D(\i_MIPS/Register/n1123 ), 
        .CK(clk), .RN(n4152), .Q(\i_MIPS/Register/register[0][15] ) );
  DFFRX1 \i_MIPS/Register/register_reg[0][16]  ( .D(\i_MIPS/Register/n1124 ), 
        .CK(clk), .RN(n4152), .Q(\i_MIPS/Register/register[0][16] ) );
  DFFRX1 \i_MIPS/Register/register_reg[0][17]  ( .D(\i_MIPS/Register/n1125 ), 
        .CK(clk), .RN(n4152), .Q(\i_MIPS/Register/register[0][17] ) );
  DFFRX1 \i_MIPS/Register/register_reg[0][18]  ( .D(\i_MIPS/Register/n1126 ), 
        .CK(clk), .RN(n4152), .Q(\i_MIPS/Register/register[0][18] ) );
  DFFRX1 \i_MIPS/Register/register_reg[0][19]  ( .D(\i_MIPS/Register/n1127 ), 
        .CK(clk), .RN(n4152), .Q(\i_MIPS/Register/register[0][19] ) );
  DFFRX1 \i_MIPS/Register/register_reg[0][20]  ( .D(\i_MIPS/Register/n1128 ), 
        .CK(clk), .RN(n4153), .Q(\i_MIPS/Register/register[0][20] ) );
  DFFRX1 \i_MIPS/Register/register_reg[0][21]  ( .D(\i_MIPS/Register/n1129 ), 
        .CK(clk), .RN(n4153), .Q(\i_MIPS/Register/register[0][21] ) );
  DFFRX1 \i_MIPS/Register/register_reg[0][22]  ( .D(\i_MIPS/Register/n1130 ), 
        .CK(clk), .RN(n4153), .Q(\i_MIPS/Register/register[0][22] ) );
  DFFRX1 \i_MIPS/Register/register_reg[0][23]  ( .D(\i_MIPS/Register/n1131 ), 
        .CK(clk), .RN(n4153), .Q(\i_MIPS/Register/register[0][23] ) );
  DFFRX1 \i_MIPS/Register/register_reg[0][25]  ( .D(\i_MIPS/Register/n1133 ), 
        .CK(clk), .RN(n4153), .Q(\i_MIPS/Register/register[0][25] ) );
  DFFRX1 \i_MIPS/Register/register_reg[0][27]  ( .D(\i_MIPS/Register/n1135 ), 
        .CK(clk), .RN(n4153), .Q(\i_MIPS/Register/register[0][27] ) );
  DFFRX1 \i_MIPS/Register/register_reg[0][28]  ( .D(\i_MIPS/Register/n1136 ), 
        .CK(clk), .RN(n4153), .Q(\i_MIPS/Register/register[0][28] ) );
  DFFRX1 \i_MIPS/Register/register_reg[0][29]  ( .D(\i_MIPS/Register/n1137 ), 
        .CK(clk), .RN(n4153), .Q(\i_MIPS/Register/register[0][29] ) );
  DFFRX1 \i_MIPS/Register/register_reg[0][30]  ( .D(\i_MIPS/Register/n1138 ), 
        .CK(clk), .RN(n4153), .Q(\i_MIPS/Register/register[0][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[0][31]  ( .D(\i_MIPS/Register/n1139 ), 
        .CK(clk), .RN(n4153), .Q(\i_MIPS/Register/register[0][31] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][0]  ( .D(\i_MIPS/Register/n532 ), 
        .CK(clk), .RN(n4103), .Q(\i_MIPS/Register/register[18][0] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][1]  ( .D(\i_MIPS/Register/n533 ), 
        .CK(clk), .RN(n4103), .Q(\i_MIPS/Register/register[18][1] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][0]  ( .D(\i_MIPS/Register/n1044 ), 
        .CK(clk), .RN(n4146), .Q(\i_MIPS/Register/register[2][0] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][1]  ( .D(\i_MIPS/Register/n1045 ), 
        .CK(clk), .RN(n4146), .Q(\i_MIPS/Register/register[2][1] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][5]  ( .D(\i_MIPS/Register/n1049 ), 
        .CK(clk), .RN(n4146), .Q(\i_MIPS/Register/register[2][5] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][12]  ( .D(\i_MIPS/Register/n1056 ), 
        .CK(clk), .RN(n4147), .Q(\i_MIPS/Register/register[2][12] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][24]  ( .D(\i_MIPS/Register/n1068 ), 
        .CK(clk), .RN(n4148), .Q(\i_MIPS/Register/register[2][24] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][26]  ( .D(\i_MIPS/Register/n1070 ), 
        .CK(clk), .RN(n4148), .Q(\i_MIPS/Register/register[2][26] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][0]  ( .D(\i_MIPS/Register/n276 ), 
        .CK(clk), .RN(n4082), .Q(\i_MIPS/Register/register[26][0] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][1]  ( .D(\i_MIPS/Register/n277 ), 
        .CK(clk), .RN(n4082), .Q(\i_MIPS/Register/register[26][1] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][0]  ( .D(\i_MIPS/Register/n788 ), 
        .CK(clk), .RN(n4124), .Q(\i_MIPS/Register/register[10][0] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][1]  ( .D(\i_MIPS/Register/n789 ), 
        .CK(clk), .RN(n4124), .Q(\i_MIPS/Register/register[10][1] ) );
  DFFRX1 \i_MIPS/IF_ID_reg[60]  ( .D(\i_MIPS/N83 ), .CK(clk), .RN(n4062), .Q(
        \i_MIPS/IR_ID[28] ), .QN(\i_MIPS/n326 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[63]  ( .D(\i_MIPS/N86 ), .CK(clk), .RN(n4062), .Q(
        \i_MIPS/IR_ID[31] ), .QN(\i_MIPS/n332 ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][2]  ( .D(\i_MIPS/Register/n534 ), 
        .CK(clk), .RN(n4103), .Q(\i_MIPS/Register/register[18][2] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][3]  ( .D(\i_MIPS/Register/n535 ), 
        .CK(clk), .RN(n4103), .Q(\i_MIPS/Register/register[18][3] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][4]  ( .D(\i_MIPS/Register/n536 ), 
        .CK(clk), .RN(n4103), .Q(\i_MIPS/Register/register[18][4] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][5]  ( .D(\i_MIPS/Register/n537 ), 
        .CK(clk), .RN(n4103), .Q(\i_MIPS/Register/register[18][5] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][6]  ( .D(\i_MIPS/Register/n538 ), 
        .CK(clk), .RN(n4103), .Q(\i_MIPS/Register/register[18][6] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][7]  ( .D(\i_MIPS/Register/n539 ), 
        .CK(clk), .RN(n4103), .Q(\i_MIPS/Register/register[18][7] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][8]  ( .D(\i_MIPS/Register/n540 ), 
        .CK(clk), .RN(n4104), .Q(\i_MIPS/Register/register[18][8] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][9]  ( .D(\i_MIPS/Register/n541 ), 
        .CK(clk), .RN(n4104), .Q(\i_MIPS/Register/register[18][9] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][10]  ( .D(\i_MIPS/Register/n542 ), 
        .CK(clk), .RN(n4104), .Q(\i_MIPS/Register/register[18][10] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][11]  ( .D(\i_MIPS/Register/n543 ), 
        .CK(clk), .RN(n4104), .Q(\i_MIPS/Register/register[18][11] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][12]  ( .D(\i_MIPS/Register/n544 ), 
        .CK(clk), .RN(n4104), .Q(\i_MIPS/Register/register[18][12] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][13]  ( .D(\i_MIPS/Register/n545 ), 
        .CK(clk), .RN(n4104), .Q(\i_MIPS/Register/register[18][13] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][14]  ( .D(\i_MIPS/Register/n546 ), 
        .CK(clk), .RN(n4104), .Q(\i_MIPS/Register/register[18][14] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][15]  ( .D(\i_MIPS/Register/n547 ), 
        .CK(clk), .RN(n4104), .Q(\i_MIPS/Register/register[18][15] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][16]  ( .D(\i_MIPS/Register/n548 ), 
        .CK(clk), .RN(n4104), .Q(\i_MIPS/Register/register[18][16] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][17]  ( .D(\i_MIPS/Register/n549 ), 
        .CK(clk), .RN(n4104), .Q(\i_MIPS/Register/register[18][17] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][18]  ( .D(\i_MIPS/Register/n550 ), 
        .CK(clk), .RN(n4104), .Q(\i_MIPS/Register/register[18][18] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][19]  ( .D(\i_MIPS/Register/n551 ), 
        .CK(clk), .RN(n4104), .Q(\i_MIPS/Register/register[18][19] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][20]  ( .D(\i_MIPS/Register/n552 ), 
        .CK(clk), .RN(n4105), .Q(\i_MIPS/Register/register[18][20] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][21]  ( .D(\i_MIPS/Register/n553 ), 
        .CK(clk), .RN(n4105), .Q(\i_MIPS/Register/register[18][21] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][22]  ( .D(\i_MIPS/Register/n554 ), 
        .CK(clk), .RN(n4105), .Q(\i_MIPS/Register/register[18][22] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][23]  ( .D(\i_MIPS/Register/n555 ), 
        .CK(clk), .RN(n4105), .Q(\i_MIPS/Register/register[18][23] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][24]  ( .D(\i_MIPS/Register/n556 ), 
        .CK(clk), .RN(n4105), .Q(\i_MIPS/Register/register[18][24] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][25]  ( .D(\i_MIPS/Register/n557 ), 
        .CK(clk), .RN(n4105), .Q(\i_MIPS/Register/register[18][25] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][26]  ( .D(\i_MIPS/Register/n558 ), 
        .CK(clk), .RN(n4105), .Q(\i_MIPS/Register/register[18][26] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][27]  ( .D(\i_MIPS/Register/n559 ), 
        .CK(clk), .RN(n4105), .Q(\i_MIPS/Register/register[18][27] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][28]  ( .D(\i_MIPS/Register/n560 ), 
        .CK(clk), .RN(n4105), .Q(\i_MIPS/Register/register[18][28] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][29]  ( .D(\i_MIPS/Register/n561 ), 
        .CK(clk), .RN(n4105), .Q(\i_MIPS/Register/register[18][29] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][30]  ( .D(\i_MIPS/Register/n562 ), 
        .CK(clk), .RN(n4105), .Q(\i_MIPS/Register/register[18][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][31]  ( .D(\i_MIPS/Register/n563 ), 
        .CK(clk), .RN(n4105), .Q(\i_MIPS/Register/register[18][31] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][2]  ( .D(\i_MIPS/Register/n1046 ), 
        .CK(clk), .RN(n4146), .Q(\i_MIPS/Register/register[2][2] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][3]  ( .D(\i_MIPS/Register/n1047 ), 
        .CK(clk), .RN(n4146), .Q(\i_MIPS/Register/register[2][3] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][4]  ( .D(\i_MIPS/Register/n1048 ), 
        .CK(clk), .RN(n4146), .Q(\i_MIPS/Register/register[2][4] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][6]  ( .D(\i_MIPS/Register/n1050 ), 
        .CK(clk), .RN(n4146), .Q(\i_MIPS/Register/register[2][6] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][7]  ( .D(\i_MIPS/Register/n1051 ), 
        .CK(clk), .RN(n4146), .Q(\i_MIPS/Register/register[2][7] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][8]  ( .D(\i_MIPS/Register/n1052 ), 
        .CK(clk), .RN(n4146), .Q(\i_MIPS/Register/register[2][8] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][9]  ( .D(\i_MIPS/Register/n1053 ), 
        .CK(clk), .RN(n4146), .Q(\i_MIPS/Register/register[2][9] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][10]  ( .D(\i_MIPS/Register/n1054 ), 
        .CK(clk), .RN(n4146), .Q(\i_MIPS/Register/register[2][10] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][11]  ( .D(\i_MIPS/Register/n1055 ), 
        .CK(clk), .RN(n4146), .Q(\i_MIPS/Register/register[2][11] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][13]  ( .D(\i_MIPS/Register/n1057 ), 
        .CK(clk), .RN(n4147), .Q(\i_MIPS/Register/register[2][13] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][14]  ( .D(\i_MIPS/Register/n1058 ), 
        .CK(clk), .RN(n4147), .Q(\i_MIPS/Register/register[2][14] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][15]  ( .D(\i_MIPS/Register/n1059 ), 
        .CK(clk), .RN(n4147), .Q(\i_MIPS/Register/register[2][15] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][16]  ( .D(\i_MIPS/Register/n1060 ), 
        .CK(clk), .RN(n4147), .Q(\i_MIPS/Register/register[2][16] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][17]  ( .D(\i_MIPS/Register/n1061 ), 
        .CK(clk), .RN(n4147), .Q(\i_MIPS/Register/register[2][17] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][18]  ( .D(\i_MIPS/Register/n1062 ), 
        .CK(clk), .RN(n4147), .Q(\i_MIPS/Register/register[2][18] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][19]  ( .D(\i_MIPS/Register/n1063 ), 
        .CK(clk), .RN(n4147), .Q(\i_MIPS/Register/register[2][19] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][20]  ( .D(\i_MIPS/Register/n1064 ), 
        .CK(clk), .RN(n4147), .Q(\i_MIPS/Register/register[2][20] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][21]  ( .D(\i_MIPS/Register/n1065 ), 
        .CK(clk), .RN(n4147), .Q(\i_MIPS/Register/register[2][21] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][22]  ( .D(\i_MIPS/Register/n1066 ), 
        .CK(clk), .RN(n4147), .Q(\i_MIPS/Register/register[2][22] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][23]  ( .D(\i_MIPS/Register/n1067 ), 
        .CK(clk), .RN(n4147), .Q(\i_MIPS/Register/register[2][23] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][25]  ( .D(\i_MIPS/Register/n1069 ), 
        .CK(clk), .RN(n4148), .Q(\i_MIPS/Register/register[2][25] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][27]  ( .D(\i_MIPS/Register/n1071 ), 
        .CK(clk), .RN(n4148), .Q(\i_MIPS/Register/register[2][27] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][28]  ( .D(\i_MIPS/Register/n1072 ), 
        .CK(clk), .RN(n4148), .Q(\i_MIPS/Register/register[2][28] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][29]  ( .D(\i_MIPS/Register/n1073 ), 
        .CK(clk), .RN(n4148), .Q(\i_MIPS/Register/register[2][29] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][30]  ( .D(\i_MIPS/Register/n1074 ), 
        .CK(clk), .RN(n4148), .Q(\i_MIPS/Register/register[2][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][31]  ( .D(\i_MIPS/Register/n1075 ), 
        .CK(clk), .RN(n4148), .Q(\i_MIPS/Register/register[2][31] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][2]  ( .D(\i_MIPS/Register/n278 ), 
        .CK(clk), .RN(n4082), .Q(\i_MIPS/Register/register[26][2] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][3]  ( .D(\i_MIPS/Register/n279 ), 
        .CK(clk), .RN(n4082), .Q(\i_MIPS/Register/register[26][3] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][4]  ( .D(\i_MIPS/Register/n280 ), 
        .CK(clk), .RN(n4082), .Q(\i_MIPS/Register/register[26][4] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][5]  ( .D(\i_MIPS/Register/n281 ), 
        .CK(clk), .RN(n4082), .Q(\i_MIPS/Register/register[26][5] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][6]  ( .D(\i_MIPS/Register/n282 ), 
        .CK(clk), .RN(n4082), .Q(\i_MIPS/Register/register[26][6] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][7]  ( .D(\i_MIPS/Register/n283 ), 
        .CK(clk), .RN(n4082), .Q(\i_MIPS/Register/register[26][7] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][8]  ( .D(\i_MIPS/Register/n284 ), 
        .CK(clk), .RN(n4082), .Q(\i_MIPS/Register/register[26][8] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][9]  ( .D(\i_MIPS/Register/n285 ), 
        .CK(clk), .RN(n4082), .Q(\i_MIPS/Register/register[26][9] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][10]  ( .D(\i_MIPS/Register/n286 ), 
        .CK(clk), .RN(n4082), .Q(\i_MIPS/Register/register[26][10] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][11]  ( .D(\i_MIPS/Register/n287 ), 
        .CK(clk), .RN(n4082), .Q(\i_MIPS/Register/register[26][11] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][12]  ( .D(\i_MIPS/Register/n288 ), 
        .CK(clk), .RN(n4083), .Q(\i_MIPS/Register/register[26][12] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][13]  ( .D(\i_MIPS/Register/n289 ), 
        .CK(clk), .RN(n4083), .Q(\i_MIPS/Register/register[26][13] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][14]  ( .D(\i_MIPS/Register/n290 ), 
        .CK(clk), .RN(n4083), .Q(\i_MIPS/Register/register[26][14] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][15]  ( .D(\i_MIPS/Register/n291 ), 
        .CK(clk), .RN(n4083), .Q(\i_MIPS/Register/register[26][15] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][16]  ( .D(\i_MIPS/Register/n292 ), 
        .CK(clk), .RN(n4083), .Q(\i_MIPS/Register/register[26][16] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][17]  ( .D(\i_MIPS/Register/n293 ), 
        .CK(clk), .RN(n4083), .Q(\i_MIPS/Register/register[26][17] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][18]  ( .D(\i_MIPS/Register/n294 ), 
        .CK(clk), .RN(n4083), .Q(\i_MIPS/Register/register[26][18] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][19]  ( .D(\i_MIPS/Register/n295 ), 
        .CK(clk), .RN(n4083), .Q(\i_MIPS/Register/register[26][19] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][20]  ( .D(\i_MIPS/Register/n296 ), 
        .CK(clk), .RN(n4083), .Q(\i_MIPS/Register/register[26][20] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][21]  ( .D(\i_MIPS/Register/n297 ), 
        .CK(clk), .RN(n4083), .Q(\i_MIPS/Register/register[26][21] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][22]  ( .D(\i_MIPS/Register/n298 ), 
        .CK(clk), .RN(n4083), .Q(\i_MIPS/Register/register[26][22] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][23]  ( .D(\i_MIPS/Register/n299 ), 
        .CK(clk), .RN(n4083), .Q(\i_MIPS/Register/register[26][23] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][24]  ( .D(\i_MIPS/Register/n300 ), 
        .CK(clk), .RN(n4084), .Q(\i_MIPS/Register/register[26][24] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][25]  ( .D(\i_MIPS/Register/n301 ), 
        .CK(clk), .RN(n4084), .Q(\i_MIPS/Register/register[26][25] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][26]  ( .D(\i_MIPS/Register/n302 ), 
        .CK(clk), .RN(n4084), .Q(\i_MIPS/Register/register[26][26] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][27]  ( .D(\i_MIPS/Register/n303 ), 
        .CK(clk), .RN(n4084), .Q(\i_MIPS/Register/register[26][27] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][28]  ( .D(\i_MIPS/Register/n304 ), 
        .CK(clk), .RN(n4084), .Q(\i_MIPS/Register/register[26][28] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][29]  ( .D(\i_MIPS/Register/n305 ), 
        .CK(clk), .RN(n4084), .Q(\i_MIPS/Register/register[26][29] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][30]  ( .D(\i_MIPS/Register/n306 ), 
        .CK(clk), .RN(n4084), .Q(\i_MIPS/Register/register[26][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][31]  ( .D(\i_MIPS/Register/n307 ), 
        .CK(clk), .RN(n4084), .Q(\i_MIPS/Register/register[26][31] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][2]  ( .D(\i_MIPS/Register/n790 ), 
        .CK(clk), .RN(n4124), .Q(\i_MIPS/Register/register[10][2] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][3]  ( .D(\i_MIPS/Register/n791 ), 
        .CK(clk), .RN(n4124), .Q(\i_MIPS/Register/register[10][3] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][4]  ( .D(\i_MIPS/Register/n792 ), 
        .CK(clk), .RN(n4125), .Q(\i_MIPS/Register/register[10][4] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][5]  ( .D(\i_MIPS/Register/n793 ), 
        .CK(clk), .RN(n4125), .Q(\i_MIPS/Register/register[10][5] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][6]  ( .D(\i_MIPS/Register/n794 ), 
        .CK(clk), .RN(n4125), .Q(\i_MIPS/Register/register[10][6] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][7]  ( .D(\i_MIPS/Register/n795 ), 
        .CK(clk), .RN(n4125), .Q(\i_MIPS/Register/register[10][7] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][8]  ( .D(\i_MIPS/Register/n796 ), 
        .CK(clk), .RN(n4125), .Q(\i_MIPS/Register/register[10][8] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][9]  ( .D(\i_MIPS/Register/n797 ), 
        .CK(clk), .RN(n4125), .Q(\i_MIPS/Register/register[10][9] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][10]  ( .D(\i_MIPS/Register/n798 ), 
        .CK(clk), .RN(n4125), .Q(\i_MIPS/Register/register[10][10] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][11]  ( .D(\i_MIPS/Register/n799 ), 
        .CK(clk), .RN(n4125), .Q(\i_MIPS/Register/register[10][11] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][12]  ( .D(\i_MIPS/Register/n800 ), 
        .CK(clk), .RN(n4125), .Q(\i_MIPS/Register/register[10][12] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][13]  ( .D(\i_MIPS/Register/n801 ), 
        .CK(clk), .RN(n4125), .Q(\i_MIPS/Register/register[10][13] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][14]  ( .D(\i_MIPS/Register/n802 ), 
        .CK(clk), .RN(n4125), .Q(\i_MIPS/Register/register[10][14] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][15]  ( .D(\i_MIPS/Register/n803 ), 
        .CK(clk), .RN(n4125), .Q(\i_MIPS/Register/register[10][15] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][16]  ( .D(\i_MIPS/Register/n804 ), 
        .CK(clk), .RN(n4126), .Q(\i_MIPS/Register/register[10][16] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][17]  ( .D(\i_MIPS/Register/n805 ), 
        .CK(clk), .RN(n4126), .Q(\i_MIPS/Register/register[10][17] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][18]  ( .D(\i_MIPS/Register/n806 ), 
        .CK(clk), .RN(n4126), .Q(\i_MIPS/Register/register[10][18] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][19]  ( .D(\i_MIPS/Register/n807 ), 
        .CK(clk), .RN(n4126), .Q(\i_MIPS/Register/register[10][19] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][20]  ( .D(\i_MIPS/Register/n808 ), 
        .CK(clk), .RN(n4126), .Q(\i_MIPS/Register/register[10][20] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][21]  ( .D(\i_MIPS/Register/n809 ), 
        .CK(clk), .RN(n4126), .Q(\i_MIPS/Register/register[10][21] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][22]  ( .D(\i_MIPS/Register/n810 ), 
        .CK(clk), .RN(n4126), .Q(\i_MIPS/Register/register[10][22] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][23]  ( .D(\i_MIPS/Register/n811 ), 
        .CK(clk), .RN(n4126), .Q(\i_MIPS/Register/register[10][23] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][24]  ( .D(\i_MIPS/Register/n812 ), 
        .CK(clk), .RN(n4126), .Q(\i_MIPS/Register/register[10][24] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][25]  ( .D(\i_MIPS/Register/n813 ), 
        .CK(clk), .RN(n4126), .Q(\i_MIPS/Register/register[10][25] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][26]  ( .D(\i_MIPS/Register/n814 ), 
        .CK(clk), .RN(n4126), .Q(\i_MIPS/Register/register[10][26] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][27]  ( .D(\i_MIPS/Register/n815 ), 
        .CK(clk), .RN(n4126), .Q(\i_MIPS/Register/register[10][27] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][28]  ( .D(\i_MIPS/Register/n816 ), 
        .CK(clk), .RN(n4127), .Q(\i_MIPS/Register/register[10][28] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][29]  ( .D(\i_MIPS/Register/n817 ), 
        .CK(clk), .RN(n4127), .Q(\i_MIPS/Register/register[10][29] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][30]  ( .D(\i_MIPS/Register/n818 ), 
        .CK(clk), .RN(n4127), .Q(\i_MIPS/Register/register[10][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][31]  ( .D(\i_MIPS/Register/n819 ), 
        .CK(clk), .RN(n4127), .Q(\i_MIPS/Register/register[10][31] ) );
  DFFRX1 \i_MIPS/IF_ID_reg[59]  ( .D(\i_MIPS/N82 ), .CK(clk), .RN(n4061), .Q(
        \i_MIPS/IR_ID[27] ), .QN(\i_MIPS/n324 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[62]  ( .D(\i_MIPS/N85 ), .CK(clk), .RN(n4062), .Q(
        \i_MIPS/IR_ID[30] ), .QN(\i_MIPS/n330 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[61]  ( .D(\i_MIPS/N84 ), .CK(clk), .RN(n4062), .Q(
        \i_MIPS/IR_ID[29] ), .QN(\i_MIPS/n328 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[0]  ( .D(\i_MIPS/n528 ), .CK(clk), .RN(n4062), .Q(
        \i_MIPS/ID_EX_0 ), .QN(\i_MIPS/n372 ) );
  DFFRX1 \i_MIPS/Register/register_reg[31][8]  ( .D(n8796), .CK(clk), .RN(
        n4069), .QN(n196) );
  DFFRX1 \i_MIPS/ID_EX_reg[67]  ( .D(\i_MIPS/n385 ), .CK(clk), .RN(n4048), .Q(
        \i_MIPS/ID_EX[67] ), .QN(\i_MIPS/n257 ) );
  DFFRX1 \i_MIPS/Register/register_reg[29][1]  ( .D(\i_MIPS/Register/n181 ), 
        .CK(clk), .RN(n4074), .Q(\i_MIPS/Register/register[29][1] ), .QN(n273)
         );
  DFFRX1 \i_MIPS/Register/register_reg[25][1]  ( .D(\i_MIPS/Register/n309 ), 
        .CK(clk), .RN(n4084), .Q(\i_MIPS/Register/register[25][1] ), .QN(n393)
         );
  DFFRX1 \i_MIPS/Register/register_reg[21][1]  ( .D(\i_MIPS/Register/n437 ), 
        .CK(clk), .RN(n4095), .Q(\i_MIPS/Register/register[21][1] ), .QN(n1167) );
  DFFRX1 \i_MIPS/Register/register_reg[19][1]  ( .D(\i_MIPS/Register/n501 ), 
        .CK(clk), .RN(n4100), .Q(\i_MIPS/Register/register[19][1] ), .QN(n1166) );
  DFFRX1 \i_MIPS/Register/register_reg[17][1]  ( .D(\i_MIPS/Register/n565 ), 
        .CK(clk), .RN(n4106), .Q(\i_MIPS/Register/register[17][1] ), .QN(n1307) );
  DFFRX1 \i_MIPS/Register/register_reg[13][1]  ( .D(\i_MIPS/Register/n693 ), 
        .CK(clk), .RN(n4116), .Q(\i_MIPS/Register/register[13][1] ), .QN(n276)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][1]  ( .D(\i_MIPS/Register/n821 ), 
        .CK(clk), .RN(n4127), .Q(\i_MIPS/Register/register[9][1] ), .QN(n394)
         );
  DFFRX1 \i_MIPS/Register/register_reg[5][1]  ( .D(\i_MIPS/Register/n949 ), 
        .CK(clk), .RN(n4138), .Q(\i_MIPS/Register/register[5][1] ), .QN(n1170)
         );
  DFFRX1 \i_MIPS/Register/register_reg[5][5]  ( .D(\i_MIPS/Register/n953 ), 
        .CK(clk), .RN(n4138), .Q(\i_MIPS/Register/register[5][5] ), .QN(n1152)
         );
  DFFRX1 \i_MIPS/Register/register_reg[5][12]  ( .D(\i_MIPS/Register/n960 ), 
        .CK(clk), .RN(n4139), .Q(\i_MIPS/Register/register[5][12] ), .QN(n1118) );
  DFFRX1 \i_MIPS/Register/register_reg[3][1]  ( .D(\i_MIPS/Register/n1013 ), 
        .CK(clk), .RN(n4143), .Q(\i_MIPS/Register/register[3][1] ), .QN(n1169)
         );
  DFFRX1 \i_MIPS/Register/register_reg[3][5]  ( .D(\i_MIPS/Register/n1017 ), 
        .CK(clk), .RN(n4143), .Q(\i_MIPS/Register/register[3][5] ), .QN(n1151)
         );
  DFFRX1 \i_MIPS/Register/register_reg[1][1]  ( .D(\i_MIPS/Register/n1077 ), 
        .CK(clk), .RN(n4148), .Q(\i_MIPS/Register/register[1][1] ), .QN(n1308)
         );
  DFFRX1 \i_MIPS/Register/register_reg[1][5]  ( .D(\i_MIPS/Register/n1081 ), 
        .CK(clk), .RN(n4149), .Q(\i_MIPS/Register/register[1][5] ), .QN(n1302)
         );
  DFFRX1 \i_MIPS/Register/register_reg[1][12]  ( .D(\i_MIPS/Register/n1088 ), 
        .CK(clk), .RN(n4149), .Q(\i_MIPS/Register/register[1][12] ), .QN(n1292) );
  DFFRX1 \D_cache/cache_reg[3][0]  ( .D(\D_cache/n1792 ), .CK(clk), .RN(n4154), 
        .Q(\D_cache/cache[3][0] ) );
  DFFRX1 \D_cache/cache_reg[7][0]  ( .D(\D_cache/n1796 ), .CK(clk), .RN(n4154), 
        .Q(\D_cache/cache[7][0] ) );
  DFFRX1 \D_cache/cache_reg[3][1]  ( .D(\D_cache/n1785 ), .CK(clk), .RN(n4154), 
        .Q(\D_cache/cache[3][1] ) );
  DFFRX1 \D_cache/cache_reg[7][1]  ( .D(\D_cache/n1781 ), .CK(clk), .RN(n4155), 
        .Q(\D_cache/cache[7][1] ) );
  DFFRX1 \D_cache/cache_reg[3][2]  ( .D(\D_cache/n1777 ), .CK(clk), .RN(n4155), 
        .Q(\D_cache/cache[3][2] ) );
  DFFRX1 \D_cache/cache_reg[7][2]  ( .D(\D_cache/n1773 ), .CK(clk), .RN(n4155), 
        .Q(\D_cache/cache[7][2] ) );
  DFFRX1 \D_cache/cache_reg[3][3]  ( .D(\D_cache/n1769 ), .CK(clk), .RN(n4156), 
        .Q(\D_cache/cache[3][3] ) );
  DFFRX1 \D_cache/cache_reg[7][3]  ( .D(\D_cache/n1765 ), .CK(clk), .RN(n4156), 
        .Q(\D_cache/cache[7][3] ) );
  DFFRX1 \D_cache/cache_reg[3][4]  ( .D(\D_cache/n1761 ), .CK(clk), .RN(n4156), 
        .Q(\D_cache/cache[3][4] ) );
  DFFRX1 \D_cache/cache_reg[7][4]  ( .D(\D_cache/n1757 ), .CK(clk), .RN(n4157), 
        .Q(\D_cache/cache[7][4] ) );
  DFFRX1 \D_cache/cache_reg[3][5]  ( .D(\D_cache/n1753 ), .CK(clk), .RN(n4157), 
        .Q(\D_cache/cache[3][5] ) );
  DFFRX1 \D_cache/cache_reg[7][5]  ( .D(\D_cache/n1749 ), .CK(clk), .RN(n4157), 
        .Q(\D_cache/cache[7][5] ) );
  DFFRX1 \D_cache/cache_reg[3][6]  ( .D(\D_cache/n1745 ), .CK(clk), .RN(n4158), 
        .Q(\D_cache/cache[3][6] ) );
  DFFRX1 \D_cache/cache_reg[7][6]  ( .D(\D_cache/n1741 ), .CK(clk), .RN(n4158), 
        .Q(\D_cache/cache[7][6] ) );
  DFFRX1 \D_cache/cache_reg[3][7]  ( .D(\D_cache/n1737 ), .CK(clk), .RN(n4158), 
        .Q(\D_cache/cache[3][7] ) );
  DFFRX1 \D_cache/cache_reg[7][7]  ( .D(\D_cache/n1733 ), .CK(clk), .RN(n4159), 
        .Q(\D_cache/cache[7][7] ) );
  DFFRX1 \D_cache/cache_reg[3][8]  ( .D(\D_cache/n1729 ), .CK(clk), .RN(n4159), 
        .Q(\D_cache/cache[3][8] ) );
  DFFRX1 \D_cache/cache_reg[7][8]  ( .D(\D_cache/n1725 ), .CK(clk), .RN(n4159), 
        .Q(\D_cache/cache[7][8] ) );
  DFFRX1 \D_cache/cache_reg[3][9]  ( .D(\D_cache/n1721 ), .CK(clk), .RN(n4160), 
        .Q(\D_cache/cache[3][9] ) );
  DFFRX1 \D_cache/cache_reg[7][9]  ( .D(\D_cache/n1717 ), .CK(clk), .RN(n4160), 
        .Q(\D_cache/cache[7][9] ) );
  DFFRX1 \D_cache/cache_reg[3][10]  ( .D(\D_cache/n1713 ), .CK(clk), .RN(n4160), .Q(\D_cache/cache[3][10] ) );
  DFFRX1 \D_cache/cache_reg[7][10]  ( .D(\D_cache/n1709 ), .CK(clk), .RN(n4161), .Q(\D_cache/cache[7][10] ) );
  DFFRX1 \D_cache/cache_reg[3][11]  ( .D(\D_cache/n1705 ), .CK(clk), .RN(n4161), .Q(\D_cache/cache[3][11] ) );
  DFFRX1 \D_cache/cache_reg[7][11]  ( .D(\D_cache/n1701 ), .CK(clk), .RN(n4161), .Q(\D_cache/cache[7][11] ) );
  DFFRX1 \D_cache/cache_reg[3][12]  ( .D(\D_cache/n1697 ), .CK(clk), .RN(n4162), .Q(\D_cache/cache[3][12] ) );
  DFFRX1 \D_cache/cache_reg[7][12]  ( .D(\D_cache/n1693 ), .CK(clk), .RN(n4162), .Q(\D_cache/cache[7][12] ) );
  DFFRX1 \D_cache/cache_reg[3][13]  ( .D(\D_cache/n1689 ), .CK(clk), .RN(n4162), .Q(\D_cache/cache[3][13] ) );
  DFFRX1 \D_cache/cache_reg[7][13]  ( .D(\D_cache/n1685 ), .CK(clk), .RN(n4163), .Q(\D_cache/cache[7][13] ) );
  DFFRX1 \D_cache/cache_reg[3][14]  ( .D(\D_cache/n1681 ), .CK(clk), .RN(n4163), .Q(\D_cache/cache[3][14] ) );
  DFFRX1 \D_cache/cache_reg[7][14]  ( .D(\D_cache/n1677 ), .CK(clk), .RN(n4163), .Q(\D_cache/cache[7][14] ) );
  DFFRX1 \D_cache/cache_reg[7][15]  ( .D(\D_cache/n1669 ), .CK(clk), .RN(n4164), .Q(\D_cache/cache[7][15] ) );
  DFFRX1 \D_cache/cache_reg[3][17]  ( .D(\D_cache/n1657 ), .CK(clk), .RN(n4165), .Q(\D_cache/cache[3][17] ) );
  DFFRX1 \D_cache/cache_reg[7][17]  ( .D(\D_cache/n1653 ), .CK(clk), .RN(n4165), .Q(\D_cache/cache[7][17] ) );
  DFFRX1 \D_cache/cache_reg[3][18]  ( .D(\D_cache/n1649 ), .CK(clk), .RN(n4166), .Q(\D_cache/cache[3][18] ) );
  DFFRX1 \D_cache/cache_reg[7][18]  ( .D(\D_cache/n1645 ), .CK(clk), .RN(n4166), .Q(\D_cache/cache[7][18] ) );
  DFFRX1 \D_cache/cache_reg[3][19]  ( .D(\D_cache/n1641 ), .CK(clk), .RN(n4166), .Q(\D_cache/cache[3][19] ) );
  DFFRX1 \D_cache/cache_reg[7][19]  ( .D(\D_cache/n1637 ), .CK(clk), .RN(n4167), .Q(\D_cache/cache[7][19] ) );
  DFFRX1 \D_cache/cache_reg[3][20]  ( .D(\D_cache/n1633 ), .CK(clk), .RN(n4167), .Q(\D_cache/cache[3][20] ) );
  DFFRX1 \D_cache/cache_reg[7][20]  ( .D(\D_cache/n1629 ), .CK(clk), .RN(n4167), .Q(\D_cache/cache[7][20] ) );
  DFFRX1 \D_cache/cache_reg[3][21]  ( .D(\D_cache/n1625 ), .CK(clk), .RN(n4168), .Q(\D_cache/cache[3][21] ) );
  DFFRX1 \D_cache/cache_reg[7][21]  ( .D(\D_cache/n1621 ), .CK(clk), .RN(n4168), .Q(\D_cache/cache[7][21] ) );
  DFFRX1 \D_cache/cache_reg[3][22]  ( .D(\D_cache/n1617 ), .CK(clk), .RN(n4168), .Q(\D_cache/cache[3][22] ) );
  DFFRX1 \D_cache/cache_reg[7][22]  ( .D(\D_cache/n1613 ), .CK(clk), .RN(n4169), .Q(\D_cache/cache[7][22] ) );
  DFFRX1 \D_cache/cache_reg[3][23]  ( .D(\D_cache/n1609 ), .CK(clk), .RN(n4169), .Q(\D_cache/cache[3][23] ) );
  DFFRX1 \D_cache/cache_reg[7][23]  ( .D(\D_cache/n1605 ), .CK(clk), .RN(n4169), .Q(\D_cache/cache[7][23] ) );
  DFFRX1 \D_cache/cache_reg[3][24]  ( .D(\D_cache/n1601 ), .CK(clk), .RN(n4170), .Q(\D_cache/cache[3][24] ) );
  DFFRX1 \D_cache/cache_reg[7][24]  ( .D(\D_cache/n1597 ), .CK(clk), .RN(n4170), .Q(\D_cache/cache[7][24] ) );
  DFFRX1 \D_cache/cache_reg[3][25]  ( .D(\D_cache/n1593 ), .CK(clk), .RN(n4170), .Q(\D_cache/cache[3][25] ) );
  DFFRX1 \D_cache/cache_reg[7][25]  ( .D(\D_cache/n1589 ), .CK(clk), .RN(n4171), .Q(\D_cache/cache[7][25] ) );
  DFFRX1 \D_cache/cache_reg[3][26]  ( .D(\D_cache/n1585 ), .CK(clk), .RN(n4171), .Q(\D_cache/cache[3][26] ) );
  DFFRX1 \D_cache/cache_reg[7][26]  ( .D(\D_cache/n1581 ), .CK(clk), .RN(n4171), .Q(\D_cache/cache[7][26] ) );
  DFFRX1 \D_cache/cache_reg[3][27]  ( .D(\D_cache/n1577 ), .CK(clk), .RN(n4172), .Q(\D_cache/cache[3][27] ) );
  DFFRX1 \D_cache/cache_reg[7][27]  ( .D(\D_cache/n1573 ), .CK(clk), .RN(n4172), .Q(\D_cache/cache[7][27] ) );
  DFFRX1 \D_cache/cache_reg[3][28]  ( .D(\D_cache/n1569 ), .CK(clk), .RN(n4172), .Q(\D_cache/cache[3][28] ) );
  DFFRX1 \D_cache/cache_reg[7][28]  ( .D(\D_cache/n1565 ), .CK(clk), .RN(n4173), .Q(\D_cache/cache[7][28] ) );
  DFFRX1 \D_cache/cache_reg[3][31]  ( .D(\D_cache/n1545 ), .CK(clk), .RN(n4174), .Q(\D_cache/cache[3][31] ) );
  DFFRX1 \D_cache/cache_reg[7][31]  ( .D(\D_cache/n1541 ), .CK(clk), .RN(n4175), .Q(\D_cache/cache[7][31] ) );
  DFFRX1 \D_cache/cache_reg[3][39]  ( .D(\D_cache/n1481 ), .CK(clk), .RN(n4180), .Q(\D_cache/cache[3][39] ) );
  DFFRX1 \D_cache/cache_reg[7][39]  ( .D(\D_cache/n1477 ), .CK(clk), .RN(n4180), .Q(\D_cache/cache[7][39] ) );
  DFFRX1 \D_cache/cache_reg[3][41]  ( .D(\D_cache/n1465 ), .CK(clk), .RN(n4181), .Q(\D_cache/cache[3][41] ) );
  DFFRX1 \D_cache/cache_reg[7][41]  ( .D(\D_cache/n1461 ), .CK(clk), .RN(n4181), .Q(\D_cache/cache[7][41] ) );
  DFFRX1 \D_cache/cache_reg[3][43]  ( .D(\D_cache/n1449 ), .CK(clk), .RN(n4182), .Q(\D_cache/cache[3][43] ) );
  DFFRX1 \D_cache/cache_reg[7][43]  ( .D(\D_cache/n1445 ), .CK(clk), .RN(n4183), .Q(\D_cache/cache[7][43] ) );
  DFFRX1 \D_cache/cache_reg[3][45]  ( .D(\D_cache/n1433 ), .CK(clk), .RN(n4184), .Q(\D_cache/cache[3][45] ) );
  DFFRX1 \D_cache/cache_reg[7][45]  ( .D(\D_cache/n1429 ), .CK(clk), .RN(n4184), .Q(\D_cache/cache[7][45] ) );
  DFFRX1 \D_cache/cache_reg[3][53]  ( .D(\D_cache/n1369 ), .CK(clk), .RN(n4189), .Q(\D_cache/cache[3][53] ) );
  DFFRX1 \D_cache/cache_reg[3][54]  ( .D(\D_cache/n1361 ), .CK(clk), .RN(n4190), .Q(\D_cache/cache[3][54] ) );
  DFFRX1 \D_cache/cache_reg[7][54]  ( .D(\D_cache/n1357 ), .CK(clk), .RN(n4190), .Q(\D_cache/cache[7][54] ) );
  DFFRX1 \D_cache/cache_reg[3][69]  ( .D(\D_cache/n1241 ), .CK(clk), .RN(n4200), .Q(\D_cache/cache[3][69] ) );
  DFFRX1 \D_cache/cache_reg[7][69]  ( .D(\D_cache/n1237 ), .CK(clk), .RN(n4200), .Q(\D_cache/cache[7][69] ) );
  DFFRX1 \D_cache/cache_reg[3][70]  ( .D(\D_cache/n1233 ), .CK(clk), .RN(n4200), .Q(\D_cache/cache[3][70] ) );
  DFFRX1 \D_cache/cache_reg[7][70]  ( .D(\D_cache/n1229 ), .CK(clk), .RN(n4201), .Q(\D_cache/cache[7][70] ) );
  DFFRX1 \D_cache/cache_reg[3][71]  ( .D(\D_cache/n1225 ), .CK(clk), .RN(n4201), .Q(\D_cache/cache[3][71] ) );
  DFFRX1 \D_cache/cache_reg[7][71]  ( .D(\D_cache/n1221 ), .CK(clk), .RN(n4201), .Q(\D_cache/cache[7][71] ) );
  DFFRX1 \D_cache/cache_reg[3][72]  ( .D(\D_cache/n1217 ), .CK(clk), .RN(n4202), .Q(\D_cache/cache[3][72] ) );
  DFFRX1 \D_cache/cache_reg[7][72]  ( .D(\D_cache/n1213 ), .CK(clk), .RN(n4202), .Q(\D_cache/cache[7][72] ) );
  DFFRX1 \D_cache/cache_reg[3][73]  ( .D(\D_cache/n1209 ), .CK(clk), .RN(n4202), .Q(\D_cache/cache[3][73] ) );
  DFFRX1 \D_cache/cache_reg[7][73]  ( .D(\D_cache/n1205 ), .CK(clk), .RN(n4203), .Q(\D_cache/cache[7][73] ) );
  DFFRX1 \D_cache/cache_reg[7][74]  ( .D(\D_cache/n1197 ), .CK(clk), .RN(n4203), .Q(\D_cache/cache[7][74] ) );
  DFFRX1 \D_cache/cache_reg[3][75]  ( .D(\D_cache/n1193 ), .CK(clk), .RN(n4204), .Q(\D_cache/cache[3][75] ) );
  DFFRX1 \D_cache/cache_reg[7][75]  ( .D(\D_cache/n1189 ), .CK(clk), .RN(n4204), .Q(\D_cache/cache[7][75] ) );
  DFFRX1 \D_cache/cache_reg[3][76]  ( .D(\D_cache/n1185 ), .CK(clk), .RN(n4204), .Q(\D_cache/cache[3][76] ) );
  DFFRX1 \D_cache/cache_reg[7][76]  ( .D(\D_cache/n1181 ), .CK(clk), .RN(n4205), .Q(\D_cache/cache[7][76] ) );
  DFFRX1 \D_cache/cache_reg[3][77]  ( .D(\D_cache/n1177 ), .CK(clk), .RN(n4205), .Q(\D_cache/cache[3][77] ) );
  DFFRX1 \D_cache/cache_reg[7][77]  ( .D(\D_cache/n1173 ), .CK(clk), .RN(n4205), .Q(\D_cache/cache[7][77] ) );
  DFFRX1 \D_cache/cache_reg[3][96]  ( .D(\D_cache/n1025 ), .CK(clk), .RN(n4218), .Q(\D_cache/cache[3][96] ) );
  DFFRX1 \D_cache/cache_reg[7][96]  ( .D(\D_cache/n1021 ), .CK(clk), .RN(n4218), .Q(\D_cache/cache[7][96] ) );
  DFFRX1 \D_cache/cache_reg[3][98]  ( .D(\D_cache/n1009 ), .CK(clk), .RN(n4219), .Q(\D_cache/cache[3][98] ) );
  DFFRX1 \D_cache/cache_reg[7][98]  ( .D(\D_cache/n1005 ), .CK(clk), .RN(n4219), .Q(\D_cache/cache[7][98] ) );
  DFFRX1 \D_cache/cache_reg[3][100]  ( .D(\D_cache/n993 ), .CK(clk), .RN(n4220), .Q(\D_cache/cache[3][100] ) );
  DFFRX1 \D_cache/cache_reg[7][100]  ( .D(\D_cache/n989 ), .CK(clk), .RN(n4221), .Q(\D_cache/cache[7][100] ) );
  DFFRX1 \D_cache/cache_reg[3][101]  ( .D(\D_cache/n985 ), .CK(clk), .RN(n4221), .Q(\D_cache/cache[3][101] ) );
  DFFRX1 \D_cache/cache_reg[7][101]  ( .D(\D_cache/n981 ), .CK(clk), .RN(n4221), .Q(\D_cache/cache[7][101] ) );
  DFFRX1 \D_cache/cache_reg[3][102]  ( .D(\D_cache/n977 ), .CK(clk), .RN(n4222), .Q(\D_cache/cache[3][102] ) );
  DFFRX1 \D_cache/cache_reg[7][102]  ( .D(\D_cache/n973 ), .CK(clk), .RN(n4222), .Q(\D_cache/cache[7][102] ) );
  DFFRX1 \D_cache/cache_reg[3][103]  ( .D(\D_cache/n969 ), .CK(clk), .RN(n4222), .Q(\D_cache/cache[3][103] ) );
  DFFRX1 \D_cache/cache_reg[7][103]  ( .D(\D_cache/n965 ), .CK(clk), .RN(n4223), .Q(\D_cache/cache[7][103] ) );
  DFFRX1 \D_cache/cache_reg[3][104]  ( .D(\D_cache/n961 ), .CK(clk), .RN(n4223), .Q(\D_cache/cache[3][104] ) );
  DFFRX1 \D_cache/cache_reg[7][104]  ( .D(\D_cache/n957 ), .CK(clk), .RN(n4223), .Q(\D_cache/cache[7][104] ) );
  DFFRX1 \D_cache/cache_reg[3][105]  ( .D(\D_cache/n953 ), .CK(clk), .RN(n4224), .Q(\D_cache/cache[3][105] ) );
  DFFRX1 \D_cache/cache_reg[7][105]  ( .D(\D_cache/n949 ), .CK(clk), .RN(n4224), .Q(\D_cache/cache[7][105] ) );
  DFFRX1 \D_cache/cache_reg[3][106]  ( .D(\D_cache/n945 ), .CK(clk), .RN(n4224), .Q(\D_cache/cache[3][106] ) );
  DFFRX1 \D_cache/cache_reg[7][106]  ( .D(\D_cache/n941 ), .CK(clk), .RN(n4225), .Q(\D_cache/cache[7][106] ) );
  DFFRX1 \D_cache/cache_reg[3][107]  ( .D(\D_cache/n937 ), .CK(clk), .RN(n4225), .Q(\D_cache/cache[3][107] ) );
  DFFRX1 \D_cache/cache_reg[7][107]  ( .D(\D_cache/n933 ), .CK(clk), .RN(n4225), .Q(\D_cache/cache[7][107] ) );
  DFFRX1 \D_cache/cache_reg[3][108]  ( .D(\D_cache/n929 ), .CK(clk), .RN(n4226), .Q(\D_cache/cache[3][108] ) );
  DFFRX1 \D_cache/cache_reg[7][108]  ( .D(\D_cache/n925 ), .CK(clk), .RN(n4226), .Q(\D_cache/cache[7][108] ) );
  DFFRX1 \D_cache/cache_reg[3][109]  ( .D(\D_cache/n921 ), .CK(clk), .RN(n4226), .Q(\D_cache/cache[3][109] ) );
  DFFRX1 \D_cache/cache_reg[7][109]  ( .D(\D_cache/n917 ), .CK(clk), .RN(n4227), .Q(\D_cache/cache[7][109] ) );
  DFFRX1 \D_cache/cache_reg[3][110]  ( .D(\D_cache/n913 ), .CK(clk), .RN(n4227), .Q(\D_cache/cache[3][110] ) );
  DFFRX1 \D_cache/cache_reg[7][110]  ( .D(\D_cache/n909 ), .CK(clk), .RN(n4227), .Q(\D_cache/cache[7][110] ) );
  DFFRX1 \D_cache/cache_reg[3][118]  ( .D(\D_cache/n849 ), .CK(clk), .RN(n4232), .Q(\D_cache/cache[3][118] ) );
  DFFRX1 \D_cache/cache_reg[7][118]  ( .D(\D_cache/n845 ), .CK(clk), .RN(n4233), .Q(\D_cache/cache[7][118] ) );
  DFFRX1 \D_cache/cache_reg[3][135]  ( .D(\D_cache/n713 ), .CK(clk), .RN(n4244), .Q(\D_cache/cache[3][135] ) );
  DFFRX1 \D_cache/cache_reg[7][135]  ( .D(\D_cache/n709 ), .CK(clk), .RN(n4244), .Q(\D_cache/cache[7][135] ) );
  DFFRX1 \D_cache/cache_reg[3][136]  ( .D(\D_cache/n705 ), .CK(clk), .RN(n4244), .Q(\D_cache/cache[3][136] ) );
  DFFRX1 \D_cache/cache_reg[7][136]  ( .D(\D_cache/n701 ), .CK(clk), .RN(n4245), .Q(\D_cache/cache[7][136] ) );
  DFFRX1 \D_cache/cache_reg[3][137]  ( .D(\D_cache/n697 ), .CK(clk), .RN(n4245), .Q(\D_cache/cache[3][137] ) );
  DFFRX1 \D_cache/cache_reg[7][137]  ( .D(\D_cache/n693 ), .CK(clk), .RN(n4245), .Q(\D_cache/cache[7][137] ) );
  DFFRX1 \D_cache/cache_reg[7][139]  ( .D(\D_cache/n677 ), .CK(clk), .RN(n4247), .Q(\D_cache/cache[7][139] ) );
  DFFRX1 \D_cache/cache_reg[3][149]  ( .D(\D_cache/n601 ), .CK(clk), .RN(n4253), .Q(\D_cache/cache[3][149] ) );
  DFFRX1 \D_cache/cache_reg[7][149]  ( .D(\D_cache/n597 ), .CK(clk), .RN(n4253), .Q(\D_cache/cache[7][149] ) );
  DFFRX1 \D_cache/cache_reg[7][151]  ( .D(\D_cache/n581 ), .CK(clk), .RN(n4255), .Q(\D_cache/cache[7][151] ) );
  DFFRX1 \D_cache/cache_reg[3][153]  ( .D(\D_cache/n569 ), .CK(clk), .RN(n4256), .Q(\D_cache/cache[3][153] ) );
  DFFRX1 \D_cache/cache_reg[7][153]  ( .D(\D_cache/n565 ), .CK(clk), .RN(n4256), .Q(\D_cache/cache[7][153] ) );
  DFFRX1 \D_cache/cache_reg[3][154]  ( .D(\D_cache/n561 ), .CK(clk), .RN(n4256), .Q(\D_cache/cache[3][154] ) );
  DFFRX1 \D_cache/cache_reg[7][154]  ( .D(\D_cache/n557 ), .CK(clk), .RN(n4257), .Q(\D_cache/cache[7][154] ) );
  DFFRX1 \D_cache/cache_reg[1][0]  ( .D(\D_cache/n1794 ), .CK(clk), .RN(n4154), 
        .Q(\D_cache/cache[1][0] ) );
  DFFRX1 \D_cache/cache_reg[5][0]  ( .D(\D_cache/n1790 ), .CK(clk), .RN(n4154), 
        .Q(\D_cache/cache[5][0] ) );
  DFFRX1 \D_cache/cache_reg[1][1]  ( .D(\D_cache/n1787 ), .CK(clk), .RN(n4154), 
        .Q(\D_cache/cache[1][1] ) );
  DFFRX1 \D_cache/cache_reg[5][1]  ( .D(\D_cache/n1783 ), .CK(clk), .RN(n4155), 
        .Q(\D_cache/cache[5][1] ) );
  DFFRX1 \D_cache/cache_reg[1][2]  ( .D(\D_cache/n1779 ), .CK(clk), .RN(n4155), 
        .Q(\D_cache/cache[1][2] ) );
  DFFRX1 \D_cache/cache_reg[5][2]  ( .D(\D_cache/n1775 ), .CK(clk), .RN(n4155), 
        .Q(\D_cache/cache[5][2] ) );
  DFFRX1 \D_cache/cache_reg[1][3]  ( .D(\D_cache/n1771 ), .CK(clk), .RN(n4156), 
        .Q(\D_cache/cache[1][3] ) );
  DFFRX1 \D_cache/cache_reg[5][3]  ( .D(\D_cache/n1767 ), .CK(clk), .RN(n4156), 
        .Q(\D_cache/cache[5][3] ) );
  DFFRX1 \D_cache/cache_reg[1][4]  ( .D(\D_cache/n1763 ), .CK(clk), .RN(n4156), 
        .Q(\D_cache/cache[1][4] ) );
  DFFRX1 \D_cache/cache_reg[5][4]  ( .D(\D_cache/n1759 ), .CK(clk), .RN(n4157), 
        .Q(\D_cache/cache[5][4] ) );
  DFFRX1 \D_cache/cache_reg[1][5]  ( .D(\D_cache/n1755 ), .CK(clk), .RN(n4157), 
        .Q(\D_cache/cache[1][5] ) );
  DFFRX1 \D_cache/cache_reg[5][5]  ( .D(\D_cache/n1751 ), .CK(clk), .RN(n4157), 
        .Q(\D_cache/cache[5][5] ) );
  DFFRX1 \D_cache/cache_reg[1][6]  ( .D(\D_cache/n1747 ), .CK(clk), .RN(n4158), 
        .Q(\D_cache/cache[1][6] ) );
  DFFRX1 \D_cache/cache_reg[5][6]  ( .D(\D_cache/n1743 ), .CK(clk), .RN(n4158), 
        .Q(\D_cache/cache[5][6] ) );
  DFFRX1 \D_cache/cache_reg[1][7]  ( .D(\D_cache/n1739 ), .CK(clk), .RN(n4158), 
        .Q(\D_cache/cache[1][7] ) );
  DFFRX1 \D_cache/cache_reg[5][7]  ( .D(\D_cache/n1735 ), .CK(clk), .RN(n4159), 
        .Q(\D_cache/cache[5][7] ) );
  DFFRX1 \D_cache/cache_reg[1][8]  ( .D(\D_cache/n1731 ), .CK(clk), .RN(n4159), 
        .Q(\D_cache/cache[1][8] ) );
  DFFRX1 \D_cache/cache_reg[5][8]  ( .D(\D_cache/n1727 ), .CK(clk), .RN(n4159), 
        .Q(\D_cache/cache[5][8] ) );
  DFFRX1 \D_cache/cache_reg[1][9]  ( .D(\D_cache/n1723 ), .CK(clk), .RN(n4160), 
        .Q(\D_cache/cache[1][9] ) );
  DFFRX1 \D_cache/cache_reg[5][9]  ( .D(\D_cache/n1719 ), .CK(clk), .RN(n4160), 
        .Q(\D_cache/cache[5][9] ) );
  DFFRX1 \D_cache/cache_reg[1][10]  ( .D(\D_cache/n1715 ), .CK(clk), .RN(n4160), .Q(\D_cache/cache[1][10] ) );
  DFFRX1 \D_cache/cache_reg[5][10]  ( .D(\D_cache/n1711 ), .CK(clk), .RN(n4161), .Q(\D_cache/cache[5][10] ) );
  DFFRX1 \D_cache/cache_reg[1][11]  ( .D(\D_cache/n1707 ), .CK(clk), .RN(n4161), .Q(\D_cache/cache[1][11] ) );
  DFFRX1 \D_cache/cache_reg[5][11]  ( .D(\D_cache/n1703 ), .CK(clk), .RN(n4161), .Q(\D_cache/cache[5][11] ) );
  DFFRX1 \D_cache/cache_reg[1][12]  ( .D(\D_cache/n1699 ), .CK(clk), .RN(n4162), .Q(\D_cache/cache[1][12] ) );
  DFFRX1 \D_cache/cache_reg[5][12]  ( .D(\D_cache/n1695 ), .CK(clk), .RN(n4162), .Q(\D_cache/cache[5][12] ) );
  DFFRX1 \D_cache/cache_reg[1][13]  ( .D(\D_cache/n1691 ), .CK(clk), .RN(n4162), .Q(\D_cache/cache[1][13] ) );
  DFFRX1 \D_cache/cache_reg[5][13]  ( .D(\D_cache/n1687 ), .CK(clk), .RN(n4163), .Q(\D_cache/cache[5][13] ) );
  DFFRX1 \D_cache/cache_reg[1][14]  ( .D(\D_cache/n1683 ), .CK(clk), .RN(n4163), .Q(\D_cache/cache[1][14] ) );
  DFFRX1 \D_cache/cache_reg[5][14]  ( .D(\D_cache/n1679 ), .CK(clk), .RN(n4163), .Q(\D_cache/cache[5][14] ) );
  DFFRX1 \D_cache/cache_reg[1][15]  ( .D(\D_cache/n1675 ), .CK(clk), .RN(n4164), .Q(\D_cache/cache[1][15] ) );
  DFFRX1 \D_cache/cache_reg[5][15]  ( .D(\D_cache/n1671 ), .CK(clk), .RN(n4164), .Q(\D_cache/cache[5][15] ) );
  DFFRX1 \D_cache/cache_reg[1][17]  ( .D(\D_cache/n1659 ), .CK(clk), .RN(n4165), .Q(\D_cache/cache[1][17] ) );
  DFFRX1 \D_cache/cache_reg[5][17]  ( .D(\D_cache/n1655 ), .CK(clk), .RN(n4165), .Q(\D_cache/cache[5][17] ) );
  DFFRX1 \D_cache/cache_reg[1][18]  ( .D(\D_cache/n1651 ), .CK(clk), .RN(n4166), .Q(\D_cache/cache[1][18] ) );
  DFFRX1 \D_cache/cache_reg[5][18]  ( .D(\D_cache/n1647 ), .CK(clk), .RN(n4166), .Q(\D_cache/cache[5][18] ) );
  DFFRX1 \D_cache/cache_reg[1][19]  ( .D(\D_cache/n1643 ), .CK(clk), .RN(n4166), .Q(\D_cache/cache[1][19] ) );
  DFFRX1 \D_cache/cache_reg[5][19]  ( .D(\D_cache/n1639 ), .CK(clk), .RN(n4167), .Q(\D_cache/cache[5][19] ) );
  DFFRX1 \D_cache/cache_reg[1][20]  ( .D(\D_cache/n1635 ), .CK(clk), .RN(n4167), .Q(\D_cache/cache[1][20] ) );
  DFFRX1 \D_cache/cache_reg[5][20]  ( .D(\D_cache/n1631 ), .CK(clk), .RN(n4167), .Q(\D_cache/cache[5][20] ) );
  DFFRX1 \D_cache/cache_reg[1][21]  ( .D(\D_cache/n1627 ), .CK(clk), .RN(n4168), .Q(\D_cache/cache[1][21] ) );
  DFFRX1 \D_cache/cache_reg[5][21]  ( .D(\D_cache/n1623 ), .CK(clk), .RN(n4168), .Q(\D_cache/cache[5][21] ) );
  DFFRX1 \D_cache/cache_reg[1][22]  ( .D(\D_cache/n1619 ), .CK(clk), .RN(n4168), .Q(\D_cache/cache[1][22] ) );
  DFFRX1 \D_cache/cache_reg[5][22]  ( .D(\D_cache/n1615 ), .CK(clk), .RN(n4169), .Q(\D_cache/cache[5][22] ) );
  DFFRX1 \D_cache/cache_reg[1][23]  ( .D(\D_cache/n1611 ), .CK(clk), .RN(n4169), .Q(\D_cache/cache[1][23] ) );
  DFFRX1 \D_cache/cache_reg[5][23]  ( .D(\D_cache/n1607 ), .CK(clk), .RN(n4169), .Q(\D_cache/cache[5][23] ) );
  DFFRX1 \D_cache/cache_reg[1][24]  ( .D(\D_cache/n1603 ), .CK(clk), .RN(n4170), .Q(\D_cache/cache[1][24] ) );
  DFFRX1 \D_cache/cache_reg[5][24]  ( .D(\D_cache/n1599 ), .CK(clk), .RN(n4170), .Q(\D_cache/cache[5][24] ) );
  DFFRX1 \D_cache/cache_reg[1][25]  ( .D(\D_cache/n1595 ), .CK(clk), .RN(n4170), .Q(\D_cache/cache[1][25] ) );
  DFFRX1 \D_cache/cache_reg[5][25]  ( .D(\D_cache/n1591 ), .CK(clk), .RN(n4171), .Q(\D_cache/cache[5][25] ) );
  DFFRX1 \D_cache/cache_reg[1][26]  ( .D(\D_cache/n1587 ), .CK(clk), .RN(n4171), .Q(\D_cache/cache[1][26] ) );
  DFFRX1 \D_cache/cache_reg[5][26]  ( .D(\D_cache/n1583 ), .CK(clk), .RN(n4171), .Q(\D_cache/cache[5][26] ) );
  DFFRX1 \D_cache/cache_reg[1][27]  ( .D(\D_cache/n1579 ), .CK(clk), .RN(n4172), .Q(\D_cache/cache[1][27] ) );
  DFFRX1 \D_cache/cache_reg[5][27]  ( .D(\D_cache/n1575 ), .CK(clk), .RN(n4172), .Q(\D_cache/cache[5][27] ) );
  DFFRX1 \D_cache/cache_reg[1][28]  ( .D(\D_cache/n1571 ), .CK(clk), .RN(n4172), .Q(\D_cache/cache[1][28] ) );
  DFFRX1 \D_cache/cache_reg[5][28]  ( .D(\D_cache/n1567 ), .CK(clk), .RN(n4173), .Q(\D_cache/cache[5][28] ) );
  DFFRX1 \D_cache/cache_reg[1][31]  ( .D(\D_cache/n1547 ), .CK(clk), .RN(n4174), .Q(\D_cache/cache[1][31] ) );
  DFFRX1 \D_cache/cache_reg[5][31]  ( .D(\D_cache/n1543 ), .CK(clk), .RN(n4175), .Q(\D_cache/cache[5][31] ) );
  DFFRX1 \D_cache/cache_reg[1][32]  ( .D(\D_cache/n1539 ), .CK(clk), .RN(n4175), .Q(\D_cache/cache[1][32] ) );
  DFFRX1 \D_cache/cache_reg[5][32]  ( .D(\D_cache/n1535 ), .CK(clk), .RN(n4175), .Q(\D_cache/cache[5][32] ) );
  DFFRX1 \D_cache/cache_reg[1][36]  ( .D(\D_cache/n1507 ), .CK(clk), .RN(n4178), .Q(\D_cache/cache[1][36] ) );
  DFFRX1 \D_cache/cache_reg[5][36]  ( .D(\D_cache/n1503 ), .CK(clk), .RN(n4178), .Q(\D_cache/cache[5][36] ) );
  DFFRX1 \D_cache/cache_reg[1][39]  ( .D(\D_cache/n1483 ), .CK(clk), .RN(n4180), .Q(\D_cache/cache[1][39] ) );
  DFFRX1 \D_cache/cache_reg[5][39]  ( .D(\D_cache/n1479 ), .CK(clk), .RN(n4180), .Q(\D_cache/cache[5][39] ) );
  DFFRX1 \D_cache/cache_reg[1][40]  ( .D(\D_cache/n1475 ), .CK(clk), .RN(n4180), .Q(\D_cache/cache[1][40] ) );
  DFFRX1 \D_cache/cache_reg[5][40]  ( .D(\D_cache/n1471 ), .CK(clk), .RN(n4181), .Q(\D_cache/cache[5][40] ) );
  DFFRX1 \D_cache/cache_reg[1][41]  ( .D(\D_cache/n1467 ), .CK(clk), .RN(n4181), .Q(\D_cache/cache[1][41] ) );
  DFFRX1 \D_cache/cache_reg[5][41]  ( .D(\D_cache/n1463 ), .CK(clk), .RN(n4181), .Q(\D_cache/cache[5][41] ) );
  DFFRX1 \D_cache/cache_reg[1][43]  ( .D(\D_cache/n1451 ), .CK(clk), .RN(n4182), .Q(\D_cache/cache[1][43] ) );
  DFFRX1 \D_cache/cache_reg[5][43]  ( .D(\D_cache/n1447 ), .CK(clk), .RN(n4183), .Q(\D_cache/cache[5][43] ) );
  DFFRX1 \D_cache/cache_reg[1][44]  ( .D(\D_cache/n1443 ), .CK(clk), .RN(n4183), .Q(\D_cache/cache[1][44] ) );
  DFFRX1 \D_cache/cache_reg[5][44]  ( .D(\D_cache/n1439 ), .CK(clk), .RN(n4183), .Q(\D_cache/cache[5][44] ) );
  DFFRX1 \D_cache/cache_reg[1][45]  ( .D(\D_cache/n1435 ), .CK(clk), .RN(n4184), .Q(\D_cache/cache[1][45] ) );
  DFFRX1 \D_cache/cache_reg[5][45]  ( .D(\D_cache/n1431 ), .CK(clk), .RN(n4184), .Q(\D_cache/cache[5][45] ) );
  DFFRX1 \D_cache/cache_reg[1][53]  ( .D(\D_cache/n1371 ), .CK(clk), .RN(n4189), .Q(\D_cache/cache[1][53] ) );
  DFFRX1 \D_cache/cache_reg[5][53]  ( .D(\D_cache/n1367 ), .CK(clk), .RN(n4189), .Q(\D_cache/cache[5][53] ) );
  DFFRX1 \D_cache/cache_reg[1][54]  ( .D(\D_cache/n1363 ), .CK(clk), .RN(n4190), .Q(\D_cache/cache[1][54] ) );
  DFFRX1 \D_cache/cache_reg[5][54]  ( .D(\D_cache/n1359 ), .CK(clk), .RN(n4190), .Q(\D_cache/cache[5][54] ) );
  DFFRX1 \D_cache/cache_reg[1][60]  ( .D(\D_cache/n1315 ), .CK(clk), .RN(n4194), .Q(\D_cache/cache[1][60] ) );
  DFFRX1 \D_cache/cache_reg[5][60]  ( .D(\D_cache/n1311 ), .CK(clk), .RN(n4194), .Q(\D_cache/cache[5][60] ) );
  DFFRX1 \D_cache/cache_reg[5][64]  ( .D(\D_cache/n1279 ), .CK(clk), .RN(n4197), .Q(\D_cache/cache[5][64] ) );
  DFFRX1 \D_cache/cache_reg[5][66]  ( .D(\D_cache/n1263 ), .CK(clk), .RN(n4198), .Q(\D_cache/cache[5][66] ) );
  DFFRX1 \D_cache/cache_reg[1][69]  ( .D(\D_cache/n1243 ), .CK(clk), .RN(n4200), .Q(\D_cache/cache[1][69] ) );
  DFFRX1 \D_cache/cache_reg[5][69]  ( .D(\D_cache/n1239 ), .CK(clk), .RN(n4200), .Q(\D_cache/cache[5][69] ) );
  DFFRX1 \D_cache/cache_reg[1][70]  ( .D(\D_cache/n1235 ), .CK(clk), .RN(n4200), .Q(\D_cache/cache[1][70] ) );
  DFFRX1 \D_cache/cache_reg[5][70]  ( .D(\D_cache/n1231 ), .CK(clk), .RN(n4201), .Q(\D_cache/cache[5][70] ) );
  DFFRX1 \D_cache/cache_reg[1][71]  ( .D(\D_cache/n1227 ), .CK(clk), .RN(n4201), .Q(\D_cache/cache[1][71] ) );
  DFFRX1 \D_cache/cache_reg[5][71]  ( .D(\D_cache/n1223 ), .CK(clk), .RN(n4201), .Q(\D_cache/cache[5][71] ) );
  DFFRX1 \D_cache/cache_reg[1][72]  ( .D(\D_cache/n1219 ), .CK(clk), .RN(n4202), .Q(\D_cache/cache[1][72] ) );
  DFFRX1 \D_cache/cache_reg[5][72]  ( .D(\D_cache/n1215 ), .CK(clk), .RN(n4202), .Q(\D_cache/cache[5][72] ) );
  DFFRX1 \D_cache/cache_reg[1][73]  ( .D(\D_cache/n1211 ), .CK(clk), .RN(n4202), .Q(\D_cache/cache[1][73] ) );
  DFFRX1 \D_cache/cache_reg[5][73]  ( .D(\D_cache/n1207 ), .CK(clk), .RN(n4203), .Q(\D_cache/cache[5][73] ) );
  DFFRX1 \D_cache/cache_reg[1][74]  ( .D(\D_cache/n1203 ), .CK(clk), .RN(n4203), .Q(\D_cache/cache[1][74] ) );
  DFFRX1 \D_cache/cache_reg[5][74]  ( .D(\D_cache/n1199 ), .CK(clk), .RN(n4203), .Q(\D_cache/cache[5][74] ) );
  DFFRX1 \D_cache/cache_reg[1][75]  ( .D(\D_cache/n1195 ), .CK(clk), .RN(n4204), .Q(\D_cache/cache[1][75] ) );
  DFFRX1 \D_cache/cache_reg[5][75]  ( .D(\D_cache/n1191 ), .CK(clk), .RN(n4204), .Q(\D_cache/cache[5][75] ) );
  DFFRX1 \D_cache/cache_reg[1][76]  ( .D(\D_cache/n1187 ), .CK(clk), .RN(n4204), .Q(\D_cache/cache[1][76] ) );
  DFFRX1 \D_cache/cache_reg[5][76]  ( .D(\D_cache/n1183 ), .CK(clk), .RN(n4205), .Q(\D_cache/cache[5][76] ) );
  DFFRX1 \D_cache/cache_reg[1][77]  ( .D(\D_cache/n1179 ), .CK(clk), .RN(n4205), .Q(\D_cache/cache[1][77] ) );
  DFFRX1 \D_cache/cache_reg[5][77]  ( .D(\D_cache/n1175 ), .CK(clk), .RN(n4205), .Q(\D_cache/cache[5][77] ) );
  DFFRX1 \D_cache/cache_reg[1][96]  ( .D(\D_cache/n1027 ), .CK(clk), .RN(n4218), .Q(\D_cache/cache[1][96] ) );
  DFFRX1 \D_cache/cache_reg[5][96]  ( .D(\D_cache/n1023 ), .CK(clk), .RN(n4218), .Q(\D_cache/cache[5][96] ) );
  DFFRX1 \D_cache/cache_reg[1][98]  ( .D(\D_cache/n1011 ), .CK(clk), .RN(n4219), .Q(\D_cache/cache[1][98] ) );
  DFFRX1 \D_cache/cache_reg[5][98]  ( .D(\D_cache/n1007 ), .CK(clk), .RN(n4219), .Q(\D_cache/cache[5][98] ) );
  DFFRX1 \D_cache/cache_reg[1][99]  ( .D(\D_cache/n1003 ), .CK(clk), .RN(n4220), .Q(\D_cache/cache[1][99] ) );
  DFFRX1 \D_cache/cache_reg[5][99]  ( .D(\D_cache/n999 ), .CK(clk), .RN(n4220), 
        .Q(\D_cache/cache[5][99] ) );
  DFFRX1 \D_cache/cache_reg[1][100]  ( .D(\D_cache/n995 ), .CK(clk), .RN(n4220), .Q(\D_cache/cache[1][100] ) );
  DFFRX1 \D_cache/cache_reg[5][100]  ( .D(\D_cache/n991 ), .CK(clk), .RN(n4221), .Q(\D_cache/cache[5][100] ) );
  DFFRX1 \D_cache/cache_reg[1][101]  ( .D(\D_cache/n987 ), .CK(clk), .RN(n4221), .Q(\D_cache/cache[1][101] ) );
  DFFRX1 \D_cache/cache_reg[5][101]  ( .D(\D_cache/n983 ), .CK(clk), .RN(n4221), .Q(\D_cache/cache[5][101] ) );
  DFFRX1 \D_cache/cache_reg[1][102]  ( .D(\D_cache/n979 ), .CK(clk), .RN(n4222), .Q(\D_cache/cache[1][102] ) );
  DFFRX1 \D_cache/cache_reg[5][102]  ( .D(\D_cache/n975 ), .CK(clk), .RN(n4222), .Q(\D_cache/cache[5][102] ) );
  DFFRX1 \D_cache/cache_reg[1][103]  ( .D(\D_cache/n971 ), .CK(clk), .RN(n4222), .Q(\D_cache/cache[1][103] ) );
  DFFRX1 \D_cache/cache_reg[5][103]  ( .D(\D_cache/n967 ), .CK(clk), .RN(n4223), .Q(\D_cache/cache[5][103] ) );
  DFFRX1 \D_cache/cache_reg[1][104]  ( .D(\D_cache/n963 ), .CK(clk), .RN(n4223), .Q(\D_cache/cache[1][104] ) );
  DFFRX1 \D_cache/cache_reg[5][104]  ( .D(\D_cache/n959 ), .CK(clk), .RN(n4223), .Q(\D_cache/cache[5][104] ) );
  DFFRX1 \D_cache/cache_reg[1][105]  ( .D(\D_cache/n955 ), .CK(clk), .RN(n4224), .Q(\D_cache/cache[1][105] ) );
  DFFRX1 \D_cache/cache_reg[5][105]  ( .D(\D_cache/n951 ), .CK(clk), .RN(n4224), .Q(\D_cache/cache[5][105] ) );
  DFFRX1 \D_cache/cache_reg[1][106]  ( .D(\D_cache/n947 ), .CK(clk), .RN(n4224), .Q(\D_cache/cache[1][106] ) );
  DFFRX1 \D_cache/cache_reg[5][106]  ( .D(\D_cache/n943 ), .CK(clk), .RN(n4225), .Q(\D_cache/cache[5][106] ) );
  DFFRX1 \D_cache/cache_reg[1][107]  ( .D(\D_cache/n939 ), .CK(clk), .RN(n4225), .Q(\D_cache/cache[1][107] ) );
  DFFRX1 \D_cache/cache_reg[5][107]  ( .D(\D_cache/n935 ), .CK(clk), .RN(n4225), .Q(\D_cache/cache[5][107] ) );
  DFFRX1 \D_cache/cache_reg[1][108]  ( .D(\D_cache/n931 ), .CK(clk), .RN(n4226), .Q(\D_cache/cache[1][108] ) );
  DFFRX1 \D_cache/cache_reg[5][108]  ( .D(\D_cache/n927 ), .CK(clk), .RN(n4226), .Q(\D_cache/cache[5][108] ) );
  DFFRX1 \D_cache/cache_reg[1][109]  ( .D(\D_cache/n923 ), .CK(clk), .RN(n4226), .Q(\D_cache/cache[1][109] ) );
  DFFRX1 \D_cache/cache_reg[5][109]  ( .D(\D_cache/n919 ), .CK(clk), .RN(n4227), .Q(\D_cache/cache[5][109] ) );
  DFFRX1 \D_cache/cache_reg[1][110]  ( .D(\D_cache/n915 ), .CK(clk), .RN(n4227), .Q(\D_cache/cache[1][110] ) );
  DFFRX1 \D_cache/cache_reg[5][110]  ( .D(\D_cache/n911 ), .CK(clk), .RN(n4227), .Q(\D_cache/cache[5][110] ) );
  DFFRX1 \D_cache/cache_reg[1][118]  ( .D(\D_cache/n851 ), .CK(clk), .RN(n4232), .Q(\D_cache/cache[1][118] ) );
  DFFRX1 \D_cache/cache_reg[5][118]  ( .D(\D_cache/n847 ), .CK(clk), .RN(n4233), .Q(\D_cache/cache[5][118] ) );
  DFFRX1 \D_cache/cache_reg[1][135]  ( .D(\D_cache/n715 ), .CK(clk), .RN(n4244), .Q(\D_cache/cache[1][135] ) );
  DFFRX1 \D_cache/cache_reg[5][135]  ( .D(\D_cache/n711 ), .CK(clk), .RN(n4244), .Q(\D_cache/cache[5][135] ) );
  DFFRX1 \D_cache/cache_reg[1][136]  ( .D(\D_cache/n707 ), .CK(clk), .RN(n4244), .Q(\D_cache/cache[1][136] ) );
  DFFRX1 \D_cache/cache_reg[5][136]  ( .D(\D_cache/n703 ), .CK(clk), .RN(n4245), .Q(\D_cache/cache[5][136] ) );
  DFFRX1 \D_cache/cache_reg[1][137]  ( .D(\D_cache/n699 ), .CK(clk), .RN(n4245), .Q(\D_cache/cache[1][137] ) );
  DFFRX1 \D_cache/cache_reg[5][137]  ( .D(\D_cache/n695 ), .CK(clk), .RN(n4245), .Q(\D_cache/cache[5][137] ) );
  DFFRX1 \D_cache/cache_reg[1][153]  ( .D(\D_cache/n571 ), .CK(clk), .RN(n4256), .Q(\D_cache/cache[1][153] ) );
  DFFRX1 \D_cache/cache_reg[5][153]  ( .D(\D_cache/n567 ), .CK(clk), .RN(n4256), .Q(\D_cache/cache[5][153] ) );
  DFFRX1 \D_cache/cache_reg[1][154]  ( .D(\D_cache/n563 ), .CK(clk), .RN(n4256), .Q(\D_cache/cache[1][154] ) );
  DFFRX1 \D_cache/cache_reg[5][154]  ( .D(\D_cache/n559 ), .CK(clk), .RN(n4257), .Q(\D_cache/cache[5][154] ) );
  DFFRX1 \D_cache/cache_reg[0][0]  ( .D(\D_cache/n1795 ), .CK(clk), .RN(n4154), 
        .Q(\D_cache/cache[0][0] ) );
  DFFRX1 \D_cache/cache_reg[4][0]  ( .D(\D_cache/n1791 ), .CK(clk), .RN(n4154), 
        .Q(\D_cache/cache[4][0] ) );
  DFFRX1 \D_cache/cache_reg[0][1]  ( .D(\D_cache/n1788 ), .CK(clk), .RN(n4154), 
        .Q(\D_cache/cache[0][1] ) );
  DFFRX1 \D_cache/cache_reg[4][1]  ( .D(\D_cache/n1784 ), .CK(clk), .RN(n4155), 
        .Q(\D_cache/cache[4][1] ) );
  DFFRX1 \D_cache/cache_reg[0][2]  ( .D(\D_cache/n1780 ), .CK(clk), .RN(n4155), 
        .Q(\D_cache/cache[0][2] ) );
  DFFRX1 \D_cache/cache_reg[4][2]  ( .D(\D_cache/n1776 ), .CK(clk), .RN(n4155), 
        .Q(\D_cache/cache[4][2] ) );
  DFFRX1 \D_cache/cache_reg[0][3]  ( .D(\D_cache/n1772 ), .CK(clk), .RN(n4156), 
        .Q(\D_cache/cache[0][3] ) );
  DFFRX1 \D_cache/cache_reg[4][3]  ( .D(\D_cache/n1768 ), .CK(clk), .RN(n4156), 
        .Q(\D_cache/cache[4][3] ) );
  DFFRX1 \D_cache/cache_reg[0][4]  ( .D(\D_cache/n1764 ), .CK(clk), .RN(n4156), 
        .Q(\D_cache/cache[0][4] ) );
  DFFRX1 \D_cache/cache_reg[4][4]  ( .D(\D_cache/n1760 ), .CK(clk), .RN(n4157), 
        .Q(\D_cache/cache[4][4] ) );
  DFFRX1 \D_cache/cache_reg[0][5]  ( .D(\D_cache/n1756 ), .CK(clk), .RN(n4157), 
        .Q(\D_cache/cache[0][5] ) );
  DFFRX1 \D_cache/cache_reg[4][5]  ( .D(\D_cache/n1752 ), .CK(clk), .RN(n4157), 
        .Q(\D_cache/cache[4][5] ) );
  DFFRX1 \D_cache/cache_reg[0][6]  ( .D(\D_cache/n1748 ), .CK(clk), .RN(n4158), 
        .Q(\D_cache/cache[0][6] ) );
  DFFRX1 \D_cache/cache_reg[4][6]  ( .D(\D_cache/n1744 ), .CK(clk), .RN(n4158), 
        .Q(\D_cache/cache[4][6] ) );
  DFFRX1 \D_cache/cache_reg[0][7]  ( .D(\D_cache/n1740 ), .CK(clk), .RN(n4158), 
        .Q(\D_cache/cache[0][7] ) );
  DFFRX1 \D_cache/cache_reg[4][7]  ( .D(\D_cache/n1736 ), .CK(clk), .RN(n4159), 
        .Q(\D_cache/cache[4][7] ) );
  DFFRX1 \D_cache/cache_reg[0][8]  ( .D(\D_cache/n1732 ), .CK(clk), .RN(n4159), 
        .Q(\D_cache/cache[0][8] ) );
  DFFRX1 \D_cache/cache_reg[4][8]  ( .D(\D_cache/n1728 ), .CK(clk), .RN(n4159), 
        .Q(\D_cache/cache[4][8] ) );
  DFFRX1 \D_cache/cache_reg[0][9]  ( .D(\D_cache/n1724 ), .CK(clk), .RN(n4160), 
        .Q(\D_cache/cache[0][9] ) );
  DFFRX1 \D_cache/cache_reg[4][9]  ( .D(\D_cache/n1720 ), .CK(clk), .RN(n4160), 
        .Q(\D_cache/cache[4][9] ) );
  DFFRX1 \D_cache/cache_reg[0][10]  ( .D(\D_cache/n1716 ), .CK(clk), .RN(n4160), .Q(\D_cache/cache[0][10] ) );
  DFFRX1 \D_cache/cache_reg[4][10]  ( .D(\D_cache/n1712 ), .CK(clk), .RN(n4161), .Q(\D_cache/cache[4][10] ) );
  DFFRX1 \D_cache/cache_reg[0][11]  ( .D(\D_cache/n1708 ), .CK(clk), .RN(n4161), .Q(\D_cache/cache[0][11] ) );
  DFFRX1 \D_cache/cache_reg[4][11]  ( .D(\D_cache/n1704 ), .CK(clk), .RN(n4161), .Q(\D_cache/cache[4][11] ) );
  DFFRX1 \D_cache/cache_reg[0][12]  ( .D(\D_cache/n1700 ), .CK(clk), .RN(n4162), .Q(\D_cache/cache[0][12] ) );
  DFFRX1 \D_cache/cache_reg[4][12]  ( .D(\D_cache/n1696 ), .CK(clk), .RN(n4162), .Q(\D_cache/cache[4][12] ) );
  DFFRX1 \D_cache/cache_reg[0][13]  ( .D(\D_cache/n1692 ), .CK(clk), .RN(n4162), .Q(\D_cache/cache[0][13] ) );
  DFFRX1 \D_cache/cache_reg[4][13]  ( .D(\D_cache/n1688 ), .CK(clk), .RN(n4163), .Q(\D_cache/cache[4][13] ) );
  DFFRX1 \D_cache/cache_reg[0][14]  ( .D(\D_cache/n1684 ), .CK(clk), .RN(n4163), .Q(\D_cache/cache[0][14] ) );
  DFFRX1 \D_cache/cache_reg[4][14]  ( .D(\D_cache/n1680 ), .CK(clk), .RN(n4163), .Q(\D_cache/cache[4][14] ) );
  DFFRX1 \D_cache/cache_reg[0][15]  ( .D(\D_cache/n1676 ), .CK(clk), .RN(n4164), .Q(\D_cache/cache[0][15] ) );
  DFFRX1 \D_cache/cache_reg[4][15]  ( .D(\D_cache/n1672 ), .CK(clk), .RN(n4164), .Q(\D_cache/cache[4][15] ) );
  DFFRX1 \D_cache/cache_reg[0][17]  ( .D(\D_cache/n1660 ), .CK(clk), .RN(n4165), .Q(\D_cache/cache[0][17] ) );
  DFFRX1 \D_cache/cache_reg[4][17]  ( .D(\D_cache/n1656 ), .CK(clk), .RN(n4165), .Q(\D_cache/cache[4][17] ) );
  DFFRX1 \D_cache/cache_reg[0][18]  ( .D(\D_cache/n1652 ), .CK(clk), .RN(n4166), .Q(\D_cache/cache[0][18] ) );
  DFFRX1 \D_cache/cache_reg[4][18]  ( .D(\D_cache/n1648 ), .CK(clk), .RN(n4166), .Q(\D_cache/cache[4][18] ) );
  DFFRX1 \D_cache/cache_reg[0][19]  ( .D(\D_cache/n1644 ), .CK(clk), .RN(n4166), .Q(\D_cache/cache[0][19] ) );
  DFFRX1 \D_cache/cache_reg[4][19]  ( .D(\D_cache/n1640 ), .CK(clk), .RN(n4167), .Q(\D_cache/cache[4][19] ) );
  DFFRX1 \D_cache/cache_reg[0][20]  ( .D(\D_cache/n1636 ), .CK(clk), .RN(n4167), .Q(\D_cache/cache[0][20] ) );
  DFFRX1 \D_cache/cache_reg[4][20]  ( .D(\D_cache/n1632 ), .CK(clk), .RN(n4167), .Q(\D_cache/cache[4][20] ) );
  DFFRX1 \D_cache/cache_reg[0][21]  ( .D(\D_cache/n1628 ), .CK(clk), .RN(n4168), .Q(\D_cache/cache[0][21] ) );
  DFFRX1 \D_cache/cache_reg[4][21]  ( .D(\D_cache/n1624 ), .CK(clk), .RN(n4168), .Q(\D_cache/cache[4][21] ) );
  DFFRX1 \D_cache/cache_reg[0][22]  ( .D(\D_cache/n1620 ), .CK(clk), .RN(n4168), .Q(\D_cache/cache[0][22] ) );
  DFFRX1 \D_cache/cache_reg[4][22]  ( .D(\D_cache/n1616 ), .CK(clk), .RN(n4169), .Q(\D_cache/cache[4][22] ) );
  DFFRX1 \D_cache/cache_reg[0][23]  ( .D(\D_cache/n1612 ), .CK(clk), .RN(n4169), .Q(\D_cache/cache[0][23] ) );
  DFFRX1 \D_cache/cache_reg[4][23]  ( .D(\D_cache/n1608 ), .CK(clk), .RN(n4169), .Q(\D_cache/cache[4][23] ) );
  DFFRX1 \D_cache/cache_reg[0][24]  ( .D(\D_cache/n1604 ), .CK(clk), .RN(n4170), .Q(\D_cache/cache[0][24] ) );
  DFFRX1 \D_cache/cache_reg[4][24]  ( .D(\D_cache/n1600 ), .CK(clk), .RN(n4170), .Q(\D_cache/cache[4][24] ) );
  DFFRX1 \D_cache/cache_reg[0][25]  ( .D(\D_cache/n1596 ), .CK(clk), .RN(n4170), .Q(\D_cache/cache[0][25] ) );
  DFFRX1 \D_cache/cache_reg[4][25]  ( .D(\D_cache/n1592 ), .CK(clk), .RN(n4171), .Q(\D_cache/cache[4][25] ) );
  DFFRX1 \D_cache/cache_reg[0][26]  ( .D(\D_cache/n1588 ), .CK(clk), .RN(n4171), .Q(\D_cache/cache[0][26] ) );
  DFFRX1 \D_cache/cache_reg[4][26]  ( .D(\D_cache/n1584 ), .CK(clk), .RN(n4171), .Q(\D_cache/cache[4][26] ) );
  DFFRX1 \D_cache/cache_reg[0][27]  ( .D(\D_cache/n1580 ), .CK(clk), .RN(n4172), .Q(\D_cache/cache[0][27] ) );
  DFFRX1 \D_cache/cache_reg[4][27]  ( .D(\D_cache/n1576 ), .CK(clk), .RN(n4172), .Q(\D_cache/cache[4][27] ) );
  DFFRX1 \D_cache/cache_reg[0][28]  ( .D(\D_cache/n1572 ), .CK(clk), .RN(n4172), .Q(\D_cache/cache[0][28] ) );
  DFFRX1 \D_cache/cache_reg[4][28]  ( .D(\D_cache/n1568 ), .CK(clk), .RN(n4173), .Q(\D_cache/cache[4][28] ) );
  DFFRX1 \D_cache/cache_reg[0][31]  ( .D(\D_cache/n1548 ), .CK(clk), .RN(n4174), .Q(\D_cache/cache[0][31] ) );
  DFFRX1 \D_cache/cache_reg[4][31]  ( .D(\D_cache/n1544 ), .CK(clk), .RN(n4175), .Q(\D_cache/cache[4][31] ) );
  DFFRX1 \D_cache/cache_reg[0][32]  ( .D(\D_cache/n1540 ), .CK(clk), .RN(n4175), .Q(\D_cache/cache[0][32] ) );
  DFFRX1 \D_cache/cache_reg[4][32]  ( .D(\D_cache/n1536 ), .CK(clk), .RN(n4175), .Q(\D_cache/cache[4][32] ) );
  DFFRX1 \D_cache/cache_reg[0][36]  ( .D(\D_cache/n1508 ), .CK(clk), .RN(n4178), .Q(\D_cache/cache[0][36] ) );
  DFFRX1 \D_cache/cache_reg[4][36]  ( .D(\D_cache/n1504 ), .CK(clk), .RN(n4178), .Q(\D_cache/cache[4][36] ) );
  DFFRX1 \D_cache/cache_reg[0][39]  ( .D(\D_cache/n1484 ), .CK(clk), .RN(n4180), .Q(\D_cache/cache[0][39] ) );
  DFFRX1 \D_cache/cache_reg[4][39]  ( .D(\D_cache/n1480 ), .CK(clk), .RN(n4180), .Q(\D_cache/cache[4][39] ) );
  DFFRX1 \D_cache/cache_reg[0][40]  ( .D(\D_cache/n1476 ), .CK(clk), .RN(n4180), .Q(\D_cache/cache[0][40] ) );
  DFFRX1 \D_cache/cache_reg[4][40]  ( .D(\D_cache/n1472 ), .CK(clk), .RN(n4181), .Q(\D_cache/cache[4][40] ) );
  DFFRX1 \D_cache/cache_reg[0][41]  ( .D(\D_cache/n1468 ), .CK(clk), .RN(n4181), .Q(\D_cache/cache[0][41] ) );
  DFFRX1 \D_cache/cache_reg[4][41]  ( .D(\D_cache/n1464 ), .CK(clk), .RN(n4181), .Q(\D_cache/cache[4][41] ) );
  DFFRX1 \D_cache/cache_reg[0][43]  ( .D(\D_cache/n1452 ), .CK(clk), .RN(n4182), .Q(\D_cache/cache[0][43] ) );
  DFFRX1 \D_cache/cache_reg[4][43]  ( .D(\D_cache/n1448 ), .CK(clk), .RN(n4183), .Q(\D_cache/cache[4][43] ) );
  DFFRX1 \D_cache/cache_reg[0][44]  ( .D(\D_cache/n1444 ), .CK(clk), .RN(n4183), .Q(\D_cache/cache[0][44] ) );
  DFFRX1 \D_cache/cache_reg[4][44]  ( .D(\D_cache/n1440 ), .CK(clk), .RN(n4183), .Q(\D_cache/cache[4][44] ) );
  DFFRX1 \D_cache/cache_reg[0][45]  ( .D(\D_cache/n1436 ), .CK(clk), .RN(n4184), .Q(\D_cache/cache[0][45] ) );
  DFFRX1 \D_cache/cache_reg[4][45]  ( .D(\D_cache/n1432 ), .CK(clk), .RN(n4184), .Q(\D_cache/cache[4][45] ) );
  DFFRX1 \D_cache/cache_reg[0][53]  ( .D(\D_cache/n1372 ), .CK(clk), .RN(n4189), .Q(\D_cache/cache[0][53] ) );
  DFFRX1 \D_cache/cache_reg[4][53]  ( .D(\D_cache/n1368 ), .CK(clk), .RN(n4189), .Q(\D_cache/cache[4][53] ) );
  DFFRX1 \D_cache/cache_reg[0][54]  ( .D(\D_cache/n1364 ), .CK(clk), .RN(n4190), .Q(\D_cache/cache[0][54] ) );
  DFFRX1 \D_cache/cache_reg[4][54]  ( .D(\D_cache/n1360 ), .CK(clk), .RN(n4190), .Q(\D_cache/cache[4][54] ) );
  DFFRX1 \D_cache/cache_reg[0][60]  ( .D(\D_cache/n1316 ), .CK(clk), .RN(n4194), .Q(\D_cache/cache[0][60] ) );
  DFFRX1 \D_cache/cache_reg[4][60]  ( .D(\D_cache/n1312 ), .CK(clk), .RN(n4194), .Q(\D_cache/cache[4][60] ) );
  DFFRX1 \D_cache/cache_reg[4][64]  ( .D(\D_cache/n1280 ), .CK(clk), .RN(n4197), .Q(\D_cache/cache[4][64] ) );
  DFFRX1 \D_cache/cache_reg[0][66]  ( .D(\D_cache/n1268 ), .CK(clk), .RN(n4198), .Q(\D_cache/cache[0][66] ) );
  DFFRX1 \D_cache/cache_reg[4][66]  ( .D(\D_cache/n1264 ), .CK(clk), .RN(n4198), .Q(\D_cache/cache[4][66] ) );
  DFFRX1 \D_cache/cache_reg[0][69]  ( .D(\D_cache/n1244 ), .CK(clk), .RN(n4200), .Q(\D_cache/cache[0][69] ) );
  DFFRX1 \D_cache/cache_reg[4][69]  ( .D(\D_cache/n1240 ), .CK(clk), .RN(n4200), .Q(\D_cache/cache[4][69] ) );
  DFFRX1 \D_cache/cache_reg[0][70]  ( .D(\D_cache/n1236 ), .CK(clk), .RN(n4200), .Q(\D_cache/cache[0][70] ) );
  DFFRX1 \D_cache/cache_reg[4][70]  ( .D(\D_cache/n1232 ), .CK(clk), .RN(n4201), .Q(\D_cache/cache[4][70] ) );
  DFFRX1 \D_cache/cache_reg[0][71]  ( .D(\D_cache/n1228 ), .CK(clk), .RN(n4201), .Q(\D_cache/cache[0][71] ) );
  DFFRX1 \D_cache/cache_reg[4][71]  ( .D(\D_cache/n1224 ), .CK(clk), .RN(n4201), .Q(\D_cache/cache[4][71] ) );
  DFFRX1 \D_cache/cache_reg[0][72]  ( .D(\D_cache/n1220 ), .CK(clk), .RN(n4202), .Q(\D_cache/cache[0][72] ) );
  DFFRX1 \D_cache/cache_reg[4][72]  ( .D(\D_cache/n1216 ), .CK(clk), .RN(n4202), .Q(\D_cache/cache[4][72] ) );
  DFFRX1 \D_cache/cache_reg[0][73]  ( .D(\D_cache/n1212 ), .CK(clk), .RN(n4202), .Q(\D_cache/cache[0][73] ) );
  DFFRX1 \D_cache/cache_reg[4][73]  ( .D(\D_cache/n1208 ), .CK(clk), .RN(n4203), .Q(\D_cache/cache[4][73] ) );
  DFFRX1 \D_cache/cache_reg[0][74]  ( .D(\D_cache/n1204 ), .CK(clk), .RN(n4203), .Q(\D_cache/cache[0][74] ) );
  DFFRX1 \D_cache/cache_reg[4][74]  ( .D(\D_cache/n1200 ), .CK(clk), .RN(n4203), .Q(\D_cache/cache[4][74] ) );
  DFFRX1 \D_cache/cache_reg[0][75]  ( .D(\D_cache/n1196 ), .CK(clk), .RN(n4204), .Q(\D_cache/cache[0][75] ) );
  DFFRX1 \D_cache/cache_reg[4][75]  ( .D(\D_cache/n1192 ), .CK(clk), .RN(n4204), .Q(\D_cache/cache[4][75] ) );
  DFFRX1 \D_cache/cache_reg[0][76]  ( .D(\D_cache/n1188 ), .CK(clk), .RN(n4204), .Q(\D_cache/cache[0][76] ) );
  DFFRX1 \D_cache/cache_reg[4][76]  ( .D(\D_cache/n1184 ), .CK(clk), .RN(n4205), .Q(\D_cache/cache[4][76] ) );
  DFFRX1 \D_cache/cache_reg[0][77]  ( .D(\D_cache/n1180 ), .CK(clk), .RN(n4205), .Q(\D_cache/cache[0][77] ) );
  DFFRX1 \D_cache/cache_reg[4][77]  ( .D(\D_cache/n1176 ), .CK(clk), .RN(n4205), .Q(\D_cache/cache[4][77] ) );
  DFFRX1 \D_cache/cache_reg[0][96]  ( .D(\D_cache/n1028 ), .CK(clk), .RN(n4218), .Q(\D_cache/cache[0][96] ) );
  DFFRX1 \D_cache/cache_reg[4][96]  ( .D(\D_cache/n1024 ), .CK(clk), .RN(n4218), .Q(\D_cache/cache[4][96] ) );
  DFFRX1 \D_cache/cache_reg[0][98]  ( .D(\D_cache/n1012 ), .CK(clk), .RN(n4219), .Q(\D_cache/cache[0][98] ) );
  DFFRX1 \D_cache/cache_reg[4][98]  ( .D(\D_cache/n1008 ), .CK(clk), .RN(n4219), .Q(\D_cache/cache[4][98] ) );
  DFFRX1 \D_cache/cache_reg[0][99]  ( .D(\D_cache/n1004 ), .CK(clk), .RN(n4220), .Q(\D_cache/cache[0][99] ) );
  DFFRX1 \D_cache/cache_reg[4][99]  ( .D(\D_cache/n1000 ), .CK(clk), .RN(n4220), .Q(\D_cache/cache[4][99] ) );
  DFFRX1 \D_cache/cache_reg[0][100]  ( .D(\D_cache/n996 ), .CK(clk), .RN(n4220), .Q(\D_cache/cache[0][100] ) );
  DFFRX1 \D_cache/cache_reg[4][100]  ( .D(\D_cache/n992 ), .CK(clk), .RN(n4221), .Q(\D_cache/cache[4][100] ) );
  DFFRX1 \D_cache/cache_reg[0][101]  ( .D(\D_cache/n988 ), .CK(clk), .RN(n4221), .Q(\D_cache/cache[0][101] ) );
  DFFRX1 \D_cache/cache_reg[4][101]  ( .D(\D_cache/n984 ), .CK(clk), .RN(n4221), .Q(\D_cache/cache[4][101] ) );
  DFFRX1 \D_cache/cache_reg[0][102]  ( .D(\D_cache/n980 ), .CK(clk), .RN(n4222), .Q(\D_cache/cache[0][102] ) );
  DFFRX1 \D_cache/cache_reg[4][102]  ( .D(\D_cache/n976 ), .CK(clk), .RN(n4222), .Q(\D_cache/cache[4][102] ) );
  DFFRX1 \D_cache/cache_reg[0][103]  ( .D(\D_cache/n972 ), .CK(clk), .RN(n4222), .Q(\D_cache/cache[0][103] ) );
  DFFRX1 \D_cache/cache_reg[4][103]  ( .D(\D_cache/n968 ), .CK(clk), .RN(n4223), .Q(\D_cache/cache[4][103] ) );
  DFFRX1 \D_cache/cache_reg[0][104]  ( .D(\D_cache/n964 ), .CK(clk), .RN(n4223), .Q(\D_cache/cache[0][104] ) );
  DFFRX1 \D_cache/cache_reg[4][104]  ( .D(\D_cache/n960 ), .CK(clk), .RN(n4223), .Q(\D_cache/cache[4][104] ) );
  DFFRX1 \D_cache/cache_reg[0][105]  ( .D(\D_cache/n956 ), .CK(clk), .RN(n4224), .Q(\D_cache/cache[0][105] ) );
  DFFRX1 \D_cache/cache_reg[4][105]  ( .D(\D_cache/n952 ), .CK(clk), .RN(n4224), .Q(\D_cache/cache[4][105] ) );
  DFFRX1 \D_cache/cache_reg[0][106]  ( .D(\D_cache/n948 ), .CK(clk), .RN(n4224), .Q(\D_cache/cache[0][106] ) );
  DFFRX1 \D_cache/cache_reg[4][106]  ( .D(\D_cache/n944 ), .CK(clk), .RN(n4225), .Q(\D_cache/cache[4][106] ) );
  DFFRX1 \D_cache/cache_reg[0][107]  ( .D(\D_cache/n940 ), .CK(clk), .RN(n4225), .Q(\D_cache/cache[0][107] ) );
  DFFRX1 \D_cache/cache_reg[4][107]  ( .D(\D_cache/n936 ), .CK(clk), .RN(n4225), .Q(\D_cache/cache[4][107] ) );
  DFFRX1 \D_cache/cache_reg[0][108]  ( .D(\D_cache/n932 ), .CK(clk), .RN(n4226), .Q(\D_cache/cache[0][108] ) );
  DFFRX1 \D_cache/cache_reg[4][108]  ( .D(\D_cache/n928 ), .CK(clk), .RN(n4226), .Q(\D_cache/cache[4][108] ) );
  DFFRX1 \D_cache/cache_reg[0][109]  ( .D(\D_cache/n924 ), .CK(clk), .RN(n4226), .Q(\D_cache/cache[0][109] ) );
  DFFRX1 \D_cache/cache_reg[4][109]  ( .D(\D_cache/n920 ), .CK(clk), .RN(n4227), .Q(\D_cache/cache[4][109] ) );
  DFFRX1 \D_cache/cache_reg[0][110]  ( .D(\D_cache/n916 ), .CK(clk), .RN(n4227), .Q(\D_cache/cache[0][110] ) );
  DFFRX1 \D_cache/cache_reg[4][110]  ( .D(\D_cache/n912 ), .CK(clk), .RN(n4227), .Q(\D_cache/cache[4][110] ) );
  DFFRX1 \D_cache/cache_reg[0][118]  ( .D(\D_cache/n852 ), .CK(clk), .RN(n4232), .Q(\D_cache/cache[0][118] ) );
  DFFRX1 \D_cache/cache_reg[4][118]  ( .D(\D_cache/n848 ), .CK(clk), .RN(n4233), .Q(\D_cache/cache[4][118] ) );
  DFFRX1 \D_cache/cache_reg[0][135]  ( .D(\D_cache/n716 ), .CK(clk), .RN(n4243), .Q(\D_cache/cache[0][135] ) );
  DFFRX1 \D_cache/cache_reg[4][135]  ( .D(\D_cache/n712 ), .CK(clk), .RN(n4244), .Q(\D_cache/cache[4][135] ) );
  DFFRX1 \D_cache/cache_reg[0][136]  ( .D(\D_cache/n708 ), .CK(clk), .RN(n4244), .Q(\D_cache/cache[0][136] ) );
  DFFRX1 \D_cache/cache_reg[4][136]  ( .D(\D_cache/n704 ), .CK(clk), .RN(n4244), .Q(\D_cache/cache[4][136] ) );
  DFFRX1 \D_cache/cache_reg[0][137]  ( .D(\D_cache/n700 ), .CK(clk), .RN(n4245), .Q(\D_cache/cache[0][137] ) );
  DFFRX1 \D_cache/cache_reg[4][137]  ( .D(\D_cache/n696 ), .CK(clk), .RN(n4245), .Q(\D_cache/cache[4][137] ) );
  DFFRX1 \D_cache/cache_reg[0][153]  ( .D(\D_cache/n572 ), .CK(clk), .RN(n4255), .Q(\D_cache/cache[0][153] ) );
  DFFRX1 \D_cache/cache_reg[4][153]  ( .D(\D_cache/n568 ), .CK(clk), .RN(n4256), .Q(\D_cache/cache[4][153] ) );
  DFFRX1 \D_cache/cache_reg[0][154]  ( .D(\D_cache/n564 ), .CK(clk), .RN(n4256), .Q(\D_cache/cache[0][154] ) );
  DFFRX1 \D_cache/cache_reg[4][154]  ( .D(\D_cache/n560 ), .CK(clk), .RN(n4257), .Q(\D_cache/cache[4][154] ) );
  DFFRX1 \D_cache/cache_reg[2][0]  ( .D(\D_cache/n1793 ), .CK(clk), .RN(n4154), 
        .Q(\D_cache/cache[2][0] ) );
  DFFRX1 \D_cache/cache_reg[6][0]  ( .D(\D_cache/n1789 ), .CK(clk), .RN(n4154), 
        .Q(\D_cache/cache[6][0] ) );
  DFFRX1 \D_cache/cache_reg[2][1]  ( .D(\D_cache/n1786 ), .CK(clk), .RN(n4154), 
        .Q(\D_cache/cache[2][1] ) );
  DFFRX1 \D_cache/cache_reg[6][1]  ( .D(\D_cache/n1782 ), .CK(clk), .RN(n4155), 
        .Q(\D_cache/cache[6][1] ) );
  DFFRX1 \D_cache/cache_reg[2][2]  ( .D(\D_cache/n1778 ), .CK(clk), .RN(n4155), 
        .Q(\D_cache/cache[2][2] ) );
  DFFRX1 \D_cache/cache_reg[6][2]  ( .D(\D_cache/n1774 ), .CK(clk), .RN(n4155), 
        .Q(\D_cache/cache[6][2] ) );
  DFFRX1 \D_cache/cache_reg[2][3]  ( .D(\D_cache/n1770 ), .CK(clk), .RN(n4156), 
        .Q(\D_cache/cache[2][3] ) );
  DFFRX1 \D_cache/cache_reg[6][3]  ( .D(\D_cache/n1766 ), .CK(clk), .RN(n4156), 
        .Q(\D_cache/cache[6][3] ) );
  DFFRX1 \D_cache/cache_reg[2][4]  ( .D(\D_cache/n1762 ), .CK(clk), .RN(n4156), 
        .Q(\D_cache/cache[2][4] ) );
  DFFRX1 \D_cache/cache_reg[6][4]  ( .D(\D_cache/n1758 ), .CK(clk), .RN(n4157), 
        .Q(\D_cache/cache[6][4] ) );
  DFFRX1 \D_cache/cache_reg[2][5]  ( .D(\D_cache/n1754 ), .CK(clk), .RN(n4157), 
        .Q(\D_cache/cache[2][5] ) );
  DFFRX1 \D_cache/cache_reg[6][5]  ( .D(\D_cache/n1750 ), .CK(clk), .RN(n4157), 
        .Q(\D_cache/cache[6][5] ) );
  DFFRX1 \D_cache/cache_reg[2][6]  ( .D(\D_cache/n1746 ), .CK(clk), .RN(n4158), 
        .Q(\D_cache/cache[2][6] ) );
  DFFRX1 \D_cache/cache_reg[6][6]  ( .D(\D_cache/n1742 ), .CK(clk), .RN(n4158), 
        .Q(\D_cache/cache[6][6] ) );
  DFFRX1 \D_cache/cache_reg[2][7]  ( .D(\D_cache/n1738 ), .CK(clk), .RN(n4158), 
        .Q(\D_cache/cache[2][7] ) );
  DFFRX1 \D_cache/cache_reg[6][7]  ( .D(\D_cache/n1734 ), .CK(clk), .RN(n4159), 
        .Q(\D_cache/cache[6][7] ) );
  DFFRX1 \D_cache/cache_reg[2][8]  ( .D(\D_cache/n1730 ), .CK(clk), .RN(n4159), 
        .Q(\D_cache/cache[2][8] ) );
  DFFRX1 \D_cache/cache_reg[6][8]  ( .D(\D_cache/n1726 ), .CK(clk), .RN(n4159), 
        .Q(\D_cache/cache[6][8] ) );
  DFFRX1 \D_cache/cache_reg[2][9]  ( .D(\D_cache/n1722 ), .CK(clk), .RN(n4160), 
        .Q(\D_cache/cache[2][9] ) );
  DFFRX1 \D_cache/cache_reg[6][9]  ( .D(\D_cache/n1718 ), .CK(clk), .RN(n4160), 
        .Q(\D_cache/cache[6][9] ) );
  DFFRX1 \D_cache/cache_reg[2][10]  ( .D(\D_cache/n1714 ), .CK(clk), .RN(n4160), .Q(\D_cache/cache[2][10] ) );
  DFFRX1 \D_cache/cache_reg[6][10]  ( .D(\D_cache/n1710 ), .CK(clk), .RN(n4161), .Q(\D_cache/cache[6][10] ) );
  DFFRX1 \D_cache/cache_reg[2][11]  ( .D(\D_cache/n1706 ), .CK(clk), .RN(n4161), .Q(\D_cache/cache[2][11] ) );
  DFFRX1 \D_cache/cache_reg[6][11]  ( .D(\D_cache/n1702 ), .CK(clk), .RN(n4161), .Q(\D_cache/cache[6][11] ) );
  DFFRX1 \D_cache/cache_reg[2][12]  ( .D(\D_cache/n1698 ), .CK(clk), .RN(n4162), .Q(\D_cache/cache[2][12] ) );
  DFFRX1 \D_cache/cache_reg[6][12]  ( .D(\D_cache/n1694 ), .CK(clk), .RN(n4162), .Q(\D_cache/cache[6][12] ) );
  DFFRX1 \D_cache/cache_reg[2][13]  ( .D(\D_cache/n1690 ), .CK(clk), .RN(n4162), .Q(\D_cache/cache[2][13] ) );
  DFFRX1 \D_cache/cache_reg[6][13]  ( .D(\D_cache/n1686 ), .CK(clk), .RN(n4163), .Q(\D_cache/cache[6][13] ) );
  DFFRX1 \D_cache/cache_reg[2][14]  ( .D(\D_cache/n1682 ), .CK(clk), .RN(n4163), .Q(\D_cache/cache[2][14] ) );
  DFFRX1 \D_cache/cache_reg[6][14]  ( .D(\D_cache/n1678 ), .CK(clk), .RN(n4163), .Q(\D_cache/cache[6][14] ) );
  DFFRX1 \D_cache/cache_reg[6][15]  ( .D(\D_cache/n1670 ), .CK(clk), .RN(n4164), .Q(\D_cache/cache[6][15] ) );
  DFFRX1 \D_cache/cache_reg[2][17]  ( .D(\D_cache/n1658 ), .CK(clk), .RN(n4165), .Q(\D_cache/cache[2][17] ) );
  DFFRX1 \D_cache/cache_reg[6][17]  ( .D(\D_cache/n1654 ), .CK(clk), .RN(n4165), .Q(\D_cache/cache[6][17] ) );
  DFFRX1 \D_cache/cache_reg[2][18]  ( .D(\D_cache/n1650 ), .CK(clk), .RN(n4166), .Q(\D_cache/cache[2][18] ) );
  DFFRX1 \D_cache/cache_reg[6][18]  ( .D(\D_cache/n1646 ), .CK(clk), .RN(n4166), .Q(\D_cache/cache[6][18] ) );
  DFFRX1 \D_cache/cache_reg[2][19]  ( .D(\D_cache/n1642 ), .CK(clk), .RN(n4166), .Q(\D_cache/cache[2][19] ) );
  DFFRX1 \D_cache/cache_reg[6][19]  ( .D(\D_cache/n1638 ), .CK(clk), .RN(n4167), .Q(\D_cache/cache[6][19] ) );
  DFFRX1 \D_cache/cache_reg[2][20]  ( .D(\D_cache/n1634 ), .CK(clk), .RN(n4167), .Q(\D_cache/cache[2][20] ) );
  DFFRX1 \D_cache/cache_reg[6][20]  ( .D(\D_cache/n1630 ), .CK(clk), .RN(n4167), .Q(\D_cache/cache[6][20] ) );
  DFFRX1 \D_cache/cache_reg[2][21]  ( .D(\D_cache/n1626 ), .CK(clk), .RN(n4168), .Q(\D_cache/cache[2][21] ) );
  DFFRX1 \D_cache/cache_reg[6][21]  ( .D(\D_cache/n1622 ), .CK(clk), .RN(n4168), .Q(\D_cache/cache[6][21] ) );
  DFFRX1 \D_cache/cache_reg[2][22]  ( .D(\D_cache/n1618 ), .CK(clk), .RN(n4168), .Q(\D_cache/cache[2][22] ) );
  DFFRX1 \D_cache/cache_reg[6][22]  ( .D(\D_cache/n1614 ), .CK(clk), .RN(n4169), .Q(\D_cache/cache[6][22] ) );
  DFFRX1 \D_cache/cache_reg[2][23]  ( .D(\D_cache/n1610 ), .CK(clk), .RN(n4169), .Q(\D_cache/cache[2][23] ) );
  DFFRX1 \D_cache/cache_reg[6][23]  ( .D(\D_cache/n1606 ), .CK(clk), .RN(n4169), .Q(\D_cache/cache[6][23] ) );
  DFFRX1 \D_cache/cache_reg[2][24]  ( .D(\D_cache/n1602 ), .CK(clk), .RN(n4170), .Q(\D_cache/cache[2][24] ) );
  DFFRX1 \D_cache/cache_reg[6][24]  ( .D(\D_cache/n1598 ), .CK(clk), .RN(n4170), .Q(\D_cache/cache[6][24] ) );
  DFFRX1 \D_cache/cache_reg[2][25]  ( .D(\D_cache/n1594 ), .CK(clk), .RN(n4170), .Q(\D_cache/cache[2][25] ) );
  DFFRX1 \D_cache/cache_reg[6][25]  ( .D(\D_cache/n1590 ), .CK(clk), .RN(n4171), .Q(\D_cache/cache[6][25] ) );
  DFFRX1 \D_cache/cache_reg[2][26]  ( .D(\D_cache/n1586 ), .CK(clk), .RN(n4171), .Q(\D_cache/cache[2][26] ) );
  DFFRX1 \D_cache/cache_reg[6][26]  ( .D(\D_cache/n1582 ), .CK(clk), .RN(n4171), .Q(\D_cache/cache[6][26] ) );
  DFFRX1 \D_cache/cache_reg[2][27]  ( .D(\D_cache/n1578 ), .CK(clk), .RN(n4172), .Q(\D_cache/cache[2][27] ) );
  DFFRX1 \D_cache/cache_reg[6][27]  ( .D(\D_cache/n1574 ), .CK(clk), .RN(n4172), .Q(\D_cache/cache[6][27] ) );
  DFFRX1 \D_cache/cache_reg[2][28]  ( .D(\D_cache/n1570 ), .CK(clk), .RN(n4172), .Q(\D_cache/cache[2][28] ) );
  DFFRX1 \D_cache/cache_reg[6][28]  ( .D(\D_cache/n1566 ), .CK(clk), .RN(n4173), .Q(\D_cache/cache[6][28] ) );
  DFFRX1 \D_cache/cache_reg[2][31]  ( .D(\D_cache/n1546 ), .CK(clk), .RN(n4174), .Q(\D_cache/cache[2][31] ) );
  DFFRX1 \D_cache/cache_reg[6][31]  ( .D(\D_cache/n1542 ), .CK(clk), .RN(n4175), .Q(\D_cache/cache[6][31] ) );
  DFFRX1 \D_cache/cache_reg[2][39]  ( .D(\D_cache/n1482 ), .CK(clk), .RN(n4180), .Q(\D_cache/cache[2][39] ) );
  DFFRX1 \D_cache/cache_reg[6][39]  ( .D(\D_cache/n1478 ), .CK(clk), .RN(n4180), .Q(\D_cache/cache[6][39] ) );
  DFFRX1 \D_cache/cache_reg[2][41]  ( .D(\D_cache/n1466 ), .CK(clk), .RN(n4181), .Q(\D_cache/cache[2][41] ) );
  DFFRX1 \D_cache/cache_reg[6][41]  ( .D(\D_cache/n1462 ), .CK(clk), .RN(n4181), .Q(\D_cache/cache[6][41] ) );
  DFFRX1 \D_cache/cache_reg[2][43]  ( .D(\D_cache/n1450 ), .CK(clk), .RN(n4182), .Q(\D_cache/cache[2][43] ) );
  DFFRX1 \D_cache/cache_reg[6][43]  ( .D(\D_cache/n1446 ), .CK(clk), .RN(n4183), .Q(\D_cache/cache[6][43] ) );
  DFFRX1 \D_cache/cache_reg[2][45]  ( .D(\D_cache/n1434 ), .CK(clk), .RN(n4184), .Q(\D_cache/cache[2][45] ) );
  DFFRX1 \D_cache/cache_reg[6][45]  ( .D(\D_cache/n1430 ), .CK(clk), .RN(n4184), .Q(\D_cache/cache[6][45] ) );
  DFFRX1 \D_cache/cache_reg[2][53]  ( .D(\D_cache/n1370 ), .CK(clk), .RN(n4189), .Q(\D_cache/cache[2][53] ) );
  DFFRX1 \D_cache/cache_reg[2][54]  ( .D(\D_cache/n1362 ), .CK(clk), .RN(n4190), .Q(\D_cache/cache[2][54] ) );
  DFFRX1 \D_cache/cache_reg[6][54]  ( .D(\D_cache/n1358 ), .CK(clk), .RN(n4190), .Q(\D_cache/cache[6][54] ) );
  DFFRX1 \D_cache/cache_reg[2][69]  ( .D(\D_cache/n1242 ), .CK(clk), .RN(n4200), .Q(\D_cache/cache[2][69] ) );
  DFFRX1 \D_cache/cache_reg[6][69]  ( .D(\D_cache/n1238 ), .CK(clk), .RN(n4200), .Q(\D_cache/cache[6][69] ) );
  DFFRX1 \D_cache/cache_reg[2][70]  ( .D(\D_cache/n1234 ), .CK(clk), .RN(n4200), .Q(\D_cache/cache[2][70] ) );
  DFFRX1 \D_cache/cache_reg[6][70]  ( .D(\D_cache/n1230 ), .CK(clk), .RN(n4201), .Q(\D_cache/cache[6][70] ) );
  DFFRX1 \D_cache/cache_reg[2][71]  ( .D(\D_cache/n1226 ), .CK(clk), .RN(n4201), .Q(\D_cache/cache[2][71] ) );
  DFFRX1 \D_cache/cache_reg[6][71]  ( .D(\D_cache/n1222 ), .CK(clk), .RN(n4201), .Q(\D_cache/cache[6][71] ) );
  DFFRX1 \D_cache/cache_reg[2][72]  ( .D(\D_cache/n1218 ), .CK(clk), .RN(n4202), .Q(\D_cache/cache[2][72] ) );
  DFFRX1 \D_cache/cache_reg[6][72]  ( .D(\D_cache/n1214 ), .CK(clk), .RN(n4202), .Q(\D_cache/cache[6][72] ) );
  DFFRX1 \D_cache/cache_reg[2][73]  ( .D(\D_cache/n1210 ), .CK(clk), .RN(n4202), .Q(\D_cache/cache[2][73] ) );
  DFFRX1 \D_cache/cache_reg[6][73]  ( .D(\D_cache/n1206 ), .CK(clk), .RN(n4203), .Q(\D_cache/cache[6][73] ) );
  DFFRX1 \D_cache/cache_reg[2][74]  ( .D(\D_cache/n1202 ), .CK(clk), .RN(n4203), .Q(\D_cache/cache[2][74] ) );
  DFFRX1 \D_cache/cache_reg[6][74]  ( .D(\D_cache/n1198 ), .CK(clk), .RN(n4203), .Q(\D_cache/cache[6][74] ) );
  DFFRX1 \D_cache/cache_reg[2][75]  ( .D(\D_cache/n1194 ), .CK(clk), .RN(n4204), .Q(\D_cache/cache[2][75] ) );
  DFFRX1 \D_cache/cache_reg[6][75]  ( .D(\D_cache/n1190 ), .CK(clk), .RN(n4204), .Q(\D_cache/cache[6][75] ) );
  DFFRX1 \D_cache/cache_reg[2][76]  ( .D(\D_cache/n1186 ), .CK(clk), .RN(n4204), .Q(\D_cache/cache[2][76] ) );
  DFFRX1 \D_cache/cache_reg[6][76]  ( .D(\D_cache/n1182 ), .CK(clk), .RN(n4205), .Q(\D_cache/cache[6][76] ) );
  DFFRX1 \D_cache/cache_reg[2][77]  ( .D(\D_cache/n1178 ), .CK(clk), .RN(n4205), .Q(\D_cache/cache[2][77] ) );
  DFFRX1 \D_cache/cache_reg[6][77]  ( .D(\D_cache/n1174 ), .CK(clk), .RN(n4205), .Q(\D_cache/cache[6][77] ) );
  DFFRX1 \D_cache/cache_reg[2][96]  ( .D(\D_cache/n1026 ), .CK(clk), .RN(n4218), .Q(\D_cache/cache[2][96] ) );
  DFFRX1 \D_cache/cache_reg[6][96]  ( .D(\D_cache/n1022 ), .CK(clk), .RN(n4218), .Q(\D_cache/cache[6][96] ) );
  DFFRX1 \D_cache/cache_reg[2][98]  ( .D(\D_cache/n1010 ), .CK(clk), .RN(n4219), .Q(\D_cache/cache[2][98] ) );
  DFFRX1 \D_cache/cache_reg[6][98]  ( .D(\D_cache/n1006 ), .CK(clk), .RN(n4219), .Q(\D_cache/cache[6][98] ) );
  DFFRX1 \D_cache/cache_reg[6][99]  ( .D(\D_cache/n998 ), .CK(clk), .RN(n4220), 
        .Q(\D_cache/cache[6][99] ) );
  DFFRX1 \D_cache/cache_reg[2][100]  ( .D(\D_cache/n994 ), .CK(clk), .RN(n4220), .Q(\D_cache/cache[2][100] ) );
  DFFRX1 \D_cache/cache_reg[6][100]  ( .D(\D_cache/n990 ), .CK(clk), .RN(n4221), .Q(\D_cache/cache[6][100] ) );
  DFFRX1 \D_cache/cache_reg[2][101]  ( .D(\D_cache/n986 ), .CK(clk), .RN(n4221), .Q(\D_cache/cache[2][101] ) );
  DFFRX1 \D_cache/cache_reg[6][101]  ( .D(\D_cache/n982 ), .CK(clk), .RN(n4221), .Q(\D_cache/cache[6][101] ) );
  DFFRX1 \D_cache/cache_reg[2][102]  ( .D(\D_cache/n978 ), .CK(clk), .RN(n4222), .Q(\D_cache/cache[2][102] ) );
  DFFRX1 \D_cache/cache_reg[6][102]  ( .D(\D_cache/n974 ), .CK(clk), .RN(n4222), .Q(\D_cache/cache[6][102] ) );
  DFFRX1 \D_cache/cache_reg[2][103]  ( .D(\D_cache/n970 ), .CK(clk), .RN(n4222), .Q(\D_cache/cache[2][103] ) );
  DFFRX1 \D_cache/cache_reg[6][103]  ( .D(\D_cache/n966 ), .CK(clk), .RN(n4223), .Q(\D_cache/cache[6][103] ) );
  DFFRX1 \D_cache/cache_reg[2][104]  ( .D(\D_cache/n962 ), .CK(clk), .RN(n4223), .Q(\D_cache/cache[2][104] ) );
  DFFRX1 \D_cache/cache_reg[6][104]  ( .D(\D_cache/n958 ), .CK(clk), .RN(n4223), .Q(\D_cache/cache[6][104] ) );
  DFFRX1 \D_cache/cache_reg[2][105]  ( .D(\D_cache/n954 ), .CK(clk), .RN(n4224), .Q(\D_cache/cache[2][105] ) );
  DFFRX1 \D_cache/cache_reg[6][105]  ( .D(\D_cache/n950 ), .CK(clk), .RN(n4224), .Q(\D_cache/cache[6][105] ) );
  DFFRX1 \D_cache/cache_reg[2][106]  ( .D(\D_cache/n946 ), .CK(clk), .RN(n4224), .Q(\D_cache/cache[2][106] ) );
  DFFRX1 \D_cache/cache_reg[6][106]  ( .D(\D_cache/n942 ), .CK(clk), .RN(n4225), .Q(\D_cache/cache[6][106] ) );
  DFFRX1 \D_cache/cache_reg[2][107]  ( .D(\D_cache/n938 ), .CK(clk), .RN(n4225), .Q(\D_cache/cache[2][107] ) );
  DFFRX1 \D_cache/cache_reg[6][107]  ( .D(\D_cache/n934 ), .CK(clk), .RN(n4225), .Q(\D_cache/cache[6][107] ) );
  DFFRX1 \D_cache/cache_reg[2][108]  ( .D(\D_cache/n930 ), .CK(clk), .RN(n4226), .Q(\D_cache/cache[2][108] ) );
  DFFRX1 \D_cache/cache_reg[6][108]  ( .D(\D_cache/n926 ), .CK(clk), .RN(n4226), .Q(\D_cache/cache[6][108] ) );
  DFFRX1 \D_cache/cache_reg[2][109]  ( .D(\D_cache/n922 ), .CK(clk), .RN(n4226), .Q(\D_cache/cache[2][109] ) );
  DFFRX1 \D_cache/cache_reg[6][109]  ( .D(\D_cache/n918 ), .CK(clk), .RN(n4227), .Q(\D_cache/cache[6][109] ) );
  DFFRX1 \D_cache/cache_reg[2][110]  ( .D(\D_cache/n914 ), .CK(clk), .RN(n4227), .Q(\D_cache/cache[2][110] ) );
  DFFRX1 \D_cache/cache_reg[6][110]  ( .D(\D_cache/n910 ), .CK(clk), .RN(n4227), .Q(\D_cache/cache[6][110] ) );
  DFFRX1 \D_cache/cache_reg[2][118]  ( .D(\D_cache/n850 ), .CK(clk), .RN(n4232), .Q(\D_cache/cache[2][118] ) );
  DFFRX1 \D_cache/cache_reg[6][118]  ( .D(\D_cache/n846 ), .CK(clk), .RN(n4233), .Q(\D_cache/cache[6][118] ) );
  DFFRX1 \D_cache/cache_reg[2][135]  ( .D(\D_cache/n714 ), .CK(clk), .RN(n4244), .Q(\D_cache/cache[2][135] ) );
  DFFRX1 \D_cache/cache_reg[6][135]  ( .D(\D_cache/n710 ), .CK(clk), .RN(n4244), .Q(\D_cache/cache[6][135] ) );
  DFFRX1 \D_cache/cache_reg[2][136]  ( .D(\D_cache/n706 ), .CK(clk), .RN(n4244), .Q(\D_cache/cache[2][136] ) );
  DFFRX1 \D_cache/cache_reg[6][136]  ( .D(\D_cache/n702 ), .CK(clk), .RN(n4245), .Q(\D_cache/cache[6][136] ) );
  DFFRX1 \D_cache/cache_reg[2][137]  ( .D(\D_cache/n698 ), .CK(clk), .RN(n4245), .Q(\D_cache/cache[2][137] ) );
  DFFRX1 \D_cache/cache_reg[6][137]  ( .D(\D_cache/n694 ), .CK(clk), .RN(n4245), .Q(\D_cache/cache[6][137] ) );
  DFFRX1 \D_cache/cache_reg[6][139]  ( .D(\D_cache/n678 ), .CK(clk), .RN(n4247), .Q(\D_cache/cache[6][139] ) );
  DFFRX1 \D_cache/cache_reg[2][149]  ( .D(\D_cache/n602 ), .CK(clk), .RN(n4253), .Q(\D_cache/cache[2][149] ) );
  DFFRX1 \D_cache/cache_reg[6][149]  ( .D(\D_cache/n598 ), .CK(clk), .RN(n4253), .Q(\D_cache/cache[6][149] ) );
  DFFRX1 \D_cache/cache_reg[6][151]  ( .D(\D_cache/n582 ), .CK(clk), .RN(n4255), .Q(\D_cache/cache[6][151] ) );
  DFFRX1 \D_cache/cache_reg[2][153]  ( .D(\D_cache/n570 ), .CK(clk), .RN(n4256), .Q(\D_cache/cache[2][153] ) );
  DFFRX1 \D_cache/cache_reg[6][153]  ( .D(\D_cache/n566 ), .CK(clk), .RN(n4256), .Q(\D_cache/cache[6][153] ) );
  DFFRX1 \D_cache/cache_reg[2][154]  ( .D(\D_cache/n562 ), .CK(clk), .RN(n4256), .Q(\D_cache/cache[2][154] ) );
  DFFRX1 \D_cache/cache_reg[6][154]  ( .D(\D_cache/n558 ), .CK(clk), .RN(n4257), .Q(\D_cache/cache[6][154] ) );
  DFFRX1 \I_cache/cache_reg[0][154]  ( .D(n8932), .CK(clk), .RN(n4360), .Q(
        \I_cache/cache[0][154] ), .QN(n1598) );
  DFFRX1 \I_cache/cache_reg[1][154]  ( .D(n8931), .CK(clk), .RN(n4360), .Q(
        \I_cache/cache[1][154] ), .QN(n177) );
  DFFRX1 \I_cache/cache_reg[2][154]  ( .D(n8930), .CK(clk), .RN(n4360), .Q(
        \I_cache/cache[2][154] ), .QN(n1599) );
  DFFRX1 \I_cache/cache_reg[3][154]  ( .D(n8929), .CK(clk), .RN(n4360), .Q(
        \I_cache/cache[3][154] ), .QN(n178) );
  DFFRX1 \I_cache/cache_reg[4][154]  ( .D(n8928), .CK(clk), .RN(n4360), .Q(
        \I_cache/cache[4][154] ), .QN(n463) );
  DFFRX1 \I_cache/cache_reg[5][154]  ( .D(n8927), .CK(clk), .RN(n4360), .Q(
        \I_cache/cache[5][154] ), .QN(n1372) );
  DFFRX1 \I_cache/cache_reg[6][154]  ( .D(n8926), .CK(clk), .RN(n4360), .Q(
        \I_cache/cache[6][154] ), .QN(n176) );
  DFFRX1 \I_cache/cache_reg[7][154]  ( .D(n8925), .CK(clk), .RN(n4360), .Q(
        \I_cache/cache[7][154] ), .QN(n1069) );
  DFFRX1 \i_MIPS/Register/register_reg[29][5]  ( .D(\i_MIPS/Register/n185 ), 
        .CK(clk), .RN(n4074), .Q(\i_MIPS/Register/register[29][5] ), .QN(n258)
         );
  DFFRX1 \i_MIPS/Register/register_reg[29][6]  ( .D(\i_MIPS/Register/n186 ), 
        .CK(clk), .RN(n4074), .Q(\i_MIPS/Register/register[29][6] ), .QN(n268)
         );
  DFFRX1 \i_MIPS/Register/register_reg[29][8]  ( .D(\i_MIPS/Register/n188 ), 
        .CK(clk), .RN(n4074), .Q(\i_MIPS/Register/register[29][8] ), .QN(n211)
         );
  DFFRX1 \i_MIPS/Register/register_reg[29][9]  ( .D(\i_MIPS/Register/n189 ), 
        .CK(clk), .RN(n4074), .Q(\i_MIPS/Register/register[29][9] ), .QN(n235)
         );
  DFFRX1 \i_MIPS/Register/register_reg[29][10]  ( .D(\i_MIPS/Register/n190 ), 
        .CK(clk), .RN(n4074), .Q(\i_MIPS/Register/register[29][10] ), .QN(n253) );
  DFFRX1 \i_MIPS/Register/register_reg[29][14]  ( .D(\i_MIPS/Register/n194 ), 
        .CK(clk), .RN(n4075), .Q(\i_MIPS/Register/register[29][14] ), .QN(n240) );
  DFFRX1 \i_MIPS/Register/register_reg[27][8]  ( .D(\i_MIPS/Register/n252 ), 
        .CK(clk), .RN(n4080), .Q(\i_MIPS/Register/register[27][8] ), .QN(n210)
         );
  DFFRX1 \i_MIPS/Register/register_reg[27][9]  ( .D(\i_MIPS/Register/n253 ), 
        .CK(clk), .RN(n4080), .Q(\i_MIPS/Register/register[27][9] ), .QN(n234)
         );
  DFFRX1 \i_MIPS/Register/register_reg[27][14]  ( .D(\i_MIPS/Register/n258 ), 
        .CK(clk), .RN(n4080), .Q(\i_MIPS/Register/register[27][14] ), .QN(n239) );
  DFFRX1 \i_MIPS/Register/register_reg[25][5]  ( .D(\i_MIPS/Register/n313 ), 
        .CK(clk), .RN(n4085), .Q(\i_MIPS/Register/register[25][5] ), .QN(n387)
         );
  DFFRX1 \i_MIPS/Register/register_reg[25][6]  ( .D(\i_MIPS/Register/n314 ), 
        .CK(clk), .RN(n4085), .Q(\i_MIPS/Register/register[25][6] ), .QN(n391)
         );
  DFFRX1 \i_MIPS/Register/register_reg[25][7]  ( .D(\i_MIPS/Register/n315 ), 
        .CK(clk), .RN(n4085), .Q(\i_MIPS/Register/register[25][7] ), .QN(n389)
         );
  DFFRX1 \i_MIPS/Register/register_reg[25][8]  ( .D(\i_MIPS/Register/n316 ), 
        .CK(clk), .RN(n4085), .Q(\i_MIPS/Register/register[25][8] ), .QN(n218)
         );
  DFFRX1 \i_MIPS/Register/register_reg[25][9]  ( .D(\i_MIPS/Register/n317 ), 
        .CK(clk), .RN(n4085), .Q(\i_MIPS/Register/register[25][9] ), .QN(n379)
         );
  DFFRX1 \i_MIPS/Register/register_reg[25][10]  ( .D(\i_MIPS/Register/n318 ), 
        .CK(clk), .RN(n4085), .Q(\i_MIPS/Register/register[25][10] ), .QN(n385) );
  DFFRX1 \i_MIPS/Register/register_reg[25][12]  ( .D(\i_MIPS/Register/n320 ), 
        .CK(clk), .RN(n4085), .Q(\i_MIPS/Register/register[25][12] ), .QN(n377) );
  DFFRX1 \i_MIPS/Register/register_reg[25][14]  ( .D(\i_MIPS/Register/n322 ), 
        .CK(clk), .RN(n4085), .Q(\i_MIPS/Register/register[25][14] ), .QN(n381) );
  DFFRX1 \i_MIPS/Register/register_reg[23][8]  ( .D(\i_MIPS/Register/n380 ), 
        .CK(clk), .RN(n4090), .Q(\i_MIPS/Register/register[23][8] ), .QN(n1093) );
  DFFRX1 \i_MIPS/Register/register_reg[21][5]  ( .D(\i_MIPS/Register/n441 ), 
        .CK(clk), .RN(n4095), .Q(\i_MIPS/Register/register[21][5] ), .QN(n1149) );
  DFFRX1 \i_MIPS/Register/register_reg[21][6]  ( .D(\i_MIPS/Register/n442 ), 
        .CK(clk), .RN(n4095), .Q(\i_MIPS/Register/register[21][6] ), .QN(n1161) );
  DFFRX1 \i_MIPS/Register/register_reg[21][7]  ( .D(\i_MIPS/Register/n443 ), 
        .CK(clk), .RN(n4095), .Q(\i_MIPS/Register/register[21][7] ), .QN(n1155) );
  DFFRX1 \i_MIPS/Register/register_reg[21][8]  ( .D(\i_MIPS/Register/n444 ), 
        .CK(clk), .RN(n4096), .Q(\i_MIPS/Register/register[21][8] ), .QN(n1095) );
  DFFRX1 \i_MIPS/Register/register_reg[21][9]  ( .D(\i_MIPS/Register/n445 ), 
        .CK(clk), .RN(n4096), .Q(\i_MIPS/Register/register[21][9] ), .QN(n1121) );
  DFFRX1 \i_MIPS/Register/register_reg[21][10]  ( .D(\i_MIPS/Register/n446 ), 
        .CK(clk), .RN(n4096), .Q(\i_MIPS/Register/register[21][10] ), .QN(
        n1143) );
  DFFRX1 \i_MIPS/Register/register_reg[21][11]  ( .D(\i_MIPS/Register/n447 ), 
        .CK(clk), .RN(n4096), .Q(\i_MIPS/Register/register[21][11] ), .QN(n224) );
  DFFRX1 \i_MIPS/Register/register_reg[21][12]  ( .D(\i_MIPS/Register/n448 ), 
        .CK(clk), .RN(n4096), .Q(\i_MIPS/Register/register[21][12] ), .QN(
        n1115) );
  DFFRX1 \i_MIPS/Register/register_reg[21][13]  ( .D(\i_MIPS/Register/n449 ), 
        .CK(clk), .RN(n4096), .Q(\i_MIPS/Register/register[21][13] ), .QN(
        n1100) );
  DFFRX1 \i_MIPS/Register/register_reg[21][14]  ( .D(\i_MIPS/Register/n450 ), 
        .CK(clk), .RN(n4096), .Q(\i_MIPS/Register/register[21][14] ), .QN(
        n1127) );
  DFFRX1 \i_MIPS/Register/register_reg[19][5]  ( .D(\i_MIPS/Register/n505 ), 
        .CK(clk), .RN(n4101), .Q(\i_MIPS/Register/register[19][5] ), .QN(n1148) );
  DFFRX1 \i_MIPS/Register/register_reg[19][6]  ( .D(\i_MIPS/Register/n506 ), 
        .CK(clk), .RN(n4101), .Q(\i_MIPS/Register/register[19][6] ), .QN(n1160) );
  DFFRX1 \i_MIPS/Register/register_reg[19][8]  ( .D(\i_MIPS/Register/n508 ), 
        .CK(clk), .RN(n4101), .Q(\i_MIPS/Register/register[19][8] ), .QN(n1094) );
  DFFRX1 \i_MIPS/Register/register_reg[19][9]  ( .D(\i_MIPS/Register/n509 ), 
        .CK(clk), .RN(n4101), .Q(\i_MIPS/Register/register[19][9] ), .QN(n1120) );
  DFFRX1 \i_MIPS/Register/register_reg[19][10]  ( .D(\i_MIPS/Register/n510 ), 
        .CK(clk), .RN(n4101), .Q(\i_MIPS/Register/register[19][10] ), .QN(
        n1142) );
  DFFRX1 \i_MIPS/Register/register_reg[19][14]  ( .D(\i_MIPS/Register/n514 ), 
        .CK(clk), .RN(n4101), .Q(\i_MIPS/Register/register[19][14] ), .QN(
        n1126) );
  DFFRX1 \i_MIPS/Register/register_reg[17][2]  ( .D(\i_MIPS/Register/n566 ), 
        .CK(clk), .RN(n4106), .Q(\i_MIPS/Register/register[17][2] ), .QN(n1310) );
  DFFRX1 \i_MIPS/Register/register_reg[17][3]  ( .D(\i_MIPS/Register/n567 ), 
        .CK(clk), .RN(n4106), .Q(\i_MIPS/Register/register[17][3] ), .QN(n1312) );
  DFFRX1 \i_MIPS/Register/register_reg[17][4]  ( .D(\i_MIPS/Register/n568 ), 
        .CK(clk), .RN(n4106), .Q(\i_MIPS/Register/register[17][4] ), .QN(n1297) );
  DFFRX1 \i_MIPS/Register/register_reg[17][5]  ( .D(\i_MIPS/Register/n569 ), 
        .CK(clk), .RN(n4106), .Q(\i_MIPS/Register/register[17][5] ), .QN(n1301) );
  DFFRX1 \i_MIPS/Register/register_reg[17][6]  ( .D(\i_MIPS/Register/n570 ), 
        .CK(clk), .RN(n4106), .Q(\i_MIPS/Register/register[17][6] ), .QN(n1305) );
  DFFRX1 \i_MIPS/Register/register_reg[17][7]  ( .D(\i_MIPS/Register/n571 ), 
        .CK(clk), .RN(n4106), .Q(\i_MIPS/Register/register[17][7] ), .QN(n1303) );
  DFFRX1 \i_MIPS/Register/register_reg[17][8]  ( .D(\i_MIPS/Register/n572 ), 
        .CK(clk), .RN(n4106), .Q(\i_MIPS/Register/register[17][8] ), .QN(n1103) );
  DFFRX1 \i_MIPS/Register/register_reg[17][9]  ( .D(\i_MIPS/Register/n573 ), 
        .CK(clk), .RN(n4106), .Q(\i_MIPS/Register/register[17][9] ), .QN(n1293) );
  DFFRX1 \i_MIPS/Register/register_reg[17][10]  ( .D(\i_MIPS/Register/n574 ), 
        .CK(clk), .RN(n4106), .Q(\i_MIPS/Register/register[17][10] ), .QN(
        n1299) );
  DFFRX1 \i_MIPS/Register/register_reg[17][11]  ( .D(\i_MIPS/Register/n575 ), 
        .CK(clk), .RN(n4106), .Q(\i_MIPS/Register/register[17][11] ), .QN(n226) );
  DFFRX1 \i_MIPS/Register/register_reg[17][12]  ( .D(\i_MIPS/Register/n576 ), 
        .CK(clk), .RN(n4107), .Q(\i_MIPS/Register/register[17][12] ), .QN(
        n1291) );
  DFFRX1 \i_MIPS/Register/register_reg[17][13]  ( .D(\i_MIPS/Register/n577 ), 
        .CK(clk), .RN(n4107), .Q(\i_MIPS/Register/register[17][13] ), .QN(
        n1105) );
  DFFRX1 \i_MIPS/Register/register_reg[17][14]  ( .D(\i_MIPS/Register/n578 ), 
        .CK(clk), .RN(n4107), .Q(\i_MIPS/Register/register[17][14] ), .QN(
        n1295) );
  DFFRX1 \i_MIPS/Register/register_reg[13][5]  ( .D(\i_MIPS/Register/n697 ), 
        .CK(clk), .RN(n4117), .Q(\i_MIPS/Register/register[13][5] ), .QN(n261)
         );
  DFFRX1 \i_MIPS/Register/register_reg[13][6]  ( .D(\i_MIPS/Register/n698 ), 
        .CK(clk), .RN(n4117), .Q(\i_MIPS/Register/register[13][6] ), .QN(n271)
         );
  DFFRX1 \i_MIPS/Register/register_reg[13][8]  ( .D(\i_MIPS/Register/n700 ), 
        .CK(clk), .RN(n4117), .Q(\i_MIPS/Register/register[13][8] ), .QN(n213)
         );
  DFFRX1 \i_MIPS/Register/register_reg[13][9]  ( .D(\i_MIPS/Register/n701 ), 
        .CK(clk), .RN(n4117), .Q(\i_MIPS/Register/register[13][9] ), .QN(n238)
         );
  DFFRX1 \i_MIPS/Register/register_reg[13][10]  ( .D(\i_MIPS/Register/n702 ), 
        .CK(clk), .RN(n4117), .Q(\i_MIPS/Register/register[13][10] ), .QN(n256) );
  DFFRX1 \i_MIPS/Register/register_reg[13][14]  ( .D(\i_MIPS/Register/n706 ), 
        .CK(clk), .RN(n4117), .Q(\i_MIPS/Register/register[13][14] ), .QN(n243) );
  DFFRX1 \i_MIPS/Register/register_reg[11][8]  ( .D(\i_MIPS/Register/n764 ), 
        .CK(clk), .RN(n4122), .Q(\i_MIPS/Register/register[11][8] ), .QN(n212)
         );
  DFFRX1 \i_MIPS/Register/register_reg[11][9]  ( .D(\i_MIPS/Register/n765 ), 
        .CK(clk), .RN(n4122), .Q(\i_MIPS/Register/register[11][9] ), .QN(n237)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][5]  ( .D(\i_MIPS/Register/n825 ), 
        .CK(clk), .RN(n4127), .Q(\i_MIPS/Register/register[9][5] ), .QN(n388)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][6]  ( .D(\i_MIPS/Register/n826 ), 
        .CK(clk), .RN(n4127), .Q(\i_MIPS/Register/register[9][6] ), .QN(n392)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][7]  ( .D(\i_MIPS/Register/n827 ), 
        .CK(clk), .RN(n4127), .Q(\i_MIPS/Register/register[9][7] ), .QN(n390)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][8]  ( .D(\i_MIPS/Register/n828 ), 
        .CK(clk), .RN(n4128), .Q(\i_MIPS/Register/register[9][8] ), .QN(n219)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][9]  ( .D(\i_MIPS/Register/n829 ), 
        .CK(clk), .RN(n4128), .Q(\i_MIPS/Register/register[9][9] ), .QN(n380)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][10]  ( .D(\i_MIPS/Register/n830 ), 
        .CK(clk), .RN(n4128), .Q(\i_MIPS/Register/register[9][10] ), .QN(n386)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][12]  ( .D(\i_MIPS/Register/n832 ), 
        .CK(clk), .RN(n4128), .Q(\i_MIPS/Register/register[9][12] ), .QN(n378)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][14]  ( .D(\i_MIPS/Register/n834 ), 
        .CK(clk), .RN(n4128), .Q(\i_MIPS/Register/register[9][14] ), .QN(n382)
         );
  DFFRX1 \i_MIPS/Register/register_reg[7][8]  ( .D(\i_MIPS/Register/n892 ), 
        .CK(clk), .RN(n4133), .Q(\i_MIPS/Register/register[7][8] ), .QN(n222)
         );
  DFFRX1 \i_MIPS/Register/register_reg[5][6]  ( .D(\i_MIPS/Register/n954 ), 
        .CK(clk), .RN(n4138), .Q(\i_MIPS/Register/register[5][6] ), .QN(n1164)
         );
  DFFRX1 \i_MIPS/Register/register_reg[5][7]  ( .D(\i_MIPS/Register/n955 ), 
        .CK(clk), .RN(n4138), .Q(\i_MIPS/Register/register[5][7] ), .QN(n1158)
         );
  DFFRX1 \i_MIPS/Register/register_reg[5][8]  ( .D(\i_MIPS/Register/n956 ), 
        .CK(clk), .RN(n4138), .Q(\i_MIPS/Register/register[5][8] ), .QN(n1097)
         );
  DFFRX1 \i_MIPS/Register/register_reg[5][9]  ( .D(\i_MIPS/Register/n957 ), 
        .CK(clk), .RN(n4138), .Q(\i_MIPS/Register/register[5][9] ), .QN(n1124)
         );
  DFFRX1 \i_MIPS/Register/register_reg[5][10]  ( .D(\i_MIPS/Register/n958 ), 
        .CK(clk), .RN(n4138), .Q(\i_MIPS/Register/register[5][10] ), .QN(n1146) );
  DFFRX1 \i_MIPS/Register/register_reg[5][11]  ( .D(\i_MIPS/Register/n959 ), 
        .CK(clk), .RN(n4138), .Q(\i_MIPS/Register/register[5][11] ), .QN(n225)
         );
  DFFRX1 \i_MIPS/Register/register_reg[5][13]  ( .D(\i_MIPS/Register/n961 ), 
        .CK(clk), .RN(n4139), .Q(\i_MIPS/Register/register[5][13] ), .QN(n1102) );
  DFFRX1 \i_MIPS/Register/register_reg[5][14]  ( .D(\i_MIPS/Register/n962 ), 
        .CK(clk), .RN(n4139), .Q(\i_MIPS/Register/register[5][14] ), .QN(n1130) );
  DFFRX1 \i_MIPS/Register/register_reg[3][6]  ( .D(\i_MIPS/Register/n1018 ), 
        .CK(clk), .RN(n4143), .Q(\i_MIPS/Register/register[3][6] ), .QN(n1163)
         );
  DFFRX1 \i_MIPS/Register/register_reg[3][8]  ( .D(\i_MIPS/Register/n1020 ), 
        .CK(clk), .RN(n4144), .Q(\i_MIPS/Register/register[3][8] ), .QN(n1096)
         );
  DFFRX1 \i_MIPS/Register/register_reg[3][9]  ( .D(\i_MIPS/Register/n1021 ), 
        .CK(clk), .RN(n4144), .Q(\i_MIPS/Register/register[3][9] ), .QN(n1123)
         );
  DFFRX1 \i_MIPS/Register/register_reg[3][10]  ( .D(\i_MIPS/Register/n1022 ), 
        .CK(clk), .RN(n4144), .Q(\i_MIPS/Register/register[3][10] ), .QN(n1145) );
  DFFRX1 \i_MIPS/Register/register_reg[3][14]  ( .D(\i_MIPS/Register/n1026 ), 
        .CK(clk), .RN(n4144), .Q(\i_MIPS/Register/register[3][14] ), .QN(n1129) );
  DFFRX1 \i_MIPS/Register/register_reg[1][2]  ( .D(\i_MIPS/Register/n1078 ), 
        .CK(clk), .RN(n4148), .Q(\i_MIPS/Register/register[1][2] ), .QN(n1311)
         );
  DFFRX1 \i_MIPS/Register/register_reg[1][3]  ( .D(\i_MIPS/Register/n1079 ), 
        .CK(clk), .RN(n4148), .Q(\i_MIPS/Register/register[1][3] ), .QN(n1313)
         );
  DFFRX1 \i_MIPS/Register/register_reg[1][6]  ( .D(\i_MIPS/Register/n1082 ), 
        .CK(clk), .RN(n4149), .Q(\i_MIPS/Register/register[1][6] ), .QN(n1306)
         );
  DFFRX1 \i_MIPS/Register/register_reg[1][7]  ( .D(\i_MIPS/Register/n1083 ), 
        .CK(clk), .RN(n4149), .Q(\i_MIPS/Register/register[1][7] ), .QN(n1304)
         );
  DFFRX1 \i_MIPS/Register/register_reg[1][8]  ( .D(\i_MIPS/Register/n1084 ), 
        .CK(clk), .RN(n4149), .Q(\i_MIPS/Register/register[1][8] ), .QN(n1104)
         );
  DFFRX1 \i_MIPS/Register/register_reg[1][9]  ( .D(\i_MIPS/Register/n1085 ), 
        .CK(clk), .RN(n4149), .Q(\i_MIPS/Register/register[1][9] ), .QN(n1294)
         );
  DFFRX1 \i_MIPS/Register/register_reg[1][10]  ( .D(\i_MIPS/Register/n1086 ), 
        .CK(clk), .RN(n4149), .Q(\i_MIPS/Register/register[1][10] ), .QN(n1300) );
  DFFRX1 \i_MIPS/Register/register_reg[1][11]  ( .D(\i_MIPS/Register/n1087 ), 
        .CK(clk), .RN(n4149), .Q(\i_MIPS/Register/register[1][11] ), .QN(n227)
         );
  DFFRX1 \i_MIPS/Register/register_reg[1][13]  ( .D(\i_MIPS/Register/n1089 ), 
        .CK(clk), .RN(n4149), .Q(\i_MIPS/Register/register[1][13] ), .QN(n1106) );
  DFFRX1 \i_MIPS/Register/register_reg[1][14]  ( .D(\i_MIPS/Register/n1090 ), 
        .CK(clk), .RN(n4149), .Q(\i_MIPS/Register/register[1][14] ), .QN(n1296) );
  DFFRX1 \I_cache/cache_reg[0][0]  ( .D(n10163), .CK(clk), .RN(n4257), .Q(
        \I_cache/cache[0][0] ), .QN(n679) );
  DFFRX1 \I_cache/cache_reg[1][0]  ( .D(n10162), .CK(clk), .RN(n4257), .Q(
        \I_cache/cache[1][0] ), .QN(n1600) );
  DFFRX1 \I_cache/cache_reg[2][0]  ( .D(n10161), .CK(clk), .RN(n4257), .Q(
        \I_cache/cache[2][0] ), .QN(n680) );
  DFFRX1 \I_cache/cache_reg[3][0]  ( .D(n10160), .CK(clk), .RN(n4257), .Q(
        \I_cache/cache[3][0] ), .QN(n1602) );
  DFFRX1 \I_cache/cache_reg[4][0]  ( .D(n10159), .CK(clk), .RN(n4257), .Q(
        \I_cache/cache[4][0] ), .QN(n684) );
  DFFRX1 \I_cache/cache_reg[5][0]  ( .D(n10158), .CK(clk), .RN(n4257), .Q(
        \I_cache/cache[5][0] ), .QN(n1601) );
  DFFRX1 \I_cache/cache_reg[6][0]  ( .D(n10157), .CK(clk), .RN(n4257), .Q(
        \I_cache/cache[6][0] ), .QN(n691) );
  DFFRX1 \I_cache/cache_reg[7][0]  ( .D(n10164), .CK(clk), .RN(n4257), .Q(
        \I_cache/cache[7][0] ), .QN(n1612) );
  DFFRX1 \I_cache/cache_reg[0][1]  ( .D(n10156), .CK(clk), .RN(n4258), .Q(
        \I_cache/cache[0][1] ), .QN(n472) );
  DFFRX1 \I_cache/cache_reg[1][1]  ( .D(n10155), .CK(clk), .RN(n4258), .Q(
        \I_cache/cache[1][1] ), .QN(n1387) );
  DFFRX1 \I_cache/cache_reg[2][1]  ( .D(n10154), .CK(clk), .RN(n4258), .Q(
        \I_cache/cache[2][1] ), .QN(n474) );
  DFFRX1 \I_cache/cache_reg[3][1]  ( .D(n10153), .CK(clk), .RN(n4258), .Q(
        \I_cache/cache[3][1] ), .QN(n1389) );
  DFFRX1 \I_cache/cache_reg[4][1]  ( .D(n10152), .CK(clk), .RN(n4258), .Q(
        \I_cache/cache[4][1] ), .QN(n473) );
  DFFRX1 \I_cache/cache_reg[5][1]  ( .D(n10151), .CK(clk), .RN(n4258), .Q(
        \I_cache/cache[5][1] ), .QN(n1388) );
  DFFRX1 \I_cache/cache_reg[6][1]  ( .D(n10150), .CK(clk), .RN(n4258), .Q(
        \I_cache/cache[6][1] ), .QN(n640) );
  DFFRX1 \I_cache/cache_reg[7][1]  ( .D(n10149), .CK(clk), .RN(n4258), .Q(
        \I_cache/cache[7][1] ), .QN(n1559) );
  DFFRX1 \I_cache/cache_reg[0][2]  ( .D(n10148), .CK(clk), .RN(n4258), .Q(
        \I_cache/cache[0][2] ), .QN(n567) );
  DFFRX1 \I_cache/cache_reg[1][2]  ( .D(n10147), .CK(clk), .RN(n4258), .Q(
        \I_cache/cache[1][2] ), .QN(n1486) );
  DFFRX1 \I_cache/cache_reg[2][2]  ( .D(n10146), .CK(clk), .RN(n4258), .Q(
        \I_cache/cache[2][2] ), .QN(n569) );
  DFFRX1 \I_cache/cache_reg[3][2]  ( .D(n10145), .CK(clk), .RN(n4258), .Q(
        \I_cache/cache[3][2] ), .QN(n1488) );
  DFFRX1 \I_cache/cache_reg[4][2]  ( .D(n10144), .CK(clk), .RN(n4259), .Q(
        \I_cache/cache[4][2] ), .QN(n568) );
  DFFRX1 \I_cache/cache_reg[5][2]  ( .D(n10143), .CK(clk), .RN(n4259), .Q(
        \I_cache/cache[5][2] ), .QN(n1487) );
  DFFRX1 \I_cache/cache_reg[6][2]  ( .D(n10142), .CK(clk), .RN(n4259), .Q(
        \I_cache/cache[6][2] ), .QN(n677) );
  DFFRX1 \I_cache/cache_reg[7][2]  ( .D(n10141), .CK(clk), .RN(n4259), .Q(
        \I_cache/cache[7][2] ), .QN(n1596) );
  DFFRX1 \I_cache/cache_reg[0][3]  ( .D(n10140), .CK(clk), .RN(n4259), .Q(
        \I_cache/cache[0][3] ), .QN(n435) );
  DFFRX1 \I_cache/cache_reg[1][3]  ( .D(n10139), .CK(clk), .RN(n4259), .Q(
        \I_cache/cache[1][3] ), .QN(n1350) );
  DFFRX1 \I_cache/cache_reg[2][3]  ( .D(n10138), .CK(clk), .RN(n4259), .Q(
        \I_cache/cache[2][3] ), .QN(n434) );
  DFFRX1 \I_cache/cache_reg[3][3]  ( .D(n10137), .CK(clk), .RN(n4259), .Q(
        \I_cache/cache[3][3] ), .QN(n1349) );
  DFFRX1 \I_cache/cache_reg[4][3]  ( .D(n10136), .CK(clk), .RN(n4259), .Q(
        \I_cache/cache[4][3] ), .QN(n448) );
  DFFRX1 \I_cache/cache_reg[5][3]  ( .D(n10135), .CK(clk), .RN(n4259), .Q(
        \I_cache/cache[5][3] ), .QN(n1362) );
  DFFRX1 \I_cache/cache_reg[6][3]  ( .D(n10134), .CK(clk), .RN(n4259), .Q(
        \I_cache/cache[6][3] ), .QN(n446) );
  DFFRX1 \I_cache/cache_reg[7][3]  ( .D(n10133), .CK(clk), .RN(n4259), .Q(
        \I_cache/cache[7][3] ), .QN(n1361) );
  DFFRX1 \I_cache/cache_reg[0][4]  ( .D(n10132), .CK(clk), .RN(n4260), .Q(
        \I_cache/cache[0][4] ), .QN(n488) );
  DFFRX1 \I_cache/cache_reg[1][4]  ( .D(n10131), .CK(clk), .RN(n4260), .Q(
        \I_cache/cache[1][4] ), .QN(n1406) );
  DFFRX1 \I_cache/cache_reg[2][4]  ( .D(n10130), .CK(clk), .RN(n4260), .Q(
        \I_cache/cache[2][4] ), .QN(n487) );
  DFFRX1 \I_cache/cache_reg[3][4]  ( .D(n10129), .CK(clk), .RN(n4260), .Q(
        \I_cache/cache[3][4] ), .QN(n1405) );
  DFFRX1 \I_cache/cache_reg[4][4]  ( .D(n10128), .CK(clk), .RN(n4260), .Q(
        \I_cache/cache[4][4] ), .QN(n641) );
  DFFRX1 \I_cache/cache_reg[5][4]  ( .D(n10127), .CK(clk), .RN(n4260), .Q(
        \I_cache/cache[5][4] ), .QN(n1560) );
  DFFRX1 \I_cache/cache_reg[6][4]  ( .D(n10126), .CK(clk), .RN(n4260), .Q(
        \I_cache/cache[6][4] ), .QN(n534) );
  DFFRX1 \I_cache/cache_reg[7][4]  ( .D(n10125), .CK(clk), .RN(n4260), .Q(
        \I_cache/cache[7][4] ), .QN(n1453) );
  DFFRX1 \I_cache/cache_reg[0][5]  ( .D(n10124), .CK(clk), .RN(n4260), .Q(
        \I_cache/cache[0][5] ), .QN(n575) );
  DFFRX1 \I_cache/cache_reg[1][5]  ( .D(n10123), .CK(clk), .RN(n4260), .Q(
        \I_cache/cache[1][5] ), .QN(n1494) );
  DFFRX1 \I_cache/cache_reg[2][5]  ( .D(n10122), .CK(clk), .RN(n4260), .Q(
        \I_cache/cache[2][5] ), .QN(n573) );
  DFFRX1 \I_cache/cache_reg[3][5]  ( .D(n10121), .CK(clk), .RN(n4260), .Q(
        \I_cache/cache[3][5] ), .QN(n1492) );
  DFFRX1 \I_cache/cache_reg[4][5]  ( .D(n10120), .CK(clk), .RN(n4261), .Q(
        \I_cache/cache[4][5] ), .QN(n655) );
  DFFRX1 \I_cache/cache_reg[5][5]  ( .D(n10119), .CK(clk), .RN(n4261), .Q(
        \I_cache/cache[5][5] ), .QN(n1574) );
  DFFRX1 \I_cache/cache_reg[6][5]  ( .D(n10118), .CK(clk), .RN(n4261), .Q(
        \I_cache/cache[6][5] ), .QN(n574) );
  DFFRX1 \I_cache/cache_reg[7][5]  ( .D(n10117), .CK(clk), .RN(n4261), .Q(
        \I_cache/cache[7][5] ), .QN(n1493) );
  DFFRX1 \I_cache/cache_reg[0][6]  ( .D(n10116), .CK(clk), .RN(n4261), .Q(
        \I_cache/cache[0][6] ), .QN(n578) );
  DFFRX1 \I_cache/cache_reg[1][6]  ( .D(n10115), .CK(clk), .RN(n4261), .Q(
        \I_cache/cache[1][6] ), .QN(n1497) );
  DFFRX1 \I_cache/cache_reg[2][6]  ( .D(n10114), .CK(clk), .RN(n4261), .Q(
        \I_cache/cache[2][6] ), .QN(n577) );
  DFFRX1 \I_cache/cache_reg[3][6]  ( .D(n10113), .CK(clk), .RN(n4261), .Q(
        \I_cache/cache[3][6] ), .QN(n1496) );
  DFFRX1 \I_cache/cache_reg[4][6]  ( .D(n10112), .CK(clk), .RN(n4261), .Q(
        \I_cache/cache[4][6] ), .QN(n647) );
  DFFRX1 \I_cache/cache_reg[5][6]  ( .D(n10111), .CK(clk), .RN(n4261), .Q(
        \I_cache/cache[5][6] ), .QN(n1566) );
  DFFRX1 \I_cache/cache_reg[6][6]  ( .D(n10110), .CK(clk), .RN(n4261), .Q(
        \I_cache/cache[6][6] ), .QN(n576) );
  DFFRX1 \I_cache/cache_reg[7][6]  ( .D(n10109), .CK(clk), .RN(n4261), .Q(
        \I_cache/cache[7][6] ), .QN(n1495) );
  DFFRX1 \I_cache/cache_reg[0][7]  ( .D(n10108), .CK(clk), .RN(n4262), .Q(
        \I_cache/cache[0][7] ), .QN(n545) );
  DFFRX1 \I_cache/cache_reg[1][7]  ( .D(n10107), .CK(clk), .RN(n4262), .Q(
        \I_cache/cache[1][7] ), .QN(n1464) );
  DFFRX1 \I_cache/cache_reg[2][7]  ( .D(n10106), .CK(clk), .RN(n4262), .Q(
        \I_cache/cache[2][7] ), .QN(n537) );
  DFFRX1 \I_cache/cache_reg[3][7]  ( .D(n10105), .CK(clk), .RN(n4262), .Q(
        \I_cache/cache[3][7] ), .QN(n1456) );
  DFFRX1 \I_cache/cache_reg[4][7]  ( .D(n10104), .CK(clk), .RN(n4262), .Q(
        \I_cache/cache[4][7] ), .QN(n546) );
  DFFRX1 \I_cache/cache_reg[5][7]  ( .D(n10103), .CK(clk), .RN(n4262), .Q(
        \I_cache/cache[5][7] ), .QN(n1465) );
  DFFRX1 \I_cache/cache_reg[6][7]  ( .D(n10102), .CK(clk), .RN(n4262), .Q(
        \I_cache/cache[6][7] ), .QN(n538) );
  DFFRX1 \I_cache/cache_reg[7][7]  ( .D(n10101), .CK(clk), .RN(n4262), .Q(
        \I_cache/cache[7][7] ), .QN(n1457) );
  DFFRX1 \I_cache/cache_reg[0][8]  ( .D(n10100), .CK(clk), .RN(n4262), .Q(
        \I_cache/cache[0][8] ), .QN(n616) );
  DFFRX1 \I_cache/cache_reg[1][8]  ( .D(n10099), .CK(clk), .RN(n4262), .Q(
        \I_cache/cache[1][8] ), .QN(n1535) );
  DFFRX1 \I_cache/cache_reg[2][8]  ( .D(n10098), .CK(clk), .RN(n4262), .Q(
        \I_cache/cache[2][8] ), .QN(n615) );
  DFFRX1 \I_cache/cache_reg[3][8]  ( .D(n10097), .CK(clk), .RN(n4262), .Q(
        \I_cache/cache[3][8] ), .QN(n1534) );
  DFFRX1 \I_cache/cache_reg[4][8]  ( .D(n10096), .CK(clk), .RN(n4263), .Q(
        \I_cache/cache[4][8] ), .QN(n663) );
  DFFRX1 \I_cache/cache_reg[5][8]  ( .D(n10095), .CK(clk), .RN(n4263), .Q(
        \I_cache/cache[5][8] ), .QN(n1582) );
  DFFRX1 \I_cache/cache_reg[6][8]  ( .D(n10094), .CK(clk), .RN(n4263), .Q(
        \I_cache/cache[6][8] ), .QN(n617) );
  DFFRX1 \I_cache/cache_reg[7][8]  ( .D(n10093), .CK(clk), .RN(n4263), .Q(
        \I_cache/cache[7][8] ), .QN(n1536) );
  DFFRX1 \I_cache/cache_reg[0][9]  ( .D(n10092), .CK(clk), .RN(n4263), .Q(
        \I_cache/cache[0][9] ), .QN(n619) );
  DFFRX1 \I_cache/cache_reg[1][9]  ( .D(n10091), .CK(clk), .RN(n4263), .Q(
        \I_cache/cache[1][9] ), .QN(n1538) );
  DFFRX1 \I_cache/cache_reg[2][9]  ( .D(n10090), .CK(clk), .RN(n4263), .Q(
        \I_cache/cache[2][9] ), .QN(n618) );
  DFFRX1 \I_cache/cache_reg[3][9]  ( .D(n10089), .CK(clk), .RN(n4263), .Q(
        \I_cache/cache[3][9] ), .QN(n1537) );
  DFFRX1 \I_cache/cache_reg[4][9]  ( .D(n10088), .CK(clk), .RN(n4263), .Q(
        \I_cache/cache[4][9] ), .QN(n666) );
  DFFRX1 \I_cache/cache_reg[5][9]  ( .D(n10087), .CK(clk), .RN(n4263), .Q(
        \I_cache/cache[5][9] ), .QN(n1585) );
  DFFRX1 \I_cache/cache_reg[6][9]  ( .D(n10086), .CK(clk), .RN(n4263), .Q(
        \I_cache/cache[6][9] ), .QN(n620) );
  DFFRX1 \I_cache/cache_reg[7][9]  ( .D(n10085), .CK(clk), .RN(n4263), .Q(
        \I_cache/cache[7][9] ), .QN(n1539) );
  DFFRX1 \I_cache/cache_reg[3][10]  ( .D(n10081), .CK(clk), .RN(n4264), .Q(
        \I_cache/cache[3][10] ), .QN(n1550) );
  DFFRX1 \I_cache/cache_reg[5][10]  ( .D(n10079), .CK(clk), .RN(n4264), .Q(
        \I_cache/cache[5][10] ), .QN(n1589) );
  DFFRX1 \I_cache/cache_reg[7][10]  ( .D(n10077), .CK(clk), .RN(n4264), .Q(
        \I_cache/cache[7][10] ), .QN(n1549) );
  DFFRX1 \I_cache/cache_reg[0][11]  ( .D(n10076), .CK(clk), .RN(n4264), .Q(
        \I_cache/cache[0][11] ), .QN(n566) );
  DFFRX1 \I_cache/cache_reg[1][11]  ( .D(n10075), .CK(clk), .RN(n4264), .Q(
        \I_cache/cache[1][11] ), .QN(n1485) );
  DFFRX1 \I_cache/cache_reg[2][11]  ( .D(n10074), .CK(clk), .RN(n4264), .Q(
        \I_cache/cache[2][11] ), .QN(n565) );
  DFFRX1 \I_cache/cache_reg[3][11]  ( .D(n10073), .CK(clk), .RN(n4264), .Q(
        \I_cache/cache[3][11] ), .QN(n1484) );
  DFFRX1 \I_cache/cache_reg[4][11]  ( .D(n10072), .CK(clk), .RN(n4265), .Q(
        \I_cache/cache[4][11] ), .QN(n673) );
  DFFRX1 \I_cache/cache_reg[5][11]  ( .D(n10071), .CK(clk), .RN(n4265), .Q(
        \I_cache/cache[5][11] ), .QN(n1592) );
  DFFRX1 \I_cache/cache_reg[6][11]  ( .D(n10070), .CK(clk), .RN(n4265), .Q(
        \I_cache/cache[6][11] ), .QN(n564) );
  DFFRX1 \I_cache/cache_reg[7][11]  ( .D(n10069), .CK(clk), .RN(n4265), .Q(
        \I_cache/cache[7][11] ), .QN(n1483) );
  DFFRX1 \I_cache/cache_reg[0][12]  ( .D(n10068), .CK(clk), .RN(n4265), .Q(
        \I_cache/cache[0][12] ), .QN(n604) );
  DFFRX1 \I_cache/cache_reg[1][12]  ( .D(n10067), .CK(clk), .RN(n4265), .Q(
        \I_cache/cache[1][12] ), .QN(n1523) );
  DFFRX1 \I_cache/cache_reg[2][12]  ( .D(n10066), .CK(clk), .RN(n4265), .Q(
        \I_cache/cache[2][12] ), .QN(n603) );
  DFFRX1 \I_cache/cache_reg[3][12]  ( .D(n10065), .CK(clk), .RN(n4265), .Q(
        \I_cache/cache[3][12] ), .QN(n1522) );
  DFFRX1 \I_cache/cache_reg[4][12]  ( .D(n10064), .CK(clk), .RN(n4265), .Q(
        \I_cache/cache[4][12] ), .QN(n659) );
  DFFRX1 \I_cache/cache_reg[5][12]  ( .D(n10063), .CK(clk), .RN(n4265), .Q(
        \I_cache/cache[5][12] ), .QN(n1578) );
  DFFRX1 \I_cache/cache_reg[6][12]  ( .D(n10062), .CK(clk), .RN(n4265), .Q(
        \I_cache/cache[6][12] ), .QN(n605) );
  DFFRX1 \I_cache/cache_reg[7][12]  ( .D(n10061), .CK(clk), .RN(n4265), .Q(
        \I_cache/cache[7][12] ), .QN(n1524) );
  DFFRX1 \I_cache/cache_reg[0][13]  ( .D(n10060), .CK(clk), .RN(n4266), .Q(
        \I_cache/cache[0][13] ), .QN(n599) );
  DFFRX1 \I_cache/cache_reg[1][13]  ( .D(n10059), .CK(clk), .RN(n4266), .Q(
        \I_cache/cache[1][13] ), .QN(n1518) );
  DFFRX1 \I_cache/cache_reg[2][13]  ( .D(n10058), .CK(clk), .RN(n4266), .Q(
        \I_cache/cache[2][13] ), .QN(n598) );
  DFFRX1 \I_cache/cache_reg[3][13]  ( .D(n10057), .CK(clk), .RN(n4266), .Q(
        \I_cache/cache[3][13] ), .QN(n1517) );
  DFFRX1 \I_cache/cache_reg[4][13]  ( .D(n10056), .CK(clk), .RN(n4266), .Q(
        \I_cache/cache[4][13] ), .QN(n657) );
  DFFRX1 \I_cache/cache_reg[5][13]  ( .D(n10055), .CK(clk), .RN(n4266), .Q(
        \I_cache/cache[5][13] ), .QN(n1576) );
  DFFRX1 \I_cache/cache_reg[6][13]  ( .D(n10054), .CK(clk), .RN(n4266), .Q(
        \I_cache/cache[6][13] ), .QN(n597) );
  DFFRX1 \I_cache/cache_reg[7][13]  ( .D(n10053), .CK(clk), .RN(n4266), .Q(
        \I_cache/cache[7][13] ), .QN(n1516) );
  DFFRX1 \I_cache/cache_reg[1][14]  ( .D(n10051), .CK(clk), .RN(n4266), .Q(
        \I_cache/cache[1][14] ), .QN(n1438) );
  DFFRX1 \I_cache/cache_reg[3][14]  ( .D(n10049), .CK(clk), .RN(n4266), .Q(
        \I_cache/cache[3][14] ), .QN(n1437) );
  DFFRX1 \I_cache/cache_reg[4][14]  ( .D(n10048), .CK(clk), .RN(n4267), .Q(
        \I_cache/cache[4][14] ), .QN(n533) );
  DFFRX1 \I_cache/cache_reg[5][14]  ( .D(n10047), .CK(clk), .RN(n4267), .Q(
        \I_cache/cache[5][14] ), .QN(n1452) );
  DFFRX1 \I_cache/cache_reg[6][14]  ( .D(n10046), .CK(clk), .RN(n4267), .Q(
        \I_cache/cache[6][14] ), .QN(n518) );
  DFFRX1 \I_cache/cache_reg[7][14]  ( .D(n10045), .CK(clk), .RN(n4267), .Q(
        \I_cache/cache[7][14] ), .QN(n1436) );
  DFFRX1 \I_cache/cache_reg[0][15]  ( .D(n10044), .CK(clk), .RN(n4267), .Q(
        \I_cache/cache[0][15] ), .QN(n1378) );
  DFFRX1 \I_cache/cache_reg[1][15]  ( .D(n10043), .CK(clk), .RN(n4267), .Q(
        \I_cache/cache[1][15] ), .QN(n455) );
  DFFRX1 \I_cache/cache_reg[2][15]  ( .D(n10042), .CK(clk), .RN(n4267), .Q(
        \I_cache/cache[2][15] ), .QN(n1377) );
  DFFRX1 \I_cache/cache_reg[3][15]  ( .D(n10041), .CK(clk), .RN(n4267), .Q(
        \I_cache/cache[3][15] ), .QN(n454) );
  DFFRX1 \I_cache/cache_reg[4][15]  ( .D(n10040), .CK(clk), .RN(n4267), .Q(
        \I_cache/cache[4][15] ), .QN(n642) );
  DFFRX1 \I_cache/cache_reg[5][15]  ( .D(n10039), .CK(clk), .RN(n4267), .Q(
        \I_cache/cache[5][15] ), .QN(n1561) );
  DFFRX1 \I_cache/cache_reg[6][15]  ( .D(n10038), .CK(clk), .RN(n4267), .Q(
        \I_cache/cache[6][15] ), .QN(n1376) );
  DFFRX1 \I_cache/cache_reg[7][15]  ( .D(n10037), .CK(clk), .RN(n4267), .Q(
        \I_cache/cache[7][15] ), .QN(n453) );
  DFFRX1 \I_cache/cache_reg[0][32]  ( .D(n9908), .CK(clk), .RN(n4278), .Q(
        \I_cache/cache[0][32] ), .QN(n683) );
  DFFRX1 \I_cache/cache_reg[1][32]  ( .D(n9907), .CK(clk), .RN(n4278), .Q(
        \I_cache/cache[1][32] ), .QN(n1609) );
  DFFRX1 \I_cache/cache_reg[2][32]  ( .D(n9906), .CK(clk), .RN(n4278), .Q(
        \I_cache/cache[2][32] ), .QN(n690) );
  DFFRX1 \I_cache/cache_reg[3][32]  ( .D(n9905), .CK(clk), .RN(n4278), .Q(
        \I_cache/cache[3][32] ), .QN(n1611) );
  DFFRX1 \I_cache/cache_reg[4][32]  ( .D(n9904), .CK(clk), .RN(n4279), .Q(
        \I_cache/cache[4][32] ), .QN(n689) );
  DFFRX1 \I_cache/cache_reg[5][32]  ( .D(n9903), .CK(clk), .RN(n4279), .Q(
        \I_cache/cache[5][32] ), .QN(n1610) );
  DFFRX1 \I_cache/cache_reg[6][32]  ( .D(n9902), .CK(clk), .RN(n4279), .Q(
        \I_cache/cache[6][32] ), .QN(n694) );
  DFFRX1 \I_cache/cache_reg[7][32]  ( .D(n9901), .CK(clk), .RN(n4279), .Q(
        \I_cache/cache[7][32] ), .QN(n1615) );
  DFFRX1 \I_cache/cache_reg[0][33]  ( .D(n9900), .CK(clk), .RN(n4279), .Q(
        \I_cache/cache[0][33] ), .QN(n481) );
  DFFRX1 \I_cache/cache_reg[1][33]  ( .D(n9899), .CK(clk), .RN(n4279), .Q(
        \I_cache/cache[1][33] ), .QN(n1396) );
  DFFRX1 \I_cache/cache_reg[2][33]  ( .D(n9898), .CK(clk), .RN(n4279), .Q(
        \I_cache/cache[2][33] ), .QN(n483) );
  DFFRX1 \I_cache/cache_reg[3][33]  ( .D(n9897), .CK(clk), .RN(n4279), .Q(
        \I_cache/cache[3][33] ), .QN(n1398) );
  DFFRX1 \I_cache/cache_reg[4][33]  ( .D(n9896), .CK(clk), .RN(n4279), .Q(
        \I_cache/cache[4][33] ), .QN(n482) );
  DFFRX1 \I_cache/cache_reg[5][33]  ( .D(n9895), .CK(clk), .RN(n4279), .Q(
        \I_cache/cache[5][33] ), .QN(n1397) );
  DFFRX1 \I_cache/cache_reg[6][33]  ( .D(n9894), .CK(clk), .RN(n4279), .Q(
        \I_cache/cache[6][33] ), .QN(n522) );
  DFFRX1 \I_cache/cache_reg[7][33]  ( .D(n9893), .CK(clk), .RN(n4279), .Q(
        \I_cache/cache[7][33] ), .QN(n1440) );
  DFFRX1 \I_cache/cache_reg[0][34]  ( .D(n9892), .CK(clk), .RN(n4280), .Q(
        \I_cache/cache[0][34] ), .QN(n561) );
  DFFRX1 \I_cache/cache_reg[1][34]  ( .D(n9891), .CK(clk), .RN(n4280), .Q(
        \I_cache/cache[1][34] ), .QN(n1480) );
  DFFRX1 \I_cache/cache_reg[2][34]  ( .D(n9890), .CK(clk), .RN(n4280), .Q(
        \I_cache/cache[2][34] ), .QN(n563) );
  DFFRX1 \I_cache/cache_reg[3][34]  ( .D(n9889), .CK(clk), .RN(n4280), .Q(
        \I_cache/cache[3][34] ), .QN(n1482) );
  DFFRX1 \I_cache/cache_reg[4][34]  ( .D(n9888), .CK(clk), .RN(n4280), .Q(
        \I_cache/cache[4][34] ), .QN(n562) );
  DFFRX1 \I_cache/cache_reg[5][34]  ( .D(n9887), .CK(clk), .RN(n4280), .Q(
        \I_cache/cache[5][34] ), .QN(n1481) );
  DFFRX1 \I_cache/cache_reg[6][34]  ( .D(n9886), .CK(clk), .RN(n4280), .Q(
        \I_cache/cache[6][34] ), .QN(n676) );
  DFFRX1 \I_cache/cache_reg[7][34]  ( .D(n9885), .CK(clk), .RN(n4280), .Q(
        \I_cache/cache[7][34] ), .QN(n1595) );
  DFFRX1 \I_cache/cache_reg[0][35]  ( .D(n9884), .CK(clk), .RN(n4280), .Q(
        \I_cache/cache[0][35] ), .QN(n444) );
  DFFRX1 \I_cache/cache_reg[1][35]  ( .D(n9883), .CK(clk), .RN(n4280), .Q(
        \I_cache/cache[1][35] ), .QN(n1359) );
  DFFRX1 \I_cache/cache_reg[2][35]  ( .D(n9882), .CK(clk), .RN(n4280), .Q(
        \I_cache/cache[2][35] ), .QN(n443) );
  DFFRX1 \I_cache/cache_reg[3][35]  ( .D(n9881), .CK(clk), .RN(n4280), .Q(
        \I_cache/cache[3][35] ), .QN(n1358) );
  DFFRX1 \I_cache/cache_reg[4][35]  ( .D(n9880), .CK(clk), .RN(n4281), .Q(
        \I_cache/cache[4][35] ), .QN(n449) );
  DFFRX1 \I_cache/cache_reg[5][35]  ( .D(n9879), .CK(clk), .RN(n4281), .Q(
        \I_cache/cache[5][35] ), .QN(n1363) );
  DFFRX1 \I_cache/cache_reg[6][35]  ( .D(n9878), .CK(clk), .RN(n4281), .Q(
        \I_cache/cache[6][35] ), .QN(n442) );
  DFFRX1 \I_cache/cache_reg[7][35]  ( .D(n9877), .CK(clk), .RN(n4281), .Q(
        \I_cache/cache[7][35] ), .QN(n1357) );
  DFFRX1 \I_cache/cache_reg[0][36]  ( .D(n9876), .CK(clk), .RN(n4281), .Q(
        \I_cache/cache[0][36] ), .QN(n552) );
  DFFRX1 \I_cache/cache_reg[1][36]  ( .D(n9875), .CK(clk), .RN(n4281), .Q(
        \I_cache/cache[1][36] ), .QN(n1471) );
  DFFRX1 \I_cache/cache_reg[2][36]  ( .D(n9874), .CK(clk), .RN(n4281), .Q(
        \I_cache/cache[2][36] ), .QN(n551) );
  DFFRX1 \I_cache/cache_reg[3][36]  ( .D(n9873), .CK(clk), .RN(n4281), .Q(
        \I_cache/cache[3][36] ), .QN(n1470) );
  DFFRX1 \I_cache/cache_reg[4][36]  ( .D(n9872), .CK(clk), .RN(n4281), .Q(
        \I_cache/cache[4][36] ), .QN(n645) );
  DFFRX1 \I_cache/cache_reg[5][36]  ( .D(n9871), .CK(clk), .RN(n4281), .Q(
        \I_cache/cache[5][36] ), .QN(n1564) );
  DFFRX1 \I_cache/cache_reg[6][36]  ( .D(n9870), .CK(clk), .RN(n4281), .Q(
        \I_cache/cache[6][36] ), .QN(n550) );
  DFFRX1 \I_cache/cache_reg[7][36]  ( .D(n9869), .CK(clk), .RN(n4281), .Q(
        \I_cache/cache[7][36] ), .QN(n1469) );
  DFFRX1 \I_cache/cache_reg[0][37]  ( .D(n9868), .CK(clk), .RN(n4282), .Q(
        \I_cache/cache[0][37] ), .QN(n572) );
  DFFRX1 \I_cache/cache_reg[1][37]  ( .D(n9867), .CK(clk), .RN(n4282), .Q(
        \I_cache/cache[1][37] ), .QN(n1491) );
  DFFRX1 \I_cache/cache_reg[2][37]  ( .D(n9866), .CK(clk), .RN(n4282), .Q(
        \I_cache/cache[2][37] ), .QN(n571) );
  DFFRX1 \I_cache/cache_reg[3][37]  ( .D(n9865), .CK(clk), .RN(n4282), .Q(
        \I_cache/cache[3][37] ), .QN(n1490) );
  DFFRX1 \I_cache/cache_reg[4][37]  ( .D(n9864), .CK(clk), .RN(n4282), .Q(
        \I_cache/cache[4][37] ), .QN(n653) );
  DFFRX1 \I_cache/cache_reg[5][37]  ( .D(n9863), .CK(clk), .RN(n4282), .Q(
        \I_cache/cache[5][37] ), .QN(n1572) );
  DFFRX1 \I_cache/cache_reg[6][37]  ( .D(n9862), .CK(clk), .RN(n4282), .Q(
        \I_cache/cache[6][37] ), .QN(n570) );
  DFFRX1 \I_cache/cache_reg[7][37]  ( .D(n9861), .CK(clk), .RN(n4282), .Q(
        \I_cache/cache[7][37] ), .QN(n1489) );
  DFFRX1 \I_cache/cache_reg[0][38]  ( .D(n9860), .CK(clk), .RN(n4282), .Q(
        \I_cache/cache[0][38] ), .QN(n499) );
  DFFRX1 \I_cache/cache_reg[1][38]  ( .D(n9859), .CK(clk), .RN(n4282), .Q(
        \I_cache/cache[1][38] ), .QN(n1417) );
  DFFRX1 \I_cache/cache_reg[2][38]  ( .D(n9858), .CK(clk), .RN(n4282), .Q(
        \I_cache/cache[2][38] ), .QN(n498) );
  DFFRX1 \I_cache/cache_reg[3][38]  ( .D(n9857), .CK(clk), .RN(n4282), .Q(
        \I_cache/cache[3][38] ), .QN(n1416) );
  DFFRX1 \I_cache/cache_reg[4][38]  ( .D(n9856), .CK(clk), .RN(n4283), .Q(
        \I_cache/cache[4][38] ), .QN(n646) );
  DFFRX1 \I_cache/cache_reg[5][38]  ( .D(n9855), .CK(clk), .RN(n4283), .Q(
        \I_cache/cache[5][38] ), .QN(n1565) );
  DFFRX1 \I_cache/cache_reg[6][38]  ( .D(n9854), .CK(clk), .RN(n4283), .Q(
        \I_cache/cache[6][38] ), .QN(n497) );
  DFFRX1 \I_cache/cache_reg[7][38]  ( .D(n9853), .CK(clk), .RN(n4283), .Q(
        \I_cache/cache[7][38] ), .QN(n1415) );
  DFFRX1 \I_cache/cache_reg[0][39]  ( .D(n9852), .CK(clk), .RN(n4283), .Q(
        \I_cache/cache[0][39] ), .QN(n614) );
  DFFRX1 \I_cache/cache_reg[1][39]  ( .D(n9851), .CK(clk), .RN(n4283), .Q(
        \I_cache/cache[1][39] ), .QN(n1533) );
  DFFRX1 \I_cache/cache_reg[2][39]  ( .D(n9850), .CK(clk), .RN(n4283), .Q(
        \I_cache/cache[2][39] ), .QN(n613) );
  DFFRX1 \I_cache/cache_reg[3][39]  ( .D(n9849), .CK(clk), .RN(n4283), .Q(
        \I_cache/cache[3][39] ), .QN(n1532) );
  DFFRX1 \I_cache/cache_reg[4][39]  ( .D(n9848), .CK(clk), .RN(n4283), .Q(
        \I_cache/cache[4][39] ), .QN(n665) );
  DFFRX1 \I_cache/cache_reg[5][39]  ( .D(n9847), .CK(clk), .RN(n4283), .Q(
        \I_cache/cache[5][39] ), .QN(n1584) );
  DFFRX1 \I_cache/cache_reg[6][39]  ( .D(n9846), .CK(clk), .RN(n4283), .Q(
        \I_cache/cache[6][39] ), .QN(n612) );
  DFFRX1 \I_cache/cache_reg[7][39]  ( .D(n9845), .CK(clk), .RN(n4283), .Q(
        \I_cache/cache[7][39] ), .QN(n1531) );
  DFFRX1 \I_cache/cache_reg[0][40]  ( .D(n9844), .CK(clk), .RN(n4284), .Q(
        \I_cache/cache[0][40] ), .QN(n610) );
  DFFRX1 \I_cache/cache_reg[1][40]  ( .D(n9843), .CK(clk), .RN(n4284), .Q(
        \I_cache/cache[1][40] ), .QN(n1529) );
  DFFRX1 \I_cache/cache_reg[2][40]  ( .D(n9842), .CK(clk), .RN(n4284), .Q(
        \I_cache/cache[2][40] ), .QN(n609) );
  DFFRX1 \I_cache/cache_reg[3][40]  ( .D(n9841), .CK(clk), .RN(n4284), .Q(
        \I_cache/cache[3][40] ), .QN(n1528) );
  DFFRX1 \I_cache/cache_reg[4][40]  ( .D(n9840), .CK(clk), .RN(n4284), .Q(
        \I_cache/cache[4][40] ), .QN(n661) );
  DFFRX1 \I_cache/cache_reg[5][40]  ( .D(n9839), .CK(clk), .RN(n4284), .Q(
        \I_cache/cache[5][40] ), .QN(n1580) );
  DFFRX1 \I_cache/cache_reg[6][40]  ( .D(n9838), .CK(clk), .RN(n4284), .Q(
        \I_cache/cache[6][40] ), .QN(n611) );
  DFFRX1 \I_cache/cache_reg[7][40]  ( .D(n9837), .CK(clk), .RN(n4284), .Q(
        \I_cache/cache[7][40] ), .QN(n1530) );
  DFFRX1 \I_cache/cache_reg[0][41]  ( .D(n9836), .CK(clk), .RN(n4284), .Q(
        \I_cache/cache[0][41] ), .QN(n508) );
  DFFRX1 \I_cache/cache_reg[1][41]  ( .D(n9835), .CK(clk), .RN(n4284), .Q(
        \I_cache/cache[1][41] ), .QN(n1426) );
  DFFRX1 \I_cache/cache_reg[2][41]  ( .D(n9834), .CK(clk), .RN(n4284), .Q(
        \I_cache/cache[2][41] ), .QN(n507) );
  DFFRX1 \I_cache/cache_reg[3][41]  ( .D(n9833), .CK(clk), .RN(n4284), .Q(
        \I_cache/cache[3][41] ), .QN(n1425) );
  DFFRX1 \I_cache/cache_reg[4][41]  ( .D(n9832), .CK(clk), .RN(n4285), .Q(
        \I_cache/cache[4][41] ), .QN(n664) );
  DFFRX1 \I_cache/cache_reg[5][41]  ( .D(n9831), .CK(clk), .RN(n4285), .Q(
        \I_cache/cache[5][41] ), .QN(n1583) );
  DFFRX1 \I_cache/cache_reg[6][41]  ( .D(n9830), .CK(clk), .RN(n4285), .Q(
        \I_cache/cache[6][41] ), .QN(n509) );
  DFFRX1 \I_cache/cache_reg[7][41]  ( .D(n9829), .CK(clk), .RN(n4285), .Q(
        \I_cache/cache[7][41] ), .QN(n1427) );
  DFFRX1 \I_cache/cache_reg[1][42]  ( .D(n9827), .CK(clk), .RN(n4285), .Q(
        \I_cache/cache[1][42] ), .QN(n1548) );
  DFFRX1 \I_cache/cache_reg[3][42]  ( .D(n9825), .CK(clk), .RN(n4285), .Q(
        \I_cache/cache[3][42] ), .QN(n1547) );
  DFFRX1 \I_cache/cache_reg[5][42]  ( .D(n9823), .CK(clk), .RN(n4285), .Q(
        \I_cache/cache[5][42] ), .QN(n1588) );
  DFFRX1 \I_cache/cache_reg[6][42]  ( .D(n9822), .CK(clk), .RN(n4285), .Q(
        \I_cache/cache[6][42] ), .QN(n627) );
  DFFRX1 \I_cache/cache_reg[7][42]  ( .D(n9821), .CK(clk), .RN(n4285), .Q(
        \I_cache/cache[7][42] ), .QN(n1546) );
  DFFRX1 \I_cache/cache_reg[0][43]  ( .D(n9820), .CK(clk), .RN(n4286), .Q(
        \I_cache/cache[0][43] ), .QN(n636) );
  DFFRX1 \I_cache/cache_reg[1][43]  ( .D(n9819), .CK(clk), .RN(n4286), .Q(
        \I_cache/cache[1][43] ), .QN(n1555) );
  DFFRX1 \I_cache/cache_reg[2][43]  ( .D(n9818), .CK(clk), .RN(n4286), .Q(
        \I_cache/cache[2][43] ), .QN(n635) );
  DFFRX1 \I_cache/cache_reg[3][43]  ( .D(n9817), .CK(clk), .RN(n4286), .Q(
        \I_cache/cache[3][43] ), .QN(n1554) );
  DFFRX1 \I_cache/cache_reg[4][43]  ( .D(n9816), .CK(clk), .RN(n4286), .Q(
        \I_cache/cache[4][43] ), .QN(n672) );
  DFFRX1 \I_cache/cache_reg[5][43]  ( .D(n9815), .CK(clk), .RN(n4286), .Q(
        \I_cache/cache[5][43] ), .QN(n1591) );
  DFFRX1 \I_cache/cache_reg[6][43]  ( .D(n9814), .CK(clk), .RN(n4286), .Q(
        \I_cache/cache[6][43] ), .QN(n634) );
  DFFRX1 \I_cache/cache_reg[7][43]  ( .D(n9813), .CK(clk), .RN(n4286), .Q(
        \I_cache/cache[7][43] ), .QN(n1553) );
  DFFRX1 \I_cache/cache_reg[0][44]  ( .D(n9812), .CK(clk), .RN(n4286), .Q(
        \I_cache/cache[0][44] ), .QN(n517) );
  DFFRX1 \I_cache/cache_reg[1][44]  ( .D(n9811), .CK(clk), .RN(n4286), .Q(
        \I_cache/cache[1][44] ), .QN(n1435) );
  DFFRX1 \I_cache/cache_reg[2][44]  ( .D(n9810), .CK(clk), .RN(n4286), .Q(
        \I_cache/cache[2][44] ), .QN(n515) );
  DFFRX1 \I_cache/cache_reg[3][44]  ( .D(n9809), .CK(clk), .RN(n4286), .Q(
        \I_cache/cache[3][44] ), .QN(n1433) );
  DFFRX1 \I_cache/cache_reg[4][44]  ( .D(n9808), .CK(clk), .RN(n4287), .Q(
        \I_cache/cache[4][44] ), .QN(n658) );
  DFFRX1 \I_cache/cache_reg[5][44]  ( .D(n9807), .CK(clk), .RN(n4287), .Q(
        \I_cache/cache[5][44] ), .QN(n1577) );
  DFFRX1 \I_cache/cache_reg[6][44]  ( .D(n9806), .CK(clk), .RN(n4287), .Q(
        \I_cache/cache[6][44] ), .QN(n516) );
  DFFRX1 \I_cache/cache_reg[7][44]  ( .D(n9805), .CK(clk), .RN(n4287), .Q(
        \I_cache/cache[7][44] ), .QN(n1434) );
  DFFRX1 \I_cache/cache_reg[0][45]  ( .D(n9804), .CK(clk), .RN(n4287), .Q(
        \I_cache/cache[0][45] ), .QN(n593) );
  DFFRX1 \I_cache/cache_reg[1][45]  ( .D(n9803), .CK(clk), .RN(n4287), .Q(
        \I_cache/cache[1][45] ), .QN(n1512) );
  DFFRX1 \I_cache/cache_reg[2][45]  ( .D(n9802), .CK(clk), .RN(n4287), .Q(
        \I_cache/cache[2][45] ), .QN(n592) );
  DFFRX1 \I_cache/cache_reg[3][45]  ( .D(n9801), .CK(clk), .RN(n4287), .Q(
        \I_cache/cache[3][45] ), .QN(n1511) );
  DFFRX1 \I_cache/cache_reg[4][45]  ( .D(n9800), .CK(clk), .RN(n4287), .Q(
        \I_cache/cache[4][45] ), .QN(n656) );
  DFFRX1 \I_cache/cache_reg[5][45]  ( .D(n9799), .CK(clk), .RN(n4287), .Q(
        \I_cache/cache[5][45] ), .QN(n1575) );
  DFFRX1 \I_cache/cache_reg[6][45]  ( .D(n9798), .CK(clk), .RN(n4287), .Q(
        \I_cache/cache[6][45] ), .QN(n591) );
  DFFRX1 \I_cache/cache_reg[7][45]  ( .D(n9797), .CK(clk), .RN(n4287), .Q(
        \I_cache/cache[7][45] ), .QN(n1510) );
  DFFRX1 \I_cache/cache_reg[1][46]  ( .D(n9795), .CK(clk), .RN(n4288), .Q(
        \I_cache/cache[1][46] ), .QN(n1515) );
  DFFRX1 \I_cache/cache_reg[2][46]  ( .D(n9794), .CK(clk), .RN(n4288), .Q(
        \I_cache/cache[2][46] ), .QN(n595) );
  DFFRX1 \I_cache/cache_reg[3][46]  ( .D(n9793), .CK(clk), .RN(n4288), .Q(
        \I_cache/cache[3][46] ), .QN(n1514) );
  DFFRX1 \I_cache/cache_reg[4][46]  ( .D(n9792), .CK(clk), .RN(n4288), .Q(
        \I_cache/cache[4][46] ), .QN(n652) );
  DFFRX1 \I_cache/cache_reg[5][46]  ( .D(n9791), .CK(clk), .RN(n4288), .Q(
        \I_cache/cache[5][46] ), .QN(n1571) );
  DFFRX1 \I_cache/cache_reg[6][46]  ( .D(n9790), .CK(clk), .RN(n4288), .Q(
        \I_cache/cache[6][46] ), .QN(n594) );
  DFFRX1 \I_cache/cache_reg[7][46]  ( .D(n9789), .CK(clk), .RN(n4288), .Q(
        \I_cache/cache[7][46] ), .QN(n1513) );
  DFFRX1 \I_cache/cache_reg[0][47]  ( .D(n9788), .CK(clk), .RN(n4288), .Q(
        \I_cache/cache[0][47] ), .QN(n1375) );
  DFFRX1 \I_cache/cache_reg[1][47]  ( .D(n9787), .CK(clk), .RN(n4288), .Q(
        \I_cache/cache[1][47] ), .QN(n452) );
  DFFRX1 \I_cache/cache_reg[2][47]  ( .D(n9786), .CK(clk), .RN(n4288), .Q(
        \I_cache/cache[2][47] ), .QN(n1374) );
  DFFRX1 \I_cache/cache_reg[3][47]  ( .D(n9785), .CK(clk), .RN(n4288), .Q(
        \I_cache/cache[3][47] ), .QN(n451) );
  DFFRX1 \I_cache/cache_reg[4][47]  ( .D(n9784), .CK(clk), .RN(n4289), .Q(
        \I_cache/cache[4][47] ), .QN(n1373) );
  DFFRX1 \I_cache/cache_reg[5][47]  ( .D(n9783), .CK(clk), .RN(n4289), .Q(
        \I_cache/cache[5][47] ), .QN(n447) );
  DFFRX1 \I_cache/cache_reg[6][47]  ( .D(n9782), .CK(clk), .RN(n4289), .Q(
        \I_cache/cache[6][47] ), .QN(n445) );
  DFFRX1 \I_cache/cache_reg[7][47]  ( .D(n9781), .CK(clk), .RN(n4289), .Q(
        \I_cache/cache[7][47] ), .QN(n1360) );
  DFFRX1 \I_cache/cache_reg[0][64]  ( .D(n9652), .CK(clk), .RN(n4300), .Q(
        \I_cache/cache[0][64] ), .QN(n682) );
  DFFRX1 \I_cache/cache_reg[1][64]  ( .D(n9651), .CK(clk), .RN(n4300), .Q(
        \I_cache/cache[1][64] ), .QN(n1606) );
  DFFRX1 \I_cache/cache_reg[2][64]  ( .D(n9650), .CK(clk), .RN(n4300), .Q(
        \I_cache/cache[2][64] ), .QN(n688) );
  DFFRX1 \I_cache/cache_reg[3][64]  ( .D(n9649), .CK(clk), .RN(n4300), .Q(
        \I_cache/cache[3][64] ), .QN(n1608) );
  DFFRX1 \I_cache/cache_reg[4][64]  ( .D(n9648), .CK(clk), .RN(n4300), .Q(
        \I_cache/cache[4][64] ), .QN(n687) );
  DFFRX1 \I_cache/cache_reg[5][64]  ( .D(n9647), .CK(clk), .RN(n4300), .Q(
        \I_cache/cache[5][64] ), .QN(n1607) );
  DFFRX1 \I_cache/cache_reg[6][64]  ( .D(n9646), .CK(clk), .RN(n4300), .Q(
        \I_cache/cache[6][64] ), .QN(n693) );
  DFFRX1 \I_cache/cache_reg[7][64]  ( .D(n9645), .CK(clk), .RN(n4300), .Q(
        \I_cache/cache[7][64] ), .QN(n1614) );
  DFFRX1 \I_cache/cache_reg[0][65]  ( .D(n9644), .CK(clk), .RN(n4300), .Q(
        \I_cache/cache[0][65] ), .QN(n478) );
  DFFRX1 \I_cache/cache_reg[1][65]  ( .D(n9643), .CK(clk), .RN(n4300), .Q(
        \I_cache/cache[1][65] ), .QN(n1393) );
  DFFRX1 \I_cache/cache_reg[2][65]  ( .D(n9642), .CK(clk), .RN(n4300), .Q(
        \I_cache/cache[2][65] ), .QN(n480) );
  DFFRX1 \I_cache/cache_reg[3][65]  ( .D(n9641), .CK(clk), .RN(n4300), .Q(
        \I_cache/cache[3][65] ), .QN(n1395) );
  DFFRX1 \I_cache/cache_reg[4][65]  ( .D(n9640), .CK(clk), .RN(n4301), .Q(
        \I_cache/cache[4][65] ), .QN(n479) );
  DFFRX1 \I_cache/cache_reg[5][65]  ( .D(n9639), .CK(clk), .RN(n4301), .Q(
        \I_cache/cache[5][65] ), .QN(n1394) );
  DFFRX1 \I_cache/cache_reg[6][65]  ( .D(n9638), .CK(clk), .RN(n4301), .Q(
        \I_cache/cache[6][65] ), .QN(n521) );
  DFFRX1 \I_cache/cache_reg[7][65]  ( .D(n9637), .CK(clk), .RN(n4301), .Q(
        \I_cache/cache[7][65] ), .QN(n1439) );
  DFFRX1 \I_cache/cache_reg[0][66]  ( .D(n9636), .CK(clk), .RN(n4301), .Q(
        \I_cache/cache[0][66] ), .QN(n553) );
  DFFRX1 \I_cache/cache_reg[1][66]  ( .D(n9635), .CK(clk), .RN(n4301), .Q(
        \I_cache/cache[1][66] ), .QN(n1472) );
  DFFRX1 \I_cache/cache_reg[2][66]  ( .D(n9634), .CK(clk), .RN(n4301), .Q(
        \I_cache/cache[2][66] ), .QN(n555) );
  DFFRX1 \I_cache/cache_reg[3][66]  ( .D(n9633), .CK(clk), .RN(n4301), .Q(
        \I_cache/cache[3][66] ), .QN(n1474) );
  DFFRX1 \I_cache/cache_reg[4][66]  ( .D(n9632), .CK(clk), .RN(n4301), .Q(
        \I_cache/cache[4][66] ), .QN(n554) );
  DFFRX1 \I_cache/cache_reg[5][66]  ( .D(n9631), .CK(clk), .RN(n4301), .Q(
        \I_cache/cache[5][66] ), .QN(n1473) );
  DFFRX1 \I_cache/cache_reg[6][66]  ( .D(n9630), .CK(clk), .RN(n4301), .Q(
        \I_cache/cache[6][66] ), .QN(n674) );
  DFFRX1 \I_cache/cache_reg[7][66]  ( .D(n9629), .CK(clk), .RN(n4301), .Q(
        \I_cache/cache[7][66] ), .QN(n1593) );
  DFFRX1 \I_cache/cache_reg[0][67]  ( .D(n9628), .CK(clk), .RN(n4302), .Q(
        \I_cache/cache[0][67] ), .QN(n441) );
  DFFRX1 \I_cache/cache_reg[1][67]  ( .D(n9627), .CK(clk), .RN(n4302), .Q(
        \I_cache/cache[1][67] ), .QN(n1356) );
  DFFRX1 \I_cache/cache_reg[2][67]  ( .D(n9626), .CK(clk), .RN(n4302), .Q(
        \I_cache/cache[2][67] ), .QN(n440) );
  DFFRX1 \I_cache/cache_reg[3][67]  ( .D(n9625), .CK(clk), .RN(n4302), .Q(
        \I_cache/cache[3][67] ), .QN(n1355) );
  DFFRX1 \I_cache/cache_reg[4][67]  ( .D(n9624), .CK(clk), .RN(n4302), .Q(
        \I_cache/cache[4][67] ), .QN(n525) );
  DFFRX1 \I_cache/cache_reg[5][67]  ( .D(n9623), .CK(clk), .RN(n4302), .Q(
        \I_cache/cache[5][67] ), .QN(n1443) );
  DFFRX1 \I_cache/cache_reg[6][67]  ( .D(n9622), .CK(clk), .RN(n4302), .Q(
        \I_cache/cache[6][67] ), .QN(n439) );
  DFFRX1 \I_cache/cache_reg[7][67]  ( .D(n9621), .CK(clk), .RN(n4302), .Q(
        \I_cache/cache[7][67] ), .QN(n1354) );
  DFFRX1 \I_cache/cache_reg[0][68]  ( .D(n9620), .CK(clk), .RN(n4302), .Q(
        \I_cache/cache[0][68] ), .QN(n549) );
  DFFRX1 \I_cache/cache_reg[1][68]  ( .D(n9619), .CK(clk), .RN(n4302), .Q(
        \I_cache/cache[1][68] ), .QN(n1468) );
  DFFRX1 \I_cache/cache_reg[2][68]  ( .D(n9618), .CK(clk), .RN(n4302), .Q(
        \I_cache/cache[2][68] ), .QN(n548) );
  DFFRX1 \I_cache/cache_reg[3][68]  ( .D(n9617), .CK(clk), .RN(n4302), .Q(
        \I_cache/cache[3][68] ), .QN(n1467) );
  DFFRX1 \I_cache/cache_reg[4][68]  ( .D(n9616), .CK(clk), .RN(n4303), .Q(
        \I_cache/cache[4][68] ), .QN(n643) );
  DFFRX1 \I_cache/cache_reg[5][68]  ( .D(n9615), .CK(clk), .RN(n4303), .Q(
        \I_cache/cache[5][68] ), .QN(n1562) );
  DFFRX1 \I_cache/cache_reg[6][68]  ( .D(n9614), .CK(clk), .RN(n4303), .Q(
        \I_cache/cache[6][68] ), .QN(n547) );
  DFFRX1 \I_cache/cache_reg[7][68]  ( .D(n9613), .CK(clk), .RN(n4303), .Q(
        \I_cache/cache[7][68] ), .QN(n1466) );
  DFFRX1 \I_cache/cache_reg[0][69]  ( .D(n9612), .CK(clk), .RN(n4303), .Q(
        \I_cache/cache[0][69] ), .QN(n491) );
  DFFRX1 \I_cache/cache_reg[1][69]  ( .D(n9611), .CK(clk), .RN(n4303), .Q(
        \I_cache/cache[1][69] ), .QN(n1409) );
  DFFRX1 \I_cache/cache_reg[2][69]  ( .D(n9610), .CK(clk), .RN(n4303), .Q(
        \I_cache/cache[2][69] ), .QN(n490) );
  DFFRX1 \I_cache/cache_reg[3][69]  ( .D(n9609), .CK(clk), .RN(n4303), .Q(
        \I_cache/cache[3][69] ), .QN(n1408) );
  DFFRX1 \I_cache/cache_reg[4][69]  ( .D(n9608), .CK(clk), .RN(n4303), .Q(
        \I_cache/cache[4][69] ), .QN(n526) );
  DFFRX1 \I_cache/cache_reg[5][69]  ( .D(n9607), .CK(clk), .RN(n4303), .Q(
        \I_cache/cache[5][69] ), .QN(n1445) );
  DFFRX1 \I_cache/cache_reg[6][69]  ( .D(n9606), .CK(clk), .RN(n4303), .Q(
        \I_cache/cache[6][69] ), .QN(n489) );
  DFFRX1 \I_cache/cache_reg[7][69]  ( .D(n9605), .CK(clk), .RN(n4303), .Q(
        \I_cache/cache[7][69] ), .QN(n1407) );
  DFFRX1 \I_cache/cache_reg[0][70]  ( .D(n9604), .CK(clk), .RN(n4304), .Q(
        \I_cache/cache[0][70] ), .QN(n496) );
  DFFRX1 \I_cache/cache_reg[1][70]  ( .D(n9603), .CK(clk), .RN(n4304), .Q(
        \I_cache/cache[1][70] ), .QN(n1414) );
  DFFRX1 \I_cache/cache_reg[2][70]  ( .D(n9602), .CK(clk), .RN(n4304), .Q(
        \I_cache/cache[2][70] ), .QN(n495) );
  DFFRX1 \I_cache/cache_reg[3][70]  ( .D(n9601), .CK(clk), .RN(n4304), .Q(
        \I_cache/cache[3][70] ), .QN(n1413) );
  DFFRX1 \I_cache/cache_reg[4][70]  ( .D(n9600), .CK(clk), .RN(n4304), .Q(
        \I_cache/cache[4][70] ), .QN(n528) );
  DFFRX1 \I_cache/cache_reg[5][70]  ( .D(n9599), .CK(clk), .RN(n4304), .Q(
        \I_cache/cache[5][70] ), .QN(n1447) );
  DFFRX1 \I_cache/cache_reg[6][70]  ( .D(n9598), .CK(clk), .RN(n4304), .Q(
        \I_cache/cache[6][70] ), .QN(n494) );
  DFFRX1 \I_cache/cache_reg[7][70]  ( .D(n9597), .CK(clk), .RN(n4304), .Q(
        \I_cache/cache[7][70] ), .QN(n1412) );
  DFFRX1 \I_cache/cache_reg[0][71]  ( .D(n9596), .CK(clk), .RN(n4304), .Q(
        \I_cache/cache[0][71] ), .QN(n542) );
  DFFRX1 \I_cache/cache_reg[1][71]  ( .D(n9595), .CK(clk), .RN(n4304), .Q(
        \I_cache/cache[1][71] ), .QN(n1461) );
  DFFRX1 \I_cache/cache_reg[2][71]  ( .D(n9594), .CK(clk), .RN(n4304), .Q(
        \I_cache/cache[2][71] ), .QN(n541) );
  DFFRX1 \I_cache/cache_reg[3][71]  ( .D(n9593), .CK(clk), .RN(n4304), .Q(
        \I_cache/cache[3][71] ), .QN(n1460) );
  DFFRX1 \I_cache/cache_reg[4][71]  ( .D(n9592), .CK(clk), .RN(n4305), .Q(
        \I_cache/cache[4][71] ), .QN(n662) );
  DFFRX1 \I_cache/cache_reg[5][71]  ( .D(n9591), .CK(clk), .RN(n4305), .Q(
        \I_cache/cache[5][71] ), .QN(n1581) );
  DFFRX1 \I_cache/cache_reg[6][71]  ( .D(n9590), .CK(clk), .RN(n4305), .Q(
        \I_cache/cache[6][71] ), .QN(n543) );
  DFFRX1 \I_cache/cache_reg[7][71]  ( .D(n9589), .CK(clk), .RN(n4305), .Q(
        \I_cache/cache[7][71] ), .QN(n1462) );
  DFFRX1 \I_cache/cache_reg[0][72]  ( .D(n9588), .CK(clk), .RN(n4305), .Q(
        \I_cache/cache[0][72] ), .QN(n462) );
  DFFRX1 \I_cache/cache_reg[1][72]  ( .D(n9587), .CK(clk), .RN(n4305), .Q(
        \I_cache/cache[1][72] ), .QN(n1371) );
  DFFRX1 \I_cache/cache_reg[2][72]  ( .D(n9586), .CK(clk), .RN(n4305), .Q(
        \I_cache/cache[2][72] ), .QN(n503) );
  DFFRX1 \I_cache/cache_reg[3][72]  ( .D(n9585), .CK(clk), .RN(n4305), .Q(
        \I_cache/cache[3][72] ), .QN(n1421) );
  DFFRX1 \I_cache/cache_reg[4][72]  ( .D(n9584), .CK(clk), .RN(n4305), .Q(
        \I_cache/cache[4][72] ), .QN(n529) );
  DFFRX1 \I_cache/cache_reg[5][72]  ( .D(n9583), .CK(clk), .RN(n4305), .Q(
        \I_cache/cache[5][72] ), .QN(n1448) );
  DFFRX1 \I_cache/cache_reg[6][72]  ( .D(n9582), .CK(clk), .RN(n4305), .Q(
        \I_cache/cache[6][72] ), .QN(n504) );
  DFFRX1 \I_cache/cache_reg[7][72]  ( .D(n9581), .CK(clk), .RN(n4305), .Q(
        \I_cache/cache[7][72] ), .QN(n1422) );
  DFFRX1 \I_cache/cache_reg[0][73]  ( .D(n9580), .CK(clk), .RN(n4306), .Q(
        \I_cache/cache[0][73] ), .QN(n607) );
  DFFRX1 \I_cache/cache_reg[1][73]  ( .D(n9579), .CK(clk), .RN(n4306), .Q(
        \I_cache/cache[1][73] ), .QN(n1526) );
  DFFRX1 \I_cache/cache_reg[2][73]  ( .D(n9578), .CK(clk), .RN(n4306), .Q(
        \I_cache/cache[2][73] ), .QN(n606) );
  DFFRX1 \I_cache/cache_reg[3][73]  ( .D(n9577), .CK(clk), .RN(n4306), .Q(
        \I_cache/cache[3][73] ), .QN(n1525) );
  DFFRX1 \I_cache/cache_reg[4][73]  ( .D(n9576), .CK(clk), .RN(n4306), .Q(
        \I_cache/cache[4][73] ), .QN(n660) );
  DFFRX1 \I_cache/cache_reg[5][73]  ( .D(n9575), .CK(clk), .RN(n4306), .Q(
        \I_cache/cache[5][73] ), .QN(n1579) );
  DFFRX1 \I_cache/cache_reg[6][73]  ( .D(n9574), .CK(clk), .RN(n4306), .Q(
        \I_cache/cache[6][73] ), .QN(n608) );
  DFFRX1 \I_cache/cache_reg[7][73]  ( .D(n9573), .CK(clk), .RN(n4306), .Q(
        \I_cache/cache[7][73] ), .QN(n1527) );
  DFFRX1 \I_cache/cache_reg[1][74]  ( .D(n9571), .CK(clk), .RN(n4306), .Q(
        \I_cache/cache[1][74] ), .QN(n1542) );
  DFFRX1 \I_cache/cache_reg[2][74]  ( .D(n9570), .CK(clk), .RN(n4306), .Q(
        \I_cache/cache[2][74] ), .QN(n622) );
  DFFRX1 \I_cache/cache_reg[3][74]  ( .D(n9569), .CK(clk), .RN(n4306), .Q(
        \I_cache/cache[3][74] ), .QN(n1541) );
  DFFRX1 \I_cache/cache_reg[4][74]  ( .D(n9568), .CK(clk), .RN(n4307), .Q(
        \I_cache/cache[4][74] ), .QN(n667) );
  DFFRX1 \I_cache/cache_reg[5][74]  ( .D(n9567), .CK(clk), .RN(n4307), .Q(
        \I_cache/cache[5][74] ), .QN(n1586) );
  DFFRX1 \I_cache/cache_reg[6][74]  ( .D(n9566), .CK(clk), .RN(n4307), .Q(
        \I_cache/cache[6][74] ), .QN(n621) );
  DFFRX1 \I_cache/cache_reg[7][74]  ( .D(n9565), .CK(clk), .RN(n4307), .Q(
        \I_cache/cache[7][74] ), .QN(n1540) );
  DFFRX1 \I_cache/cache_reg[0][75]  ( .D(n9564), .CK(clk), .RN(n4307), .Q(
        \I_cache/cache[0][75] ), .QN(n633) );
  DFFRX1 \I_cache/cache_reg[1][75]  ( .D(n9563), .CK(clk), .RN(n4307), .Q(
        \I_cache/cache[1][75] ), .QN(n1552) );
  DFFRX1 \I_cache/cache_reg[2][75]  ( .D(n9562), .CK(clk), .RN(n4307), .Q(
        \I_cache/cache[2][75] ), .QN(n539) );
  DFFRX1 \I_cache/cache_reg[3][75]  ( .D(n9561), .CK(clk), .RN(n4307), .Q(
        \I_cache/cache[3][75] ), .QN(n1458) );
  DFFRX1 \I_cache/cache_reg[4][75]  ( .D(n9560), .CK(clk), .RN(n4307), .Q(
        \I_cache/cache[4][75] ), .QN(n671) );
  DFFRX1 \I_cache/cache_reg[5][75]  ( .D(n9559), .CK(clk), .RN(n4307), .Q(
        \I_cache/cache[5][75] ), .QN(n1590) );
  DFFRX1 \I_cache/cache_reg[6][75]  ( .D(n9558), .CK(clk), .RN(n4307), .Q(
        \I_cache/cache[6][75] ), .QN(n540) );
  DFFRX1 \I_cache/cache_reg[7][75]  ( .D(n9557), .CK(clk), .RN(n4307), .Q(
        \I_cache/cache[7][75] ), .QN(n1459) );
  DFFRX1 \I_cache/cache_reg[0][76]  ( .D(n9556), .CK(clk), .RN(n4308), .Q(
        \I_cache/cache[0][76] ), .QN(n514) );
  DFFRX1 \I_cache/cache_reg[1][76]  ( .D(n9555), .CK(clk), .RN(n4308), .Q(
        \I_cache/cache[1][76] ), .QN(n1432) );
  DFFRX1 \I_cache/cache_reg[2][76]  ( .D(n9554), .CK(clk), .RN(n4308), .Q(
        \I_cache/cache[2][76] ), .QN(n512) );
  DFFRX1 \I_cache/cache_reg[3][76]  ( .D(n9553), .CK(clk), .RN(n4308), .Q(
        \I_cache/cache[3][76] ), .QN(n1430) );
  DFFRX1 \I_cache/cache_reg[4][76]  ( .D(n9552), .CK(clk), .RN(n4308), .Q(
        \I_cache/cache[4][76] ), .QN(n532) );
  DFFRX1 \I_cache/cache_reg[5][76]  ( .D(n9551), .CK(clk), .RN(n4308), .Q(
        \I_cache/cache[5][76] ), .QN(n1451) );
  DFFRX1 \I_cache/cache_reg[6][76]  ( .D(n9550), .CK(clk), .RN(n4308), .Q(
        \I_cache/cache[6][76] ), .QN(n513) );
  DFFRX1 \I_cache/cache_reg[7][76]  ( .D(n9549), .CK(clk), .RN(n4308), .Q(
        \I_cache/cache[7][76] ), .QN(n1431) );
  DFFRX1 \I_cache/cache_reg[0][77]  ( .D(n9548), .CK(clk), .RN(n4308), .Q(
        \I_cache/cache[0][77] ), .QN(n581) );
  DFFRX1 \I_cache/cache_reg[1][77]  ( .D(n9547), .CK(clk), .RN(n4308), .Q(
        \I_cache/cache[1][77] ), .QN(n1500) );
  DFFRX1 \I_cache/cache_reg[2][77]  ( .D(n9546), .CK(clk), .RN(n4308), .Q(
        \I_cache/cache[2][77] ), .QN(n580) );
  DFFRX1 \I_cache/cache_reg[3][77]  ( .D(n9545), .CK(clk), .RN(n4308), .Q(
        \I_cache/cache[3][77] ), .QN(n1499) );
  DFFRX1 \I_cache/cache_reg[4][77]  ( .D(n9544), .CK(clk), .RN(n4309), .Q(
        \I_cache/cache[4][77] ), .QN(n651) );
  DFFRX1 \I_cache/cache_reg[5][77]  ( .D(n9543), .CK(clk), .RN(n4309), .Q(
        \I_cache/cache[5][77] ), .QN(n1570) );
  DFFRX1 \I_cache/cache_reg[6][77]  ( .D(n9542), .CK(clk), .RN(n4309), .Q(
        \I_cache/cache[6][77] ), .QN(n579) );
  DFFRX1 \I_cache/cache_reg[7][77]  ( .D(n9541), .CK(clk), .RN(n4309), .Q(
        \I_cache/cache[7][77] ), .QN(n1498) );
  DFFRX1 \I_cache/cache_reg[0][78]  ( .D(n9540), .CK(clk), .RN(n4309), .Q(
        \I_cache/cache[0][78] ), .QN(n584) );
  DFFRX1 \I_cache/cache_reg[1][78]  ( .D(n9539), .CK(clk), .RN(n4309), .Q(
        \I_cache/cache[1][78] ), .QN(n1503) );
  DFFRX1 \I_cache/cache_reg[2][78]  ( .D(n9538), .CK(clk), .RN(n4309), .Q(
        \I_cache/cache[2][78] ), .QN(n583) );
  DFFRX1 \I_cache/cache_reg[3][78]  ( .D(n9537), .CK(clk), .RN(n4309), .Q(
        \I_cache/cache[3][78] ), .QN(n1502) );
  DFFRX1 \I_cache/cache_reg[4][78]  ( .D(n9536), .CK(clk), .RN(n4309), .Q(
        \I_cache/cache[4][78] ), .QN(n648) );
  DFFRX1 \I_cache/cache_reg[5][78]  ( .D(n9535), .CK(clk), .RN(n4309), .Q(
        \I_cache/cache[5][78] ), .QN(n1567) );
  DFFRX1 \I_cache/cache_reg[6][78]  ( .D(n9534), .CK(clk), .RN(n4309), .Q(
        \I_cache/cache[6][78] ), .QN(n582) );
  DFFRX1 \I_cache/cache_reg[7][78]  ( .D(n9533), .CK(clk), .RN(n4309), .Q(
        \I_cache/cache[7][78] ), .QN(n1501) );
  DFFRX1 \I_cache/cache_reg[0][79]  ( .D(n9532), .CK(clk), .RN(n4310), .Q(
        \I_cache/cache[0][79] ), .QN(n458) );
  DFFRX1 \I_cache/cache_reg[1][79]  ( .D(n9531), .CK(clk), .RN(n4310), .Q(
        \I_cache/cache[1][79] ), .QN(n1367) );
  DFFRX1 \I_cache/cache_reg[2][79]  ( .D(n9530), .CK(clk), .RN(n4310), .Q(
        \I_cache/cache[2][79] ), .QN(n457) );
  DFFRX1 \I_cache/cache_reg[3][79]  ( .D(n9529), .CK(clk), .RN(n4310), .Q(
        \I_cache/cache[3][79] ), .QN(n1366) );
  DFFRX1 \I_cache/cache_reg[4][79]  ( .D(n9528), .CK(clk), .RN(n4310), .Q(
        \I_cache/cache[4][79] ), .QN(n523) );
  DFFRX1 \I_cache/cache_reg[5][79]  ( .D(n9527), .CK(clk), .RN(n4310), .Q(
        \I_cache/cache[5][79] ), .QN(n1441) );
  DFFRX1 \I_cache/cache_reg[6][79]  ( .D(n9526), .CK(clk), .RN(n4310), .Q(
        \I_cache/cache[6][79] ), .QN(n459) );
  DFFRX1 \I_cache/cache_reg[7][79]  ( .D(n9525), .CK(clk), .RN(n4310), .Q(
        \I_cache/cache[7][79] ), .QN(n1368) );
  DFFRX1 \I_cache/cache_reg[0][96]  ( .D(n9396), .CK(clk), .RN(n4321), .Q(
        \I_cache/cache[0][96] ), .QN(n681) );
  DFFRX1 \I_cache/cache_reg[1][96]  ( .D(n9395), .CK(clk), .RN(n4321), .Q(
        \I_cache/cache[1][96] ), .QN(n1603) );
  DFFRX1 \I_cache/cache_reg[2][96]  ( .D(n9394), .CK(clk), .RN(n4321), .Q(
        \I_cache/cache[2][96] ), .QN(n686) );
  DFFRX1 \I_cache/cache_reg[3][96]  ( .D(n9393), .CK(clk), .RN(n4321), .Q(
        \I_cache/cache[3][96] ), .QN(n1605) );
  DFFRX1 \I_cache/cache_reg[4][96]  ( .D(n9392), .CK(clk), .RN(n4321), .Q(
        \I_cache/cache[4][96] ), .QN(n685) );
  DFFRX1 \I_cache/cache_reg[5][96]  ( .D(n9391), .CK(clk), .RN(n4321), .Q(
        \I_cache/cache[5][96] ), .QN(n1604) );
  DFFRX1 \I_cache/cache_reg[6][96]  ( .D(n9390), .CK(clk), .RN(n4321), .Q(
        \I_cache/cache[6][96] ), .QN(n692) );
  DFFRX1 \I_cache/cache_reg[7][96]  ( .D(n9389), .CK(clk), .RN(n4321), .Q(
        \I_cache/cache[7][96] ), .QN(n1613) );
  DFFRX1 \I_cache/cache_reg[0][97]  ( .D(n9388), .CK(clk), .RN(n4322), .Q(
        \I_cache/cache[0][97] ), .QN(n475) );
  DFFRX1 \I_cache/cache_reg[1][97]  ( .D(n9387), .CK(clk), .RN(n4322), .Q(
        \I_cache/cache[1][97] ), .QN(n1390) );
  DFFRX1 \I_cache/cache_reg[2][97]  ( .D(n9386), .CK(clk), .RN(n4322), .Q(
        \I_cache/cache[2][97] ), .QN(n477) );
  DFFRX1 \I_cache/cache_reg[3][97]  ( .D(n9385), .CK(clk), .RN(n4322), .Q(
        \I_cache/cache[3][97] ), .QN(n1392) );
  DFFRX1 \I_cache/cache_reg[4][97]  ( .D(n9384), .CK(clk), .RN(n4322), .Q(
        \I_cache/cache[4][97] ), .QN(n476) );
  DFFRX1 \I_cache/cache_reg[5][97]  ( .D(n9383), .CK(clk), .RN(n4322), .Q(
        \I_cache/cache[5][97] ), .QN(n1391) );
  DFFRX1 \I_cache/cache_reg[6][97]  ( .D(n9382), .CK(clk), .RN(n4322), .Q(
        \I_cache/cache[6][97] ), .QN(n536) );
  DFFRX1 \I_cache/cache_reg[7][97]  ( .D(n9381), .CK(clk), .RN(n4322), .Q(
        \I_cache/cache[7][97] ), .QN(n1455) );
  DFFRX1 \I_cache/cache_reg[0][98]  ( .D(n9380), .CK(clk), .RN(n4322), .Q(
        \I_cache/cache[0][98] ), .QN(n556) );
  DFFRX1 \I_cache/cache_reg[1][98]  ( .D(n9379), .CK(clk), .RN(n4322), .Q(
        \I_cache/cache[1][98] ), .QN(n1475) );
  DFFRX1 \I_cache/cache_reg[2][98]  ( .D(n9378), .CK(clk), .RN(n4322), .Q(
        \I_cache/cache[2][98] ), .QN(n558) );
  DFFRX1 \I_cache/cache_reg[3][98]  ( .D(n9377), .CK(clk), .RN(n4322), .Q(
        \I_cache/cache[3][98] ), .QN(n1477) );
  DFFRX1 \I_cache/cache_reg[4][98]  ( .D(n9376), .CK(clk), .RN(n4323), .Q(
        \I_cache/cache[4][98] ), .QN(n557) );
  DFFRX1 \I_cache/cache_reg[5][98]  ( .D(n9375), .CK(clk), .RN(n4323), .Q(
        \I_cache/cache[5][98] ), .QN(n1476) );
  DFFRX1 \I_cache/cache_reg[6][98]  ( .D(n9374), .CK(clk), .RN(n4323), .Q(
        \I_cache/cache[6][98] ), .QN(n675) );
  DFFRX1 \I_cache/cache_reg[7][98]  ( .D(n9373), .CK(clk), .RN(n4323), .Q(
        \I_cache/cache[7][98] ), .QN(n1594) );
  DFFRX1 \I_cache/cache_reg[0][99]  ( .D(n9372), .CK(clk), .RN(n4323), .Q(
        \I_cache/cache[0][99] ), .QN(n438) );
  DFFRX1 \I_cache/cache_reg[1][99]  ( .D(n9371), .CK(clk), .RN(n4323), .Q(
        \I_cache/cache[1][99] ), .QN(n1353) );
  DFFRX1 \I_cache/cache_reg[2][99]  ( .D(n9370), .CK(clk), .RN(n4323), .Q(
        \I_cache/cache[2][99] ), .QN(n437) );
  DFFRX1 \I_cache/cache_reg[3][99]  ( .D(n9369), .CK(clk), .RN(n4323), .Q(
        \I_cache/cache[3][99] ), .QN(n1352) );
  DFFRX1 \I_cache/cache_reg[4][99]  ( .D(n9368), .CK(clk), .RN(n4323), .Q(
        \I_cache/cache[4][99] ), .QN(n450) );
  DFFRX1 \I_cache/cache_reg[5][99]  ( .D(n9367), .CK(clk), .RN(n4323), .Q(
        \I_cache/cache[5][99] ), .QN(n1364) );
  DFFRX1 \I_cache/cache_reg[6][99]  ( .D(n9366), .CK(clk), .RN(n4323), .Q(
        \I_cache/cache[6][99] ), .QN(n436) );
  DFFRX1 \I_cache/cache_reg[7][99]  ( .D(n9365), .CK(clk), .RN(n4323), .Q(
        \I_cache/cache[7][99] ), .QN(n1351) );
  DFFRX1 \I_cache/cache_reg[0][100]  ( .D(n9364), .CK(clk), .RN(n4324), .Q(
        \I_cache/cache[0][100] ), .QN(n560) );
  DFFRX1 \I_cache/cache_reg[1][100]  ( .D(n9363), .CK(clk), .RN(n4324), .Q(
        \I_cache/cache[1][100] ), .QN(n1479) );
  DFFRX1 \I_cache/cache_reg[2][100]  ( .D(n9362), .CK(clk), .RN(n4324), .Q(
        \I_cache/cache[2][100] ), .QN(n559) );
  DFFRX1 \I_cache/cache_reg[3][100]  ( .D(n9361), .CK(clk), .RN(n4324), .Q(
        \I_cache/cache[3][100] ), .QN(n1478) );
  DFFRX1 \I_cache/cache_reg[4][100]  ( .D(n9360), .CK(clk), .RN(n4324), .Q(
        \I_cache/cache[4][100] ), .QN(n644) );
  DFFRX1 \I_cache/cache_reg[5][100]  ( .D(n9359), .CK(clk), .RN(n4324), .Q(
        \I_cache/cache[5][100] ), .QN(n1563) );
  DFFRX1 \I_cache/cache_reg[6][100]  ( .D(n9358), .CK(clk), .RN(n4324), .Q(
        \I_cache/cache[6][100] ), .QN(n470) );
  DFFRX1 \I_cache/cache_reg[7][100]  ( .D(n9357), .CK(clk), .RN(n4324), .Q(
        \I_cache/cache[7][100] ), .QN(n1385) );
  DFFRX1 \I_cache/cache_reg[0][101]  ( .D(n9356), .CK(clk), .RN(n4324), .Q(
        \I_cache/cache[0][101] ), .QN(n587) );
  DFFRX1 \I_cache/cache_reg[1][101]  ( .D(n9355), .CK(clk), .RN(n4324), .Q(
        \I_cache/cache[1][101] ), .QN(n1506) );
  DFFRX1 \I_cache/cache_reg[2][101]  ( .D(n9354), .CK(clk), .RN(n4324), .Q(
        \I_cache/cache[2][101] ), .QN(n586) );
  DFFRX1 \I_cache/cache_reg[3][101]  ( .D(n9353), .CK(clk), .RN(n4324), .Q(
        \I_cache/cache[3][101] ), .QN(n1505) );
  DFFRX1 \I_cache/cache_reg[4][101]  ( .D(n9352), .CK(clk), .RN(n4325), .Q(
        \I_cache/cache[4][101] ), .QN(n649) );
  DFFRX1 \I_cache/cache_reg[5][101]  ( .D(n9351), .CK(clk), .RN(n4325), .Q(
        \I_cache/cache[5][101] ), .QN(n1568) );
  DFFRX1 \I_cache/cache_reg[6][101]  ( .D(n9350), .CK(clk), .RN(n4325), .Q(
        \I_cache/cache[6][101] ), .QN(n585) );
  DFFRX1 \I_cache/cache_reg[7][101]  ( .D(n9349), .CK(clk), .RN(n4325), .Q(
        \I_cache/cache[7][101] ), .QN(n1504) );
  DFFRX1 \I_cache/cache_reg[0][102]  ( .D(n9348), .CK(clk), .RN(n4325), .Q(
        \I_cache/cache[0][102] ), .QN(n460) );
  DFFRX1 \I_cache/cache_reg[1][102]  ( .D(n9347), .CK(clk), .RN(n4325), .Q(
        \I_cache/cache[1][102] ), .QN(n1369) );
  DFFRX1 \I_cache/cache_reg[2][102]  ( .D(n9346), .CK(clk), .RN(n4325), .Q(
        \I_cache/cache[2][102] ), .QN(n493) );
  DFFRX1 \I_cache/cache_reg[3][102]  ( .D(n9345), .CK(clk), .RN(n4325), .Q(
        \I_cache/cache[3][102] ), .QN(n1411) );
  DFFRX1 \I_cache/cache_reg[4][102]  ( .D(n9344), .CK(clk), .RN(n4325), .Q(
        \I_cache/cache[4][102] ), .QN(n527) );
  DFFRX1 \I_cache/cache_reg[5][102]  ( .D(n9343), .CK(clk), .RN(n4325), .Q(
        \I_cache/cache[5][102] ), .QN(n1446) );
  DFFRX1 \I_cache/cache_reg[6][102]  ( .D(n9342), .CK(clk), .RN(n4325), .Q(
        \I_cache/cache[6][102] ), .QN(n492) );
  DFFRX1 \I_cache/cache_reg[7][102]  ( .D(n9341), .CK(clk), .RN(n4325), .Q(
        \I_cache/cache[7][102] ), .QN(n1410) );
  DFFRX1 \I_cache/cache_reg[0][103]  ( .D(n9340), .CK(clk), .RN(n4326), .Q(
        \I_cache/cache[0][103] ), .QN(n544) );
  DFFRX1 \I_cache/cache_reg[1][103]  ( .D(n9339), .CK(clk), .RN(n4326), .Q(
        \I_cache/cache[1][103] ), .QN(n1463) );
  DFFRX1 \I_cache/cache_reg[2][103]  ( .D(n9338), .CK(clk), .RN(n4326), .Q(
        \I_cache/cache[2][103] ), .QN(n464) );
  DFFRX1 \I_cache/cache_reg[3][103]  ( .D(n9337), .CK(clk), .RN(n4326), .Q(
        \I_cache/cache[3][103] ), .QN(n1379) );
  DFFRX1 \I_cache/cache_reg[4][103]  ( .D(n9336), .CK(clk), .RN(n4326), .Q(
        \I_cache/cache[4][103] ), .QN(n466) );
  DFFRX1 \I_cache/cache_reg[5][103]  ( .D(n9335), .CK(clk), .RN(n4326), .Q(
        \I_cache/cache[5][103] ), .QN(n1381) );
  DFFRX1 \I_cache/cache_reg[6][103]  ( .D(n9334), .CK(clk), .RN(n4326), .Q(
        \I_cache/cache[6][103] ), .QN(n465) );
  DFFRX1 \I_cache/cache_reg[7][103]  ( .D(n9333), .CK(clk), .RN(n4326), .Q(
        \I_cache/cache[7][103] ), .QN(n1380) );
  DFFRX1 \I_cache/cache_reg[0][104]  ( .D(n9332), .CK(clk), .RN(n4326), .Q(
        \I_cache/cache[0][104] ), .QN(n502) );
  DFFRX1 \I_cache/cache_reg[1][104]  ( .D(n9331), .CK(clk), .RN(n4326), .Q(
        \I_cache/cache[1][104] ), .QN(n1420) );
  DFFRX1 \I_cache/cache_reg[2][104]  ( .D(n9330), .CK(clk), .RN(n4326), .Q(
        \I_cache/cache[2][104] ), .QN(n500) );
  DFFRX1 \I_cache/cache_reg[3][104]  ( .D(n9329), .CK(clk), .RN(n4326), .Q(
        \I_cache/cache[3][104] ), .QN(n1418) );
  DFFRX1 \I_cache/cache_reg[4][104]  ( .D(n9328), .CK(clk), .RN(n4327), .Q(
        \I_cache/cache[4][104] ), .QN(n535) );
  DFFRX1 \I_cache/cache_reg[5][104]  ( .D(n9327), .CK(clk), .RN(n4327), .Q(
        \I_cache/cache[5][104] ), .QN(n1454) );
  DFFRX1 \I_cache/cache_reg[6][104]  ( .D(n9326), .CK(clk), .RN(n4327), .Q(
        \I_cache/cache[6][104] ), .QN(n501) );
  DFFRX1 \I_cache/cache_reg[7][104]  ( .D(n9325), .CK(clk), .RN(n4327), .Q(
        \I_cache/cache[7][104] ), .QN(n1419) );
  DFFRX1 \I_cache/cache_reg[0][105]  ( .D(n9324), .CK(clk), .RN(n4327), .Q(
        \I_cache/cache[0][105] ), .QN(n456) );
  DFFRX1 \I_cache/cache_reg[1][105]  ( .D(n9323), .CK(clk), .RN(n4327), .Q(
        \I_cache/cache[1][105] ), .QN(n1365) );
  DFFRX1 \I_cache/cache_reg[2][105]  ( .D(n9322), .CK(clk), .RN(n4327), .Q(
        \I_cache/cache[2][105] ), .QN(n505) );
  DFFRX1 \I_cache/cache_reg[3][105]  ( .D(n9321), .CK(clk), .RN(n4327), .Q(
        \I_cache/cache[3][105] ), .QN(n1423) );
  DFFRX1 \I_cache/cache_reg[4][105]  ( .D(n9320), .CK(clk), .RN(n4327), .Q(
        \I_cache/cache[4][105] ), .QN(n530) );
  DFFRX1 \I_cache/cache_reg[5][105]  ( .D(n9319), .CK(clk), .RN(n4327), .Q(
        \I_cache/cache[5][105] ), .QN(n1449) );
  DFFRX1 \I_cache/cache_reg[6][105]  ( .D(n9318), .CK(clk), .RN(n4327), .Q(
        \I_cache/cache[6][105] ), .QN(n506) );
  DFFRX1 \I_cache/cache_reg[7][105]  ( .D(n9317), .CK(clk), .RN(n4327), .Q(
        \I_cache/cache[7][105] ), .QN(n1424) );
  DFFRX1 \I_cache/cache_reg[1][106]  ( .D(n9315), .CK(clk), .RN(n4328), .Q(
        \I_cache/cache[1][106] ), .QN(n1545) );
  DFFRX1 \I_cache/cache_reg[3][106]  ( .D(n9313), .CK(clk), .RN(n4328), .Q(
        \I_cache/cache[3][106] ), .QN(n1544) );
  DFFRX1 \I_cache/cache_reg[4][106]  ( .D(n9312), .CK(clk), .RN(n4328), .Q(
        \I_cache/cache[4][106] ), .QN(n668) );
  DFFRX1 \I_cache/cache_reg[5][106]  ( .D(n9311), .CK(clk), .RN(n4328), .Q(
        \I_cache/cache[5][106] ), .QN(n1587) );
  DFFRX1 \I_cache/cache_reg[6][106]  ( .D(n9310), .CK(clk), .RN(n4328), .Q(
        \I_cache/cache[6][106] ), .QN(n624) );
  DFFRX1 \I_cache/cache_reg[7][106]  ( .D(n9309), .CK(clk), .RN(n4328), .Q(
        \I_cache/cache[7][106] ), .QN(n1543) );
  DFFRX1 \I_cache/cache_reg[0][107]  ( .D(n9308), .CK(clk), .RN(n4328), .Q(
        \I_cache/cache[0][107] ), .QN(n467) );
  DFFRX1 \I_cache/cache_reg[1][107]  ( .D(n9307), .CK(clk), .RN(n4328), .Q(
        \I_cache/cache[1][107] ), .QN(n1382) );
  DFFRX1 \I_cache/cache_reg[2][107]  ( .D(n9306), .CK(clk), .RN(n4328), .Q(
        \I_cache/cache[2][107] ), .QN(n469) );
  DFFRX1 \I_cache/cache_reg[3][107]  ( .D(n9305), .CK(clk), .RN(n4328), .Q(
        \I_cache/cache[3][107] ), .QN(n1384) );
  DFFRX1 \I_cache/cache_reg[4][107]  ( .D(n9304), .CK(clk), .RN(n4329), .Q(
        \I_cache/cache[4][107] ), .QN(n471) );
  DFFRX1 \I_cache/cache_reg[5][107]  ( .D(n9303), .CK(clk), .RN(n4329), .Q(
        \I_cache/cache[5][107] ), .QN(n1386) );
  DFFRX1 \I_cache/cache_reg[6][107]  ( .D(n9302), .CK(clk), .RN(n4329), .Q(
        \I_cache/cache[6][107] ), .QN(n468) );
  DFFRX1 \I_cache/cache_reg[7][107]  ( .D(n9301), .CK(clk), .RN(n4329), .Q(
        \I_cache/cache[7][107] ), .QN(n1383) );
  DFFRX1 \I_cache/cache_reg[0][108]  ( .D(n9300), .CK(clk), .RN(n4329), .Q(
        \I_cache/cache[0][108] ), .QN(n461) );
  DFFRX1 \I_cache/cache_reg[1][108]  ( .D(n9299), .CK(clk), .RN(n4329), .Q(
        \I_cache/cache[1][108] ), .QN(n1370) );
  DFFRX1 \I_cache/cache_reg[2][108]  ( .D(n9298), .CK(clk), .RN(n4329), .Q(
        \I_cache/cache[2][108] ), .QN(n510) );
  DFFRX1 \I_cache/cache_reg[3][108]  ( .D(n9297), .CK(clk), .RN(n4329), .Q(
        \I_cache/cache[3][108] ), .QN(n1428) );
  DFFRX1 \I_cache/cache_reg[4][108]  ( .D(n9296), .CK(clk), .RN(n4329), .Q(
        \I_cache/cache[4][108] ), .QN(n531) );
  DFFRX1 \I_cache/cache_reg[5][108]  ( .D(n9295), .CK(clk), .RN(n4329), .Q(
        \I_cache/cache[5][108] ), .QN(n1450) );
  DFFRX1 \I_cache/cache_reg[6][108]  ( .D(n9294), .CK(clk), .RN(n4329), .Q(
        \I_cache/cache[6][108] ), .QN(n511) );
  DFFRX1 \I_cache/cache_reg[7][108]  ( .D(n9293), .CK(clk), .RN(n4329), .Q(
        \I_cache/cache[7][108] ), .QN(n1429) );
  DFFRX1 \I_cache/cache_reg[0][109]  ( .D(n9292), .CK(clk), .RN(n4330), .Q(
        \I_cache/cache[0][109] ), .QN(n602) );
  DFFRX1 \I_cache/cache_reg[1][109]  ( .D(n9291), .CK(clk), .RN(n4330), .Q(
        \I_cache/cache[1][109] ), .QN(n1521) );
  DFFRX1 \I_cache/cache_reg[2][109]  ( .D(n9290), .CK(clk), .RN(n4330), .Q(
        \I_cache/cache[2][109] ), .QN(n601) );
  DFFRX1 \I_cache/cache_reg[3][109]  ( .D(n9289), .CK(clk), .RN(n4330), .Q(
        \I_cache/cache[3][109] ), .QN(n1520) );
  DFFRX1 \I_cache/cache_reg[4][109]  ( .D(n9288), .CK(clk), .RN(n4330), .Q(
        \I_cache/cache[4][109] ), .QN(n654) );
  DFFRX1 \I_cache/cache_reg[5][109]  ( .D(n9287), .CK(clk), .RN(n4330), .Q(
        \I_cache/cache[5][109] ), .QN(n1573) );
  DFFRX1 \I_cache/cache_reg[6][109]  ( .D(n9286), .CK(clk), .RN(n4330), .Q(
        \I_cache/cache[6][109] ), .QN(n600) );
  DFFRX1 \I_cache/cache_reg[7][109]  ( .D(n9285), .CK(clk), .RN(n4330), .Q(
        \I_cache/cache[7][109] ), .QN(n1519) );
  DFFRX1 \I_cache/cache_reg[0][110]  ( .D(n9284), .CK(clk), .RN(n4330), .Q(
        \I_cache/cache[0][110] ), .QN(n590) );
  DFFRX1 \I_cache/cache_reg[1][110]  ( .D(n9283), .CK(clk), .RN(n4330), .Q(
        \I_cache/cache[1][110] ), .QN(n1509) );
  DFFRX1 \I_cache/cache_reg[2][110]  ( .D(n9282), .CK(clk), .RN(n4330), .Q(
        \I_cache/cache[2][110] ), .QN(n589) );
  DFFRX1 \I_cache/cache_reg[3][110]  ( .D(n9281), .CK(clk), .RN(n4330), .Q(
        \I_cache/cache[3][110] ), .QN(n1508) );
  DFFRX1 \I_cache/cache_reg[4][110]  ( .D(n9280), .CK(clk), .RN(n4331), .Q(
        \I_cache/cache[4][110] ), .QN(n650) );
  DFFRX1 \I_cache/cache_reg[5][110]  ( .D(n9279), .CK(clk), .RN(n4331), .Q(
        \I_cache/cache[5][110] ), .QN(n1569) );
  DFFRX1 \I_cache/cache_reg[6][110]  ( .D(n9278), .CK(clk), .RN(n4331), .Q(
        \I_cache/cache[6][110] ), .QN(n588) );
  DFFRX1 \I_cache/cache_reg[7][110]  ( .D(n9277), .CK(clk), .RN(n4331), .Q(
        \I_cache/cache[7][110] ), .QN(n1507) );
  DFFRX1 \I_cache/cache_reg[0][111]  ( .D(n9276), .CK(clk), .RN(n4331), .Q(
        \I_cache/cache[0][111] ), .QN(n484) );
  DFFRX1 \I_cache/cache_reg[1][111]  ( .D(n9275), .CK(clk), .RN(n4331), .Q(
        \I_cache/cache[1][111] ), .QN(n1399) );
  DFFRX1 \I_cache/cache_reg[2][111]  ( .D(n9274), .CK(clk), .RN(n4331), .Q(
        \I_cache/cache[2][111] ), .QN(n485) );
  DFFRX1 \I_cache/cache_reg[3][111]  ( .D(n9273), .CK(clk), .RN(n4331), .Q(
        \I_cache/cache[3][111] ), .QN(n1400) );
  DFFRX1 \I_cache/cache_reg[4][111]  ( .D(n9272), .CK(clk), .RN(n4331), .Q(
        \I_cache/cache[4][111] ), .QN(n524) );
  DFFRX1 \I_cache/cache_reg[5][111]  ( .D(n9271), .CK(clk), .RN(n4331), .Q(
        \I_cache/cache[5][111] ), .QN(n1442) );
  DFFRX1 \I_cache/cache_reg[6][111]  ( .D(n9270), .CK(clk), .RN(n4331), .Q(
        \I_cache/cache[6][111] ), .QN(n486) );
  DFFRX1 \I_cache/cache_reg[7][111]  ( .D(n9269), .CK(clk), .RN(n4331), .Q(
        \I_cache/cache[7][111] ), .QN(n1401) );
  DFFRX1 \I_cache/cache_reg[0][153]  ( .D(n8940), .CK(clk), .RN(n4359), .Q(
        \I_cache/cache[0][153] ), .QN(n172) );
  DFFRX1 \I_cache/cache_reg[1][153]  ( .D(n8939), .CK(clk), .RN(n4359), .Q(
        \I_cache/cache[1][153] ), .QN(n1402) );
  DFFRX1 \I_cache/cache_reg[2][153]  ( .D(n8938), .CK(clk), .RN(n4359), .Q(
        \I_cache/cache[2][153] ), .QN(n174) );
  DFFRX1 \I_cache/cache_reg[3][153]  ( .D(n8937), .CK(clk), .RN(n4359), .Q(
        \I_cache/cache[3][153] ), .QN(n1404) );
  DFFRX1 \I_cache/cache_reg[4][153]  ( .D(n8936), .CK(clk), .RN(n4359), .Q(
        \I_cache/cache[4][153] ), .QN(n173) );
  DFFRX1 \I_cache/cache_reg[5][153]  ( .D(n8935), .CK(clk), .RN(n4359), .Q(
        \I_cache/cache[5][153] ), .QN(n1403) );
  DFFRX1 \I_cache/cache_reg[6][153]  ( .D(n8934), .CK(clk), .RN(n4359), .Q(
        \I_cache/cache[6][153] ), .QN(n175) );
  DFFRX1 \I_cache/cache_reg[7][153]  ( .D(n8933), .CK(clk), .RN(n4359), .Q(
        \I_cache/cache[7][153] ), .QN(n1444) );
  DFFRX1 \i_MIPS/ID_EX_reg[99]  ( .D(\i_MIPS/n486 ), .CK(clk), .RN(n4056), .Q(
        \i_MIPS/ID_EX[99] ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[0]  ( .D(\i_MIPS/n563 ), .CK(clk), .RN(n4065), .Q(
        \i_MIPS/EX_MEM_0 ), .QN(\i_MIPS/n373 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[48]  ( .D(\i_MIPS/N71 ), .CK(clk), .RN(n4060), .Q(
        \i_MIPS/IR_ID[16] ), .QN(\i_MIPS/n312 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[55]  ( .D(\i_MIPS/N78 ), .CK(clk), .RN(n4061), .Q(
        \i_MIPS/IR_ID[23] ), .QN(\i_MIPS/n230 ) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[25]  ( .D(\i_MIPS/PC/n59 ), .CK(clk), .RN(n4068), 
        .Q(ICACHE_addr[23]), .QN(\i_MIPS/PC/n27 ) );
  DFFRX2 \i_MIPS/EX_MEM_reg[69]  ( .D(\i_MIPS/n477 ), .CK(clk), .RN(n4056), 
        .Q(\i_MIPS/Reg_W[0] ), .QN(n963) );
  DFFRX2 \i_MIPS/EX_MEM_reg[70]  ( .D(\i_MIPS/n476 ), .CK(clk), .RN(n4056), 
        .Q(\i_MIPS/Reg_W[1] ), .QN(n78) );
  DFFRX2 \i_MIPS/EX_MEM_reg[71]  ( .D(\i_MIPS/n475 ), .CK(clk), .RN(n4055), 
        .Q(\i_MIPS/Reg_W[2] ), .QN(n53) );
  DFFRX2 \i_MIPS/EX_MEM_reg[73]  ( .D(\i_MIPS/n473 ), .CK(clk), .RN(n4055), 
        .Q(\i_MIPS/Reg_W[4] ), .QN(n2996) );
  DFFRX2 \i_MIPS/EX_MEM_reg[72]  ( .D(\i_MIPS/n474 ), .CK(clk), .RN(n4055), 
        .Q(\i_MIPS/Reg_W[3] ), .QN(n2997) );
  DFFRX1 \i_MIPS/ID_EX_reg[108]  ( .D(\i_MIPS/n521 ), .CK(clk), .RN(n4062), 
        .QN(\i_MIPS/n329 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[72]  ( .D(\i_MIPS/n375 ), .CK(clk), .RN(n4047), .Q(
        n1885), .QN(\i_MIPS/n247 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[71]  ( .D(\i_MIPS/n377 ), .CK(clk), .RN(n4047), .Q(
        \i_MIPS/ID_EX[71] ), .QN(\i_MIPS/n249 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[70]  ( .D(\i_MIPS/n379 ), .CK(clk), .RN(n4047), .Q(
        \i_MIPS/ID_EX[70] ), .QN(\i_MIPS/n251 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[69]  ( .D(\i_MIPS/n381 ), .CK(clk), .RN(n4048), .Q(
        \i_MIPS/ID_EX[69] ), .QN(\i_MIPS/n253 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[68]  ( .D(\i_MIPS/n383 ), .CK(clk), .RN(n4048), .Q(
        \i_MIPS/ID_EX[68] ), .QN(\i_MIPS/n255 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[66]  ( .D(\i_MIPS/n387 ), .CK(clk), .RN(n4048), .Q(
        \i_MIPS/ID_EX[66] ), .QN(\i_MIPS/n259 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[65]  ( .D(\i_MIPS/n389 ), .CK(clk), .RN(n4048), .Q(
        \i_MIPS/ID_EX[65] ), .QN(\i_MIPS/n261 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[64]  ( .D(\i_MIPS/n391 ), .CK(clk), .RN(n4048), .Q(
        \i_MIPS/ID_EX[64] ), .QN(\i_MIPS/n263 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[63]  ( .D(\i_MIPS/n393 ), .CK(clk), .RN(n4049), .Q(
        \i_MIPS/ID_EX[63] ), .QN(\i_MIPS/n265 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[62]  ( .D(\i_MIPS/n395 ), .CK(clk), .RN(n4049), .Q(
        \i_MIPS/ID_EX[62] ), .QN(\i_MIPS/n267 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[61]  ( .D(\i_MIPS/n397 ), .CK(clk), .RN(n4049), .Q(
        \i_MIPS/ID_EX[61] ), .QN(\i_MIPS/n269 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[60]  ( .D(\i_MIPS/n399 ), .CK(clk), .RN(n4049), .Q(
        \i_MIPS/ID_EX[60] ), .QN(\i_MIPS/n271 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[59]  ( .D(\i_MIPS/n401 ), .CK(clk), .RN(n4049), .Q(
        \i_MIPS/ID_EX[59] ), .QN(\i_MIPS/n273 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[58]  ( .D(\i_MIPS/n403 ), .CK(clk), .RN(n4049), .Q(
        \i_MIPS/ID_EX[58] ), .QN(\i_MIPS/n275 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[56]  ( .D(\i_MIPS/n407 ), .CK(clk), .RN(n4050), .Q(
        n1882), .QN(\i_MIPS/n279 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[55]  ( .D(\i_MIPS/n409 ), .CK(clk), .RN(n4050), .Q(
        n1883), .QN(\i_MIPS/n281 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[53]  ( .D(\i_MIPS/n413 ), .CK(clk), .RN(n4050), .Q(
        n1891), .QN(\i_MIPS/n285 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[52]  ( .D(\i_MIPS/n415 ), .CK(clk), .RN(n4050), .Q(
        \i_MIPS/ID_EX[52] ), .QN(\i_MIPS/n287 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[51]  ( .D(\i_MIPS/n417 ), .CK(clk), .RN(n4051), .Q(
        n1890), .QN(\i_MIPS/n289 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[49]  ( .D(\i_MIPS/n421 ), .CK(clk), .RN(n4051), .Q(
        \i_MIPS/ID_EX[49] ), .QN(\i_MIPS/n293 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[45]  ( .D(\i_MIPS/n429 ), .CK(clk), .RN(n4052), .Q(
        n1881), .QN(\i_MIPS/n301 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[47]  ( .D(\i_MIPS/n425 ), .CK(clk), .RN(n4051), .Q(
        \i_MIPS/ID_EX[47] ), .QN(\i_MIPS/n297 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[110]  ( .D(\i_MIPS/n523 ), .CK(clk), .RN(n4062), 
        .Q(\i_MIPS/ID_EX[110] ), .QN(\i_MIPS/n333 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[109]  ( .D(\i_MIPS/n522 ), .CK(clk), .RN(n4062), 
        .Q(\i_MIPS/ID_EX[109] ), .QN(\i_MIPS/n331 ) );
  DFFRX1 \D_cache/cache_reg[3][128]  ( .D(\D_cache/n769 ), .CK(clk), .RN(n4239), .Q(\D_cache/cache[3][128] ) );
  DFFRX1 \D_cache/cache_reg[3][129]  ( .D(\D_cache/n761 ), .CK(clk), .RN(n4240), .Q(\D_cache/cache[3][129] ) );
  DFFRX1 \D_cache/cache_reg[7][129]  ( .D(\D_cache/n757 ), .CK(clk), .RN(n4240), .Q(\D_cache/cache[7][129] ) );
  DFFRX1 \D_cache/cache_reg[3][130]  ( .D(\D_cache/n753 ), .CK(clk), .RN(n4240), .Q(\D_cache/cache[3][130] ) );
  DFFRX1 \D_cache/cache_reg[7][130]  ( .D(\D_cache/n749 ), .CK(clk), .RN(n4241), .Q(\D_cache/cache[7][130] ) );
  DFFRX1 \D_cache/cache_reg[3][131]  ( .D(\D_cache/n745 ), .CK(clk), .RN(n4241), .Q(\D_cache/cache[3][131] ) );
  DFFRX1 \D_cache/cache_reg[7][131]  ( .D(\D_cache/n741 ), .CK(clk), .RN(n4241), .Q(\D_cache/cache[7][131] ) );
  DFFRX1 \D_cache/cache_reg[3][132]  ( .D(\D_cache/n737 ), .CK(clk), .RN(n4242), .Q(\D_cache/cache[3][132] ) );
  DFFRX1 \D_cache/cache_reg[7][132]  ( .D(\D_cache/n733 ), .CK(clk), .RN(n4242), .Q(\D_cache/cache[7][132] ) );
  DFFRX1 \D_cache/cache_reg[3][133]  ( .D(\D_cache/n729 ), .CK(clk), .RN(n4242), .Q(\D_cache/cache[3][133] ) );
  DFFRX1 \D_cache/cache_reg[7][133]  ( .D(\D_cache/n725 ), .CK(clk), .RN(n4243), .Q(\D_cache/cache[7][133] ) );
  DFFRX1 \D_cache/cache_reg[3][134]  ( .D(\D_cache/n721 ), .CK(clk), .RN(n4243), .Q(\D_cache/cache[3][134] ) );
  DFFRX1 \D_cache/cache_reg[7][134]  ( .D(\D_cache/n717 ), .CK(clk), .RN(n4243), .Q(\D_cache/cache[7][134] ) );
  DFFRX1 \D_cache/cache_reg[3][138]  ( .D(\D_cache/n689 ), .CK(clk), .RN(n4246), .Q(\D_cache/cache[3][138] ) );
  DFFRX1 \D_cache/cache_reg[7][138]  ( .D(\D_cache/n685 ), .CK(clk), .RN(n4246), .Q(\D_cache/cache[7][138] ) );
  DFFRX1 \D_cache/cache_reg[3][139]  ( .D(\D_cache/n681 ), .CK(clk), .RN(n4246), .Q(\D_cache/cache[3][139] ) );
  DFFRX1 \D_cache/cache_reg[3][140]  ( .D(\D_cache/n673 ), .CK(clk), .RN(n4247), .Q(\D_cache/cache[3][140] ) );
  DFFRX1 \D_cache/cache_reg[7][140]  ( .D(\D_cache/n669 ), .CK(clk), .RN(n4247), .Q(\D_cache/cache[7][140] ) );
  DFFRX1 \D_cache/cache_reg[3][141]  ( .D(\D_cache/n665 ), .CK(clk), .RN(n4248), .Q(\D_cache/cache[3][141] ) );
  DFFRX1 \D_cache/cache_reg[7][141]  ( .D(\D_cache/n661 ), .CK(clk), .RN(n4248), .Q(\D_cache/cache[7][141] ) );
  DFFRX1 \D_cache/cache_reg[3][142]  ( .D(\D_cache/n657 ), .CK(clk), .RN(n4248), .Q(\D_cache/cache[3][142] ) );
  DFFRX1 \D_cache/cache_reg[7][142]  ( .D(\D_cache/n653 ), .CK(clk), .RN(n4249), .Q(\D_cache/cache[7][142] ) );
  DFFRX1 \D_cache/cache_reg[3][143]  ( .D(\D_cache/n649 ), .CK(clk), .RN(n4249), .Q(\D_cache/cache[3][143] ) );
  DFFRX1 \D_cache/cache_reg[7][143]  ( .D(\D_cache/n645 ), .CK(clk), .RN(n4249), .Q(\D_cache/cache[7][143] ) );
  DFFRX1 \D_cache/cache_reg[3][144]  ( .D(\D_cache/n641 ), .CK(clk), .RN(n4250), .Q(\D_cache/cache[3][144] ) );
  DFFRX1 \D_cache/cache_reg[7][144]  ( .D(\D_cache/n637 ), .CK(clk), .RN(n4250), .Q(\D_cache/cache[7][144] ) );
  DFFRX1 \D_cache/cache_reg[3][145]  ( .D(\D_cache/n633 ), .CK(clk), .RN(n4250), .Q(\D_cache/cache[3][145] ) );
  DFFRX1 \D_cache/cache_reg[7][145]  ( .D(\D_cache/n629 ), .CK(clk), .RN(n4251), .Q(\D_cache/cache[7][145] ) );
  DFFRX1 \D_cache/cache_reg[3][146]  ( .D(\D_cache/n625 ), .CK(clk), .RN(n4251), .Q(\D_cache/cache[3][146] ) );
  DFFRX1 \D_cache/cache_reg[7][146]  ( .D(\D_cache/n621 ), .CK(clk), .RN(n4251), .Q(\D_cache/cache[7][146] ) );
  DFFRX1 \D_cache/cache_reg[3][147]  ( .D(\D_cache/n617 ), .CK(clk), .RN(n4252), .Q(\D_cache/cache[3][147] ) );
  DFFRX1 \D_cache/cache_reg[7][147]  ( .D(\D_cache/n613 ), .CK(clk), .RN(n4252), .Q(\D_cache/cache[7][147] ) );
  DFFRX1 \D_cache/cache_reg[3][148]  ( .D(\D_cache/n609 ), .CK(clk), .RN(n4252), .Q(\D_cache/cache[3][148] ) );
  DFFRX1 \D_cache/cache_reg[7][148]  ( .D(\D_cache/n605 ), .CK(clk), .RN(n4253), .Q(\D_cache/cache[7][148] ) );
  DFFRX1 \D_cache/cache_reg[3][150]  ( .D(\D_cache/n593 ), .CK(clk), .RN(n4254), .Q(\D_cache/cache[3][150] ) );
  DFFRX1 \D_cache/cache_reg[7][150]  ( .D(\D_cache/n589 ), .CK(clk), .RN(n4254), .Q(\D_cache/cache[7][150] ) );
  DFFRX1 \D_cache/cache_reg[3][151]  ( .D(\D_cache/n585 ), .CK(clk), .RN(n4254), .Q(\D_cache/cache[3][151] ) );
  DFFRX1 \D_cache/cache_reg[3][152]  ( .D(\D_cache/n577 ), .CK(clk), .RN(n4255), .Q(\D_cache/cache[3][152] ) );
  DFFRX1 \D_cache/cache_reg[7][152]  ( .D(\D_cache/n573 ), .CK(clk), .RN(n4255), .Q(\D_cache/cache[7][152] ) );
  DFFRX1 \D_cache/cache_reg[7][128]  ( .D(\D_cache/n765 ), .CK(clk), .RN(n4256), .Q(\D_cache/cache[7][128] ) );
  DFFRX1 \D_cache/cache_reg[1][128]  ( .D(\D_cache/n771 ), .CK(clk), .RN(n4239), .Q(\D_cache/cache[1][128] ) );
  DFFRX1 \D_cache/cache_reg[5][128]  ( .D(\D_cache/n767 ), .CK(clk), .RN(n4239), .Q(\D_cache/cache[5][128] ) );
  DFFRX1 \D_cache/cache_reg[1][129]  ( .D(\D_cache/n763 ), .CK(clk), .RN(n4240), .Q(\D_cache/cache[1][129] ) );
  DFFRX1 \D_cache/cache_reg[5][129]  ( .D(\D_cache/n759 ), .CK(clk), .RN(n4240), .Q(\D_cache/cache[5][129] ) );
  DFFRX1 \D_cache/cache_reg[1][130]  ( .D(\D_cache/n755 ), .CK(clk), .RN(n4240), .Q(\D_cache/cache[1][130] ) );
  DFFRX1 \D_cache/cache_reg[5][130]  ( .D(\D_cache/n751 ), .CK(clk), .RN(n4241), .Q(\D_cache/cache[5][130] ) );
  DFFRX1 \D_cache/cache_reg[1][131]  ( .D(\D_cache/n747 ), .CK(clk), .RN(n4241), .Q(\D_cache/cache[1][131] ) );
  DFFRX1 \D_cache/cache_reg[5][131]  ( .D(\D_cache/n743 ), .CK(clk), .RN(n4241), .Q(\D_cache/cache[5][131] ) );
  DFFRX1 \D_cache/cache_reg[1][132]  ( .D(\D_cache/n739 ), .CK(clk), .RN(n4242), .Q(\D_cache/cache[1][132] ) );
  DFFRX1 \D_cache/cache_reg[5][132]  ( .D(\D_cache/n735 ), .CK(clk), .RN(n4242), .Q(\D_cache/cache[5][132] ) );
  DFFRX1 \D_cache/cache_reg[1][133]  ( .D(\D_cache/n731 ), .CK(clk), .RN(n4242), .Q(\D_cache/cache[1][133] ) );
  DFFRX1 \D_cache/cache_reg[5][133]  ( .D(\D_cache/n727 ), .CK(clk), .RN(n4243), .Q(\D_cache/cache[5][133] ) );
  DFFRX1 \D_cache/cache_reg[1][134]  ( .D(\D_cache/n723 ), .CK(clk), .RN(n4243), .Q(\D_cache/cache[1][134] ) );
  DFFRX1 \D_cache/cache_reg[5][134]  ( .D(\D_cache/n719 ), .CK(clk), .RN(n4243), .Q(\D_cache/cache[5][134] ) );
  DFFRX1 \D_cache/cache_reg[1][138]  ( .D(\D_cache/n691 ), .CK(clk), .RN(n4246), .Q(\D_cache/cache[1][138] ) );
  DFFRX1 \D_cache/cache_reg[5][138]  ( .D(\D_cache/n687 ), .CK(clk), .RN(n4246), .Q(\D_cache/cache[5][138] ) );
  DFFRX1 \D_cache/cache_reg[1][139]  ( .D(\D_cache/n683 ), .CK(clk), .RN(n4246), .Q(\D_cache/cache[1][139] ) );
  DFFRX1 \D_cache/cache_reg[5][139]  ( .D(\D_cache/n679 ), .CK(clk), .RN(n4247), .Q(\D_cache/cache[5][139] ) );
  DFFRX1 \D_cache/cache_reg[1][140]  ( .D(\D_cache/n675 ), .CK(clk), .RN(n4247), .Q(\D_cache/cache[1][140] ) );
  DFFRX1 \D_cache/cache_reg[5][140]  ( .D(\D_cache/n671 ), .CK(clk), .RN(n4247), .Q(\D_cache/cache[5][140] ) );
  DFFRX1 \D_cache/cache_reg[1][141]  ( .D(\D_cache/n667 ), .CK(clk), .RN(n4248), .Q(\D_cache/cache[1][141] ) );
  DFFRX1 \D_cache/cache_reg[5][141]  ( .D(\D_cache/n663 ), .CK(clk), .RN(n4248), .Q(\D_cache/cache[5][141] ) );
  DFFRX1 \D_cache/cache_reg[1][142]  ( .D(\D_cache/n659 ), .CK(clk), .RN(n4248), .Q(\D_cache/cache[1][142] ) );
  DFFRX1 \D_cache/cache_reg[5][142]  ( .D(\D_cache/n655 ), .CK(clk), .RN(n4249), .Q(\D_cache/cache[5][142] ) );
  DFFRX1 \D_cache/cache_reg[1][143]  ( .D(\D_cache/n651 ), .CK(clk), .RN(n4249), .Q(\D_cache/cache[1][143] ) );
  DFFRX1 \D_cache/cache_reg[5][143]  ( .D(\D_cache/n647 ), .CK(clk), .RN(n4249), .Q(\D_cache/cache[5][143] ) );
  DFFRX1 \D_cache/cache_reg[1][144]  ( .D(\D_cache/n643 ), .CK(clk), .RN(n4250), .Q(\D_cache/cache[1][144] ) );
  DFFRX1 \D_cache/cache_reg[5][144]  ( .D(\D_cache/n639 ), .CK(clk), .RN(n4250), .Q(\D_cache/cache[5][144] ) );
  DFFRX1 \D_cache/cache_reg[1][145]  ( .D(\D_cache/n635 ), .CK(clk), .RN(n4250), .Q(\D_cache/cache[1][145] ) );
  DFFRX1 \D_cache/cache_reg[5][145]  ( .D(\D_cache/n631 ), .CK(clk), .RN(n4251), .Q(\D_cache/cache[5][145] ) );
  DFFRX1 \D_cache/cache_reg[1][146]  ( .D(\D_cache/n627 ), .CK(clk), .RN(n4251), .Q(\D_cache/cache[1][146] ) );
  DFFRX1 \D_cache/cache_reg[5][146]  ( .D(\D_cache/n623 ), .CK(clk), .RN(n4251), .Q(\D_cache/cache[5][146] ) );
  DFFRX1 \D_cache/cache_reg[1][147]  ( .D(\D_cache/n619 ), .CK(clk), .RN(n4252), .Q(\D_cache/cache[1][147] ) );
  DFFRX1 \D_cache/cache_reg[5][147]  ( .D(\D_cache/n615 ), .CK(clk), .RN(n4252), .Q(\D_cache/cache[5][147] ) );
  DFFRX1 \D_cache/cache_reg[1][148]  ( .D(\D_cache/n611 ), .CK(clk), .RN(n4252), .Q(\D_cache/cache[1][148] ) );
  DFFRX1 \D_cache/cache_reg[5][148]  ( .D(\D_cache/n607 ), .CK(clk), .RN(n4253), .Q(\D_cache/cache[5][148] ) );
  DFFRX1 \D_cache/cache_reg[1][149]  ( .D(\D_cache/n603 ), .CK(clk), .RN(n4253), .Q(\D_cache/cache[1][149] ) );
  DFFRX1 \D_cache/cache_reg[5][149]  ( .D(\D_cache/n599 ), .CK(clk), .RN(n4253), .Q(\D_cache/cache[5][149] ) );
  DFFRX1 \D_cache/cache_reg[1][150]  ( .D(\D_cache/n595 ), .CK(clk), .RN(n4254), .Q(\D_cache/cache[1][150] ) );
  DFFRX1 \D_cache/cache_reg[5][150]  ( .D(\D_cache/n591 ), .CK(clk), .RN(n4254), .Q(\D_cache/cache[5][150] ) );
  DFFRX1 \D_cache/cache_reg[1][151]  ( .D(\D_cache/n587 ), .CK(clk), .RN(n4254), .Q(\D_cache/cache[1][151] ) );
  DFFRX1 \D_cache/cache_reg[5][151]  ( .D(\D_cache/n583 ), .CK(clk), .RN(n4255), .Q(\D_cache/cache[5][151] ) );
  DFFRX1 \D_cache/cache_reg[1][152]  ( .D(\D_cache/n579 ), .CK(clk), .RN(n4255), .Q(\D_cache/cache[1][152] ) );
  DFFRX1 \D_cache/cache_reg[5][152]  ( .D(\D_cache/n575 ), .CK(clk), .RN(n4255), .Q(\D_cache/cache[5][152] ) );
  DFFRX1 \D_cache/cache_reg[0][128]  ( .D(\D_cache/n772 ), .CK(clk), .RN(n4239), .Q(\D_cache/cache[0][128] ) );
  DFFRX1 \D_cache/cache_reg[4][128]  ( .D(\D_cache/n768 ), .CK(clk), .RN(n4239), .Q(\D_cache/cache[4][128] ) );
  DFFRX1 \D_cache/cache_reg[0][129]  ( .D(\D_cache/n764 ), .CK(clk), .RN(n4239), .Q(\D_cache/cache[0][129] ) );
  DFFRX1 \D_cache/cache_reg[4][129]  ( .D(\D_cache/n760 ), .CK(clk), .RN(n4240), .Q(\D_cache/cache[4][129] ) );
  DFFRX1 \D_cache/cache_reg[0][130]  ( .D(\D_cache/n756 ), .CK(clk), .RN(n4240), .Q(\D_cache/cache[0][130] ) );
  DFFRX1 \D_cache/cache_reg[4][130]  ( .D(\D_cache/n752 ), .CK(clk), .RN(n4240), .Q(\D_cache/cache[4][130] ) );
  DFFRX1 \D_cache/cache_reg[0][131]  ( .D(\D_cache/n748 ), .CK(clk), .RN(n4241), .Q(\D_cache/cache[0][131] ) );
  DFFRX1 \D_cache/cache_reg[4][131]  ( .D(\D_cache/n744 ), .CK(clk), .RN(n4241), .Q(\D_cache/cache[4][131] ) );
  DFFRX1 \D_cache/cache_reg[0][132]  ( .D(\D_cache/n740 ), .CK(clk), .RN(n4241), .Q(\D_cache/cache[0][132] ) );
  DFFRX1 \D_cache/cache_reg[4][132]  ( .D(\D_cache/n736 ), .CK(clk), .RN(n4242), .Q(\D_cache/cache[4][132] ) );
  DFFRX1 \D_cache/cache_reg[0][133]  ( .D(\D_cache/n732 ), .CK(clk), .RN(n4242), .Q(\D_cache/cache[0][133] ) );
  DFFRX1 \D_cache/cache_reg[4][133]  ( .D(\D_cache/n728 ), .CK(clk), .RN(n4242), .Q(\D_cache/cache[4][133] ) );
  DFFRX1 \D_cache/cache_reg[0][134]  ( .D(\D_cache/n724 ), .CK(clk), .RN(n4243), .Q(\D_cache/cache[0][134] ) );
  DFFRX1 \D_cache/cache_reg[4][134]  ( .D(\D_cache/n720 ), .CK(clk), .RN(n4243), .Q(\D_cache/cache[4][134] ) );
  DFFRX1 \D_cache/cache_reg[0][138]  ( .D(\D_cache/n692 ), .CK(clk), .RN(n4245), .Q(\D_cache/cache[0][138] ) );
  DFFRX1 \D_cache/cache_reg[4][138]  ( .D(\D_cache/n688 ), .CK(clk), .RN(n4246), .Q(\D_cache/cache[4][138] ) );
  DFFRX1 \D_cache/cache_reg[0][139]  ( .D(\D_cache/n684 ), .CK(clk), .RN(n4246), .Q(\D_cache/cache[0][139] ) );
  DFFRX1 \D_cache/cache_reg[4][139]  ( .D(\D_cache/n680 ), .CK(clk), .RN(n4246), .Q(\D_cache/cache[4][139] ) );
  DFFRX1 \D_cache/cache_reg[0][140]  ( .D(\D_cache/n676 ), .CK(clk), .RN(n4247), .Q(\D_cache/cache[0][140] ) );
  DFFRX1 \D_cache/cache_reg[4][140]  ( .D(\D_cache/n672 ), .CK(clk), .RN(n4247), .Q(\D_cache/cache[4][140] ) );
  DFFRX1 \D_cache/cache_reg[0][141]  ( .D(\D_cache/n668 ), .CK(clk), .RN(n4247), .Q(\D_cache/cache[0][141] ) );
  DFFRX1 \D_cache/cache_reg[4][141]  ( .D(\D_cache/n664 ), .CK(clk), .RN(n4248), .Q(\D_cache/cache[4][141] ) );
  DFFRX1 \D_cache/cache_reg[0][142]  ( .D(\D_cache/n660 ), .CK(clk), .RN(n4248), .Q(\D_cache/cache[0][142] ) );
  DFFRX1 \D_cache/cache_reg[4][142]  ( .D(\D_cache/n656 ), .CK(clk), .RN(n4248), .Q(\D_cache/cache[4][142] ) );
  DFFRX1 \D_cache/cache_reg[0][143]  ( .D(\D_cache/n652 ), .CK(clk), .RN(n4249), .Q(\D_cache/cache[0][143] ) );
  DFFRX1 \D_cache/cache_reg[4][143]  ( .D(\D_cache/n648 ), .CK(clk), .RN(n4249), .Q(\D_cache/cache[4][143] ) );
  DFFRX1 \D_cache/cache_reg[0][144]  ( .D(\D_cache/n644 ), .CK(clk), .RN(n4249), .Q(\D_cache/cache[0][144] ) );
  DFFRX1 \D_cache/cache_reg[4][144]  ( .D(\D_cache/n640 ), .CK(clk), .RN(n4250), .Q(\D_cache/cache[4][144] ) );
  DFFRX1 \D_cache/cache_reg[0][145]  ( .D(\D_cache/n636 ), .CK(clk), .RN(n4250), .Q(\D_cache/cache[0][145] ) );
  DFFRX1 \D_cache/cache_reg[4][145]  ( .D(\D_cache/n632 ), .CK(clk), .RN(n4250), .Q(\D_cache/cache[4][145] ) );
  DFFRX1 \D_cache/cache_reg[0][146]  ( .D(\D_cache/n628 ), .CK(clk), .RN(n4251), .Q(\D_cache/cache[0][146] ) );
  DFFRX1 \D_cache/cache_reg[4][146]  ( .D(\D_cache/n624 ), .CK(clk), .RN(n4251), .Q(\D_cache/cache[4][146] ) );
  DFFRX1 \D_cache/cache_reg[0][147]  ( .D(\D_cache/n620 ), .CK(clk), .RN(n4251), .Q(\D_cache/cache[0][147] ) );
  DFFRX1 \D_cache/cache_reg[4][147]  ( .D(\D_cache/n616 ), .CK(clk), .RN(n4252), .Q(\D_cache/cache[4][147] ) );
  DFFRX1 \D_cache/cache_reg[0][148]  ( .D(\D_cache/n612 ), .CK(clk), .RN(n4252), .Q(\D_cache/cache[0][148] ) );
  DFFRX1 \D_cache/cache_reg[4][148]  ( .D(\D_cache/n608 ), .CK(clk), .RN(n4252), .Q(\D_cache/cache[4][148] ) );
  DFFRX1 \D_cache/cache_reg[0][149]  ( .D(\D_cache/n604 ), .CK(clk), .RN(n4253), .Q(\D_cache/cache[0][149] ) );
  DFFRX1 \D_cache/cache_reg[4][149]  ( .D(\D_cache/n600 ), .CK(clk), .RN(n4253), .Q(\D_cache/cache[4][149] ) );
  DFFRX1 \D_cache/cache_reg[0][150]  ( .D(\D_cache/n596 ), .CK(clk), .RN(n4253), .Q(\D_cache/cache[0][150] ) );
  DFFRX1 \D_cache/cache_reg[4][150]  ( .D(\D_cache/n592 ), .CK(clk), .RN(n4254), .Q(\D_cache/cache[4][150] ) );
  DFFRX1 \D_cache/cache_reg[0][151]  ( .D(\D_cache/n588 ), .CK(clk), .RN(n4254), .Q(\D_cache/cache[0][151] ) );
  DFFRX1 \D_cache/cache_reg[4][151]  ( .D(\D_cache/n584 ), .CK(clk), .RN(n4254), .Q(\D_cache/cache[4][151] ) );
  DFFRX1 \D_cache/cache_reg[0][152]  ( .D(\D_cache/n580 ), .CK(clk), .RN(n4255), .Q(\D_cache/cache[0][152] ) );
  DFFRX1 \D_cache/cache_reg[4][152]  ( .D(\D_cache/n576 ), .CK(clk), .RN(n4255), .Q(\D_cache/cache[4][152] ) );
  DFFRX1 \D_cache/cache_reg[2][128]  ( .D(\D_cache/n770 ), .CK(clk), .RN(n4239), .Q(\D_cache/cache[2][128] ) );
  DFFRX1 \D_cache/cache_reg[6][128]  ( .D(\D_cache/n766 ), .CK(clk), .RN(n4239), .Q(\D_cache/cache[6][128] ) );
  DFFRX1 \D_cache/cache_reg[2][129]  ( .D(\D_cache/n762 ), .CK(clk), .RN(n4240), .Q(\D_cache/cache[2][129] ) );
  DFFRX1 \D_cache/cache_reg[6][129]  ( .D(\D_cache/n758 ), .CK(clk), .RN(n4240), .Q(\D_cache/cache[6][129] ) );
  DFFRX1 \D_cache/cache_reg[2][130]  ( .D(\D_cache/n754 ), .CK(clk), .RN(n4240), .Q(\D_cache/cache[2][130] ) );
  DFFRX1 \D_cache/cache_reg[6][130]  ( .D(\D_cache/n750 ), .CK(clk), .RN(n4241), .Q(\D_cache/cache[6][130] ) );
  DFFRX1 \D_cache/cache_reg[2][131]  ( .D(\D_cache/n746 ), .CK(clk), .RN(n4241), .Q(\D_cache/cache[2][131] ) );
  DFFRX1 \D_cache/cache_reg[6][131]  ( .D(\D_cache/n742 ), .CK(clk), .RN(n4241), .Q(\D_cache/cache[6][131] ) );
  DFFRX1 \D_cache/cache_reg[2][132]  ( .D(\D_cache/n738 ), .CK(clk), .RN(n4242), .Q(\D_cache/cache[2][132] ) );
  DFFRX1 \D_cache/cache_reg[6][132]  ( .D(\D_cache/n734 ), .CK(clk), .RN(n4242), .Q(\D_cache/cache[6][132] ) );
  DFFRX1 \D_cache/cache_reg[2][133]  ( .D(\D_cache/n730 ), .CK(clk), .RN(n4242), .Q(\D_cache/cache[2][133] ) );
  DFFRX1 \D_cache/cache_reg[6][133]  ( .D(\D_cache/n726 ), .CK(clk), .RN(n4243), .Q(\D_cache/cache[6][133] ) );
  DFFRX1 \D_cache/cache_reg[2][134]  ( .D(\D_cache/n722 ), .CK(clk), .RN(n4243), .Q(\D_cache/cache[2][134] ) );
  DFFRX1 \D_cache/cache_reg[6][134]  ( .D(\D_cache/n718 ), .CK(clk), .RN(n4243), .Q(\D_cache/cache[6][134] ) );
  DFFRX1 \D_cache/cache_reg[2][138]  ( .D(\D_cache/n690 ), .CK(clk), .RN(n4246), .Q(\D_cache/cache[2][138] ) );
  DFFRX1 \D_cache/cache_reg[6][138]  ( .D(\D_cache/n686 ), .CK(clk), .RN(n4246), .Q(\D_cache/cache[6][138] ) );
  DFFRX1 \D_cache/cache_reg[2][139]  ( .D(\D_cache/n682 ), .CK(clk), .RN(n4246), .Q(\D_cache/cache[2][139] ) );
  DFFRX1 \D_cache/cache_reg[2][140]  ( .D(\D_cache/n674 ), .CK(clk), .RN(n4247), .Q(\D_cache/cache[2][140] ) );
  DFFRX1 \D_cache/cache_reg[6][140]  ( .D(\D_cache/n670 ), .CK(clk), .RN(n4247), .Q(\D_cache/cache[6][140] ) );
  DFFRX1 \D_cache/cache_reg[2][141]  ( .D(\D_cache/n666 ), .CK(clk), .RN(n4248), .Q(\D_cache/cache[2][141] ) );
  DFFRX1 \D_cache/cache_reg[6][141]  ( .D(\D_cache/n662 ), .CK(clk), .RN(n4248), .Q(\D_cache/cache[6][141] ) );
  DFFRX1 \D_cache/cache_reg[2][142]  ( .D(\D_cache/n658 ), .CK(clk), .RN(n4248), .Q(\D_cache/cache[2][142] ) );
  DFFRX1 \D_cache/cache_reg[6][142]  ( .D(\D_cache/n654 ), .CK(clk), .RN(n4249), .Q(\D_cache/cache[6][142] ) );
  DFFRX1 \D_cache/cache_reg[2][143]  ( .D(\D_cache/n650 ), .CK(clk), .RN(n4249), .Q(\D_cache/cache[2][143] ) );
  DFFRX1 \D_cache/cache_reg[6][143]  ( .D(\D_cache/n646 ), .CK(clk), .RN(n4249), .Q(\D_cache/cache[6][143] ) );
  DFFRX1 \D_cache/cache_reg[2][144]  ( .D(\D_cache/n642 ), .CK(clk), .RN(n4250), .Q(\D_cache/cache[2][144] ) );
  DFFRX1 \D_cache/cache_reg[6][144]  ( .D(\D_cache/n638 ), .CK(clk), .RN(n4250), .Q(\D_cache/cache[6][144] ) );
  DFFRX1 \D_cache/cache_reg[2][145]  ( .D(\D_cache/n634 ), .CK(clk), .RN(n4250), .Q(\D_cache/cache[2][145] ) );
  DFFRX1 \D_cache/cache_reg[6][145]  ( .D(\D_cache/n630 ), .CK(clk), .RN(n4251), .Q(\D_cache/cache[6][145] ) );
  DFFRX1 \D_cache/cache_reg[2][146]  ( .D(\D_cache/n626 ), .CK(clk), .RN(n4251), .Q(\D_cache/cache[2][146] ) );
  DFFRX1 \D_cache/cache_reg[6][146]  ( .D(\D_cache/n622 ), .CK(clk), .RN(n4251), .Q(\D_cache/cache[6][146] ) );
  DFFRX1 \D_cache/cache_reg[2][147]  ( .D(\D_cache/n618 ), .CK(clk), .RN(n4252), .Q(\D_cache/cache[2][147] ) );
  DFFRX1 \D_cache/cache_reg[6][147]  ( .D(\D_cache/n614 ), .CK(clk), .RN(n4252), .Q(\D_cache/cache[6][147] ) );
  DFFRX1 \D_cache/cache_reg[2][148]  ( .D(\D_cache/n610 ), .CK(clk), .RN(n4252), .Q(\D_cache/cache[2][148] ) );
  DFFRX1 \D_cache/cache_reg[6][148]  ( .D(\D_cache/n606 ), .CK(clk), .RN(n4253), .Q(\D_cache/cache[6][148] ) );
  DFFRX1 \D_cache/cache_reg[2][150]  ( .D(\D_cache/n594 ), .CK(clk), .RN(n4254), .Q(\D_cache/cache[2][150] ) );
  DFFRX1 \D_cache/cache_reg[6][150]  ( .D(\D_cache/n590 ), .CK(clk), .RN(n4254), .Q(\D_cache/cache[6][150] ) );
  DFFRX1 \D_cache/cache_reg[2][151]  ( .D(\D_cache/n586 ), .CK(clk), .RN(n4254), .Q(\D_cache/cache[2][151] ) );
  DFFRX1 \D_cache/cache_reg[2][152]  ( .D(\D_cache/n578 ), .CK(clk), .RN(n4255), .Q(\D_cache/cache[2][152] ) );
  DFFRX1 \D_cache/cache_reg[6][152]  ( .D(\D_cache/n574 ), .CK(clk), .RN(n4255), .Q(\D_cache/cache[6][152] ) );
  DFFRX1 \I_cache/cache_reg[0][128]  ( .D(n9140), .CK(clk), .RN(n4342), .Q(
        \I_cache/cache[0][128] ), .QN(n969) );
  DFFRX1 \I_cache/cache_reg[1][128]  ( .D(n9139), .CK(clk), .RN(n4342), .Q(
        \I_cache/cache[1][128] ), .QN(n80) );
  DFFRX1 \I_cache/cache_reg[2][128]  ( .D(n9138), .CK(clk), .RN(n4342), .Q(
        \I_cache/cache[2][128] ), .QN(n158) );
  DFFRX1 \I_cache/cache_reg[3][128]  ( .D(n9137), .CK(clk), .RN(n4342), .Q(
        \I_cache/cache[3][128] ), .QN(n1049) );
  DFFRX1 \I_cache/cache_reg[4][128]  ( .D(n9136), .CK(clk), .RN(n4343), .Q(
        \I_cache/cache[4][128] ), .QN(n170) );
  DFFRX1 \I_cache/cache_reg[5][128]  ( .D(n9135), .CK(clk), .RN(n4343), .Q(
        \I_cache/cache[5][128] ), .QN(n1067) );
  DFFRX1 \I_cache/cache_reg[6][128]  ( .D(n9134), .CK(clk), .RN(n4343), .Q(
        \I_cache/cache[6][128] ), .QN(n129) );
  DFFRX1 \I_cache/cache_reg[0][129]  ( .D(n9132), .CK(clk), .RN(n4343), .Q(
        \I_cache/cache[0][129] ), .QN(n155) );
  DFFRX1 \I_cache/cache_reg[1][129]  ( .D(n9131), .CK(clk), .RN(n4343), .Q(
        \I_cache/cache[1][129] ), .QN(n1046) );
  DFFRX1 \I_cache/cache_reg[2][129]  ( .D(n9130), .CK(clk), .RN(n4343), .Q(
        \I_cache/cache[2][129] ), .QN(n136) );
  DFFRX1 \I_cache/cache_reg[3][129]  ( .D(n9129), .CK(clk), .RN(n4343), .Q(
        \I_cache/cache[3][129] ), .QN(n1026) );
  DFFRX1 \I_cache/cache_reg[4][129]  ( .D(n9128), .CK(clk), .RN(n4343), .Q(
        \I_cache/cache[4][129] ), .QN(n998) );
  DFFRX1 \I_cache/cache_reg[5][129]  ( .D(n9127), .CK(clk), .RN(n4343), .Q(
        \I_cache/cache[5][129] ), .QN(n110) );
  DFFRX1 \I_cache/cache_reg[6][129]  ( .D(n9126), .CK(clk), .RN(n4343), .Q(
        \I_cache/cache[6][129] ), .QN(n135) );
  DFFRX1 \I_cache/cache_reg[7][129]  ( .D(n9125), .CK(clk), .RN(n4343), .Q(
        \I_cache/cache[7][129] ), .QN(n1025) );
  DFFRX1 \I_cache/cache_reg[0][130]  ( .D(n9124), .CK(clk), .RN(n4343), .Q(
        \I_cache/cache[0][130] ), .QN(n1006) );
  DFFRX1 \I_cache/cache_reg[1][130]  ( .D(n9123), .CK(clk), .RN(n4344), .Q(
        \I_cache/cache[1][130] ), .QN(n118) );
  DFFRX1 \I_cache/cache_reg[2][130]  ( .D(n9122), .CK(clk), .RN(n4344), .Q(
        \I_cache/cache[2][130] ), .QN(n982) );
  DFFRX1 \I_cache/cache_reg[3][130]  ( .D(n9121), .CK(clk), .RN(n4344), .Q(
        \I_cache/cache[3][130] ), .QN(n94) );
  DFFRX1 \I_cache/cache_reg[4][130]  ( .D(n9120), .CK(clk), .RN(n4344), .Q(
        \I_cache/cache[4][130] ), .QN(n995) );
  DFFRX1 \I_cache/cache_reg[5][130]  ( .D(n9119), .CK(clk), .RN(n4344), .Q(
        \I_cache/cache[5][130] ), .QN(n107) );
  DFFRX1 \I_cache/cache_reg[6][130]  ( .D(n9118), .CK(clk), .RN(n4344), .Q(
        \I_cache/cache[6][130] ), .QN(n981) );
  DFFRX1 \I_cache/cache_reg[7][130]  ( .D(n9117), .CK(clk), .RN(n4344), .Q(
        \I_cache/cache[7][130] ), .QN(n93) );
  DFFRX1 \I_cache/cache_reg[0][131]  ( .D(n9116), .CK(clk), .RN(n4344), .Q(
        \I_cache/cache[0][131] ), .QN(n1007) );
  DFFRX1 \I_cache/cache_reg[1][131]  ( .D(n9115), .CK(clk), .RN(n4344), .Q(
        \I_cache/cache[1][131] ), .QN(n119) );
  DFFRX1 \I_cache/cache_reg[2][131]  ( .D(n9114), .CK(clk), .RN(n4344), .Q(
        \I_cache/cache[2][131] ), .QN(n980) );
  DFFRX1 \I_cache/cache_reg[3][131]  ( .D(n9113), .CK(clk), .RN(n4344), .Q(
        \I_cache/cache[3][131] ), .QN(n92) );
  DFFRX1 \I_cache/cache_reg[4][131]  ( .D(n9112), .CK(clk), .RN(n4344), .Q(
        \I_cache/cache[4][131] ), .QN(n996) );
  DFFRX1 \I_cache/cache_reg[5][131]  ( .D(n9111), .CK(clk), .RN(n4345), .Q(
        \I_cache/cache[5][131] ), .QN(n108) );
  DFFRX1 \I_cache/cache_reg[6][131]  ( .D(n9110), .CK(clk), .RN(n4345), .Q(
        \I_cache/cache[6][131] ), .QN(n979) );
  DFFRX1 \I_cache/cache_reg[7][131]  ( .D(n9109), .CK(clk), .RN(n4345), .Q(
        \I_cache/cache[7][131] ), .QN(n91) );
  DFFRX1 \I_cache/cache_reg[0][132]  ( .D(n9108), .CK(clk), .RN(n4345), .Q(
        \I_cache/cache[0][132] ), .QN(n985) );
  DFFRX1 \I_cache/cache_reg[1][132]  ( .D(n9107), .CK(clk), .RN(n4345), .Q(
        \I_cache/cache[1][132] ), .QN(n97) );
  DFFRX1 \I_cache/cache_reg[2][132]  ( .D(n9106), .CK(clk), .RN(n4345), .Q(
        \I_cache/cache[2][132] ), .QN(n983) );
  DFFRX1 \I_cache/cache_reg[3][132]  ( .D(n9105), .CK(clk), .RN(n4345), .Q(
        \I_cache/cache[3][132] ), .QN(n95) );
  DFFRX1 \I_cache/cache_reg[4][132]  ( .D(n9104), .CK(clk), .RN(n4345), .Q(
        \I_cache/cache[4][132] ), .QN(n1001) );
  DFFRX1 \I_cache/cache_reg[5][132]  ( .D(n9103), .CK(clk), .RN(n4345), .Q(
        \I_cache/cache[5][132] ), .QN(n113) );
  DFFRX1 \I_cache/cache_reg[6][132]  ( .D(n9102), .CK(clk), .RN(n4345), .Q(
        \I_cache/cache[6][132] ), .QN(n984) );
  DFFRX1 \I_cache/cache_reg[7][132]  ( .D(n9101), .CK(clk), .RN(n4345), .Q(
        \I_cache/cache[7][132] ), .QN(n96) );
  DFFRX1 \I_cache/cache_reg[0][133]  ( .D(n9100), .CK(clk), .RN(n4345), .Q(
        \I_cache/cache[0][133] ), .QN(n988) );
  DFFRX1 \I_cache/cache_reg[1][133]  ( .D(n9099), .CK(clk), .RN(n4346), .Q(
        \I_cache/cache[1][133] ), .QN(n100) );
  DFFRX1 \I_cache/cache_reg[2][133]  ( .D(n9098), .CK(clk), .RN(n4346), .Q(
        \I_cache/cache[2][133] ), .QN(n986) );
  DFFRX1 \I_cache/cache_reg[3][133]  ( .D(n9097), .CK(clk), .RN(n4346), .Q(
        \I_cache/cache[3][133] ), .QN(n98) );
  DFFRX1 \I_cache/cache_reg[4][133]  ( .D(n9096), .CK(clk), .RN(n4346), .Q(
        \I_cache/cache[4][133] ), .QN(n1003) );
  DFFRX1 \I_cache/cache_reg[5][133]  ( .D(n9095), .CK(clk), .RN(n4346), .Q(
        \I_cache/cache[5][133] ), .QN(n115) );
  DFFRX1 \I_cache/cache_reg[6][133]  ( .D(n9094), .CK(clk), .RN(n4346), .Q(
        \I_cache/cache[6][133] ), .QN(n987) );
  DFFRX1 \I_cache/cache_reg[7][133]  ( .D(n9093), .CK(clk), .RN(n4346), .Q(
        \I_cache/cache[7][133] ), .QN(n99) );
  DFFRX1 \I_cache/cache_reg[0][134]  ( .D(n9092), .CK(clk), .RN(n4346), .Q(
        \I_cache/cache[0][134] ), .QN(n991) );
  DFFRX1 \I_cache/cache_reg[1][134]  ( .D(n9091), .CK(clk), .RN(n4346), .Q(
        \I_cache/cache[1][134] ), .QN(n103) );
  DFFRX1 \I_cache/cache_reg[2][134]  ( .D(n9090), .CK(clk), .RN(n4346), .Q(
        \I_cache/cache[2][134] ), .QN(n989) );
  DFFRX1 \I_cache/cache_reg[3][134]  ( .D(n9089), .CK(clk), .RN(n4346), .Q(
        \I_cache/cache[3][134] ), .QN(n101) );
  DFFRX1 \I_cache/cache_reg[4][134]  ( .D(n9088), .CK(clk), .RN(n4346), .Q(
        \I_cache/cache[4][134] ), .QN(n1004) );
  DFFRX1 \I_cache/cache_reg[5][134]  ( .D(n9087), .CK(clk), .RN(n4347), .Q(
        \I_cache/cache[5][134] ), .QN(n116) );
  DFFRX1 \I_cache/cache_reg[6][134]  ( .D(n9086), .CK(clk), .RN(n4347), .Q(
        \I_cache/cache[6][134] ), .QN(n990) );
  DFFRX1 \I_cache/cache_reg[7][134]  ( .D(n9085), .CK(clk), .RN(n4347), .Q(
        \I_cache/cache[7][134] ), .QN(n102) );
  DFFRX1 \I_cache/cache_reg[0][135]  ( .D(n9084), .CK(clk), .RN(n4347), .Q(
        \I_cache/cache[0][135] ), .QN(n150) );
  DFFRX1 \I_cache/cache_reg[1][135]  ( .D(n9083), .CK(clk), .RN(n4347), .Q(
        \I_cache/cache[1][135] ), .QN(n1041) );
  DFFRX1 \I_cache/cache_reg[2][135]  ( .D(n9082), .CK(clk), .RN(n4347), .Q(
        \I_cache/cache[2][135] ), .QN(n149) );
  DFFRX1 \I_cache/cache_reg[3][135]  ( .D(n9081), .CK(clk), .RN(n4347), .Q(
        \I_cache/cache[3][135] ), .QN(n1040) );
  DFFRX1 \I_cache/cache_reg[4][135]  ( .D(n9080), .CK(clk), .RN(n4347), .Q(
        \I_cache/cache[4][135] ), .QN(n163) );
  DFFRX1 \I_cache/cache_reg[5][135]  ( .D(n9079), .CK(clk), .RN(n4347), .Q(
        \I_cache/cache[5][135] ), .QN(n1053) );
  DFFRX1 \I_cache/cache_reg[6][135]  ( .D(n9078), .CK(clk), .RN(n4347), .Q(
        \I_cache/cache[6][135] ), .QN(n148) );
  DFFRX1 \I_cache/cache_reg[7][135]  ( .D(n9077), .CK(clk), .RN(n4347), .Q(
        \I_cache/cache[7][135] ), .QN(n1039) );
  DFFRX1 \I_cache/cache_reg[0][136]  ( .D(n9076), .CK(clk), .RN(n4347), .Q(
        \I_cache/cache[0][136] ), .QN(n1056) );
  DFFRX1 \I_cache/cache_reg[1][136]  ( .D(n9075), .CK(clk), .RN(n4348), .Q(
        \I_cache/cache[1][136] ), .QN(n1057) );
  DFFRX1 \I_cache/cache_reg[2][136]  ( .D(n9074), .CK(clk), .RN(n4348), .Q(
        \I_cache/cache[2][136] ), .QN(n145) );
  DFFRX1 \I_cache/cache_reg[3][136]  ( .D(n9073), .CK(clk), .RN(n4348), .Q(
        \I_cache/cache[3][136] ), .QN(n1036) );
  DFFRX1 \I_cache/cache_reg[4][136]  ( .D(n9072), .CK(clk), .RN(n4348), .Q(
        \I_cache/cache[4][136] ), .QN(n144) );
  DFFRX1 \I_cache/cache_reg[5][136]  ( .D(n9071), .CK(clk), .RN(n4348), .Q(
        \I_cache/cache[5][136] ), .QN(n1035) );
  DFFRX1 \I_cache/cache_reg[6][136]  ( .D(n9070), .CK(clk), .RN(n4348), .Q(
        \I_cache/cache[6][136] ), .QN(n1058) );
  DFFRX1 \I_cache/cache_reg[7][136]  ( .D(n9069), .CK(clk), .RN(n4348), .Q(
        \I_cache/cache[7][136] ), .QN(n1059) );
  DFFRX1 \I_cache/cache_reg[0][137]  ( .D(n9068), .CK(clk), .RN(n4348), .Q(
        \I_cache/cache[0][137] ), .QN(n147) );
  DFFRX1 \I_cache/cache_reg[1][137]  ( .D(n9067), .CK(clk), .RN(n4348), .Q(
        \I_cache/cache[1][137] ), .QN(n1038) );
  DFFRX1 \I_cache/cache_reg[2][137]  ( .D(n9066), .CK(clk), .RN(n4348), .Q(
        \I_cache/cache[2][137] ), .QN(n146) );
  DFFRX1 \I_cache/cache_reg[3][137]  ( .D(n9065), .CK(clk), .RN(n4348), .Q(
        \I_cache/cache[3][137] ), .QN(n1037) );
  DFFRX1 \I_cache/cache_reg[4][137]  ( .D(n9064), .CK(clk), .RN(n4348), .Q(
        \I_cache/cache[4][137] ), .QN(n974) );
  DFFRX1 \I_cache/cache_reg[5][137]  ( .D(n9063), .CK(clk), .RN(n4349), .Q(
        \I_cache/cache[5][137] ), .QN(n86) );
  DFFRX1 \I_cache/cache_reg[6][137]  ( .D(n9062), .CK(clk), .RN(n4349), .Q(
        \I_cache/cache[6][137] ), .QN(n1055) );
  DFFRX1 \I_cache/cache_reg[7][137]  ( .D(n9061), .CK(clk), .RN(n4349), .Q(
        \I_cache/cache[7][137] ), .QN(n1066) );
  DFFRX1 \I_cache/cache_reg[0][138]  ( .D(n9060), .CK(clk), .RN(n4349), .Q(
        \I_cache/cache[0][138] ), .QN(n978) );
  DFFRX1 \I_cache/cache_reg[1][138]  ( .D(n9059), .CK(clk), .RN(n4349), .Q(
        \I_cache/cache[1][138] ), .QN(n90) );
  DFFRX1 \I_cache/cache_reg[2][138]  ( .D(n9058), .CK(clk), .RN(n4349), .Q(
        \I_cache/cache[2][138] ), .QN(n976) );
  DFFRX1 \I_cache/cache_reg[3][138]  ( .D(n9057), .CK(clk), .RN(n4349), .Q(
        \I_cache/cache[3][138] ), .QN(n88) );
  DFFRX1 \I_cache/cache_reg[4][138]  ( .D(n9056), .CK(clk), .RN(n4349), .Q(
        \I_cache/cache[4][138] ), .QN(n1002) );
  DFFRX1 \I_cache/cache_reg[5][138]  ( .D(n9055), .CK(clk), .RN(n4349), .Q(
        \I_cache/cache[5][138] ), .QN(n114) );
  DFFRX1 \I_cache/cache_reg[6][138]  ( .D(n9054), .CK(clk), .RN(n4349), .Q(
        \I_cache/cache[6][138] ), .QN(n977) );
  DFFRX1 \I_cache/cache_reg[7][138]  ( .D(n9053), .CK(clk), .RN(n4349), .Q(
        \I_cache/cache[7][138] ), .QN(n89) );
  DFFRX1 \I_cache/cache_reg[0][139]  ( .D(n9052), .CK(clk), .RN(n4349), .Q(
        \I_cache/cache[0][139] ), .QN(n152) );
  DFFRX1 \I_cache/cache_reg[1][139]  ( .D(n9051), .CK(clk), .RN(n4350), .Q(
        \I_cache/cache[1][139] ), .QN(n1043) );
  DFFRX1 \I_cache/cache_reg[2][139]  ( .D(n9050), .CK(clk), .RN(n4350), .Q(
        \I_cache/cache[2][139] ), .QN(n151) );
  DFFRX1 \I_cache/cache_reg[3][139]  ( .D(n9049), .CK(clk), .RN(n4350), .Q(
        \I_cache/cache[3][139] ), .QN(n1042) );
  DFFRX1 \I_cache/cache_reg[4][139]  ( .D(n9048), .CK(clk), .RN(n4350), .Q(
        \I_cache/cache[4][139] ), .QN(n162) );
  DFFRX1 \I_cache/cache_reg[5][139]  ( .D(n9047), .CK(clk), .RN(n4350), .Q(
        \I_cache/cache[5][139] ), .QN(n1052) );
  DFFRX1 \I_cache/cache_reg[6][139]  ( .D(n9046), .CK(clk), .RN(n4350), .Q(
        \I_cache/cache[6][139] ), .QN(n1031) );
  DFFRX1 \I_cache/cache_reg[7][139]  ( .D(n9045), .CK(clk), .RN(n4350), .Q(
        \I_cache/cache[7][139] ), .QN(n1032) );
  DFFRX1 \I_cache/cache_reg[0][140]  ( .D(n9044), .CK(clk), .RN(n4350), .Q(
        \I_cache/cache[0][140] ), .QN(n160) );
  DFFRX1 \I_cache/cache_reg[1][140]  ( .D(n9043), .CK(clk), .RN(n4350), .Q(
        \I_cache/cache[1][140] ), .QN(n1051) );
  DFFRX1 \I_cache/cache_reg[2][140]  ( .D(n9042), .CK(clk), .RN(n4350), .Q(
        \I_cache/cache[2][140] ), .QN(n159) );
  DFFRX1 \I_cache/cache_reg[3][140]  ( .D(n9041), .CK(clk), .RN(n4350), .Q(
        \I_cache/cache[3][140] ), .QN(n1050) );
  DFFRX1 \I_cache/cache_reg[4][140]  ( .D(n9040), .CK(clk), .RN(n4350), .Q(
        \I_cache/cache[4][140] ), .QN(n975) );
  DFFRX1 \I_cache/cache_reg[5][140]  ( .D(n9039), .CK(clk), .RN(n4351), .Q(
        \I_cache/cache[5][140] ), .QN(n87) );
  DFFRX1 \I_cache/cache_reg[6][140]  ( .D(n9038), .CK(clk), .RN(n4351), .Q(
        \I_cache/cache[6][140] ), .QN(n1060) );
  DFFRX1 \I_cache/cache_reg[7][140]  ( .D(n9037), .CK(clk), .RN(n4351), .Q(
        \I_cache/cache[7][140] ), .QN(n1033) );
  DFFRX1 \I_cache/cache_reg[0][141]  ( .D(n9036), .CK(clk), .RN(n4351), .Q(
        \I_cache/cache[0][141] ), .QN(n971) );
  DFFRX1 \I_cache/cache_reg[1][141]  ( .D(n9035), .CK(clk), .RN(n4351), .Q(
        \I_cache/cache[1][141] ), .QN(n82) );
  DFFRX1 \I_cache/cache_reg[2][141]  ( .D(n9034), .CK(clk), .RN(n4351), .Q(
        \I_cache/cache[2][141] ), .QN(n138) );
  DFFRX1 \I_cache/cache_reg[3][141]  ( .D(n9033), .CK(clk), .RN(n4351), .Q(
        \I_cache/cache[3][141] ), .QN(n1028) );
  DFFRX1 \I_cache/cache_reg[4][141]  ( .D(n9032), .CK(clk), .RN(n4351), .Q(
        \I_cache/cache[4][141] ), .QN(n1000) );
  DFFRX1 \I_cache/cache_reg[5][141]  ( .D(n9031), .CK(clk), .RN(n4351), .Q(
        \I_cache/cache[5][141] ), .QN(n112) );
  DFFRX1 \I_cache/cache_reg[6][141]  ( .D(n9030), .CK(clk), .RN(n4351), .Q(
        \I_cache/cache[6][141] ), .QN(n137) );
  DFFRX1 \I_cache/cache_reg[7][141]  ( .D(n9029), .CK(clk), .RN(n4351), .Q(
        \I_cache/cache[7][141] ), .QN(n1027) );
  DFFRX1 \I_cache/cache_reg[0][142]  ( .D(n9028), .CK(clk), .RN(n4351), .Q(
        \I_cache/cache[0][142] ), .QN(n972) );
  DFFRX1 \I_cache/cache_reg[1][142]  ( .D(n9027), .CK(clk), .RN(n4352), .Q(
        \I_cache/cache[1][142] ), .QN(n83) );
  DFFRX1 \I_cache/cache_reg[2][142]  ( .D(n9026), .CK(clk), .RN(n4352), .Q(
        \I_cache/cache[2][142] ), .QN(n134) );
  DFFRX1 \I_cache/cache_reg[3][142]  ( .D(n9025), .CK(clk), .RN(n4352), .Q(
        \I_cache/cache[3][142] ), .QN(n1023) );
  DFFRX1 \I_cache/cache_reg[4][142]  ( .D(n9024), .CK(clk), .RN(n4352), .Q(
        \I_cache/cache[4][142] ), .QN(n999) );
  DFFRX1 \I_cache/cache_reg[5][142]  ( .D(n9023), .CK(clk), .RN(n4352), .Q(
        \I_cache/cache[5][142] ), .QN(n111) );
  DFFRX1 \I_cache/cache_reg[6][142]  ( .D(n9022), .CK(clk), .RN(n4352), .Q(
        \I_cache/cache[6][142] ), .QN(n133) );
  DFFRX1 \I_cache/cache_reg[7][142]  ( .D(n9021), .CK(clk), .RN(n4352), .Q(
        \I_cache/cache[7][142] ), .QN(n1022) );
  DFFRX1 \I_cache/cache_reg[0][143]  ( .D(n9020), .CK(clk), .RN(n4352), .Q(
        \I_cache/cache[0][143] ), .QN(n970) );
  DFFRX1 \I_cache/cache_reg[1][143]  ( .D(n9019), .CK(clk), .RN(n4352), .Q(
        \I_cache/cache[1][143] ), .QN(n81) );
  DFFRX1 \I_cache/cache_reg[2][143]  ( .D(n9018), .CK(clk), .RN(n4352), .Q(
        \I_cache/cache[2][143] ), .QN(n132) );
  DFFRX1 \I_cache/cache_reg[3][143]  ( .D(n9017), .CK(clk), .RN(n4352), .Q(
        \I_cache/cache[3][143] ), .QN(n1021) );
  DFFRX1 \I_cache/cache_reg[4][143]  ( .D(n9016), .CK(clk), .RN(n4352), .Q(
        \I_cache/cache[4][143] ), .QN(n997) );
  DFFRX1 \I_cache/cache_reg[5][143]  ( .D(n9015), .CK(clk), .RN(n4353), .Q(
        \I_cache/cache[5][143] ), .QN(n109) );
  DFFRX1 \I_cache/cache_reg[6][143]  ( .D(n9014), .CK(clk), .RN(n4353), .Q(
        \I_cache/cache[6][143] ), .QN(n131) );
  DFFRX1 \I_cache/cache_reg[7][143]  ( .D(n9013), .CK(clk), .RN(n4353), .Q(
        \I_cache/cache[7][143] ), .QN(n1020) );
  DFFRX1 \I_cache/cache_reg[0][144]  ( .D(n9012), .CK(clk), .RN(n4353), .Q(
        \I_cache/cache[0][144] ), .QN(n154) );
  DFFRX1 \I_cache/cache_reg[1][144]  ( .D(n9011), .CK(clk), .RN(n4353), .Q(
        \I_cache/cache[1][144] ), .QN(n1045) );
  DFFRX1 \I_cache/cache_reg[2][144]  ( .D(n9010), .CK(clk), .RN(n4353), .Q(
        \I_cache/cache[2][144] ), .QN(n153) );
  DFFRX1 \I_cache/cache_reg[3][144]  ( .D(n9009), .CK(clk), .RN(n4353), .Q(
        \I_cache/cache[3][144] ), .QN(n1044) );
  DFFRX1 \I_cache/cache_reg[4][144]  ( .D(n9008), .CK(clk), .RN(n4353), .Q(
        \I_cache/cache[4][144] ), .QN(n164) );
  DFFRX1 \I_cache/cache_reg[5][144]  ( .D(n9007), .CK(clk), .RN(n4353), .Q(
        \I_cache/cache[5][144] ), .QN(n1054) );
  DFFRX1 \I_cache/cache_reg[6][144]  ( .D(n9006), .CK(clk), .RN(n4353), .Q(
        \I_cache/cache[6][144] ), .QN(n130) );
  DFFRX1 \I_cache/cache_reg[7][144]  ( .D(n9005), .CK(clk), .RN(n4353), .Q(
        \I_cache/cache[7][144] ), .QN(n1019) );
  DFFRX1 \I_cache/cache_reg[0][145]  ( .D(n9004), .CK(clk), .RN(n4353), .Q(
        \I_cache/cache[0][145] ), .QN(n1008) );
  DFFRX1 \I_cache/cache_reg[1][145]  ( .D(n9003), .CK(clk), .RN(n4354), .Q(
        \I_cache/cache[1][145] ), .QN(n120) );
  DFFRX1 \I_cache/cache_reg[2][145]  ( .D(n9002), .CK(clk), .RN(n4354), .Q(
        \I_cache/cache[2][145] ), .QN(n1073) );
  DFFRX1 \I_cache/cache_reg[3][145]  ( .D(n9001), .CK(clk), .RN(n4354), .Q(
        \I_cache/cache[3][145] ), .QN(n84) );
  DFFRX1 \I_cache/cache_reg[4][145]  ( .D(n9000), .CK(clk), .RN(n4354), .Q(
        \I_cache/cache[4][145] ), .QN(n1080) );
  DFFRX1 \I_cache/cache_reg[5][145]  ( .D(n8999), .CK(clk), .RN(n4354), .Q(
        \I_cache/cache[5][145] ), .QN(n168) );
  DFFRX1 \I_cache/cache_reg[6][145]  ( .D(n8998), .CK(clk), .RN(n4354), .Q(
        \I_cache/cache[6][145] ), .QN(n1009) );
  DFFRX1 \I_cache/cache_reg[7][145]  ( .D(n8997), .CK(clk), .RN(n4354), .Q(
        \I_cache/cache[7][145] ), .QN(n121) );
  DFFRX1 \I_cache/cache_reg[0][146]  ( .D(n8996), .CK(clk), .RN(n4354), .Q(
        \I_cache/cache[0][146] ), .QN(n994) );
  DFFRX1 \I_cache/cache_reg[1][146]  ( .D(n8995), .CK(clk), .RN(n4354), .Q(
        \I_cache/cache[1][146] ), .QN(n106) );
  DFFRX1 \I_cache/cache_reg[2][146]  ( .D(n8994), .CK(clk), .RN(n4354), .Q(
        \I_cache/cache[2][146] ), .QN(n992) );
  DFFRX1 \I_cache/cache_reg[3][146]  ( .D(n8993), .CK(clk), .RN(n4354), .Q(
        \I_cache/cache[3][146] ), .QN(n104) );
  DFFRX1 \I_cache/cache_reg[4][146]  ( .D(n8992), .CK(clk), .RN(n4354), .Q(
        \I_cache/cache[4][146] ), .QN(n1005) );
  DFFRX1 \I_cache/cache_reg[5][146]  ( .D(n8991), .CK(clk), .RN(n4355), .Q(
        \I_cache/cache[5][146] ), .QN(n117) );
  DFFRX1 \I_cache/cache_reg[6][146]  ( .D(n8990), .CK(clk), .RN(n4355), .Q(
        \I_cache/cache[6][146] ), .QN(n993) );
  DFFRX1 \I_cache/cache_reg[7][146]  ( .D(n8989), .CK(clk), .RN(n4355), .Q(
        \I_cache/cache[7][146] ), .QN(n105) );
  DFFRX1 \I_cache/cache_reg[0][147]  ( .D(n8988), .CK(clk), .RN(n4355), .Q(
        \I_cache/cache[0][147] ), .QN(n1011) );
  DFFRX1 \I_cache/cache_reg[1][147]  ( .D(n8987), .CK(clk), .RN(n4355), .Q(
        \I_cache/cache[1][147] ), .QN(n123) );
  DFFRX1 \I_cache/cache_reg[2][147]  ( .D(n8986), .CK(clk), .RN(n4355), .Q(
        \I_cache/cache[2][147] ), .QN(n1075) );
  DFFRX1 \I_cache/cache_reg[3][147]  ( .D(n8985), .CK(clk), .RN(n4355), .Q(
        \I_cache/cache[3][147] ), .QN(n141) );
  DFFRX1 \I_cache/cache_reg[4][147]  ( .D(n8984), .CK(clk), .RN(n4355), .Q(
        \I_cache/cache[4][147] ), .QN(n1079) );
  DFFRX1 \I_cache/cache_reg[5][147]  ( .D(n8983), .CK(clk), .RN(n4355), .Q(
        \I_cache/cache[5][147] ), .QN(n167) );
  DFFRX1 \I_cache/cache_reg[6][147]  ( .D(n8982), .CK(clk), .RN(n4355), .Q(
        \I_cache/cache[6][147] ), .QN(n142) );
  DFFRX1 \I_cache/cache_reg[7][147]  ( .D(n8981), .CK(clk), .RN(n4355), .Q(
        \I_cache/cache[7][147] ), .QN(n1034) );
  DFFRX1 \I_cache/cache_reg[0][148]  ( .D(n8980), .CK(clk), .RN(n4355), .Q(
        \I_cache/cache[0][148] ), .QN(n1013) );
  DFFRX1 \I_cache/cache_reg[1][148]  ( .D(n8979), .CK(clk), .RN(n4356), .Q(
        \I_cache/cache[1][148] ), .QN(n1061) );
  DFFRX1 \I_cache/cache_reg[2][148]  ( .D(n8978), .CK(clk), .RN(n4356), .Q(
        \I_cache/cache[2][148] ), .QN(n156) );
  DFFRX1 \I_cache/cache_reg[3][148]  ( .D(n8977), .CK(clk), .RN(n4356), .Q(
        \I_cache/cache[3][148] ), .QN(n1047) );
  DFFRX1 \I_cache/cache_reg[4][148]  ( .D(n8976), .CK(clk), .RN(n4356), .Q(
        \I_cache/cache[4][148] ), .QN(n143) );
  DFFRX1 \I_cache/cache_reg[5][148]  ( .D(n8975), .CK(clk), .RN(n4356), .Q(
        \I_cache/cache[5][148] ), .QN(n1024) );
  DFFRX1 \I_cache/cache_reg[6][148]  ( .D(n8974), .CK(clk), .RN(n4356), .Q(
        \I_cache/cache[6][148] ), .QN(n139) );
  DFFRX1 \I_cache/cache_reg[7][148]  ( .D(n8973), .CK(clk), .RN(n4356), .Q(
        \I_cache/cache[7][148] ), .QN(n1029) );
  DFFRX1 \I_cache/cache_reg[0][149]  ( .D(n8972), .CK(clk), .RN(n4356), .Q(
        \I_cache/cache[0][149] ), .QN(n1012) );
  DFFRX1 \I_cache/cache_reg[1][149]  ( .D(n8971), .CK(clk), .RN(n4356), .Q(
        \I_cache/cache[1][149] ), .QN(n124) );
  DFFRX1 \I_cache/cache_reg[2][149]  ( .D(n8970), .CK(clk), .RN(n4356), .Q(
        \I_cache/cache[2][149] ), .QN(n1076) );
  DFFRX1 \I_cache/cache_reg[3][149]  ( .D(n8969), .CK(clk), .RN(n4356), .Q(
        \I_cache/cache[3][149] ), .QN(n161) );
  DFFRX1 \I_cache/cache_reg[4][149]  ( .D(n8968), .CK(clk), .RN(n4356), .Q(
        \I_cache/cache[4][149] ), .QN(n1078) );
  DFFRX1 \I_cache/cache_reg[5][149]  ( .D(n8967), .CK(clk), .RN(n4357), .Q(
        \I_cache/cache[5][149] ), .QN(n166) );
  DFFRX1 \I_cache/cache_reg[6][149]  ( .D(n8966), .CK(clk), .RN(n4357), .Q(
        \I_cache/cache[6][149] ), .QN(n125) );
  DFFRX1 \I_cache/cache_reg[7][149]  ( .D(n8965), .CK(clk), .RN(n4357), .Q(
        \I_cache/cache[7][149] ), .QN(n1014) );
  DFFRX1 \I_cache/cache_reg[0][150]  ( .D(n8964), .CK(clk), .RN(n4357), .Q(
        \I_cache/cache[0][150] ), .QN(n1010) );
  DFFRX1 \I_cache/cache_reg[1][150]  ( .D(n8963), .CK(clk), .RN(n4357), .Q(
        \I_cache/cache[1][150] ), .QN(n122) );
  DFFRX1 \I_cache/cache_reg[2][150]  ( .D(n8962), .CK(clk), .RN(n4357), .Q(
        \I_cache/cache[2][150] ), .QN(n1077) );
  DFFRX1 \I_cache/cache_reg[3][150]  ( .D(n8961), .CK(clk), .RN(n4357), .Q(
        \I_cache/cache[3][150] ), .QN(n165) );
  DFFRX1 \I_cache/cache_reg[4][150]  ( .D(n8960), .CK(clk), .RN(n4357), .Q(
        \I_cache/cache[4][150] ), .QN(n1081) );
  DFFRX1 \I_cache/cache_reg[5][150]  ( .D(n8959), .CK(clk), .RN(n4357), .Q(
        \I_cache/cache[5][150] ), .QN(n169) );
  DFFRX1 \I_cache/cache_reg[6][150]  ( .D(n8958), .CK(clk), .RN(n4357), .Q(
        \I_cache/cache[6][150] ), .QN(n973) );
  DFFRX1 \I_cache/cache_reg[7][150]  ( .D(n8957), .CK(clk), .RN(n4357), .Q(
        \I_cache/cache[7][150] ), .QN(n85) );
  DFFRX1 \I_cache/cache_reg[0][151]  ( .D(n8956), .CK(clk), .RN(n4357), .Q(
        \I_cache/cache[0][151] ), .QN(n127) );
  DFFRX1 \I_cache/cache_reg[1][151]  ( .D(n8955), .CK(clk), .RN(n4358), .Q(
        \I_cache/cache[1][151] ), .QN(n1016) );
  DFFRX1 \I_cache/cache_reg[2][151]  ( .D(n8954), .CK(clk), .RN(n4358), .Q(
        \I_cache/cache[2][151] ), .QN(n126) );
  DFFRX1 \I_cache/cache_reg[3][151]  ( .D(n8953), .CK(clk), .RN(n4358), .Q(
        \I_cache/cache[3][151] ), .QN(n1015) );
  DFFRX1 \I_cache/cache_reg[4][151]  ( .D(n8952), .CK(clk), .RN(n4358), .Q(
        \I_cache/cache[4][151] ), .QN(n171) );
  DFFRX1 \I_cache/cache_reg[5][151]  ( .D(n8951), .CK(clk), .RN(n4358), .Q(
        \I_cache/cache[5][151] ), .QN(n1068) );
  DFFRX1 \I_cache/cache_reg[6][151]  ( .D(n8950), .CK(clk), .RN(n4358), .Q(
        \I_cache/cache[6][151] ), .QN(n128) );
  DFFRX1 \I_cache/cache_reg[7][151]  ( .D(n8949), .CK(clk), .RN(n4358), .Q(
        \I_cache/cache[7][151] ), .QN(n1017) );
  DFFRX1 \I_cache/cache_reg[0][152]  ( .D(n8948), .CK(clk), .RN(n4358), .Q(
        \I_cache/cache[0][152] ), .QN(n1064) );
  DFFRX1 \I_cache/cache_reg[1][152]  ( .D(n8947), .CK(clk), .RN(n4358), .Q(
        \I_cache/cache[1][152] ), .QN(n1065) );
  DFFRX1 \I_cache/cache_reg[2][152]  ( .D(n8946), .CK(clk), .RN(n4358), .Q(
        \I_cache/cache[2][152] ), .QN(n1062) );
  DFFRX1 \I_cache/cache_reg[3][152]  ( .D(n8945), .CK(clk), .RN(n4358), .Q(
        \I_cache/cache[3][152] ), .QN(n1063) );
  DFFRX1 \I_cache/cache_reg[4][152]  ( .D(n8944), .CK(clk), .RN(n4358), .Q(
        \I_cache/cache[4][152] ), .QN(n157) );
  DFFRX1 \I_cache/cache_reg[5][152]  ( .D(n8943), .CK(clk), .RN(n4359), .Q(
        \I_cache/cache[5][152] ), .QN(n1048) );
  DFFRX1 \I_cache/cache_reg[6][152]  ( .D(n8942), .CK(clk), .RN(n4359), .Q(
        \I_cache/cache[6][152] ), .QN(n140) );
  DFFRX1 \I_cache/cache_reg[7][152]  ( .D(n8941), .CK(clk), .RN(n4359), .Q(
        \I_cache/cache[7][152] ), .QN(n1030) );
  DFFRX1 \I_cache/cache_reg[7][128]  ( .D(n9133), .CK(clk), .RN(n4359), .Q(
        \I_cache/cache[7][128] ), .QN(n1018) );
  DFFRX1 \i_MIPS/ID_EX_reg[104]  ( .D(\i_MIPS/n481 ), .CK(clk), .RN(n4056), 
        .Q(\i_MIPS/ID_EX[104] ), .QN(n2884) );
  DFFRX1 \i_MIPS/ID_EX_reg[103]  ( .D(\i_MIPS/n482 ), .CK(clk), .RN(n4056), 
        .Q(\i_MIPS/ID_EX[103] ) );
  DFFRX1 \i_MIPS/ID_EX_reg[102]  ( .D(\i_MIPS/n483 ), .CK(clk), .RN(n4056), 
        .Q(\i_MIPS/ID_EX[102] ) );
  DFFRX1 \i_MIPS/ID_EX_reg[101]  ( .D(\i_MIPS/n484 ), .CK(clk), .RN(n4056), 
        .Q(\i_MIPS/ID_EX[101] ) );
  DFFRX1 \i_MIPS/ID_EX_reg[100]  ( .D(\i_MIPS/n485 ), .CK(clk), .RN(n4056), 
        .Q(\i_MIPS/ID_EX[100] ) );
  DFFRX1 \i_MIPS/ID_EX_reg[98]  ( .D(\i_MIPS/n487 ), .CK(clk), .RN(n4056), .Q(
        \i_MIPS/ID_EX[98] ) );
  DFFRX1 \i_MIPS/ID_EX_reg[97]  ( .D(\i_MIPS/n488 ), .CK(clk), .RN(n4057), .Q(
        \i_MIPS/ID_EX[97] ) );
  DFFRX1 \i_MIPS/ID_EX_reg[96]  ( .D(\i_MIPS/n489 ), .CK(clk), .RN(n4057), .Q(
        \i_MIPS/ID_EX[96] ) );
  DFFRX1 \i_MIPS/ID_EX_reg[95]  ( .D(\i_MIPS/n490 ), .CK(clk), .RN(n4057), .Q(
        \i_MIPS/ID_EX[95] ) );
  DFFRX1 \i_MIPS/ID_EX_reg[94]  ( .D(\i_MIPS/n491 ), .CK(clk), .RN(n4057), .Q(
        \i_MIPS/ID_EX[94] ) );
  DFFRX1 \i_MIPS/ID_EX_reg[93]  ( .D(\i_MIPS/n492 ), .CK(clk), .RN(n4057), .Q(
        \i_MIPS/ID_EX[93] ) );
  DFFRX1 \i_MIPS/ID_EX_reg[92]  ( .D(\i_MIPS/n493 ), .CK(clk), .RN(n4057), .Q(
        \i_MIPS/ID_EX[92] ) );
  DFFRX1 \i_MIPS/ID_EX_reg[91]  ( .D(\i_MIPS/n494 ), .CK(clk), .RN(n4057), .Q(
        \i_MIPS/ID_EX[91] ) );
  DFFRX1 \i_MIPS/ID_EX_reg[90]  ( .D(\i_MIPS/n495 ), .CK(clk), .RN(n4057), .Q(
        \i_MIPS/ID_EX[90] ) );
  DFFRX1 \i_MIPS/ID_EX_reg[105]  ( .D(\i_MIPS/n518 ), .CK(clk), .RN(n4061), 
        .Q(\i_MIPS/ID_EX[105] ), .QN(\i_MIPS/n323 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[107]  ( .D(\i_MIPS/n520 ), .CK(clk), .RN(n4061), 
        .Q(\i_MIPS/ID_EX[107] ), .QN(\i_MIPS/n327 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[114]  ( .D(\i_MIPS/n516 ), .CK(clk), .RN(n4060), 
        .Q(\i_MIPS/ID_EX[114] ), .QN(\i_MIPS/n319 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[115]  ( .D(\i_MIPS/n517 ), .CK(clk), .RN(n4061), 
        .Q(\i_MIPS/ID_EX[115] ), .QN(\i_MIPS/n321 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[113]  ( .D(\i_MIPS/n515 ), .CK(clk), .RN(n4060), 
        .Q(\i_MIPS/ID_EX[113] ), .QN(\i_MIPS/n317 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[88]  ( .D(\i_MIPS/n497 ), .CK(clk), .RN(n4057), .Q(
        \i_MIPS/ID_EX[88] ), .QN(n2889) );
  DFFRX1 \i_MIPS/ID_EX_reg[86]  ( .D(\i_MIPS/n499 ), .CK(clk), .RN(n4057), .Q(
        \i_MIPS/ID_EX[86] ), .QN(n2993) );
  DFFRX1 \i_MIPS/ID_EX_reg[84]  ( .D(\i_MIPS/n501 ), .CK(clk), .RN(n4058), .Q(
        \i_MIPS/ID_EX[84] ), .QN(n2991) );
  DFFRX1 \i_MIPS/IF_ID_reg[52]  ( .D(\i_MIPS/N75 ), .CK(clk), .RN(n4061), .Q(
        \i_MIPS/IR_ID[20] ), .QN(\i_MIPS/n320 ) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[23]  ( .D(\i_MIPS/PC/n57 ), .CK(clk), .RN(n4067), 
        .Q(ICACHE_addr[21]), .QN(\i_MIPS/PC/n25 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[17]  ( .D(\i_MIPS/n554 ), .CK(clk), .RN(n4065), .Q(
        \i_MIPS/ALUin1[8] ), .QN(\i_MIPS/n363 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[28]  ( .D(\i_MIPS/n543 ), .CK(clk), .RN(n4064), .Q(
        \i_MIPS/ALUin1[19] ), .QN(\i_MIPS/n352 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[21]  ( .D(\i_MIPS/n550 ), .CK(clk), .RN(n4064), .Q(
        \i_MIPS/ALUin1[12] ), .QN(\i_MIPS/n359 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[33]  ( .D(\i_MIPS/n538 ), .CK(clk), .RN(n4063), .Q(
        \i_MIPS/ALUin1[24] ), .QN(\i_MIPS/n347 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[32]  ( .D(\i_MIPS/n539 ), .CK(clk), .RN(n4063), .Q(
        \i_MIPS/ALUin1[23] ), .QN(\i_MIPS/n348 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[31]  ( .D(\i_MIPS/n540 ), .CK(clk), .RN(n4064), .Q(
        \i_MIPS/ALUin1[22] ), .QN(\i_MIPS/n349 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[18]  ( .D(\i_MIPS/n553 ), .CK(clk), .RN(n4065), .Q(
        \i_MIPS/ALUin1[9] ), .QN(\i_MIPS/n362 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[30]  ( .D(\i_MIPS/n541 ), .CK(clk), .RN(n4064), .Q(
        \i_MIPS/ALUin1[21] ), .QN(\i_MIPS/n350 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[19]  ( .D(\i_MIPS/n552 ), .CK(clk), .RN(n4065), .Q(
        \i_MIPS/ALUin1[10] ), .QN(\i_MIPS/n361 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[29]  ( .D(\i_MIPS/n542 ), .CK(clk), .RN(n4064), .Q(
        \i_MIPS/ALUin1[20] ), .QN(\i_MIPS/n351 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[20]  ( .D(\i_MIPS/n551 ), .CK(clk), .RN(n4064), .Q(
        \i_MIPS/ALUin1[11] ), .QN(\i_MIPS/n360 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[40]  ( .D(\i_MIPS/n531 ), .CK(clk), .RN(n4063), .Q(
        \i_MIPS/ALU/N303 ), .QN(\i_MIPS/n340 ) );
  MXI2X1 \D_cache/U2073  ( .A(\D_cache/n1971 ), .B(\D_cache/n1972 ), .S0(n3065), .Y(\D_cache/N97 ) );
  MXI4X1 \D_cache/U2154  ( .A(\D_cache/cache[0][6] ), .B(\D_cache/cache[1][6] ), .C(\D_cache/cache[2][6] ), .D(\D_cache/cache[3][6] ), .S0(n2106), .S1(n2383), 
        .Y(\D_cache/n1809 ) );
  MXI4X1 \D_cache/U2153  ( .A(\D_cache/cache[4][6] ), .B(\D_cache/cache[5][6] ), .C(\D_cache/cache[6][6] ), .D(\D_cache/cache[7][6] ), .S0(n2105), .S1(n2377), 
        .Y(\D_cache/n1810 ) );
  MXI2X1 \D_cache/U1992  ( .A(\D_cache/n1809 ), .B(\D_cache/n1810 ), .S0(n2147), .Y(\D_cache/N178 ) );
  MXI4X1 \D_cache/U2155  ( .A(\D_cache/cache[4][7] ), .B(\D_cache/cache[5][7] ), .C(\D_cache/cache[6][7] ), .D(\D_cache/cache[7][7] ), .S0(n2084), .S1(n2228), 
        .Y(\D_cache/n1812 ) );
  MXI4X1 \D_cache/U2156  ( .A(\D_cache/cache[0][7] ), .B(\D_cache/cache[1][7] ), .C(\D_cache/cache[2][7] ), .D(\D_cache/cache[3][7] ), .S0(n2114), .S1(n2233), 
        .Y(\D_cache/n1811 ) );
  MXI2X1 \D_cache/U1993  ( .A(\D_cache/n1811 ), .B(\D_cache/n1812 ), .S0(n4041), .Y(\D_cache/N177 ) );
  MXI4X1 \D_cache/U2157  ( .A(\D_cache/cache[4][8] ), .B(\D_cache/cache[5][8] ), .C(\D_cache/cache[6][8] ), .D(\D_cache/cache[7][8] ), .S0(n2066), .S1(n2260), 
        .Y(\D_cache/n1814 ) );
  MXI4X1 \D_cache/U2158  ( .A(\D_cache/cache[0][8] ), .B(\D_cache/cache[1][8] ), .C(\D_cache/cache[2][8] ), .D(\D_cache/cache[3][8] ), .S0(n2069), .S1(n2255), 
        .Y(\D_cache/n1813 ) );
  MXI2X1 \D_cache/U1994  ( .A(\D_cache/n1813 ), .B(\D_cache/n1814 ), .S0(n2147), .Y(\D_cache/N176 ) );
  MXI4X1 \D_cache/U2160  ( .A(\D_cache/cache[0][9] ), .B(\D_cache/cache[1][9] ), .C(\D_cache/cache[2][9] ), .D(\D_cache/cache[3][9] ), .S0(n2122), .S1(n2365), 
        .Y(\D_cache/n1815 ) );
  MXI4X1 \D_cache/U2159  ( .A(\D_cache/cache[4][9] ), .B(\D_cache/cache[5][9] ), .C(\D_cache/cache[6][9] ), .D(\D_cache/cache[7][9] ), .S0(n2121), .S1(n2360), 
        .Y(\D_cache/n1816 ) );
  MXI2X1 \D_cache/U1995  ( .A(\D_cache/n1815 ), .B(\D_cache/n1816 ), .S0(n3062), .Y(\D_cache/N175 ) );
  MXI2X1 \D_cache/U1996  ( .A(\D_cache/n1817 ), .B(\D_cache/n1818 ), .S0(n3066), .Y(\D_cache/N174 ) );
  MXI4X1 \D_cache/U2187  ( .A(\D_cache/cache[4][23] ), .B(
        \D_cache/cache[5][23] ), .C(\D_cache/cache[6][23] ), .D(
        \D_cache/cache[7][23] ), .S0(n2133), .S1(n2224), .Y(\D_cache/n1844 )
         );
  MXI4X1 \D_cache/U2188  ( .A(\D_cache/cache[0][23] ), .B(
        \D_cache/cache[1][23] ), .C(\D_cache/cache[2][23] ), .D(
        \D_cache/cache[3][23] ), .S0(n2122), .S1(n2225), .Y(\D_cache/n1843 )
         );
  MXI2X1 \D_cache/U2009  ( .A(\D_cache/n1843 ), .B(\D_cache/n1844 ), .S0(n3067), .Y(\D_cache/N161 ) );
  MXI2X1 \D_cache/U2062  ( .A(\D_cache/n1949 ), .B(\D_cache/n1950 ), .S0(n3066), .Y(\D_cache/N108 ) );
  MXI2X1 \D_cache/U2068  ( .A(\D_cache/n1961 ), .B(\D_cache/n1962 ), .S0(
        DCACHE_addr[4]), .Y(\D_cache/N102 ) );
  MXI2X1 \D_cache/U2089  ( .A(\D_cache/n2003 ), .B(\D_cache/n2004 ), .S0(n3063), .Y(\D_cache/N81 ) );
  MXI4X1 \D_cache/U2333  ( .A(\D_cache/cache[4][96] ), .B(
        \D_cache/cache[5][96] ), .C(\D_cache/cache[6][96] ), .D(
        \D_cache/cache[7][96] ), .S0(n2144), .S1(n2196), .Y(\D_cache/n1990 )
         );
  MXI4X1 \D_cache/U2334  ( .A(\D_cache/cache[0][96] ), .B(
        \D_cache/cache[1][96] ), .C(\D_cache/cache[2][96] ), .D(
        \D_cache/cache[3][96] ), .S0(n2117), .S1(n2197), .Y(\D_cache/n1989 )
         );
  MXI2X1 \D_cache/U2082  ( .A(\D_cache/n1989 ), .B(\D_cache/n1990 ), .S0(n3064), .Y(\D_cache/N88 ) );
  MXI2X1 \D_cache/U2067  ( .A(\D_cache/n1959 ), .B(\D_cache/n1960 ), .S0(n4041), .Y(\D_cache/N103 ) );
  MXI4X1 \D_cache/U2181  ( .A(\D_cache/cache[4][20] ), .B(
        \D_cache/cache[5][20] ), .C(\D_cache/cache[6][20] ), .D(
        \D_cache/cache[7][20] ), .S0(n2076), .S1(n2180), .Y(\D_cache/n1838 )
         );
  MXI4X1 \D_cache/U2182  ( .A(\D_cache/cache[0][20] ), .B(
        \D_cache/cache[1][20] ), .C(\D_cache/cache[2][20] ), .D(
        \D_cache/cache[3][20] ), .S0(n2139), .S1(n2185), .Y(\D_cache/n1837 )
         );
  MXI2X1 \D_cache/U2006  ( .A(\D_cache/n1837 ), .B(\D_cache/n1838 ), .S0(n2147), .Y(\D_cache/N164 ) );
  MXI2X1 \D_cache/U2003  ( .A(\D_cache/n1831 ), .B(\D_cache/n1832 ), .S0(n2146), .Y(\D_cache/N167 ) );
  MXI2X1 \D_cache/U2066  ( .A(\D_cache/n1957 ), .B(\D_cache/n1958 ), .S0(n3064), .Y(\D_cache/N104 ) );
  MXI2X1 \D_cache/U2065  ( .A(\D_cache/n1955 ), .B(\D_cache/n1956 ), .S0(
        DCACHE_addr[4]), .Y(\D_cache/N105 ) );
  MXI2X1 \D_cache/U2002  ( .A(\D_cache/n1829 ), .B(\D_cache/n1830 ), .S0(
        DCACHE_addr[4]), .Y(\D_cache/N168 ) );
  MXI4X1 \D_cache/U2172  ( .A(\D_cache/cache[0][15] ), .B(
        \D_cache/cache[1][15] ), .C(\D_cache/cache[2][15] ), .D(
        \D_cache/cache[3][15] ), .S0(n2140), .S1(n2364), .Y(\D_cache/n1827 )
         );
  MXI4X1 \D_cache/U2171  ( .A(\D_cache/cache[4][15] ), .B(
        \D_cache/cache[5][15] ), .C(\D_cache/cache[6][15] ), .D(
        \D_cache/cache[7][15] ), .S0(n2138), .S1(n2322), .Y(\D_cache/n1828 )
         );
  MXI2X1 \D_cache/U2001  ( .A(\D_cache/n1827 ), .B(\D_cache/n1828 ), .S0(n3065), .Y(\D_cache/N169 ) );
  MXI2X1 \D_cache/U2005  ( .A(\D_cache/n1835 ), .B(\D_cache/n1836 ), .S0(
        DCACHE_addr[4]), .Y(\D_cache/N165 ) );
  MXI2X1 \D_cache/U2083  ( .A(\D_cache/n1991 ), .B(\D_cache/n1992 ), .S0(n3064), .Y(\D_cache/N87 ) );
  MXI2X1 \D_cache/U2088  ( .A(\D_cache/n2001 ), .B(\D_cache/n2002 ), .S0(n2146), .Y(\D_cache/N82 ) );
  MXI4X1 \D_cache/U2343  ( .A(\D_cache/cache[4][101] ), .B(
        \D_cache/cache[5][101] ), .C(\D_cache/cache[6][101] ), .D(
        \D_cache/cache[7][101] ), .S0(n2138), .S1(n2347), .Y(\D_cache/n2000 )
         );
  MXI4X1 \D_cache/U2344  ( .A(\D_cache/cache[0][101] ), .B(
        \D_cache/cache[1][101] ), .C(\D_cache/cache[2][101] ), .D(
        \D_cache/cache[3][101] ), .S0(n2122), .S1(n2349), .Y(\D_cache/n1999 )
         );
  MXI2X1 \D_cache/U2087  ( .A(\D_cache/n1999 ), .B(\D_cache/n2000 ), .S0(n3064), .Y(\D_cache/N83 ) );
  MXI2X1 \D_cache/U2010  ( .A(\D_cache/n1845 ), .B(\D_cache/n1846 ), .S0(n3065), .Y(\D_cache/N160 ) );
  MXI2X1 \D_cache/U1989  ( .A(\D_cache/n1803 ), .B(\D_cache/n1804 ), .S0(n2147), .Y(\D_cache/N181 ) );
  MXI2X1 \D_cache/U2064  ( .A(\D_cache/n1953 ), .B(\D_cache/n1954 ), .S0(
        DCACHE_addr[4]), .Y(\D_cache/N106 ) );
  MXI2X1 \D_cache/U2013  ( .A(\D_cache/n1851 ), .B(\D_cache/n1852 ), .S0(n3067), .Y(\D_cache/N157 ) );
  MXI2X1 \D_cache/U2011  ( .A(\D_cache/n1847 ), .B(\D_cache/n1848 ), .S0(n3067), .Y(\D_cache/N159 ) );
  MXI4X1 \D_cache/U2151  ( .A(\D_cache/cache[4][5] ), .B(\D_cache/cache[5][5] ), .C(\D_cache/cache[6][5] ), .D(\D_cache/cache[7][5] ), .S0(n2132), .S1(n2355), 
        .Y(\D_cache/n1808 ) );
  MXI4X1 \D_cache/U2152  ( .A(\D_cache/cache[0][5] ), .B(\D_cache/cache[1][5] ), .C(\D_cache/cache[2][5] ), .D(\D_cache/cache[3][5] ), .S0(n2093), .S1(n2358), 
        .Y(\D_cache/n1807 ) );
  MXI2X1 \D_cache/U1991  ( .A(\D_cache/n1807 ), .B(\D_cache/n1808 ), .S0(n3064), .Y(\D_cache/N179 ) );
  MXI2X1 \D_cache/U2086  ( .A(\D_cache/n1997 ), .B(\D_cache/n1998 ), .S0(n3066), .Y(\D_cache/N84 ) );
  MXI4X1 \D_cache/U2178  ( .A(\D_cache/cache[0][18] ), .B(
        \D_cache/cache[1][18] ), .C(\D_cache/cache[2][18] ), .D(
        \D_cache/cache[3][18] ), .S0(n2085), .S1(n2253), .Y(\D_cache/n1833 )
         );
  MXI4X1 \D_cache/U2177  ( .A(\D_cache/cache[4][18] ), .B(
        \D_cache/cache[5][18] ), .C(\D_cache/cache[6][18] ), .D(
        \D_cache/cache[7][18] ), .S0(n2084), .S1(n2259), .Y(\D_cache/n1834 )
         );
  MXI2X1 \D_cache/U2004  ( .A(\D_cache/n1833 ), .B(\D_cache/n1834 ), .S0(n3067), .Y(\D_cache/N166 ) );
  MXI2X1 \D_cache/U2012  ( .A(\D_cache/n1849 ), .B(\D_cache/n1850 ), .S0(n3064), .Y(\D_cache/N158 ) );
  MXI4X1 \D_cache/U2169  ( .A(\D_cache/cache[4][14] ), .B(
        \D_cache/cache[5][14] ), .C(\D_cache/cache[6][14] ), .D(
        \D_cache/cache[7][14] ), .S0(n2094), .S1(n2285), .Y(\D_cache/n1826 )
         );
  MXI4X1 \D_cache/U2170  ( .A(\D_cache/cache[0][14] ), .B(
        \D_cache/cache[1][14] ), .C(\D_cache/cache[2][14] ), .D(
        \D_cache/cache[3][14] ), .S0(n2097), .S1(n2301), .Y(\D_cache/n1825 )
         );
  MXI2X1 \D_cache/U2000  ( .A(\D_cache/n1825 ), .B(\D_cache/n1826 ), .S0(
        DCACHE_addr[4]), .Y(\D_cache/N170 ) );
  MXI2X1 \D_cache/U2007  ( .A(\D_cache/n1839 ), .B(\D_cache/n1840 ), .S0(n2146), .Y(\D_cache/N163 ) );
  MXI4X1 \D_cache/U2166  ( .A(\D_cache/cache[0][12] ), .B(
        \D_cache/cache[1][12] ), .C(\D_cache/cache[2][12] ), .D(
        \D_cache/cache[3][12] ), .S0(n2089), .S1(n2324), .Y(\D_cache/n1821 )
         );
  MXI4X1 \D_cache/U2165  ( .A(\D_cache/cache[4][12] ), .B(
        \D_cache/cache[5][12] ), .C(\D_cache/cache[6][12] ), .D(
        \D_cache/cache[7][12] ), .S0(n2088), .S1(n2320), .Y(\D_cache/n1822 )
         );
  MXI2X1 \D_cache/U1998  ( .A(\D_cache/n1821 ), .B(\D_cache/n1822 ), .S0(n3064), .Y(\D_cache/N172 ) );
  MXI2X1 \D_cache/U1999  ( .A(\D_cache/n1823 ), .B(\D_cache/n1824 ), .S0(
        DCACHE_addr[4]), .Y(\D_cache/N171 ) );
  MXI2X1 \D_cache/U1997  ( .A(\D_cache/n1819 ), .B(\D_cache/n1820 ), .S0(n2146), .Y(\D_cache/N173 ) );
  MXI2X1 \D_cache/U2052  ( .A(\D_cache/n1929 ), .B(\D_cache/n1930 ), .S0(n3064), .Y(\D_cache/N118 ) );
  MXI2X1 \D_cache/U2057  ( .A(\D_cache/n1939 ), .B(\D_cache/n1940 ), .S0(n3064), .Y(\D_cache/N113 ) );
  MXI2X1 \D_cache/U2050  ( .A(\D_cache/n1925 ), .B(\D_cache/n1926 ), .S0(n3065), .Y(\D_cache/N120 ) );
  MXI2X1 \D_cache/U2053  ( .A(\D_cache/n1931 ), .B(\D_cache/n1932 ), .S0(n2147), .Y(\D_cache/N117 ) );
  MXI2X1 \D_cache/U2051  ( .A(\D_cache/n1927 ), .B(\D_cache/n1928 ), .S0(n3067), .Y(\D_cache/N119 ) );
  MXI2X1 \D_cache/U2056  ( .A(\D_cache/n1937 ), .B(\D_cache/n1938 ), .S0(n3064), .Y(\D_cache/N114 ) );
  MXI2X1 \D_cache/U2055  ( .A(\D_cache/n1935 ), .B(\D_cache/n1936 ), .S0(n3062), .Y(\D_cache/N115 ) );
  MXI2X1 \D_cache/U2060  ( .A(\D_cache/n1945 ), .B(\D_cache/n1946 ), .S0(
        DCACHE_addr[4]), .Y(\D_cache/N110 ) );
  MXI2X1 \D_cache/U2054  ( .A(\D_cache/n1933 ), .B(\D_cache/n1934 ), .S0(n2147), .Y(\D_cache/N116 ) );
  MXI2X1 \D_cache/U2059  ( .A(\D_cache/n1943 ), .B(\D_cache/n1944 ), .S0(n4041), .Y(\D_cache/N111 ) );
  MXI2X1 \D_cache/U2058  ( .A(\D_cache/n1941 ), .B(\D_cache/n1942 ), .S0(n3067), .Y(\D_cache/N112 ) );
  MXI4X1 \D_cache/U2142  ( .A(\D_cache/cache[0][0] ), .B(\D_cache/cache[1][0] ), .C(\D_cache/cache[2][0] ), .D(\D_cache/cache[3][0] ), .S0(n2116), .S1(n2385), 
        .Y(\D_cache/n1797 ) );
  MXI4X1 \D_cache/U2141  ( .A(\D_cache/cache[4][0] ), .B(\D_cache/cache[5][0] ), .C(\D_cache/cache[6][0] ), .D(\D_cache/cache[7][0] ), .S0(n2113), .S1(n2382), 
        .Y(\D_cache/n1798 ) );
  MXI2X1 \D_cache/U1986  ( .A(\D_cache/n1797 ), .B(\D_cache/n1798 ), .S0(
        n10321), .Y(\D_cache/N184 ) );
  MXI4X1 \D_cache/U2145  ( .A(\D_cache/cache[4][2] ), .B(\D_cache/cache[5][2] ), .C(\D_cache/cache[6][2] ), .D(\D_cache/cache[7][2] ), .S0(n2087), .S1(n2247), 
        .Y(\D_cache/n1802 ) );
  MXI4X1 \D_cache/U2146  ( .A(\D_cache/cache[0][2] ), .B(\D_cache/cache[1][2] ), .C(\D_cache/cache[2][2] ), .D(\D_cache/cache[3][2] ), .S0(n2090), .S1(n2242), 
        .Y(\D_cache/n1801 ) );
  MXI2X1 \D_cache/U1988  ( .A(\D_cache/n1801 ), .B(\D_cache/n1802 ), .S0(n3065), .Y(\D_cache/N182 ) );
  MXI4X1 \D_cache/U2143  ( .A(\D_cache/cache[4][1] ), .B(\D_cache/cache[5][1] ), .C(\D_cache/cache[6][1] ), .D(\D_cache/cache[7][1] ), .S0(n2123), .S1(n2279), 
        .Y(\D_cache/n1800 ) );
  MXI4X1 \D_cache/U2144  ( .A(\D_cache/cache[0][1] ), .B(\D_cache/cache[1][1] ), .C(\D_cache/cache[2][1] ), .D(\D_cache/cache[3][1] ), .S0(n2118), .S1(n2295), 
        .Y(\D_cache/n1799 ) );
  MXI2X1 \D_cache/U1987  ( .A(\D_cache/n1799 ), .B(\D_cache/n1800 ), .S0(n3063), .Y(\D_cache/N183 ) );
  MXI4X1 \D_cache/U2149  ( .A(\D_cache/cache[4][4] ), .B(\D_cache/cache[5][4] ), .C(\D_cache/cache[6][4] ), .D(\D_cache/cache[7][4] ), .S0(n2098), .S1(n2257), 
        .Y(\D_cache/n1806 ) );
  MXI4X1 \D_cache/U2150  ( .A(\D_cache/cache[0][4] ), .B(\D_cache/cache[1][4] ), .C(\D_cache/cache[2][4] ), .D(\D_cache/cache[3][4] ), .S0(n2089), .S1(n2251), 
        .Y(\D_cache/n1805 ) );
  MXI2X1 \D_cache/U1990  ( .A(\D_cache/n1805 ), .B(\D_cache/n1806 ), .S0(n3065), .Y(\D_cache/N180 ) );
  MXI2X1 \D_cache/U2072  ( .A(\D_cache/n1969 ), .B(\D_cache/n1970 ), .S0(
        DCACHE_addr[4]), .Y(\D_cache/N98 ) );
  MXI4X1 \D_cache/U2428  ( .A(\D_cache/cache[0][143] ), .B(
        \D_cache/cache[1][143] ), .C(\D_cache/cache[2][143] ), .D(
        \D_cache/cache[3][143] ), .S0(n2126), .S1(n2415), .Y(\D_cache/n2083 )
         );
  MXI4X1 \D_cache/U2426  ( .A(\D_cache/cache[0][142] ), .B(
        \D_cache/cache[1][142] ), .C(\D_cache/cache[2][142] ), .D(
        \D_cache/cache[3][142] ), .S0(n2068), .S1(n2408), .Y(\D_cache/n2081 )
         );
  MXI4X1 \D_cache/U2425  ( .A(\D_cache/cache[4][142] ), .B(
        \D_cache/cache[5][142] ), .C(\D_cache/cache[6][142] ), .D(
        \D_cache/cache[7][142] ), .S0(n2061), .S1(n2405), .Y(\D_cache/n2082 )
         );
  MXI4X1 \D_cache/U2424  ( .A(\D_cache/cache[0][141] ), .B(
        \D_cache/cache[1][141] ), .C(\D_cache/cache[2][141] ), .D(
        \D_cache/cache[3][141] ), .S0(n2137), .S1(n2411), .Y(\D_cache/n2079 )
         );
  MXI4X1 \D_cache/U2404  ( .A(\D_cache/cache[0][131] ), .B(
        \D_cache/cache[1][131] ), .C(\D_cache/cache[2][131] ), .D(
        \D_cache/cache[3][131] ), .S0(n2128), .S1(n2440), .Y(\D_cache/n2059 )
         );
  MXI4X1 \D_cache/U2403  ( .A(\D_cache/cache[4][131] ), .B(
        \D_cache/cache[5][131] ), .C(\D_cache/cache[6][131] ), .D(
        \D_cache/cache[7][131] ), .S0(n2128), .S1(n2439), .Y(\D_cache/n2060 )
         );
  MXI4X1 \D_cache/U2399  ( .A(\D_cache/cache[4][129] ), .B(
        \D_cache/cache[5][129] ), .C(\D_cache/cache[6][129] ), .D(
        \D_cache/cache[7][129] ), .S0(n2130), .S1(n2170), .Y(\D_cache/n2056 )
         );
  MXI4X1 \D_cache/U2400  ( .A(\D_cache/cache[0][129] ), .B(
        \D_cache/cache[1][129] ), .C(\D_cache/cache[2][129] ), .D(
        \D_cache/cache[3][129] ), .S0(n2126), .S1(n2171), .Y(\D_cache/n2055 )
         );
  MXI4X1 \D_cache/U2410  ( .A(\D_cache/cache[0][134] ), .B(
        \D_cache/cache[1][134] ), .C(\D_cache/cache[2][134] ), .D(
        \D_cache/cache[3][134] ), .S0(n2069), .S1(n2421), .Y(\D_cache/n2065 )
         );
  MXI4X1 \D_cache/U2409  ( .A(\D_cache/cache[4][134] ), .B(
        \D_cache/cache[5][134] ), .C(\D_cache/cache[6][134] ), .D(
        \D_cache/cache[7][134] ), .S0(n2107), .S1(n2418), .Y(\D_cache/n2066 )
         );
  MXI4X1 \D_cache/U2417  ( .A(\D_cache/cache[4][138] ), .B(
        \D_cache/cache[5][138] ), .C(\D_cache/cache[6][138] ), .D(
        \D_cache/cache[7][138] ), .S0(n2093), .S1(n2417), .Y(\D_cache/n2074 )
         );
  MXI4X1 \D_cache/U2418  ( .A(\D_cache/cache[0][138] ), .B(
        \D_cache/cache[1][138] ), .C(\D_cache/cache[2][138] ), .D(
        \D_cache/cache[3][138] ), .S0(n2096), .S1(n2420), .Y(\D_cache/n2073 )
         );
  MXI4X1 \D_cache/U2405  ( .A(\D_cache/cache[4][132] ), .B(
        \D_cache/cache[5][132] ), .C(\D_cache/cache[6][132] ), .D(
        \D_cache/cache[7][132] ), .S0(n2142), .S1(n2419), .Y(\D_cache/n2062 )
         );
  MXI4X1 \D_cache/U2406  ( .A(\D_cache/cache[0][132] ), .B(
        \D_cache/cache[1][132] ), .C(\D_cache/cache[2][132] ), .D(
        \D_cache/cache[3][132] ), .S0(n2141), .S1(n2423), .Y(\D_cache/n2061 )
         );
  MXI4X1 \D_cache/U2431  ( .A(\D_cache/cache[4][145] ), .B(
        \D_cache/cache[5][145] ), .C(\D_cache/cache[6][145] ), .D(
        \D_cache/cache[7][145] ), .S0(n2128), .S1(n2430), .Y(\D_cache/n2088 )
         );
  MXI4X1 \D_cache/U2441  ( .A(\D_cache/cache[4][150] ), .B(
        \D_cache/cache[5][150] ), .C(\D_cache/cache[6][150] ), .D(
        \D_cache/cache[7][150] ), .S0(n2129), .S1(n2427), .Y(\D_cache/n2098 )
         );
  MXI4X1 \D_cache/U2442  ( .A(\D_cache/cache[0][150] ), .B(
        \D_cache/cache[1][150] ), .C(\D_cache/cache[2][150] ), .D(
        \D_cache/cache[3][150] ), .S0(n2109), .S1(n2432), .Y(\D_cache/n2097 )
         );
  MXI4X1 \D_cache/U2433  ( .A(\D_cache/cache[4][146] ), .B(
        \D_cache/cache[5][146] ), .C(\D_cache/cache[6][146] ), .D(
        \D_cache/cache[7][146] ), .S0(n2074), .S1(n2426), .Y(\D_cache/n2090 )
         );
  MXI4X1 \D_cache/U2434  ( .A(\D_cache/cache[0][146] ), .B(
        \D_cache/cache[1][146] ), .C(\D_cache/cache[2][146] ), .D(
        \D_cache/cache[3][146] ), .S0(n2100), .S1(n2431), .Y(\D_cache/n2089 )
         );
  MXI4X1 \D_cache/U2435  ( .A(\D_cache/cache[4][147] ), .B(
        \D_cache/cache[5][147] ), .C(\D_cache/cache[6][147] ), .D(
        \D_cache/cache[7][147] ), .S0(n2129), .S1(n2179), .Y(\D_cache/n2092 )
         );
  MXI4X1 \D_cache/U2436  ( .A(\D_cache/cache[0][147] ), .B(
        \D_cache/cache[1][147] ), .C(\D_cache/cache[2][147] ), .D(
        \D_cache/cache[3][147] ), .S0(n2127), .S1(n2402), .Y(\D_cache/n2091 )
         );
  MXI2X1 \D_cache/U2133  ( .A(\D_cache/n2091 ), .B(\D_cache/n2092 ), .S0(n3067), .Y(\D_cache/N37 ) );
  MXI4X1 \D_cache/U2437  ( .A(\D_cache/cache[4][148] ), .B(
        \D_cache/cache[5][148] ), .C(\D_cache/cache[6][148] ), .D(
        \D_cache/cache[7][148] ), .S0(n2127), .S1(n2174), .Y(\D_cache/n2094 )
         );
  MXI4X1 \D_cache/U2438  ( .A(\D_cache/cache[0][148] ), .B(
        \D_cache/cache[1][148] ), .C(\D_cache/cache[2][148] ), .D(
        \D_cache/cache[3][148] ), .S0(n2099), .S1(n2177), .Y(\D_cache/n2093 )
         );
  MXI4X1 \D_cache/U2430  ( .A(\D_cache/cache[0][144] ), .B(
        \D_cache/cache[1][144] ), .C(\D_cache/cache[2][144] ), .D(
        \D_cache/cache[3][144] ), .S0(n2072), .S1(n2412), .Y(\D_cache/n2085 )
         );
  MXI4X1 \D_cache/U2420  ( .A(\D_cache/cache[0][139] ), .B(
        \D_cache/cache[1][139] ), .C(\D_cache/cache[2][139] ), .D(
        \D_cache/cache[3][139] ), .S0(n2073), .S1(n2416), .Y(\D_cache/n2075 )
         );
  MXI4X1 \D_cache/U2419  ( .A(\D_cache/cache[4][139] ), .B(
        \D_cache/cache[5][139] ), .C(\D_cache/cache[6][139] ), .D(
        \D_cache/cache[7][139] ), .S0(n2143), .S1(n2414), .Y(\D_cache/n2076 )
         );
  MXI2X1 \D_cache/U2137  ( .A(\D_cache/n2099 ), .B(\D_cache/n2100 ), .S0(n3063), .Y(\D_cache/N33 ) );
  MXI4X1 \D_cache/U2450  ( .A(\D_cache/cache[0][154] ), .B(
        \D_cache/cache[1][154] ), .C(\D_cache/cache[2][154] ), .D(
        \D_cache/cache[3][154] ), .S0(n2111), .S1(n2181), .Y(\D_cache/n2105 )
         );
  MXI4X1 \D_cache/U2449  ( .A(\D_cache/cache[4][154] ), .B(
        \D_cache/cache[5][154] ), .C(\D_cache/cache[6][154] ), .D(
        \D_cache/cache[7][154] ), .S0(n2109), .S1(n2180), .Y(\D_cache/n2106 )
         );
  MXI2X1 \D_cache/U2140  ( .A(\D_cache/n2105 ), .B(\D_cache/n2106 ), .S0(n3065), .Y(\D_cache/N30 ) );
  DFFRX4 \i_MIPS/ID_EX_reg[79]  ( .D(\i_MIPS/n506 ), .CK(clk), .RN(n4058), .Q(
        \i_MIPS/ID_EX[79] ), .QN(n54) );
  MXI4XL \D_cache/U2330  ( .A(\D_cache/cache[0][94] ), .B(
        \D_cache/cache[1][94] ), .C(\D_cache/cache[2][94] ), .D(
        \D_cache/cache[3][94] ), .S0(n2119), .S1(n2187), .Y(\D_cache/n1985 )
         );
  MXI4XL \D_cache/U2329  ( .A(\D_cache/cache[4][94] ), .B(
        \D_cache/cache[5][94] ), .C(\D_cache/cache[6][94] ), .D(
        \D_cache/cache[7][94] ), .S0(n2077), .S1(n2184), .Y(\D_cache/n1986 )
         );
  MXI2XL \D_cache/U2080  ( .A(\D_cache/n1985 ), .B(\D_cache/n1986 ), .S0(n3063), .Y(\D_cache/N90 ) );
  MXI4XL \D_cache/U2324  ( .A(\D_cache/cache[0][91] ), .B(
        \D_cache/cache[1][91] ), .C(\D_cache/cache[2][91] ), .D(
        \D_cache/cache[3][91] ), .S0(n2090), .S1(n2332), .Y(\D_cache/n1979 )
         );
  MXI4XL \D_cache/U2323  ( .A(\D_cache/cache[4][91] ), .B(
        \D_cache/cache[5][91] ), .C(\D_cache/cache[6][91] ), .D(
        \D_cache/cache[7][91] ), .S0(n2074), .S1(n2184), .Y(\D_cache/n1980 )
         );
  MXI2XL \D_cache/U2077  ( .A(\D_cache/n1979 ), .B(\D_cache/n1980 ), .S0(n2146), .Y(\D_cache/N93 ) );
  MXI4XL \D_cache/U2312  ( .A(\D_cache/cache[0][85] ), .B(
        \D_cache/cache[1][85] ), .C(\D_cache/cache[2][85] ), .D(
        \D_cache/cache[3][85] ), .S0(n2064), .S1(n2305), .Y(\D_cache/n1967 )
         );
  MXI4XL \D_cache/U2311  ( .A(\D_cache/cache[4][85] ), .B(
        \D_cache/cache[5][85] ), .C(\D_cache/cache[6][85] ), .D(
        \D_cache/cache[7][85] ), .S0(n2104), .S1(n2298), .Y(\D_cache/n1968 )
         );
  MXI2XL \D_cache/U2071  ( .A(\D_cache/n1967 ), .B(\D_cache/n1968 ), .S0(n3063), .Y(\D_cache/N99 ) );
  MXI4XL \D_cache/U2318  ( .A(\D_cache/cache[0][88] ), .B(
        \D_cache/cache[1][88] ), .C(\D_cache/cache[2][88] ), .D(
        \D_cache/cache[3][88] ), .S0(n2108), .S1(n2183), .Y(\D_cache/n1973 )
         );
  MXI4XL \D_cache/U2317  ( .A(\D_cache/cache[4][88] ), .B(
        \D_cache/cache[5][88] ), .C(\D_cache/cache[6][88] ), .D(
        \D_cache/cache[7][88] ), .S0(n2140), .S1(n2178), .Y(\D_cache/n1974 )
         );
  MXI2XL \D_cache/U2074  ( .A(\D_cache/n1973 ), .B(\D_cache/n1974 ), .S0(n3065), .Y(\D_cache/N96 ) );
  MXI4XL \D_cache/U2354  ( .A(\D_cache/cache[0][106] ), .B(
        \D_cache/cache[1][106] ), .C(\D_cache/cache[2][106] ), .D(
        \D_cache/cache[3][106] ), .S0(n2066), .S1(n2184), .Y(\D_cache/n2009 )
         );
  MXI4XL \D_cache/U2353  ( .A(\D_cache/cache[4][106] ), .B(
        \D_cache/cache[5][106] ), .C(\D_cache/cache[6][106] ), .D(
        \D_cache/cache[7][106] ), .S0(n2061), .S1(n2392), .Y(\D_cache/n2010 )
         );
  MXI2XL \D_cache/U2092  ( .A(\D_cache/n2009 ), .B(\D_cache/n2010 ), .S0(n3067), .Y(\D_cache/N78 ) );
  MXI4XL \D_cache/U2336  ( .A(\D_cache/cache[0][97] ), .B(
        \D_cache/cache[1][97] ), .C(\D_cache/cache[2][97] ), .D(
        \D_cache/cache[3][97] ), .S0(n2121), .S1(n2306), .Y(\D_cache/n1991 )
         );
  MXI4XL \D_cache/U2335  ( .A(\D_cache/cache[4][97] ), .B(
        \D_cache/cache[5][97] ), .C(\D_cache/cache[6][97] ), .D(
        \D_cache/cache[7][97] ), .S0(n2116), .S1(n2290), .Y(\D_cache/n1992 )
         );
  MXI4XL \D_cache/U2342  ( .A(\D_cache/cache[0][100] ), .B(
        \D_cache/cache[1][100] ), .C(\D_cache/cache[2][100] ), .D(
        \D_cache/cache[3][100] ), .S0(n2082), .S1(n2181), .Y(\D_cache/n1997 )
         );
  MXI4XL \D_cache/U2341  ( .A(\D_cache/cache[4][100] ), .B(
        \D_cache/cache[5][100] ), .C(\D_cache/cache[6][100] ), .D(
        \D_cache/cache[7][100] ), .S0(n2097), .S1(n2176), .Y(\D_cache/n1998 )
         );
  MXI4XL \D_cache/U2300  ( .A(\D_cache/cache[0][79] ), .B(
        \D_cache/cache[1][79] ), .C(\D_cache/cache[2][79] ), .D(
        \D_cache/cache[3][79] ), .S0(n2085), .S1(n2304), .Y(\D_cache/n1955 )
         );
  MXI4XL \D_cache/U2299  ( .A(\D_cache/cache[4][79] ), .B(
        \D_cache/cache[5][79] ), .C(\D_cache/cache[6][79] ), .D(
        \D_cache/cache[7][79] ), .S0(n2144), .S1(n2282), .Y(\D_cache/n1956 )
         );
  MXI4XL \D_cache/U2306  ( .A(\D_cache/cache[0][82] ), .B(
        \D_cache/cache[1][82] ), .C(\D_cache/cache[2][82] ), .D(
        \D_cache/cache[3][82] ), .S0(n2124), .S1(n2431), .Y(\D_cache/n1961 )
         );
  MXI4XL \D_cache/U2305  ( .A(\D_cache/cache[4][82] ), .B(
        \D_cache/cache[5][82] ), .C(\D_cache/cache[6][82] ), .D(
        \D_cache/cache[7][82] ), .S0(n2101), .S1(n2420), .Y(\D_cache/n1962 )
         );
  MXI4XL \D_cache/U2294  ( .A(\D_cache/cache[0][76] ), .B(
        \D_cache/cache[1][76] ), .C(\D_cache/cache[2][76] ), .D(
        \D_cache/cache[3][76] ), .S0(n2088), .S1(n2300), .Y(\D_cache/n1949 )
         );
  MXI4XL \D_cache/U2293  ( .A(\D_cache/cache[4][76] ), .B(
        \D_cache/cache[5][76] ), .C(\D_cache/cache[6][76] ), .D(
        \D_cache/cache[7][76] ), .S0(n2112), .S1(n2273), .Y(\D_cache/n1950 )
         );
  MXI4XL \D_cache/U2313  ( .A(\D_cache/cache[4][86] ), .B(
        \D_cache/cache[5][86] ), .C(\D_cache/cache[6][86] ), .D(
        \D_cache/cache[7][86] ), .S0(n2139), .S1(n2407), .Y(\D_cache/n1970 )
         );
  MXI4XL \D_cache/U2314  ( .A(\D_cache/cache[0][86] ), .B(
        \D_cache/cache[1][86] ), .C(\D_cache/cache[2][86] ), .D(
        \D_cache/cache[3][86] ), .S0(n2116), .S1(n2408), .Y(\D_cache/n1969 )
         );
  MXI4XL \D_cache/U2331  ( .A(\D_cache/cache[4][95] ), .B(
        \D_cache/cache[5][95] ), .C(\D_cache/cache[6][95] ), .D(
        \D_cache/cache[7][95] ), .S0(n2141), .S1(n2404), .Y(\D_cache/n1988 )
         );
  MXI4XL \D_cache/U2332  ( .A(\D_cache/cache[0][95] ), .B(
        \D_cache/cache[1][95] ), .C(\D_cache/cache[2][95] ), .D(
        \D_cache/cache[3][95] ), .S0(n2062), .S1(n2403), .Y(\D_cache/n1987 )
         );
  MXI2XL \D_cache/U2081  ( .A(\D_cache/n1987 ), .B(\D_cache/n1988 ), .S0(
        DCACHE_addr[4]), .Y(\D_cache/N89 ) );
  MXI4XL \D_cache/U2327  ( .A(\D_cache/cache[4][93] ), .B(
        \D_cache/cache[5][93] ), .C(\D_cache/cache[6][93] ), .D(
        \D_cache/cache[7][93] ), .S0(n2071), .S1(n2189), .Y(\D_cache/n1984 )
         );
  MXI4XL \D_cache/U2328  ( .A(\D_cache/cache[0][93] ), .B(
        \D_cache/cache[1][93] ), .C(\D_cache/cache[2][93] ), .D(
        \D_cache/cache[3][93] ), .S0(n2072), .S1(n2195), .Y(\D_cache/n1983 )
         );
  MXI2XL \D_cache/U2079  ( .A(\D_cache/n1983 ), .B(\D_cache/n1984 ), .S0(n2146), .Y(\D_cache/N91 ) );
  MXI4XL \D_cache/U2325  ( .A(\D_cache/cache[4][92] ), .B(
        \D_cache/cache[5][92] ), .C(\D_cache/cache[6][92] ), .D(
        \D_cache/cache[7][92] ), .S0(n2138), .S1(n2170), .Y(\D_cache/n1982 )
         );
  MXI4XL \D_cache/U2326  ( .A(\D_cache/cache[0][92] ), .B(
        \D_cache/cache[1][92] ), .C(\D_cache/cache[2][92] ), .D(
        \D_cache/cache[3][92] ), .S0(n2137), .S1(n2433), .Y(\D_cache/n1981 )
         );
  MXI2XL \D_cache/U2078  ( .A(\D_cache/n1981 ), .B(\D_cache/n1982 ), .S0(n4041), .Y(\D_cache/N92 ) );
  MXI4XL \D_cache/U2321  ( .A(\D_cache/cache[4][90] ), .B(
        \D_cache/cache[5][90] ), .C(\D_cache/cache[6][90] ), .D(
        \D_cache/cache[7][90] ), .S0(n2124), .S1(n2337), .Y(\D_cache/n1978 )
         );
  MXI4XL \D_cache/U2322  ( .A(\D_cache/cache[0][90] ), .B(
        \D_cache/cache[1][90] ), .C(\D_cache/cache[2][90] ), .D(
        \D_cache/cache[3][90] ), .S0(n2139), .S1(n2369), .Y(\D_cache/n1977 )
         );
  MXI2XL \D_cache/U2076  ( .A(\D_cache/n1977 ), .B(\D_cache/n1978 ), .S0(n3062), .Y(\D_cache/N94 ) );
  MXI4XL \D_cache/U2307  ( .A(\D_cache/cache[4][83] ), .B(
        \D_cache/cache[5][83] ), .C(\D_cache/cache[6][83] ), .D(
        \D_cache/cache[7][83] ), .S0(n2109), .S1(n2223), .Y(\D_cache/n1964 )
         );
  MXI4XL \D_cache/U2308  ( .A(\D_cache/cache[0][83] ), .B(
        \D_cache/cache[1][83] ), .C(\D_cache/cache[2][83] ), .D(
        \D_cache/cache[3][83] ), .S0(n2071), .S1(n2218), .Y(\D_cache/n1963 )
         );
  MXI2XL \D_cache/U2069  ( .A(\D_cache/n1963 ), .B(\D_cache/n1964 ), .S0(n3064), .Y(\D_cache/N101 ) );
  MXI4XL \D_cache/U2319  ( .A(\D_cache/cache[4][89] ), .B(
        \D_cache/cache[5][89] ), .C(\D_cache/cache[6][89] ), .D(
        \D_cache/cache[7][89] ), .S0(n2101), .S1(n2336), .Y(\D_cache/n1976 )
         );
  MXI4XL \D_cache/U2320  ( .A(\D_cache/cache[0][89] ), .B(
        \D_cache/cache[1][89] ), .C(\D_cache/cache[2][89] ), .D(
        \D_cache/cache[3][89] ), .S0(n2137), .S1(n2183), .Y(\D_cache/n1975 )
         );
  MXI2XL \D_cache/U2075  ( .A(\D_cache/n1975 ), .B(\D_cache/n1976 ), .S0(n2146), .Y(\D_cache/N95 ) );
  MXI4XL \D_cache/U2339  ( .A(\D_cache/cache[4][99] ), .B(
        \D_cache/cache[5][99] ), .C(\D_cache/cache[6][99] ), .D(
        \D_cache/cache[7][99] ), .S0(n2076), .S1(n2183), .Y(\D_cache/n1996 )
         );
  MXI4XL \D_cache/U2340  ( .A(\D_cache/cache[0][99] ), .B(
        \D_cache/cache[1][99] ), .C(\D_cache/cache[2][99] ), .D(
        \D_cache/cache[3][99] ), .S0(n2113), .S1(n2184), .Y(\D_cache/n1995 )
         );
  MXI2XL \D_cache/U2085  ( .A(\D_cache/n1995 ), .B(\D_cache/n1996 ), .S0(n2146), .Y(\D_cache/N85 ) );
  MXI4XL \D_cache/U2337  ( .A(\D_cache/cache[4][98] ), .B(
        \D_cache/cache[5][98] ), .C(\D_cache/cache[6][98] ), .D(
        \D_cache/cache[7][98] ), .S0(n2082), .S1(n2186), .Y(\D_cache/n1994 )
         );
  MXI4XL \D_cache/U2338  ( .A(\D_cache/cache[0][98] ), .B(
        \D_cache/cache[1][98] ), .C(\D_cache/cache[2][98] ), .D(
        \D_cache/cache[3][98] ), .S0(n2115), .S1(n2185), .Y(\D_cache/n1993 )
         );
  MXI2XL \D_cache/U2084  ( .A(\D_cache/n1993 ), .B(\D_cache/n1994 ), .S0(
        n10321), .Y(\D_cache/N86 ) );
  MXI4XL \D_cache/U2303  ( .A(\D_cache/cache[4][81] ), .B(
        \D_cache/cache[5][81] ), .C(\D_cache/cache[6][81] ), .D(
        \D_cache/cache[7][81] ), .S0(n2102), .S1(n2430), .Y(\D_cache/n1960 )
         );
  MXI4XL \D_cache/U2304  ( .A(\D_cache/cache[0][81] ), .B(
        \D_cache/cache[1][81] ), .C(\D_cache/cache[2][81] ), .D(
        \D_cache/cache[3][81] ), .S0(n2139), .S1(n2440), .Y(\D_cache/n1959 )
         );
  MXI4XL \D_cache/U2309  ( .A(\D_cache/cache[4][84] ), .B(
        \D_cache/cache[5][84] ), .C(\D_cache/cache[6][84] ), .D(
        \D_cache/cache[7][84] ), .S0(n2143), .S1(n2435), .Y(\D_cache/n1966 )
         );
  MXI4XL \D_cache/U2310  ( .A(\D_cache/cache[0][84] ), .B(
        \D_cache/cache[1][84] ), .C(\D_cache/cache[2][84] ), .D(
        \D_cache/cache[3][84] ), .S0(n2063), .S1(n2437), .Y(\D_cache/n1965 )
         );
  MXI2XL \D_cache/U2070  ( .A(\D_cache/n1965 ), .B(\D_cache/n1966 ), .S0(n3064), .Y(\D_cache/N100 ) );
  MXI4XL \D_cache/U2297  ( .A(\D_cache/cache[4][78] ), .B(
        \D_cache/cache[5][78] ), .C(\D_cache/cache[6][78] ), .D(
        \D_cache/cache[7][78] ), .S0(n2125), .S1(n2248), .Y(\D_cache/n1954 )
         );
  MXI4XL \D_cache/U2298  ( .A(\D_cache/cache[0][78] ), .B(
        \D_cache/cache[1][78] ), .C(\D_cache/cache[2][78] ), .D(
        \D_cache/cache[3][78] ), .S0(n2067), .S1(n2254), .Y(\D_cache/n1953 )
         );
  MXI4XL \D_cache/U2349  ( .A(\D_cache/cache[4][104] ), .B(
        \D_cache/cache[5][104] ), .C(\D_cache/cache[6][104] ), .D(
        \D_cache/cache[7][104] ), .S0(n2064), .S1(n2391), .Y(\D_cache/n2006 )
         );
  MXI4XL \D_cache/U2350  ( .A(\D_cache/cache[0][104] ), .B(
        \D_cache/cache[1][104] ), .C(\D_cache/cache[2][104] ), .D(
        \D_cache/cache[3][104] ), .S0(n2062), .S1(n2390), .Y(\D_cache/n2005 )
         );
  MXI2XL \D_cache/U2090  ( .A(\D_cache/n2005 ), .B(\D_cache/n2006 ), .S0(
        n10321), .Y(\D_cache/N80 ) );
  MXI4XL \D_cache/U2355  ( .A(\D_cache/cache[4][107] ), .B(
        \D_cache/cache[5][107] ), .C(\D_cache/cache[6][107] ), .D(
        \D_cache/cache[7][107] ), .S0(n2080), .S1(n2213), .Y(\D_cache/n2012 )
         );
  MXI4XL \D_cache/U2356  ( .A(\D_cache/cache[0][107] ), .B(
        \D_cache/cache[1][107] ), .C(\D_cache/cache[2][107] ), .D(
        \D_cache/cache[3][107] ), .S0(DCACHE_addr[2]), .S1(n2210), .Y(
        \D_cache/n2011 ) );
  MXI2XL \D_cache/U2093  ( .A(\D_cache/n2011 ), .B(\D_cache/n2012 ), .S0(n3063), .Y(\D_cache/N77 ) );
  MXI4XL \D_cache/U2357  ( .A(\D_cache/cache[4][108] ), .B(
        \D_cache/cache[5][108] ), .C(\D_cache/cache[6][108] ), .D(
        \D_cache/cache[7][108] ), .S0(n2067), .S1(n2198), .Y(\D_cache/n2014 )
         );
  MXI4XL \D_cache/U2358  ( .A(\D_cache/cache[0][108] ), .B(
        \D_cache/cache[1][108] ), .C(\D_cache/cache[2][108] ), .D(
        \D_cache/cache[3][108] ), .S0(n2068), .S1(n2197), .Y(\D_cache/n2013 )
         );
  MXI2XL \D_cache/U2094  ( .A(\D_cache/n2013 ), .B(\D_cache/n2014 ), .S0(n3062), .Y(\D_cache/N76 ) );
  MXI4XL \D_cache/U2295  ( .A(\D_cache/cache[4][77] ), .B(
        \D_cache/cache[5][77] ), .C(\D_cache/cache[6][77] ), .D(
        \D_cache/cache[7][77] ), .S0(n2083), .S1(n2205), .Y(\D_cache/n1952 )
         );
  MXI4XL \D_cache/U2296  ( .A(\D_cache/cache[0][77] ), .B(
        \D_cache/cache[1][77] ), .C(\D_cache/cache[2][77] ), .D(
        \D_cache/cache[3][77] ), .S0(n2077), .S1(n2204), .Y(\D_cache/n1951 )
         );
  MXI2XL \D_cache/U2063  ( .A(\D_cache/n1951 ), .B(\D_cache/n1952 ), .S0(
        n10321), .Y(\D_cache/N107 ) );
  MXI4XL \D_cache/U2372  ( .A(\D_cache/cache[0][115] ), .B(
        \D_cache/cache[1][115] ), .C(\D_cache/cache[2][115] ), .D(
        \D_cache/cache[3][115] ), .S0(n2086), .S1(n2200), .Y(\D_cache/n2027 )
         );
  MXI4XL \D_cache/U2371  ( .A(\D_cache/cache[4][115] ), .B(
        \D_cache/cache[5][115] ), .C(\D_cache/cache[6][115] ), .D(
        \D_cache/cache[7][115] ), .S0(n2073), .S1(n2199), .Y(\D_cache/n2028 )
         );
  MXI2XL \D_cache/U2101  ( .A(\D_cache/n2027 ), .B(\D_cache/n2028 ), .S0(n3063), .Y(\D_cache/N69 ) );
  MXI4XL \D_cache/U2275  ( .A(\D_cache/cache[4][67] ), .B(
        \D_cache/cache[5][67] ), .C(\D_cache/cache[6][67] ), .D(
        \D_cache/cache[7][67] ), .S0(n2095), .S1(n2271), .Y(\D_cache/n1932 )
         );
  MXI4XL \D_cache/U2276  ( .A(\D_cache/cache[0][67] ), .B(
        \D_cache/cache[1][67] ), .C(\D_cache/cache[2][67] ), .D(
        \D_cache/cache[3][67] ), .S0(n2064), .S1(n2281), .Y(\D_cache/n1931 )
         );
  MXI4XL \D_cache/U2273  ( .A(\D_cache/cache[4][66] ), .B(
        \D_cache/cache[5][66] ), .C(\D_cache/cache[6][66] ), .D(
        \D_cache/cache[7][66] ), .S0(n2077), .S1(n2299), .Y(\D_cache/n1930 )
         );
  MXI4XL \D_cache/U2274  ( .A(\D_cache/cache[0][66] ), .B(
        \D_cache/cache[1][66] ), .C(\D_cache/cache[2][66] ), .D(
        \D_cache/cache[3][66] ), .S0(n2115), .S1(n2303), .Y(\D_cache/n1929 )
         );
  MXI4XL \D_cache/U2392  ( .A(\D_cache/cache[0][125] ), .B(
        \D_cache/cache[1][125] ), .C(\D_cache/cache[2][125] ), .D(
        \D_cache/cache[3][125] ), .S0(n2075), .S1(n2427), .Y(\D_cache/n2047 )
         );
  MXI4XL \D_cache/U2391  ( .A(\D_cache/cache[4][125] ), .B(
        \D_cache/cache[5][125] ), .C(\D_cache/cache[6][125] ), .D(
        \D_cache/cache[7][125] ), .S0(n2089), .S1(n2424), .Y(\D_cache/n2048 )
         );
  MXI2XL \D_cache/U2111  ( .A(\D_cache/n2047 ), .B(\D_cache/n2048 ), .S0(
        DCACHE_addr[4]), .Y(\D_cache/N59 ) );
  MXI4XL \D_cache/U2386  ( .A(\D_cache/cache[0][122] ), .B(
        \D_cache/cache[1][122] ), .C(\D_cache/cache[2][122] ), .D(
        \D_cache/cache[3][122] ), .S0(n2064), .S1(n2277), .Y(\D_cache/n2041 )
         );
  MXI4XL \D_cache/U2385  ( .A(\D_cache/cache[4][122] ), .B(
        \D_cache/cache[5][122] ), .C(\D_cache/cache[6][122] ), .D(
        \D_cache/cache[7][122] ), .S0(n2083), .S1(n2275), .Y(\D_cache/n2042 )
         );
  MXI2XL \D_cache/U2108  ( .A(\D_cache/n2041 ), .B(\D_cache/n2042 ), .S0(n4041), .Y(\D_cache/N62 ) );
  MXI4XL \D_cache/U2374  ( .A(\D_cache/cache[0][116] ), .B(
        \D_cache/cache[1][116] ), .C(\D_cache/cache[2][116] ), .D(
        \D_cache/cache[3][116] ), .S0(n2113), .S1(n2375), .Y(\D_cache/n2029 )
         );
  MXI4XL \D_cache/U2373  ( .A(\D_cache/cache[4][116] ), .B(
        \D_cache/cache[5][116] ), .C(\D_cache/cache[6][116] ), .D(
        \D_cache/cache[7][116] ), .S0(n2086), .S1(n2182), .Y(\D_cache/n2030 )
         );
  MXI2XL \D_cache/U2102  ( .A(\D_cache/n2029 ), .B(\D_cache/n2030 ), .S0(n3063), .Y(\D_cache/N68 ) );
  MXI4XL \D_cache/U2360  ( .A(\D_cache/cache[0][109] ), .B(
        \D_cache/cache[1][109] ), .C(\D_cache/cache[2][109] ), .D(
        \D_cache/cache[3][109] ), .S0(n2079), .S1(n2195), .Y(\D_cache/n2015 )
         );
  MXI4XL \D_cache/U2359  ( .A(\D_cache/cache[4][109] ), .B(
        \D_cache/cache[5][109] ), .C(\D_cache/cache[6][109] ), .D(
        \D_cache/cache[7][109] ), .S0(n2070), .S1(n2196), .Y(\D_cache/n2016 )
         );
  MXI2XL \D_cache/U2095  ( .A(\D_cache/n2015 ), .B(\D_cache/n2016 ), .S0(n3062), .Y(\D_cache/N75 ) );
  MXI4XL \D_cache/U2393  ( .A(\D_cache/cache[4][126] ), .B(
        \D_cache/cache[5][126] ), .C(\D_cache/cache[6][126] ), .D(
        \D_cache/cache[7][126] ), .S0(n2138), .S1(n2418), .Y(\D_cache/n2050 )
         );
  MXI4XL \D_cache/U2394  ( .A(\D_cache/cache[0][126] ), .B(
        \D_cache/cache[1][126] ), .C(\D_cache/cache[2][126] ), .D(
        \D_cache/cache[3][126] ), .S0(n2079), .S1(n2419), .Y(\D_cache/n2049 )
         );
  MXI2XL \D_cache/U2112  ( .A(\D_cache/n2049 ), .B(\D_cache/n2050 ), .S0(n4041), .Y(\D_cache/N58 ) );
  MXI4XL \D_cache/U2381  ( .A(\D_cache/cache[4][120] ), .B(
        \D_cache/cache[5][120] ), .C(\D_cache/cache[6][120] ), .D(
        \D_cache/cache[7][120] ), .S0(n2107), .S1(n2422), .Y(\D_cache/n2038 )
         );
  MXI4XL \D_cache/U2382  ( .A(\D_cache/cache[0][120] ), .B(
        \D_cache/cache[1][120] ), .C(\D_cache/cache[2][120] ), .D(
        \D_cache/cache[3][120] ), .S0(n2096), .S1(n2423), .Y(\D_cache/n2037 )
         );
  MXI2XL \D_cache/U2106  ( .A(\D_cache/n2037 ), .B(\D_cache/n2038 ), .S0(n2146), .Y(\D_cache/N64 ) );
  MXI4XL \D_cache/U2387  ( .A(\D_cache/cache[4][123] ), .B(
        \D_cache/cache[5][123] ), .C(\D_cache/cache[6][123] ), .D(
        \D_cache/cache[7][123] ), .S0(n2078), .S1(n2267), .Y(\D_cache/n2044 )
         );
  MXI4XL \D_cache/U2388  ( .A(\D_cache/cache[0][123] ), .B(
        \D_cache/cache[1][123] ), .C(\D_cache/cache[2][123] ), .D(
        \D_cache/cache[3][123] ), .S0(n2075), .S1(n2269), .Y(\D_cache/n2043 )
         );
  MXI2XL \D_cache/U2109  ( .A(\D_cache/n2043 ), .B(\D_cache/n2044 ), .S0(n4041), .Y(\D_cache/N61 ) );
  MXI4XL \D_cache/U2375  ( .A(\D_cache/cache[4][117] ), .B(
        \D_cache/cache[5][117] ), .C(\D_cache/cache[6][117] ), .D(
        \D_cache/cache[7][117] ), .S0(n2099), .S1(n2243), .Y(\D_cache/n2032 )
         );
  MXI4XL \D_cache/U2376  ( .A(\D_cache/cache[0][117] ), .B(
        \D_cache/cache[1][117] ), .C(\D_cache/cache[2][117] ), .D(
        \D_cache/cache[3][117] ), .S0(n2106), .S1(n2245), .Y(\D_cache/n2031 )
         );
  MXI2XL \D_cache/U2103  ( .A(\D_cache/n2031 ), .B(\D_cache/n2032 ), .S0(
        DCACHE_addr[4]), .Y(\D_cache/N67 ) );
  MXI4XL \D_cache/U2447  ( .A(\D_cache/cache[4][153] ), .B(
        \D_cache/cache[5][153] ), .C(\D_cache/cache[6][153] ), .D(
        \D_cache/cache[7][153] ), .S0(n2134), .S1(n2410), .Y(\D_cache/n2104 )
         );
  MXI4XL \D_cache/U2448  ( .A(\D_cache/cache[0][153] ), .B(
        \D_cache/cache[1][153] ), .C(\D_cache/cache[2][153] ), .D(
        \D_cache/cache[3][153] ), .S0(n2135), .S1(n2325), .Y(\D_cache/n2103 )
         );
  MXI2XL \D_cache/U2139  ( .A(\D_cache/n2103 ), .B(\D_cache/n2104 ), .S0(
        DCACHE_addr[4]), .Y(\D_cache/N31 ) );
  MXI4XL \D_cache/U2361  ( .A(\D_cache/cache[4][110] ), .B(
        \D_cache/cache[5][110] ), .C(\D_cache/cache[6][110] ), .D(
        \D_cache/cache[7][110] ), .S0(n2065), .S1(n2388), .Y(\D_cache/n2018 )
         );
  MXI4XL \D_cache/U2362  ( .A(\D_cache/cache[0][110] ), .B(
        \D_cache/cache[1][110] ), .C(\D_cache/cache[2][110] ), .D(
        \D_cache/cache[3][110] ), .S0(n2143), .S1(n2389), .Y(\D_cache/n2017 )
         );
  MXI2XL \D_cache/U2096  ( .A(\D_cache/n2017 ), .B(\D_cache/n2018 ), .S0(n3065), .Y(\D_cache/N74 ) );
  MXI4XL \D_cache/U2367  ( .A(\D_cache/cache[4][113] ), .B(
        \D_cache/cache[5][113] ), .C(\D_cache/cache[6][113] ), .D(
        \D_cache/cache[7][113] ), .S0(n2085), .S1(n2207), .Y(\D_cache/n2024 )
         );
  MXI4XL \D_cache/U2368  ( .A(\D_cache/cache[0][113] ), .B(
        \D_cache/cache[1][113] ), .C(\D_cache/cache[2][113] ), .D(
        \D_cache/cache[3][113] ), .S0(n2078), .S1(n2208), .Y(\D_cache/n2023 )
         );
  MXI2XL \D_cache/U2099  ( .A(\D_cache/n2023 ), .B(\D_cache/n2024 ), .S0(n3064), .Y(\D_cache/N71 ) );
  MXI4XL \D_cache/U2378  ( .A(\D_cache/cache[0][118] ), .B(
        \D_cache/cache[1][118] ), .C(\D_cache/cache[2][118] ), .D(
        \D_cache/cache[3][118] ), .S0(n2121), .S1(n2175), .Y(\D_cache/n2033 )
         );
  MXI4XL \D_cache/U2377  ( .A(\D_cache/cache[4][118] ), .B(
        \D_cache/cache[5][118] ), .C(\D_cache/cache[6][118] ), .D(
        \D_cache/cache[7][118] ), .S0(n2099), .S1(n2174), .Y(\D_cache/n2034 )
         );
  MXI4XL \D_cache/U2204  ( .A(\D_cache/cache[0][31] ), .B(
        \D_cache/cache[1][31] ), .C(\D_cache/cache[2][31] ), .D(
        \D_cache/cache[3][31] ), .S0(n2125), .S1(n2199), .Y(\D_cache/n1859 )
         );
  MXI4XL \D_cache/U2203  ( .A(\D_cache/cache[4][31] ), .B(
        \D_cache/cache[5][31] ), .C(\D_cache/cache[6][31] ), .D(
        \D_cache/cache[7][31] ), .S0(n2104), .S1(n2198), .Y(\D_cache/n1860 )
         );
  MXI2XL \D_cache/U2017  ( .A(\D_cache/n1859 ), .B(\D_cache/n1860 ), .S0(n3062), .Y(\D_cache/N153 ) );
  MXI4XL \D_cache/U2175  ( .A(\D_cache/cache[4][17] ), .B(
        \D_cache/cache[5][17] ), .C(\D_cache/cache[6][17] ), .D(
        \D_cache/cache[7][17] ), .S0(n2093), .S1(n2329), .Y(\D_cache/n1832 )
         );
  MXI4XL \D_cache/U2176  ( .A(\D_cache/cache[0][17] ), .B(
        \D_cache/cache[1][17] ), .C(\D_cache/cache[2][17] ), .D(
        \D_cache/cache[3][17] ), .S0(n2068), .S1(n2328), .Y(\D_cache/n1831 )
         );
  MXI4XL \D_cache/U2196  ( .A(\D_cache/cache[0][27] ), .B(
        \D_cache/cache[1][27] ), .C(\D_cache/cache[2][27] ), .D(
        \D_cache/cache[3][27] ), .S0(n2094), .S1(n2369), .Y(\D_cache/n1851 )
         );
  MXI4XL \D_cache/U2195  ( .A(\D_cache/cache[4][27] ), .B(
        \D_cache/cache[5][27] ), .C(\D_cache/cache[6][27] ), .D(
        \D_cache/cache[7][27] ), .S0(n2095), .S1(n2374), .Y(\D_cache/n1852 )
         );
  MXI4XL \D_cache/U2197  ( .A(\D_cache/cache[4][28] ), .B(
        \D_cache/cache[5][28] ), .C(\D_cache/cache[6][28] ), .D(
        \D_cache/cache[7][28] ), .S0(n2103), .S1(n2366), .Y(\D_cache/n1854 )
         );
  MXI4XL \D_cache/U2198  ( .A(\D_cache/cache[0][28] ), .B(
        \D_cache/cache[1][28] ), .C(\D_cache/cache[2][28] ), .D(
        \D_cache/cache[3][28] ), .S0(n2067), .S1(n2367), .Y(\D_cache/n1853 )
         );
  MXI2XL \D_cache/U2014  ( .A(\D_cache/n1853 ), .B(\D_cache/n1854 ), .S0(n3066), .Y(\D_cache/N156 ) );
  MXI4XL \D_cache/U2185  ( .A(\D_cache/cache[4][22] ), .B(
        \D_cache/cache[5][22] ), .C(\D_cache/cache[6][22] ), .D(
        \D_cache/cache[7][22] ), .S0(n2069), .S1(n2202), .Y(\D_cache/n1842 )
         );
  MXI4XL \D_cache/U2186  ( .A(\D_cache/cache[0][22] ), .B(
        \D_cache/cache[1][22] ), .C(\D_cache/cache[2][22] ), .D(
        \D_cache/cache[3][22] ), .S0(n2071), .S1(n2203), .Y(\D_cache/n1841 )
         );
  MXI2XL \D_cache/U2008  ( .A(\D_cache/n1841 ), .B(\D_cache/n1842 ), .S0(n4041), .Y(\D_cache/N162 ) );
  MXI4XL \D_cache/U2179  ( .A(\D_cache/cache[4][19] ), .B(
        \D_cache/cache[5][19] ), .C(\D_cache/cache[6][19] ), .D(
        \D_cache/cache[7][19] ), .S0(n2068), .S1(n2340), .Y(\D_cache/n1836 )
         );
  MXI4XL \D_cache/U2180  ( .A(\D_cache/cache[0][19] ), .B(
        \D_cache/cache[1][19] ), .C(\D_cache/cache[2][19] ), .D(
        \D_cache/cache[3][19] ), .S0(n2065), .S1(n2333), .Y(\D_cache/n1835 )
         );
  MXI4XL \D_cache/U2167  ( .A(\D_cache/cache[4][13] ), .B(
        \D_cache/cache[5][13] ), .C(\D_cache/cache[6][13] ), .D(
        \D_cache/cache[7][13] ), .S0(n2100), .S1(n2335), .Y(\D_cache/n1824 )
         );
  MXI4XL \D_cache/U2168  ( .A(\D_cache/cache[0][13] ), .B(
        \D_cache/cache[1][13] ), .C(\D_cache/cache[2][13] ), .D(
        \D_cache/cache[3][13] ), .S0(n2092), .S1(n2342), .Y(\D_cache/n1823 )
         );
  MXI4XL \D_cache/U2191  ( .A(\D_cache/cache[4][25] ), .B(
        \D_cache/cache[5][25] ), .C(\D_cache/cache[6][25] ), .D(
        \D_cache/cache[7][25] ), .S0(n2111), .S1(n2358), .Y(\D_cache/n1848 )
         );
  MXI4XL \D_cache/U2192  ( .A(\D_cache/cache[0][25] ), .B(
        \D_cache/cache[1][25] ), .C(\D_cache/cache[2][25] ), .D(
        \D_cache/cache[3][25] ), .S0(n2083), .S1(n2323), .Y(\D_cache/n1847 )
         );
  MXI4XL \D_cache/U2199  ( .A(\D_cache/cache[4][29] ), .B(
        \D_cache/cache[5][29] ), .C(\D_cache/cache[6][29] ), .D(
        \D_cache/cache[7][29] ), .S0(n2112), .S1(n2182), .Y(\D_cache/n1856 )
         );
  MXI4XL \D_cache/U2200  ( .A(\D_cache/cache[0][29] ), .B(
        \D_cache/cache[1][29] ), .C(\D_cache/cache[2][29] ), .D(
        \D_cache/cache[3][29] ), .S0(n2067), .S1(n2186), .Y(\D_cache/n1855 )
         );
  MXI4XL \D_cache/U2395  ( .A(\D_cache/cache[4][127] ), .B(
        \D_cache/cache[5][127] ), .C(\D_cache/cache[6][127] ), .D(
        \D_cache/cache[7][127] ), .S0(n2136), .S1(n2201), .Y(\D_cache/n2052 )
         );
  MXI4XL \D_cache/U2396  ( .A(\D_cache/cache[0][127] ), .B(
        \D_cache/cache[1][127] ), .C(\D_cache/cache[2][127] ), .D(
        \D_cache/cache[3][127] ), .S0(n2142), .S1(n2402), .Y(\D_cache/n2051 )
         );
  MXI2XL \D_cache/U2113  ( .A(\D_cache/n2051 ), .B(\D_cache/n2052 ), .S0(n2146), .Y(\D_cache/N57 ) );
  MXI4XL \D_cache/U2389  ( .A(\D_cache/cache[4][124] ), .B(
        \D_cache/cache[5][124] ), .C(\D_cache/cache[6][124] ), .D(
        \D_cache/cache[7][124] ), .S0(n2064), .S1(n2411), .Y(\D_cache/n2046 )
         );
  MXI4XL \D_cache/U2390  ( .A(\D_cache/cache[0][124] ), .B(
        \D_cache/cache[1][124] ), .C(\D_cache/cache[2][124] ), .D(
        \D_cache/cache[3][124] ), .S0(n2069), .S1(n2412), .Y(\D_cache/n2045 )
         );
  MXI2XL \D_cache/U2110  ( .A(\D_cache/n2045 ), .B(\D_cache/n2046 ), .S0(n3063), .Y(\D_cache/N60 ) );
  MXI4XL \D_cache/U2383  ( .A(\D_cache/cache[4][121] ), .B(
        \D_cache/cache[5][121] ), .C(\D_cache/cache[6][121] ), .D(
        \D_cache/cache[7][121] ), .S0(n2084), .S1(n2274), .Y(\D_cache/n2040 )
         );
  MXI4XL \D_cache/U2384  ( .A(\D_cache/cache[0][121] ), .B(
        \D_cache/cache[1][121] ), .C(\D_cache/cache[2][121] ), .D(
        \D_cache/cache[3][121] ), .S0(n2108), .S1(n2276), .Y(\D_cache/n2039 )
         );
  MXI2XL \D_cache/U2107  ( .A(\D_cache/n2039 ), .B(\D_cache/n2040 ), .S0(n3065), .Y(\D_cache/N63 ) );
  MXI4XL \D_cache/U2291  ( .A(\D_cache/cache[4][75] ), .B(
        \D_cache/cache[5][75] ), .C(\D_cache/cache[6][75] ), .D(
        \D_cache/cache[7][75] ), .S0(n2119), .S1(n2201), .Y(\D_cache/n1948 )
         );
  MXI4XL \D_cache/U2292  ( .A(\D_cache/cache[0][75] ), .B(
        \D_cache/cache[1][75] ), .C(\D_cache/cache[2][75] ), .D(
        \D_cache/cache[3][75] ), .S0(n2120), .S1(n2182), .Y(\D_cache/n1947 )
         );
  MXI2XL \D_cache/U2061  ( .A(\D_cache/n1947 ), .B(\D_cache/n1948 ), .S0(n2147), .Y(\D_cache/N109 ) );
  MXI4XL \D_cache/U2285  ( .A(\D_cache/cache[4][72] ), .B(
        \D_cache/cache[5][72] ), .C(\D_cache/cache[6][72] ), .D(
        \D_cache/cache[7][72] ), .S0(n2098), .S1(n2237), .Y(\D_cache/n1942 )
         );
  MXI4XL \D_cache/U2286  ( .A(\D_cache/cache[0][72] ), .B(
        \D_cache/cache[1][72] ), .C(\D_cache/cache[2][72] ), .D(
        \D_cache/cache[3][72] ), .S0(n2078), .S1(n2246), .Y(\D_cache/n1941 )
         );
  MXI4XL \D_cache/U2363  ( .A(\D_cache/cache[4][111] ), .B(
        \D_cache/cache[5][111] ), .C(\D_cache/cache[6][111] ), .D(
        \D_cache/cache[7][111] ), .S0(n2073), .S1(n2211), .Y(\D_cache/n2020 )
         );
  MXI4XL \D_cache/U2364  ( .A(\D_cache/cache[0][111] ), .B(
        \D_cache/cache[1][111] ), .C(\D_cache/cache[2][111] ), .D(
        \D_cache/cache[3][111] ), .S0(n2074), .S1(n2212), .Y(\D_cache/n2019 )
         );
  MXI2XL \D_cache/U2097  ( .A(\D_cache/n2019 ), .B(\D_cache/n2020 ), .S0(
        DCACHE_addr[4]), .Y(\D_cache/N73 ) );
  MXI4XL \D_cache/U2369  ( .A(\D_cache/cache[4][114] ), .B(
        \D_cache/cache[5][114] ), .C(\D_cache/cache[6][114] ), .D(
        \D_cache/cache[7][114] ), .S0(n2081), .S1(n2293), .Y(\D_cache/n2026 )
         );
  MXI4XL \D_cache/U2370  ( .A(\D_cache/cache[0][114] ), .B(
        \D_cache/cache[1][114] ), .C(\D_cache/cache[2][114] ), .D(
        \D_cache/cache[3][114] ), .S0(n2134), .S1(n2297), .Y(\D_cache/n2025 )
         );
  MXI2XL \D_cache/U2100  ( .A(\D_cache/n2025 ), .B(\D_cache/n2026 ), .S0(n2147), .Y(\D_cache/N70 ) );
  MXI4XL \D_cache/U2289  ( .A(\D_cache/cache[4][74] ), .B(
        \D_cache/cache[5][74] ), .C(\D_cache/cache[6][74] ), .D(
        \D_cache/cache[7][74] ), .S0(n2139), .S1(n2252), .Y(\D_cache/n1946 )
         );
  MXI4XL \D_cache/U2290  ( .A(\D_cache/cache[0][74] ), .B(
        \D_cache/cache[1][74] ), .C(\D_cache/cache[2][74] ), .D(
        \D_cache/cache[3][74] ), .S0(n2143), .S1(n2266), .Y(\D_cache/n1945 )
         );
  MXI4XL \D_cache/U2283  ( .A(\D_cache/cache[4][71] ), .B(
        \D_cache/cache[5][71] ), .C(\D_cache/cache[6][71] ), .D(
        \D_cache/cache[7][71] ), .S0(n2080), .S1(n2302), .Y(\D_cache/n1940 )
         );
  MXI4XL \D_cache/U2284  ( .A(\D_cache/cache[0][71] ), .B(
        \D_cache/cache[1][71] ), .C(\D_cache/cache[2][71] ), .D(
        \D_cache/cache[3][71] ), .S0(n2111), .S1(n2360), .Y(\D_cache/n1939 )
         );
  MXI4XL \D_cache/U2277  ( .A(\D_cache/cache[4][68] ), .B(
        \D_cache/cache[5][68] ), .C(\D_cache/cache[6][68] ), .D(
        \D_cache/cache[7][68] ), .S0(n2132), .S1(n2188), .Y(\D_cache/n1934 )
         );
  MXI4XL \D_cache/U2278  ( .A(\D_cache/cache[0][68] ), .B(
        \D_cache/cache[1][68] ), .C(\D_cache/cache[2][68] ), .D(
        \D_cache/cache[3][68] ), .S0(n2120), .S1(n2194), .Y(\D_cache/n1933 )
         );
  MXI4XL \D_cache/U2287  ( .A(\D_cache/cache[4][73] ), .B(
        \D_cache/cache[5][73] ), .C(\D_cache/cache[6][73] ), .D(
        \D_cache/cache[7][73] ), .S0(n2065), .S1(n2341), .Y(\D_cache/n1944 )
         );
  MXI4XL \D_cache/U2288  ( .A(\D_cache/cache[0][73] ), .B(
        \D_cache/cache[1][73] ), .C(\D_cache/cache[2][73] ), .D(
        \D_cache/cache[3][73] ), .S0(n2062), .S1(n2354), .Y(\D_cache/n1943 )
         );
  MXI4XL \D_cache/U2201  ( .A(\D_cache/cache[4][30] ), .B(
        \D_cache/cache[5][30] ), .C(\D_cache/cache[6][30] ), .D(
        \D_cache/cache[7][30] ), .S0(n2103), .S1(n2368), .Y(\D_cache/n1858 )
         );
  MXI4XL \D_cache/U2202  ( .A(\D_cache/cache[0][30] ), .B(
        \D_cache/cache[1][30] ), .C(\D_cache/cache[2][30] ), .D(
        \D_cache/cache[3][30] ), .S0(n2133), .S1(n2226), .Y(\D_cache/n1857 )
         );
  MXI2XL \D_cache/U2016  ( .A(\D_cache/n1857 ), .B(\D_cache/n1858 ), .S0(n3066), .Y(\D_cache/N154 ) );
  MXI4XL \D_cache/U2190  ( .A(\D_cache/cache[0][24] ), .B(
        \D_cache/cache[1][24] ), .C(\D_cache/cache[2][24] ), .D(
        \D_cache/cache[3][24] ), .S0(n2141), .S1(n2414), .Y(\D_cache/n1845 )
         );
  MXI4XL \D_cache/U2189  ( .A(\D_cache/cache[4][24] ), .B(
        \D_cache/cache[5][24] ), .C(\D_cache/cache[6][24] ), .D(
        \D_cache/cache[7][24] ), .S0(n2140), .S1(n2413), .Y(\D_cache/n1846 )
         );
  MXI4XL \D_cache/U2184  ( .A(\D_cache/cache[0][21] ), .B(
        \D_cache/cache[1][21] ), .C(\D_cache/cache[2][21] ), .D(
        \D_cache/cache[3][21] ), .S0(n2124), .S1(n2421), .Y(\D_cache/n1839 )
         );
  MXI4XL \D_cache/U2183  ( .A(\D_cache/cache[4][21] ), .B(
        \D_cache/cache[5][21] ), .C(\D_cache/cache[6][21] ), .D(
        \D_cache/cache[7][21] ), .S0(n2123), .S1(n2387), .Y(\D_cache/n1840 )
         );
  MXI4XL \D_cache/U2148  ( .A(\D_cache/cache[0][3] ), .B(\D_cache/cache[1][3] ), .C(\D_cache/cache[2][3] ), .D(\D_cache/cache[3][3] ), .S0(DCACHE_addr[2]), 
        .S1(n2227), .Y(\D_cache/n1803 ) );
  MXI4XL \D_cache/U2147  ( .A(\D_cache/cache[4][3] ), .B(\D_cache/cache[5][3] ), .C(\D_cache/cache[6][3] ), .D(\D_cache/cache[7][3] ), .S0(n2139), .S1(n2363), 
        .Y(\D_cache/n1804 ) );
  MXI4XL \D_cache/U2163  ( .A(\D_cache/cache[4][11] ), .B(
        \D_cache/cache[5][11] ), .C(\D_cache/cache[6][11] ), .D(
        \D_cache/cache[7][11] ), .S0(n2131), .S1(DCACHE_addr[3]), .Y(
        \D_cache/n1820 ) );
  MXI4XL \D_cache/U2164  ( .A(\D_cache/cache[0][11] ), .B(
        \D_cache/cache[1][11] ), .C(\D_cache/cache[2][11] ), .D(
        \D_cache/cache[3][11] ), .S0(n2112), .S1(n2219), .Y(\D_cache/n1819 )
         );
  MXI4XL \D_cache/U2193  ( .A(\D_cache/cache[4][26] ), .B(
        \D_cache/cache[5][26] ), .C(\D_cache/cache[6][26] ), .D(
        \D_cache/cache[7][26] ), .S0(n2132), .S1(n2378), .Y(\D_cache/n1850 )
         );
  MXI4XL \D_cache/U2194  ( .A(\D_cache/cache[0][26] ), .B(
        \D_cache/cache[1][26] ), .C(\D_cache/cache[2][26] ), .D(
        \D_cache/cache[3][26] ), .S0(n2133), .S1(n2384), .Y(\D_cache/n1849 )
         );
  MXI4XL \D_cache/U2348  ( .A(\D_cache/cache[0][103] ), .B(
        \D_cache/cache[1][103] ), .C(\D_cache/cache[2][103] ), .D(
        \D_cache/cache[3][103] ), .S0(n2115), .S1(n2284), .Y(\D_cache/n2003 )
         );
  MXI4XL \D_cache/U2347  ( .A(\D_cache/cache[4][103] ), .B(
        \D_cache/cache[5][103] ), .C(\D_cache/cache[6][103] ), .D(
        \D_cache/cache[7][103] ), .S0(n2105), .S1(n2261), .Y(\D_cache/n2004 )
         );
  MXI4XL \D_cache/U2351  ( .A(\D_cache/cache[4][105] ), .B(
        \D_cache/cache[5][105] ), .C(\D_cache/cache[6][105] ), .D(
        \D_cache/cache[7][105] ), .S0(n2063), .S1(n2187), .Y(\D_cache/n2008 )
         );
  MXI4XL \D_cache/U2352  ( .A(\D_cache/cache[0][105] ), .B(
        \D_cache/cache[1][105] ), .C(\D_cache/cache[2][105] ), .D(
        \D_cache/cache[3][105] ), .S0(n2144), .S1(n2189), .Y(\D_cache/n2007 )
         );
  MXI2XL \D_cache/U2091  ( .A(\D_cache/n2007 ), .B(\D_cache/n2008 ), .S0(n3063), .Y(\D_cache/N79 ) );
  MXI4XL \D_cache/U2301  ( .A(\D_cache/cache[4][80] ), .B(
        \D_cache/cache[5][80] ), .C(\D_cache/cache[6][80] ), .D(
        \D_cache/cache[7][80] ), .S0(n2142), .S1(n2343), .Y(\D_cache/n1958 )
         );
  MXI4XL \D_cache/U2302  ( .A(\D_cache/cache[0][80] ), .B(
        \D_cache/cache[1][80] ), .C(\D_cache/cache[2][80] ), .D(
        \D_cache/cache[3][80] ), .S0(n2139), .S1(n2345), .Y(\D_cache/n1957 )
         );
  MXI4XL \D_cache/U2315  ( .A(\D_cache/cache[4][87] ), .B(
        \D_cache/cache[5][87] ), .C(\D_cache/cache[6][87] ), .D(
        \D_cache/cache[7][87] ), .S0(n2137), .S1(n2341), .Y(\D_cache/n1972 )
         );
  MXI4XL \D_cache/U2316  ( .A(\D_cache/cache[0][87] ), .B(
        \D_cache/cache[1][87] ), .C(\D_cache/cache[2][87] ), .D(
        \D_cache/cache[3][87] ), .S0(n2139), .S1(n2349), .Y(\D_cache/n1971 )
         );
  MXI4XL \D_cache/U2345  ( .A(\D_cache/cache[4][102] ), .B(
        \D_cache/cache[5][102] ), .C(\D_cache/cache[6][102] ), .D(
        \D_cache/cache[7][102] ), .S0(n2097), .S1(n2376), .Y(\D_cache/n2002 )
         );
  MXI4XL \D_cache/U2346  ( .A(\D_cache/cache[0][102] ), .B(
        \D_cache/cache[1][102] ), .C(\D_cache/cache[2][102] ), .D(
        \D_cache/cache[3][102] ), .S0(n2124), .S1(n2379), .Y(\D_cache/n2001 )
         );
  MXI4XL \D_cache/U2271  ( .A(\D_cache/cache[4][65] ), .B(
        \D_cache/cache[5][65] ), .C(\D_cache/cache[6][65] ), .D(
        \D_cache/cache[7][65] ), .S0(n2131), .S1(n2322), .Y(\D_cache/n1928 )
         );
  MXI4XL \D_cache/U2272  ( .A(\D_cache/cache[0][65] ), .B(
        \D_cache/cache[1][65] ), .C(\D_cache/cache[2][65] ), .D(
        \D_cache/cache[3][65] ), .S0(n2136), .S1(n2327), .Y(\D_cache/n1927 )
         );
  MXI4XL \D_cache/U2269  ( .A(\D_cache/cache[4][64] ), .B(
        \D_cache/cache[5][64] ), .C(\D_cache/cache[6][64] ), .D(
        \D_cache/cache[7][64] ), .S0(n2066), .S1(n2426), .Y(\D_cache/n1926 )
         );
  MXI4XL \D_cache/U2270  ( .A(\D_cache/cache[0][64] ), .B(
        \D_cache/cache[1][64] ), .C(\D_cache/cache[2][64] ), .D(
        \D_cache/cache[3][64] ), .S0(n2063), .S1(n2436), .Y(\D_cache/n1925 )
         );
  MXI4XL \D_cache/U2380  ( .A(\D_cache/cache[0][119] ), .B(
        \D_cache/cache[1][119] ), .C(\D_cache/cache[2][119] ), .D(
        \D_cache/cache[3][119] ), .S0(n2092), .S1(n2381), .Y(\D_cache/n2035 )
         );
  MXI4XL \D_cache/U2379  ( .A(\D_cache/cache[4][119] ), .B(
        \D_cache/cache[5][119] ), .C(\D_cache/cache[6][119] ), .D(
        \D_cache/cache[7][119] ), .S0(n2067), .S1(n2380), .Y(\D_cache/n2036 )
         );
  MXI2XL \D_cache/U2105  ( .A(\D_cache/n2035 ), .B(\D_cache/n2036 ), .S0(n3065), .Y(\D_cache/N65 ) );
  MXI4XL \D_cache/U2366  ( .A(\D_cache/cache[0][112] ), .B(
        \D_cache/cache[1][112] ), .C(\D_cache/cache[2][112] ), .D(
        \D_cache/cache[3][112] ), .S0(n2072), .S1(n2194), .Y(\D_cache/n2021 )
         );
  MXI4XL \D_cache/U2365  ( .A(\D_cache/cache[4][112] ), .B(
        \D_cache/cache[5][112] ), .C(\D_cache/cache[6][112] ), .D(
        \D_cache/cache[7][112] ), .S0(n2075), .S1(n2188), .Y(\D_cache/n2022 )
         );
  MXI2XL \D_cache/U2098  ( .A(\D_cache/n2021 ), .B(\D_cache/n2022 ), .S0(n4041), .Y(\D_cache/N72 ) );
  MXI4XL \D_cache/U2279  ( .A(\D_cache/cache[4][69] ), .B(
        \D_cache/cache[5][69] ), .C(\D_cache/cache[6][69] ), .D(
        \D_cache/cache[7][69] ), .S0(n2139), .S1(n2307), .Y(\D_cache/n1936 )
         );
  MXI4XL \D_cache/U2280  ( .A(\D_cache/cache[0][69] ), .B(
        \D_cache/cache[1][69] ), .C(\D_cache/cache[2][69] ), .D(
        \D_cache/cache[3][69] ), .S0(n2142), .S1(n2317), .Y(\D_cache/n1935 )
         );
  MXI4XL \D_cache/U2161  ( .A(\D_cache/cache[4][10] ), .B(
        \D_cache/cache[5][10] ), .C(\D_cache/cache[6][10] ), .D(
        \D_cache/cache[7][10] ), .S0(n2139), .S1(n2250), .Y(\D_cache/n1818 )
         );
  MXI4XL \D_cache/U2162  ( .A(\D_cache/cache[0][10] ), .B(
        \D_cache/cache[1][10] ), .C(\D_cache/cache[2][10] ), .D(
        \D_cache/cache[3][10] ), .S0(n2143), .S1(n2249), .Y(\D_cache/n1817 )
         );
  MXI4XL \D_cache/U2173  ( .A(\D_cache/cache[4][16] ), .B(
        \D_cache/cache[5][16] ), .C(\D_cache/cache[6][16] ), .D(
        \D_cache/cache[7][16] ), .S0(n2076), .S1(n2309), .Y(\D_cache/n1830 )
         );
  MXI4XL \D_cache/U2174  ( .A(\D_cache/cache[0][16] ), .B(
        \D_cache/cache[1][16] ), .C(\D_cache/cache[2][16] ), .D(
        \D_cache/cache[3][16] ), .S0(n2101), .S1(n2318), .Y(\D_cache/n1829 )
         );
  MXI4XL \D_cache/U2281  ( .A(\D_cache/cache[4][70] ), .B(
        \D_cache/cache[5][70] ), .C(\D_cache/cache[6][70] ), .D(
        \D_cache/cache[7][70] ), .S0(n2141), .S1(n2386), .Y(\D_cache/n1938 )
         );
  MXI4XL \D_cache/U2282  ( .A(\D_cache/cache[0][70] ), .B(
        \D_cache/cache[1][70] ), .C(\D_cache/cache[2][70] ), .D(
        \D_cache/cache[3][70] ), .S0(n2106), .S1(n2417), .Y(\D_cache/n1937 )
         );
  MXI4XL \D_cache/U2443  ( .A(\D_cache/cache[4][151] ), .B(
        \D_cache/cache[5][151] ), .C(\D_cache/cache[6][151] ), .D(
        \D_cache/cache[7][151] ), .S0(n2130), .S1(n2434), .Y(\D_cache/n2100 )
         );
  MXI4XL \D_cache/U2444  ( .A(\D_cache/cache[0][151] ), .B(
        \D_cache/cache[1][151] ), .C(\D_cache/cache[2][151] ), .D(
        \D_cache/cache[3][151] ), .S0(n2137), .S1(n2437), .Y(\D_cache/n2099 )
         );
  MXI4XL \D_cache/U2415  ( .A(\D_cache/cache[4][137] ), .B(
        \D_cache/cache[5][137] ), .C(\D_cache/cache[6][137] ), .D(
        \D_cache/cache[7][137] ), .S0(n2102), .S1(n2403), .Y(\D_cache/n2072 )
         );
  MXI4XL \D_cache/U2416  ( .A(\D_cache/cache[0][137] ), .B(
        \D_cache/cache[1][137] ), .C(\D_cache/cache[2][137] ), .D(
        \D_cache/cache[3][137] ), .S0(n2142), .S1(n2406), .Y(\D_cache/n2071 )
         );
  MXI4XL \D_cache/U2398  ( .A(\D_cache/cache[0][128] ), .B(
        \D_cache/cache[1][128] ), .C(\D_cache/cache[2][128] ), .D(
        \D_cache/cache[3][128] ), .S0(n2130), .S1(n2429), .Y(\D_cache/n2053 )
         );
  DFFRHQX8 \i_MIPS/EX_MEM_reg[9]  ( .D(\i_MIPS/n465 ), .CK(clk), .RN(n4055), 
        .Q(n2750) );
  MXI2X1 \D_cache/U2015  ( .A(\D_cache/n1855 ), .B(\D_cache/n1856 ), .S0(
        DCACHE_addr[4]), .Y(\D_cache/N155 ) );
  MXI4XL \D_cache/U2440  ( .A(\D_cache/cache[0][149] ), .B(
        \D_cache/cache[1][149] ), .C(\D_cache/cache[2][149] ), .D(
        \D_cache/cache[3][149] ), .S0(n2092), .S1(n2175), .Y(\D_cache/n2095 )
         );
  MXI4XL \D_cache/U2439  ( .A(\D_cache/cache[4][149] ), .B(
        \D_cache/cache[5][149] ), .C(\D_cache/cache[6][149] ), .D(
        \D_cache/cache[7][149] ), .S0(n2129), .S1(n2172), .Y(\D_cache/n2096 )
         );
  DFFRHQX8 \i_MIPS/EX_MEM_reg[10]  ( .D(\i_MIPS/n464 ), .CK(clk), .RN(n4055), 
        .Q(n2747) );
  DFFRX4 \i_MIPS/ID_EX_reg[80]  ( .D(\i_MIPS/n505 ), .CK(clk), .RN(n4058), .Q(
        \i_MIPS/ID_EX[80] ), .QN(n2988) );
  DFFRX1 \i_MIPS/EX_MEM_reg[18]  ( .D(\i_MIPS/n456 ), .CK(clk), .RN(n4054), 
        .Q(n10315), .QN(n1621) );
  DFFRHQX8 \i_MIPS/ID_EX_reg[8]  ( .D(\i_MIPS/n470 ), .CK(clk), .RN(n4055), 
        .Q(n2730) );
  DFFRX4 \i_MIPS/ID_EX_reg[73]  ( .D(\i_MIPS/n512 ), .CK(clk), .RN(n4059), .Q(
        \i_MIPS/ID_EX[73] ), .QN(n964) );
  DFFRX1 \i_MIPS/ID_EX_reg[38]  ( .D(\i_MIPS/n533 ), .CK(clk), .RN(n4063), .Q(
        \i_MIPS/ALUin1[29] ), .QN(\i_MIPS/n342 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[82]  ( .D(\i_MIPS/n503 ), .CK(clk), .RN(n4058), .Q(
        \i_MIPS/ID_EX[82] ), .QN(n2990) );
  DFFRX1 \i_MIPS/ID_EX_reg[46]  ( .D(\i_MIPS/n427 ), .CK(clk), .RN(n4051), .Q(
        n1884), .QN(\i_MIPS/n299 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[37]  ( .D(\i_MIPS/n534 ), .CK(clk), .RN(n4063), .Q(
        \i_MIPS/ALUin1[28] ), .QN(\i_MIPS/n343 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[57]  ( .D(\i_MIPS/N80 ), .CK(clk), .RN(n4061), .Q(
        \i_MIPS/IR_ID[25] ), .QN(\i_MIPS/n232 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[36]  ( .D(\i_MIPS/n535 ), .CK(clk), .RN(n4063), .Q(
        \i_MIPS/ALUin1[27] ), .QN(\i_MIPS/n344 ) );
  DFFRX4 \i_MIPS/EX_MEM_reg[11]  ( .D(\i_MIPS/n463 ), .CK(clk), .RN(n4054), 
        .Q(n10321), .QN(n2722) );
  DFFRX4 \i_MIPS/ID_EX_reg[5]  ( .D(\i_MIPS/n478 ), .CK(clk), .RN(n4056), .Q(
        \i_MIPS/ID_EX_5 ) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[1]  ( .D(\i_MIPS/PC/n35 ), .CK(clk), .RN(n4066), 
        .Q(\i_MIPS/PC_o[1] ), .QN(\i_MIPS/PC/n3 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[106]  ( .D(\i_MIPS/n519 ), .CK(clk), .RN(n4061), 
        .Q(\i_MIPS/ID_EX[106] ), .QN(\i_MIPS/n325 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[37]  ( .D(\i_MIPS/n436 ), .CK(clk), .RN(n4052), 
        .Q(n10355), .QN(\i_MIPS/n308 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[38]  ( .D(\i_MIPS/n434 ), .CK(clk), .RN(n4052), 
        .Q(n10354), .QN(\i_MIPS/n306 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[39]  ( .D(\i_MIPS/n432 ), .CK(clk), .RN(n4052), 
        .Q(n10353), .QN(\i_MIPS/n304 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[40]  ( .D(\i_MIPS/n430 ), .CK(clk), .RN(n4052), 
        .Q(n10352), .QN(\i_MIPS/n302 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[41]  ( .D(\i_MIPS/n428 ), .CK(clk), .RN(n4052), 
        .Q(n10351), .QN(\i_MIPS/n300 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[42]  ( .D(\i_MIPS/n426 ), .CK(clk), .RN(n4051), 
        .Q(n10350), .QN(\i_MIPS/n298 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[43]  ( .D(\i_MIPS/n424 ), .CK(clk), .RN(n4051), 
        .Q(n10349), .QN(\i_MIPS/n296 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[44]  ( .D(\i_MIPS/n422 ), .CK(clk), .RN(n4051), 
        .Q(n10348), .QN(\i_MIPS/n294 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[45]  ( .D(\i_MIPS/n420 ), .CK(clk), .RN(n4051), 
        .Q(n10347), .QN(\i_MIPS/n292 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[46]  ( .D(\i_MIPS/n418 ), .CK(clk), .RN(n4051), 
        .Q(n10346), .QN(\i_MIPS/n290 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[47]  ( .D(\i_MIPS/n416 ), .CK(clk), .RN(n4051), 
        .Q(n10345), .QN(\i_MIPS/n288 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[48]  ( .D(\i_MIPS/n414 ), .CK(clk), .RN(n4050), 
        .Q(n10344), .QN(\i_MIPS/n286 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[49]  ( .D(\i_MIPS/n412 ), .CK(clk), .RN(n4050), 
        .Q(n10343), .QN(\i_MIPS/n284 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[50]  ( .D(\i_MIPS/n410 ), .CK(clk), .RN(n4050), 
        .Q(n10342), .QN(\i_MIPS/n282 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[51]  ( .D(\i_MIPS/n408 ), .CK(clk), .RN(n4050), 
        .Q(n10341), .QN(\i_MIPS/n280 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[52]  ( .D(\i_MIPS/n406 ), .CK(clk), .RN(n4050), 
        .Q(n10340), .QN(\i_MIPS/n278 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[53]  ( .D(\i_MIPS/n404 ), .CK(clk), .RN(n4050), 
        .Q(n10339), .QN(\i_MIPS/n276 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[54]  ( .D(\i_MIPS/n402 ), .CK(clk), .RN(n4049), 
        .Q(n10338), .QN(\i_MIPS/n274 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[55]  ( .D(\i_MIPS/n400 ), .CK(clk), .RN(n4049), 
        .Q(n10337), .QN(\i_MIPS/n272 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[56]  ( .D(\i_MIPS/n398 ), .CK(clk), .RN(n4049), 
        .Q(n10336), .QN(\i_MIPS/n270 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[57]  ( .D(\i_MIPS/n396 ), .CK(clk), .RN(n4049), 
        .Q(n10335), .QN(\i_MIPS/n268 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[58]  ( .D(\i_MIPS/n394 ), .CK(clk), .RN(n4049), 
        .Q(n10334), .QN(\i_MIPS/n266 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[59]  ( .D(\i_MIPS/n392 ), .CK(clk), .RN(n4049), 
        .Q(n10333), .QN(\i_MIPS/n264 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[60]  ( .D(\i_MIPS/n390 ), .CK(clk), .RN(n4048), 
        .Q(n10332), .QN(\i_MIPS/n262 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[61]  ( .D(\i_MIPS/n388 ), .CK(clk), .RN(n4048), 
        .Q(n10331), .QN(\i_MIPS/n260 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[62]  ( .D(\i_MIPS/n386 ), .CK(clk), .RN(n4048), 
        .Q(n10330), .QN(\i_MIPS/n258 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[63]  ( .D(\i_MIPS/n384 ), .CK(clk), .RN(n4048), 
        .Q(n10329), .QN(\i_MIPS/n256 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[64]  ( .D(\i_MIPS/n382 ), .CK(clk), .RN(n4048), 
        .Q(n10328), .QN(\i_MIPS/n254 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[65]  ( .D(\i_MIPS/n380 ), .CK(clk), .RN(n4048), 
        .Q(n10327), .QN(\i_MIPS/n252 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[66]  ( .D(\i_MIPS/n378 ), .CK(clk), .RN(n4047), 
        .Q(n10326), .QN(\i_MIPS/n250 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[67]  ( .D(\i_MIPS/n376 ), .CK(clk), .RN(n4047), 
        .Q(n10325), .QN(\i_MIPS/n248 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[68]  ( .D(\i_MIPS/n374 ), .CK(clk), .RN(n4047), 
        .Q(n10324), .QN(\i_MIPS/n246 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[4]  ( .D(\i_MIPS/n479 ), .CK(clk), .RN(n4056), .Q(
        n10356), .QN(\i_MIPS/n310 ) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[24]  ( .D(\i_MIPS/PC/n58 ), .CK(clk), .RN(n4068), 
        .Q(ICACHE_addr[22]), .QN(\i_MIPS/PC/n26 ) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[26]  ( .D(\i_MIPS/PC/n60 ), .CK(clk), .RN(n4068), 
        .Q(ICACHE_addr[24]), .QN(\i_MIPS/PC/n28 ) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[29]  ( .D(\i_MIPS/PC/n63 ), .CK(clk), .RN(n4068), 
        .Q(ICACHE_addr[27]), .QN(\i_MIPS/PC/n31 ) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[18]  ( .D(\i_MIPS/PC/n52 ), .CK(clk), .RN(n4067), 
        .Q(ICACHE_addr[16]), .QN(\i_MIPS/PC/n20 ) );
  MXI2X2 \D_cache/U2135  ( .A(\D_cache/n2095 ), .B(\D_cache/n2096 ), .S0(n4041), .Y(\D_cache/N35 ) );
  MXI2X2 \D_cache/U2138  ( .A(\D_cache/n2101 ), .B(\D_cache/n2102 ), .S0(n2146), .Y(\D_cache/N32 ) );
  MXI2X2 \D_cache/U2120  ( .A(\D_cache/n2065 ), .B(\D_cache/n2066 ), .S0(n2147), .Y(\D_cache/N50 ) );
  MXI2X2 \D_cache/U2129  ( .A(\D_cache/n2083 ), .B(\D_cache/n2084 ), .S0(n2146), .Y(\D_cache/N41 ) );
  DFFRX4 \i_MIPS/PC/PC_o_reg[16]  ( .D(\i_MIPS/PC/n50 ), .CK(clk), .RN(n4067), 
        .Q(ICACHE_addr[14]), .QN(\i_MIPS/PC/n18 ) );
  DFFRX4 \i_MIPS/PC/PC_o_reg[8]  ( .D(\i_MIPS/PC/n42 ), .CK(clk), .RN(n4066), 
        .Q(ICACHE_addr[6]), .QN(\i_MIPS/PC/n10 ) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[27]  ( .D(\i_MIPS/PC/n61 ), .CK(clk), .RN(n4068), 
        .Q(ICACHE_addr[25]), .QN(\i_MIPS/PC/n29 ) );
  DFFRX4 \i_MIPS/PC/PC_o_reg[14]  ( .D(\i_MIPS/PC/n48 ), .CK(clk), .RN(n4067), 
        .Q(ICACHE_addr[12]), .QN(\i_MIPS/PC/n16 ) );
  DFFRX4 \i_MIPS/PC/PC_o_reg[11]  ( .D(\i_MIPS/PC/n45 ), .CK(clk), .RN(n4066), 
        .Q(ICACHE_addr[9]), .QN(\i_MIPS/PC/n13 ) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[22]  ( .D(\i_MIPS/PC/n56 ), .CK(clk), .RN(n4067), 
        .Q(ICACHE_addr[20]), .QN(\i_MIPS/PC/n24 ) );
  DFFRX4 \i_MIPS/PC/PC_o_reg[9]  ( .D(\i_MIPS/PC/n43 ), .CK(clk), .RN(n4066), 
        .Q(ICACHE_addr[7]), .QN(\i_MIPS/PC/n11 ) );
  DFFRX4 \i_MIPS/PC/PC_o_reg[13]  ( .D(\i_MIPS/PC/n47 ), .CK(clk), .RN(n4067), 
        .Q(ICACHE_addr[11]), .QN(\i_MIPS/PC/n15 ) );
  DFFRX4 \i_MIPS/PC/PC_o_reg[10]  ( .D(\i_MIPS/PC/n44 ), .CK(clk), .RN(n4066), 
        .Q(ICACHE_addr[8]), .QN(\i_MIPS/PC/n12 ) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[20]  ( .D(\i_MIPS/PC/n54 ), .CK(clk), .RN(n4067), 
        .Q(ICACHE_addr[18]), .QN(\i_MIPS/PC/n22 ) );
  DFFRX4 \i_MIPS/PC/PC_o_reg[17]  ( .D(\i_MIPS/PC/n51 ), .CK(clk), .RN(n4067), 
        .Q(ICACHE_addr[15]), .QN(\i_MIPS/PC/n19 ) );
  DFFRX4 \i_MIPS/PC/PC_o_reg[19]  ( .D(\i_MIPS/PC/n53 ), .CK(clk), .RN(n4067), 
        .Q(ICACHE_addr[17]), .QN(\i_MIPS/PC/n21 ) );
  MXI4X4 \D_cache/U2423  ( .A(\D_cache/cache[4][141] ), .B(
        \D_cache/cache[5][141] ), .C(\D_cache/cache[6][141] ), .D(
        \D_cache/cache[7][141] ), .S0(n2135), .S1(n2409), .Y(\D_cache/n2080 )
         );
  MXI2X4 \D_cache/U2127  ( .A(\D_cache/n2079 ), .B(\D_cache/n2080 ), .S0(n4041), .Y(\D_cache/N43 ) );
  MXI4X2 \D_cache/U2445  ( .A(\D_cache/cache[4][152] ), .B(
        \D_cache/cache[5][152] ), .C(\D_cache/cache[6][152] ), .D(
        \D_cache/cache[7][152] ), .S0(n2123), .S1(n2435), .Y(\D_cache/n2102 )
         );
  MXI4X1 \D_cache/U2412  ( .A(\D_cache/cache[0][135] ), .B(
        \D_cache/cache[1][135] ), .C(\D_cache/cache[2][135] ), .D(
        \D_cache/cache[3][135] ), .S0(n2144), .S1(n2401), .Y(\D_cache/n2067 )
         );
  DFFRX4 \i_MIPS/PC/PC_o_reg[0]  ( .D(\i_MIPS/PC/n34 ), .CK(clk), .RN(n4066), 
        .Q(\i_MIPS/BranchAddr[0] ), .QN(\i_MIPS/PC/n2 ) );
  MXI4X1 \D_cache/U2414  ( .A(\D_cache/cache[0][136] ), .B(
        \D_cache/cache[1][136] ), .C(\D_cache/cache[2][136] ), .D(
        \D_cache/cache[3][136] ), .S0(n2091), .S1(n2176), .Y(\D_cache/n2069 )
         );
  MXI4X1 \D_cache/U2413  ( .A(\D_cache/cache[4][136] ), .B(
        \D_cache/cache[5][136] ), .C(\D_cache/cache[6][136] ), .D(
        \D_cache/cache[7][136] ), .S0(n2090), .S1(n2173), .Y(\D_cache/n2070 )
         );
  DFFRX2 \i_MIPS/PC/PC_o_reg[31]  ( .D(\i_MIPS/PC/n65 ), .CK(clk), .RN(n4068), 
        .Q(ICACHE_addr[29]), .QN(\i_MIPS/PC/n33 ) );
  MXI2X2 \D_cache/U2118  ( .A(\D_cache/n2061 ), .B(\D_cache/n2062 ), .S0(n2147), .Y(\D_cache/N52 ) );
  MXI2X2 \D_cache/U2134  ( .A(\D_cache/n2093 ), .B(\D_cache/n2094 ), .S0(n4041), .Y(\D_cache/N36 ) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[30]  ( .D(\i_MIPS/PC/n64 ), .CK(clk), .RN(n4068), 
        .Q(ICACHE_addr[28]), .QN(\i_MIPS/PC/n32 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[1]  ( .D(\i_MIPS/N24 ), .CK(clk), .RN(n4047), .Q(
        \i_MIPS/IF_ID_1 ), .QN(\i_MIPS/n181 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[30]  ( .D(\i_MIPS/N53 ), .CK(clk), .RN(n4044), .Q(
        \i_MIPS/IF_ID_30 ), .QN(\i_MIPS/n210 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[54]  ( .D(\i_MIPS/n411 ), .CK(clk), .RN(n4050), .Q(
        n1889), .QN(\i_MIPS/n283 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[48]  ( .D(\i_MIPS/n423 ), .CK(clk), .RN(n4051), .Q(
        n1888), .QN(\i_MIPS/n295 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[42]  ( .D(\i_MIPS/n435 ), .CK(clk), .RN(n4052), .Q(
        n1887), .QN(\i_MIPS/n307 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[44]  ( .D(\i_MIPS/n431 ), .CK(clk), .RN(n4052), .Q(
        n1886), .QN(\i_MIPS/n303 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[43]  ( .D(\i_MIPS/n433 ), .CK(clk), .RN(n4052), .Q(
        n2717), .QN(\i_MIPS/n305 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[36]  ( .D(\i_MIPS/n438 ), .CK(clk), .RN(n4052), 
        .Q(n10297), .QN(n1847) );
  DFFRX1 \i_MIPS/PC/PC_o_reg[28]  ( .D(\i_MIPS/PC/n62 ), .CK(clk), .RN(n4068), 
        .Q(ICACHE_addr[26]), .QN(\i_MIPS/PC/n30 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[17]  ( .D(\i_MIPS/n457 ), .CK(clk), .RN(n4054), 
        .Q(n10316), .QN(n3037) );
  DFFRX1 \i_MIPS/EX_MEM_reg[23]  ( .D(\i_MIPS/n451 ), .CK(clk), .RN(n4053), 
        .Q(n10310), .QN(n1620) );
  DFFRX2 \i_MIPS/EX_MEM_reg[28]  ( .D(\i_MIPS/n446 ), .CK(clk), .RN(n4053), 
        .Q(n10305), .QN(n1619) );
  DFFRX2 \i_MIPS/EX_MEM_reg[31]  ( .D(\i_MIPS/n443 ), .CK(clk), .RN(n4053), 
        .Q(n10302), .QN(n1618) );
  DFFRX2 \i_MIPS/EX_MEM_reg[24]  ( .D(\i_MIPS/n450 ), .CK(clk), .RN(n4053), 
        .Q(n10309), .QN(n1617) );
  DFFRX2 \i_MIPS/EX_MEM_reg[35]  ( .D(\i_MIPS/n439 ), .CK(clk), .RN(n4052), 
        .Q(n10298), .QN(n1616) );
  DFFRX1 \i_MIPS/EX_MEM_reg[12]  ( .D(\i_MIPS/n462 ), .CK(clk), .RN(n4054), 
        .QN(n2703) );
  DFFRX1 \i_MIPS/EX_MEM_reg[20]  ( .D(\i_MIPS/n454 ), .CK(clk), .RN(n4054), 
        .Q(n10313), .QN(n1085) );
  DFFRX2 \i_MIPS/EX_MEM_reg[32]  ( .D(\i_MIPS/n442 ), .CK(clk), .RN(n4053), 
        .Q(n10301), .QN(n1084) );
  DFFRX2 \i_MIPS/ID_EX_reg[6]  ( .D(\i_MIPS/n472 ), .CK(clk), .RN(n4055), .Q(
        \i_MIPS/ALUOp[0] ), .QN(n1083) );
  DFFRX2 \i_MIPS/ID_EX_reg[78]  ( .D(\i_MIPS/n507 ), .CK(clk), .RN(n4058), .Q(
        \i_MIPS/ID_EX[78] ), .QN(n2885) );
  DFFRX1 \i_MIPS/ID_EX_reg[23]  ( .D(\i_MIPS/n548 ), .CK(clk), .RN(n4064), .Q(
        \i_MIPS/ALUin1[14] ), .QN(\i_MIPS/n357 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[27]  ( .D(\i_MIPS/n544 ), .CK(clk), .RN(n4064), .Q(
        \i_MIPS/ALUin1[18] ), .QN(\i_MIPS/n353 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[13]  ( .D(\i_MIPS/n558 ), .CK(clk), .RN(n4065), .Q(
        \i_MIPS/ALUin1[4] ), .QN(\i_MIPS/n367 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[34]  ( .D(\i_MIPS/n537 ), .CK(clk), .RN(n4063), .Q(
        \i_MIPS/ALUin1[25] ), .QN(\i_MIPS/n346 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[10]  ( .D(\i_MIPS/n561 ), .CK(clk), .RN(n4065), .Q(
        \i_MIPS/ALUin1[1] ), .QN(\i_MIPS/n370 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[53]  ( .D(\i_MIPS/N76 ), .CK(clk), .RN(n4061), .Q(
        \i_MIPS/IR_ID[21] ), .QN(\i_MIPS/n228 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[50]  ( .D(\i_MIPS/N73 ), .CK(clk), .RN(n4060), .Q(
        \i_MIPS/IR_ID[18] ), .QN(\i_MIPS/n316 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[15]  ( .D(\i_MIPS/n556 ), .CK(clk), .RN(n4065), .Q(
        \i_MIPS/ALUin1[6] ), .QN(\i_MIPS/n365 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[33]  ( .D(\i_MIPS/n441 ), .CK(clk), .RN(n4053), 
        .Q(n10300) );
  DFFRX1 \i_MIPS/IF_ID_reg[49]  ( .D(\i_MIPS/N72 ), .CK(clk), .RN(n4060), .Q(
        \i_MIPS/IR_ID[17] ), .QN(\i_MIPS/n314 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[25]  ( .D(\i_MIPS/n546 ), .CK(clk), .RN(n4064), .Q(
        \i_MIPS/ALUin1[16] ), .QN(\i_MIPS/n355 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[76]  ( .D(\i_MIPS/n509 ), .CK(clk), .RN(n4058), .Q(
        \i_MIPS/ID_EX[76] ), .QN(n2887) );
  DFFRX2 \i_MIPS/ID_EX_reg[26]  ( .D(\i_MIPS/n545 ), .CK(clk), .RN(n4064), .Q(
        \i_MIPS/ALUin1[17] ), .QN(\i_MIPS/n354 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[9]  ( .D(\i_MIPS/n562 ), .CK(clk), .RN(n4065), .Q(
        \i_MIPS/ALUin1[0] ), .QN(\i_MIPS/n371 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[14]  ( .D(\i_MIPS/n557 ), .CK(clk), .RN(n4065), .Q(
        \i_MIPS/ALUin1[5] ), .QN(\i_MIPS/n366 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[35]  ( .D(\i_MIPS/n536 ), .CK(clk), .RN(n4063), .Q(
        \i_MIPS/ALUin1[26] ), .QN(\i_MIPS/n345 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[12]  ( .D(\i_MIPS/n559 ), .CK(clk), .RN(n4065), .Q(
        \i_MIPS/ALUin1[3] ), .QN(\i_MIPS/n368 ) );
  MXI2X1 \D_cache/U2104  ( .A(\D_cache/n2033 ), .B(\D_cache/n2034 ), .S0(n3063), .Y(\D_cache/N66 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[39]  ( .D(\i_MIPS/n532 ), .CK(clk), .RN(n4063), .Q(
        \i_MIPS/ALUin1[30] ), .QN(\i_MIPS/n341 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[8]  ( .D(\i_MIPS/n466 ), .CK(clk), .RN(n4055), .Q(
        n10322), .QN(n2701) );
  DFFRX1 \i_MIPS/EX_MEM_reg[7]  ( .D(\i_MIPS/n467 ), .CK(clk), .RN(n4055), .Q(
        n10323), .QN(n2712) );
  DFFRX2 \i_MIPS/ID_EX_reg[77]  ( .D(\i_MIPS/n508 ), .CK(clk), .RN(n4058), .Q(
        \i_MIPS/ID_EX[77] ), .QN(n2888) );
  DFFRX1 \i_MIPS/ID_EX_reg[83]  ( .D(\i_MIPS/n502 ), .CK(clk), .RN(n4058), .Q(
        \i_MIPS/ID_EX[83] ), .QN(n2989) );
  DFFRX1 \i_MIPS/ID_EX_reg[85]  ( .D(\i_MIPS/n500 ), .CK(clk), .RN(n4058), .Q(
        \i_MIPS/ID_EX[85] ), .QN(n2992) );
  DFFRX1 \i_MIPS/ID_EX_reg[87]  ( .D(\i_MIPS/n498 ), .CK(clk), .RN(n4057), .Q(
        \i_MIPS/ID_EX[87] ), .QN(n2994) );
  DFFRX1 \i_MIPS/ID_EX_reg[111]  ( .D(\i_MIPS/n513 ), .CK(clk), .RN(n4060), 
        .Q(\i_MIPS/ID_EX[111] ), .QN(\i_MIPS/n313 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[112]  ( .D(\i_MIPS/n514 ), .CK(clk), .RN(n4060), 
        .Q(\i_MIPS/ID_EX[112] ), .QN(\i_MIPS/n315 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[3]  ( .D(\i_MIPS/n524 ), .CK(clk), .RN(n4062), .Q(
        DCACHE_ren), .QN(\i_MIPS/n334 ) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[15]  ( .D(\i_MIPS/PC/n49 ), .CK(clk), .RN(n4067), 
        .Q(ICACHE_addr[13]), .QN(\i_MIPS/PC/n17 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[66]  ( .D(\i_MIPS/N89 ), .CK(clk), .RN(n4044), .Q(
        \i_MIPS/IF_ID[66] ), .QN(\i_MIPS/n235 ) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[7]  ( .D(\i_MIPS/PC/n41 ), .CK(clk), .RN(n4066), 
        .Q(ICACHE_addr[5]), .QN(\i_MIPS/PC/n9 ) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[12]  ( .D(\i_MIPS/PC/n46 ), .CK(clk), .RN(n4067), 
        .Q(ICACHE_addr[10]), .QN(\i_MIPS/PC/n14 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[95]  ( .D(\i_MIPS/N118 ), .CK(clk), .RN(n4042), .Q(
        \i_MIPS/IF_ID[95] ), .QN(\i_MIPS/n177 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[85]  ( .D(\i_MIPS/N108 ), .CK(clk), .RN(n4043), .Q(
        \i_MIPS/IF_ID[85] ), .QN(\i_MIPS/n167 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[51]  ( .D(\i_MIPS/N74 ), .CK(clk), .RN(n4060), .Q(
        \i_MIPS/IR_ID[19] ), .QN(\i_MIPS/n318 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[54]  ( .D(\i_MIPS/N77 ), .CK(clk), .RN(n4061), .Q(
        \i_MIPS/IR_ID[22] ), .QN(\i_MIPS/n229 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[56]  ( .D(\i_MIPS/N79 ), .CK(clk), .RN(n4061), .Q(
        \i_MIPS/IR_ID[24] ), .QN(\i_MIPS/n231 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[41]  ( .D(\i_MIPS/n437 ), .CK(clk), .RN(n4052), .Q(
        n2799), .QN(\i_MIPS/n309 ) );
  MXI4X1 \D_cache/U2432  ( .A(\D_cache/cache[0][145] ), .B(
        \D_cache/cache[1][145] ), .C(\D_cache/cache[2][145] ), .D(
        \D_cache/cache[3][145] ), .S0(n2143), .S1(n2436), .Y(\D_cache/n2087 )
         );
  MXI4X1 \D_cache/U2429  ( .A(\D_cache/cache[4][144] ), .B(
        \D_cache/cache[5][144] ), .C(\D_cache/cache[6][144] ), .D(
        \D_cache/cache[7][144] ), .S0(n2142), .S1(n2410), .Y(\D_cache/n2086 )
         );
  MXI4X2 \D_cache/U2427  ( .A(\D_cache/cache[4][143] ), .B(
        \D_cache/cache[5][143] ), .C(\D_cache/cache[6][143] ), .D(
        \D_cache/cache[7][143] ), .S0(n2070), .S1(n2413), .Y(\D_cache/n2084 )
         );
  MXI2X2 \D_cache/U2128  ( .A(\D_cache/n2081 ), .B(\D_cache/n2082 ), .S0(n3066), .Y(\D_cache/N42 ) );
  MXI4X1 \D_cache/U2421  ( .A(\D_cache/cache[4][140] ), .B(
        \D_cache/cache[5][140] ), .C(\D_cache/cache[6][140] ), .D(
        \D_cache/cache[7][140] ), .S0(n2141), .S1(n2404), .Y(\D_cache/n2078 )
         );
  MXI2X2 \D_cache/U2124  ( .A(\D_cache/n2073 ), .B(\D_cache/n2074 ), .S0(n3066), .Y(\D_cache/N46 ) );
  MXI2X1 \D_cache/U2122  ( .A(\D_cache/n2069 ), .B(\D_cache/n2070 ), .S0(n3067), .Y(\D_cache/N48 ) );
  MXI2X1 \D_cache/U2121  ( .A(\D_cache/n2067 ), .B(\D_cache/n2068 ), .S0(
        DCACHE_addr[4]), .Y(\D_cache/N49 ) );
  MXI4X1 \D_cache/U2408  ( .A(\D_cache/cache[0][133] ), .B(
        \D_cache/cache[1][133] ), .C(\D_cache/cache[2][133] ), .D(
        \D_cache/cache[3][133] ), .S0(n2094), .S1(n2424), .Y(\D_cache/n2063 )
         );
  MXI4X1 \D_cache/U2407  ( .A(\D_cache/cache[4][133] ), .B(
        \D_cache/cache[5][133] ), .C(\D_cache/cache[6][133] ), .D(
        \D_cache/cache[7][133] ), .S0(n2104), .S1(n2422), .Y(\D_cache/n2064 )
         );
  MXI2X2 \D_cache/U2119  ( .A(\D_cache/n2063 ), .B(\D_cache/n2064 ), .S0(n3065), .Y(\D_cache/N51 ) );
  MXI4X2 \D_cache/U2401  ( .A(\D_cache/cache[4][130] ), .B(
        \D_cache/cache[5][130] ), .C(\D_cache/cache[6][130] ), .D(
        \D_cache/cache[7][130] ), .S0(n2131), .S1(n2428), .Y(\D_cache/n2058 )
         );
  MXI4X2 \D_cache/U2402  ( .A(\D_cache/cache[0][130] ), .B(
        \D_cache/cache[1][130] ), .C(\D_cache/cache[2][130] ), .D(
        \D_cache/cache[3][130] ), .S0(n2136), .S1(n2433), .Y(\D_cache/n2057 )
         );
  MXI2X2 \D_cache/U2116  ( .A(\D_cache/n2057 ), .B(\D_cache/n2058 ), .S0(
        n10321), .Y(\D_cache/N54 ) );
  DFFRX4 \i_MIPS/PC/PC_o_reg[2]  ( .D(\i_MIPS/PC/n36 ), .CK(clk), .RN(n4066), 
        .Q(ICACHE_addr[0]), .QN(\i_MIPS/PC/n4 ) );
  DFFRX4 \i_MIPS/PC/PC_o_reg[3]  ( .D(\i_MIPS/PC/n37 ), .CK(clk), .RN(n4066), 
        .Q(ICACHE_addr[1]), .QN(\i_MIPS/PC/n5 ) );
  DFFRX4 \i_MIPS/ID_EX_reg[74]  ( .D(\i_MIPS/n511 ), .CK(clk), .RN(n4058), .Q(
        \i_MIPS/ID_EX[74] ), .QN(n2886) );
  DFFRX4 \i_MIPS/ID_EX_reg[81]  ( .D(\i_MIPS/n504 ), .CK(clk), .RN(n4058), .Q(
        n55), .QN(n1082) );
  MXI4X1 \D_cache/U2397  ( .A(\D_cache/cache[4][128] ), .B(
        \D_cache/cache[5][128] ), .C(\D_cache/cache[6][128] ), .D(
        \D_cache/cache[7][128] ), .S0(n2144), .S1(n2425), .Y(\D_cache/n2054 )
         );
  MXI2X4 \D_cache/U2114  ( .A(\D_cache/n2053 ), .B(\D_cache/n2054 ), .S0(n3065), .Y(\D_cache/N56 ) );
  MXI2X4 \D_cache/U2117  ( .A(\D_cache/n2059 ), .B(\D_cache/n2060 ), .S0(n2146), .Y(\D_cache/N53 ) );
  MXI2X4 \D_cache/U2123  ( .A(\D_cache/n2071 ), .B(\D_cache/n2072 ), .S0(n4041), .Y(\D_cache/N47 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[57]  ( .D(\i_MIPS/n405 ), .CK(clk), .RN(n4050), .Q(
        \i_MIPS/ID_EX[57] ), .QN(\i_MIPS/n277 ) );
  DFFRX4 \i_MIPS/ID_EX_reg[11]  ( .D(\i_MIPS/n560 ), .CK(clk), .RN(n4065), .Q(
        \i_MIPS/ALUin1[2] ), .QN(\i_MIPS/n369 ) );
  MXI4X2 \D_cache/U2422  ( .A(\D_cache/cache[0][140] ), .B(
        \D_cache/cache[1][140] ), .C(\D_cache/cache[2][140] ), .D(
        \D_cache/cache[3][140] ), .S0(n2134), .S1(n2407), .Y(\D_cache/n2077 )
         );
  MXI2X2 \D_cache/U2126  ( .A(\D_cache/n2077 ), .B(\D_cache/n2078 ), .S0(
        DCACHE_addr[4]), .Y(\D_cache/N44 ) );
  MXI2X4 \D_cache/U2130  ( .A(\D_cache/n2085 ), .B(\D_cache/n2086 ), .S0(n2147), .Y(\D_cache/N40 ) );
  MXI2X4 \D_cache/U2131  ( .A(\D_cache/n2087 ), .B(\D_cache/n2088 ), .S0(
        DCACHE_addr[4]), .Y(\D_cache/N39 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[16]  ( .D(\i_MIPS/n555 ), .CK(clk), .RN(n4065), .Q(
        \i_MIPS/ALUin1[7] ), .QN(\i_MIPS/n364 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[89]  ( .D(\i_MIPS/n496 ), .CK(clk), .RN(n4057), .Q(
        \i_MIPS/ID_EX[89] ) );
  MXI4X2 \D_cache/U2411  ( .A(\D_cache/cache[4][135] ), .B(
        \D_cache/cache[5][135] ), .C(\D_cache/cache[6][135] ), .D(
        \D_cache/cache[7][135] ), .S0(n2063), .S1(n2178), .Y(\D_cache/n2068 )
         );
  MXI2X2 \D_cache/U2125  ( .A(\D_cache/n2075 ), .B(\D_cache/n2076 ), .S0(n2147), .Y(\D_cache/N45 ) );
  MXI2X2 \D_cache/U2115  ( .A(\D_cache/n2055 ), .B(\D_cache/n2056 ), .S0(
        n10321), .Y(\D_cache/N55 ) );
  DFFRX4 \i_MIPS/ID_EX_reg[75]  ( .D(\i_MIPS/n510 ), .CK(clk), .RN(n4058), .Q(
        \i_MIPS/ID_EX[75] ), .QN(n79) );
  DFFRX4 \i_MIPS/ID_EX_reg[24]  ( .D(\i_MIPS/n547 ), .CK(clk), .RN(n4064), .Q(
        \i_MIPS/ALUin1[15] ), .QN(\i_MIPS/n356 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[22]  ( .D(\i_MIPS/n549 ), .CK(clk), .RN(n4064), .Q(
        \i_MIPS/ALUin1[13] ), .QN(\i_MIPS/n358 ) );
  MXI2X2 \D_cache/U2136  ( .A(\D_cache/n2097 ), .B(\D_cache/n2098 ), .S0(n3063), .Y(\D_cache/N34 ) );
  DFFRX4 \i_MIPS/ID_EX_reg[7]  ( .D(\i_MIPS/n471 ), .CK(clk), .RN(n4055), .Q(
        \i_MIPS/ALUOp[1] ), .QN(n967) );
  MXI2X4 \D_cache/U2132  ( .A(\D_cache/n2089 ), .B(\D_cache/n2090 ), .S0(n2147), .Y(\D_cache/N38 ) );
  MXI4X2 \D_cache/U2446  ( .A(\D_cache/cache[0][152] ), .B(
        \D_cache/cache[1][152] ), .C(\D_cache/cache[2][152] ), .D(
        \D_cache/cache[3][152] ), .S0(n2071), .S1(n2438), .Y(\D_cache/n2101 )
         );
  NAND2X4 U2 ( .A(n8148), .B(n3577), .Y(n8190) );
  NAND3BX2 U3 ( .AN(n8220), .B(n8219), .C(n8218), .Y(\i_MIPS/PC/n46 ) );
  INVX4 U4 ( .A(\D_cache/N35 ), .Y(n2751) );
  CLKMX2X4 U5 ( .A(DCACHE_addr[7]), .B(DCACHE_rdata[9]), .S0(n4021), .Y(n3027)
         );
  AO21X4 U6 ( .A0(n5673), .A1(n6323), .B0(n5672), .Y(n6910) );
  OAI221X1 U7 ( .A0(n3107), .A1(n6911), .B0(n6912), .B1(n3098), .C0(n3096), 
        .Y(n6923) );
  BUFX6 U8 ( .A(n8308), .Y(n22) );
  NAND3BX2 U9 ( .AN(n7845), .B(n7844), .C(n7843), .Y(\i_MIPS/PC/n41 ) );
  OAI221X1 U10 ( .A0(n3106), .A1(n6324), .B0(n6325), .B1(n3098), .C0(n3096), 
        .Y(n6328) );
  INVX3 U11 ( .A(n8251), .Y(n6388) );
  INVX4 U12 ( .A(n5675), .Y(n4649) );
  NAND3X8 U13 ( .A(n6981), .B(n6980), .C(n6979), .Y(n7789) );
  NOR2X1 U14 ( .A(n2538), .B(n2539), .Y(n2537) );
  NAND2X2 U15 ( .A(n5484), .B(\i_MIPS/ID_EX[83] ), .Y(n6136) );
  NAND2X2 U16 ( .A(n4835), .B(n5483), .Y(n5904) );
  OAI31XL U17 ( .A0(n6920), .A1(\i_MIPS/ID_EX[83] ), .A2(n6919), .B0(n7014), 
        .Y(n6921) );
  NAND2X2 U18 ( .A(n6468), .B(n21), .Y(n6691) );
  CLKINVX4 U19 ( .A(n8225), .Y(n6747) );
  NOR2X1 U20 ( .A(n2600), .B(n2601), .Y(n2599) );
  INVXL U21 ( .A(n7073), .Y(n2) );
  INVX6 U22 ( .A(n7633), .Y(n7073) );
  NAND4X2 U23 ( .A(n4423), .B(n4422), .C(n4421), .D(n4420), .Y(n8690) );
  OA22X2 U24 ( .A0(n3458), .A1(n995), .B0(n3411), .B1(n107), .Y(n4421) );
  BUFX4 U25 ( .A(n2793), .Y(n3264) );
  BUFX4 U26 ( .A(n7048), .Y(n3164) );
  NAND4X1 U27 ( .A(n4743), .B(n4742), .C(n4741), .D(n4740), .Y(n7048) );
  INVX3 U28 ( .A(n2716), .Y(n4682) );
  NAND2BX4 U29 ( .AN(\i_MIPS/PC/n8 ), .B(n2902), .Y(n2800) );
  AND2X4 U30 ( .A(n10), .B(ICACHE_addr[2]), .Y(n2902) );
  AOI2BB2X1 U31 ( .B0(\D_cache/N150 ), .B1(n2153), .A0N(n23), .A1N(n8900), .Y(
        \D_cache/n177 ) );
  INVX1 U32 ( .A(n4680), .Y(n4677) );
  AOI222X1 U33 ( .A0(n2811), .A1(n6135), .B0(n6134), .B1(n6133), .C0(n6132), 
        .C1(n6131), .Y(n6143) );
  INVX3 U34 ( .A(n4774), .Y(\i_MIPS/EX_MEM_next[71] ) );
  NAND2X1 U35 ( .A(\i_MIPS/ALUin1[15] ), .B(n4646), .Y(n8477) );
  CLKMX2X8 U36 ( .A(\i_MIPS/n279 ), .B(n2889), .S0(n4018), .Y(n4646) );
  OA22X2 U37 ( .A0(n3309), .A1(n155), .B0(n3231), .B1(n1046), .Y(n4406) );
  AND3X2 U38 ( .A(\i_MIPS/ID_EX[76] ), .B(\i_MIPS/ALUOp[1] ), .C(n1083), .Y(
        n4608) );
  AND4X6 U39 ( .A(\i_MIPS/ALUOp[1] ), .B(n1083), .C(n2887), .D(n2888), .Y(
        n2893) );
  NAND3BX4 U40 ( .AN(n4388), .B(ICACHE_addr[4]), .C(n4387), .Y(n8114) );
  AND2X4 U41 ( .A(n1968), .B(n1969), .Y(n4479) );
  OAI222X1 U42 ( .A0(n6334), .A1(n5748), .B0(n3068), .B1(n5747), .C0(n5746), 
        .C1(n3069), .Y(n5753) );
  INVX2 U43 ( .A(n6022), .Y(n3) );
  INVX1 U44 ( .A(n6022), .Y(n4) );
  INVXL U45 ( .A(n6022), .Y(n8738) );
  CLKBUFX3 U46 ( .A(n8738), .Y(n3674) );
  OAI221X4 U47 ( .A0(n8766), .A1(n7044), .B0(n8753), .B1(n7043), .C0(n6021), 
        .Y(n6022) );
  CLKBUFX3 U48 ( .A(n6073), .Y(n5) );
  OAI221XL U49 ( .A0(n8759), .A1(n7044), .B0(n8746), .B1(n7043), .C0(n4771), 
        .Y(n4772) );
  NAND4X4 U50 ( .A(n4451), .B(n4450), .C(n4449), .D(n4448), .Y(n4463) );
  XNOR2X4 U51 ( .A(ICACHE_addr[11]), .B(n8694), .Y(n4451) );
  AOI2BB2X1 U52 ( .B0(\D_cache/N140 ), .B1(n2153), .A0N(n24), .A1N(n8890), .Y(
        \D_cache/n196 ) );
  BUFX8 U53 ( .A(n3039), .Y(n24) );
  INVX6 U54 ( .A(n4867), .Y(n8744) );
  NAND2BX2 U55 ( .AN(n3001), .B(n8591), .Y(n7407) );
  OAI221X4 U56 ( .A0(n3106), .A1(n5737), .B0(n5736), .B1(n3098), .C0(n3097), 
        .Y(n5741) );
  AO21X4 U57 ( .A0(n7896), .A1(n7895), .B0(n2857), .Y(n7913) );
  NAND4X6 U58 ( .A(n7330), .B(n7329), .C(n7328), .D(n7327), .Y(n8367) );
  NAND2BX2 U59 ( .AN(n2163), .B(n8653), .Y(n7330) );
  INVX3 U60 ( .A(n4727), .Y(n4725) );
  NAND2X1 U61 ( .A(\i_MIPS/ALUin1[1] ), .B(n4681), .Y(n6535) );
  MXI2X2 U62 ( .A(\i_MIPS/ID_EX[112] ), .B(\i_MIPS/ID_EX[85] ), .S0(
        \i_MIPS/ID_EX_5 ), .Y(n7632) );
  MXI2X4 U63 ( .A(DCACHE_addr[5]), .B(DCACHE_rdata[7]), .S0(n4023), .Y(n8740)
         );
  OAI221X4 U64 ( .A0(\D_cache/n164 ), .A1(n8863), .B0(n3074), .B1(n8844), .C0(
        \D_cache/n170 ), .Y(DCACHE_rdata[7]) );
  NAND2X1 U65 ( .A(n7998), .B(n3577), .Y(n8022) );
  INVX6 U66 ( .A(n2762), .Y(n3112) );
  BUFX4 U67 ( .A(n3112), .Y(n3109) );
  NAND2X6 U68 ( .A(n6974), .B(n6973), .Y(n6975) );
  XOR2X4 U69 ( .A(n2441), .B(n8228), .Y(n6974) );
  NAND2BX2 U70 ( .AN(n3576), .B(n8558), .Y(n7344) );
  NOR4X2 U71 ( .A(n5831), .B(n5830), .C(n6766), .D(n5829), .Y(n5836) );
  NAND2X1 U72 ( .A(n8535), .B(n8547), .Y(n5975) );
  NAND2X1 U73 ( .A(n4639), .B(\i_MIPS/n351 ), .Y(n8547) );
  NAND3X2 U74 ( .A(ICACHE_addr[14]), .B(ICACHE_addr[13]), .C(n7978), .Y(n7994)
         );
  INVX3 U75 ( .A(n7963), .Y(n7978) );
  NAND2X8 U76 ( .A(n3580), .B(n8146), .Y(n2001) );
  AND4X2 U77 ( .A(n7608), .B(n7632), .C(\i_MIPS/forward_unit/n32 ), .D(n4774), 
        .Y(\i_MIPS/forward_unit/n15 ) );
  OAI221X2 U78 ( .A0(\D_cache/n164 ), .A1(n8870), .B0(n3074), .B1(n8851), .C0(
        \D_cache/n199 ), .Y(DCACHE_rdata[0]) );
  OAI221X2 U79 ( .A0(\D_cache/n164 ), .A1(n8864), .B0(n3074), .B1(n8845), .C0(
        \D_cache/n171 ), .Y(DCACHE_rdata[6]) );
  OAI221X2 U80 ( .A0(\D_cache/n164 ), .A1(n8866), .B0(n3074), .B1(n8847), .C0(
        \D_cache/n173 ), .Y(DCACHE_rdata[4]) );
  OAI221X2 U81 ( .A0(\D_cache/n164 ), .A1(n8865), .B0(n3074), .B1(n8846), .C0(
        \D_cache/n172 ), .Y(DCACHE_rdata[5]) );
  OAI221X1 U82 ( .A0(\D_cache/n164 ), .A1(n8868), .B0(n3074), .B1(n8849), .C0(
        \D_cache/n177 ), .Y(DCACHE_rdata[2]) );
  BUFX8 U83 ( .A(\D_cache/n165 ), .Y(n3074) );
  INVX6 U84 ( .A(n8086), .Y(n8188) );
  OAI221X4 U85 ( .A0(n3106), .A1(n6536), .B0(n2821), .B1(n3098), .C0(n3096), 
        .Y(n6540) );
  NAND4X4 U86 ( .A(n7731), .B(n7730), .C(n7729), .D(n7728), .Y(n7898) );
  NAND2BX1 U87 ( .AN(n2163), .B(n8658), .Y(n7731) );
  NAND2X2 U88 ( .A(n6258), .B(n6390), .Y(n5536) );
  OA22XL U89 ( .A0(n6402), .A1(n6268), .B0(n3070), .B1(n6390), .Y(n6275) );
  OAI2BB1X1 U90 ( .A0N(n6392), .A1N(n6391), .B0(n6390), .Y(n6395) );
  AOI2BB1XL U91 ( .A0N(n5188), .A1N(n5187), .B0(n5186), .Y(n5189) );
  NAND2X4 U92 ( .A(n6127), .B(n6188), .Y(n5187) );
  OR2X8 U93 ( .A(n4597), .B(n6260), .Y(n4822) );
  NAND2X2 U94 ( .A(n8473), .B(n8480), .Y(n4597) );
  INVX1 U95 ( .A(n6879), .Y(n6) );
  CLKBUFX6 U96 ( .A(n8730), .Y(n3660) );
  NAND2X2 U97 ( .A(n7909), .B(n7908), .Y(n8207) );
  XOR3XL U98 ( .A(n7909), .B(n8209), .C(n7908), .Y(n7904) );
  NAND4X4 U99 ( .A(n7708), .B(n7707), .C(n7706), .D(n7705), .Y(n7908) );
  INVX3 U100 ( .A(n5190), .Y(n2759) );
  NAND3X4 U101 ( .A(n7386), .B(n7385), .C(n7383), .Y(n2714) );
  NAND2BX2 U102 ( .AN(n3001), .B(n8586), .Y(n7383) );
  BUFX4 U103 ( .A(n8512), .Y(n7) );
  NAND2XL U104 ( .A(\i_MIPS/ALUin1[9] ), .B(n11), .Y(n8512) );
  OAI221X4 U105 ( .A0(n7009), .A1(n6461), .B0(n6460), .B1(n6824), .C0(n6459), 
        .Y(n6481) );
  BUFX20 U106 ( .A(n2988), .Y(n8) );
  INVX6 U107 ( .A(ICACHE_addr[2]), .Y(n4388) );
  OAI221X4 U108 ( .A0(n3107), .A1(n6838), .B0(n6835), .B1(n3098), .C0(n3096), 
        .Y(n6852) );
  INVX2 U109 ( .A(n6839), .Y(n6835) );
  CLKBUFX3 U110 ( .A(n2766), .Y(n3351) );
  NAND3BX4 U111 ( .AN(n4603), .B(n5977), .C(n5976), .Y(n4601) );
  INVX8 U112 ( .A(n8300), .Y(n7072) );
  NAND2X4 U113 ( .A(n8470), .B(n8471), .Y(n6259) );
  AOI211X2 U114 ( .A0(n5130), .A1(n5401), .B0(n5129), .C0(n5128), .Y(n5131) );
  OAI2BB2X1 U115 ( .B0(n5127), .B1(n6610), .A0N(n5126), .A1N(n5125), .Y(n5128)
         );
  BUFX6 U116 ( .A(n4821), .Y(n9) );
  NAND2X2 U117 ( .A(n4653), .B(\i_MIPS/n358 ), .Y(n6404) );
  OAI221X4 U118 ( .A0(\i_MIPS/n359 ), .A1(n3092), .B0(\i_MIPS/n358 ), .B1(
        n3087), .C0(n4716), .Y(n6829) );
  OA22X2 U119 ( .A0(\i_MIPS/n349 ), .A1(n14), .B0(\i_MIPS/n350 ), .B1(n3078), 
        .Y(n5113) );
  OA22XL U120 ( .A0(n5900), .A1(n3082), .B0(\i_MIPS/n344 ), .B1(n3078), .Y(
        n4968) );
  OA22X2 U121 ( .A0(\i_MIPS/n344 ), .A1(n3082), .B0(\i_MIPS/n345 ), .B1(n3078), 
        .Y(n4895) );
  OA22XL U122 ( .A0(\i_MIPS/n351 ), .A1(n3082), .B0(\i_MIPS/n352 ), .B1(n3078), 
        .Y(n4986) );
  INVX6 U123 ( .A(n3079), .Y(n3078) );
  NAND2X2 U124 ( .A(n4646), .B(\i_MIPS/n356 ), .Y(n5549) );
  INVXL U125 ( .A(n2728), .Y(n5036) );
  CLKAND2X8 U126 ( .A(\i_MIPS/ALUin1[0] ), .B(n2728), .Y(n2892) );
  AND2X4 U127 ( .A(n2728), .B(\i_MIPS/n371 ), .Y(n2839) );
  NAND2X4 U128 ( .A(n2726), .B(n2727), .Y(n2728) );
  CLKBUFX6 U129 ( .A(n3022), .Y(n3017) );
  NAND3BX4 U130 ( .AN(\i_MIPS/ID_EX[75] ), .B(n2893), .C(n964), .Y(n4618) );
  CLKMX2X8 U131 ( .A(\i_MIPS/ID_EX[75] ), .B(n2717), .S0(n4020), .Y(n2716) );
  NAND4X1 U132 ( .A(\i_MIPS/ID_EX[75] ), .B(\i_MIPS/ID_EX[78] ), .C(
        \i_MIPS/ID_EX[73] ), .D(n2893), .Y(n4619) );
  MX2X2 U133 ( .A(n4609), .B(n2893), .S0(\i_MIPS/ID_EX[75] ), .Y(n4610) );
  BUFX20 U134 ( .A(ICACHE_addr[3]), .Y(n10) );
  AO21X4 U135 ( .A0(n5106), .A1(\i_MIPS/n370 ), .B0(n2839), .Y(n6534) );
  INVX3 U136 ( .A(n4681), .Y(n5106) );
  OAI222X1 U137 ( .A0(n3070), .A1(n5255), .B0(n5183), .B1(n6125), .C0(n5182), 
        .C1(n6201), .Y(n5210) );
  OAI211X2 U138 ( .A0(n4690), .A1(n5186), .B0(n5255), .C0(n6194), .Y(n4693) );
  NAND2X2 U139 ( .A(\i_MIPS/ALUin1[10] ), .B(n4688), .Y(n5255) );
  BUFX8 U140 ( .A(n4668), .Y(n11) );
  NAND4X4 U141 ( .A(\D_cache/n532 ), .B(\D_cache/n533 ), .C(\D_cache/n534 ), 
        .D(\D_cache/n535 ), .Y(\D_cache/n528 ) );
  CLKXOR2X2 U142 ( .A(\D_cache/N51 ), .B(n3037), .Y(\D_cache/n533 ) );
  NAND3BX2 U143 ( .AN(n10), .B(ICACHE_addr[2]), .C(\i_MIPS/PC/n8 ), .Y(n2793)
         );
  CLKBUFX3 U144 ( .A(n8457), .Y(n12) );
  CLKBUFX3 U145 ( .A(n8457), .Y(n13) );
  INVX6 U146 ( .A(n3073), .Y(n8457) );
  CLKBUFX6 U147 ( .A(n8457), .Y(n3615) );
  BUFX4 U148 ( .A(n3615), .Y(n3610) );
  BUFX8 U149 ( .A(n3615), .Y(n3611) );
  CLKBUFX8 U150 ( .A(n3612), .Y(n3614) );
  OAI221X4 U151 ( .A0(\D_cache/n164 ), .A1(n8855), .B0(n3074), .B1(n8836), 
        .C0(\D_cache/n193 ), .Y(DCACHE_rdata[15]) );
  BUFX8 U152 ( .A(n7840), .Y(n20) );
  AOI2BB1X2 U153 ( .A0N(n2758), .A1N(n4822), .B0(n9), .Y(n4823) );
  BUFX12 U154 ( .A(n3081), .Y(n14) );
  INVXL U155 ( .A(n2863), .Y(n3081) );
  XNOR2X4 U156 ( .A(n8275), .B(n8265), .Y(n6980) );
  CLKMX2X6 U157 ( .A(\i_MIPS/ID_EX[57] ), .B(\i_MIPS/ID_EX[89] ), .S0(n4018), 
        .Y(n52) );
  AOI22X1 U158 ( .A0(\D_cache/N126 ), .A1(n2153), .B0(n3032), .B1(
        \D_cache/N158 ), .Y(\D_cache/n181 ) );
  INVX8 U159 ( .A(n3040), .Y(n3032) );
  OAI222X4 U160 ( .A0(n2796), .A1(n6678), .B0(n6612), .B1(n5203), .C0(n6550), 
        .C1(n6338), .Y(n4918) );
  BUFX8 U161 ( .A(n8490), .Y(n15) );
  NAND2XL U162 ( .A(n2716), .B(n5381), .Y(n8490) );
  XNOR2X4 U163 ( .A(n8243), .B(n7782), .Y(n5449) );
  OAI222X4 U164 ( .A0(n5448), .A1(n3218), .B0(n5447), .B1(n3216), .C0(n2748), 
        .C1(n3215), .Y(n7782) );
  INVX3 U165 ( .A(n6503), .Y(n8743) );
  OAI222X4 U166 ( .A0(n6454), .A1(n3166), .B0(n6432), .B1(n2761), .C0(n8726), 
        .C1(n3162), .Y(n7923) );
  XNOR2X4 U167 ( .A(ICACHE_addr[7]), .B(n8690), .Y(n4429) );
  AOI221X2 U168 ( .A0(n5479), .A1(n5478), .B0(n5477), .B1(n5476), .C0(n6766), 
        .Y(n5486) );
  OAI221X4 U169 ( .A0(n3106), .A1(n6062), .B0(n5475), .B1(n3098), .C0(n3097), 
        .Y(n5476) );
  OA22X4 U170 ( .A0(n3461), .A1(n1003), .B0(n3413), .B1(n115), .Y(n4437) );
  OA22X2 U171 ( .A0(n3457), .A1(n1005), .B0(n3435), .B1(n117), .Y(n4414) );
  BUFX4 U172 ( .A(n3442), .Y(n3435) );
  OAI221X4 U173 ( .A0(n3106), .A1(n6691), .B0(n6469), .B1(n3098), .C0(n3096), 
        .Y(n6470) );
  INVX6 U174 ( .A(n6984), .Y(n3104) );
  CLKINVX4 U175 ( .A(n2869), .Y(n6984) );
  AND3X6 U176 ( .A(n8206), .B(n7946), .C(n2861), .Y(n7950) );
  NAND3X1 U177 ( .A(n7949), .B(n8206), .C(n7946), .Y(n7918) );
  NAND2X2 U178 ( .A(n7915), .B(n7914), .Y(n8206) );
  AOI221X2 U179 ( .A0(n4839), .A1(n4838), .B0(n4837), .B1(n4836), .C0(n6766), 
        .Y(n4843) );
  OAI221X4 U180 ( .A0(n3106), .A1(n4834), .B0(n2848), .B1(n3099), .C0(n3096), 
        .Y(n4836) );
  CLKBUFX20 U181 ( .A(n8131), .Y(n3000) );
  BUFX3 U182 ( .A(n2906), .Y(n3094) );
  BUFX2 U183 ( .A(n2906), .Y(n3093) );
  AND2XL U184 ( .A(n2906), .B(\i_MIPS/ALUin1[25] ), .Y(n2894) );
  AND2X1 U185 ( .A(n3075), .B(\i_MIPS/ID_EX[80] ), .Y(n2906) );
  BUFX20 U186 ( .A(n8133), .Y(n3001) );
  NAND3BX2 U187 ( .AN(n8426), .B(ICACHE_addr[0]), .C(\i_MIPS/PC/n5 ), .Y(n8133) );
  MX2X1 U188 ( .A(n5107), .B(n6993), .S0(n5106), .Y(n5108) );
  OAI221X4 U189 ( .A0(n2892), .A1(n3107), .B0(n2839), .B1(n3099), .C0(n3097), 
        .Y(n5107) );
  BUFX12 U190 ( .A(n2783), .Y(n16) );
  NAND2XL U191 ( .A(n2978), .B(n2974), .Y(n2783) );
  NAND2BX1 U192 ( .AN(n3576), .B(n8562), .Y(n7729) );
  CLKBUFX16 U193 ( .A(n8132), .Y(n3576) );
  CLKAND2X2 U194 ( .A(n7979), .B(n7981), .Y(n2806) );
  NAND2X6 U195 ( .A(n5385), .B(n5398), .Y(n4896) );
  XOR3XL U196 ( .A(n3580), .B(n7998), .C(n7997), .Y(n7990) );
  INVX6 U197 ( .A(n7997), .Y(n8000) );
  NAND2BX4 U198 ( .AN(n7987), .B(n8021), .Y(n7997) );
  AOI2BB1X2 U199 ( .A0N(n8065), .A1N(n8058), .B0(n8061), .Y(n8027) );
  INVX4 U200 ( .A(n8088), .Y(n8065) );
  XOR2X4 U201 ( .A(n8174), .B(n8180), .Y(n8175) );
  INVX8 U202 ( .A(n7994), .Y(n8016) );
  XNOR2X2 U203 ( .A(n8175), .B(n3577), .Y(n8178) );
  BUFX16 U204 ( .A(n3593), .Y(n17) );
  CLKBUFX16 U205 ( .A(n3593), .Y(n18) );
  INVX6 U206 ( .A(n8189), .Y(n8193) );
  AOI2BB1X1 U207 ( .A0N(n8147), .A1N(n8189), .B0(n8192), .Y(n8149) );
  NAND2X8 U208 ( .A(n8145), .B(n8144), .Y(n8189) );
  OAI2BB2X1 U209 ( .B0(\i_MIPS/n211 ), .B1(n3612), .A0N(n966), .A1N(n2161), 
        .Y(\i_MIPS/N54 ) );
  XNOR2X4 U210 ( .A(n8317), .B(ICACHE_addr[29]), .Y(n966) );
  INVX6 U211 ( .A(n8051), .Y(n8066) );
  INVX3 U212 ( .A(n8146), .Y(n8148) );
  NAND3X8 U213 ( .A(n1999), .B(n2000), .C(n8194), .Y(n8287) );
  OR2X2 U214 ( .A(n8197), .B(n3577), .Y(n1999) );
  AND2X4 U215 ( .A(n8277), .B(n12), .Y(n3046) );
  CLKINVX12 U216 ( .A(n20), .Y(n8277) );
  CLKAND2X6 U217 ( .A(n3579), .B(n8122), .Y(n2860) );
  XOR2X4 U218 ( .A(n1070), .B(\D_cache/N47 ), .Y(n3043) );
  XNOR2X4 U219 ( .A(\D_cache/N53 ), .B(DCACHE_addr[8]), .Y(n2769) );
  AOI2BB1X4 U220 ( .A0N(n8210), .A1N(n8209), .B0(n8208), .Y(n8212) );
  CLKINVX4 U221 ( .A(n7901), .Y(n8209) );
  OA22XL U222 ( .A0(n8181), .A1(n3599), .B0(n2158), .B1(n8180), .Y(n8182) );
  CLKINVX8 U223 ( .A(n8180), .Y(n8197) );
  BUFX6 U224 ( .A(n4830), .Y(n19) );
  OA22X2 U225 ( .A0(n8032), .A1(n3598), .B0(n2158), .B1(n8042), .Y(n8033) );
  INVX6 U226 ( .A(n8042), .Y(n8043) );
  OAI222X2 U227 ( .A0(n4965), .A1(n3219), .B0(n4964), .B1(n3216), .C0(n8734), 
        .C1(n3214), .Y(n7801) );
  INVX8 U228 ( .A(n8159), .Y(n4965) );
  INVX4 U229 ( .A(n6600), .Y(n8494) );
  NAND2X2 U230 ( .A(\i_MIPS/ALUin1[2] ), .B(n4682), .Y(n6600) );
  NAND2X2 U231 ( .A(n8320), .B(n8319), .Y(n8304) );
  AOI21X4 U232 ( .A0(n8291), .A1(n8270), .B0(n8269), .Y(n8272) );
  NAND2X2 U233 ( .A(n3579), .B(n8267), .Y(n8291) );
  XOR3X2 U234 ( .A(n3580), .B(n8126), .C(n8146), .Y(n8129) );
  OA21X2 U235 ( .A0(n2860), .A1(n8125), .B0(n8145), .Y(n8126) );
  OA22XL U236 ( .A0(n8138), .A1(n3599), .B0(n2158), .B1(n8146), .Y(n8139) );
  NAND2X4 U237 ( .A(n3579), .B(n8170), .Y(n8194) );
  OA22X4 U238 ( .A0(n8154), .A1(n3599), .B0(n2158), .B1(n8170), .Y(n8155) );
  INVX8 U239 ( .A(n8170), .Y(n8171) );
  XOR2X4 U240 ( .A(n8168), .B(ICACHE_addr[23]), .Y(n8170) );
  OAI222X2 U241 ( .A0(n5883), .A1(n3164), .B0(n5861), .B1(n2761), .C0(n8720), 
        .C1(n3163), .Y(n8295) );
  INVX6 U242 ( .A(n8284), .Y(n5883) );
  NAND3BX4 U243 ( .AN(n4922), .B(n4921), .C(n4920), .Y(n8159) );
  AOI222X1 U244 ( .A0(n2809), .A1(n6686), .B0(n4908), .B1(n4907), .C0(n4906), 
        .C1(n4905), .Y(n4921) );
  AOI222X2 U245 ( .A0(\i_MIPS/IF_ID[94] ), .A1(n2157), .B0(n8302), .B1(n8330), 
        .C0(\i_MIPS/IF_ID_29 ), .C1(n3596), .Y(n8297) );
  NAND2X4 U246 ( .A(n8302), .B(n3577), .Y(n8321) );
  INVX8 U247 ( .A(n8301), .Y(n8302) );
  OA22X4 U248 ( .A0(n8095), .A1(n3599), .B0(n2158), .B1(n8122), .Y(n8096) );
  XOR2X4 U249 ( .A(n8120), .B(ICACHE_addr[21]), .Y(n8122) );
  NAND3BX2 U250 ( .AN(ICACHE_addr[1]), .B(\i_MIPS/PC/n4 ), .C(n8684), .Y(n8132) );
  OAI222X4 U251 ( .A0(n5253), .A1(n3166), .B0(n5231), .B1(n2761), .C0(n8742), 
        .C1(n3162), .Y(n7887) );
  OAI211X2 U252 ( .A0(n4675), .A1(n4679), .B0(n4987), .C0(n4972), .Y(n4676) );
  INVX3 U253 ( .A(n4896), .Y(n4675) );
  INVX4 U254 ( .A(n8061), .Y(n8064) );
  AOI2BB1X2 U255 ( .A0N(\i_MIPS/ID_EX[74] ), .A1N(n2885), .B0(n4618), .Y(n4621) );
  NAND4X6 U256 ( .A(\i_MIPS/ID_EX[74] ), .B(n2893), .C(n79), .D(n2885), .Y(
        n5048) );
  MX2XL U257 ( .A(\i_MIPS/ID_EX[75] ), .B(n2885), .S0(\i_MIPS/ID_EX[74] ), .Y(
        n4615) );
  CLKMX2X6 U258 ( .A(n4612), .B(n4611), .S0(\i_MIPS/ID_EX[74] ), .Y(n4613) );
  OAI222X2 U259 ( .A0(n5533), .A1(n3164), .B0(n5511), .B1(n2761), .C0(n8739), 
        .C1(n3163), .Y(n8151) );
  INVX6 U260 ( .A(n8039), .Y(n5533) );
  CLKINVX8 U261 ( .A(n6748), .Y(n8226) );
  AOI222X2 U262 ( .A0(\i_MIPS/IF_ID[96] ), .A1(n2157), .B0(n8330), .B1(n966), 
        .C0(\i_MIPS/IF_ID_31 ), .C1(n3597), .Y(n8331) );
  NAND2BX2 U263 ( .AN(n8067), .B(n8082), .Y(n8412) );
  NAND2X4 U264 ( .A(n8083), .B(n8082), .Y(n8087) );
  NAND2X1 U265 ( .A(n8066), .B(n3577), .Y(n8082) );
  INVX4 U266 ( .A(n8352), .Y(n8359) );
  NAND4X4 U267 ( .A(n7346), .B(n7345), .C(n7344), .D(n7343), .Y(n8352) );
  XNOR2X4 U268 ( .A(n8256), .B(n7809), .Y(n5805) );
  OAI222X4 U269 ( .A0(n5731), .A1(n3218), .B0(n5730), .B1(n3217), .C0(n27), 
        .C1(n3215), .Y(n7809) );
  NAND3BX2 U270 ( .AN(n5336), .B(n5335), .C(n5334), .Y(n8229) );
  AOI222X2 U271 ( .A0(n2809), .A1(n6267), .B0(n5327), .B1(n5326), .C0(n5325), 
        .C1(n5324), .Y(n5335) );
  BUFX8 U272 ( .A(n6467), .Y(n21) );
  NAND2X8 U273 ( .A(\i_MIPS/PC_o[1] ), .B(n2160), .Y(n8238) );
  NAND2X8 U274 ( .A(\i_MIPS/BranchAddr[0] ), .B(n2159), .Y(n8261) );
  CLKINVX8 U275 ( .A(n8246), .Y(n5318) );
  NAND3BX4 U276 ( .AN(n5275), .B(n5274), .C(n5273), .Y(n8246) );
  MXI2X4 U277 ( .A(\i_MIPS/EX_MEM[5] ), .B(DCACHE_rdata[0]), .S0(n4022), .Y(
        n8727) );
  OAI221X4 U278 ( .A0(n3106), .A1(n6392), .B0(n6262), .B1(n3098), .C0(n3096), 
        .Y(n6265) );
  AO21X4 U279 ( .A0(n6324), .A1(n6339), .B0(n5539), .Y(n5540) );
  AOI21X1 U280 ( .A0(n6323), .A1(n8485), .B0(n5534), .Y(n2823) );
  NAND2X1 U281 ( .A(n4658), .B(\i_MIPS/n353 ), .Y(n5739) );
  NAND2XL U282 ( .A(\i_MIPS/ALUin1[18] ), .B(n4658), .Y(n4826) );
  INVX4 U283 ( .A(n4658), .Y(n4643) );
  MXI2X2 U284 ( .A(\i_MIPS/ID_EX[59] ), .B(\i_MIPS/ID_EX[91] ), .S0(n4018), 
        .Y(n4658) );
  OAI222X2 U285 ( .A0(n5318), .A1(n3164), .B0(n5296), .B1(n2761), .C0(n2795), 
        .C1(n3163), .Y(n7903) );
  MXI2X4 U286 ( .A(\i_MIPS/ID_EX[58] ), .B(\i_MIPS/ID_EX[90] ), .S0(n4018), 
        .Y(n4657) );
  INVX20 U287 ( .A(n4020), .Y(n4018) );
  XNOR2X1 U288 ( .A(n8071), .B(n3577), .Y(n8073) );
  XOR2X4 U289 ( .A(n8070), .B(n8075), .Y(n8071) );
  CLKXOR2X1 U290 ( .A(n7821), .B(n10), .Y(n8372) );
  INVX4 U291 ( .A(n7821), .Y(n7822) );
  NAND2X4 U292 ( .A(n7815), .B(ICACHE_addr[2]), .Y(n7821) );
  NAND2X8 U293 ( .A(ICACHE_addr[1]), .B(ICACHE_addr[0]), .Y(n7819) );
  NAND3BX4 U294 ( .AN(n8426), .B(ICACHE_addr[1]), .C(\i_MIPS/PC/n4 ), .Y(n8131) );
  XOR3X2 U295 ( .A(n3580), .B(n8268), .C(n8270), .Y(n8200) );
  NAND2X2 U296 ( .A(n8289), .B(n3002), .Y(n8270) );
  OAI2BB2X4 U297 ( .B0(\i_MIPS/n177 ), .B1(n13), .A0N(n2159), .A1N(n8307), .Y(
        \i_MIPS/N118 ) );
  AOI32X2 U298 ( .A0(n8321), .A1(n8320), .A2(n8319), .B0(n3579), .B1(n8318), 
        .Y(n8323) );
  OAI2BB2X1 U299 ( .B0(\i_MIPS/n207 ), .B1(n12), .A0N(n8268), .A1N(n2161), .Y(
        \i_MIPS/N50 ) );
  NAND2X4 U300 ( .A(n8268), .B(n3577), .Y(n8288) );
  CLKINVX6 U301 ( .A(n8267), .Y(n8268) );
  OAI2BB2X1 U302 ( .B0(\i_MIPS/n175 ), .B1(n3615), .A0N(n2159), .A1N(n8274), 
        .Y(\i_MIPS/N116 ) );
  CLKINVX3 U303 ( .A(n8276), .Y(n8274) );
  CLKINVX8 U304 ( .A(n8122), .Y(n8124) );
  INVX4 U305 ( .A(n8083), .Y(n8069) );
  NAND2X4 U306 ( .A(n8413), .B(n3577), .Y(n8083) );
  XOR2X4 U307 ( .A(n2802), .B(ICACHE_addr[26]), .Y(n8286) );
  NAND2X2 U308 ( .A(n8285), .B(ICACHE_addr[25]), .Y(n2802) );
  NAND2BX4 U309 ( .AN(n8149), .B(n8190), .Y(n8173) );
  OA22XL U310 ( .A0(n8076), .A1(n3599), .B0(n2158), .B1(n8075), .Y(n8077) );
  CLKINVX12 U311 ( .A(n8075), .Y(n8091) );
  XOR2X4 U312 ( .A(n8057), .B(ICACHE_addr[20]), .Y(n8075) );
  NAND2X1 U313 ( .A(n8293), .B(n3577), .Y(n8319) );
  INVX4 U314 ( .A(n8288), .Y(n8269) );
  NAND3X6 U315 ( .A(n8289), .B(n8288), .C(n3002), .Y(n8290) );
  CLKXOR2X2 U316 ( .A(n8068), .B(ICACHE_addr[19]), .Y(n8420) );
  NAND3X4 U317 ( .A(ICACHE_addr[18]), .B(ICACHE_addr[17]), .C(n8056), .Y(n8068) );
  INVX4 U318 ( .A(n8191), .Y(n8172) );
  OAI211X2 U319 ( .A0(n8193), .A1(n8192), .B0(n8191), .C0(n8190), .Y(n8195) );
  NAND2X2 U320 ( .A(n8171), .B(n3577), .Y(n8191) );
  NAND2X4 U321 ( .A(n8185), .B(ICACHE_addr[23]), .Y(n8169) );
  INVX3 U322 ( .A(n8168), .Y(n8185) );
  NAND3X6 U323 ( .A(ICACHE_addr[26]), .B(ICACHE_addr[25]), .C(n8285), .Y(n8305) );
  INVX4 U324 ( .A(n8271), .Y(n8285) );
  CLKXOR2X2 U325 ( .A(n8271), .B(ICACHE_addr[25]), .Y(n8267) );
  NAND3X4 U326 ( .A(ICACHE_addr[24]), .B(ICACHE_addr[23]), .C(n8185), .Y(n8271) );
  XOR2X4 U327 ( .A(n8169), .B(ICACHE_addr[24]), .Y(n8180) );
  NAND2X1 U328 ( .A(n8197), .B(n3577), .Y(n8289) );
  XOR2X2 U329 ( .A(n8315), .B(ICACHE_addr[28]), .Y(n8318) );
  NAND2BX2 U330 ( .AN(n8305), .B(ICACHE_addr[27]), .Y(n8315) );
  INVX4 U331 ( .A(n7977), .Y(n5803) );
  OAI2BB1X2 U332 ( .A0N(n8493), .A1N(n8492), .B0(n8491), .Y(n8496) );
  INVXL U333 ( .A(n15), .Y(n8493) );
  CLKINVX1 U334 ( .A(n8711), .Y(n1960) );
  INVX3 U335 ( .A(n4034), .Y(n3061) );
  CLKINVX6 U336 ( .A(n4032), .Y(n3059) );
  CLKINVX6 U337 ( .A(n4033), .Y(n3060) );
  CLKINVX4 U338 ( .A(n3061), .Y(n2372) );
  INVX1 U339 ( .A(n3056), .Y(n2122) );
  CLKINVX2 U340 ( .A(n3061), .Y(n2370) );
  CLKMX2X4 U341 ( .A(n5747), .B(n5748), .S0(n4016), .Y(n6685) );
  CLKINVX1 U342 ( .A(n6334), .Y(n5480) );
  CLKINVX1 U343 ( .A(n3069), .Y(n6337) );
  NAND4X4 U344 ( .A(\i_MIPS/IF_ID[97] ), .B(\i_MIPS/n233 ), .C(n7831), .D(
        n7830), .Y(n7080) );
  INVX3 U345 ( .A(n2149), .Y(n3062) );
  NAND2X2 U346 ( .A(n7822), .B(n2155), .Y(n7818) );
  NAND2X4 U347 ( .A(\i_MIPS/ALUin1[13] ), .B(n4651), .Y(n6400) );
  BUFX4 U348 ( .A(n4030), .Y(n4027) );
  INVX3 U349 ( .A(n8255), .Y(n5731) );
  CLKMX2X2 U350 ( .A(n1092), .B(\D_cache/n178 ), .S0(n4023), .Y(n5859) );
  INVX6 U351 ( .A(n8324), .Y(n3581) );
  INVX1 U352 ( .A(n8665), .Y(n7559) );
  INVX1 U353 ( .A(n8633), .Y(n7558) );
  AOI222X1 U354 ( .A0(n5757), .A1(n6619), .B0(n2826), .B1(n5756), .C0(n5755), 
        .C1(n6993), .Y(n5758) );
  XOR2X1 U355 ( .A(n7995), .B(ICACHE_addr[16]), .Y(n8025) );
  NAND4X1 U356 ( .A(n7236), .B(n7235), .C(n7234), .D(n7233), .Y(n7838) );
  INVX1 U357 ( .A(n8467), .Y(n8469) );
  INVXL U358 ( .A(n8498), .Y(n8505) );
  NAND2XL U359 ( .A(n8466), .B(n8473), .Y(n8514) );
  NAND2X6 U360 ( .A(n4525), .B(n4524), .Y(n4526) );
  NAND2X6 U361 ( .A(n1961), .B(n1962), .Y(n4524) );
  INVX1 U362 ( .A(n4625), .Y(n4703) );
  CLKINVX1 U363 ( .A(n8524), .Y(n6058) );
  INVX3 U364 ( .A(n4629), .Y(n4630) );
  INVX3 U365 ( .A(n8192), .Y(n8187) );
  AOI21X1 U366 ( .A0(n6688), .A1(n8548), .B0(n6687), .Y(n2853) );
  INVXL U367 ( .A(n8549), .Y(n6687) );
  INVX3 U368 ( .A(n4031), .Y(n3058) );
  INVX3 U369 ( .A(n4038), .Y(n4031) );
  XNOR2X2 U370 ( .A(n1617), .B(\D_cache/N44 ), .Y(\D_cache/n531 ) );
  XNOR2X2 U371 ( .A(n1620), .B(\D_cache/N45 ), .Y(\D_cache/n529 ) );
  INVXL U372 ( .A(n8507), .Y(n4969) );
  OR2X1 U373 ( .A(n6846), .B(n6845), .Y(n2744) );
  NAND4BX1 U374 ( .AN(n7039), .B(n7038), .C(n7037), .D(n7036), .Y(n7040) );
  NAND2X2 U375 ( .A(n4670), .B(\i_MIPS/n366 ), .Y(n5398) );
  NAND2X2 U376 ( .A(n4669), .B(\i_MIPS/n367 ), .Y(n5385) );
  NAND4BX2 U377 ( .AN(n6285), .B(n6284), .C(n6283), .D(n6282), .Y(n6296) );
  OR2X1 U378 ( .A(n3507), .B(n1033), .Y(n1959) );
  BUFX8 U379 ( .A(n3351), .Y(n3330) );
  BUFX12 U380 ( .A(n3397), .Y(n3373) );
  BUFX16 U381 ( .A(n3306), .Y(n3286) );
  CLKBUFX8 U382 ( .A(n3264), .Y(n3238) );
  CLKBUFX3 U383 ( .A(n2370), .Y(n2376) );
  BUFX4 U384 ( .A(n2395), .Y(n2413) );
  CLKBUFX3 U385 ( .A(n2311), .Y(n2320) );
  CLKBUFX3 U386 ( .A(n2370), .Y(n2377) );
  INVX3 U387 ( .A(n3056), .Y(n2123) );
  NAND2X2 U388 ( .A(n4681), .B(\i_MIPS/n370 ), .Y(n5124) );
  NAND4X1 U389 ( .A(n4535), .B(n4534), .C(n4533), .D(n4532), .Y(n4538) );
  OA22XL U390 ( .A0(n3480), .A1(n463), .B0(n3415), .B1(n1372), .Y(n4533) );
  BUFX4 U391 ( .A(n2395), .Y(n2412) );
  CLKBUFX2 U392 ( .A(n2371), .Y(n2380) );
  INVX3 U393 ( .A(n3056), .Y(n2134) );
  INVX1 U394 ( .A(n3056), .Y(n2113) );
  BUFX4 U395 ( .A(n2393), .Y(n2404) );
  BUFX4 U396 ( .A(n2393), .Y(n2403) );
  CLKBUFX3 U397 ( .A(n2332), .Y(n2343) );
  INVX2 U398 ( .A(n3056), .Y(n2131) );
  INVX2 U399 ( .A(n3056), .Y(n2136) );
  BUFX4 U400 ( .A(n2394), .Y(n2408) );
  BUFX4 U401 ( .A(n2394), .Y(n2407) );
  INVX3 U402 ( .A(n2059), .Y(n2116) );
  CLKBUFX3 U403 ( .A(n2313), .Y(n2328) );
  NAND2X4 U404 ( .A(n8091), .B(n3577), .Y(n8144) );
  CLKINVX1 U405 ( .A(n8569), .Y(n7556) );
  AO22X1 U406 ( .A0(n2853), .A1(n3100), .B0(n3110), .B1(n6692), .Y(n6697) );
  BUFX4 U407 ( .A(n5965), .Y(n3069) );
  OAI221X1 U408 ( .A0(n6334), .A1(n5462), .B0(n3076), .B1(n6464), .C0(n5614), 
        .Y(n6462) );
  BUFX12 U409 ( .A(\i_MIPS/ID_EX[82] ), .Y(n3076) );
  INVX3 U410 ( .A(n2145), .Y(n4661) );
  NAND2X2 U411 ( .A(\i_MIPS/ALUin1[17] ), .B(n4648), .Y(n5681) );
  BUFX8 U412 ( .A(n3261), .Y(n3237) );
  BUFX16 U413 ( .A(n3397), .Y(n3372) );
  BUFX8 U414 ( .A(n2766), .Y(n3331) );
  BUFX4 U415 ( .A(n3531), .Y(n3507) );
  BUFX6 U416 ( .A(n3574), .Y(n3548) );
  CLKBUFX3 U417 ( .A(n2313), .Y(n2326) );
  CLKBUFX3 U418 ( .A(n2310), .Y(n2314) );
  CLKBUFX3 U419 ( .A(n2333), .Y(n2346) );
  INVX1 U420 ( .A(n3056), .Y(n2125) );
  CLKBUFX3 U421 ( .A(n2310), .Y(n2315) );
  CLKBUFX3 U422 ( .A(n2350), .Y(n2356) );
  CLKBUFX3 U423 ( .A(n2350), .Y(n2357) );
  BUFX4 U424 ( .A(n2395), .Y(n2415) );
  CLKBUFX3 U425 ( .A(n2332), .Y(n2344) );
  BUFX4 U426 ( .A(n2393), .Y(n2401) );
  BUFX4 U427 ( .A(n2393), .Y(n2405) );
  BUFX4 U428 ( .A(n2394), .Y(n2406) );
  INVX2 U429 ( .A(n3056), .Y(n2135) );
  AOI221X1 U430 ( .A0(n5544), .A1(n5543), .B0(n5542), .B1(n5541), .C0(n6766), 
        .Y(n5555) );
  NAND3X2 U431 ( .A(ICACHE_addr[6]), .B(ICACHE_addr[5]), .C(n7846), .Y(n7861)
         );
  CLKMX2X2 U432 ( .A(n6798), .B(n6797), .S0(n4012), .Y(n6801) );
  MX2XL U433 ( .A(n5931), .B(n5930), .S0(n4013), .Y(n5934) );
  INVX3 U434 ( .A(n8242), .Y(n5448) );
  MX2X1 U435 ( .A(n5858), .B(n5857), .S0(n4013), .Y(n5861) );
  NAND3X2 U436 ( .A(ICACHE_addr[12]), .B(ICACHE_addr[11]), .C(n7943), .Y(n7963) );
  AO22X2 U437 ( .A0(n2850), .A1(n3101), .B0(n3108), .B1(n6395), .Y(n6397) );
  MX2XL U438 ( .A(n4763), .B(n4762), .S0(n4013), .Y(n4773) );
  NAND4BX1 U439 ( .AN(n4752), .B(n4751), .C(n4750), .D(n4749), .Y(n4763) );
  NAND4BX1 U440 ( .AN(n4761), .B(n4760), .C(n4759), .D(n4758), .Y(n4762) );
  INVX3 U441 ( .A(n8231), .Y(n6187) );
  NAND4BX1 U442 ( .AN(n4799), .B(n4798), .C(n4797), .D(n4796), .Y(n4800) );
  INVX4 U443 ( .A(n8314), .Y(n4810) );
  INVX1 U444 ( .A(\D_cache/N30 ), .Y(n8808) );
  CLKBUFX2 U445 ( .A(n2372), .Y(n2388) );
  CLKBUFX2 U446 ( .A(n2373), .Y(n2390) );
  CLKBUFX3 U447 ( .A(n2350), .Y(n2354) );
  CLKBUFX2 U448 ( .A(n2353), .Y(n2367) );
  CLKBUFX3 U449 ( .A(n2370), .Y(n2378) );
  CLKBUFX3 U450 ( .A(n2330), .Y(n2335) );
  CLKBUFX3 U451 ( .A(n2352), .Y(n2365) );
  INVX3 U452 ( .A(n2867), .Y(n3040) );
  CLKBUFX3 U453 ( .A(n2330), .Y(n2337) );
  BUFX16 U454 ( .A(n3039), .Y(n23) );
  INVX4 U455 ( .A(n2868), .Y(n7043) );
  INVX3 U456 ( .A(n3031), .Y(n8742) );
  MXI2X4 U457 ( .A(n2204), .B(DCACHE_rdata[5]), .S0(n4023), .Y(n2748) );
  NAND2X2 U458 ( .A(\i_MIPS/ALUin1[14] ), .B(n4645), .Y(n6335) );
  CLKMX2X2 U459 ( .A(n3072), .B(n2865), .S0(n6207), .Y(n6208) );
  OAI221X1 U460 ( .A0(n3106), .A1(n5260), .B0(n2849), .B1(n3098), .C0(n3097), 
        .Y(n5263) );
  INVX8 U461 ( .A(n6824), .Y(n6905) );
  NAND2XL U462 ( .A(n6337), .B(n6682), .Y(n5752) );
  CLKBUFX3 U463 ( .A(n2351), .Y(n2361) );
  OAI222X1 U464 ( .A0(n5731), .A1(n3164), .B0(n5709), .B1(n2761), .C0(n27), 
        .C1(n3163), .Y(n7989) );
  OR2X4 U465 ( .A(n5781), .B(n2761), .Y(n1949) );
  OR2X1 U466 ( .A(n8731), .B(n3163), .Y(n1950) );
  OR2X2 U467 ( .A(n5803), .B(n3164), .Y(n1948) );
  CLKMX2X2 U468 ( .A(n5954), .B(n5953), .S0(n4014), .Y(n5955) );
  CLKINVX1 U469 ( .A(n7797), .Y(n7798) );
  NOR3X1 U470 ( .A(n7796), .B(n7794), .C(n7795), .Y(n2830) );
  NAND4X4 U471 ( .A(n7414), .B(n7413), .C(n7412), .D(n7411), .Y(n8335) );
  XOR3XL U472 ( .A(n7863), .B(n7854), .C(n7862), .Y(n7857) );
  XOR3XL U473 ( .A(n7883), .B(n2827), .C(n7882), .Y(n7876) );
  NAND2BX1 U474 ( .AN(n2163), .B(n8661), .Y(n7607) );
  INVX4 U475 ( .A(n8367), .Y(n8373) );
  OAI21XL U476 ( .A0(\i_MIPS/n235 ), .A1(n3611), .B0(n8238), .Y(\i_MIPS/N89 )
         );
  NAND2X1 U477 ( .A(n8498), .B(n8507), .Y(n4592) );
  CLKINVX1 U478 ( .A(n8492), .Y(n8495) );
  NAND2X4 U479 ( .A(\i_MIPS/PC/n33 ), .B(n1981), .Y(n1983) );
  INVX3 U480 ( .A(n8712), .Y(n1981) );
  NAND2X2 U481 ( .A(ICACHE_addr[29]), .B(n8712), .Y(n1982) );
  XOR2X2 U482 ( .A(n8701), .B(ICACHE_addr[18]), .Y(n4402) );
  CLKINVX1 U483 ( .A(n8547), .Y(n8550) );
  NAND2X2 U484 ( .A(n4429), .B(n4428), .Y(n4430) );
  CLKINVX1 U485 ( .A(n5048), .Y(n4710) );
  AO21X2 U486 ( .A0(n5534), .A1(n8488), .B0(n8486), .Y(n5672) );
  INVX3 U487 ( .A(n6335), .Y(n5539) );
  OAI211X1 U488 ( .A0(n4665), .A1(n4655), .B0(n6913), .C0(n2825), .Y(n4656) );
  CLKINVX1 U489 ( .A(n5536), .Y(n4663) );
  NAND2X1 U490 ( .A(n4707), .B(\i_MIPS/n340 ), .Y(n8528) );
  NAND2BX1 U491 ( .AN(n4903), .B(n8498), .Y(n4970) );
  MXI2X4 U492 ( .A(\i_MIPS/ID_EX[47] ), .B(n3075), .S0(n4019), .Y(n4674) );
  CLKMX2X2 U493 ( .A(\i_MIPS/n301 ), .B(n2888), .S0(n4019), .Y(n4669) );
  OAI221XL U494 ( .A0(\i_MIPS/Register/register[2][12] ), .A1(n3124), .B0(
        \i_MIPS/Register/register[10][12] ), .B1(n3121), .C0(n6277), .Y(n6285)
         );
  AND2X2 U495 ( .A(\i_MIPS/IR_ID[17] ), .B(\i_MIPS/n312 ), .Y(n2978) );
  OAI22X1 U496 ( .A0(n8906), .A1(n8905), .B0(n8904), .B1(n8906), .Y(n8923) );
  OAI211X1 U497 ( .A0(n8489), .A1(n8513), .B0(n8488), .C0(n8487), .Y(n8906) );
  NAND2X2 U498 ( .A(\i_MIPS/n307 ), .B(n4020), .Y(n2731) );
  NAND2X1 U499 ( .A(n8217), .B(n8216), .Y(n7946) );
  NAND2X1 U500 ( .A(n2807), .B(n7913), .Y(n7949) );
  CLKINVX1 U501 ( .A(n52), .Y(n2154) );
  NAND2X2 U502 ( .A(n6391), .B(n6404), .Y(n5535) );
  CLKINVX1 U503 ( .A(n5187), .Y(n4690) );
  CLKINVX1 U504 ( .A(n11), .Y(n4689) );
  CLKINVX1 U505 ( .A(n8545), .Y(n5983) );
  CLKINVX1 U506 ( .A(n4635), .Y(n4627) );
  INVX1 U507 ( .A(n4642), .Y(n4639) );
  MXI2X4 U508 ( .A(\i_MIPS/ID_EX[49] ), .B(n55), .S0(n4019), .Y(n4667) );
  NAND2X1 U509 ( .A(n6466), .B(n8465), .Y(n6688) );
  NAND2X2 U510 ( .A(n6189), .B(n6207), .Y(n5186) );
  NAND2X1 U511 ( .A(n5470), .B(n5469), .Y(n6059) );
  CLKINVX1 U512 ( .A(n4628), .Y(n4626) );
  NAND2BX1 U513 ( .AN(n5195), .B(n7), .Y(n5259) );
  CLKBUFX3 U514 ( .A(n4692), .Y(n2145) );
  CLKINVX1 U515 ( .A(n6909), .Y(n5674) );
  CLKINVX1 U516 ( .A(n4657), .Y(n4648) );
  NAND2X4 U517 ( .A(n2892), .B(n5124), .Y(n6532) );
  NAND2X1 U518 ( .A(n4677), .B(\i_MIPS/n368 ), .Y(n8491) );
  NAND2X1 U519 ( .A(\i_MIPS/ALUin1[3] ), .B(n4680), .Y(n8492) );
  CLKINVX8 U520 ( .A(n2747), .Y(n4040) );
  NAND2X2 U521 ( .A(n2752), .B(n2753), .Y(\D_cache/n551 ) );
  NAND2X1 U522 ( .A(n8722), .B(\D_cache/N35 ), .Y(n2752) );
  XNOR2X1 U523 ( .A(n1618), .B(\D_cache/N37 ), .Y(\D_cache/n552 ) );
  XOR2X1 U524 ( .A(\D_cache/N32 ), .B(n10297), .Y(\D_cache/n539 ) );
  XNOR2X1 U525 ( .A(n1616), .B(\D_cache/N33 ), .Y(\D_cache/n537 ) );
  NAND2X1 U526 ( .A(\i_MIPS/ALUin1[28] ), .B(n4624), .Y(n5891) );
  CLKINVX1 U527 ( .A(n4624), .Y(n4704) );
  AND2X2 U528 ( .A(n3084), .B(\i_MIPS/ALUin1[14] ), .Y(n2987) );
  CLKINVX1 U529 ( .A(n5732), .Y(n5736) );
  NAND2X1 U530 ( .A(\i_MIPS/ALUin1[18] ), .B(n4643), .Y(n5738) );
  NAND2BX1 U531 ( .AN(n4899), .B(n5390), .Y(n4973) );
  AOI2BB1X1 U532 ( .A0N(n4898), .A1N(n4897), .B0(n4896), .Y(n4899) );
  NAND2X1 U533 ( .A(\i_MIPS/ALUin1[6] ), .B(n4674), .Y(n8507) );
  NOR2X1 U534 ( .A(n2718), .B(n6393), .Y(n2850) );
  AND2X2 U535 ( .A(n6394), .B(n8482), .Y(n2718) );
  NAND2X1 U536 ( .A(n4651), .B(\i_MIPS/n358 ), .Y(n8481) );
  AND4X1 U537 ( .A(n963), .B(n78), .C(\i_MIPS/forward_unit/n25 ), .D(n53), .Y(
        \i_MIPS/forward_unit/n10 ) );
  AND2X2 U538 ( .A(\i_MIPS/EX_MEM_0 ), .B(n3219), .Y(n4806) );
  CLKBUFX3 U539 ( .A(n2373), .Y(n2389) );
  CLKBUFX3 U540 ( .A(n2373), .Y(n2391) );
  CLKBUFX3 U541 ( .A(n2310), .Y(n2317) );
  CLKBUFX3 U542 ( .A(n2353), .Y(n2366) );
  CLKBUFX3 U543 ( .A(n2372), .Y(n2384) );
  CLKBUFX3 U544 ( .A(n2395), .Y(n2414) );
  CLKBUFX3 U545 ( .A(n2332), .Y(n2342) );
  AND3X2 U546 ( .A(n3099), .B(n3107), .C(n3097), .Y(n5045) );
  CLKBUFX3 U547 ( .A(n2393), .Y(n2402) );
  CLKBUFX3 U548 ( .A(n2396), .Y(n2418) );
  CLKBUFX3 U549 ( .A(n2396), .Y(n2419) );
  CLKBUFX3 U550 ( .A(n2397), .Y(n2424) );
  CLKBUFX3 U551 ( .A(n2398), .Y(n2427) );
  CLKBUFX3 U552 ( .A(n2395), .Y(n2411) );
  CLKBUFX3 U553 ( .A(n2397), .Y(n2423) );
  CLKBUFX3 U554 ( .A(n2397), .Y(n2422) );
  CLKINVX1 U555 ( .A(\D_cache/n316 ), .Y(n8903) );
  CLKBUFX3 U556 ( .A(n2399), .Y(n2433) );
  CLKBUFX3 U557 ( .A(n2400), .Y(n2437) );
  CLKBUFX3 U558 ( .A(n2399), .Y(n2435) );
  CLKBUFX3 U559 ( .A(n2399), .Y(n2431) );
  CLKINVX1 U560 ( .A(n3056), .Y(n2115) );
  CLKBUFX3 U561 ( .A(n2398), .Y(n2426) );
  CLKINVX1 U562 ( .A(n3056), .Y(n2133) );
  CLKBUFX3 U563 ( .A(n2353), .Y(n2368) );
  CLKBUFX3 U564 ( .A(n2311), .Y(n2318) );
  CLKINVX1 U565 ( .A(n3056), .Y(n2121) );
  INVX3 U566 ( .A(n7787), .Y(n7832) );
  NAND2X1 U567 ( .A(n2807), .B(n7912), .Y(n7954) );
  INVX1 U568 ( .A(n7871), .Y(n7869) );
  OR2X4 U569 ( .A(n8058), .B(n8063), .Y(n8090) );
  BUFX12 U570 ( .A(n8287), .Y(n3002) );
  NAND2X2 U571 ( .A(n2154), .B(\i_MIPS/n355 ), .Y(n6913) );
  NAND2X1 U572 ( .A(n52), .B(\i_MIPS/n355 ), .Y(n8539) );
  OAI221X1 U573 ( .A0(n5204), .A1(n6334), .B0(n3076), .B1(n6685), .C0(n5614), 
        .Y(n6678) );
  NAND2X2 U574 ( .A(n4689), .B(\i_MIPS/n362 ), .Y(n8468) );
  CLKINVX1 U575 ( .A(n8537), .Y(n4828) );
  NAND2X1 U576 ( .A(n3080), .B(\i_MIPS/ALUin1[13] ), .Y(n5457) );
  INVX3 U577 ( .A(n3094), .Y(n3092) );
  NAND2X1 U578 ( .A(n3080), .B(\i_MIPS/ALUin1[18] ), .Y(n5744) );
  OAI221XL U579 ( .A0(n5204), .A1(n3068), .B0(n3069), .B1(n5748), .C0(n5964), 
        .Y(n6050) );
  NAND2X2 U580 ( .A(n4648), .B(\i_MIPS/n354 ), .Y(n8540) );
  NAND2X1 U581 ( .A(\i_MIPS/ALUin1[17] ), .B(n4657), .Y(n8541) );
  CLKINVX1 U582 ( .A(n7819), .Y(n7815) );
  AND2X2 U583 ( .A(n3093), .B(\i_MIPS/ALUin1[5] ), .Y(n2984) );
  AND2X2 U584 ( .A(n3088), .B(\i_MIPS/ALUin1[4] ), .Y(n2898) );
  AND4X1 U585 ( .A(\i_MIPS/n323 ), .B(\i_MIPS/ALUOp[1] ), .C(
        \i_MIPS/ALU_Control/n11 ), .D(\i_MIPS/ID_EX[106] ), .Y(
        \i_MIPS/ALU_Control/n10 ) );
  OA22X2 U586 ( .A0(n3459), .A1(n996), .B0(n3412), .B1(n108), .Y(n4425) );
  OA22X2 U587 ( .A0(n3460), .A1(n1004), .B0(n3442), .B1(n116), .Y(n4433) );
  CLKBUFX3 U588 ( .A(n2400), .Y(n2438) );
  CLKBUFX3 U589 ( .A(n2310), .Y(n2316) );
  CLKBUFX3 U590 ( .A(n2398), .Y(n2428) );
  CLKINVX1 U591 ( .A(n2058), .Y(n2119) );
  CLKBUFX3 U592 ( .A(n2399), .Y(n2432) );
  CLKBUFX3 U593 ( .A(n2352), .Y(n2362) );
  CLKINVX1 U594 ( .A(n2060), .Y(n2120) );
  CLKBUFX3 U595 ( .A(n2396), .Y(n2416) );
  CLKBUFX3 U596 ( .A(n2399), .Y(n2434) );
  CLKINVX1 U597 ( .A(n3056), .Y(n2117) );
  CLKINVX1 U598 ( .A(n2057), .Y(n2118) );
  CLKBUFX3 U599 ( .A(n2394), .Y(n2409) );
  NOR4X1 U600 ( .A(n5097), .B(n5096), .C(n5095), .D(n5094), .Y(n5098) );
  OAI222X1 U601 ( .A0(n5448), .A1(n3166), .B0(n5426), .B1(n2761), .C0(n2748), 
        .C1(n3163), .Y(n8243) );
  NAND2X1 U602 ( .A(n2824), .B(n2832), .Y(n7010) );
  OAI222X1 U603 ( .A0(n4965), .A1(n3165), .B0(n4943), .B1(n2761), .C0(n8734), 
        .C1(n3162), .Y(n8160) );
  INVX8 U604 ( .A(n8426), .Y(n8684) );
  AND3X4 U605 ( .A(n1974), .B(n1975), .C(n7014), .Y(n6776) );
  NAND2X1 U606 ( .A(n6770), .B(n6769), .Y(n1974) );
  INVX3 U607 ( .A(n6982), .Y(n6987) );
  NAND2X1 U608 ( .A(n6988), .B(n7002), .Y(n7018) );
  OAI221X1 U609 ( .A0(n3106), .A1(n5604), .B0(n5603), .B1(n3098), .C0(n3097), 
        .Y(n5605) );
  AOI222X1 U610 ( .A0(n6680), .A1(n6773), .B0(n5618), .B1(n6993), .C0(n5617), 
        .C1(n6990), .Y(n5624) );
  CLKMX2X4 U611 ( .A(n6068), .B(n6067), .S0(n6066), .Y(n6069) );
  OAI31XL U612 ( .A0(n6849), .A1(n6848), .A2(n6847), .B0(n7014), .Y(n6850) );
  OAI221XL U613 ( .A0(n5888), .A1(n6754), .B0(n4721), .B1(n6996), .C0(n4720), 
        .Y(n4733) );
  CLKINVX1 U614 ( .A(n8459), .Y(n4607) );
  CLKINVX1 U615 ( .A(n8235), .Y(n5177) );
  CLKMX2X2 U616 ( .A(n7041), .B(n7040), .S0(n4012), .Y(n7047) );
  NAND4BX1 U617 ( .AN(n7030), .B(n7029), .C(n7028), .D(n7027), .Y(n7041) );
  CLKINVX1 U618 ( .A(n8040), .Y(n8056) );
  CLKINVX1 U619 ( .A(n7861), .Y(n7816) );
  CLKINVX1 U620 ( .A(n7892), .Y(n7916) );
  CLKINVX1 U621 ( .A(n8068), .Y(n8080) );
  CLKINVX1 U622 ( .A(n7928), .Y(n7943) );
  CLKINVX1 U623 ( .A(n7818), .Y(n7846) );
  CLKINVX1 U624 ( .A(n8120), .Y(n8142) );
  OAI222X1 U625 ( .A0(n6526), .A1(n3166), .B0(n6504), .B1(n2761), .C0(n8743), 
        .C1(n3162), .Y(n8163) );
  CLKINVX6 U626 ( .A(n8227), .Y(n6902) );
  OR2X1 U627 ( .A(n6319), .B(n3166), .Y(n1977) );
  NAND4X2 U628 ( .A(n4491), .B(n4490), .C(n4489), .D(n4488), .Y(n8709) );
  OA22X1 U629 ( .A0(n3286), .A1(n1012), .B0(n3238), .B1(n124), .Y(n4491) );
  OA22X1 U630 ( .A0(n3548), .A1(n125), .B0(n3507), .B1(n1014), .Y(n4488) );
  NAND4X2 U631 ( .A(n4487), .B(n4486), .C(n4485), .D(n4484), .Y(n8707) );
  OA22X1 U632 ( .A0(n3286), .A1(n1011), .B0(n3238), .B1(n123), .Y(n4487) );
  OA22X1 U633 ( .A0(n3373), .A1(n1075), .B0(n3330), .B1(n141), .Y(n4486) );
  AND2X2 U634 ( .A(n1958), .B(n1959), .Y(n4504) );
  AND2X2 U635 ( .A(n3979), .B(n3957), .Y(n2808) );
  OR2X1 U636 ( .A(n6902), .B(n3219), .Y(n1930) );
  INVX3 U637 ( .A(n3057), .Y(n2128) );
  OR2X2 U638 ( .A(n2757), .B(\D_cache/n204 ), .Y(n8807) );
  CLKBUFX3 U639 ( .A(n2312), .Y(n2325) );
  CLKBUFX3 U640 ( .A(n2373), .Y(n2392) );
  CLKBUFX3 U641 ( .A(n2371), .Y(n2379) );
  CLKBUFX3 U642 ( .A(n2333), .Y(n2347) );
  CLKBUFX3 U643 ( .A(n2372), .Y(n2386) );
  CLKBUFX3 U644 ( .A(n2370), .Y(n2374) );
  CLKBUFX3 U645 ( .A(n2312), .Y(n2323) );
  CLKBUFX3 U646 ( .A(n2372), .Y(n2387) );
  CLKBUFX3 U647 ( .A(n2331), .Y(n2340) );
  CLKBUFX3 U648 ( .A(n2312), .Y(n2324) );
  CLKBUFX3 U649 ( .A(n2371), .Y(n2383) );
  CLKBUFX3 U650 ( .A(n2350), .Y(n2355) );
  CLKBUFX3 U651 ( .A(n2352), .Y(n2363) );
  CLKBUFX3 U652 ( .A(n2371), .Y(n2382) );
  INVX3 U653 ( .A(n3057), .Y(n2129) );
  CLKMX2X2 U654 ( .A(DCACHE_rdata[13]), .B(n10315), .S0(\i_MIPS/n336 ), .Y(
        n3041) );
  OAI221X1 U655 ( .A0(\D_cache/n164 ), .A1(n8857), .B0(n3074), .B1(n8838), 
        .C0(\D_cache/n195 ), .Y(DCACHE_rdata[13]) );
  MXI2X2 U656 ( .A(DCACHE_addr[6]), .B(DCACHE_rdata[8]), .S0(n4021), .Y(n8745)
         );
  OAI221X1 U657 ( .A0(\D_cache/n164 ), .A1(n8862), .B0(n3074), .B1(n8843), 
        .C0(\D_cache/n169 ), .Y(DCACHE_rdata[8]) );
  MXI2X2 U658 ( .A(n10313), .B(DCACHE_rdata[15]), .S0(n4021), .Y(n8724) );
  CLKBUFX3 U659 ( .A(n2371), .Y(n2381) );
  CLKBUFX3 U660 ( .A(n2370), .Y(n2375) );
  CLKBUFX3 U661 ( .A(n2330), .Y(n2336) );
  CLKBUFX3 U662 ( .A(n2332), .Y(n2345) );
  CLKBUFX3 U663 ( .A(n2313), .Y(n2327) );
  CLKBUFX3 U664 ( .A(n2352), .Y(n2364) );
  NOR3BX2 U665 ( .AN(\i_MIPS/Register/n120 ), .B(\i_MIPS/Reg_W[3] ), .C(
        \i_MIPS/Reg_W[4] ), .Y(\i_MIPS/Register/n140 ) );
  CLKINVX1 U666 ( .A(n6097), .Y(n8737) );
  AOI2BB2X1 U667 ( .B0(\D_cache/N128 ), .B1(n2153), .A0N(n23), .A1N(n8878), 
        .Y(\D_cache/n183 ) );
  CLKBUFX3 U668 ( .A(n2313), .Y(n2329) );
  OAI221X1 U669 ( .A0(\D_cache/n164 ), .A1(n8856), .B0(n3074), .B1(n8837), 
        .C0(\D_cache/n194 ), .Y(DCACHE_rdata[14]) );
  AOI2BB2X1 U670 ( .B0(\D_cache/N152 ), .B1(n2153), .A0N(n24), .A1N(n8902), 
        .Y(\D_cache/n199 ) );
  NAND2BX1 U671 ( .AN(n3000), .B(n8618), .Y(n7385) );
  NAND2BX2 U672 ( .AN(n2163), .B(n8650), .Y(n7386) );
  NAND2BX1 U673 ( .AN(n3000), .B(n8619), .Y(n7413) );
  CLKINVX6 U674 ( .A(n7789), .Y(n7831) );
  INVX4 U675 ( .A(n7830), .Y(n7788) );
  CLKINVX1 U676 ( .A(n7305), .Y(n7306) );
  AND2X4 U677 ( .A(n8402), .B(\i_MIPS/PC/n4 ), .Y(n2840) );
  AND2X4 U678 ( .A(n8373), .B(n8372), .Y(n2855) );
  NAND2X1 U679 ( .A(n8368), .B(n8367), .Y(n8350) );
  AND2X2 U680 ( .A(n7849), .B(n7848), .Y(n2854) );
  AND2X2 U681 ( .A(n7881), .B(n7880), .Y(n2857) );
  AND2X2 U682 ( .A(n7931), .B(n7930), .Y(n2858) );
  AOI2BB1X1 U683 ( .A0N(n7984), .A1N(n8020), .B0(n8023), .Y(n7987) );
  NAND2BX1 U684 ( .AN(n8027), .B(n8059), .Y(n8045) );
  BUFX8 U685 ( .A(n3581), .Y(n3579) );
  NAND2X1 U686 ( .A(n8143), .B(n8144), .Y(n8123) );
  INVX1 U687 ( .A(n6141), .Y(n6906) );
  CLKMX2X2 U688 ( .A(n3072), .B(n2865), .S0(n6339), .Y(n6340) );
  AOI222X1 U689 ( .A0(n2810), .A1(n6686), .B0(n6329), .B1(n6328), .C0(n6327), 
        .C1(n6326), .Y(n6345) );
  CLKMX2X3 U690 ( .A(n6697), .B(n6696), .S0(n6695), .Y(n6698) );
  CLKINVX1 U691 ( .A(n5960), .Y(n5961) );
  CLKINVX1 U692 ( .A(n5888), .Y(n7006) );
  CLKINVX1 U693 ( .A(n6056), .Y(n5756) );
  AOI2BB2X1 U694 ( .B0(\D_cache/N143 ), .B1(n2153), .A0N(n3040), .A1N(n8893), 
        .Y(\D_cache/n166 ) );
  NAND4X1 U695 ( .A(\i_MIPS/Pred_1bit/current_state ), .B(n2830), .C(n7827), 
        .D(n2829), .Y(n7842) );
  OAI22XL U696 ( .A0(n3298), .A1(n456), .B0(n3251), .B1(n1365), .Y(n2781) );
  OA22X1 U697 ( .A0(n3295), .A1(n458), .B0(n3248), .B1(n1367), .Y(n7553) );
  OA22X1 U698 ( .A0(n3559), .A1(n459), .B0(n3517), .B1(n1368), .Y(n7550) );
  OA22X1 U699 ( .A0(n3382), .A1(n457), .B0(n3340), .B1(n1366), .Y(n7552) );
  NAND4X2 U700 ( .A(n4406), .B(n4405), .C(n4404), .D(n4403), .Y(n8689) );
  OA22X1 U701 ( .A0(n3575), .A1(n135), .B0(n3498), .B1(n1025), .Y(n4403) );
  OA22X1 U702 ( .A0(n3364), .A1(n136), .B0(n3321), .B1(n1026), .Y(n4405) );
  OA22X1 U703 ( .A0(n3575), .A1(n981), .B0(n3501), .B1(n93), .Y(n4420) );
  OA22X2 U704 ( .A0(n3279), .A1(n1006), .B0(n3230), .B1(n118), .Y(n4423) );
  OA22X2 U705 ( .A0(n3367), .A1(n982), .B0(n3324), .B1(n94), .Y(n4422) );
  NAND4X4 U706 ( .A(n4439), .B(n4438), .C(n4437), .D(n4436), .Y(n8693) );
  OA22X2 U707 ( .A0(n3544), .A1(n987), .B0(n3503), .B1(n99), .Y(n4436) );
  OA22X2 U708 ( .A0(n3282), .A1(n988), .B0(n3234), .B1(n100), .Y(n4439) );
  OA22X2 U709 ( .A0(n3369), .A1(n986), .B0(n3326), .B1(n98), .Y(n4438) );
  NAND4X2 U710 ( .A(n4467), .B(n4466), .C(n4465), .D(n4464), .Y(n8695) );
  NAND4X4 U711 ( .A(n4475), .B(n4474), .C(n4473), .D(n4472), .Y(n8696) );
  AND2X2 U712 ( .A(n1938), .B(n1939), .Y(n4468) );
  NAND4X4 U713 ( .A(n4447), .B(n4446), .C(n4445), .D(n4444), .Y(n8698) );
  OA22X2 U714 ( .A0(n3546), .A1(n977), .B0(n3505), .B1(n89), .Y(n4444) );
  NAND4X2 U715 ( .A(n4410), .B(n4409), .C(n4408), .D(n4407), .Y(n8703) );
  OA22X2 U716 ( .A0(n3277), .A1(n970), .B0(n3232), .B1(n81), .Y(n4410) );
  NAND4X4 U717 ( .A(n4416), .B(n4415), .C(n4414), .D(n4413), .Y(n8706) );
  OA22X1 U718 ( .A0(n3575), .A1(n993), .B0(n3500), .B1(n105), .Y(n4413) );
  OA22X1 U719 ( .A0(n3278), .A1(n994), .B0(n3232), .B1(n106), .Y(n4416) );
  OA22X1 U720 ( .A0(n3366), .A1(n992), .B0(n3323), .B1(n104), .Y(n4415) );
  NAND4X2 U721 ( .A(n4479), .B(n4478), .C(n4477), .D(n4476), .Y(n8708) );
  NAND4X4 U722 ( .A(n4523), .B(n4522), .C(n4521), .D(n4520), .Y(n8711) );
  OA22X1 U723 ( .A0(n3374), .A1(n126), .B0(n3331), .B1(n1015), .Y(n4522) );
  CLKINVX1 U724 ( .A(\D_cache/N88 ), .Y(n8851) );
  CLKINVX1 U725 ( .A(\D_cache/N87 ), .Y(n8850) );
  CLKINVX1 U726 ( .A(\D_cache/N84 ), .Y(n8847) );
  CLKINVX1 U727 ( .A(\D_cache/N83 ), .Y(n8846) );
  CLKINVX1 U728 ( .A(\D_cache/N82 ), .Y(n8845) );
  CLKINVX1 U729 ( .A(\D_cache/N120 ), .Y(n8870) );
  CLKINVX1 U730 ( .A(\D_cache/N119 ), .Y(n8869) );
  CLKINVX1 U731 ( .A(\D_cache/N116 ), .Y(n8866) );
  CLKINVX1 U732 ( .A(\D_cache/N115 ), .Y(n8865) );
  CLKINVX1 U733 ( .A(\D_cache/N114 ), .Y(n8864) );
  CLKINVX1 U734 ( .A(\D_cache/N112 ), .Y(n8862) );
  CLKINVX1 U735 ( .A(\D_cache/N111 ), .Y(n8861) );
  CLKINVX1 U736 ( .A(\D_cache/N110 ), .Y(n8860) );
  CLKINVX1 U737 ( .A(\D_cache/N106 ), .Y(n8856) );
  CLKINVX1 U738 ( .A(\D_cache/N104 ), .Y(n8854) );
  CLKINVX1 U739 ( .A(\D_cache/N103 ), .Y(n8853) );
  CLKINVX1 U740 ( .A(\D_cache/N97 ), .Y(n8767) );
  CLKBUFX3 U741 ( .A(n2330), .Y(n2334) );
  CLKBUFX3 U742 ( .A(n2311), .Y(n2319) );
  CLKBUFX3 U743 ( .A(n2331), .Y(n2339) );
  CLKBUFX3 U744 ( .A(n2311), .Y(n2321) );
  CLKBUFX3 U745 ( .A(n2333), .Y(n2348) );
  CLKBUFX3 U746 ( .A(n2351), .Y(n2359) );
  CLKBUFX3 U747 ( .A(n2331), .Y(n2338) );
  CLKINVX1 U748 ( .A(\D_cache/N184 ), .Y(n8902) );
  CLKINVX1 U749 ( .A(\D_cache/N183 ), .Y(n8901) );
  CLKINVX1 U750 ( .A(\D_cache/N181 ), .Y(n8899) );
  CLKINVX1 U751 ( .A(\D_cache/N180 ), .Y(n8898) );
  CLKINVX1 U752 ( .A(\D_cache/N179 ), .Y(n8897) );
  CLKINVX1 U753 ( .A(\D_cache/N178 ), .Y(n8896) );
  CLKINVX1 U754 ( .A(\D_cache/N177 ), .Y(n8895) );
  CLKINVX1 U755 ( .A(\D_cache/N176 ), .Y(n8894) );
  CLKINVX1 U756 ( .A(\D_cache/N175 ), .Y(n8893) );
  CLKINVX1 U757 ( .A(\D_cache/N174 ), .Y(n8892) );
  CLKINVX1 U758 ( .A(\D_cache/N170 ), .Y(n8888) );
  CLKINVX1 U759 ( .A(\D_cache/N168 ), .Y(n8886) );
  CLKINVX1 U760 ( .A(\D_cache/N165 ), .Y(n8883) );
  CLKINVX1 U761 ( .A(\D_cache/N164 ), .Y(n8882) );
  CLKINVX1 U762 ( .A(\D_cache/N163 ), .Y(n8881) );
  CLKINVX1 U763 ( .A(\D_cache/N161 ), .Y(n8879) );
  CLKINVX1 U764 ( .A(\D_cache/N160 ), .Y(n8878) );
  CLKINVX1 U765 ( .A(\D_cache/N159 ), .Y(n8877) );
  NAND4X1 U766 ( .A(n5555), .B(n5554), .C(n5553), .D(n5552), .Y(n8253) );
  NAND3BX2 U767 ( .AN(n4992), .B(n4991), .C(n4990), .Y(n8009) );
  NAND4X2 U768 ( .A(n6276), .B(n6275), .C(n6274), .D(n6273), .Y(n7786) );
  OR2X2 U769 ( .A(n8733), .B(n3214), .Y(n2740) );
  OR2X1 U770 ( .A(n3214), .B(n8736), .Y(n2711) );
  CLKINVX1 U771 ( .A(n8318), .Y(n8325) );
  BUFX12 U772 ( .A(n8415), .Y(n3593) );
  XOR2X2 U773 ( .A(n7836), .B(\i_MIPS/IF_ID[64] ), .Y(n7834) );
  NAND4X1 U774 ( .A(n6411), .B(n6410), .C(n6409), .D(n6408), .Y(n8249) );
  OAI222XL U775 ( .A0(n3070), .A1(n5390), .B0(n6461), .B1(n6402), .C0(n6407), 
        .C1(n5548), .Y(n5405) );
  OAI222XL U776 ( .A0(n6272), .A1(n5548), .B0(n3070), .B1(n5384), .C0(n6612), 
        .C1(n5320), .Y(n5336) );
  INVX3 U777 ( .A(n8229), .Y(n5379) );
  CLKMX2X2 U778 ( .A(n5251), .B(n5250), .S0(n4014), .Y(n5252) );
  OAI222X4 U779 ( .A0(n5318), .A1(n3219), .B0(n5317), .B1(n3216), .C0(n2795), 
        .C1(n3214), .Y(n7804) );
  INVX3 U780 ( .A(n8253), .Y(n5598) );
  CLKINVX4 U781 ( .A(n7814), .Y(n6971) );
  NAND3X2 U782 ( .A(n2754), .B(n2755), .C(n2756), .Y(n7810) );
  OR2X1 U783 ( .A(n8731), .B(n3215), .Y(n2756) );
  OR2X1 U784 ( .A(n6525), .B(n3216), .Y(n1944) );
  OR2X1 U785 ( .A(n6526), .B(n3219), .Y(n1943) );
  BUFX4 U786 ( .A(n7799), .Y(n2441) );
  NAND3X2 U787 ( .A(n1930), .B(n1931), .C(n1932), .Y(n7799) );
  OR2X1 U788 ( .A(n6880), .B(n3217), .Y(n1931) );
  OR2X1 U789 ( .A(n6), .B(n3214), .Y(n1932) );
  CLKMX2X2 U790 ( .A(n6821), .B(n6820), .S0(\i_MIPS/IR_ID[20] ), .Y(n6822) );
  CLKMX2X2 U791 ( .A(n5881), .B(n5880), .S0(n4014), .Y(n5882) );
  CLKMX2X2 U792 ( .A(n7068), .B(n7067), .S0(\i_MIPS/IR_ID[20] ), .Y(n7070) );
  NAND4BX1 U793 ( .AN(n7066), .B(n7065), .C(n7064), .D(n7063), .Y(n7067) );
  NAND4BX1 U794 ( .AN(n7057), .B(n7056), .C(n7055), .D(n7054), .Y(n7068) );
  CLKMX2X2 U795 ( .A(n4801), .B(n4800), .S0(n4015), .Y(n4809) );
  NAND4BX1 U796 ( .AN(n4790), .B(n4789), .C(n4788), .D(n4787), .Y(n4801) );
  CLKMX2X2 U797 ( .A(\i_MIPS/ID_EX[114] ), .B(\i_MIPS/ID_EX[87] ), .S0(
        \i_MIPS/ID_EX_5 ), .Y(n2890) );
  CLKMX2X2 U798 ( .A(\i_MIPS/ID_EX[115] ), .B(\i_MIPS/ID_EX[88] ), .S0(
        \i_MIPS/ID_EX_5 ), .Y(n2891) );
  INVX4 U799 ( .A(n3616), .Y(n3622) );
  NAND2X4 U800 ( .A(n1072), .B(n5134), .Y(n8235) );
  AND3X2 U801 ( .A(n5131), .B(n5132), .C(n5133), .Y(n1072) );
  CLKMX2X2 U802 ( .A(n5110), .B(n5109), .S0(\i_MIPS/ALUin1[1] ), .Y(n5134) );
  OA22X1 U803 ( .A0(n6202), .A1(n6996), .B0(n6136), .B1(n5680), .Y(n5132) );
  CLKMX2X2 U804 ( .A(n1847), .B(\D_cache/n175 ), .S0(n4021), .Y(n4771) );
  OAI221X1 U805 ( .A0(n8762), .A1(n7044), .B0(n8749), .B1(n7043), .C0(n5932), 
        .Y(n5933) );
  CLKMX2X2 U806 ( .A(n8722), .B(\D_cache/n179 ), .S0(n4021), .Y(n5932) );
  AOI2BB2X1 U807 ( .B0(\D_cache/N124 ), .B1(n2153), .A0N(n23), .A1N(n8874), 
        .Y(\D_cache/n179 ) );
  MXI2X1 U808 ( .A(n1091), .B(\D_cache/n185 ), .S0(n4022), .Y(n3024) );
  AOI2BB2X1 U809 ( .B0(\D_cache/N130 ), .B1(n2153), .A0N(n23), .A1N(n8880), 
        .Y(\D_cache/n185 ) );
  BUFX8 U810 ( .A(n8727), .Y(n3654) );
  AND4X1 U811 ( .A(\i_MIPS/IR_ID[31] ), .B(\i_MIPS/IR_ID[29] ), .C(n2995), .D(
        n7634), .Y(n2803) );
  CLKINVX1 U812 ( .A(n8216), .Y(n8221) );
  CLKINVX1 U813 ( .A(n7944), .Y(n7956) );
  CLKINVX1 U814 ( .A(n7965), .Y(n7968) );
  CLKINVX1 U815 ( .A(n7982), .Y(n7986) );
  CLKINVX1 U816 ( .A(n7996), .Y(n7998) );
  CLKINVX1 U817 ( .A(n8420), .Y(n8413) );
  BUFX16 U818 ( .A(n3046), .Y(n2160) );
  BUFX12 U819 ( .A(n3046), .Y(n2161) );
  BUFX16 U820 ( .A(n3046), .Y(n2159) );
  AOI2BB1X1 U821 ( .A0N(n6209), .A1N(n6824), .B0(n6208), .Y(n6210) );
  AOI222XL U822 ( .A0(n6830), .A1(n5960), .B0(n6774), .B1(n5898), .C0(n6832), 
        .C1(n5319), .Y(n4844) );
  OAI222XL U823 ( .A0(n3070), .A1(n6188), .B0(n6126), .B1(n6125), .C0(n2796), 
        .C1(n6124), .Y(n6144) );
  NAND3BX1 U824 ( .AN(n5210), .B(n5209), .C(n5208), .Y(n8012) );
  AOI222X1 U825 ( .A0(n2811), .A1(n5746), .B0(n5200), .B1(n5199), .C0(n5198), 
        .C1(n5197), .Y(n5209) );
  OAI222XL U826 ( .A0(n3070), .A1(n6258), .B0(n5610), .B1(n6125), .C0(n5612), 
        .C1(n5548), .Y(n5275) );
  NAND4X1 U827 ( .A(n5688), .B(n5687), .C(n5686), .D(n5685), .Y(n8255) );
  AOI222XL U828 ( .A0(n6680), .A1(n6206), .B0(n5733), .B1(n6993), .C0(n2818), 
        .C1(n6990), .Y(n5686) );
  AOI2BB1X1 U829 ( .A0N(n6824), .A1N(n5684), .B0(n5683), .Y(n5685) );
  BUFX12 U830 ( .A(n2724), .Y(n2157) );
  AND2X2 U831 ( .A(n3047), .B(n2862), .Y(n2724) );
  NAND4BX2 U832 ( .AN(n6626), .B(n6625), .C(n6624), .D(n6623), .Y(n8233) );
  NAND3X1 U833 ( .A(n1963), .B(n1964), .C(n6609), .Y(n6626) );
  OR4X4 U834 ( .A(n6554), .B(n2835), .C(n2836), .D(n2837), .Y(n8240) );
  NAND3BX1 U835 ( .AN(n8406), .B(n8405), .C(n8404), .Y(\i_MIPS/PC/n36 ) );
  OA22X2 U836 ( .A0(n8403), .A1(n3599), .B0(ICACHE_addr[0]), .B1(n2158), .Y(
        n8404) );
  AOI222X1 U837 ( .A0(\i_MIPS/IF_ID[93] ), .A1(n2157), .B0(n8293), .B1(n8330), 
        .C0(\i_MIPS/IF_ID_28 ), .C1(n3597), .Y(n8280) );
  OAI221XL U838 ( .A0(n8262), .A1(n18), .B0(\i_MIPS/PC/n2 ), .B1(n8457), .C0(
        n8260), .Y(\i_MIPS/PC/n34 ) );
  CLKINVX1 U839 ( .A(n8309), .Y(n8307) );
  NAND3BX2 U840 ( .AN(n8035), .B(n8034), .C(n8033), .Y(\i_MIPS/PC/n53 ) );
  NAND3BX2 U841 ( .AN(n7993), .B(n7992), .C(n7991), .Y(\i_MIPS/PC/n51 ) );
  NAND3BX2 U842 ( .AN(n8055), .B(n8054), .C(n8053), .Y(\i_MIPS/PC/n54 ) );
  NAND3BX2 U843 ( .AN(n7891), .B(n7890), .C(n7889), .Y(\i_MIPS/PC/n44 ) );
  NAND3BX2 U844 ( .AN(n7927), .B(n7926), .C(n7925), .Y(\i_MIPS/PC/n47 ) );
  NAND3BX2 U845 ( .AN(n7879), .B(n7878), .C(n7877), .Y(\i_MIPS/PC/n43 ) );
  NAND3X1 U846 ( .A(n2033), .B(n2034), .C(n2035), .Y(n8220) );
  NAND3BX2 U847 ( .AN(n8079), .B(n8078), .C(n8077), .Y(\i_MIPS/PC/n56 ) );
  AOI2BB2X1 U848 ( .B0(\i_MIPS/IF_ID[72] ), .B1(n2157), .A0N(n3594), .A1N(
        \i_MIPS/n187 ), .Y(n7844) );
  NAND3X1 U849 ( .A(n2039), .B(n2040), .C(n2041), .Y(n7845) );
  NAND3BX2 U850 ( .AN(n7907), .B(n7906), .C(n7905), .Y(\i_MIPS/PC/n45 ) );
  NAND3BX2 U851 ( .AN(n7942), .B(n7941), .C(n7940), .Y(\i_MIPS/PC/n48 ) );
  NAND3BX2 U852 ( .AN(n8205), .B(n8204), .C(n8203), .Y(\i_MIPS/PC/n61 ) );
  NAND3BX2 U853 ( .AN(n7860), .B(n7859), .C(n7858), .Y(\i_MIPS/PC/n42 ) );
  NAND3BX2 U854 ( .AN(n7975), .B(n7974), .C(n7973), .Y(\i_MIPS/PC/n50 ) );
  NAND3BX2 U855 ( .AN(n8008), .B(n8007), .C(n8006), .Y(\i_MIPS/PC/n52 ) );
  NAND3BX2 U856 ( .AN(n8141), .B(n8140), .C(n8139), .Y(\i_MIPS/PC/n58 ) );
  AND2X2 U857 ( .A(\i_MIPS/IF_ID[66] ), .B(n2157), .Y(n2719) );
  AO22X1 U858 ( .A0(n3612), .A1(n7075), .B0(\i_MIPS/ID_EX_5 ), .B1(n3629), .Y(
        \i_MIPS/n478 ) );
  NAND3BX1 U859 ( .AN(n7962), .B(n7961), .C(n7960), .Y(\i_MIPS/PC/n49 ) );
  NAND3X1 U860 ( .A(n2741), .B(n2742), .C(n2743), .Y(n7962) );
  NAND3BX2 U861 ( .AN(n8098), .B(n8097), .C(n8096), .Y(\i_MIPS/PC/n57 ) );
  NAND3BX2 U862 ( .AN(n8157), .B(n8156), .C(n8155), .Y(\i_MIPS/PC/n59 ) );
  OAI222XL U863 ( .A0(n3584), .A1(n195), .B0(n3645), .B1(n3582), .C0(n3689), 
        .C1(\i_MIPS/n207 ), .Y(n8777) );
  OAI222XL U864 ( .A0(n3585), .A1(n193), .B0(n3676), .B1(n3582), .C0(n3689), 
        .C1(\i_MIPS/n205 ), .Y(n8779) );
  OAI222XL U865 ( .A0(n3585), .A1(n194), .B0(n3636), .B1(n3582), .C0(n3689), 
        .C1(\i_MIPS/n199 ), .Y(n8785) );
  AO22X2 U866 ( .A0(n2904), .A1(n2829), .B0(\i_MIPS/IF_ID[97] ), .B1(n3073), 
        .Y(\i_MIPS/N120 ) );
  OAI2BB2XL U867 ( .B0(\i_MIPS/n212 ), .B1(n3613), .A0N(n2161), .A1N(n8402), 
        .Y(\i_MIPS/N55 ) );
  OAI2BB2XL U868 ( .B0(\i_MIPS/n214 ), .B1(n3611), .A0N(n2160), .A1N(n8381), 
        .Y(\i_MIPS/N57 ) );
  OAI2BB2XL U869 ( .B0(\i_MIPS/n176 ), .B1(n3612), .A0N(n2160), .A1N(n8294), 
        .Y(\i_MIPS/N117 ) );
  CLKINVX1 U870 ( .A(n8296), .Y(n8294) );
  OAI2BB2X1 U871 ( .B0(\i_MIPS/n178 ), .B1(n13), .A0N(n2159), .A1N(n8327), .Y(
        \i_MIPS/N119 ) );
  OAI2BB2XL U872 ( .B0(\i_MIPS/n165 ), .B1(n12), .A0N(n2160), .A1N(n8002), .Y(
        \i_MIPS/N106 ) );
  CLKINVX1 U873 ( .A(n8003), .Y(n8002) );
  OAI2BB2X1 U874 ( .B0(\i_MIPS/n169 ), .B1(n8457), .A0N(n2161), .A1N(n8072), 
        .Y(\i_MIPS/N110 ) );
  OAI2BB2XL U875 ( .B0(\i_MIPS/n171 ), .B1(n3613), .A0N(n2161), .A1N(n8127), 
        .Y(\i_MIPS/N112 ) );
  CLKINVX1 U876 ( .A(n8129), .Y(n8127) );
  OAI2BB2XL U877 ( .B0(\i_MIPS/n172 ), .B1(n3614), .A0N(n2159), .A1N(n8150), 
        .Y(\i_MIPS/N113 ) );
  CLKINVX1 U878 ( .A(n8152), .Y(n8150) );
  OAI2BB2XL U879 ( .B0(\i_MIPS/n173 ), .B1(n13), .A0N(n2161), .A1N(n8176), .Y(
        \i_MIPS/N114 ) );
  CLKINVX1 U880 ( .A(n8178), .Y(n8176) );
  NAND3BX2 U881 ( .AN(n8425), .B(n8424), .C(n8423), .Y(\i_MIPS/PC/n55 ) );
  NAND3BX2 U882 ( .AN(n8376), .B(n8375), .C(n8374), .Y(\i_MIPS/PC/n39 ) );
  NAND3BX2 U883 ( .AN(n8391), .B(n8390), .C(n8389), .Y(\i_MIPS/PC/n38 ) );
  NAND3BX1 U884 ( .AN(n8344), .B(n8343), .C(n8342), .Y(\i_MIPS/PC/n37 ) );
  NAND3X1 U885 ( .A(n1990), .B(n1991), .C(n1992), .Y(n8344) );
  NOR2X6 U886 ( .A(n6122), .B(n6121), .Y(n6978) );
  INVX4 U887 ( .A(n4650), .Y(n4664) );
  XNOR2X4 U888 ( .A(n8236), .B(n7733), .Y(n5178) );
  CLKINVX4 U889 ( .A(n8223), .Y(n4890) );
  AOI22X1 U890 ( .A0(\D_cache/N125 ), .A1(n2153), .B0(n3032), .B1(
        \D_cache/N157 ), .Y(\D_cache/n180 ) );
  MXI2X2 U891 ( .A(n10323), .B(DCACHE_rdata[2]), .S0(n4021), .Y(n8733) );
  CLKBUFX6 U892 ( .A(n8733), .Y(n3663) );
  INVX16 U893 ( .A(n4024), .Y(n3056) );
  OA22XL U894 ( .A0(\i_MIPS/ALUin1[8] ), .A1(n3082), .B0(\i_MIPS/ALUin1[7] ), 
        .B1(n3078), .Y(n4981) );
  NAND2X2 U895 ( .A(\i_MIPS/ALUin1[7] ), .B(n4686), .Y(n6127) );
  CLKMX2X4 U896 ( .A(\i_MIPS/n299 ), .B(n2885), .S0(n4019), .Y(n4670) );
  CLKINVX8 U897 ( .A(n8164), .Y(n6045) );
  AO22XL U898 ( .A0(n6469), .A1(n3101), .B0(n3108), .B1(n6691), .Y(n6473) );
  MXI2X4 U899 ( .A(DCACHE_addr[14]), .B(DCACHE_rdata[16]), .S0(n4023), .Y(
        n8728) );
  OAI221X4 U900 ( .A0(\D_cache/n164 ), .A1(n8854), .B0(n3074), .B1(n8835), 
        .C0(\D_cache/n192 ), .Y(DCACHE_rdata[16]) );
  BUFX4 U901 ( .A(n8313), .Y(n25) );
  INVX3 U902 ( .A(n5510), .Y(n8739) );
  CLKBUFX6 U903 ( .A(n8721), .Y(n3643) );
  INVX3 U904 ( .A(n5648), .Y(n8717) );
  INVX3 U905 ( .A(n8015), .Y(n5671) );
  NAND2X6 U906 ( .A(n6618), .B(\i_MIPS/ALU/N303 ), .Y(n7014) );
  CLKINVX1 U907 ( .A(n3061), .Y(n2373) );
  INVX3 U908 ( .A(n2722), .Y(n3063) );
  NAND2X1 U909 ( .A(n26), .B(n10), .Y(n2156) );
  BUFX4 U910 ( .A(n3306), .Y(n3285) );
  CLKINVX1 U911 ( .A(n3059), .Y(n2351) );
  CLKBUFX3 U912 ( .A(n2312), .Y(n2322) );
  CLKBUFX3 U913 ( .A(n3257), .Y(n3244) );
  CLKBUFX3 U914 ( .A(n2766), .Y(n3329) );
  BUFX4 U915 ( .A(n3487), .Y(n3463) );
  CLKINVX1 U916 ( .A(n3058), .Y(n2310) );
  CLKBUFX3 U917 ( .A(n2351), .Y(n2360) );
  INVX3 U918 ( .A(n2722), .Y(n3067) );
  INVX1 U919 ( .A(n4028), .Y(n2105) );
  NAND2X2 U920 ( .A(n2902), .B(\i_MIPS/PC/n8 ), .Y(n2766) );
  BUFX4 U921 ( .A(n3486), .Y(n3462) );
  CLKBUFX3 U922 ( .A(n3442), .Y(n3434) );
  CLKINVX1 U923 ( .A(n3058), .Y(n2311) );
  CLKBUFX3 U924 ( .A(n2351), .Y(n2358) );
  BUFX4 U925 ( .A(n3574), .Y(n3549) );
  BUFX4 U926 ( .A(n8114), .Y(n3440) );
  BUFX2 U927 ( .A(n2793), .Y(n3263) );
  CLKBUFX3 U928 ( .A(n3264), .Y(n3256) );
  INVX3 U929 ( .A(n3058), .Y(n2312) );
  CLKBUFX3 U930 ( .A(n2394), .Y(n2410) );
  INVX3 U931 ( .A(n2151), .Y(n3064) );
  BUFX4 U932 ( .A(n3308), .Y(n3306) );
  CLKINVX1 U933 ( .A(n3058), .Y(n2313) );
  CLKINVX1 U934 ( .A(n10321), .Y(n2150) );
  INVX1 U935 ( .A(n3056), .Y(n2112) );
  CLKBUFX3 U936 ( .A(n2767), .Y(n3573) );
  CLKBUFX3 U937 ( .A(n3573), .Y(n3571) );
  CLKINVX1 U938 ( .A(n3060), .Y(n2330) );
  INVX3 U939 ( .A(n2722), .Y(n3065) );
  INVX3 U940 ( .A(n2150), .Y(n3066) );
  CLKINVX1 U941 ( .A(n3056), .Y(n2124) );
  AND2X4 U942 ( .A(\i_MIPS/PC/n6 ), .B(\i_MIPS/PC/n8 ), .Y(n26) );
  CLKINVX1 U943 ( .A(n3060), .Y(n2332) );
  CLKBUFX3 U944 ( .A(n3482), .Y(n3469) );
  NAND3BXL U945 ( .AN(n8684), .B(n8553), .C(n3051), .Y(n8410) );
  INVX1 U946 ( .A(n4027), .Y(n2097) );
  NAND3X2 U947 ( .A(\i_MIPS/PC/n6 ), .B(ICACHE_addr[4]), .C(n4387), .Y(n2798)
         );
  CLKINVX1 U948 ( .A(n3060), .Y(n2333) );
  CLKBUFX3 U949 ( .A(n3526), .Y(n3513) );
  BUFX4 U950 ( .A(n8114), .Y(n3441) );
  CLKINVX1 U951 ( .A(n3059), .Y(n2353) );
  INVX1 U952 ( .A(n3056), .Y(n2114) );
  CLKINVX1 U953 ( .A(n3060), .Y(n2331) );
  CLKBUFX3 U954 ( .A(n2353), .Y(n2369) );
  AND2X2 U955 ( .A(n2980), .B(n2973), .Y(n187) );
  AND2X2 U956 ( .A(n2979), .B(n2870), .Y(n2775) );
  AND2X2 U957 ( .A(n2981), .B(n2871), .Y(n2774) );
  INVX3 U958 ( .A(n3080), .Y(n3077) );
  INVX4 U959 ( .A(n2869), .Y(n3098) );
  INVX3 U960 ( .A(n2869), .Y(n3099) );
  INVX3 U961 ( .A(n2722), .Y(n2147) );
  INVX3 U962 ( .A(n2722), .Y(n2146) );
  INVX16 U963 ( .A(n2722), .Y(DCACHE_addr[4]) );
  CLKINVX1 U964 ( .A(n3056), .Y(n2132) );
  MXI2X4 U965 ( .A(DCACHE_addr[15]), .B(DCACHE_rdata[17]), .S0(n4021), .Y(n27)
         );
  CLKBUFX3 U966 ( .A(n3397), .Y(n3391) );
  NAND2X1 U967 ( .A(\i_MIPS/Register/n122 ), .B(\i_MIPS/Register/n105 ), .Y(
        n28) );
  NAND2X1 U968 ( .A(\i_MIPS/Register/n122 ), .B(\i_MIPS/Register/n107 ), .Y(
        n29) );
  NAND2X1 U969 ( .A(\i_MIPS/Register/n122 ), .B(\i_MIPS/Register/n109 ), .Y(
        n30) );
  NAND2X1 U970 ( .A(\i_MIPS/Register/n122 ), .B(\i_MIPS/Register/n111 ), .Y(
        n31) );
  NAND2X1 U971 ( .A(\i_MIPS/Register/n122 ), .B(\i_MIPS/Register/n113 ), .Y(
        n32) );
  NAND2X1 U972 ( .A(\i_MIPS/Register/n122 ), .B(\i_MIPS/Register/n115 ), .Y(
        n33) );
  NAND2X1 U973 ( .A(\i_MIPS/Register/n122 ), .B(\i_MIPS/Register/n117 ), .Y(
        n34) );
  NAND2X1 U974 ( .A(\i_MIPS/Register/n122 ), .B(\i_MIPS/Register/n119 ), .Y(
        n35) );
  NAND2X1 U975 ( .A(\i_MIPS/Register/n131 ), .B(\i_MIPS/Register/n105 ), .Y(
        n36) );
  NAND2X1 U976 ( .A(\i_MIPS/Register/n131 ), .B(\i_MIPS/Register/n107 ), .Y(
        n37) );
  NAND2X1 U977 ( .A(\i_MIPS/Register/n131 ), .B(\i_MIPS/Register/n109 ), .Y(
        n38) );
  NAND2X1 U978 ( .A(\i_MIPS/Register/n131 ), .B(\i_MIPS/Register/n111 ), .Y(
        n39) );
  NAND2X1 U979 ( .A(\i_MIPS/Register/n131 ), .B(\i_MIPS/Register/n113 ), .Y(
        n40) );
  NAND2X1 U980 ( .A(\i_MIPS/Register/n131 ), .B(\i_MIPS/Register/n115 ), .Y(
        n41) );
  NAND2X1 U981 ( .A(\i_MIPS/Register/n131 ), .B(\i_MIPS/Register/n117 ), .Y(
        n42) );
  NAND2X1 U982 ( .A(\i_MIPS/Register/n131 ), .B(\i_MIPS/Register/n119 ), .Y(
        n43) );
  NAND2X1 U983 ( .A(\i_MIPS/Register/n140 ), .B(\i_MIPS/Register/n105 ), .Y(
        n44) );
  NAND2X1 U984 ( .A(\i_MIPS/Register/n140 ), .B(\i_MIPS/Register/n107 ), .Y(
        n45) );
  NAND2X1 U985 ( .A(\i_MIPS/Register/n140 ), .B(\i_MIPS/Register/n109 ), .Y(
        n46) );
  NAND2X1 U986 ( .A(\i_MIPS/Register/n140 ), .B(\i_MIPS/Register/n111 ), .Y(
        n47) );
  NAND2X1 U987 ( .A(\i_MIPS/Register/n140 ), .B(\i_MIPS/Register/n113 ), .Y(
        n48) );
  NAND2X1 U988 ( .A(\i_MIPS/Register/n140 ), .B(\i_MIPS/Register/n115 ), .Y(
        n49) );
  NAND2X1 U989 ( .A(\i_MIPS/Register/n140 ), .B(\i_MIPS/Register/n117 ), .Y(
        n50) );
  NAND2X1 U990 ( .A(\i_MIPS/Register/n140 ), .B(\i_MIPS/Register/n119 ), .Y(
        n51) );
  BUFX12 U991 ( .A(n7071), .Y(n3219) );
  INVX3 U992 ( .A(n3089), .Y(n3086) );
  NAND2X1 U993 ( .A(n2983), .B(n2977), .Y(n2790) );
  CLKINVX1 U994 ( .A(\D_cache/N66 ), .Y(n8755) );
  CLKINVX1 U995 ( .A(n3059), .Y(n2352) );
  CLKBUFX3 U996 ( .A(n2333), .Y(n2349) );
  NAND2X1 U997 ( .A(n2974), .B(n2872), .Y(n2784) );
  NAND2X1 U998 ( .A(n2975), .B(n2873), .Y(n2789) );
  NAND2X1 U999 ( .A(n2976), .B(n2873), .Y(n2787) );
  NAND2X1 U1000 ( .A(n2983), .B(n2871), .Y(n2791) );
  NAND2X1 U1001 ( .A(n2973), .B(n2872), .Y(n2786) );
  NAND2X1 U1002 ( .A(n2978), .B(n2972), .Y(n2773) );
  NAND2X1 U1003 ( .A(n2978), .B(n2973), .Y(n2777) );
  NAND2X1 U1004 ( .A(n2873), .B(n2871), .Y(n2763) );
  NAND2X1 U1005 ( .A(n2977), .B(n2873), .Y(n2788) );
  NAND2X1 U1006 ( .A(n2872), .B(n2870), .Y(n2764) );
  NAND2X1 U1007 ( .A(n2978), .B(n2870), .Y(n2792) );
  INVX6 U1008 ( .A(n3093), .Y(n3091) );
  INVX3 U1009 ( .A(n8714), .Y(n3052) );
  BUFX12 U1010 ( .A(\i_MIPS/ID_EX[79] ), .Y(n3075) );
  CLKBUFX3 U1011 ( .A(n2790), .Y(n3121) );
  INVX6 U1012 ( .A(n1082), .Y(n4016) );
  MXI2X1 U1013 ( .A(\i_MIPS/ID_EX[113] ), .B(\i_MIPS/ID_EX[86] ), .S0(
        \i_MIPS/ID_EX_5 ), .Y(n4774) );
  CLKAND2X3 U1014 ( .A(n1972), .B(n1973), .Y(n56) );
  CLKBUFX3 U1015 ( .A(n3309), .Y(n3304) );
  CLKBUFX3 U1016 ( .A(n3575), .Y(n3568) );
  CLKBUFX3 U1017 ( .A(n3327), .Y(n3349) );
  NAND3XL U1018 ( .A(n2126), .B(n2164), .C(n3062), .Y(\D_cache/n208 ) );
  NAND3XL U1019 ( .A(n2130), .B(n2149), .C(n2208), .Y(\D_cache/n210 ) );
  INVX4 U1020 ( .A(n3041), .Y(n8726) );
  OA22X1 U1021 ( .A0(n8812), .A1(n4006), .B0(n1084), .B1(n4011), .Y(n72) );
  OA22XL U1022 ( .A0(n2751), .A1(n4006), .B0(n8722), .B1(n4010), .Y(n73) );
  OA22X1 U1023 ( .A0(n8811), .A1(n4006), .B0(n1092), .B1(n4010), .Y(n74) );
  OA22X1 U1024 ( .A0(n8810), .A1(n4006), .B0(n1616), .B1(n4010), .Y(n75) );
  AOI22X1 U1025 ( .A0(ICACHE_addr[5]), .A1(mem_read_I), .B0(n3053), .B1(n8688), 
        .Y(n76) );
  AOI22X1 U1026 ( .A0(ICACHE_addr[29]), .A1(mem_read_I), .B0(mem_write_I), 
        .B1(n8712), .Y(n77) );
  CLKBUFX3 U1027 ( .A(n8732), .Y(n3662) );
  BUFX4 U1028 ( .A(n3095), .Y(n3097) );
  BUFX16 U1029 ( .A(n8713), .Y(mem_read_I) );
  INVX12 U1030 ( .A(\D_cache/n522 ), .Y(mem_read_D) );
  BUFX4 U1031 ( .A(n2760), .Y(n3216) );
  BUFX4 U1032 ( .A(n2760), .Y(n3217) );
  AND2X2 U1033 ( .A(n4622), .B(n4724), .Y(n2869) );
  AND2X2 U1034 ( .A(n2979), .B(n2973), .Y(n179) );
  AND2X2 U1035 ( .A(n2982), .B(n2975), .Y(n180) );
  AND2X2 U1036 ( .A(n2982), .B(n2976), .Y(n181) );
  AND2X2 U1037 ( .A(n2981), .B(n2975), .Y(n182) );
  AND2X2 U1038 ( .A(n2981), .B(n2976), .Y(n183) );
  AND2X2 U1039 ( .A(n2982), .B(n2871), .Y(n184) );
  AND2X2 U1040 ( .A(n2982), .B(n2977), .Y(n185) );
  AND2X2 U1041 ( .A(n2981), .B(n2977), .Y(n186) );
  AND2X2 U1042 ( .A(n2980), .B(n2972), .Y(n188) );
  AND2X2 U1043 ( .A(n2980), .B(n2974), .Y(n189) );
  AND2X2 U1044 ( .A(n2979), .B(n2972), .Y(n190) );
  AND2X2 U1045 ( .A(n2979), .B(n2974), .Y(n191) );
  AND2X2 U1046 ( .A(n2980), .B(n2870), .Y(n192) );
  CLKINVX1 U1047 ( .A(n7608), .Y(\i_MIPS/EX_MEM_next[69] ) );
  INVX12 U1048 ( .A(n2730), .Y(n4020) );
  NAND3X2 U1049 ( .A(n1943), .B(n1944), .C(n1945), .Y(n8161) );
  INVX1 U1050 ( .A(n6879), .Y(n8730) );
  CLKINVX1 U1051 ( .A(n3059), .Y(n2350) );
  CLKBUFX3 U1052 ( .A(n2331), .Y(n2341) );
  CLKBUFX3 U1053 ( .A(n3646), .Y(n3647) );
  NAND2X1 U1054 ( .A(n10), .B(n8686), .Y(n947) );
  AOI22X1 U1055 ( .A0(ICACHE_addr[6]), .A1(mem_read_I), .B0(n3054), .B1(n8689), 
        .Y(n948) );
  AOI22X1 U1056 ( .A0(ICACHE_addr[7]), .A1(mem_read_I), .B0(n3055), .B1(n8690), 
        .Y(n949) );
  AOI22X1 U1057 ( .A0(ICACHE_addr[8]), .A1(mem_read_I), .B0(n3053), .B1(n8691), 
        .Y(n950) );
  AOI22X1 U1058 ( .A0(ICACHE_addr[9]), .A1(mem_read_I), .B0(n3054), .B1(n8692), 
        .Y(n951) );
  AOI22X1 U1059 ( .A0(ICACHE_addr[10]), .A1(mem_read_I), .B0(n3055), .B1(n8693), .Y(n952) );
  AOI22X1 U1060 ( .A0(ICACHE_addr[11]), .A1(mem_read_I), .B0(n3053), .B1(n8694), .Y(n953) );
  AOI22X1 U1061 ( .A0(ICACHE_addr[12]), .A1(mem_read_I), .B0(n3054), .B1(n8695), .Y(n954) );
  AOI22X1 U1062 ( .A0(ICACHE_addr[13]), .A1(mem_read_I), .B0(n3055), .B1(n8696), .Y(n955) );
  AOI22X1 U1063 ( .A0(ICACHE_addr[14]), .A1(mem_read_I), .B0(n3053), .B1(n8697), .Y(n956) );
  AOI22X1 U1064 ( .A0(ICACHE_addr[18]), .A1(mem_read_I), .B0(mem_write_I), 
        .B1(n8701), .Y(n957) );
  AOI22X1 U1065 ( .A0(ICACHE_addr[19]), .A1(mem_read_I), .B0(mem_write_I), 
        .B1(n8702), .Y(n958) );
  AOI22X1 U1066 ( .A0(ICACHE_addr[20]), .A1(mem_read_I), .B0(mem_write_I), 
        .B1(n8703), .Y(n959) );
  AOI22X1 U1067 ( .A0(ICACHE_addr[25]), .A1(mem_read_I), .B0(mem_write_I), 
        .B1(n8708), .Y(n960) );
  AOI22X1 U1068 ( .A0(ICACHE_addr[28]), .A1(mem_read_I), .B0(mem_write_I), 
        .B1(n8711), .Y(n961) );
  AOI22X1 U1069 ( .A0(ICACHE_addr[15]), .A1(mem_read_I), .B0(n3054), .B1(n8698), .Y(n962) );
  CLKINVX1 U1070 ( .A(n7045), .Y(n8719) );
  INVX1 U1071 ( .A(n3041), .Y(n3019) );
  NOR2BX1 U1072 ( .AN(\D_cache/n202 ), .B(\D_cache/n216 ), .Y(\D_cache/n251 )
         );
  CLKBUFX3 U1073 ( .A(\D_cache/n251 ), .Y(n3987) );
  CLKBUFX3 U1074 ( .A(\D_cache/n251 ), .Y(n3988) );
  AND2X4 U1075 ( .A(n8903), .B(\D_cache/n200 ), .Y(n2867) );
  INVX6 U1076 ( .A(n2867), .Y(n3039) );
  NOR2BX1 U1077 ( .AN(\D_cache/n201 ), .B(\D_cache/n216 ), .Y(\D_cache/n388 )
         );
  CLKBUFX3 U1078 ( .A(\D_cache/n388 ), .Y(n3994) );
  CLKBUFX3 U1079 ( .A(\D_cache/n388 ), .Y(n3993) );
  NOR2BX1 U1080 ( .AN(\D_cache/n203 ), .B(\D_cache/n216 ), .Y(\D_cache/n320 )
         );
  CLKBUFX3 U1081 ( .A(\D_cache/n320 ), .Y(n3990) );
  CLKBUFX3 U1082 ( .A(\D_cache/n320 ), .Y(n3991) );
  AOI22X2 U1083 ( .A0(n10297), .A1(n2808), .B0(\D_cache/N32 ), .B1(n8551), .Y(
        n965) );
  INVX3 U1084 ( .A(n10300), .Y(n8722) );
  AND2X2 U1085 ( .A(\D_cache/n201 ), .B(\D_cache/n200 ), .Y(n968) );
  NAND2X1 U1086 ( .A(\i_MIPS/ALUin1[27] ), .B(n4703), .Y(n6763) );
  NAND3X1 U1087 ( .A(n3957), .B(n8772), .C(\D_cache/n518 ), .Y(\D_cache/n522 )
         );
  INVX16 U1088 ( .A(n3578), .Y(n3577) );
  CLKINVX1 U1089 ( .A(\D_cache/N171 ), .Y(n8889) );
  CLKBUFX3 U1090 ( .A(n2907), .Y(n3088) );
  CLKINVX1 U1091 ( .A(\D_cache/N167 ), .Y(n8885) );
  CLKINVX1 U1092 ( .A(\D_cache/N158 ), .Y(n8876) );
  CLKINVX1 U1093 ( .A(\D_cache/N173 ), .Y(n8891) );
  CLKINVX1 U1094 ( .A(\D_cache/N157 ), .Y(n8875) );
  CLKMX2X2 U1095 ( .A(\i_MIPS/n283 ), .B(n2993), .S0(n4019), .Y(n4653) );
  NAND4BX1 U1096 ( .AN(n2794), .B(n3165), .C(n4770), .D(n4769), .Y(n7046) );
  CLKBUFX3 U1097 ( .A(n3104), .Y(n3102) );
  INVX3 U1098 ( .A(n3112), .Y(n3107) );
  INVX6 U1099 ( .A(n3112), .Y(n3106) );
  NAND3X2 U1100 ( .A(n1976), .B(n1977), .C(n1978), .Y(n8214) );
  NAND2X1 U1101 ( .A(\D_cache/N30 ), .B(DCACHE_ren), .Y(n1074) );
  CLKMX2X2 U1102 ( .A(\i_MIPS/n295 ), .B(n8), .S0(n4019), .Y(n4673) );
  CLKINVX1 U1103 ( .A(n8685), .Y(n8714) );
  CLKBUFX6 U1104 ( .A(n2828), .Y(n3597) );
  BUFX4 U1105 ( .A(n7069), .Y(n3214) );
  CLKBUFX3 U1106 ( .A(n2774), .Y(n3157) );
  CLKBUFX3 U1107 ( .A(n180), .Y(n3138) );
  CLKBUFX3 U1108 ( .A(n184), .Y(n3144) );
  CLKBUFX3 U1109 ( .A(n182), .Y(n3150) );
  AND3X4 U1110 ( .A(n1948), .B(n1949), .C(n1950), .Y(n1086) );
  INVX16 U1111 ( .A(n4020), .Y(n4019) );
  NAND3X2 U1112 ( .A(n1935), .B(n1936), .C(n1937), .Y(n8258) );
  INVX3 U1113 ( .A(n2722), .Y(n4041) );
  CLKMX2X2 U1114 ( .A(\i_MIPS/n303 ), .B(n2887), .S0(n4019), .Y(n4680) );
  OA22X1 U1115 ( .A0(n3462), .A1(n143), .B0(n3441), .B1(n1024), .Y(n4477) );
  CLKINVX1 U1116 ( .A(n4772), .Y(n8718) );
  BUFX4 U1117 ( .A(n8718), .Y(n3638) );
  CLKINVX1 U1118 ( .A(n5933), .Y(n8721) );
  BUFX4 U1119 ( .A(\i_MIPS/IR_ID[25] ), .Y(n4013) );
  CLKINVX1 U1120 ( .A(n5860), .Y(n8720) );
  CLKINVX1 U1121 ( .A(n6800), .Y(n8723) );
  BUFX4 U1122 ( .A(n3664), .Y(n3665) );
  INVX3 U1123 ( .A(mem_write_D), .Y(n4007) );
  INVX3 U1124 ( .A(mem_write_D), .Y(n4006) );
  CLKINVX1 U1125 ( .A(n6972), .Y(n7976) );
  INVX3 U1126 ( .A(n4027), .Y(n2109) );
  NAND2X6 U1127 ( .A(n7046), .B(n3164), .Y(n2761) );
  NAND4X4 U1128 ( .A(n6075), .B(n6074), .C(n5), .D(n6072), .Y(n8263) );
  NAND2X1 U1129 ( .A(\i_MIPS/ALUin1[29] ), .B(n4705), .Y(n5821) );
  NAND3X6 U1130 ( .A(n8292), .B(n8291), .C(n8290), .Y(n8320) );
  CLKAND2X12 U1131 ( .A(ICACHE_addr[2]), .B(n8686), .Y(mem_addr_I[4]) );
  AO22X2 U1132 ( .A0(n3602), .A1(ICACHE_addr[16]), .B0(n3601), .B1(n8699), .Y(
        n8450) );
  AO22X2 U1133 ( .A0(n3606), .A1(ICACHE_addr[17]), .B0(n3600), .B1(n8700), .Y(
        n8454) );
  INVX12 U1134 ( .A(n76), .Y(mem_addr_I[7]) );
  INVX12 U1135 ( .A(n948), .Y(mem_addr_I[8]) );
  INVX12 U1136 ( .A(n949), .Y(mem_addr_I[9]) );
  INVX12 U1137 ( .A(n950), .Y(mem_addr_I[10]) );
  INVX12 U1138 ( .A(n951), .Y(mem_addr_I[11]) );
  INVX12 U1139 ( .A(n952), .Y(mem_addr_I[12]) );
  INVX12 U1140 ( .A(n953), .Y(mem_addr_I[13]) );
  INVX12 U1141 ( .A(n954), .Y(mem_addr_I[14]) );
  INVX12 U1142 ( .A(n955), .Y(mem_addr_I[15]) );
  INVX12 U1143 ( .A(n956), .Y(mem_addr_I[16]) );
  INVX12 U1144 ( .A(n957), .Y(mem_addr_I[20]) );
  INVX12 U1145 ( .A(n958), .Y(mem_addr_I[21]) );
  INVX12 U1146 ( .A(n959), .Y(mem_addr_I[22]) );
  INVX12 U1147 ( .A(n960), .Y(mem_addr_I[27]) );
  INVX12 U1148 ( .A(n961), .Y(mem_addr_I[30]) );
  INVX12 U1149 ( .A(n77), .Y(mem_addr_I[31]) );
  INVX12 U1150 ( .A(n75), .Y(mem_addr_D[30]) );
  INVX12 U1151 ( .A(n74), .Y(mem_addr_D[29]) );
  INVX12 U1152 ( .A(n73), .Y(mem_addr_D[28]) );
  INVX12 U1153 ( .A(n72), .Y(mem_addr_D[27]) );
  CLKAND2X12 U1154 ( .A(n3633), .B(n8554), .Y(mem_wdata_I[0]) );
  CLKAND2X12 U1155 ( .A(n3633), .B(n8555), .Y(mem_wdata_I[1]) );
  CLKAND2X12 U1156 ( .A(n3633), .B(n8556), .Y(mem_wdata_I[2]) );
  CLKAND2X12 U1157 ( .A(n3633), .B(n8557), .Y(mem_wdata_I[3]) );
  CLKAND2X12 U1158 ( .A(n3633), .B(n8558), .Y(mem_wdata_I[4]) );
  CLKAND2X12 U1159 ( .A(n3633), .B(n8559), .Y(mem_wdata_I[5]) );
  CLKAND2X12 U1160 ( .A(n3633), .B(n8560), .Y(mem_wdata_I[6]) );
  CLKAND2X12 U1161 ( .A(n3633), .B(n8561), .Y(mem_wdata_I[7]) );
  CLKAND2X12 U1162 ( .A(n3633), .B(n8562), .Y(mem_wdata_I[8]) );
  CLKAND2X12 U1163 ( .A(n3633), .B(n8563), .Y(mem_wdata_I[9]) );
  CLKAND2X12 U1164 ( .A(n3633), .B(n8564), .Y(mem_wdata_I[10]) );
  CLKAND2X12 U1165 ( .A(n3633), .B(n8565), .Y(mem_wdata_I[11]) );
  CLKAND2X12 U1166 ( .A(n3633), .B(n8566), .Y(mem_wdata_I[12]) );
  CLKAND2X12 U1167 ( .A(n3633), .B(n8567), .Y(mem_wdata_I[13]) );
  CLKAND2X12 U1168 ( .A(n3633), .B(n8568), .Y(mem_wdata_I[14]) );
  CLKAND2X12 U1169 ( .A(n3633), .B(n8569), .Y(mem_wdata_I[15]) );
  CLKAND2X12 U1170 ( .A(n3633), .B(n8570), .Y(mem_wdata_I[16]) );
  CLKAND2X12 U1171 ( .A(n3633), .B(n8571), .Y(mem_wdata_I[17]) );
  CLKAND2X12 U1172 ( .A(n3633), .B(n8572), .Y(mem_wdata_I[18]) );
  CLKAND2X12 U1173 ( .A(n3633), .B(n8573), .Y(mem_wdata_I[19]) );
  CLKAND2X12 U1174 ( .A(n3633), .B(n8574), .Y(mem_wdata_I[20]) );
  CLKAND2X12 U1175 ( .A(n3633), .B(n8575), .Y(mem_wdata_I[21]) );
  CLKAND2X12 U1176 ( .A(n3633), .B(n8576), .Y(mem_wdata_I[22]) );
  CLKAND2X12 U1177 ( .A(n3633), .B(n8577), .Y(mem_wdata_I[23]) );
  CLKAND2X12 U1178 ( .A(n3633), .B(n8578), .Y(mem_wdata_I[24]) );
  CLKAND2X12 U1179 ( .A(n3633), .B(n8579), .Y(mem_wdata_I[25]) );
  CLKAND2X12 U1180 ( .A(n3633), .B(n8580), .Y(mem_wdata_I[26]) );
  CLKAND2X12 U1181 ( .A(n3633), .B(n8581), .Y(mem_wdata_I[27]) );
  CLKAND2X12 U1182 ( .A(n3633), .B(n8582), .Y(mem_wdata_I[28]) );
  CLKAND2X12 U1183 ( .A(n3633), .B(n8583), .Y(mem_wdata_I[29]) );
  CLKAND2X12 U1184 ( .A(n3633), .B(n8584), .Y(mem_wdata_I[30]) );
  CLKAND2X12 U1185 ( .A(n3633), .B(n8585), .Y(mem_wdata_I[31]) );
  CLKAND2X12 U1186 ( .A(n3633), .B(n8586), .Y(mem_wdata_I[32]) );
  CLKAND2X12 U1187 ( .A(n3633), .B(n8587), .Y(mem_wdata_I[33]) );
  CLKAND2X12 U1188 ( .A(n3633), .B(n8588), .Y(mem_wdata_I[34]) );
  CLKAND2X12 U1189 ( .A(n3633), .B(n8589), .Y(mem_wdata_I[35]) );
  CLKAND2X12 U1190 ( .A(n3633), .B(n8590), .Y(mem_wdata_I[36]) );
  CLKAND2X12 U1191 ( .A(n3633), .B(n8591), .Y(mem_wdata_I[37]) );
  CLKAND2X12 U1192 ( .A(n3633), .B(n8592), .Y(mem_wdata_I[38]) );
  CLKAND2X12 U1193 ( .A(n3633), .B(n8593), .Y(mem_wdata_I[39]) );
  CLKAND2X12 U1194 ( .A(n3633), .B(n8594), .Y(mem_wdata_I[40]) );
  CLKAND2X12 U1195 ( .A(n3633), .B(n8595), .Y(mem_wdata_I[41]) );
  BUFX12 U1196 ( .A(n8714), .Y(n3633) );
  CLKAND2X12 U1197 ( .A(n3633), .B(n8596), .Y(mem_wdata_I[42]) );
  CLKAND2X12 U1198 ( .A(n3633), .B(n8597), .Y(mem_wdata_I[43]) );
  CLKAND2X12 U1199 ( .A(n3633), .B(n8598), .Y(mem_wdata_I[44]) );
  CLKAND2X12 U1200 ( .A(n3633), .B(n8599), .Y(mem_wdata_I[45]) );
  CLKAND2X12 U1201 ( .A(n3633), .B(n8600), .Y(mem_wdata_I[46]) );
  CLKAND2X12 U1202 ( .A(n3633), .B(n8601), .Y(mem_wdata_I[47]) );
  CLKAND2X12 U1203 ( .A(n3055), .B(n8602), .Y(mem_wdata_I[48]) );
  CLKAND2X12 U1204 ( .A(n3055), .B(n8603), .Y(mem_wdata_I[49]) );
  CLKAND2X12 U1205 ( .A(n3053), .B(n8604), .Y(mem_wdata_I[50]) );
  CLKAND2X12 U1206 ( .A(n3054), .B(n8605), .Y(mem_wdata_I[51]) );
  CLKAND2X12 U1207 ( .A(n3055), .B(n8606), .Y(mem_wdata_I[52]) );
  CLKAND2X12 U1208 ( .A(n3053), .B(n8607), .Y(mem_wdata_I[53]) );
  CLKAND2X12 U1209 ( .A(n3054), .B(n8608), .Y(mem_wdata_I[54]) );
  CLKAND2X12 U1210 ( .A(n3055), .B(n8609), .Y(mem_wdata_I[55]) );
  CLKAND2X12 U1211 ( .A(n3053), .B(n8610), .Y(mem_wdata_I[56]) );
  CLKAND2X12 U1212 ( .A(n3054), .B(n8611), .Y(mem_wdata_I[57]) );
  CLKAND2X12 U1213 ( .A(n3055), .B(n8612), .Y(mem_wdata_I[58]) );
  CLKAND2X12 U1214 ( .A(n3053), .B(n8613), .Y(mem_wdata_I[59]) );
  CLKAND2X12 U1215 ( .A(n3054), .B(n8614), .Y(mem_wdata_I[60]) );
  CLKAND2X12 U1216 ( .A(n3055), .B(n8615), .Y(mem_wdata_I[61]) );
  CLKAND2X12 U1217 ( .A(n3053), .B(n8616), .Y(mem_wdata_I[62]) );
  CLKAND2X12 U1218 ( .A(n3054), .B(n8617), .Y(mem_wdata_I[63]) );
  CLKAND2X12 U1219 ( .A(n3055), .B(n8618), .Y(mem_wdata_I[64]) );
  CLKAND2X12 U1220 ( .A(n3053), .B(n8619), .Y(mem_wdata_I[65]) );
  CLKAND2X12 U1221 ( .A(n3054), .B(n8620), .Y(mem_wdata_I[66]) );
  CLKAND2X12 U1222 ( .A(n3055), .B(n8621), .Y(mem_wdata_I[67]) );
  CLKAND2X12 U1223 ( .A(n3053), .B(n8622), .Y(mem_wdata_I[68]) );
  CLKAND2X12 U1224 ( .A(n3054), .B(n8623), .Y(mem_wdata_I[69]) );
  CLKAND2X12 U1225 ( .A(n3055), .B(n8624), .Y(mem_wdata_I[70]) );
  CLKAND2X12 U1226 ( .A(n3053), .B(n8625), .Y(mem_wdata_I[71]) );
  CLKAND2X12 U1227 ( .A(n3054), .B(n8626), .Y(mem_wdata_I[72]) );
  CLKAND2X12 U1228 ( .A(n3055), .B(n8627), .Y(mem_wdata_I[73]) );
  CLKAND2X12 U1229 ( .A(n3053), .B(n8628), .Y(mem_wdata_I[74]) );
  CLKAND2X12 U1230 ( .A(n3054), .B(n8629), .Y(mem_wdata_I[75]) );
  CLKAND2X12 U1231 ( .A(n3055), .B(n8630), .Y(mem_wdata_I[76]) );
  CLKAND2X12 U1232 ( .A(n3053), .B(n8631), .Y(mem_wdata_I[77]) );
  CLKAND2X12 U1233 ( .A(n3054), .B(n8632), .Y(mem_wdata_I[78]) );
  INVX8 U1234 ( .A(n3052), .Y(n3054) );
  CLKAND2X12 U1235 ( .A(n3055), .B(n8633), .Y(mem_wdata_I[79]) );
  CLKAND2X12 U1236 ( .A(n3053), .B(n8634), .Y(mem_wdata_I[80]) );
  INVX8 U1237 ( .A(n3052), .Y(n3053) );
  CLKAND2X12 U1238 ( .A(n3054), .B(n8635), .Y(mem_wdata_I[81]) );
  CLKAND2X12 U1239 ( .A(n3055), .B(n8636), .Y(mem_wdata_I[82]) );
  CLKAND2X12 U1240 ( .A(n3053), .B(n8637), .Y(mem_wdata_I[83]) );
  CLKAND2X12 U1241 ( .A(n3054), .B(n8638), .Y(mem_wdata_I[84]) );
  CLKAND2X12 U1242 ( .A(n3055), .B(n8639), .Y(mem_wdata_I[85]) );
  CLKAND2X12 U1243 ( .A(n3053), .B(n8640), .Y(mem_wdata_I[86]) );
  CLKAND2X12 U1244 ( .A(n3054), .B(n8641), .Y(mem_wdata_I[87]) );
  CLKAND2X12 U1245 ( .A(n3055), .B(n8642), .Y(mem_wdata_I[88]) );
  INVX8 U1246 ( .A(n3052), .Y(n3055) );
  CLKAND2X12 U1247 ( .A(n3053), .B(n8643), .Y(mem_wdata_I[89]) );
  CLKAND2X12 U1248 ( .A(n3054), .B(n8644), .Y(mem_wdata_I[90]) );
  CLKAND2X12 U1249 ( .A(n3055), .B(n8645), .Y(mem_wdata_I[91]) );
  CLKAND2X12 U1250 ( .A(n3053), .B(n8646), .Y(mem_wdata_I[92]) );
  CLKAND2X12 U1251 ( .A(n3054), .B(n8647), .Y(mem_wdata_I[93]) );
  CLKAND2X12 U1252 ( .A(n3055), .B(n8648), .Y(mem_wdata_I[94]) );
  CLKAND2X12 U1253 ( .A(n3053), .B(n8649), .Y(mem_wdata_I[95]) );
  CLKAND2X12 U1254 ( .A(n3054), .B(n8650), .Y(mem_wdata_I[96]) );
  CLKAND2X12 U1255 ( .A(n3055), .B(n8651), .Y(mem_wdata_I[97]) );
  CLKAND2X12 U1256 ( .A(n3053), .B(n8652), .Y(mem_wdata_I[98]) );
  CLKAND2X12 U1257 ( .A(n3054), .B(n8653), .Y(mem_wdata_I[99]) );
  CLKAND2X12 U1258 ( .A(n3055), .B(n8654), .Y(mem_wdata_I[100]) );
  CLKAND2X12 U1259 ( .A(n3053), .B(n8655), .Y(mem_wdata_I[101]) );
  CLKAND2X12 U1260 ( .A(n3054), .B(n8656), .Y(mem_wdata_I[102]) );
  CLKAND2X12 U1261 ( .A(n3055), .B(n8657), .Y(mem_wdata_I[103]) );
  CLKAND2X12 U1262 ( .A(n3053), .B(n8658), .Y(mem_wdata_I[104]) );
  CLKAND2X12 U1263 ( .A(n3054), .B(n8659), .Y(mem_wdata_I[105]) );
  CLKAND2X12 U1264 ( .A(n3055), .B(n8660), .Y(mem_wdata_I[106]) );
  CLKAND2X12 U1265 ( .A(n3053), .B(n8661), .Y(mem_wdata_I[107]) );
  CLKAND2X12 U1266 ( .A(n3054), .B(n8662), .Y(mem_wdata_I[108]) );
  CLKAND2X12 U1267 ( .A(n3055), .B(n8663), .Y(mem_wdata_I[109]) );
  CLKAND2X12 U1268 ( .A(n3053), .B(n8664), .Y(mem_wdata_I[110]) );
  CLKAND2X12 U1269 ( .A(n3054), .B(n8665), .Y(mem_wdata_I[111]) );
  CLKAND2X12 U1270 ( .A(n3055), .B(n8666), .Y(mem_wdata_I[112]) );
  CLKAND2X12 U1271 ( .A(n3053), .B(n8667), .Y(mem_wdata_I[113]) );
  CLKAND2X12 U1272 ( .A(n3054), .B(n8668), .Y(mem_wdata_I[114]) );
  CLKAND2X12 U1273 ( .A(n3055), .B(n8669), .Y(mem_wdata_I[115]) );
  CLKAND2X12 U1274 ( .A(n3053), .B(n8670), .Y(mem_wdata_I[116]) );
  CLKAND2X12 U1275 ( .A(n3054), .B(n8671), .Y(mem_wdata_I[117]) );
  CLKAND2X12 U1276 ( .A(n3055), .B(n8672), .Y(mem_wdata_I[118]) );
  CLKAND2X12 U1277 ( .A(n3053), .B(n8673), .Y(mem_wdata_I[119]) );
  CLKAND2X12 U1278 ( .A(n3054), .B(n8674), .Y(mem_wdata_I[120]) );
  CLKAND2X12 U1279 ( .A(n3055), .B(n8675), .Y(mem_wdata_I[121]) );
  CLKAND2X12 U1280 ( .A(n3053), .B(n8676), .Y(mem_wdata_I[122]) );
  CLKAND2X12 U1281 ( .A(n3054), .B(n8677), .Y(mem_wdata_I[123]) );
  CLKAND2X12 U1282 ( .A(n3055), .B(n8678), .Y(mem_wdata_I[124]) );
  CLKAND2X12 U1283 ( .A(n3053), .B(n8679), .Y(mem_wdata_I[125]) );
  CLKAND2X12 U1284 ( .A(n3054), .B(n8680), .Y(mem_wdata_I[126]) );
  CLKAND2X12 U1285 ( .A(n3055), .B(n8681), .Y(mem_wdata_I[127]) );
  INVXL U1286 ( .A(n10211), .Y(n1915) );
  INVX12 U1287 ( .A(n1915), .Y(mem_wdata_D[84]) );
  NOR2BX1 U1288 ( .AN(\D_cache/N132 ), .B(n4006), .Y(n10211) );
  INVXL U1289 ( .A(n10212), .Y(n1917) );
  INVX12 U1290 ( .A(n1917), .Y(mem_wdata_D[83]) );
  NOR2BX1 U1291 ( .AN(\D_cache/N133 ), .B(n4007), .Y(n10212) );
  INVXL U1292 ( .A(n10213), .Y(n1919) );
  INVX12 U1293 ( .A(n1919), .Y(mem_wdata_D[82]) );
  NOR2BX1 U1294 ( .AN(\D_cache/N134 ), .B(n4006), .Y(n10213) );
  INVXL U1295 ( .A(n10227), .Y(n1921) );
  INVX12 U1296 ( .A(n1921), .Y(mem_wdata_D[68]) );
  NOR2BX1 U1297 ( .AN(\D_cache/N148 ), .B(n3998), .Y(n10227) );
  INVXL U1298 ( .A(n10229), .Y(n1923) );
  INVX12 U1299 ( .A(n1923), .Y(mem_wdata_D[66]) );
  NOR2BX1 U1300 ( .AN(\D_cache/N150 ), .B(n4004), .Y(n10229) );
  INVXL U1301 ( .A(n10230), .Y(n1925) );
  INVX12 U1302 ( .A(n1925), .Y(mem_wdata_D[65]) );
  NOR2BX1 U1303 ( .AN(\D_cache/N151 ), .B(n4005), .Y(n10230) );
  INVXL U1304 ( .A(n10231), .Y(n1927) );
  INVX12 U1305 ( .A(n1927), .Y(mem_wdata_D[64]) );
  NOR2BX1 U1306 ( .AN(\D_cache/N152 ), .B(n4000), .Y(n10231) );
  INVX12 U1307 ( .A(n947), .Y(mem_addr_I[5]) );
  AOI211X2 U1308 ( .A0(n8922), .A1(n5051), .B0(n5050), .C0(n5049), .Y(n5057)
         );
  XOR3X1 U1309 ( .A(n7899), .B(n7885), .C(n7898), .Y(n7888) );
  INVX1 U1310 ( .A(n7898), .Y(n7896) );
  OR2X1 U1311 ( .A(n7835), .B(n3049), .Y(n2039) );
  OR2X1 U1312 ( .A(n8386), .B(n3049), .Y(n1987) );
  INVX1 U1313 ( .A(n7908), .Y(n7915) );
  AND3X8 U1314 ( .A(n7787), .B(n7831), .C(n7830), .Y(n3047) );
  CLKXOR2X8 U1315 ( .A(n22), .B(n7073), .Y(n7830) );
  NAND2BX2 U1316 ( .AN(n3576), .B(n8559), .Y(n7408) );
  NAND2X2 U1317 ( .A(n7851), .B(n7850), .Y(n7865) );
  AND2X8 U1318 ( .A(n6993), .B(n4724), .Y(n2865) );
  OR2X1 U1319 ( .A(n8371), .B(n3049), .Y(n1993) );
  CLKMX2X2 U1320 ( .A(n5254), .B(n5616), .S0(n4016), .Y(n6831) );
  OAI221X1 U1321 ( .A0(\i_MIPS/n347 ), .A1(n14), .B0(\i_MIPS/n348 ), .B1(n3077), .C0(n4967), .Y(n5254) );
  NAND2BX4 U1322 ( .AN(n5538), .B(n6400), .Y(n6324) );
  INVX3 U1323 ( .A(n4674), .Y(n4672) );
  AND2X6 U1324 ( .A(n2862), .B(n7836), .Y(n2828) );
  NAND3BX4 U1325 ( .AN(n4728), .B(n4725), .C(n2819), .Y(n6848) );
  MX2XL U1326 ( .A(n2799), .B(n7732), .S0(n3623), .Y(\i_MIPS/n437 ) );
  NAND2XL U1327 ( .A(n8481), .B(n6389), .Y(n6399) );
  INVX4 U1328 ( .A(n6389), .Y(n8479) );
  NOR2X8 U1329 ( .A(n5454), .B(n5453), .Y(n5809) );
  NAND4X6 U1330 ( .A(n5181), .B(n5180), .C(n5179), .D(n5178), .Y(n5454) );
  INVX1 U1331 ( .A(n4632), .Y(n4633) );
  OA22X1 U1332 ( .A0(n6549), .A1(n5752), .B0(n6056), .B1(n6547), .Y(n5625) );
  AO21X1 U1333 ( .A0(n5612), .A1(n3076), .B0(n5613), .Y(n6547) );
  OAI22X2 U1334 ( .A0(n8909), .A1(n8805), .B0(n2841), .B1(n8909), .Y(n8910) );
  INVX3 U1335 ( .A(n7862), .Y(n7867) );
  NAND2X2 U1336 ( .A(n8504), .B(n8502), .Y(n4900) );
  CLKINVX1 U1337 ( .A(n4900), .Y(n4591) );
  NAND3BX1 U1338 ( .AN(n5834), .B(n5833), .C(n3102), .Y(n5835) );
  XNOR2X2 U1339 ( .A(n8163), .B(n8161), .Y(n6751) );
  NAND4X4 U1340 ( .A(n6752), .B(n6751), .C(n6750), .D(n6749), .Y(n6977) );
  NAND2X1 U1341 ( .A(\D_cache/n202 ), .B(\D_cache/n200 ), .Y(\D_cache/n165 )
         );
  NAND4X4 U1342 ( .A(n7685), .B(n7684), .C(n7683), .D(n7682), .Y(n8211) );
  NAND2X4 U1343 ( .A(n2731), .B(n2732), .Y(n4681) );
  MXI2X2 U1344 ( .A(DCACHE_addr[12]), .B(DCACHE_rdata[14]), .S0(n4022), .Y(
        n8725) );
  OAI221X4 U1345 ( .A0(\i_MIPS/n364 ), .A1(n3091), .B0(\i_MIPS/n363 ), .B1(
        n3085), .C0(n5201), .Y(n6330) );
  CLKMX2X2 U1346 ( .A(n6331), .B(n6330), .S0(n4016), .Y(n6679) );
  OAI2BB1X4 U1347 ( .A0N(n6762), .A1N(n6765), .B0(n6763), .Y(n5893) );
  AND2X4 U1348 ( .A(ICACHE_addr[4]), .B(n10), .Y(n2901) );
  CLKINVX4 U1349 ( .A(n10), .Y(n4387) );
  NAND2X2 U1350 ( .A(n7981), .B(n7980), .Y(n8020) );
  INVX3 U1351 ( .A(n4652), .Y(n4662) );
  OAI2BB1X4 U1352 ( .A0N(n5810), .A1N(n8531), .B0(n8533), .Y(n6982) );
  NAND2X1 U1353 ( .A(n8488), .B(n8485), .Y(n4824) );
  CLKAND2X12 U1354 ( .A(n2733), .B(n2734), .Y(n8382) );
  CLKINVX8 U1355 ( .A(n8130), .Y(n2162) );
  CLKXOR2X1 U1356 ( .A(n7819), .B(ICACHE_addr[2]), .Y(n8387) );
  OR2X2 U1357 ( .A(n8339), .B(n3049), .Y(n1990) );
  OR2X2 U1358 ( .A(n7959), .B(n3049), .Y(n2741) );
  OR2XL U1359 ( .A(n7990), .B(n3049), .Y(n2009) );
  NAND2X1 U1360 ( .A(n4686), .B(\i_MIPS/n364 ), .Y(n8509) );
  NAND4X4 U1361 ( .A(n7583), .B(n7582), .C(n7581), .D(n7580), .Y(n7967) );
  OA22X1 U1362 ( .A0(n8359), .A1(n3599), .B0(n2158), .B1(n8358), .Y(n8360) );
  NOR4X1 U1363 ( .A(n4659), .B(n5682), .C(n4816), .D(n5749), .Y(n4697) );
  INVX3 U1364 ( .A(n4829), .Y(n4659) );
  INVX3 U1365 ( .A(n6400), .Y(n4665) );
  CLKINVX1 U1366 ( .A(n5535), .Y(n4655) );
  XOR2X4 U1367 ( .A(n8295), .B(n8283), .Y(n5884) );
  CLKINVX1 U1368 ( .A(n7010), .Y(n5817) );
  OA22X1 U1369 ( .A0(n7011), .A1(n7010), .B0(n7009), .B1(n7008), .Y(n7012) );
  AOI22X1 U1370 ( .A0(\D_cache/N139 ), .A1(n2153), .B0(n3032), .B1(
        \D_cache/N171 ), .Y(\D_cache/n195 ) );
  OAI222X2 U1371 ( .A0(n5598), .A1(n3164), .B0(n5576), .B1(n2761), .C0(n8724), 
        .C1(n3163), .Y(n7958) );
  XNOR2X1 U1372 ( .A(n1084), .B(\D_cache/N36 ), .Y(\D_cache/n553 ) );
  OAI222X2 U1373 ( .A0(n6319), .A1(n3219), .B0(n6318), .B1(n3217), .C0(n8729), 
        .C1(n3214), .Y(n8222) );
  NAND2X2 U1374 ( .A(n8060), .B(n8059), .Y(n8063) );
  NAND2X2 U1375 ( .A(n8043), .B(n3577), .Y(n8060) );
  NAND2X2 U1376 ( .A(n8026), .B(n3577), .Y(n8059) );
  NAND2BX4 U1377 ( .AN(n3576), .B(n8555), .Y(n7412) );
  CLKAND2X3 U1378 ( .A(n3579), .B(n7996), .Y(n2859) );
  OAI222X2 U1379 ( .A0(n5671), .A1(n3218), .B0(n5670), .B1(n3217), .C0(n8717), 
        .C1(n3215), .Y(n8014) );
  OAI221X4 U1380 ( .A0(\i_MIPS/n341 ), .A1(n3091), .B0(\i_MIPS/n342 ), .B1(
        n3086), .C0(n4968), .Y(n5616) );
  CLKMX2X2 U1381 ( .A(n5103), .B(n5102), .S0(n4015), .Y(n5104) );
  INVX4 U1382 ( .A(n8257), .Y(n5105) );
  CLKINVX6 U1383 ( .A(n5470), .Y(n4605) );
  OAI221X1 U1384 ( .A0(n6332), .A1(n6772), .B0(n3068), .B1(n6836), .C0(n4717), 
        .Y(n5546) );
  OAI221X4 U1385 ( .A0(\i_MIPS/n371 ), .A1(n3092), .B0(\i_MIPS/n370 ), .B1(
        n3087), .C0(n4713), .Y(n6772) );
  MXI2X8 U1386 ( .A(n10316), .B(DCACHE_rdata[12]), .S0(n4021), .Y(n8729) );
  INVX3 U1387 ( .A(n8266), .Y(n5956) );
  INVX1 U1388 ( .A(n5889), .Y(n5892) );
  AOI221X1 U1389 ( .A0(n5897), .A1(n5896), .B0(n5895), .B1(n5894), .C0(n6766), 
        .Y(n5910) );
  AND3X8 U1390 ( .A(n8188), .B(n8187), .C(n8186), .Y(n8196) );
  NAND3X6 U1391 ( .A(n8017), .B(n8019), .C(n8018), .Y(n8088) );
  NAND2X6 U1392 ( .A(n2715), .B(n7384), .Y(n8402) );
  INVX4 U1393 ( .A(n6257), .Y(n5537) );
  XNOR2X4 U1394 ( .A(n1086), .B(n7810), .Y(n5804) );
  NAND4X8 U1395 ( .A(n4396), .B(n4395), .C(n4394), .D(n4393), .Y(n8701) );
  INVX4 U1396 ( .A(n6848), .Y(n5484) );
  NAND2XL U1397 ( .A(n8465), .B(n8547), .Y(n4837) );
  NAND2X1 U1398 ( .A(n4642), .B(\i_MIPS/n351 ), .Y(n4833) );
  OA22X1 U1399 ( .A0(n8217), .A1(n3599), .B0(n2158), .B1(n8216), .Y(n8218) );
  OR2X1 U1400 ( .A(n8416), .B(n18), .Y(n2013) );
  OAI222X2 U1401 ( .A0(n6747), .A1(n3166), .B0(n6746), .B1(n2761), .C0(n3022), 
        .C1(n3162), .Y(n6748) );
  NAND2X2 U1402 ( .A(n4682), .B(n5381), .Y(n6621) );
  INVX12 U1403 ( .A(n4539), .Y(n4537) );
  NAND2X2 U1404 ( .A(n7894), .B(n7893), .Y(n7911) );
  NAND2X4 U1405 ( .A(n7863), .B(n7862), .Y(n7893) );
  XNOR2X4 U1406 ( .A(ICACHE_addr[23]), .B(n8706), .Y(n4417) );
  OAI2BB2X1 U1407 ( .B0(\i_MIPS/n167 ), .B1(n12), .A0N(n2160), .A1N(n8048), 
        .Y(\i_MIPS/N108 ) );
  CLKINVX1 U1408 ( .A(n8049), .Y(n8048) );
  NAND2BX1 U1409 ( .AN(n3576), .B(n8560), .Y(n7779) );
  AOI2BB1XL U1410 ( .A0N(n8065), .A1N(n8090), .B0(n8081), .Y(n8067) );
  OA22X1 U1411 ( .A0(n3548), .A1(n142), .B0(n3507), .B1(n1034), .Y(n4484) );
  NAND4X8 U1412 ( .A(n4435), .B(n4434), .C(n4433), .D(n4432), .Y(n8694) );
  AND2X2 U1413 ( .A(n8539), .B(n8540), .Y(n2812) );
  OAI221X2 U1414 ( .A0(n4589), .A1(n4599), .B0(n8538), .B1(n2815), .C0(n2838), 
        .Y(n4590) );
  INVX4 U1415 ( .A(n4590), .Y(n5977) );
  OA22X1 U1416 ( .A0(n3373), .A1(n1076), .B0(n3330), .B1(n161), .Y(n4490) );
  OAI222X2 U1417 ( .A0(n5105), .A1(n3219), .B0(n5104), .B1(n3216), .C0(n3654), 
        .C1(n3214), .Y(n7732) );
  OAI221X1 U1418 ( .A0(n6332), .A1(n6267), .B0(n3068), .B1(n6123), .C0(n5053), 
        .Y(n6919) );
  OAI221X4 U1419 ( .A0(\i_MIPS/n340 ), .A1(n3091), .B0(\i_MIPS/n341 ), .B1(
        n3087), .C0(n4811), .Y(n6267) );
  OA22X1 U1420 ( .A0(n6334), .A1(n5969), .B0(n6135), .B1(n3069), .Y(n5053) );
  AOI2BB1XL U1421 ( .A0N(n5900), .A1N(n3078), .B0(n2899), .Y(n4811) );
  XOR2X1 U1422 ( .A(n1071), .B(\D_cache/N49 ), .Y(n3044) );
  MXI2X4 U1423 ( .A(DCACHE_addr[1]), .B(DCACHE_rdata[3]), .S0(n4021), .Y(n8736) );
  OAI221X4 U1424 ( .A0(\D_cache/n164 ), .A1(n8867), .B0(n3074), .B1(n8848), 
        .C0(\D_cache/n174 ), .Y(DCACHE_rdata[3]) );
  INVX6 U1425 ( .A(n7989), .Y(n8256) );
  OAI221X4 U1426 ( .A0(\D_cache/n164 ), .A1(n8853), .B0(n3074), .B1(n8834), 
        .C0(\D_cache/n191 ), .Y(DCACHE_rdata[17]) );
  AO22X2 U1427 ( .A0(n2846), .A1(n3102), .B0(n3109), .B1(n5988), .Y(n5993) );
  NAND2X2 U1428 ( .A(n2799), .B(n2725), .Y(n2726) );
  INVX1 U1429 ( .A(n4019), .Y(n2725) );
  NAND4X4 U1430 ( .A(n6000), .B(n5999), .C(n5998), .D(n5997), .Y(n8164) );
  NOR4X4 U1431 ( .A(n5996), .B(n5995), .C(n6766), .D(n5994), .Y(n5997) );
  CLKMX2X4 U1432 ( .A(n5993), .B(n5992), .S0(n5991), .Y(n5994) );
  OAI221X1 U1433 ( .A0(n8763), .A1(n7044), .B0(n8750), .B1(n7043), .C0(n6799), 
        .Y(n6800) );
  NOR2X1 U1434 ( .A(\D_cache/n216 ), .B(\D_cache/n316 ), .Y(\D_cache/n455 ) );
  NAND2BX1 U1435 ( .AN(DCACHE_ren), .B(\D_cache/n204 ), .Y(\D_cache/n216 ) );
  NOR2X2 U1436 ( .A(n8808), .B(\D_cache/n520 ), .Y(\D_cache/n204 ) );
  NAND4X6 U1437 ( .A(n2771), .B(\D_cache/n525 ), .C(\D_cache/n526 ), .D(
        \D_cache/n527 ), .Y(\D_cache/n520 ) );
  NOR2X8 U1438 ( .A(n6458), .B(n6457), .Y(n6752) );
  NAND2X8 U1439 ( .A(n6456), .B(n6455), .Y(n6457) );
  AND3X8 U1440 ( .A(n2759), .B(n4595), .C(n5191), .Y(n2758) );
  AOI211X2 U1441 ( .A0(n9), .A1(n6389), .B0(n4824), .C0(n4599), .Y(n4600) );
  OA22X1 U1442 ( .A0(n8341), .A1(n3599), .B0(n2158), .B1(n8340), .Y(n8342) );
  OR2X8 U1443 ( .A(n8196), .B(n8195), .Y(n2000) );
  NAND2BX2 U1444 ( .AN(n3000), .B(n8621), .Y(n7329) );
  XOR2X4 U1445 ( .A(n7808), .B(n8037), .Y(n6122) );
  MXI2X2 U1446 ( .A(\i_MIPS/ID_EX[60] ), .B(\i_MIPS/ID_EX[92] ), .S0(n4018), 
        .Y(n4660) );
  AOI222X2 U1447 ( .A0(n2810), .A1(n6477), .B0(n6399), .B1(n6398), .C0(n6397), 
        .C1(n6396), .Y(n6411) );
  AND2X1 U1448 ( .A(n6614), .B(n6337), .Y(n2810) );
  XOR3XL U1449 ( .A(n7851), .B(n7853), .C(n7850), .Y(n7835) );
  AOI21XL U1450 ( .A0(n7919), .A1(n7952), .B0(n7918), .Y(n7921) );
  INVX1 U1451 ( .A(n7952), .Y(n7897) );
  OA22X1 U1452 ( .A0(n8388), .A1(n3599), .B0(n2158), .B1(n8387), .Y(n8389) );
  OA22X1 U1453 ( .A0(n7881), .A1(n3598), .B0(n2158), .B1(n7880), .Y(n7877) );
  OAI221X4 U1454 ( .A0(\i_MIPS/n351 ), .A1(n3091), .B0(\i_MIPS/n352 ), .B1(
        n3085), .C0(n5112), .Y(n5395) );
  CLKMX2X4 U1455 ( .A(n5395), .B(n5383), .S0(n4016), .Y(n6203) );
  NAND4BX4 U1456 ( .AN(n6481), .B(n6480), .C(n6479), .D(n6478), .Y(n8162) );
  AOI221X2 U1457 ( .A0(n6473), .A1(n6472), .B0(n6471), .B1(n6470), .C0(n6766), 
        .Y(n6479) );
  INVX3 U1458 ( .A(n4909), .Y(n4835) );
  NAND2X2 U1459 ( .A(n2819), .B(n2816), .Y(n4909) );
  AO21X4 U1460 ( .A0(n5473), .A1(n5472), .B0(n5471), .Y(n6062) );
  AO22X1 U1461 ( .A0(n5475), .A1(n3102), .B0(n3110), .B1(n6062), .Y(n5479) );
  NAND2X1 U1462 ( .A(\i_MIPS/ALUin1[16] ), .B(n52), .Y(n6914) );
  NAND2BX2 U1463 ( .AN(n3001), .B(n8589), .Y(n7327) );
  XNOR2X4 U1464 ( .A(n7829), .B(n7807), .Y(n5180) );
  NAND3X4 U1465 ( .A(n2705), .B(n2706), .C(n2707), .Y(n7807) );
  OAI222X4 U1466 ( .A0(n5035), .A1(n3166), .B0(n5013), .B1(n2761), .C0(n8740), 
        .C1(n3162), .Y(n7829) );
  CLKINVX1 U1467 ( .A(n8009), .Y(n5035) );
  XNOR2X4 U1468 ( .A(n8230), .B(n7784), .Y(n5450) );
  CLKMX2X4 U1469 ( .A(n6296), .B(n6295), .S0(n4012), .Y(n6297) );
  XNOR2X4 U1470 ( .A(n8214), .B(n8222), .Y(n6320) );
  NAND4X4 U1471 ( .A(n6857), .B(n6856), .C(n6855), .D(n6854), .Y(n8227) );
  AOI211X2 U1472 ( .A0(n6853), .A1(n6852), .B0(n6851), .C0(n6850), .Y(n6854)
         );
  NAND3X6 U1473 ( .A(n2744), .B(n2745), .C(n2746), .Y(n6851) );
  NAND2X2 U1474 ( .A(n4652), .B(\i_MIPS/n359 ), .Y(n6391) );
  OA22X1 U1475 ( .A0(n8373), .A1(n3599), .B0(n2158), .B1(n8372), .Y(n8374) );
  OAI222X2 U1476 ( .A0(n6256), .A1(n3166), .B0(n6234), .B1(n2761), .C0(n3020), 
        .C1(n3162), .Y(n7875) );
  INVX2 U1477 ( .A(n3027), .Y(n3020) );
  CLKINVX4 U1478 ( .A(n8244), .Y(n6256) );
  XOR3X4 U1479 ( .A(n3580), .B(n966), .C(n8326), .Y(n8328) );
  AOI222X4 U1480 ( .A0(n6990), .A1(n6760), .B0(n6832), .B1(n6759), .C0(n7006), 
        .C1(n6758), .Y(n6777) );
  INVX8 U1481 ( .A(n8167), .Y(n6823) );
  NAND2X1 U1482 ( .A(\i_MIPS/ALUin1[16] ), .B(n2154), .Y(n6909) );
  NAND2BX2 U1483 ( .AN(n2163), .B(n8651), .Y(n7414) );
  NAND2BX2 U1484 ( .AN(n3001), .B(n8587), .Y(n7411) );
  AOI2BB1X4 U1485 ( .A0N(n2859), .A1N(n8000), .B0(n7999), .Y(n8001) );
  OR2X1 U1486 ( .A(n8215), .B(n3049), .Y(n2033) );
  INVX12 U1487 ( .A(n5904), .Y(n6990) );
  XNOR2X4 U1488 ( .A(ICACHE_addr[10]), .B(n8693), .Y(n4450) );
  INVX3 U1489 ( .A(n5546), .Y(n4718) );
  CLKINVX6 U1490 ( .A(n8335), .Y(n8341) );
  OA22X4 U1491 ( .A0(n3305), .A1(n969), .B0(n3239), .B1(n80), .Y(n4519) );
  NAND3BX2 U1492 ( .AN(n4710), .B(n5049), .C(n4727), .Y(n4617) );
  XNOR2X4 U1493 ( .A(ICACHE_addr[9]), .B(n8692), .Y(n4449) );
  NAND4X8 U1494 ( .A(n4443), .B(n4442), .C(n4441), .D(n4440), .Y(n8692) );
  INVX4 U1495 ( .A(n8081), .Y(n8085) );
  OAI222X2 U1496 ( .A0(n6388), .A1(n3219), .B0(n6387), .B1(n3217), .C0(n8725), 
        .C1(n3214), .Y(n7812) );
  OAI222X4 U1497 ( .A0(n6388), .A1(n3166), .B0(n6366), .B1(n2761), .C0(n8725), 
        .C1(n3162), .Y(n7938) );
  INVX12 U1498 ( .A(n6136), .Y(n6614) );
  NAND3X2 U1499 ( .A(n1965), .B(n1966), .C(n1967), .Y(n7803) );
  AOI21X4 U1500 ( .A0(n5601), .A1(n8535), .B0(n4828), .Y(n2848) );
  AOI32X4 U1501 ( .A0(n2812), .A1(n6323), .A2(n5673), .B0(n2812), .B1(n5672), 
        .Y(n4825) );
  AO21X4 U1502 ( .A0(n5117), .A1(n5754), .B0(n5123), .Y(n5680) );
  NAND3BX4 U1503 ( .AN(n4901), .B(n4594), .C(n5322), .Y(n5191) );
  NAND3X6 U1504 ( .A(n15), .B(n4593), .C(n8491), .Y(n5322) );
  AOI222X4 U1505 ( .A0(n2811), .A1(n5265), .B0(n5264), .B1(n5263), .C0(n5262), 
        .C1(n5261), .Y(n5274) );
  MXI2X4 U1506 ( .A(DCACHE_rdata[11]), .B(DCACHE_addr[9]), .S0(\i_MIPS/n336 ), 
        .Y(n2795) );
  OAI222X2 U1507 ( .A0(n6454), .A1(n3219), .B0(n6453), .B1(n3217), .C0(n8726), 
        .C1(n3214), .Y(n7785) );
  NAND3BX4 U1508 ( .AN(n8090), .B(n8089), .C(n8088), .Y(n8186) );
  NAND2BX2 U1509 ( .AN(n3576), .B(n8561), .Y(n7756) );
  INVX4 U1510 ( .A(n7882), .Y(n7881) );
  NAND3X8 U1511 ( .A(n6322), .B(n6321), .C(n6320), .Y(n6458) );
  INVX8 U1512 ( .A(n3047), .Y(n7836) );
  NOR2BX2 U1513 ( .AN(n4022), .B(\D_cache/n165 ), .Y(n2868) );
  INVX3 U1514 ( .A(n8286), .Y(n8293) );
  NAND2X1 U1515 ( .A(n8685), .B(n8687), .Y(n8686) );
  XNOR2X4 U1516 ( .A(n8160), .B(n7801), .Y(n5181) );
  NAND2X1 U1517 ( .A(n3050), .B(n2158), .Y(n8259) );
  CLKBUFX3 U1518 ( .A(n3105), .Y(n3100) );
  CLKAND2X3 U1519 ( .A(n7966), .B(n7965), .Y(n2856) );
  INVX2 U1520 ( .A(n7967), .Y(n7966) );
  CLKBUFX2 U1521 ( .A(n3309), .Y(n3277) );
  NAND2X1 U1522 ( .A(n8336), .B(n8335), .Y(n2734) );
  AOI21X2 U1523 ( .A0(n8412), .A1(n8084), .B0(n8069), .Y(n8070) );
  NAND4X4 U1524 ( .A(n7410), .B(n7409), .C(n7408), .D(n7407), .Y(n7850) );
  NOR2X6 U1525 ( .A(n4431), .B(n4430), .Y(n4531) );
  NOR2X6 U1526 ( .A(n4527), .B(n4526), .Y(n4528) );
  XNOR2X4 U1527 ( .A(n7887), .B(n8011), .Y(n5452) );
  NAND4X8 U1528 ( .A(n4531), .B(n4530), .C(n4529), .D(n4528), .Y(n4539) );
  NAND4X4 U1529 ( .A(n8277), .B(n3615), .C(n7842), .D(n7841), .Y(n2772) );
  NOR4X4 U1530 ( .A(n6071), .B(n6070), .C(n6766), .D(n6069), .Y(n6072) );
  XNOR2X4 U1531 ( .A(\D_cache/N42 ), .B(DCACHE_addr[19]), .Y(\D_cache/n554 )
         );
  OAI222X2 U1532 ( .A0(n5379), .A1(n3218), .B0(n5378), .B1(n3216), .C0(n56), 
        .C1(n3215), .Y(n7784) );
  INVX16 U1533 ( .A(n2152), .Y(\D_cache/n164 ) );
  NOR2X8 U1534 ( .A(n4412), .B(n4411), .Y(n4418) );
  NAND3BX4 U1535 ( .AN(n3073), .B(n8278), .C(n8277), .Y(n8417) );
  BUFX20 U1536 ( .A(n8417), .Y(n3049) );
  NAND2X2 U1537 ( .A(n4680), .B(\i_MIPS/n368 ), .Y(n6552) );
  OR2X1 U1538 ( .A(n8357), .B(n3049), .Y(n1984) );
  OAI222X2 U1539 ( .A0(n5598), .A1(n3218), .B0(n5597), .B1(n3216), .C0(n8724), 
        .C1(n3215), .Y(n7811) );
  AND2X4 U1540 ( .A(n8259), .B(\i_MIPS/PC_o[1] ), .Y(n2720) );
  OAI222X2 U1541 ( .A0(n5533), .A1(n3218), .B0(n5532), .B1(n3216), .C0(n8739), 
        .C1(n3215), .Y(n8038) );
  OA22X4 U1542 ( .A0(n3275), .A1(n971), .B0(n3230), .B1(n82), .Y(n4396) );
  NAND4X4 U1543 ( .A(n7607), .B(n7606), .C(n7605), .D(n7604), .Y(n7932) );
  AOI21X4 U1544 ( .A0(n7945), .A1(n7944), .B0(n2858), .Y(n2861) );
  AOI221X2 U1545 ( .A0(n5608), .A1(n5607), .B0(n5606), .B1(n5605), .C0(n6766), 
        .Y(n5626) );
  NAND4X4 U1546 ( .A(n5452), .B(n5451), .C(n5450), .D(n5449), .Y(n5453) );
  NAND2X6 U1547 ( .A(n4912), .B(n2834), .Y(n7001) );
  AND4X4 U1548 ( .A(n4726), .B(n5048), .C(n4724), .D(n4727), .Y(n2834) );
  XNOR2X2 U1549 ( .A(ICACHE_addr[15]), .B(n8698), .Y(n4448) );
  OAI211X2 U1550 ( .A0(\i_MIPS/PC/n30 ), .A1(n12), .B0(n8281), .C0(n8280), .Y(
        \i_MIPS/PC/n62 ) );
  OA22X4 U1551 ( .A0(n8282), .A1(n18), .B0(n8276), .B1(n3050), .Y(n8281) );
  NAND2X4 U1552 ( .A(n8354), .B(n8352), .Y(n7864) );
  CLKINVX3 U1553 ( .A(n8328), .Y(n8327) );
  NAND3BX2 U1554 ( .AN(n20), .B(n7839), .C(n3610), .Y(n8421) );
  OAI221X1 U1555 ( .A0(n3107), .A1(n4974), .B0(n2852), .B1(n3099), .C0(n3097), 
        .Y(n4977) );
  XOR3X2 U1556 ( .A(n3580), .B(n8302), .C(n8304), .Y(n8296) );
  XOR2X4 U1557 ( .A(n7813), .B(n7976), .Y(n6973) );
  OAI222X4 U1558 ( .A0(n6971), .A1(n3219), .B0(n6949), .B1(n3216), .C0(n8728), 
        .C1(n3214), .Y(n7813) );
  NAND2X6 U1559 ( .A(n2832), .B(n2834), .Y(n6824) );
  NAND2BX4 U1560 ( .AN(\i_MIPS/ALU_Control/n10 ), .B(n4613), .Y(n4726) );
  CLKBUFX3 U1561 ( .A(n3104), .Y(n3103) );
  AO22XL U1562 ( .A0(n5323), .A1(n3103), .B0(n3111), .B1(n5386), .Y(n5325) );
  NAND2X6 U1563 ( .A(n4667), .B(\i_MIPS/n363 ), .Y(n6189) );
  OA22X2 U1564 ( .A0(n3305), .A1(n127), .B0(n3239), .B1(n1016), .Y(n4523) );
  OA22X2 U1565 ( .A0(n3549), .A1(n128), .B0(n3508), .B1(n1017), .Y(n4520) );
  NAND4X4 U1566 ( .A(n7781), .B(n7780), .C(n7779), .D(n7778), .Y(n7862) );
  NAND2X4 U1567 ( .A(n8188), .B(n8186), .Y(n8143) );
  OAI211X2 U1568 ( .A0(\i_MIPS/PC/n31 ), .A1(n13), .B0(n8298), .C0(n8297), .Y(
        \i_MIPS/PC/n63 ) );
  OA22X1 U1569 ( .A0(n8299), .A1(n18), .B0(n8296), .B1(n3050), .Y(n8298) );
  NAND4X4 U1570 ( .A(n7758), .B(n7757), .C(n7756), .D(n7755), .Y(n7882) );
  OA22XL U1571 ( .A0(n3549), .A1(n446), .B0(n3508), .B1(n1361), .Y(n4540) );
  OA22XL U1572 ( .A0(n3549), .A1(n534), .B0(n3508), .B1(n1453), .Y(n4544) );
  OA22XL U1573 ( .A0(n3549), .A1(n176), .B0(n3508), .B1(n1069), .Y(n4532) );
  OA22X2 U1574 ( .A0(n3549), .A1(n129), .B0(n3508), .B1(n1018), .Y(n4516) );
  INVX8 U1575 ( .A(n8279), .Y(n8330) );
  NAND3BX4 U1576 ( .AN(n8278), .B(n8277), .C(n3610), .Y(n8279) );
  OA22X1 U1577 ( .A0(n6202), .A1(n5752), .B0(n6056), .B1(n5680), .Y(n5687) );
  AOI221X2 U1578 ( .A0(n5679), .A1(n5678), .B0(n5677), .B1(n5676), .C0(n6766), 
        .Y(n5688) );
  AO22X1 U1579 ( .A0(n2822), .A1(n3102), .B0(n3110), .B1(n5735), .Y(n5679) );
  NOR2X8 U1580 ( .A(n5804), .B(n5805), .Y(n5806) );
  NAND4X4 U1581 ( .A(n5809), .B(n5806), .C(n5807), .D(n5808), .Y(n5885) );
  OAI221X2 U1582 ( .A0(n8085), .A1(n8087), .B0(n8091), .B1(n3577), .C0(n8084), 
        .Y(n8086) );
  XNOR2X4 U1583 ( .A(ICACHE_addr[24]), .B(n8707), .Y(n4493) );
  CLKINVX8 U1584 ( .A(n7009), .Y(n6682) );
  INVXL U1585 ( .A(n5752), .Y(n5757) );
  OA22X4 U1586 ( .A0(n8312), .A1(n18), .B0(n8309), .B1(n3050), .Y(n8311) );
  OAI221X4 U1587 ( .A0(\i_MIPS/n345 ), .A1(n3082), .B0(\i_MIPS/n346 ), .B1(
        n3077), .C0(n5114), .Y(n5481) );
  CLKMX2X8 U1588 ( .A(n5383), .B(n5481), .S0(n4016), .Y(n6464) );
  XOR2X4 U1589 ( .A(n7800), .B(n8226), .Y(n6749) );
  OAI222X4 U1590 ( .A0(n6747), .A1(n3219), .B0(n6725), .B1(n3217), .C0(n3022), 
        .C1(n3214), .Y(n7800) );
  NOR4X4 U1591 ( .A(n4734), .B(n4733), .C(n4732), .D(n4731), .Y(n4735) );
  OAI2BB1X4 U1592 ( .A0N(n4737), .A1N(n4736), .B0(n4735), .Y(n8314) );
  NOR3X2 U1593 ( .A(n1996), .B(n1997), .C(n1998), .Y(n8310) );
  AND2X4 U1594 ( .A(\i_MIPS/IF_ID[95] ), .B(n2157), .Y(n1996) );
  NAND3BX4 U1595 ( .AN(n19), .B(n4695), .C(n6257), .Y(n4696) );
  NAND2X4 U1596 ( .A(\i_MIPS/ALUin1[11] ), .B(n4661), .Y(n6258) );
  OAI221X4 U1597 ( .A0(n3106), .A1(n5735), .B0(n2822), .B1(n3098), .C0(n3097), 
        .Y(n5676) );
  XNOR2X4 U1598 ( .A(n8258), .B(n7732), .Y(n5179) );
  OAI221X2 U1599 ( .A0(n8239), .A1(n18), .B0(\i_MIPS/PC/n3 ), .B1(n8457), .C0(
        n8237), .Y(\i_MIPS/PC/n35 ) );
  NAND4X2 U1600 ( .A(n5062), .B(n5061), .C(n5060), .D(n5059), .Y(n8257) );
  NOR2X1 U1601 ( .A(n8224), .B(n18), .Y(n2022) );
  AO22XL U1602 ( .A0(n191), .A1(n228), .B0(n3207), .B1(n1348), .Y(n5094) );
  NAND4X1 U1603 ( .A(n7830), .B(n7787), .C(n7831), .D(\i_MIPS/IF_ID[64] ), .Y(
        n7792) );
  NAND2X4 U1604 ( .A(n2840), .B(n7820), .Y(n2733) );
  NAND4X8 U1605 ( .A(n4400), .B(n4399), .C(n4398), .D(n4397), .Y(n8702) );
  OA22X4 U1606 ( .A0(n3276), .A1(n972), .B0(n3230), .B1(n83), .Y(n4400) );
  CLKBUFX2 U1607 ( .A(n3309), .Y(n3276) );
  INVX4 U1608 ( .A(n2714), .Y(n2715) );
  NAND2BX1 U1609 ( .AN(n3576), .B(n8554), .Y(n7384) );
  NOR2X2 U1610 ( .A(n8049), .B(n3050), .Y(n2021) );
  XNOR2X4 U1611 ( .A(n8047), .B(n3577), .Y(n8049) );
  NAND2X4 U1612 ( .A(n8467), .B(n8468), .Y(n5192) );
  NAND2X2 U1613 ( .A(n2815), .B(n4825), .Y(n5732) );
  OAI222X2 U1614 ( .A0(n5671), .A1(n3164), .B0(n5649), .B1(n2761), .C0(n8717), 
        .C1(n3163), .Y(n8029) );
  OA22X4 U1615 ( .A0(n8329), .A1(n18), .B0(n8328), .B1(n3050), .Y(n8332) );
  NAND2X4 U1616 ( .A(n8124), .B(n3577), .Y(n8145) );
  OAI222X2 U1617 ( .A0(n5253), .A1(n3219), .B0(n5252), .B1(n3216), .C0(n8742), 
        .C1(n3214), .Y(n8011) );
  AO22X2 U1618 ( .A0(n6987), .A1(n3103), .B0(n3109), .B1(n6986), .Y(n7019) );
  OAI221X4 U1619 ( .A0(n7021), .A1(n8459), .B0(n7021), .B1(n8525), .C0(n7020), 
        .Y(n8300) );
  AOI211X1 U1620 ( .A0(n7019), .A1(n7018), .B0(n7017), .C0(n7016), .Y(n7020)
         );
  OAI211X2 U1621 ( .A0(n4598), .A1(n4597), .B0(n8481), .C0(n8482), .Y(n4821)
         );
  INVX3 U1622 ( .A(n6259), .Y(n4598) );
  BUFX12 U1623 ( .A(n8421), .Y(n3599) );
  AOI21X4 U1624 ( .A0(n8194), .A1(n8173), .B0(n8172), .Y(n8174) );
  OAI221X4 U1625 ( .A0(n7559), .A1(n2163), .B0(n7558), .B1(n3000), .C0(n7557), 
        .Y(n8324) );
  AO22X1 U1626 ( .A0(n2843), .A1(n3100), .B0(n3109), .B1(n4708), .Y(n4736) );
  INVX6 U1627 ( .A(n4726), .Y(n5049) );
  NAND2X4 U1628 ( .A(n8017), .B(n8018), .Y(n7979) );
  NAND3BX4 U1629 ( .AN(n7954), .B(n7953), .C(n7952), .Y(n8018) );
  XNOR2X4 U1630 ( .A(\D_cache/N43 ), .B(DCACHE_addr[18]), .Y(\D_cache/n555 )
         );
  NOR2X1 U1631 ( .A(n8264), .B(n18), .Y(n2736) );
  INVX16 U1632 ( .A(n3026), .Y(n7044) );
  AND2X8 U1633 ( .A(n2152), .B(n4022), .Y(n3026) );
  OR2X1 U1634 ( .A(n3106), .B(n6063), .Y(n1933) );
  OR2X1 U1635 ( .A(n2847), .B(n3098), .Y(n1934) );
  NAND3X2 U1636 ( .A(n1933), .B(n1934), .C(n3097), .Y(n6067) );
  AO21X4 U1637 ( .A0(n6062), .A1(n6061), .B0(n6060), .Y(n6063) );
  OR2X4 U1638 ( .A(n5105), .B(n3165), .Y(n1935) );
  OR2X2 U1639 ( .A(n5083), .B(n2761), .Y(n1936) );
  OR2X2 U1640 ( .A(n3654), .B(n3162), .Y(n1937) );
  OR2X1 U1641 ( .A(n3547), .B(n1055), .Y(n1938) );
  OR2XL U1642 ( .A(n3506), .B(n1066), .Y(n1939) );
  BUFX12 U1643 ( .A(n3574), .Y(n3547) );
  CLKBUFX4 U1644 ( .A(n3530), .Y(n3506) );
  OR2X1 U1645 ( .A(n3285), .B(n1056), .Y(n1940) );
  OR2X1 U1646 ( .A(n3237), .B(n1057), .Y(n1941) );
  AND2X2 U1647 ( .A(n1940), .B(n1941), .Y(n4475) );
  AND2XL U1648 ( .A(n5259), .B(n8470), .Y(n1942) );
  NOR2X2 U1649 ( .A(n1942), .B(n5258), .Y(n2849) );
  NAND2X4 U1650 ( .A(n4688), .B(\i_MIPS/n361 ), .Y(n8470) );
  INVXL U1651 ( .A(n8466), .Y(n5258) );
  AO22X4 U1652 ( .A0(n2849), .A1(n3103), .B0(n3111), .B1(n5260), .Y(n5262) );
  OR2X4 U1653 ( .A(n8743), .B(n3214), .Y(n1945) );
  INVX4 U1654 ( .A(n8162), .Y(n6526) );
  OR2XL U1655 ( .A(n3106), .B(n5386), .Y(n1946) );
  OR2X1 U1656 ( .A(n5323), .B(n3098), .Y(n1947) );
  NAND3X1 U1657 ( .A(n1946), .B(n1947), .C(n3097), .Y(n5326) );
  INVXL U1658 ( .A(n5388), .Y(n5323) );
  OR2X1 U1659 ( .A(n6615), .B(n6544), .Y(n1951) );
  OR2XL U1660 ( .A(n2796), .B(n6050), .Y(n1952) );
  OR2X1 U1661 ( .A(n6057), .B(n6136), .Y(n1953) );
  NAND3X2 U1662 ( .A(n1951), .B(n1952), .C(n1953), .Y(n5207) );
  MX2X1 U1663 ( .A(n5203), .B(n5202), .S0(n4016), .Y(n6615) );
  NOR2X1 U1664 ( .A(n3548), .B(n1031), .Y(n1954) );
  NOR2X1 U1665 ( .A(n3507), .B(n1032), .Y(n1955) );
  NOR2X1 U1666 ( .A(n1954), .B(n1955), .Y(n4500) );
  OR2X1 U1667 ( .A(n3547), .B(n1058), .Y(n1956) );
  OR2X1 U1668 ( .A(n3506), .B(n1059), .Y(n1957) );
  AND2X2 U1669 ( .A(n1956), .B(n1957), .Y(n4472) );
  OR2X1 U1670 ( .A(n3548), .B(n1060), .Y(n1958) );
  NAND2X2 U1671 ( .A(ICACHE_addr[28]), .B(n8711), .Y(n1961) );
  NAND2X8 U1672 ( .A(\i_MIPS/PC/n32 ), .B(n1960), .Y(n1962) );
  OR2X1 U1673 ( .A(n6613), .B(n6612), .Y(n1963) );
  OR2X1 U1674 ( .A(n6611), .B(n6610), .Y(n1964) );
  NAND2X6 U1675 ( .A(n6204), .B(n4016), .Y(n6612) );
  AOI211XL U1676 ( .A0(n6599), .A1(n8), .B0(n2898), .C0(n2984), .Y(n6611) );
  NAND2X6 U1677 ( .A(n6204), .B(n4017), .Y(n6610) );
  OR2X1 U1678 ( .A(n4890), .B(n3219), .Y(n1965) );
  OR2XL U1679 ( .A(n4868), .B(n3216), .Y(n1966) );
  OR2XL U1680 ( .A(n8744), .B(n3214), .Y(n1967) );
  MX2XL U1681 ( .A(n4865), .B(n4864), .S0(n4015), .Y(n4868) );
  XOR2X4 U1682 ( .A(n7803), .B(n8224), .Y(n5886) );
  OR2X4 U1683 ( .A(n3285), .B(n1013), .Y(n1968) );
  OR2X1 U1684 ( .A(n3237), .B(n1061), .Y(n1969) );
  OR2X1 U1685 ( .A(n3373), .B(n1062), .Y(n1970) );
  OR2X1 U1686 ( .A(n3330), .B(n1063), .Y(n1971) );
  CLKAND2X3 U1687 ( .A(n1970), .B(n1971), .Y(n4510) );
  NAND4X4 U1688 ( .A(n4511), .B(n4510), .C(n4509), .D(n4508), .Y(n8712) );
  NAND2X1 U1689 ( .A(n2075), .B(\i_MIPS/n336 ), .Y(n1972) );
  NAND2X2 U1690 ( .A(DCACHE_rdata[4]), .B(n4021), .Y(n1973) );
  INVX1 U1691 ( .A(n4029), .Y(n2075) );
  BUFX4 U1692 ( .A(\i_MIPS/EX_MEM_1 ), .Y(n4021) );
  NAND2X1 U1693 ( .A(n6768), .B(n6767), .Y(n1975) );
  AO22X1 U1694 ( .A0(n6764), .A1(n3101), .B0(n3108), .B1(n6765), .Y(n6770) );
  INVX12 U1695 ( .A(n7014), .Y(n6766) );
  NAND4BX4 U1696 ( .AN(n6778), .B(n6777), .C(n6776), .D(n6775), .Y(n8167) );
  OR2X2 U1697 ( .A(n8729), .B(n3162), .Y(n1976) );
  OR2X1 U1698 ( .A(n6297), .B(n2761), .Y(n1978) );
  CLKINVX8 U1699 ( .A(n7786), .Y(n6319) );
  OR2X1 U1700 ( .A(n3286), .B(n1064), .Y(n1979) );
  OR2X1 U1701 ( .A(n3238), .B(n1065), .Y(n1980) );
  AND2X2 U1702 ( .A(n1979), .B(n1980), .Y(n4511) );
  NAND2X8 U1703 ( .A(n1982), .B(n1983), .Y(n4512) );
  NAND4X6 U1704 ( .A(n4515), .B(n4514), .C(n4513), .D(n4512), .Y(n4527) );
  OR2XL U1705 ( .A(n8356), .B(n18), .Y(n1985) );
  OR2XL U1706 ( .A(\i_MIPS/PC/n8 ), .B(n13), .Y(n1986) );
  NAND3X2 U1707 ( .A(n1984), .B(n1985), .C(n1986), .Y(n8362) );
  XOR3XL U1708 ( .A(n8354), .B(n8353), .C(n8352), .Y(n8357) );
  OR2XL U1709 ( .A(n8385), .B(n18), .Y(n1988) );
  OR2X1 U1710 ( .A(\i_MIPS/PC/n6 ), .B(n13), .Y(n1989) );
  NAND3X2 U1711 ( .A(n1987), .B(n1988), .C(n1989), .Y(n8391) );
  INVXL U1712 ( .A(n8230), .Y(n8385) );
  OR2XL U1713 ( .A(n8338), .B(n17), .Y(n1991) );
  OR2X1 U1714 ( .A(\i_MIPS/PC/n5 ), .B(n3615), .Y(n1992) );
  OR2XL U1715 ( .A(n8370), .B(n18), .Y(n1994) );
  OR2X1 U1716 ( .A(\i_MIPS/PC/n7 ), .B(n3612), .Y(n1995) );
  NAND3X2 U1717 ( .A(n1993), .B(n1994), .C(n1995), .Y(n8376) );
  AND2XL U1718 ( .A(n8325), .B(n8330), .Y(n1997) );
  AND2XL U1719 ( .A(\i_MIPS/IF_ID_30 ), .B(n3597), .Y(n1998) );
  OAI211X2 U1720 ( .A0(\i_MIPS/PC/n32 ), .A1(n3613), .B0(n8311), .C0(n8310), 
        .Y(\i_MIPS/PC/n64 ) );
  CLKINVX1 U1721 ( .A(n2860), .Y(n2002) );
  NAND2X4 U1722 ( .A(n2001), .B(n2002), .Y(n8192) );
  BUFX20 U1723 ( .A(n3581), .Y(n3580) );
  XOR2X4 U1724 ( .A(n8121), .B(ICACHE_addr[22]), .Y(n8146) );
  OR2XL U1725 ( .A(n8030), .B(n3049), .Y(n2003) );
  OR2XL U1726 ( .A(n8036), .B(n18), .Y(n2004) );
  OR2X1 U1727 ( .A(\i_MIPS/PC/n21 ), .B(n3612), .Y(n2005) );
  NAND3X2 U1728 ( .A(n2003), .B(n2004), .C(n2005), .Y(n8035) );
  XOR3X1 U1729 ( .A(n3580), .B(n8043), .C(n8045), .Y(n8030) );
  OR2X1 U1730 ( .A(n8152), .B(n3049), .Y(n2006) );
  OR2XL U1731 ( .A(n8158), .B(n18), .Y(n2007) );
  OR2X1 U1732 ( .A(\i_MIPS/PC/n27 ), .B(n3610), .Y(n2008) );
  NAND3X2 U1733 ( .A(n2006), .B(n2007), .C(n2008), .Y(n8157) );
  XOR3X1 U1734 ( .A(n3580), .B(n8171), .C(n8173), .Y(n8152) );
  OR2XL U1735 ( .A(n8256), .B(n18), .Y(n2010) );
  OR2X1 U1736 ( .A(\i_MIPS/PC/n19 ), .B(n3615), .Y(n2011) );
  NAND3X2 U1737 ( .A(n2009), .B(n2010), .C(n2011), .Y(n7993) );
  OR2X1 U1738 ( .A(n8418), .B(n3050), .Y(n2012) );
  OR2X1 U1739 ( .A(\i_MIPS/PC/n23 ), .B(n3611), .Y(n2014) );
  NAND3X2 U1740 ( .A(n2012), .B(n2013), .C(n2014), .Y(n8425) );
  XOR3X2 U1741 ( .A(n8413), .B(n3579), .C(n8412), .Y(n8418) );
  OR2X1 U1742 ( .A(n8129), .B(n3049), .Y(n2015) );
  OR2XL U1743 ( .A(n8128), .B(n18), .Y(n2016) );
  OR2X1 U1744 ( .A(\i_MIPS/PC/n26 ), .B(n13), .Y(n2017) );
  NAND3X2 U1745 ( .A(n2015), .B(n2016), .C(n2017), .Y(n8141) );
  INVXL U1746 ( .A(n7808), .Y(n8128) );
  OR2X1 U1747 ( .A(n8093), .B(n3049), .Y(n2018) );
  OR2XL U1748 ( .A(n8228), .B(n18), .Y(n2019) );
  OR2X1 U1749 ( .A(\i_MIPS/PC/n25 ), .B(n3614), .Y(n2020) );
  NAND3X2 U1750 ( .A(n2018), .B(n2019), .C(n2020), .Y(n8098) );
  XOR3X1 U1751 ( .A(n3579), .B(n8124), .C(n8123), .Y(n8093) );
  INVX6 U1752 ( .A(n6903), .Y(n8228) );
  NOR2XL U1753 ( .A(\i_MIPS/PC/n22 ), .B(n3611), .Y(n2023) );
  OR3X2 U1754 ( .A(n2021), .B(n2022), .C(n2023), .Y(n8055) );
  OR2XL U1755 ( .A(n7888), .B(n3049), .Y(n2024) );
  OR2XL U1756 ( .A(n8013), .B(n18), .Y(n2025) );
  OR2X1 U1757 ( .A(\i_MIPS/PC/n12 ), .B(n3614), .Y(n2026) );
  NAND3X2 U1758 ( .A(n2024), .B(n2025), .C(n2026), .Y(n7891) );
  OR2XL U1759 ( .A(n7924), .B(n3049), .Y(n2027) );
  OR2XL U1760 ( .A(n8250), .B(n18), .Y(n2028) );
  OR2X1 U1761 ( .A(\i_MIPS/PC/n15 ), .B(n12), .Y(n2029) );
  NAND3X2 U1762 ( .A(n2027), .B(n2028), .C(n2029), .Y(n7927) );
  XOR3X2 U1763 ( .A(n7933), .B(n7935), .C(n7932), .Y(n7924) );
  INVXL U1764 ( .A(n7923), .Y(n8250) );
  OR2XL U1765 ( .A(n7876), .B(n3049), .Y(n2030) );
  OR2XL U1766 ( .A(n8245), .B(n18), .Y(n2031) );
  OR2X1 U1767 ( .A(\i_MIPS/PC/n11 ), .B(n3614), .Y(n2032) );
  NAND3X2 U1768 ( .A(n2030), .B(n2031), .C(n2032), .Y(n7879) );
  OR2XL U1769 ( .A(n8248), .B(n17), .Y(n2034) );
  OR2X1 U1770 ( .A(\i_MIPS/PC/n14 ), .B(n3615), .Y(n2035) );
  XOR3X2 U1771 ( .A(n8221), .B(n8212), .C(n8211), .Y(n8215) );
  OR2X1 U1772 ( .A(n8073), .B(n3049), .Y(n2036) );
  OR2XL U1773 ( .A(n8226), .B(n18), .Y(n2037) );
  OR2X1 U1774 ( .A(\i_MIPS/PC/n24 ), .B(n8457), .Y(n2038) );
  NAND3X2 U1775 ( .A(n2036), .B(n2037), .C(n2038), .Y(n8079) );
  OR2XL U1776 ( .A(n8010), .B(n17), .Y(n2040) );
  OR2X1 U1777 ( .A(\i_MIPS/PC/n9 ), .B(n3614), .Y(n2041) );
  OR2XL U1778 ( .A(n7904), .B(n3049), .Y(n2042) );
  OR2XL U1779 ( .A(n8247), .B(n18), .Y(n2043) );
  OR2X1 U1780 ( .A(\i_MIPS/PC/n13 ), .B(n8457), .Y(n2044) );
  NAND3X2 U1781 ( .A(n2042), .B(n2043), .C(n2044), .Y(n7907) );
  INVXL U1782 ( .A(n7903), .Y(n8247) );
  OR2XL U1783 ( .A(n7939), .B(n3049), .Y(n2045) );
  OR2XL U1784 ( .A(n8252), .B(n18), .Y(n2046) );
  OR2X1 U1785 ( .A(\i_MIPS/PC/n16 ), .B(n3613), .Y(n2047) );
  NAND3X2 U1786 ( .A(n2045), .B(n2046), .C(n2047), .Y(n7942) );
  XOR3X2 U1787 ( .A(n7956), .B(n7936), .C(n7955), .Y(n7939) );
  OR2X1 U1788 ( .A(n8200), .B(n3049), .Y(n2048) );
  OR2XL U1789 ( .A(n8458), .B(n18), .Y(n2049) );
  OR2X1 U1790 ( .A(\i_MIPS/PC/n29 ), .B(n3610), .Y(n2050) );
  NAND3X2 U1791 ( .A(n2048), .B(n2049), .C(n2050), .Y(n8205) );
  OR2XL U1792 ( .A(n7857), .B(n3049), .Y(n2051) );
  OR2XL U1793 ( .A(n8232), .B(n18), .Y(n2052) );
  OR2X1 U1794 ( .A(\i_MIPS/PC/n10 ), .B(n3615), .Y(n2053) );
  NAND3X2 U1795 ( .A(n2051), .B(n2052), .C(n2053), .Y(n7860) );
  INVXL U1796 ( .A(n7856), .Y(n8232) );
  OR2XL U1797 ( .A(n7972), .B(n3050), .Y(n2054) );
  OR2XL U1798 ( .A(n7976), .B(n18), .Y(n2055) );
  OR2XL U1799 ( .A(\i_MIPS/PC/n18 ), .B(n8457), .Y(n2056) );
  NAND3X2 U1800 ( .A(n2054), .B(n2055), .C(n2056), .Y(n7975) );
  XOR3X2 U1801 ( .A(n7986), .B(n7970), .C(n7985), .Y(n7972) );
  BUFX12 U1802 ( .A(n8417), .Y(n3050) );
  OAI222X4 U1803 ( .A0(n2796), .A1(n6756), .B0(n6549), .B1(n6201), .C0(n6551), 
        .C1(n6544), .Y(n5272) );
  AOI21X1 U1804 ( .A0(n6059), .A1(n8522), .B0(n6058), .Y(n2847) );
  OR4X2 U1805 ( .A(n5047), .B(n5674), .C(n8923), .D(n8924), .Y(n5051) );
  OAI22X1 U1806 ( .A0(n8921), .A1(n8920), .B0(n8716), .B1(n8921), .Y(n8922) );
  OAI221X4 U1807 ( .A0(n3068), .A1(n6267), .B0(n3069), .B1(n5969), .C0(n5964), 
        .Y(n6124) );
  CLKMX2X2 U1808 ( .A(n5969), .B(n6267), .S0(n4016), .Y(n5971) );
  CLKMX2X4 U1809 ( .A(n6123), .B(n5969), .S0(n4016), .Y(n5319) );
  OAI221X4 U1810 ( .A0(\i_MIPS/n346 ), .A1(n14), .B0(\i_MIPS/n347 ), .B1(n3077), .C0(n4813), .Y(n5969) );
  XNOR2X4 U1811 ( .A(n7875), .B(n7805), .Y(n6321) );
  OAI222X4 U1812 ( .A0(n6256), .A1(n3218), .B0(n6255), .B1(n3217), .C0(n3020), 
        .C1(n3214), .Y(n7805) );
  XNOR2X4 U1813 ( .A(n7856), .B(n7806), .Y(n6322) );
  OAI222X4 U1814 ( .A0(n6187), .A1(n3166), .B0(n6165), .B1(n2761), .C0(n3162), 
        .C1(n8745), .Y(n7856) );
  XNOR2X4 U1815 ( .A(n7938), .B(n7812), .Y(n6456) );
  NAND3BX2 U1816 ( .AN(n10), .B(n4388), .C(\i_MIPS/PC/n8 ), .Y(n2797) );
  OAI2BB1X4 U1817 ( .A0N(n5539), .A1N(n5549), .B0(n5545), .Y(n5675) );
  XNOR2X4 U1818 ( .A(ICACHE_addr[12]), .B(n8695), .Y(n4483) );
  XNOR2X4 U1819 ( .A(ICACHE_addr[13]), .B(n8696), .Y(n4481) );
  INVX8 U1820 ( .A(n6544), .Y(n6204) );
  NAND4BX2 U1821 ( .AN(n5488), .B(n5487), .C(n5486), .D(n5485), .Y(n8039) );
  AOI222X4 U1822 ( .A0(n5468), .A1(n6990), .B0(n6774), .B1(n6206), .C0(n5467), 
        .C1(n7006), .Y(n5487) );
  XNOR2X4 U1823 ( .A(n8029), .B(n8014), .Y(n5807) );
  AND2X4 U1824 ( .A(n3084), .B(\i_MIPS/ALUin1[17] ), .Y(n2905) );
  OAI222X4 U1825 ( .A0(n8003), .A1(n3049), .B0(n1086), .B1(n18), .C0(
        \i_MIPS/PC/n20 ), .C1(n3610), .Y(n8008) );
  XNOR2X4 U1826 ( .A(\D_cache/N46 ), .B(DCACHE_addr[15]), .Y(\D_cache/n532 )
         );
  CLKMX2X2 U1827 ( .A(n3072), .B(n2865), .S0(n5256), .Y(n5206) );
  CLKMX2X2 U1828 ( .A(n3072), .B(n2865), .S0(n6404), .Y(n6406) );
  CLKMX2X2 U1829 ( .A(n3072), .B(n2865), .S0(n4972), .Y(n4917) );
  BUFX12 U1830 ( .A(n6405), .Y(n3072) );
  XOR2X4 U1831 ( .A(n8272), .B(n8286), .Y(n8273) );
  NAND2X4 U1832 ( .A(n6680), .B(n4017), .Y(n6201) );
  AOI22XL U1833 ( .A0(\D_cache/N135 ), .A1(n2153), .B0(n3032), .B1(
        \D_cache/N167 ), .Y(\D_cache/n191 ) );
  OAI211X2 U1834 ( .A0(\i_MIPS/PC/n33 ), .A1(n3612), .B0(n8332), .C0(n8331), 
        .Y(\i_MIPS/PC/n65 ) );
  OAI222X2 U1835 ( .A0(n6187), .A1(n3218), .B0(n6186), .B1(n3217), .C0(n3215), 
        .C1(n8745), .Y(n7806) );
  OAI222X2 U1836 ( .A0(n5379), .A1(n3164), .B0(n5357), .B1(n2761), .C0(n56), 
        .C1(n3163), .Y(n8230) );
  INVXL U1837 ( .A(n2076), .Y(n2057) );
  INVXL U1838 ( .A(n2066), .Y(n2058) );
  INVXL U1839 ( .A(n2141), .Y(n2059) );
  INVXL U1840 ( .A(n2065), .Y(n2060) );
  CLKINVX1 U1841 ( .A(n4030), .Y(n2061) );
  CLKINVX1 U1842 ( .A(n4030), .Y(n2062) );
  CLKINVX1 U1843 ( .A(n4030), .Y(n2063) );
  CLKINVX1 U1844 ( .A(n4030), .Y(n2064) );
  CLKINVX1 U1845 ( .A(n4030), .Y(n2065) );
  CLKINVX1 U1846 ( .A(n4030), .Y(n2066) );
  CLKINVX1 U1847 ( .A(n4030), .Y(n2067) );
  CLKINVX1 U1848 ( .A(n4030), .Y(n2068) );
  CLKINVX1 U1849 ( .A(n4029), .Y(n2069) );
  CLKINVX1 U1850 ( .A(n4029), .Y(n2070) );
  CLKINVX1 U1851 ( .A(n4029), .Y(n2071) );
  CLKINVX1 U1852 ( .A(n4029), .Y(n2072) );
  CLKINVX1 U1853 ( .A(n4029), .Y(n2073) );
  CLKINVX1 U1854 ( .A(n4029), .Y(n2074) );
  CLKINVX1 U1855 ( .A(n4029), .Y(n2076) );
  CLKINVX1 U1856 ( .A(n3056), .Y(n2077) );
  CLKINVX1 U1857 ( .A(n3056), .Y(n2078) );
  CLKINVX1 U1858 ( .A(n3056), .Y(n2079) );
  INVX1 U1859 ( .A(n3056), .Y(n2080) );
  CLKINVX1 U1860 ( .A(n3056), .Y(n2081) );
  CLKINVX1 U1861 ( .A(n3056), .Y(n2082) );
  CLKINVX1 U1862 ( .A(n3056), .Y(n2083) );
  CLKINVX1 U1863 ( .A(n3056), .Y(n2084) );
  CLKINVX1 U1864 ( .A(n4026), .Y(n2085) );
  CLKINVX1 U1865 ( .A(n4026), .Y(n2086) );
  INVX1 U1866 ( .A(n4026), .Y(n2087) );
  INVX1 U1867 ( .A(n4026), .Y(n2088) );
  CLKINVX1 U1868 ( .A(n4026), .Y(n2089) );
  CLKINVX1 U1869 ( .A(n4026), .Y(n2090) );
  CLKINVX1 U1870 ( .A(n4026), .Y(n2091) );
  CLKINVX1 U1871 ( .A(n4026), .Y(n2092) );
  CLKINVX1 U1872 ( .A(n4027), .Y(n2093) );
  CLKINVX1 U1873 ( .A(n4027), .Y(n2094) );
  INVX1 U1874 ( .A(n4027), .Y(n2095) );
  CLKINVX1 U1875 ( .A(n4027), .Y(n2096) );
  CLKINVX1 U1876 ( .A(n4027), .Y(n2098) );
  CLKINVX1 U1877 ( .A(n4027), .Y(n2099) );
  CLKINVX1 U1878 ( .A(n4027), .Y(n2100) );
  CLKINVX1 U1879 ( .A(n4028), .Y(n2101) );
  CLKINVX1 U1880 ( .A(n4028), .Y(n2102) );
  INVX1 U1881 ( .A(n4028), .Y(n2103) );
  CLKINVX1 U1882 ( .A(n4028), .Y(n2104) );
  CLKINVX1 U1883 ( .A(n4028), .Y(n2106) );
  CLKINVX1 U1884 ( .A(n4028), .Y(n2107) );
  CLKINVX1 U1885 ( .A(n4028), .Y(n2108) );
  INVX16 U1886 ( .A(n3056), .Y(DCACHE_addr[2]) );
  INVX3 U1887 ( .A(n3056), .Y(n2111) );
  INVX4 U1888 ( .A(n3057), .Y(n2126) );
  INVX4 U1889 ( .A(n3057), .Y(n2127) );
  INVX4 U1890 ( .A(n3057), .Y(n2130) );
  CLKBUFX2 U1891 ( .A(n2750), .Y(n2137) );
  CLKBUFX2 U1892 ( .A(n2750), .Y(n2138) );
  CLKBUFX2 U1893 ( .A(n2750), .Y(n2139) );
  CLKBUFX2 U1894 ( .A(n2750), .Y(n2140) );
  CLKBUFX2 U1895 ( .A(n2750), .Y(n2141) );
  CLKBUFX2 U1896 ( .A(n2750), .Y(n2142) );
  CLKBUFX2 U1897 ( .A(n2750), .Y(n2143) );
  CLKBUFX2 U1898 ( .A(n2750), .Y(n2144) );
  INVX8 U1899 ( .A(n4026), .Y(n4024) );
  INVX20 U1900 ( .A(n2750), .Y(n4030) );
  BUFX12 U1901 ( .A(n4030), .Y(n4029) );
  BUFX6 U1902 ( .A(n4030), .Y(n4026) );
  CLKBUFX6 U1903 ( .A(n4030), .Y(n4028) );
  INVX12 U1904 ( .A(n4025), .Y(n3057) );
  AO21X4 U1905 ( .A0(n5889), .A1(n8530), .B0(n8460), .Y(n5810) );
  OAI2BB1X2 U1906 ( .A0N(n6761), .A1N(n8518), .B0(n8520), .Y(n5889) );
  INVX4 U1907 ( .A(n3597), .Y(n3594) );
  INVX8 U1908 ( .A(n6550), .Y(n6617) );
  NOR2X2 U1909 ( .A(n3076), .B(n5482), .Y(n6205) );
  OAI221X4 U1910 ( .A0(n2796), .A1(n6546), .B0(n6545), .B1(n6544), .C0(n6543), 
        .Y(n6554) );
  AOI211X2 U1911 ( .A0(n6924), .A1(n6923), .B0(n6922), .C0(n6921), .Y(n6925)
         );
  AO22X4 U1912 ( .A0(n6917), .A1(n6993), .B0(n6916), .B1(n6915), .Y(n6922) );
  AOI221X1 U1913 ( .A0(n8476), .A1(n8475), .B0(n8474), .B1(n8473), .C0(n8472), 
        .Y(n8489) );
  NAND2X2 U1914 ( .A(\i_MIPS/ALUin1[11] ), .B(n2145), .Y(n8473) );
  OR2X4 U1915 ( .A(n5803), .B(n3218), .Y(n2754) );
  NAND2BX4 U1916 ( .AN(n5189), .B(n6194), .Y(n5257) );
  NAND2X2 U1917 ( .A(\i_MIPS/ALUin1[9] ), .B(n4689), .Y(n6194) );
  XOR2X2 U1918 ( .A(n8151), .B(n8038), .Y(n5600) );
  AOI2BB1X1 U1919 ( .A0N(\i_MIPS/ALUin1[14] ), .A1N(n3078), .B0(n2844), .Y(
        n4913) );
  NAND2XL U1920 ( .A(\i_MIPS/ALUin1[14] ), .B(n4654), .Y(n8478) );
  OA21X1 U1921 ( .A0(\i_MIPS/ALUin1[18] ), .A1(n3086), .B0(n4914), .Y(n4814)
         );
  XNOR2X4 U1922 ( .A(n2765), .B(n8318), .Y(n8306) );
  AOI211X2 U1923 ( .A0(n5402), .A1(n6529), .B0(n4989), .C0(n4988), .Y(n4990)
         );
  XNOR2X4 U1924 ( .A(n8273), .B(n3577), .Y(n8276) );
  NOR4X2 U1925 ( .A(n6700), .B(n6699), .C(n6766), .D(n6698), .Y(n6701) );
  OAI221X4 U1926 ( .A0(n6334), .A1(n6267), .B0(n3076), .B1(n5319), .C0(n5614), 
        .Y(n5331) );
  XNOR2X4 U1927 ( .A(ICACHE_addr[5]), .B(n8688), .Y(n4525) );
  XNOR2X4 U1928 ( .A(ICACHE_addr[25]), .B(n8708), .Y(n4480) );
  OAI221X4 U1929 ( .A0(n3107), .A1(n5257), .B0(n5196), .B1(n3098), .C0(n3097), 
        .Y(n5199) );
  XNOR2X4 U1930 ( .A(ICACHE_addr[14]), .B(n8697), .Y(n4482) );
  NAND4X4 U1931 ( .A(n4499), .B(n4498), .C(n4497), .D(n4496), .Y(n8704) );
  OA22X2 U1932 ( .A0(n3548), .A1(n130), .B0(n3507), .B1(n1019), .Y(n4496) );
  OA22X4 U1933 ( .A0(n3372), .A1(n1073), .B0(n3329), .B1(n84), .Y(n4454) );
  NAND2X6 U1934 ( .A(n4493), .B(n4492), .Y(n4494) );
  XNOR2X4 U1935 ( .A(ICACHE_addr[26]), .B(n8709), .Y(n4492) );
  NAND4X4 U1936 ( .A(n4503), .B(n4502), .C(n4501), .D(n4500), .Y(n8699) );
  XNOR2X4 U1937 ( .A(ICACHE_addr[21]), .B(n8704), .Y(n4515) );
  AOI222X1 U1938 ( .A0(n6465), .A1(n6990), .B0(n6832), .B1(n6464), .C0(n6830), 
        .C1(n6463), .Y(n6480) );
  AOI222X1 U1939 ( .A0(n6833), .A1(n6990), .B0(n6832), .B1(n6831), .C0(n6830), 
        .C1(n6829), .Y(n6855) );
  CLKINVX1 U1940 ( .A(n6201), .Y(n6830) );
  OAI222X4 U1941 ( .A0(n2796), .A1(n6828), .B0(n6612), .B1(n5269), .C0(n6550), 
        .C1(n5547), .Y(n4989) );
  XOR3X2 U1942 ( .A(n8026), .B(n8001), .C(n3577), .Y(n8003) );
  XNOR2X4 U1943 ( .A(n7923), .B(n7785), .Y(n6455) );
  XNOR2X4 U1944 ( .A(n7903), .B(n7804), .Y(n5451) );
  NAND2X4 U1945 ( .A(\i_MIPS/ALUin1[4] ), .B(n4669), .Y(n8499) );
  OA22X1 U1946 ( .A0(\i_MIPS/ALUin1[5] ), .A1(n14), .B0(\i_MIPS/ALUin1[4] ), 
        .B1(n3078), .Y(n5038) );
  NAND2X6 U1947 ( .A(\i_MIPS/ALUin1[4] ), .B(n4678), .Y(n5384) );
  INVXL U1948 ( .A(n3064), .Y(n2148) );
  INVXL U1949 ( .A(n3067), .Y(n2149) );
  INVXL U1950 ( .A(n3063), .Y(n2151) );
  INVXL U1951 ( .A(n6688), .Y(n6469) );
  AOI2BB1X4 U1952 ( .A0N(n5537), .A1N(n5536), .B0(n5535), .Y(n5538) );
  INVX6 U1953 ( .A(n2796), .Y(n6618) );
  OAI222X4 U1954 ( .A0(n2796), .A1(n6462), .B0(n6612), .B1(n5397), .C0(n2831), 
        .C1(n6550), .Y(n5400) );
  NAND2X4 U1955 ( .A(n8492), .B(n8499), .Y(n4901) );
  XOR2X1 U1956 ( .A(n7608), .B(\i_MIPS/IR_ID[21] ), .Y(n4742) );
  XOR2X1 U1957 ( .A(n7608), .B(\i_MIPS/IR_ID[16] ), .Y(n4781) );
  OAI33X1 U1958 ( .A0(n3098), .A1(n5833), .A2(n2876), .B0(n3106), .B1(n2876), 
        .B2(n5811), .Y(n5838) );
  INVX1 U1959 ( .A(n5810), .Y(n5833) );
  NAND2X6 U1960 ( .A(\i_MIPS/ALUin1[5] ), .B(n4670), .Y(n8498) );
  NAND2X6 U1961 ( .A(\i_MIPS/ALUin1[5] ), .B(n4671), .Y(n5390) );
  AOI2BB1XL U1962 ( .A0N(n2728), .A1N(\i_MIPS/n371 ), .B0(n2839), .Y(n5044) );
  OAI222X4 U1963 ( .A0(n5177), .A1(n3164), .B0(n5155), .B1(n2761), .C0(n8732), 
        .C1(n3162), .Y(n8236) );
  BUFX6 U1964 ( .A(n3033), .Y(n2152) );
  OA22X4 U1965 ( .A0(n3547), .A1(n973), .B0(n3506), .B1(n85), .Y(n4456) );
  NAND4X4 U1966 ( .A(n4507), .B(n4506), .C(n4505), .D(n4504), .Y(n8700) );
  XNOR2X4 U1967 ( .A(ICACHE_addr[16]), .B(n8699), .Y(n4514) );
  NAND2X1 U1968 ( .A(\i_MIPS/ID_EX[73] ), .B(n4019), .Y(n2727) );
  NAND4X4 U1969 ( .A(n4483), .B(n4482), .C(n4481), .D(n4480), .Y(n4495) );
  XNOR2X4 U1970 ( .A(ICACHE_addr[17]), .B(n8700), .Y(n4513) );
  OAI222X4 U1971 ( .A0(n6120), .A1(n3166), .B0(n6098), .B1(n2761), .C0(n8737), 
        .C1(n3162), .Y(n8177) );
  XOR2X4 U1972 ( .A(n8234), .B(n7734), .Y(n6670) );
  OAI222X4 U1973 ( .A0(n6669), .A1(n3166), .B0(n6647), .B1(n2761), .C0(n8733), 
        .C1(n3162), .Y(n8234) );
  NAND2X2 U1974 ( .A(n4461), .B(n4460), .Y(n4462) );
  XNOR2X2 U1975 ( .A(ICACHE_addr[27]), .B(n8710), .Y(n4460) );
  BUFX20 U1976 ( .A(n968), .Y(n2153) );
  AO22X4 U1977 ( .A0(n8325), .A1(n3577), .B0(n8323), .B1(n8322), .Y(n8326) );
  NOR4X4 U1978 ( .A(\i_MIPS/n329 ), .B(\i_MIPS/ID_EX[110] ), .C(
        \i_MIPS/ID_EX[109] ), .D(n1083), .Y(\i_MIPS/ALU_Control/n11 ) );
  OAI221X4 U1979 ( .A0(n8771), .A1(n7044), .B0(n8758), .B1(n7043), .C0(n5647), 
        .Y(n5648) );
  OAI222X4 U1980 ( .A0(n5177), .A1(n3219), .B0(n5176), .B1(n3216), .C0(n8732), 
        .C1(n3214), .Y(n7733) );
  XNOR2X4 U1981 ( .A(n8306), .B(n3577), .Y(n8309) );
  OAI221X4 U1982 ( .A0(n3106), .A1(n6692), .B0(n2853), .B1(n3098), .C0(n3096), 
        .Y(n6696) );
  NAND2X2 U1983 ( .A(n11), .B(\i_MIPS/n362 ), .Y(n6207) );
  MXI2X2 U1984 ( .A(\i_MIPS/ID_EX[50] ), .B(n3076), .S0(n4019), .Y(n4668) );
  AOI21X2 U1985 ( .A0(n5824), .A1(n5754), .B0(n5123), .Y(n2818) );
  INVX4 U1986 ( .A(n4670), .Y(n4671) );
  OAI221X1 U1987 ( .A0(\D_cache/n164 ), .A1(n8860), .B0(n3074), .B1(n8841), 
        .C0(\D_cache/n198 ), .Y(DCACHE_rdata[10]) );
  OAI221X2 U1988 ( .A0(\D_cache/n164 ), .A1(n8869), .B0(n3074), .B1(n8850), 
        .C0(\D_cache/n188 ), .Y(DCACHE_rdata[1]) );
  AOI21X1 U1989 ( .A0(n6910), .A1(n8539), .B0(n5674), .Y(n2822) );
  NAND4X4 U1990 ( .A(n5626), .B(n5625), .C(n5624), .D(n5623), .Y(n8015) );
  OAI222X2 U1991 ( .A0(n6971), .A1(n3166), .B0(n6970), .B1(n2761), .C0(n8728), 
        .C1(n3162), .Y(n6972) );
  NAND3BX4 U1992 ( .AN(n4897), .B(n4684), .C(n5321), .Y(n5184) );
  NAND3X6 U1993 ( .A(n6552), .B(n4683), .C(n6621), .Y(n5321) );
  OAI222X1 U1994 ( .A0(n3050), .A1(n8401), .B0(n8400), .B1(n18), .C0(
        \i_MIPS/PC/n4 ), .C1(n8457), .Y(n8406) );
  BUFX6 U1995 ( .A(n2901), .Y(n2155) );
  INVX8 U1996 ( .A(n3596), .Y(n3595) );
  OA22X4 U1997 ( .A0(n3462), .A1(n974), .B0(n3434), .B1(n86), .Y(n4469) );
  OA22X4 U1998 ( .A0(n3463), .A1(n975), .B0(n3436), .B1(n87), .Y(n4505) );
  OA22X2 U1999 ( .A0(n3549), .A1(n131), .B0(n3499), .B1(n1020), .Y(n4407) );
  OA22X2 U2000 ( .A0(n3365), .A1(n132), .B0(n3322), .B1(n1021), .Y(n4409) );
  OA22X2 U2001 ( .A0(n3575), .A1(n133), .B0(n3527), .B1(n1022), .Y(n4397) );
  OA22X2 U2002 ( .A0(n3374), .A1(n134), .B0(n3329), .B1(n1023), .Y(n4399) );
  OA22X2 U2003 ( .A0(n3575), .A1(n137), .B0(n3498), .B1(n1027), .Y(n4393) );
  OA22X2 U2004 ( .A0(n3363), .A1(n138), .B0(n3320), .B1(n1028), .Y(n4395) );
  NAND4X2 U2005 ( .A(n4519), .B(n4518), .C(n4517), .D(n4516), .Y(n8688) );
  XOR2X4 U2006 ( .A(n8177), .B(n8165), .Y(n6121) );
  OAI222X4 U2007 ( .A0(n6120), .A1(n3218), .B0(n6119), .B1(n3217), .C0(n8737), 
        .C1(n3215), .Y(n8165) );
  NAND4X4 U2008 ( .A(n4471), .B(n4470), .C(n4469), .D(n4468), .Y(n8697) );
  AOI222X2 U2009 ( .A0(\i_MIPS/IF_ID[65] ), .A1(n2157), .B0(n3048), .B1(
        \i_MIPS/BranchAddr[0] ), .C0(\i_MIPS/IF_ID_0 ), .C1(n3596), .Y(n8260)
         );
  NAND2X2 U2010 ( .A(n3050), .B(n2158), .Y(n3048) );
  BUFX20 U2011 ( .A(n2772), .Y(n2158) );
  OAI2BB1X4 U2012 ( .A0N(n6838), .A1N(n6837), .B0(n6841), .Y(n5988) );
  NAND2BX4 U2013 ( .AN(n5987), .B(n6693), .Y(n6838) );
  NAND4BX2 U2014 ( .AN(n8501), .B(n8500), .C(n8499), .D(n8498), .Y(n8503) );
  INVX6 U2015 ( .A(\i_MIPS/ALUin1[2] ), .Y(n5381) );
  NAND2X2 U2016 ( .A(\i_MIPS/ID_EX[78] ), .B(n4610), .Y(n4611) );
  CLKINVX1 U2017 ( .A(n8499), .Y(n5387) );
  AOI222X2 U2018 ( .A0(n6542), .A1(n6993), .B0(n6541), .B1(n6540), .C0(n6539), 
        .C1(n6538), .Y(n6543) );
  OAI222X2 U2019 ( .A0(n6902), .A1(n3166), .B0(n6901), .B1(n2761), .C0(n8730), 
        .C1(n3162), .Y(n6903) );
  AOI222X2 U2020 ( .A0(n6199), .A1(n6993), .B0(n6198), .B1(n6197), .C0(n6196), 
        .C1(n6195), .Y(n6213) );
  OAI221X4 U2021 ( .A0(n3106), .A1(n6193), .B0(n2820), .B1(n3098), .C0(n3097), 
        .Y(n6197) );
  AO22X1 U2022 ( .A0(n5603), .A1(n3102), .B0(n3110), .B1(n5604), .Y(n5608) );
  OAI222X4 U2023 ( .A0(n6597), .A1(n3166), .B0(n6575), .B1(n2761), .C0(n3162), 
        .C1(n8736), .Y(n8241) );
  AOI222X2 U2024 ( .A0(n2810), .A1(n6267), .B0(n6266), .B1(n6265), .C0(n6264), 
        .C1(n6263), .Y(n6276) );
  OA21X1 U2025 ( .A0(\i_MIPS/ALUin1[13] ), .A1(n3087), .B0(n5456), .Y(n4984)
         );
  OAI221X4 U2026 ( .A0(\i_MIPS/ALUin1[13] ), .A1(n3082), .B0(
        \i_MIPS/ALUin1[12] ), .B1(n3078), .C0(n5041), .Y(n5329) );
  OAI221X2 U2027 ( .A0(n8767), .A1(n7044), .B0(n8754), .B1(n7043), .C0(n6878), 
        .Y(n6879) );
  OAI221X4 U2028 ( .A0(n3106), .A1(n6986), .B0(n6987), .B1(n3099), .C0(n3097), 
        .Y(n6985) );
  OAI2BB1X4 U2029 ( .A0N(n5828), .A1N(n5811), .B0(n5821), .Y(n6986) );
  AOI222X2 U2030 ( .A0(n6608), .A1(n6993), .B0(n6607), .B1(n6606), .C0(n6605), 
        .C1(n6604), .Y(n6609) );
  OAI221X4 U2031 ( .A0(n3106), .A1(n6601), .B0(n6602), .B1(n3098), .C0(n3096), 
        .Y(n6606) );
  CLKINVX16 U2032 ( .A(n2162), .Y(n2163) );
  NAND2X2 U2033 ( .A(n7815), .B(n8684), .Y(n8130) );
  AOI211X4 U2034 ( .A0(n7789), .A1(\i_MIPS/n233 ), .B0(n7828), .C0(n1627), .Y(
        n7790) );
  INVX4 U2035 ( .A(n4669), .Y(n4678) );
  OAI33X4 U2036 ( .A0(n2843), .A1(n2875), .A2(n3099), .B0(n4708), .B1(n2875), 
        .B2(n2762), .Y(n4734) );
  INVXL U2037 ( .A(n2210), .Y(n2164) );
  INVXL U2038 ( .A(n2213), .Y(n2165) );
  CLKINVX1 U2039 ( .A(n4040), .Y(n2166) );
  CLKINVX1 U2040 ( .A(n4040), .Y(n2167) );
  CLKINVX1 U2041 ( .A(n4040), .Y(n2168) );
  CLKINVX1 U2042 ( .A(n4040), .Y(n2169) );
  CLKBUFX3 U2043 ( .A(n2166), .Y(n2170) );
  CLKBUFX3 U2044 ( .A(n2166), .Y(n2171) );
  CLKBUFX3 U2045 ( .A(n2166), .Y(n2172) );
  CLKBUFX3 U2046 ( .A(n2166), .Y(n2173) );
  CLKBUFX3 U2047 ( .A(n2166), .Y(n2174) );
  CLKBUFX3 U2048 ( .A(n2167), .Y(n2175) );
  CLKBUFX3 U2049 ( .A(n2167), .Y(n2176) );
  CLKBUFX3 U2050 ( .A(n2167), .Y(n2177) );
  CLKBUFX3 U2051 ( .A(n2167), .Y(n2178) );
  CLKBUFX3 U2052 ( .A(n2167), .Y(n2179) );
  CLKBUFX3 U2053 ( .A(n2168), .Y(n2180) );
  CLKBUFX3 U2054 ( .A(n2168), .Y(n2181) );
  CLKBUFX3 U2055 ( .A(n2168), .Y(n2182) );
  CLKBUFX3 U2056 ( .A(n2168), .Y(n2183) );
  CLKBUFX3 U2057 ( .A(n2168), .Y(n2184) );
  CLKBUFX3 U2058 ( .A(n2169), .Y(n2185) );
  CLKBUFX3 U2059 ( .A(n2169), .Y(n2186) );
  CLKBUFX3 U2060 ( .A(n2169), .Y(n2187) );
  CLKBUFX3 U2061 ( .A(n2169), .Y(n2188) );
  CLKBUFX3 U2062 ( .A(n2169), .Y(n2189) );
  CLKINVX1 U2063 ( .A(n4039), .Y(n2190) );
  CLKINVX1 U2064 ( .A(n4039), .Y(n2191) );
  CLKINVX1 U2065 ( .A(n4039), .Y(n2192) );
  CLKINVX1 U2066 ( .A(n4039), .Y(n2193) );
  CLKBUFX3 U2067 ( .A(n2190), .Y(n2194) );
  CLKBUFX3 U2068 ( .A(n2190), .Y(n2195) );
  CLKBUFX3 U2069 ( .A(n2190), .Y(n2196) );
  CLKBUFX3 U2070 ( .A(n2190), .Y(n2197) );
  CLKBUFX3 U2071 ( .A(n2190), .Y(n2198) );
  CLKBUFX3 U2072 ( .A(n2191), .Y(n2199) );
  CLKBUFX3 U2073 ( .A(n2191), .Y(n2200) );
  CLKBUFX3 U2074 ( .A(n2191), .Y(n2201) );
  CLKBUFX3 U2075 ( .A(n2191), .Y(n2202) );
  CLKBUFX3 U2076 ( .A(n2191), .Y(n2203) );
  CLKBUFX3 U2077 ( .A(n2192), .Y(n2204) );
  CLKBUFX3 U2078 ( .A(n2192), .Y(n2205) );
  CLKBUFX3 U2079 ( .A(n2192), .Y(n2206) );
  CLKBUFX3 U2080 ( .A(n2192), .Y(n2207) );
  CLKBUFX3 U2081 ( .A(n2192), .Y(n2208) );
  CLKBUFX3 U2082 ( .A(n2193), .Y(n2209) );
  CLKBUFX3 U2083 ( .A(n2193), .Y(n2210) );
  CLKBUFX3 U2084 ( .A(n2193), .Y(n2211) );
  CLKBUFX3 U2085 ( .A(n2193), .Y(n2212) );
  CLKBUFX3 U2086 ( .A(n2193), .Y(n2213) );
  CLKINVX1 U2087 ( .A(n4035), .Y(n2214) );
  CLKINVX1 U2088 ( .A(n4035), .Y(n2215) );
  CLKINVX1 U2089 ( .A(n4035), .Y(n2216) );
  CLKINVX1 U2090 ( .A(n4035), .Y(n2217) );
  CLKBUFX3 U2091 ( .A(n2214), .Y(n2218) );
  CLKBUFX3 U2092 ( .A(n2214), .Y(n2219) );
  CLKBUFX3 U2093 ( .A(n2214), .Y(n2220) );
  CLKBUFX3 U2094 ( .A(n2214), .Y(n2221) );
  BUFX12 U2095 ( .A(n2214), .Y(DCACHE_addr[3]) );
  CLKBUFX3 U2096 ( .A(n2215), .Y(n2223) );
  CLKBUFX3 U2097 ( .A(n2215), .Y(n2224) );
  CLKBUFX3 U2098 ( .A(n2215), .Y(n2225) );
  CLKBUFX3 U2099 ( .A(n2215), .Y(n2226) );
  CLKBUFX3 U2100 ( .A(n2215), .Y(n2227) );
  CLKBUFX3 U2101 ( .A(n2216), .Y(n2228) );
  CLKBUFX3 U2102 ( .A(n2216), .Y(n2229) );
  CLKBUFX3 U2103 ( .A(n2216), .Y(n2230) );
  CLKBUFX3 U2104 ( .A(n2216), .Y(n2231) );
  CLKBUFX3 U2105 ( .A(n2216), .Y(n2232) );
  CLKBUFX3 U2106 ( .A(n2217), .Y(n2233) );
  CLKBUFX3 U2107 ( .A(n2217), .Y(n2234) );
  CLKBUFX3 U2108 ( .A(n2217), .Y(n2235) );
  CLKBUFX3 U2109 ( .A(n2217), .Y(n2236) );
  CLKBUFX3 U2110 ( .A(n2217), .Y(n2237) );
  CLKINVX1 U2111 ( .A(n4036), .Y(n2238) );
  CLKINVX1 U2112 ( .A(n4036), .Y(n2239) );
  CLKINVX1 U2113 ( .A(n4036), .Y(n2240) );
  CLKINVX1 U2114 ( .A(n4036), .Y(n2241) );
  CLKBUFX3 U2115 ( .A(n2238), .Y(n2242) );
  CLKBUFX3 U2116 ( .A(n2238), .Y(n2243) );
  CLKBUFX3 U2117 ( .A(n2238), .Y(n2244) );
  CLKBUFX3 U2118 ( .A(n2238), .Y(n2245) );
  CLKBUFX3 U2119 ( .A(n2238), .Y(n2246) );
  CLKBUFX3 U2120 ( .A(n2239), .Y(n2247) );
  CLKBUFX3 U2121 ( .A(n2239), .Y(n2248) );
  CLKBUFX3 U2122 ( .A(n2239), .Y(n2249) );
  CLKBUFX3 U2123 ( .A(n2239), .Y(n2250) );
  CLKBUFX3 U2124 ( .A(n2239), .Y(n2251) );
  CLKBUFX3 U2125 ( .A(n2240), .Y(n2252) );
  CLKBUFX3 U2126 ( .A(n2240), .Y(n2253) );
  CLKBUFX3 U2127 ( .A(n2240), .Y(n2254) );
  CLKBUFX3 U2128 ( .A(n2240), .Y(n2255) );
  CLKBUFX3 U2129 ( .A(n2240), .Y(n2256) );
  CLKBUFX3 U2130 ( .A(n2241), .Y(n2257) );
  CLKBUFX3 U2131 ( .A(n2241), .Y(n2258) );
  CLKBUFX3 U2132 ( .A(n2241), .Y(n2259) );
  CLKBUFX3 U2133 ( .A(n2241), .Y(n2260) );
  CLKBUFX3 U2134 ( .A(n2241), .Y(n2261) );
  CLKINVX1 U2135 ( .A(n4038), .Y(n2262) );
  CLKINVX1 U2136 ( .A(n4038), .Y(n2263) );
  CLKINVX1 U2137 ( .A(n4038), .Y(n2264) );
  CLKINVX1 U2138 ( .A(n4038), .Y(n2265) );
  CLKBUFX3 U2139 ( .A(n2262), .Y(n2266) );
  CLKBUFX3 U2140 ( .A(n2262), .Y(n2267) );
  CLKBUFX3 U2141 ( .A(n2262), .Y(n2268) );
  CLKBUFX3 U2142 ( .A(n2262), .Y(n2269) );
  CLKBUFX3 U2143 ( .A(n2262), .Y(n2270) );
  CLKBUFX3 U2144 ( .A(n2263), .Y(n2271) );
  CLKBUFX3 U2145 ( .A(n2263), .Y(n2272) );
  CLKBUFX3 U2146 ( .A(n2263), .Y(n2273) );
  CLKBUFX3 U2147 ( .A(n2263), .Y(n2274) );
  CLKBUFX3 U2148 ( .A(n2263), .Y(n2275) );
  CLKBUFX3 U2149 ( .A(n2264), .Y(n2276) );
  CLKBUFX3 U2150 ( .A(n2264), .Y(n2277) );
  CLKBUFX3 U2151 ( .A(n2264), .Y(n2278) );
  CLKBUFX3 U2152 ( .A(n2264), .Y(n2279) );
  CLKBUFX3 U2153 ( .A(n2264), .Y(n2280) );
  CLKBUFX3 U2154 ( .A(n2265), .Y(n2281) );
  CLKBUFX3 U2155 ( .A(n2265), .Y(n2282) );
  CLKBUFX3 U2156 ( .A(n2265), .Y(n2283) );
  CLKBUFX3 U2157 ( .A(n2265), .Y(n2284) );
  CLKBUFX3 U2158 ( .A(n2265), .Y(n2285) );
  CLKINVX1 U2159 ( .A(n4037), .Y(n2286) );
  CLKINVX1 U2160 ( .A(n4037), .Y(n2287) );
  CLKINVX1 U2161 ( .A(n4037), .Y(n2288) );
  CLKINVX1 U2162 ( .A(n4037), .Y(n2289) );
  CLKBUFX3 U2163 ( .A(n2286), .Y(n2290) );
  CLKBUFX3 U2164 ( .A(n2286), .Y(n2291) );
  CLKBUFX3 U2165 ( .A(n2286), .Y(n2292) );
  CLKBUFX3 U2166 ( .A(n2286), .Y(n2293) );
  CLKBUFX3 U2167 ( .A(n2286), .Y(n2294) );
  CLKBUFX3 U2168 ( .A(n2287), .Y(n2295) );
  CLKBUFX3 U2169 ( .A(n2287), .Y(n2296) );
  CLKBUFX3 U2170 ( .A(n2287), .Y(n2297) );
  CLKBUFX3 U2171 ( .A(n2287), .Y(n2298) );
  CLKBUFX3 U2172 ( .A(n2287), .Y(n2299) );
  CLKBUFX3 U2173 ( .A(n2288), .Y(n2300) );
  CLKBUFX3 U2174 ( .A(n2288), .Y(n2301) );
  CLKBUFX3 U2175 ( .A(n2288), .Y(n2302) );
  CLKBUFX3 U2176 ( .A(n2288), .Y(n2303) );
  CLKBUFX3 U2177 ( .A(n2288), .Y(n2304) );
  CLKBUFX3 U2178 ( .A(n2289), .Y(n2305) );
  CLKBUFX3 U2179 ( .A(n2289), .Y(n2306) );
  CLKBUFX3 U2180 ( .A(n2289), .Y(n2307) );
  CLKBUFX3 U2181 ( .A(n2289), .Y(n2308) );
  CLKBUFX3 U2182 ( .A(n2289), .Y(n2309) );
  CLKINVX8 U2183 ( .A(n3061), .Y(n2371) );
  BUFX6 U2184 ( .A(n2372), .Y(n2385) );
  CLKBUFX4 U2185 ( .A(n2747), .Y(n2393) );
  CLKBUFX4 U2186 ( .A(n2747), .Y(n2394) );
  CLKBUFX4 U2187 ( .A(n2747), .Y(n2395) );
  CLKBUFX3 U2188 ( .A(n2747), .Y(n2396) );
  CLKBUFX3 U2189 ( .A(n2747), .Y(n2397) );
  CLKBUFX3 U2190 ( .A(n2747), .Y(n2398) );
  CLKBUFX3 U2191 ( .A(n2747), .Y(n2399) );
  CLKBUFX3 U2192 ( .A(n2747), .Y(n2400) );
  BUFX4 U2193 ( .A(n2396), .Y(n2417) );
  BUFX4 U2194 ( .A(n2396), .Y(n2420) );
  BUFX4 U2195 ( .A(n2397), .Y(n2421) );
  BUFX4 U2196 ( .A(n2397), .Y(n2425) );
  BUFX4 U2197 ( .A(n2398), .Y(n2429) );
  BUFX4 U2198 ( .A(n2398), .Y(n2430) );
  BUFX4 U2199 ( .A(n2400), .Y(n2436) );
  BUFX4 U2200 ( .A(n2400), .Y(n2439) );
  BUFX4 U2201 ( .A(n2400), .Y(n2440) );
  INVXL U2202 ( .A(n4035), .Y(n4034) );
  CLKINVX4 U2203 ( .A(n4036), .Y(n4033) );
  CLKINVX4 U2204 ( .A(n4037), .Y(n4032) );
  CLKBUFX2 U2205 ( .A(n4040), .Y(n4039) );
  CLKBUFX2 U2206 ( .A(n4040), .Y(n4035) );
  CLKBUFX2 U2207 ( .A(n4040), .Y(n4036) );
  CLKBUFX2 U2208 ( .A(n4040), .Y(n4038) );
  CLKBUFX2 U2209 ( .A(n4040), .Y(n4037) );
  MXI2X4 U2210 ( .A(n10310), .B(DCACHE_rdata[18]), .S0(n4023), .Y(n8731) );
  CLKINVX4 U2211 ( .A(n8381), .Y(n8388) );
  NAND2X4 U2212 ( .A(n8383), .B(n8381), .Y(n8349) );
  NAND4X4 U2213 ( .A(n7366), .B(n7365), .C(n7364), .D(n7363), .Y(n8381) );
  OAI2BB1X4 U2214 ( .A0N(n5732), .A1N(n4827), .B0(n4826), .Y(n5601) );
  OAI221X4 U2215 ( .A0(\D_cache/n164 ), .A1(n8858), .B0(n3074), .B1(n8839), 
        .C0(\D_cache/n196 ), .Y(DCACHE_rdata[12]) );
  OR2X1 U2216 ( .A(n8871), .B(n4002), .Y(n10168) );
  INVX12 U2217 ( .A(n10168), .Y(mem_wdata_D[127]) );
  CLKINVX2 U2218 ( .A(n2866), .Y(n4002) );
  OR2X1 U2219 ( .A(n8878), .B(n4001), .Y(n10175) );
  INVX12 U2220 ( .A(n10175), .Y(mem_wdata_D[120]) );
  CLKINVX2 U2221 ( .A(mem_write_D), .Y(n4001) );
  OR2X1 U2222 ( .A(n8853), .B(n4005), .Y(n10246) );
  INVX12 U2223 ( .A(n10246), .Y(mem_wdata_D[49]) );
  CLKINVX2 U2224 ( .A(n2866), .Y(n4005) );
  OR2X1 U2225 ( .A(n8899), .B(n3998), .Y(n10196) );
  INVX12 U2226 ( .A(n10196), .Y(mem_wdata_D[99]) );
  CLKINVX2 U2227 ( .A(mem_write_D), .Y(n3998) );
  BUFX12 U2228 ( .A(n10200), .Y(mem_wdata_D[95]) );
  NOR2BX1 U2229 ( .AN(\D_cache/N121 ), .B(n4007), .Y(n10200) );
  BUFX12 U2230 ( .A(n10215), .Y(mem_wdata_D[80]) );
  NOR2BXL U2231 ( .AN(\D_cache/N136 ), .B(n4007), .Y(n10215) );
  INVX12 U2232 ( .A(n2448), .Y(mem_addr_D[26]) );
  NOR2XL U2233 ( .A(n1618), .B(n4011), .Y(n2449) );
  NOR2XL U2234 ( .A(n8813), .B(n4006), .Y(n2450) );
  NOR2XL U2235 ( .A(n2449), .B(n2450), .Y(n2448) );
  INVX12 U2236 ( .A(n2451), .Y(mem_addr_D[25]) );
  NOR2X1 U2237 ( .A(n1089), .B(n4011), .Y(n2452) );
  NOR2XL U2238 ( .A(n8814), .B(n4007), .Y(n2453) );
  NOR2XL U2239 ( .A(n2452), .B(n2453), .Y(n2451) );
  OR2X1 U2240 ( .A(n8872), .B(n4002), .Y(n10169) );
  INVX12 U2241 ( .A(n10169), .Y(mem_wdata_D[126]) );
  OR2X1 U2242 ( .A(n8873), .B(n4002), .Y(n10170) );
  INVX12 U2243 ( .A(n10170), .Y(mem_wdata_D[125]) );
  OR2X1 U2244 ( .A(n8874), .B(n4002), .Y(n10171) );
  INVX12 U2245 ( .A(n10171), .Y(mem_wdata_D[124]) );
  OR2X1 U2246 ( .A(n8879), .B(n4001), .Y(n10176) );
  INVX12 U2247 ( .A(n10176), .Y(mem_wdata_D[119]) );
  OR2X1 U2248 ( .A(n8885), .B(n3999), .Y(n10182) );
  INVX12 U2249 ( .A(n10182), .Y(mem_wdata_D[113]) );
  CLKINVX2 U2250 ( .A(mem_write_D), .Y(n3999) );
  OR2X1 U2251 ( .A(n8854), .B(n4005), .Y(n10247) );
  INVX12 U2252 ( .A(n10247), .Y(mem_wdata_D[48]) );
  OR2X1 U2253 ( .A(n8900), .B(n3998), .Y(n10197) );
  INVX12 U2254 ( .A(n10197), .Y(mem_wdata_D[98]) );
  BUFX12 U2255 ( .A(n10216), .Y(mem_wdata_D[79]) );
  NOR2BXL U2256 ( .AN(\D_cache/N137 ), .B(n4002), .Y(n10216) );
  BUFX12 U2257 ( .A(n10202), .Y(mem_wdata_D[93]) );
  NOR2BXL U2258 ( .AN(\D_cache/N123 ), .B(n4007), .Y(n10202) );
  BUFX12 U2259 ( .A(n10203), .Y(mem_wdata_D[92]) );
  NOR2BXL U2260 ( .AN(\D_cache/N124 ), .B(n4007), .Y(n10203) );
  INVX12 U2261 ( .A(n2464), .Y(mem_addr_D[13]) );
  NOR2X1 U2262 ( .A(n1621), .B(n4011), .Y(n2465) );
  NOR2XL U2263 ( .A(n8826), .B(n4006), .Y(n2466) );
  NOR2XL U2264 ( .A(n2465), .B(n2466), .Y(n2464) );
  INVX12 U2265 ( .A(n2467), .Y(mem_addr_D[24]) );
  NOR2X1 U2266 ( .A(n1090), .B(n4010), .Y(n2468) );
  NOR2XL U2267 ( .A(n8815), .B(n4004), .Y(n2469) );
  NOR2XL U2268 ( .A(n2468), .B(n2469), .Y(n2467) );
  OR2X1 U2269 ( .A(n8875), .B(n4002), .Y(n10172) );
  INVX12 U2270 ( .A(n10172), .Y(mem_wdata_D[123]) );
  OR2X1 U2271 ( .A(n8880), .B(n4001), .Y(n10177) );
  INVX12 U2272 ( .A(n10177), .Y(mem_wdata_D[118]) );
  OR2X1 U2273 ( .A(n8889), .B(n4000), .Y(n10186) );
  INVX12 U2274 ( .A(n10186), .Y(mem_wdata_D[109]) );
  CLKINVX2 U2275 ( .A(n2866), .Y(n4000) );
  OR2X1 U2276 ( .A(n8762), .B(n3999), .Y(n10235) );
  INVX12 U2277 ( .A(n10235), .Y(mem_wdata_D[60]) );
  OR2X1 U2278 ( .A(n8855), .B(n4005), .Y(n10248) );
  INVX12 U2279 ( .A(n10248), .Y(mem_wdata_D[47]) );
  OR2X1 U2280 ( .A(n8856), .B(n4005), .Y(n10249) );
  INVX12 U2281 ( .A(n10249), .Y(mem_wdata_D[46]) );
  OR2X1 U2282 ( .A(n8864), .B(n4004), .Y(n10257) );
  INVX12 U2283 ( .A(n10257), .Y(mem_wdata_D[38]) );
  CLKINVX2 U2284 ( .A(n2866), .Y(n4004) );
  OR2X1 U2285 ( .A(n8750), .B(n4003), .Y(n10268) );
  INVX12 U2286 ( .A(n10268), .Y(mem_wdata_D[27]) );
  CLKINVX2 U2287 ( .A(mem_write_D), .Y(n4003) );
  OR2X1 U2288 ( .A(n8751), .B(n4003), .Y(n10269) );
  INVX12 U2289 ( .A(n10269), .Y(mem_wdata_D[26]) );
  OR2X1 U2290 ( .A(n8752), .B(n4003), .Y(n10270) );
  INVX12 U2291 ( .A(n10270), .Y(mem_wdata_D[25]) );
  BUFX12 U2292 ( .A(n10271), .Y(mem_wdata_D[24]) );
  NOR2XL U2293 ( .A(n8753), .B(n4003), .Y(n10271) );
  OR2X1 U2294 ( .A(n8754), .B(n4003), .Y(n10272) );
  INVX12 U2295 ( .A(n10272), .Y(mem_wdata_D[23]) );
  OR2X1 U2296 ( .A(n8901), .B(n3998), .Y(n10198) );
  INVX12 U2297 ( .A(n10198), .Y(mem_wdata_D[97]) );
  BUFX12 U2298 ( .A(n10206), .Y(mem_wdata_D[89]) );
  NOR2BXL U2299 ( .AN(\D_cache/N127 ), .B(n4007), .Y(n10206) );
  BUFX12 U2300 ( .A(n10218), .Y(mem_wdata_D[77]) );
  NOR2BXL U2301 ( .AN(\D_cache/N139 ), .B(n4003), .Y(n10218) );
  INVX12 U2302 ( .A(n2485), .Y(mem_addr_D[12]) );
  NOR2X1 U2303 ( .A(n3037), .B(n4010), .Y(n2486) );
  NOR2XL U2304 ( .A(n8827), .B(n4006), .Y(n2487) );
  NOR2XL U2305 ( .A(n2486), .B(n2487), .Y(n2485) );
  INVX12 U2306 ( .A(n2488), .Y(mem_addr_D[23]) );
  NOR2XL U2307 ( .A(n1619), .B(n4011), .Y(n2489) );
  NOR2XL U2308 ( .A(n8816), .B(n4005), .Y(n2490) );
  NOR2XL U2309 ( .A(n2489), .B(n2490), .Y(n2488) );
  INVX12 U2310 ( .A(n2491), .Y(mem_addr_I[23]) );
  INVXL U2311 ( .A(n8704), .Y(n2492) );
  NOR2X1 U2312 ( .A(n2492), .B(n3052), .Y(n2493) );
  NOR2XL U2313 ( .A(n2516), .B(\i_MIPS/PC/n25 ), .Y(n2494) );
  NOR2XL U2314 ( .A(n2493), .B(n2494), .Y(n2491) );
  OR2X1 U2315 ( .A(n8876), .B(n4002), .Y(n10173) );
  INVX12 U2316 ( .A(n10173), .Y(mem_wdata_D[122]) );
  OR2X1 U2317 ( .A(n8881), .B(n4001), .Y(n10178) );
  INVX12 U2318 ( .A(n10178), .Y(mem_wdata_D[117]) );
  OR2X1 U2319 ( .A(n8890), .B(n4000), .Y(n10187) );
  INVX12 U2320 ( .A(n10187), .Y(mem_wdata_D[108]) );
  OR2X1 U2321 ( .A(n8891), .B(n4000), .Y(n10188) );
  INVX12 U2322 ( .A(n10188), .Y(mem_wdata_D[107]) );
  OR2X1 U2323 ( .A(n8763), .B(n3999), .Y(n10236) );
  INVX12 U2324 ( .A(n10236), .Y(mem_wdata_D[59]) );
  OR2X1 U2325 ( .A(n8764), .B(n3999), .Y(n10237) );
  INVX12 U2326 ( .A(n10237), .Y(mem_wdata_D[58]) );
  OR2X1 U2327 ( .A(n8857), .B(n4005), .Y(n10250) );
  INVX12 U2328 ( .A(n10250), .Y(mem_wdata_D[45]) );
  OR2X1 U2329 ( .A(n8865), .B(n4004), .Y(n10258) );
  INVX12 U2330 ( .A(n10258), .Y(mem_wdata_D[37]) );
  OR2X1 U2331 ( .A(n8866), .B(n4004), .Y(n10259) );
  INVX12 U2332 ( .A(n10259), .Y(mem_wdata_D[36]) );
  BUFX12 U2333 ( .A(n10273), .Y(mem_wdata_D[22]) );
  NOR2XL U2334 ( .A(n8755), .B(n4003), .Y(n10273) );
  OR2X1 U2335 ( .A(n8902), .B(n3998), .Y(n10199) );
  INVX12 U2336 ( .A(n10199), .Y(mem_wdata_D[96]) );
  BUFX12 U2337 ( .A(n10219), .Y(mem_wdata_D[76]) );
  NOR2BXL U2338 ( .AN(\D_cache/N140 ), .B(n4006), .Y(n10219) );
  BUFX12 U2339 ( .A(n10201), .Y(mem_wdata_D[94]) );
  NOR2BXL U2340 ( .AN(\D_cache/N122 ), .B(n4007), .Y(n10201) );
  INVX12 U2341 ( .A(n2508), .Y(mem_addr_D[11]) );
  NOR2X1 U2342 ( .A(n1622), .B(n4010), .Y(n2509) );
  NOR2XL U2343 ( .A(n8828), .B(n4006), .Y(n2510) );
  NOR2XL U2344 ( .A(n2509), .B(n2510), .Y(n2508) );
  INVX12 U2345 ( .A(n2511), .Y(mem_addr_D[22]) );
  NOR2XL U2346 ( .A(n1091), .B(n4010), .Y(n2512) );
  NOR2XL U2347 ( .A(n8817), .B(n4000), .Y(n2513) );
  NOR2XL U2348 ( .A(n2512), .B(n2513), .Y(n2511) );
  INVX12 U2349 ( .A(n2514), .Y(mem_addr_I[19]) );
  INVXL U2350 ( .A(n8700), .Y(n2515) );
  CLKINVX1 U2351 ( .A(mem_read_I), .Y(n2516) );
  NOR2X1 U2352 ( .A(n2515), .B(n3052), .Y(n2517) );
  NOR2XL U2353 ( .A(n2516), .B(\i_MIPS/PC/n21 ), .Y(n2518) );
  NOR2XL U2354 ( .A(n2517), .B(n2518), .Y(n2514) );
  OR2X1 U2355 ( .A(n8877), .B(n4002), .Y(n10174) );
  INVX12 U2356 ( .A(n10174), .Y(mem_wdata_D[121]) );
  OR2X1 U2357 ( .A(n8882), .B(n4001), .Y(n10179) );
  INVX12 U2358 ( .A(n10179), .Y(mem_wdata_D[116]) );
  OR2X1 U2359 ( .A(n8883), .B(n4001), .Y(n10180) );
  INVX12 U2360 ( .A(n10180), .Y(mem_wdata_D[115]) );
  OR2X1 U2361 ( .A(n8884), .B(n4001), .Y(n10181) );
  INVX12 U2362 ( .A(n10181), .Y(mem_wdata_D[114]) );
  BUFX12 U2363 ( .A(n10183), .Y(mem_wdata_D[112]) );
  NOR2XL U2364 ( .A(n8886), .B(n4001), .Y(n10183) );
  OR2X1 U2365 ( .A(n8892), .B(n4000), .Y(n10189) );
  INVX12 U2366 ( .A(n10189), .Y(mem_wdata_D[106]) );
  OR2X1 U2367 ( .A(n8765), .B(n3999), .Y(n10238) );
  INVX12 U2368 ( .A(n10238), .Y(mem_wdata_D[57]) );
  OR2X1 U2369 ( .A(n8858), .B(n4005), .Y(n10251) );
  INVX12 U2370 ( .A(n10251), .Y(mem_wdata_D[44]) );
  OR2X1 U2371 ( .A(n8867), .B(n4004), .Y(n10260) );
  INVX12 U2372 ( .A(n10260), .Y(mem_wdata_D[35]) );
  BUFX12 U2373 ( .A(n10263), .Y(mem_wdata_D[32]) );
  NOR2XL U2374 ( .A(n8870), .B(n4002), .Y(n10263) );
  OR2X1 U2375 ( .A(n8756), .B(n4003), .Y(n10274) );
  INVX12 U2376 ( .A(n10274), .Y(mem_wdata_D[21]) );
  OR2X1 U2377 ( .A(n8757), .B(n4003), .Y(n10275) );
  INVX12 U2378 ( .A(n10275), .Y(mem_wdata_D[20]) );
  OR2X1 U2379 ( .A(n8759), .B(n3998), .Y(n10232) );
  INVX12 U2380 ( .A(n10232), .Y(mem_wdata_D[63]) );
  BUFX12 U2381 ( .A(n10220), .Y(mem_wdata_D[75]) );
  NOR2BXL U2382 ( .AN(\D_cache/N141 ), .B(n4001), .Y(n10220) );
  BUFX12 U2383 ( .A(n10205), .Y(mem_wdata_D[90]) );
  NOR2BXL U2384 ( .AN(\D_cache/N126 ), .B(n4007), .Y(n10205) );
  INVX12 U2385 ( .A(n2534), .Y(mem_addr_D[10]) );
  NOR2XL U2386 ( .A(n1626), .B(n4011), .Y(n2535) );
  NOR2XL U2387 ( .A(n8829), .B(n4006), .Y(n2536) );
  NOR2XL U2388 ( .A(n2535), .B(n2536), .Y(n2534) );
  INVX12 U2389 ( .A(n2537), .Y(mem_addr_D[21]) );
  NOR2X1 U2390 ( .A(n1088), .B(n4011), .Y(n2538) );
  NOR2XL U2391 ( .A(n8818), .B(n4003), .Y(n2539) );
  CLKBUFX2 U2392 ( .A(\D_cache/n522 ), .Y(n4011) );
  INVX12 U2393 ( .A(n2540), .Y(mem_addr_I[18]) );
  INVXL U2394 ( .A(n8699), .Y(n2541) );
  NOR2X1 U2395 ( .A(n2541), .B(n3052), .Y(n2542) );
  NOR2XL U2396 ( .A(n2516), .B(\i_MIPS/PC/n20 ), .Y(n2543) );
  NOR2XL U2397 ( .A(n2542), .B(n2543), .Y(n2540) );
  OR2X1 U2398 ( .A(n8887), .B(n4001), .Y(n10184) );
  INVX12 U2399 ( .A(n10184), .Y(mem_wdata_D[111]) );
  OR2X1 U2400 ( .A(n8893), .B(n4000), .Y(n10190) );
  INVX12 U2401 ( .A(n10190), .Y(mem_wdata_D[105]) );
  OR2X1 U2402 ( .A(n8766), .B(n3999), .Y(n10239) );
  INVX12 U2403 ( .A(n10239), .Y(mem_wdata_D[56]) );
  OR2X1 U2404 ( .A(n8767), .B(n3999), .Y(n10240) );
  INVX12 U2405 ( .A(n10240), .Y(mem_wdata_D[55]) );
  BUFX12 U2406 ( .A(n10241), .Y(mem_wdata_D[54]) );
  NOR2XL U2407 ( .A(n8768), .B(n3999), .Y(n10241) );
  OR2X1 U2408 ( .A(n8770), .B(n3999), .Y(n10243) );
  INVX12 U2409 ( .A(n10243), .Y(mem_wdata_D[52]) );
  OR2X1 U2410 ( .A(n8859), .B(n4005), .Y(n10252) );
  INVX12 U2411 ( .A(n10252), .Y(mem_wdata_D[43]) );
  OR2X1 U2412 ( .A(n8860), .B(n4005), .Y(n10253) );
  INVX12 U2413 ( .A(n10253), .Y(mem_wdata_D[42]) );
  OR2X1 U2414 ( .A(n8868), .B(n4004), .Y(n10261) );
  INVX12 U2415 ( .A(n10261), .Y(mem_wdata_D[34]) );
  OR2X1 U2416 ( .A(n8869), .B(n4004), .Y(n10262) );
  INVX12 U2417 ( .A(n10262), .Y(mem_wdata_D[33]) );
  BUFX12 U2418 ( .A(n10264), .Y(mem_wdata_D[31]) );
  NOR2XL U2419 ( .A(n8746), .B(n4004), .Y(n10264) );
  OR2X1 U2420 ( .A(n8747), .B(n4004), .Y(n10265) );
  INVX12 U2421 ( .A(n10265), .Y(mem_wdata_D[30]) );
  OR2X1 U2422 ( .A(n8758), .B(n4003), .Y(n10276) );
  INVX12 U2423 ( .A(n10276), .Y(mem_wdata_D[19]) );
  OR2X1 U2424 ( .A(n8835), .B(n4002), .Y(n10279) );
  INVX12 U2425 ( .A(n10279), .Y(mem_wdata_D[16]) );
  OR2X1 U2426 ( .A(n8760), .B(n3998), .Y(n10233) );
  INVX12 U2427 ( .A(n10233), .Y(mem_wdata_D[62]) );
  OR2X1 U2428 ( .A(n8761), .B(n3998), .Y(n10234) );
  INVX12 U2429 ( .A(n10234), .Y(mem_wdata_D[61]) );
  OR2X1 U2430 ( .A(n8769), .B(n3998), .Y(n10242) );
  INVX12 U2431 ( .A(n10242), .Y(mem_wdata_D[53]) );
  OR2X1 U2432 ( .A(n8842), .B(n3998), .Y(n10286) );
  INVX12 U2433 ( .A(n10286), .Y(mem_wdata_D[9]) );
  BUFX12 U2434 ( .A(n10221), .Y(mem_wdata_D[74]) );
  NOR2BXL U2435 ( .AN(\D_cache/N142 ), .B(n4007), .Y(n10221) );
  BUFX12 U2436 ( .A(n10207), .Y(mem_wdata_D[88]) );
  NOR2BXL U2437 ( .AN(\D_cache/N128 ), .B(n4007), .Y(n10207) );
  BUFX12 U2438 ( .A(n10208), .Y(mem_wdata_D[87]) );
  NOR2BXL U2439 ( .AN(\D_cache/N129 ), .B(n4007), .Y(n10208) );
  BUFX12 U2440 ( .A(n10210), .Y(mem_wdata_D[85]) );
  NOR2BXL U2441 ( .AN(\D_cache/N131 ), .B(n4007), .Y(n10210) );
  INVX12 U2442 ( .A(n2566), .Y(mem_addr_D[9]) );
  NOR2X1 U2443 ( .A(n1624), .B(n4010), .Y(n2567) );
  NOR2XL U2444 ( .A(n8830), .B(n4006), .Y(n2568) );
  NOR2XL U2445 ( .A(n2567), .B(n2568), .Y(n2566) );
  INVX12 U2446 ( .A(n2569), .Y(mem_addr_D[20]) );
  NOR2X1 U2447 ( .A(n1087), .B(n4011), .Y(n2570) );
  NOR2XL U2448 ( .A(n8819), .B(n4002), .Y(n2571) );
  NOR2XL U2449 ( .A(n2570), .B(n2571), .Y(n2569) );
  INVX12 U2450 ( .A(n2572), .Y(mem_addr_I[29]) );
  INVXL U2451 ( .A(n8710), .Y(n2573) );
  NOR2X1 U2452 ( .A(n2573), .B(n3052), .Y(n2574) );
  NOR2XL U2453 ( .A(n2516), .B(\i_MIPS/PC/n31 ), .Y(n2575) );
  NOR2XL U2454 ( .A(n2574), .B(n2575), .Y(n2572) );
  INVX12 U2455 ( .A(n2576), .Y(mem_addr_I[28]) );
  INVXL U2456 ( .A(n8709), .Y(n2577) );
  NOR2X1 U2457 ( .A(n2577), .B(n3052), .Y(n2578) );
  NOR2XL U2458 ( .A(n2516), .B(\i_MIPS/PC/n30 ), .Y(n2579) );
  NOR2XL U2459 ( .A(n2578), .B(n2579), .Y(n2576) );
  BUFX16 U2460 ( .A(n8714), .Y(mem_write_I) );
  OR2X1 U2461 ( .A(n8888), .B(n4001), .Y(n10185) );
  INVX12 U2462 ( .A(n10185), .Y(mem_wdata_D[110]) );
  OR2X1 U2463 ( .A(n8894), .B(n4000), .Y(n10191) );
  INVX12 U2464 ( .A(n10191), .Y(mem_wdata_D[104]) );
  OR2X1 U2465 ( .A(n8895), .B(n4000), .Y(n10192) );
  INVX12 U2466 ( .A(n10192), .Y(mem_wdata_D[103]) );
  BUFX12 U2467 ( .A(n10193), .Y(mem_wdata_D[102]) );
  NOR2XL U2468 ( .A(n8896), .B(n4000), .Y(n10193) );
  OR2X1 U2469 ( .A(n8897), .B(n4000), .Y(n10194) );
  INVX12 U2470 ( .A(n10194), .Y(mem_wdata_D[101]) );
  BUFX12 U2471 ( .A(n10195), .Y(mem_wdata_D[100]) );
  NOR2XL U2472 ( .A(n8898), .B(n4000), .Y(n10195) );
  OR2X1 U2473 ( .A(n8771), .B(n3999), .Y(n10244) );
  INVX12 U2474 ( .A(n10244), .Y(mem_wdata_D[51]) );
  BUFX12 U2475 ( .A(n10254), .Y(mem_wdata_D[41]) );
  NOR2XL U2476 ( .A(n8861), .B(n4005), .Y(n10254) );
  BUFX12 U2477 ( .A(n10255), .Y(mem_wdata_D[40]) );
  NOR2XL U2478 ( .A(n8862), .B(n4005), .Y(n10255) );
  BUFX12 U2479 ( .A(n10266), .Y(mem_wdata_D[29]) );
  NOR2XL U2480 ( .A(n8748), .B(n4004), .Y(n10266) );
  OR2X1 U2481 ( .A(n8833), .B(n4003), .Y(n10277) );
  INVX12 U2482 ( .A(n10277), .Y(mem_wdata_D[18]) );
  OR2X1 U2483 ( .A(n8837), .B(n4002), .Y(n10281) );
  INVX12 U2484 ( .A(n10281), .Y(mem_wdata_D[14]) );
  OR2X1 U2485 ( .A(n8843), .B(n3998), .Y(n10287) );
  INVX12 U2486 ( .A(n10287), .Y(mem_wdata_D[8]) );
  BUFX12 U2487 ( .A(n10204), .Y(mem_wdata_D[91]) );
  NOR2BXL U2488 ( .AN(\D_cache/N125 ), .B(n4007), .Y(n10204) );
  BUFX12 U2489 ( .A(n10225), .Y(mem_wdata_D[70]) );
  NOR2BXL U2490 ( .AN(\D_cache/N146 ), .B(n4007), .Y(n10225) );
  BUFX12 U2491 ( .A(n10228), .Y(mem_wdata_D[67]) );
  NOR2BXL U2492 ( .AN(\D_cache/N149 ), .B(n4007), .Y(n10228) );
  INVX12 U2493 ( .A(n2596), .Y(mem_addr_D[8]) );
  NOR2X1 U2494 ( .A(n1623), .B(n4011), .Y(n2597) );
  NOR2XL U2495 ( .A(n8831), .B(n4006), .Y(n2598) );
  NOR2XL U2496 ( .A(n2597), .B(n2598), .Y(n2596) );
  INVX12 U2497 ( .A(n2599), .Y(mem_addr_D[19]) );
  NOR2XL U2498 ( .A(n1617), .B(n4011), .Y(n2600) );
  NOR2XL U2499 ( .A(n8820), .B(n4001), .Y(n2601) );
  INVX12 U2500 ( .A(n2602), .Y(mem_addr_I[26]) );
  INVXL U2501 ( .A(n8707), .Y(n2603) );
  NOR2X1 U2502 ( .A(n2603), .B(n3052), .Y(n2604) );
  NOR2XL U2503 ( .A(n2516), .B(\i_MIPS/PC/n28 ), .Y(n2605) );
  NOR2XL U2504 ( .A(n2604), .B(n2605), .Y(n2602) );
  INVX12 U2505 ( .A(n2606), .Y(mem_addr_I[24]) );
  INVXL U2506 ( .A(n8705), .Y(n2607) );
  NOR2X1 U2507 ( .A(n2607), .B(n3052), .Y(n2608) );
  NOR2XL U2508 ( .A(n8687), .B(\i_MIPS/PC/n26 ), .Y(n2609) );
  NOR2X1 U2509 ( .A(n2608), .B(n2609), .Y(n2606) );
  OR2X1 U2510 ( .A(n8852), .B(n3999), .Y(n10245) );
  INVX12 U2511 ( .A(n10245), .Y(mem_wdata_D[50]) );
  OR2X1 U2512 ( .A(n8863), .B(n4005), .Y(n10256) );
  INVX12 U2513 ( .A(n10256), .Y(mem_wdata_D[39]) );
  BUFX12 U2514 ( .A(n10267), .Y(mem_wdata_D[28]) );
  NOR2XL U2515 ( .A(n8749), .B(n4004), .Y(n10267) );
  OR2X1 U2516 ( .A(n8834), .B(n4003), .Y(n10278) );
  INVX12 U2517 ( .A(n10278), .Y(mem_wdata_D[17]) );
  OR2X1 U2518 ( .A(n8836), .B(n4001), .Y(n10280) );
  INVX12 U2519 ( .A(n10280), .Y(mem_wdata_D[15]) );
  OR2X1 U2520 ( .A(n8838), .B(n4002), .Y(n10282) );
  INVX12 U2521 ( .A(n10282), .Y(mem_wdata_D[13]) );
  OR2X1 U2522 ( .A(n8841), .B(n4000), .Y(n10285) );
  INVX12 U2523 ( .A(n10285), .Y(mem_wdata_D[10]) );
  BUFX12 U2524 ( .A(n10291), .Y(mem_wdata_D[4]) );
  NOR2XL U2525 ( .A(n8847), .B(n4004), .Y(n10291) );
  BUFX12 U2526 ( .A(n10165), .Y(mem_addr_D[6]) );
  NOR2XL U2527 ( .A(\D_cache/n523 ), .B(n2151), .Y(n10165) );
  NOR2X1 U2528 ( .A(mem_write_D), .B(mem_read_D), .Y(\D_cache/n523 ) );
  OR2X1 U2529 ( .A(n8844), .B(n3998), .Y(n10288) );
  INVX12 U2530 ( .A(n10288), .Y(mem_wdata_D[7]) );
  CLKAND2X12 U2531 ( .A(ICACHE_addr[4]), .B(n8686), .Y(mem_addr_I[6]) );
  BUFX12 U2532 ( .A(n10222), .Y(mem_wdata_D[73]) );
  NOR2BXL U2533 ( .AN(\D_cache/N143 ), .B(n4006), .Y(n10222) );
  BUFX12 U2534 ( .A(n10223), .Y(mem_wdata_D[72]) );
  NOR2BXL U2535 ( .AN(\D_cache/N144 ), .B(n3998), .Y(n10223) );
  BUFX12 U2536 ( .A(n10209), .Y(mem_wdata_D[86]) );
  NOR2BXL U2537 ( .AN(\D_cache/N130 ), .B(n4007), .Y(n10209) );
  INVX12 U2538 ( .A(n2623), .Y(mem_addr_D[14]) );
  NOR2XL U2539 ( .A(n1071), .B(n4010), .Y(n2624) );
  NOR2XL U2540 ( .A(n8825), .B(n4006), .Y(n2625) );
  NOR2XL U2541 ( .A(n2624), .B(n2625), .Y(n2623) );
  CLKBUFX2 U2542 ( .A(\D_cache/n522 ), .Y(n4010) );
  INVX12 U2543 ( .A(n2626), .Y(mem_addr_D[16]) );
  NOR2XL U2544 ( .A(n1070), .B(n4010), .Y(n2627) );
  NOR2XL U2545 ( .A(n8823), .B(n3999), .Y(n2628) );
  NOR2XL U2546 ( .A(n2627), .B(n2628), .Y(n2626) );
  CLKBUFX3 U2547 ( .A(n8723), .Y(n3644) );
  CLKBUFX3 U2548 ( .A(n8737), .Y(n3671) );
  CLKBUFX3 U2549 ( .A(n8719), .Y(n3639) );
  CLKBUFX3 U2550 ( .A(n8717), .Y(n3635) );
  CLKBUFX3 U2551 ( .A(n8743), .Y(n3684) );
  CLKBUFX3 U2552 ( .A(n8720), .Y(n3641) );
  CLKBUFX3 U2553 ( .A(n8739), .Y(n3675) );
  CLKBUFX3 U2554 ( .A(n8738), .Y(n3673) );
  CLKBUFX3 U2555 ( .A(n8734), .Y(n3666) );
  MXI2X4 U2556 ( .A(n3063), .B(DCACHE_rdata[6]), .S0(n4023), .Y(n8734) );
  MXI2X1 U2557 ( .A(n2129), .B(DCACHE_rdata[4]), .S0(n4023), .Y(n8735) );
  BUFX12 U2558 ( .A(n10356), .Y(DCACHE_wen) );
  INVX12 U2559 ( .A(n2630), .Y(mem_addr_D[31]) );
  INVXL U2560 ( .A(\D_cache/N32 ), .Y(n2631) );
  NOR2X1 U2561 ( .A(n4007), .B(n2631), .Y(n2632) );
  NOR2XL U2562 ( .A(n4011), .B(n1847), .Y(n2633) );
  NOR2XL U2563 ( .A(n2632), .B(n2633), .Y(n2630) );
  BUFX16 U2564 ( .A(n2866), .Y(mem_write_D) );
  INVX12 U2565 ( .A(n962), .Y(mem_addr_I[17]) );
  BUFX12 U2566 ( .A(n10296), .Y(mem_addr_I[25]) );
  AO22XL U2567 ( .A0(ICACHE_addr[23]), .A1(mem_read_I), .B0(mem_write_I), .B1(
        n8706), .Y(n10296) );
  OR2X1 U2568 ( .A(n8839), .B(n4002), .Y(n10283) );
  INVX12 U2569 ( .A(n10283), .Y(mem_wdata_D[12]) );
  OR2X1 U2570 ( .A(n8840), .B(n4001), .Y(n10284) );
  INVX12 U2571 ( .A(n10284), .Y(mem_wdata_D[11]) );
  OR2X1 U2572 ( .A(n8846), .B(n3999), .Y(n10290) );
  INVX12 U2573 ( .A(n10290), .Y(mem_wdata_D[5]) );
  OR2X1 U2574 ( .A(n8848), .B(n4005), .Y(n10292) );
  INVX12 U2575 ( .A(n10292), .Y(mem_wdata_D[3]) );
  OR2X1 U2576 ( .A(n8849), .B(n4004), .Y(n10293) );
  INVX12 U2577 ( .A(n10293), .Y(mem_wdata_D[2]) );
  OR2X1 U2578 ( .A(n8850), .B(n4003), .Y(n10294) );
  INVX12 U2579 ( .A(n10294), .Y(mem_wdata_D[1]) );
  OR2X1 U2580 ( .A(n8851), .B(n4000), .Y(n10295) );
  INVX12 U2581 ( .A(n10295), .Y(mem_wdata_D[0]) );
  OR2X1 U2582 ( .A(\D_cache/n523 ), .B(n2165), .Y(n10166) );
  INVX12 U2583 ( .A(n10166), .Y(mem_addr_D[5]) );
  OR2X1 U2584 ( .A(\D_cache/n523 ), .B(n2059), .Y(n10167) );
  INVX12 U2585 ( .A(n10167), .Y(mem_addr_D[4]) );
  OR2X1 U2586 ( .A(n8845), .B(n3998), .Y(n10289) );
  INVX12 U2587 ( .A(n10289), .Y(mem_wdata_D[6]) );
  BUFX12 U2588 ( .A(n10224), .Y(mem_wdata_D[71]) );
  NOR2BXL U2589 ( .AN(\D_cache/N145 ), .B(n4006), .Y(n10224) );
  BUFX12 U2590 ( .A(n10226), .Y(mem_wdata_D[69]) );
  NOR2BXL U2591 ( .AN(\D_cache/N147 ), .B(n4006), .Y(n10226) );
  BUFX12 U2592 ( .A(n10214), .Y(mem_wdata_D[81]) );
  NOR2BXL U2593 ( .AN(\D_cache/N135 ), .B(n4007), .Y(n10214) );
  BUFX12 U2594 ( .A(n10217), .Y(mem_wdata_D[78]) );
  NOR2BXL U2595 ( .AN(\D_cache/N138 ), .B(n4007), .Y(n10217) );
  INVX12 U2596 ( .A(n2650), .Y(mem_addr_D[7]) );
  NOR2XL U2597 ( .A(n2703), .B(n4010), .Y(n2651) );
  NOR2XL U2598 ( .A(n8832), .B(n4006), .Y(n2652) );
  NOR2XL U2599 ( .A(n2651), .B(n2652), .Y(n2650) );
  INVX12 U2600 ( .A(n2653), .Y(mem_addr_D[15]) );
  NOR2XL U2601 ( .A(n1085), .B(n4010), .Y(n2654) );
  NOR2XL U2602 ( .A(n8824), .B(n4006), .Y(n2655) );
  NOR2XL U2603 ( .A(n2654), .B(n2655), .Y(n2653) );
  INVX12 U2604 ( .A(n2656), .Y(mem_addr_D[18]) );
  NOR2XL U2605 ( .A(n1620), .B(n4011), .Y(n2657) );
  NOR2XL U2606 ( .A(n8821), .B(n4006), .Y(n2658) );
  NOR2XL U2607 ( .A(n2657), .B(n2658), .Y(n2656) );
  INVX12 U2608 ( .A(n2659), .Y(mem_addr_D[17]) );
  NOR2XL U2609 ( .A(n1625), .B(n4010), .Y(n2660) );
  NOR2XL U2610 ( .A(n8822), .B(n4007), .Y(n2661) );
  NOR2XL U2611 ( .A(n2660), .B(n2661), .Y(n2659) );
  INVX12 U2612 ( .A(n1618), .Y(DCACHE_addr[24]) );
  INVX12 U2613 ( .A(n1619), .Y(DCACHE_addr[21]) );
  INVX12 U2614 ( .A(n1617), .Y(DCACHE_addr[17]) );
  INVX12 U2615 ( .A(n1084), .Y(DCACHE_addr[25]) );
  INVX12 U2616 ( .A(n3037), .Y(DCACHE_addr[10]) );
  INVX12 U2617 ( .A(n1620), .Y(DCACHE_addr[16]) );
  INVX12 U2618 ( .A(n1085), .Y(DCACHE_addr[13]) );
  BUFX12 U2619 ( .A(n10324), .Y(DCACHE_wdata[31]) );
  BUFX12 U2620 ( .A(n10325), .Y(DCACHE_wdata[30]) );
  BUFX12 U2621 ( .A(n10326), .Y(DCACHE_wdata[29]) );
  BUFX12 U2622 ( .A(n10327), .Y(DCACHE_wdata[28]) );
  BUFX12 U2623 ( .A(n10328), .Y(DCACHE_wdata[27]) );
  BUFX12 U2624 ( .A(n10329), .Y(DCACHE_wdata[26]) );
  BUFX12 U2625 ( .A(n10330), .Y(DCACHE_wdata[25]) );
  BUFX12 U2626 ( .A(n10331), .Y(DCACHE_wdata[24]) );
  BUFX12 U2627 ( .A(n10332), .Y(DCACHE_wdata[23]) );
  BUFX12 U2628 ( .A(n10333), .Y(DCACHE_wdata[22]) );
  BUFX12 U2629 ( .A(n10334), .Y(DCACHE_wdata[21]) );
  BUFX12 U2630 ( .A(n10335), .Y(DCACHE_wdata[20]) );
  BUFX12 U2631 ( .A(n10336), .Y(DCACHE_wdata[19]) );
  BUFX12 U2632 ( .A(n10337), .Y(DCACHE_wdata[18]) );
  BUFX12 U2633 ( .A(n10338), .Y(DCACHE_wdata[17]) );
  BUFX12 U2634 ( .A(n10339), .Y(DCACHE_wdata[16]) );
  BUFX12 U2635 ( .A(n10340), .Y(DCACHE_wdata[15]) );
  BUFX12 U2636 ( .A(n10341), .Y(DCACHE_wdata[14]) );
  BUFX12 U2637 ( .A(n10342), .Y(DCACHE_wdata[13]) );
  BUFX12 U2638 ( .A(n10343), .Y(DCACHE_wdata[12]) );
  BUFX12 U2639 ( .A(n10344), .Y(DCACHE_wdata[11]) );
  BUFX12 U2640 ( .A(n10345), .Y(DCACHE_wdata[10]) );
  BUFX12 U2641 ( .A(n10346), .Y(DCACHE_wdata[9]) );
  BUFX12 U2642 ( .A(n10347), .Y(DCACHE_wdata[8]) );
  BUFX12 U2643 ( .A(n10348), .Y(DCACHE_wdata[7]) );
  BUFX12 U2644 ( .A(n10349), .Y(DCACHE_wdata[6]) );
  BUFX12 U2645 ( .A(n10350), .Y(DCACHE_wdata[5]) );
  BUFX12 U2646 ( .A(n10351), .Y(DCACHE_wdata[4]) );
  BUFX12 U2647 ( .A(n10352), .Y(DCACHE_wdata[3]) );
  BUFX12 U2648 ( .A(n10353), .Y(DCACHE_wdata[2]) );
  BUFX12 U2649 ( .A(n10354), .Y(DCACHE_wdata[1]) );
  BUFX12 U2650 ( .A(n10355), .Y(DCACHE_wdata[0]) );
  INVX16 U2651 ( .A(n2701), .Y(DCACHE_addr[1]) );
  NAND2XL U2652 ( .A(n10322), .B(n10323), .Y(\D_cache/n316 ) );
  INVX16 U2653 ( .A(n2703), .Y(DCACHE_addr[5]) );
  XNOR2X1 U2654 ( .A(\i_MIPS/ID_EX[106] ), .B(\i_MIPS/ID_EX[107] ), .Y(
        \i_MIPS/ALU_Control/n18 ) );
  NAND4BX1 U2655 ( .AN(\i_MIPS/ID_EX[106] ), .B(\i_MIPS/ID_EX[105] ), .C(
        \i_MIPS/ID_EX[107] ), .D(\i_MIPS/ALU_Control/n11 ), .Y(
        \i_MIPS/ALU_Control/n20 ) );
  OR2X1 U2656 ( .A(n5035), .B(n3219), .Y(n2705) );
  OR2XL U2657 ( .A(n5034), .B(n3216), .Y(n2706) );
  OR2X1 U2658 ( .A(n8740), .B(n3214), .Y(n2707) );
  MX2XL U2659 ( .A(n5033), .B(n5032), .S0(n4015), .Y(n5034) );
  BUFX8 U2660 ( .A(n6918), .Y(n2708) );
  NAND2X2 U2661 ( .A(n4622), .B(n4728), .Y(n2762) );
  OR2X2 U2662 ( .A(n6597), .B(n3219), .Y(n2709) );
  OR2X1 U2663 ( .A(n6596), .B(n3216), .Y(n2710) );
  NAND3X2 U2664 ( .A(n2709), .B(n2710), .C(n2711), .Y(n7783) );
  CLKINVX4 U2665 ( .A(n8240), .Y(n6597) );
  XOR2X4 U2666 ( .A(n8241), .B(n7783), .Y(n6671) );
  NAND2X4 U2667 ( .A(n8341), .B(n8340), .Y(n7820) );
  INVX12 U2668 ( .A(n2712), .Y(DCACHE_addr[0]) );
  INVXL U2669 ( .A(n8402), .Y(n8403) );
  NAND2BX2 U2670 ( .AN(n6261), .B(n8473), .Y(n6394) );
  NAND2X4 U2671 ( .A(n4662), .B(\i_MIPS/n359 ), .Y(n8482) );
  INVXL U2672 ( .A(n8480), .Y(n6393) );
  OAI221X4 U2673 ( .A0(n3106), .A1(n6395), .B0(n2850), .B1(n3098), .C0(n3096), 
        .Y(n6398) );
  AND2X2 U2674 ( .A(\i_MIPS/IF_ID_1 ), .B(n3596), .Y(n2721) );
  NOR3X4 U2675 ( .A(n2719), .B(n2720), .C(n2721), .Y(n8237) );
  BUFX6 U2676 ( .A(n2828), .Y(n3596) );
  OAI221X1 U2677 ( .A0(\D_cache/n164 ), .A1(n8852), .B0(n3074), .B1(n8833), 
        .C0(\D_cache/n190 ), .Y(DCACHE_rdata[18]) );
  OAI221X1 U2678 ( .A0(\D_cache/n164 ), .A1(n8861), .B0(n3074), .B1(n8842), 
        .C0(\D_cache/n166 ), .Y(DCACHE_rdata[9]) );
  CLKBUFX3 U2679 ( .A(n3105), .Y(n3101) );
  CLKBUFX2 U2680 ( .A(n3485), .Y(n3461) );
  CLKBUFX2 U2681 ( .A(n3437), .Y(n3413) );
  INVXL U2682 ( .A(n4641), .Y(n4699) );
  BUFX12 U2683 ( .A(n8421), .Y(n3598) );
  CLKBUFX3 U2684 ( .A(n7069), .Y(n3215) );
  CLKBUFX3 U2685 ( .A(n3309), .Y(n3303) );
  NAND2X1 U2686 ( .A(n4632), .B(\i_MIPS/n349 ), .Y(n6694) );
  OA22XL U2687 ( .A0(\i_MIPS/Register/register[6][12] ), .A1(n3172), .B0(
        \i_MIPS/Register/register[14][12] ), .B1(n3169), .Y(n6298) );
  AND2X2 U2688 ( .A(n3094), .B(\i_MIPS/ALUin1[26] ), .Y(n2896) );
  NOR2XL U2689 ( .A(\i_MIPS/PC/n28 ), .B(n3611), .Y(n2737) );
  OA22XL U2690 ( .A0(\i_MIPS/Register/register[22][0] ), .A1(n3170), .B0(
        \i_MIPS/Register/register[30][0] ), .B1(n3168), .Y(n5093) );
  NAND2X4 U2691 ( .A(n2886), .B(n4019), .Y(n2732) );
  OA22XL U2692 ( .A0(\i_MIPS/Register/register[6][0] ), .A1(n3116), .B0(
        \i_MIPS/Register/register[14][0] ), .B1(n3113), .Y(n5063) );
  OA22XL U2693 ( .A0(\i_MIPS/Register/register[16][0] ), .A1(n3186), .B0(
        \i_MIPS/Register/register[24][0] ), .B1(n3182), .Y(n5099) );
  OA22XL U2694 ( .A0(n3477), .A1(n535), .B0(n3430), .B1(n1454), .Y(n7720) );
  OA22XL U2695 ( .A0(\i_MIPS/Register/register[22][23] ), .A1(n3170), .B0(
        \i_MIPS/Register/register[30][23] ), .B1(n3169), .Y(n6867) );
  AND2XL U2696 ( .A(n5036), .B(\i_MIPS/n371 ), .Y(n5037) );
  AO21X4 U2697 ( .A0(n8388), .A1(n8387), .B0(n8382), .Y(n8348) );
  OA22X1 U2698 ( .A0(n3387), .A1(n464), .B0(n3345), .B1(n1379), .Y(n7747) );
  OR3X2 U2699 ( .A(n2735), .B(n2736), .C(n2737), .Y(n8184) );
  NAND3BX2 U2700 ( .AN(n8184), .B(n8183), .C(n8182), .Y(\i_MIPS/PC/n60 ) );
  XOR2X2 U2701 ( .A(n8305), .B(ICACHE_addr[27]), .Y(n8301) );
  NAND3X4 U2702 ( .A(ICACHE_addr[20]), .B(ICACHE_addr[19]), .C(n8080), .Y(
        n8120) );
  INVX12 U2703 ( .A(n8722), .Y(DCACHE_addr[26]) );
  CLKBUFX2 U2704 ( .A(n3109), .Y(n3108) );
  CLKBUFX2 U2705 ( .A(n3485), .Y(n3454) );
  CLKBUFX2 U2706 ( .A(n3439), .Y(n3410) );
  AND2XL U2707 ( .A(n6682), .B(n5480), .Y(n2813) );
  AO22XL U2708 ( .A0(n2881), .A1(n6617), .B0(n2818), .B1(n6618), .Y(n5129) );
  INVX1 U2709 ( .A(n7850), .Y(n7849) );
  CLKBUFX2 U2710 ( .A(n2863), .Y(n3083) );
  INVX1 U2711 ( .A(n8522), .Y(n8523) );
  AO21X1 U2712 ( .A0(n8521), .A1(n8520), .B0(n8519), .Y(n8908) );
  NAND2X4 U2713 ( .A(n5390), .B(n4971), .Y(n4679) );
  OR2XL U2714 ( .A(\i_MIPS/PC/n17 ), .B(n8457), .Y(n2743) );
  OR2XL U2715 ( .A(n8254), .B(n17), .Y(n2742) );
  NAND2X2 U2716 ( .A(\i_MIPS/ALUin1[22] ), .B(n4633), .Y(n6693) );
  AND2X1 U2717 ( .A(n3089), .B(\i_MIPS/ALUin1[26] ), .Y(n2897) );
  AO22X1 U2718 ( .A0(\i_MIPS/control_out[7] ), .A1(n3610), .B0(
        \i_MIPS/ALUOp[1] ), .B1(n8552), .Y(\i_MIPS/n471 ) );
  OA22XL U2719 ( .A0(n3550), .A1(n536), .B0(n3509), .B1(n1455), .Y(n4559) );
  NOR2X1 U2720 ( .A(n8178), .B(n3049), .Y(n2735) );
  CLKBUFX2 U2721 ( .A(n3575), .Y(n3567) );
  CLKINVX3 U2722 ( .A(n8233), .Y(n6669) );
  INVX3 U2723 ( .A(n4676), .Y(n5185) );
  MX2XL U2724 ( .A(n3072), .B(n2865), .S0(n6391), .Y(n6271) );
  XOR3XL U2725 ( .A(n7968), .B(n2806), .C(n7967), .Y(n7959) );
  OR2X4 U2726 ( .A(n6844), .B(n6843), .Y(n2745) );
  INVX1 U2727 ( .A(n3028), .Y(n8254) );
  OAI31X4 U2728 ( .A0(n4616), .A1(\i_MIPS/ID_EX[73] ), .A2(n4615), .B0(n4614), 
        .Y(n4727) );
  OA22X1 U2729 ( .A0(\i_MIPS/Register/register[20][0] ), .A1(n3179), .B0(
        \i_MIPS/Register/register[28][0] ), .B1(n3177), .Y(n5100) );
  OA22X1 U2730 ( .A0(\i_MIPS/Register/register[4][12] ), .A1(n3179), .B0(
        \i_MIPS/Register/register[12][12] ), .B1(n3178), .Y(n6305) );
  OA22X1 U2731 ( .A0(\i_MIPS/Register/register[20][23] ), .A1(n3181), .B0(
        \i_MIPS/Register/register[28][23] ), .B1(n3178), .Y(n6874) );
  OA22X1 U2732 ( .A0(\i_MIPS/Register/register[16][23] ), .A1(n3187), .B0(
        \i_MIPS/Register/register[24][23] ), .B1(n3182), .Y(n6873) );
  OR2X2 U2733 ( .A(n6669), .B(n3219), .Y(n2738) );
  OR2X1 U2734 ( .A(n6668), .B(n3216), .Y(n2739) );
  NAND3X2 U2735 ( .A(n2738), .B(n2739), .C(n2740), .Y(n7734) );
  CLKMX2X2 U2736 ( .A(n2717), .B(n7734), .S0(n3623), .Y(\i_MIPS/n433 ) );
  AND2X2 U2737 ( .A(\i_MIPS/ALU_Control/n15 ), .B(\i_MIPS/ALUOp[1] ), .Y(n4614) );
  NAND2XL U2738 ( .A(n6680), .B(n4016), .Y(n6845) );
  NAND3XL U2739 ( .A(n8716), .B(n8913), .C(n2838), .Y(n8924) );
  NAND2X8 U2740 ( .A(n2832), .B(n2708), .Y(n6544) );
  AND2X1 U2741 ( .A(n6617), .B(n4017), .Y(n2811) );
  INVXL U2742 ( .A(n5254), .Y(n5610) );
  CLKBUFX2 U2743 ( .A(n3324), .Y(n3348) );
  NAND2X2 U2744 ( .A(n10300), .B(n2751), .Y(n2753) );
  CLKINVX1 U2745 ( .A(n4660), .Y(n4644) );
  OA22XL U2746 ( .A0(n3386), .A1(n537), .B0(n3344), .B1(n1456), .Y(n7737) );
  OA22XL U2747 ( .A0(n3563), .A1(n538), .B0(n3521), .B1(n1457), .Y(n7735) );
  INVX1 U2748 ( .A(n6673), .Y(n6674) );
  INVX1 U2749 ( .A(n7866), .Y(n7863) );
  INVX1 U2750 ( .A(n7895), .Y(n7899) );
  NAND2X1 U2751 ( .A(\i_MIPS/ALUin1[23] ), .B(n4634), .Y(n6841) );
  OR2XL U2752 ( .A(n3070), .B(n6841), .Y(n2746) );
  INVXL U2753 ( .A(n6836), .Y(n6846) );
  AND2XL U2754 ( .A(n6837), .B(n6841), .Y(n6844) );
  MX2X4 U2755 ( .A(\i_MIPS/n281 ), .B(n2994), .S0(n4018), .Y(n4654) );
  CLKBUFX4 U2756 ( .A(n3095), .Y(n3096) );
  BUFX2 U2757 ( .A(n3481), .Y(n3473) );
  AOI21X1 U2758 ( .A0(n5674), .A1(n8540), .B0(n5047), .Y(n2815) );
  NAND2X1 U2759 ( .A(n6682), .B(n5970), .Y(n6908) );
  CLKINVX1 U2760 ( .A(n8517), .Y(n8521) );
  INVXL U2761 ( .A(n5481), .Y(n5115) );
  OAI211X1 U2762 ( .A0(n6334), .A1(n5616), .B0(n5615), .C0(n5614), .Y(n6546)
         );
  CLKBUFX2 U2763 ( .A(n2863), .Y(n3084) );
  OAI222X2 U2764 ( .A0(n5956), .A1(n3164), .B0(n5934), .B1(n2761), .C0(n8721), 
        .C1(n3163), .Y(n8275) );
  NAND3BX1 U2765 ( .AN(n8479), .B(n8478), .C(n8477), .Y(n8483) );
  AND2X2 U2766 ( .A(n8), .B(n54), .Y(n2864) );
  INVX2 U2767 ( .A(n4706), .Y(n6992) );
  INVX1 U2768 ( .A(n4623), .Y(n4705) );
  INVX1 U2769 ( .A(n8478), .Y(n5534) );
  CLKBUFX2 U2770 ( .A(n2907), .Y(n3089) );
  OA22X1 U2771 ( .A0(n3564), .A1(n465), .B0(n3522), .B1(n1380), .Y(n7745) );
  OA22X1 U2772 ( .A0(n3462), .A1(n144), .B0(n3441), .B1(n1035), .Y(n4473) );
  NAND2X1 U2773 ( .A(\i_MIPS/ALUin1[26] ), .B(n4629), .Y(n8461) );
  CLKAND2X3 U2774 ( .A(\i_MIPS/Sign_Extend_ID[31] ), .B(n3627), .Y(n2804) );
  OA22X1 U2775 ( .A0(n3478), .A1(n466), .B0(n3431), .B1(n1381), .Y(n7746) );
  OA22X1 U2776 ( .A0(\i_MIPS/Register/register[0][12] ), .A1(n3187), .B0(
        \i_MIPS/Register/register[8][12] ), .B1(n3184), .Y(n6304) );
  NOR2X8 U2777 ( .A(\D_cache/n520 ), .B(n1074), .Y(\D_cache/n200 ) );
  INVX1 U2778 ( .A(n6124), .Y(n5967) );
  NAND2X8 U2779 ( .A(n4912), .B(n2708), .Y(n6550) );
  INVXL U2780 ( .A(n6677), .Y(n6683) );
  CLKBUFX2 U2781 ( .A(n3575), .Y(n3566) );
  OAI221X1 U2782 ( .A0(n3106), .A1(n5988), .B0(n2846), .B1(n3098), .C0(n3097), 
        .Y(n5992) );
  NAND3BX1 U2783 ( .AN(n4665), .B(n4664), .C(n4663), .Y(n4830) );
  CLKINVX3 U2784 ( .A(n5672), .Y(n4589) );
  NAND2X1 U2785 ( .A(n2812), .B(n4827), .Y(n4599) );
  NAND2X4 U2786 ( .A(n4664), .B(n4656), .Y(n4829) );
  INVX1 U2787 ( .A(n4827), .Y(n8538) );
  INVX1 U2788 ( .A(n5265), .Y(n5611) );
  INVX12 U2789 ( .A(n3070), .Y(n6993) );
  INVX1 U2790 ( .A(n5259), .Y(n5196) );
  OAI211X2 U2791 ( .A0(n4591), .A1(n4592), .B0(n8509), .C0(n8506), .Y(n5190)
         );
  INVXL U2792 ( .A(n5616), .Y(n5267) );
  INVX1 U2793 ( .A(n6332), .Y(n5754) );
  MX2XL U2794 ( .A(n6836), .B(n5266), .S0(n55), .Y(n6773) );
  CLKBUFX2 U2795 ( .A(n3309), .Y(n3302) );
  CLKBUFX3 U2796 ( .A(n3397), .Y(n3390) );
  BUFX2 U2797 ( .A(n3974), .Y(n3973) );
  MX2XL U2798 ( .A(n5973), .B(n5972), .S0(n4016), .Y(n6141) );
  OAI2BB1X4 U2799 ( .A0N(n5905), .A1N(n5893), .B0(n5890), .Y(n5811) );
  OAI2BB1X1 U2800 ( .A0N(n8511), .A1N(n8510), .B0(n8509), .Y(n8905) );
  AND2X2 U2801 ( .A(n5483), .B(n5970), .Y(n2832) );
  INVX3 U2802 ( .A(n4636), .Y(n4634) );
  INVX1 U2803 ( .A(n8543), .Y(n8546) );
  AND2X4 U2804 ( .A(n5981), .B(n8545), .Y(n2833) );
  OAI221X1 U2805 ( .A0(\i_MIPS/n347 ), .A1(n3091), .B0(\i_MIPS/n348 ), .B1(
        n3085), .C0(n5113), .Y(n5383) );
  CLKBUFX2 U2806 ( .A(n2907), .Y(n3090) );
  OA22XL U2807 ( .A0(n3383), .A1(n539), .B0(n3341), .B1(n1458), .Y(n7601) );
  OA22XL U2808 ( .A0(n3560), .A1(n540), .B0(n3518), .B1(n1459), .Y(n7599) );
  INVX1 U2809 ( .A(n7914), .Y(n7909) );
  MX2XL U2810 ( .A(n5963), .B(n5962), .S0(n4016), .Y(n5902) );
  INVXL U2811 ( .A(n5462), .Y(n5824) );
  OA22XL U2812 ( .A0(n3387), .A1(n541), .B0(n3345), .B1(n1460), .Y(n7752) );
  OA22XL U2813 ( .A0(n3300), .A1(n542), .B0(n3253), .B1(n1461), .Y(n7753) );
  OA22XL U2814 ( .A0(n3564), .A1(n543), .B0(n3522), .B1(n1462), .Y(n7750) );
  OA22XL U2815 ( .A0(n3300), .A1(n544), .B0(n3253), .B1(n1463), .Y(n7748) );
  OA22XL U2816 ( .A0(n3299), .A1(n545), .B0(n3252), .B1(n1464), .Y(n7738) );
  XOR2X1 U2817 ( .A(\i_MIPS/IR_ID[19] ), .B(n2890), .Y(n4775) );
  NAND2X2 U2818 ( .A(\i_MIPS/ALUin1[7] ), .B(n4673), .Y(n8510) );
  NAND2XL U2819 ( .A(\i_MIPS/ALUin1[24] ), .B(n4635), .Y(n5469) );
  AND2XL U2820 ( .A(n3090), .B(\i_MIPS/ALUin1[27] ), .Y(n2895) );
  AND2X1 U2821 ( .A(\i_MIPS/IR_ID[18] ), .B(\i_MIPS/n318 ), .Y(n2973) );
  OA22XL U2822 ( .A0(\i_MIPS/Register/register[20][12] ), .A1(n3181), .B0(
        \i_MIPS/Register/register[28][12] ), .B1(n3178), .Y(n6314) );
  OA22X1 U2823 ( .A0(\i_MIPS/Register/register[16][12] ), .A1(n3187), .B0(
        \i_MIPS/Register/register[24][12] ), .B1(n3184), .Y(n6313) );
  NAND2X1 U2824 ( .A(\i_MIPS/ALUin1[19] ), .B(n4660), .Y(n8537) );
  AO21XL U2825 ( .A0(n3080), .A1(\i_MIPS/ALUin1[29] ), .B0(n2903), .Y(n5122)
         );
  AND2X2 U2826 ( .A(\i_MIPS/IR_ID[24] ), .B(\i_MIPS/n230 ), .Y(n2977) );
  OA22XL U2827 ( .A0(\i_MIPS/Register/register[22][4] ), .A1(n3171), .B0(
        \i_MIPS/Register/register[30][4] ), .B1(n3167), .Y(n5367) );
  OA22XL U2828 ( .A0(\i_MIPS/Register/register[22][18] ), .A1(n3172), .B0(
        \i_MIPS/Register/register[30][18] ), .B1(n3168), .Y(n5791) );
  OA22XL U2829 ( .A0(\i_MIPS/Register/register[20][0] ), .A1(n3128), .B0(
        \i_MIPS/Register/register[28][0] ), .B1(n3125), .Y(n5079) );
  OA22XL U2830 ( .A0(\i_MIPS/Register/register[16][0] ), .A1(n3134), .B0(
        \i_MIPS/Register/register[24][0] ), .B1(n3131), .Y(n5078) );
  OA22XL U2831 ( .A0(\i_MIPS/Register/register[20][4] ), .A1(n3180), .B0(
        \i_MIPS/Register/register[28][4] ), .B1(n3176), .Y(n5374) );
  OA22XL U2832 ( .A0(\i_MIPS/Register/register[4][0] ), .A1(n3128), .B0(
        \i_MIPS/Register/register[12][0] ), .B1(n3125), .Y(n5070) );
  OA22XL U2833 ( .A0(\i_MIPS/Register/register[20][18] ), .A1(n3181), .B0(
        \i_MIPS/Register/register[28][18] ), .B1(n3177), .Y(n5798) );
  OA22XL U2834 ( .A0(\i_MIPS/Register/register[16][4] ), .A1(n3185), .B0(
        \i_MIPS/Register/register[24][4] ), .B1(n3182), .Y(n5373) );
  OA22XL U2835 ( .A0(\i_MIPS/Register/register[0][0] ), .A1(n3134), .B0(
        \i_MIPS/Register/register[8][0] ), .B1(n3131), .Y(n5069) );
  OA22XL U2836 ( .A0(\i_MIPS/Register/register[16][18] ), .A1(n3186), .B0(
        \i_MIPS/Register/register[24][18] ), .B1(n3183), .Y(n5797) );
  OA22XL U2837 ( .A0(n3477), .A1(n546), .B0(n3430), .B1(n1465), .Y(n7736) );
  MX2XL U2838 ( .A(\i_MIPS/ID_EX[59] ), .B(n7810), .S0(n3626), .Y(
        \i_MIPS/n401 ) );
  INVX12 U2839 ( .A(n1616), .Y(DCACHE_addr[28]) );
  CLKBUFX3 U2840 ( .A(n3586), .Y(n3592) );
  INVX1 U2841 ( .A(n6910), .Y(n6912) );
  CLKINVX1 U2842 ( .A(n3955), .Y(n2757) );
  INVXL U2843 ( .A(n6054), .Y(n6055) );
  CLKINVX6 U2844 ( .A(n4029), .Y(n4025) );
  AO21X4 U2845 ( .A0(n5977), .A1(n5976), .B0(n5975), .Y(n6466) );
  INVX3 U2846 ( .A(n7932), .Y(n7931) );
  AND3XL U2847 ( .A(n5739), .B(n4829), .C(n5734), .Y(n4832) );
  INVX1 U2848 ( .A(n8143), .Y(n8147) );
  AOI211X2 U2849 ( .A0(n2833), .A1(n5978), .B0(n8544), .C0(n2845), .Y(n4602)
         );
  AO22X1 U2850 ( .A0(n5196), .A1(n2869), .B0(n3111), .B1(n5257), .Y(n5198) );
  CLKBUFX3 U2851 ( .A(n3486), .Y(n3484) );
  CLKBUFX3 U2852 ( .A(n3440), .Y(n3438) );
  CLKINVX12 U2853 ( .A(n2865), .Y(n7005) );
  MX2XL U2854 ( .A(n7005), .B(n3071), .S0(n6672), .Y(n6704) );
  NAND2X8 U2855 ( .A(n4537), .B(n4538), .Y(n8426) );
  MX2XL U2856 ( .A(n3072), .B(n2865), .S0(n4987), .Y(n4988) );
  NAND2XL U2857 ( .A(n7069), .B(n3219), .Y(n2760) );
  INVX3 U2858 ( .A(n8012), .Y(n5253) );
  NAND2BXL U2859 ( .AN(n3576), .B(n8567), .Y(n7581) );
  NAND2X2 U2860 ( .A(n6905), .B(n1082), .Y(n6996) );
  AO21X1 U2861 ( .A0(n5604), .A1(n5621), .B0(n5618), .Y(n4834) );
  AO21X4 U2862 ( .A0(n6691), .A1(n6690), .B0(n6689), .Y(n6692) );
  AND2X1 U2863 ( .A(n4833), .B(n4666), .Y(n4698) );
  AOI21X1 U2864 ( .A0(n7011), .A1(n5754), .B0(n5753), .Y(n2826) );
  CLKBUFX3 U2865 ( .A(n7046), .Y(n3163) );
  CLKINVX3 U2866 ( .A(n6849), .Y(n4912) );
  CLKINVX1 U2867 ( .A(n8462), .Y(n8463) );
  NAND3BX1 U2868 ( .AN(n8912), .B(n2842), .C(n8463), .Y(n8464) );
  AO21XL U2869 ( .A0(n6601), .A1(n6621), .B0(n6608), .Y(n6536) );
  INVXL U2870 ( .A(n6761), .Y(n6764) );
  BUFX2 U2871 ( .A(n3662), .Y(n3015) );
  INVX1 U2872 ( .A(n7002), .Y(n7003) );
  CLKBUFX3 U2873 ( .A(n3975), .Y(n3972) );
  CLKBUFX3 U2874 ( .A(n3219), .Y(n3218) );
  MX2X2 U2875 ( .A(DCACHE_addr[8]), .B(DCACHE_rdata[10]), .S0(n4023), .Y(n3031) );
  AO21X4 U2876 ( .A0(n8322), .A1(n8304), .B0(n8303), .Y(n2765) );
  OAI2BB1X1 U2877 ( .A0N(n6190), .A1N(n6189), .B0(n6188), .Y(n6193) );
  BUFX8 U2878 ( .A(n7004), .Y(n3071) );
  NAND2BXL U2879 ( .AN(n3000), .B(n8624), .Y(n7780) );
  NAND2BXL U2880 ( .AN(n2163), .B(n8656), .Y(n7781) );
  NAND2BXL U2881 ( .AN(n3001), .B(n8592), .Y(n7778) );
  NAND2BXL U2882 ( .AN(n3000), .B(n8628), .Y(n7684) );
  NAND2BXL U2883 ( .AN(n2163), .B(n8660), .Y(n7685) );
  NAND2BXL U2884 ( .AN(n3001), .B(n8596), .Y(n7682) );
  NAND2BXL U2885 ( .AN(n3000), .B(n8630), .Y(n7630) );
  NAND2BXL U2886 ( .AN(n2163), .B(n8662), .Y(n7631) );
  NAND2BXL U2887 ( .AN(n3001), .B(n8598), .Y(n7628) );
  NAND2BXL U2888 ( .AN(n3000), .B(n8632), .Y(n7533) );
  NAND2BXL U2889 ( .AN(n2163), .B(n8664), .Y(n7534) );
  NAND2BXL U2890 ( .AN(n3001), .B(n8600), .Y(n7531) );
  NAND2BXL U2891 ( .AN(n3000), .B(n8626), .Y(n7730) );
  NAND2BXL U2892 ( .AN(n3000), .B(n8627), .Y(n7707) );
  NAND2BXL U2893 ( .AN(n2163), .B(n8659), .Y(n7708) );
  NAND2BXL U2894 ( .AN(n3001), .B(n8595), .Y(n7705) );
  INVX3 U2895 ( .A(n5193), .Y(n4596) );
  CLKINVX3 U2896 ( .A(n8123), .Y(n8125) );
  AOI211X1 U2897 ( .A0(n5402), .A1(n4919), .B0(n4918), .C0(n4917), .Y(n4920)
         );
  INVXL U2898 ( .A(n7841), .Y(n7839) );
  AOI211X1 U2899 ( .A0(n5402), .A1(n5401), .B0(n5400), .C0(n5399), .Y(n5403)
         );
  OAI2BB1X1 U2900 ( .A0N(n8508), .A1N(n8507), .B0(n8506), .Y(n8511) );
  AOI2BB1X4 U2901 ( .A0N(n6060), .A1N(n5471), .B0(n4700), .Y(n4702) );
  NAND2X6 U2902 ( .A(n6061), .B(n6065), .Y(n4700) );
  AND2XL U2903 ( .A(\D_cache/n203 ), .B(\D_cache/n200 ), .Y(n3033) );
  NAND2X1 U2904 ( .A(n4629), .B(\i_MIPS/n345 ), .Y(n6065) );
  OAI222XL U2905 ( .A0(n6334), .A1(n6333), .B0(n6332), .B1(n6619), .C0(n3076), 
        .C1(n6679), .Y(n7008) );
  AND2X2 U2906 ( .A(n8520), .B(n8461), .Y(n2842) );
  NAND2X1 U2907 ( .A(n4654), .B(\i_MIPS/n357 ), .Y(n6339) );
  MX2XL U2908 ( .A(n5268), .B(n5611), .S0(n4016), .Y(n5547) );
  NAND2X1 U2909 ( .A(n4634), .B(\i_MIPS/n348 ), .Y(n6834) );
  NAND2X1 U2910 ( .A(n3076), .B(\i_MIPS/n340 ), .Y(n5964) );
  INVX6 U2911 ( .A(\i_MIPS/n320 ), .Y(n4015) );
  OA22X1 U2912 ( .A0(n3296), .A1(n467), .B0(n3249), .B1(n1382), .Y(n7597) );
  OA22X1 U2913 ( .A0(n3560), .A1(n468), .B0(n3518), .B1(n1383), .Y(n7594) );
  OA22X1 U2914 ( .A0(n3383), .A1(n469), .B0(n3341), .B1(n1384), .Y(n7596) );
  NAND2BXL U2915 ( .AN(n3000), .B(n8637), .Y(n7138) );
  NAND2BXL U2916 ( .AN(n3000), .B(n8636), .Y(n7162) );
  NAND2BXL U2917 ( .AN(n3000), .B(n8634), .Y(n7114) );
  NAND2BXL U2918 ( .AN(n3001), .B(n8609), .Y(n7459) );
  NAND2BXL U2919 ( .AN(n3001), .B(n8610), .Y(n7435) );
  NAND2BXL U2920 ( .AN(n3001), .B(n8608), .Y(n8134) );
  OA22X1 U2921 ( .A0(n3553), .A1(n470), .B0(n3511), .B1(n1385), .Y(n7335) );
  NAND2BXL U2922 ( .AN(n3576), .B(n8581), .Y(n7210) );
  NAND2BX1 U2923 ( .AN(n3576), .B(n8580), .Y(n7186) );
  NAND4X1 U2924 ( .A(n7188), .B(n7187), .C(n7186), .D(n7185), .Y(n7797) );
  INVXL U2925 ( .A(n6675), .Y(n6052) );
  NAND4X1 U2926 ( .A(n7553), .B(n7552), .C(n7551), .D(n7550), .Y(n8601) );
  AOI22XL U2927 ( .A0(\D_cache/N141 ), .A1(n2153), .B0(n3032), .B1(
        \D_cache/N173 ), .Y(\D_cache/n197 ) );
  XOR2X4 U2928 ( .A(n8703), .B(ICACHE_addr[20]), .Y(n4411) );
  XOR2X4 U2929 ( .A(n8689), .B(ICACHE_addr[6]), .Y(n4412) );
  XOR2X4 U2930 ( .A(n8702), .B(ICACHE_addr[19]), .Y(n4401) );
  INVXL U2931 ( .A(\i_MIPS/forward_unit/n15 ), .Y(n4779) );
  CLKMX2X3 U2932 ( .A(\i_MIPS/n285 ), .B(n2992), .S0(n4018), .Y(n4652) );
  NAND3XL U2933 ( .A(\i_MIPS/ALU_Control/n11 ), .B(\i_MIPS/n323 ), .C(
        \i_MIPS/ALU_Control/n18 ), .Y(\i_MIPS/ALU_Control/n15 ) );
  NAND3BXL U2934 ( .AN(\i_MIPS/ID_EX[76] ), .B(n1083), .C(n2888), .Y(n4616) );
  CLKMX2X2 U2935 ( .A(n2966), .B(n2967), .S0(DCACHE_addr[4]), .Y(
        \D_cache/N134 ) );
  OA22X1 U2936 ( .A0(\i_MIPS/Register/register[20][22] ), .A1(n3128), .B0(
        \i_MIPS/Register/register[28][22] ), .B1(n3126), .Y(n6742) );
  BUFX16 U2937 ( .A(n7828), .Y(n3073) );
  OA22X1 U2938 ( .A0(\i_MIPS/Register/register[4][4] ), .A1(n3180), .B0(
        \i_MIPS/Register/register[12][4] ), .B1(n3176), .Y(n5365) );
  NOR2X1 U2939 ( .A(\i_MIPS/Reg_W[4] ), .B(\i_MIPS/Reg_W[3] ), .Y(
        \i_MIPS/forward_unit/n25 ) );
  MX2X1 U2940 ( .A(n1881), .B(n3036), .S0(n3626), .Y(\i_MIPS/n429 ) );
  XOR2X1 U2941 ( .A(n8040), .B(ICACHE_addr[17]), .Y(n8042) );
  MXI2XL U2942 ( .A(n2992), .B(\i_MIPS/n224 ), .S0(n3623), .Y(\i_MIPS/n500 )
         );
  MXI2XL U2943 ( .A(\i_MIPS/n284 ), .B(\i_MIPS/n285 ), .S0(n3621), .Y(
        \i_MIPS/n412 ) );
  MXI2XL U2944 ( .A(\i_MIPS/n288 ), .B(\i_MIPS/n289 ), .S0(n3619), .Y(
        \i_MIPS/n416 ) );
  OA22X1 U2945 ( .A0(n3474), .A1(n471), .B0(n3427), .B1(n1386), .Y(n7595) );
  OA22X1 U2946 ( .A0(n3472), .A1(n1373), .B0(n3425), .B1(n447), .Y(n7541) );
  NAND2BX1 U2947 ( .AN(DCACHE_ren), .B(\i_MIPS/n310 ), .Y(n2801) );
  CLKINVX1 U2948 ( .A(n2801), .Y(\D_cache/n214 ) );
  OR2XL U2949 ( .A(n5802), .B(n3217), .Y(n2755) );
  CLKINVX3 U2950 ( .A(n3630), .Y(n3625) );
  CLKINVX3 U2951 ( .A(n3630), .Y(n3626) );
  CLKINVX3 U2952 ( .A(n3630), .Y(n3623) );
  CLKINVX3 U2953 ( .A(n3630), .Y(n3624) );
  BUFX2 U2954 ( .A(n3616), .Y(n3630) );
  CLKINVX2 U2955 ( .A(n3551), .Y(n3540) );
  CLKINVX2 U2956 ( .A(n3341), .Y(n3318) );
  CLKINVX3 U2957 ( .A(n3551), .Y(n3539) );
  CLKINVX3 U2958 ( .A(n3322), .Y(n3316) );
  CLKINVX3 U2959 ( .A(n3552), .Y(n3541) );
  CLKINVX3 U2960 ( .A(n3320), .Y(n3319) );
  BUFX2 U2961 ( .A(n3352), .Y(n3321) );
  NAND2XL U2962 ( .A(n8684), .B(n8807), .Y(n8552) );
  INVX1 U2963 ( .A(n7911), .Y(n7912) );
  INVXL U2964 ( .A(n6612), .Y(n5130) );
  CLKBUFX2 U2965 ( .A(n3112), .Y(n3110) );
  CLKBUFX2 U2966 ( .A(n3112), .Y(n3111) );
  CLKINVX2 U2967 ( .A(n3380), .Y(n3361) );
  CLKINVX2 U2968 ( .A(n3244), .Y(n3228) );
  CLKINVX2 U2969 ( .A(n3276), .Y(n3273) );
  CLKINVX3 U2970 ( .A(n3365), .Y(n3359) );
  CLKINVX3 U2971 ( .A(n3242), .Y(n3226) );
  CLKINVX3 U2972 ( .A(n3277), .Y(n3272) );
  CLKINVX3 U2973 ( .A(n3280), .Y(n3269) );
  CLKINVX3 U2974 ( .A(n3246), .Y(n3224) );
  CLKINVX3 U2975 ( .A(n3279), .Y(n3270) );
  CLKINVX3 U2976 ( .A(n3230), .Y(n3229) );
  CLKINVX3 U2977 ( .A(n3275), .Y(n3274) );
  CLKINVX3 U2978 ( .A(n3363), .Y(n3362) );
  CLKINVX2 U2979 ( .A(n3521), .Y(n3496) );
  CLKINVX3 U2980 ( .A(n3499), .Y(n3494) );
  CLKINVX3 U2981 ( .A(n3518), .Y(n3497) );
  INVX3 U2982 ( .A(n8087), .Y(n8089) );
  BUFX2 U2983 ( .A(n2766), .Y(n3352) );
  MX2XL U2984 ( .A(n2865), .B(n3072), .S0(n5682), .Y(n5683) );
  NAND2X2 U2985 ( .A(n6617), .B(n4016), .Y(n6125) );
  CLKINVX8 U2986 ( .A(n7001), .Y(n6680) );
  BUFX2 U2987 ( .A(n3573), .Y(n3572) );
  AO22XL U2988 ( .A0(n6680), .A1(n6054), .B0(n2817), .B1(n6990), .Y(n5751) );
  AO22XL U2989 ( .A0(n5736), .A1(n3102), .B0(n3110), .B1(n5737), .Y(n5742) );
  CLKBUFX2 U2990 ( .A(n3485), .Y(n3453) );
  CLKBUFX2 U2991 ( .A(n3485), .Y(n3460) );
  CLKBUFX2 U2992 ( .A(n3439), .Y(n3409) );
  BUFX2 U2993 ( .A(n3395), .Y(n3364) );
  BUFX2 U2994 ( .A(n3262), .Y(n3231) );
  BUFX2 U2995 ( .A(n3529), .Y(n3498) );
  MX2XL U2996 ( .A(n2865), .B(n3072), .S0(n5749), .Y(n5750) );
  INVXL U2997 ( .A(n3068), .Y(n5609) );
  INVX1 U2998 ( .A(n6919), .Y(n5054) );
  INVXL U2999 ( .A(n6050), .Y(n6051) );
  CLKBUFX2 U3000 ( .A(n3352), .Y(n3350) );
  CLKBUFX2 U3001 ( .A(n3574), .Y(n3569) );
  INVXL U3002 ( .A(n6828), .Y(n6833) );
  INVXL U3003 ( .A(n6756), .Y(n6760) );
  CLKBUFX2 U3004 ( .A(n3482), .Y(n3470) );
  CLKBUFX2 U3005 ( .A(n3482), .Y(n3471) );
  CLKBUFX2 U3006 ( .A(n3481), .Y(n3475) );
  CLKBUFX2 U3007 ( .A(n3481), .Y(n3474) );
  CLKBUFX2 U3008 ( .A(n3525), .Y(n3517) );
  CLKBUFX2 U3009 ( .A(n3257), .Y(n3245) );
  CLKBUFX2 U3010 ( .A(n3257), .Y(n3246) );
  CLKBUFX2 U3011 ( .A(n3526), .Y(n3514) );
  CLKBUFX2 U3012 ( .A(n3526), .Y(n3515) );
  CLKBUFX2 U3013 ( .A(n3525), .Y(n3519) );
  CLKBUFX2 U3014 ( .A(n3525), .Y(n3518) );
  CLKBUFX2 U3015 ( .A(n3350), .Y(n3347) );
  CLKBUFX2 U3016 ( .A(n3574), .Y(n3570) );
  CLKBUFX2 U3017 ( .A(n3439), .Y(n3408) );
  NAND3X1 U3018 ( .A(n2206), .B(n2127), .C(n3066), .Y(\D_cache/n206 ) );
  INVX3 U3019 ( .A(n7951), .Y(n7953) );
  CLKINVX3 U3020 ( .A(n8249), .Y(n6454) );
  INVX3 U3021 ( .A(n8348), .Y(n7873) );
  MX2XL U3022 ( .A(n3072), .B(n2865), .S0(n5398), .Y(n5399) );
  OAI221X2 U3023 ( .A0(n8064), .A1(n8063), .B0(n8066), .B1(n3577), .C0(n8062), 
        .Y(n8081) );
  XOR2X2 U3024 ( .A(n8199), .B(n8166), .Y(n6976) );
  OAI211X2 U3025 ( .A0(n8024), .A1(n8023), .B0(n8022), .C0(n8021), .Y(n8058)
         );
  INVX3 U3026 ( .A(n8020), .Y(n8024) );
  NAND4BX2 U3027 ( .AN(n4845), .B(n4844), .C(n4843), .D(n4842), .Y(n8223) );
  NAND4BX2 U3028 ( .AN(n5838), .B(n5837), .C(n5836), .D(n5835), .Y(n8284) );
  NAND3BXL U3029 ( .AN(n5812), .B(n5832), .C(n3109), .Y(n5837) );
  NAND4X2 U3030 ( .A(n6928), .B(n6927), .C(n6926), .D(n6925), .Y(n7814) );
  NAND2XL U3031 ( .A(n2877), .B(n6905), .Y(n6927) );
  OA22XL U3032 ( .A0(n6908), .A1(n6907), .B0(n6906), .B1(n7001), .Y(n6926) );
  NAND2XL U3033 ( .A(n5959), .B(n6620), .Y(n5999) );
  NAND4X2 U3034 ( .A(n6704), .B(n6703), .C(n6702), .D(n6701), .Y(n8225) );
  NAND2XL U3035 ( .A(n6676), .B(n6905), .Y(n6703) );
  AOI2BB1XL U3036 ( .A0N(n6824), .A1N(n6755), .B0(n5622), .Y(n5623) );
  NAND2BXL U3037 ( .AN(n3576), .B(n8565), .Y(n7605) );
  INVX3 U3038 ( .A(n8263), .Y(n6120) );
  NAND2BXL U3039 ( .AN(n3576), .B(n8568), .Y(n7532) );
  NAND2BXL U3040 ( .AN(n3576), .B(n8566), .Y(n7629) );
  NAND2BXL U3041 ( .AN(n3576), .B(n8563), .Y(n7706) );
  NAND2BXL U3042 ( .AN(n3576), .B(n8564), .Y(n7683) );
  INVXL U3043 ( .A(n6323), .Y(n6325) );
  BUFX2 U3044 ( .A(n3263), .Y(n3261) );
  BUFX2 U3045 ( .A(n3396), .Y(n3394) );
  BUFX2 U3046 ( .A(n2800), .Y(n3529) );
  CLKBUFX2 U3047 ( .A(n3263), .Y(n3260) );
  CLKBUFX2 U3048 ( .A(n3396), .Y(n3393) );
  CLKBUFX2 U3049 ( .A(n3308), .Y(n3307) );
  CLKBUFX2 U3050 ( .A(n2800), .Y(n3528) );
  INVXL U3051 ( .A(n5975), .Y(n4604) );
  INVX1 U3052 ( .A(n6838), .Y(n6840) );
  MX2XL U3053 ( .A(n3072), .B(n2865), .S0(n5828), .Y(n5829) );
  MX2XL U3054 ( .A(n3072), .B(n2865), .S0(n5905), .Y(n5906) );
  MX2XL U3055 ( .A(n3072), .B(n2865), .S0(n5549), .Y(n5550) );
  MX2XL U3056 ( .A(n3072), .B(n2865), .S0(n5621), .Y(n5622) );
  MX2XL U3057 ( .A(n7005), .B(n3071), .S0(n4816), .Y(n4817) );
  MX2XL U3058 ( .A(n3071), .B(n7005), .S0(n6690), .Y(n6459) );
  MX2XL U3059 ( .A(n3071), .B(n7005), .S0(n6061), .Y(n5461) );
  OAI222X1 U3060 ( .A0(n5960), .A1(n3069), .B0(n3068), .B1(n5973), .C0(n5970), 
        .C1(n5898), .Y(n6268) );
  MXI2XL U3061 ( .A(n5396), .B(n5395), .S0(n4016), .Y(n2831) );
  AOI21XL U3062 ( .A0(n8497), .A1(n15), .B0(n8494), .Y(n2821) );
  AOI21XL U3063 ( .A0(n6192), .A1(n8467), .B0(n8516), .Y(n2820) );
  NAND2BXL U3064 ( .AN(n19), .B(n6257), .Y(n4831) );
  INVX3 U3065 ( .A(n6772), .Y(n6549) );
  INVXL U3066 ( .A(n6267), .Y(n5899) );
  INVX1 U3067 ( .A(n4638), .Y(n5473) );
  INVX1 U3068 ( .A(n5984), .Y(n4637) );
  MX2XL U3069 ( .A(n5266), .B(n6772), .S0(n4016), .Y(n4966) );
  XOR3XL U3070 ( .A(n8368), .B(n2814), .C(n8367), .Y(n8371) );
  NAND2XL U3071 ( .A(n5484), .B(n2832), .Y(n4820) );
  INVX3 U3072 ( .A(n5734), .Y(n5682) );
  INVX1 U3073 ( .A(n6203), .Y(n5116) );
  AO21XL U3074 ( .A0(n5824), .A1(n6337), .B0(n2874), .Y(n6403) );
  INVXL U3075 ( .A(n6123), .Y(n6126) );
  INVXL U3076 ( .A(n5747), .Y(n5183) );
  MX2XL U3077 ( .A(n6475), .B(n5813), .S0(n4016), .Y(n6206) );
  INVXL U3078 ( .A(n8539), .Y(n8542) );
  CLKBUFX2 U3079 ( .A(n3264), .Y(n3258) );
  CLKBUFX2 U3080 ( .A(n3394), .Y(n3392) );
  CLKBUFX2 U3081 ( .A(n3308), .Y(n3305) );
  CLKBUFX2 U3082 ( .A(n3441), .Y(n3436) );
  INVX1 U3083 ( .A(n8525), .Y(n8529) );
  INVX1 U3084 ( .A(n8530), .Y(n8534) );
  AND2XL U3085 ( .A(n8349), .B(n8348), .Y(n2814) );
  AND2XL U3086 ( .A(n7893), .B(n7952), .Y(n2827) );
  INVX1 U3087 ( .A(n4666), .Y(n4695) );
  MX2XL U3088 ( .A(n6673), .B(n6331), .S0(n55), .Y(n6053) );
  AND2XL U3089 ( .A(n5484), .B(n4017), .Y(n2824) );
  CLKBUFX2 U3090 ( .A(\D_cache/n455 ), .Y(n3996) );
  CLKBUFX2 U3091 ( .A(n8718), .Y(n3637) );
  CLKBUFX2 U3092 ( .A(n8744), .Y(n3686) );
  NAND3BXL U3093 ( .AN(n8684), .B(n8683), .C(n8682), .Y(n8687) );
  NAND2XL U3094 ( .A(n8392), .B(n4538), .Y(n8683) );
  XOR3XL U3095 ( .A(n8383), .B(n8382), .C(n8381), .Y(n8386) );
  NAND2XL U3096 ( .A(n8427), .B(n4539), .Y(n8553) );
  AO21XL U3097 ( .A0(n6337), .A1(n6336), .B0(n2874), .Y(n6989) );
  XOR3XL U3098 ( .A(n2840), .B(n8336), .C(n8335), .Y(n8337) );
  INVXL U3099 ( .A(n8243), .Y(n8370) );
  INVXL U3100 ( .A(n8163), .Y(n8416) );
  INVXL U3101 ( .A(n8234), .Y(n8400) );
  INVXL U3102 ( .A(n8160), .Y(n8356) );
  INVXL U3103 ( .A(n8029), .Y(n8036) );
  INVXL U3104 ( .A(n8177), .Y(n8264) );
  INVXL U3105 ( .A(n8151), .Y(n8158) );
  INVXL U3106 ( .A(n7938), .Y(n8252) );
  INVXL U3107 ( .A(n7875), .Y(n8245) );
  INVXL U3108 ( .A(n7829), .Y(n8010) );
  INVXL U3109 ( .A(n7887), .Y(n8013) );
  INVXL U3110 ( .A(n8236), .Y(n8239) );
  INVXL U3111 ( .A(n7661), .Y(n8329) );
  INVXL U3112 ( .A(n22), .Y(n8312) );
  INVXL U3113 ( .A(n8199), .Y(n8458) );
  INVXL U3114 ( .A(n8295), .Y(n8299) );
  INVXL U3115 ( .A(n6619), .Y(n5182) );
  INVXL U3116 ( .A(n6621), .Y(n6622) );
  NAND2BXL U3117 ( .AN(n3576), .B(n8574), .Y(n7508) );
  NAND2BXL U3118 ( .AN(n3576), .B(n8579), .Y(n7658) );
  NAND2BXL U3119 ( .AN(n3576), .B(n8575), .Y(n7484) );
  NAND2BXL U3120 ( .AN(n3576), .B(n8571), .Y(n7088) );
  INVXL U3121 ( .A(n6837), .Y(n6827) );
  INVXL U3122 ( .A(n6907), .Y(n5974) );
  CLKBUFX2 U3123 ( .A(n3264), .Y(n3255) );
  CLKBUFX2 U3124 ( .A(n3442), .Y(n3433) );
  CLKBUFX2 U3125 ( .A(n3397), .Y(n3389) );
  CLKBUFX2 U3126 ( .A(n3487), .Y(n3480) );
  CLKBUFX2 U3127 ( .A(n3531), .Y(n3524) );
  CLKBUFX2 U3128 ( .A(n3463), .Y(n3483) );
  CLKBUFX2 U3129 ( .A(n3530), .Y(n3527) );
  CLKBUFX2 U3130 ( .A(n3256), .Y(n3259) );
  INVXL U3131 ( .A(n5990), .Y(n5957) );
  INVX1 U3132 ( .A(n8074), .Y(n8076) );
  INVX1 U3133 ( .A(n8179), .Y(n8181) );
  INVX1 U3134 ( .A(n8456), .Y(n8138) );
  INVX1 U3135 ( .A(n8201), .Y(n8202) );
  MX2XL U3136 ( .A(n2098), .B(n8229), .S0(n3625), .Y(\i_MIPS/n465 ) );
  MX2XL U3137 ( .A(n2221), .B(n8242), .S0(n3624), .Y(\i_MIPS/n464 ) );
  MX2XL U3138 ( .A(n10321), .B(n8159), .S0(n3624), .Y(\i_MIPS/n463 ) );
  CLKBUFX2 U3139 ( .A(n3975), .Y(n3971) );
  NAND3X1 U3140 ( .A(n2057), .B(n2150), .C(n2209), .Y(\D_cache/n211 ) );
  NAND3X1 U3141 ( .A(n2207), .B(n2058), .C(n3065), .Y(\D_cache/n207 ) );
  NAND3X1 U3142 ( .A(n2060), .B(n2164), .C(n3063), .Y(\D_cache/n209 ) );
  NAND3X1 U3143 ( .A(n2165), .B(n2148), .C(n2128), .Y(\D_cache/n212 ) );
  NAND3X1 U3144 ( .A(n2165), .B(n2148), .C(n2059), .Y(\D_cache/n213 ) );
  BUFX12 U3145 ( .A(n6842), .Y(n3070) );
  NAND3BX2 U3146 ( .AN(n5405), .B(n5404), .C(n5403), .Y(n8242) );
  AO21X4 U3147 ( .A0(n8359), .A1(n8358), .B0(n2855), .Y(n7868) );
  AOI221X2 U3148 ( .A0(n7869), .A1(n7868), .B0(n7867), .B1(n7866), .C0(n2854), 
        .Y(n7870) );
  NAND2X4 U3149 ( .A(n2155), .B(n4388), .Y(n2767) );
  NAND2XL U3150 ( .A(n8518), .B(n8520), .Y(n6768) );
  NAND2XL U3151 ( .A(n8485), .B(n8478), .Y(n6329) );
  AO22XL U3152 ( .A0(n6325), .A1(n3104), .B0(n3109), .B1(n6324), .Y(n6327) );
  NAND2XL U3153 ( .A(n5621), .B(n5602), .Y(n5607) );
  NAND4X2 U3154 ( .A(n7534), .B(n7533), .C(n7532), .D(n7531), .Y(n7985) );
  NAND4X2 U3155 ( .A(n7631), .B(n7630), .C(n7629), .D(n7628), .Y(n7955) );
  OAI222X2 U3156 ( .A0(n6045), .A1(n3164), .B0(n6023), .B1(n2761), .C0(n4), 
        .C1(n3163), .Y(n7808) );
  NAND2X4 U3157 ( .A(n4678), .B(\i_MIPS/n367 ), .Y(n8504) );
  NAND2X2 U3158 ( .A(n4644), .B(\i_MIPS/n352 ), .Y(n8535) );
  XNOR2X2 U3159 ( .A(n1619), .B(\D_cache/N40 ), .Y(\D_cache/n530 ) );
  AOI2BB2XL U3160 ( .B0(\D_cache/N148 ), .B1(n2153), .A0N(n23), .A1N(n8898), 
        .Y(\D_cache/n173 ) );
  OA22X4 U3161 ( .A0(n3371), .A1(n976), .B0(n3328), .B1(n88), .Y(n4446) );
  OA22X4 U3162 ( .A0(n3284), .A1(n978), .B0(n3236), .B1(n90), .Y(n4447) );
  NAND2XL U3163 ( .A(n6533), .B(n5124), .Y(n5125) );
  INVXL U3164 ( .A(n8060), .Y(n8044) );
  NAND3X2 U3165 ( .A(n6535), .B(n6600), .C(n6534), .Y(n4593) );
  AO21X4 U3166 ( .A0(n7983), .A1(n7982), .B0(n2856), .Y(n8023) );
  NAND2X2 U3167 ( .A(n4671), .B(\i_MIPS/n366 ), .Y(n8502) );
  NAND2X2 U3168 ( .A(n4661), .B(\i_MIPS/n360 ), .Y(n8471) );
  NAND2XL U3169 ( .A(n6128), .B(n6127), .Y(n6190) );
  NAND2XL U3170 ( .A(n6258), .B(n6257), .Y(n6392) );
  AND3X2 U3171 ( .A(n2768), .B(n2769), .C(n2770), .Y(n3042) );
  XNOR2X1 U3172 ( .A(\D_cache/N55 ), .B(DCACHE_addr[6]), .Y(n2768) );
  XNOR2X1 U3173 ( .A(\D_cache/N54 ), .B(DCACHE_addr[7]), .Y(n2770) );
  OA22XL U3174 ( .A0(n6612), .A1(n5330), .B0(n6138), .B1(n6550), .Y(n5060) );
  MX2XL U3175 ( .A(n7005), .B(n3071), .S0(n5037), .Y(n5062) );
  NAND4X2 U3176 ( .A(n6213), .B(n6212), .C(n6211), .D(n6210), .Y(n8244) );
  OA22XL U3177 ( .A0(n6202), .A1(n6201), .B0(n2796), .B1(n6200), .Y(n6212) );
  OA22XL U3178 ( .A0(n7009), .A1(n6826), .B0(n6825), .B1(n6824), .Y(n6857) );
  MX2XL U3179 ( .A(n7005), .B(n3071), .S0(n6827), .Y(n6856) );
  NAND2XL U3180 ( .A(n5734), .B(n5681), .Y(n5678) );
  NAND2XL U3181 ( .A(n8541), .B(n8540), .Y(n5677) );
  MX2XL U3182 ( .A(n7005), .B(n3071), .S0(n5111), .Y(n5133) );
  NAND2XL U3183 ( .A(n3579), .B(n8420), .Y(n8084) );
  CLKXOR2X2 U3184 ( .A(n1085), .B(\D_cache/N48 ), .Y(n3045) );
  AOI2BB2XL U3185 ( .B0(\D_cache/N147 ), .B1(n2153), .A0N(n23), .A1N(n8897), 
        .Y(\D_cache/n172 ) );
  NAND3X2 U3186 ( .A(n6533), .B(n6603), .C(n6532), .Y(n4683) );
  NAND2X2 U3187 ( .A(n6537), .B(n5384), .Y(n4897) );
  OA22XL U3188 ( .A0(n3372), .A1(n1077), .B0(n3329), .B1(n165), .Y(n4458) );
  OA22X4 U3189 ( .A0(n3542), .A1(n979), .B0(n3531), .B1(n91), .Y(n4424) );
  NAND4X4 U3190 ( .A(n4427), .B(n4426), .C(n4425), .D(n4424), .Y(n8691) );
  OA22X4 U3191 ( .A0(n3397), .A1(n980), .B0(n3324), .B1(n92), .Y(n4426) );
  AOI222XL U3192 ( .A0(n6774), .A1(n6773), .B0(n2813), .B1(n6772), .C0(n6771), 
        .C1(n6993), .Y(n6775) );
  NAND2XL U3193 ( .A(n7007), .B(n6620), .Y(n6074) );
  MX2XL U3194 ( .A(n7005), .B(n3071), .S0(n6046), .Y(n6075) );
  AOI2BB1XL U3195 ( .A0N(n2758), .A1N(n6260), .B0(n6259), .Y(n6261) );
  NAND2BX4 U3196 ( .AN(n5982), .B(n5981), .Y(n6839) );
  AOI2BB1X2 U3197 ( .A0N(n5980), .A1N(n5979), .B0(n5978), .Y(n5982) );
  INVX3 U3198 ( .A(n6466), .Y(n5980) );
  MX2X2 U3199 ( .A(n5742), .B(n5741), .S0(n5740), .Y(n5760) );
  AOI211X2 U3200 ( .A0(n6905), .A1(n6053), .B0(n5751), .C0(n5750), .Y(n5759)
         );
  NOR4X4 U3201 ( .A(\D_cache/n550 ), .B(\D_cache/n551 ), .C(\D_cache/n552 ), 
        .D(\D_cache/n553 ), .Y(n2771) );
  AND4X4 U3202 ( .A(n7793), .B(n7792), .C(n7791), .D(n7790), .Y(n2862) );
  NAND2XL U3203 ( .A(n7832), .B(\i_MIPS/n233 ), .Y(n7793) );
  OA22X4 U3204 ( .A0(n3370), .A1(n983), .B0(n3327), .B1(n95), .Y(n4442) );
  OA22X4 U3205 ( .A0(n3545), .A1(n984), .B0(n3504), .B1(n96), .Y(n4440) );
  OA22X4 U3206 ( .A0(n3283), .A1(n985), .B0(n3235), .B1(n97), .Y(n4443) );
  OA22X4 U3207 ( .A0(n3368), .A1(n989), .B0(n3325), .B1(n101), .Y(n4434) );
  OA22X4 U3208 ( .A0(n3543), .A1(n990), .B0(n3502), .B1(n102), .Y(n4432) );
  OA22X4 U3209 ( .A0(n3281), .A1(n991), .B0(n3233), .B1(n103), .Y(n4435) );
  AOI2BB2XL U3210 ( .B0(\D_cache/N142 ), .B1(n2153), .A0N(n24), .A1N(n8892), 
        .Y(\D_cache/n198 ) );
  OAI211X2 U3211 ( .A0(n6904), .A1(n4649), .B0(n5681), .C0(n6914), .Y(n4650)
         );
  OA22X4 U3212 ( .A0(n7556), .A1(n3576), .B0(n7555), .B1(n3001), .Y(n7557) );
  OA22XL U3213 ( .A0(\i_MIPS/n368 ), .A1(n3082), .B0(\i_MIPS/n367 ), .B1(n3078), .Y(n4819) );
  OA22XL U3214 ( .A0(\i_MIPS/n358 ), .A1(n14), .B0(\i_MIPS/n357 ), .B1(n3077), 
        .Y(n5745) );
  AOI2BB1XL U3215 ( .A0N(\i_MIPS/n368 ), .A1N(n3078), .B0(n2900), .Y(n4713) );
  OA21XL U3216 ( .A0(\i_MIPS/n365 ), .A1(n3092), .B0(n5463), .Y(n5464) );
  OA21XL U3217 ( .A0(\i_MIPS/n352 ), .A1(n3082), .B0(n5744), .Y(n4915) );
  AOI2BB1XL U3218 ( .A0N(\i_MIPS/n368 ), .A1N(n3092), .B0(n2898), .Y(n4892) );
  OA22XL U3219 ( .A0(\i_MIPS/n367 ), .A1(n14), .B0(\i_MIPS/n366 ), .B1(n3078), 
        .Y(n5380) );
  OA21XL U3220 ( .A0(\i_MIPS/n362 ), .A1(n3086), .B0(n5118), .Y(n4714) );
  AOI2BB1XL U3221 ( .A0N(\i_MIPS/n356 ), .A1N(n3078), .B0(n2987), .Y(n4716) );
  AOI2BB1XL U3222 ( .A0N(\i_MIPS/n365 ), .A1N(n3087), .B0(n2984), .Y(n4840) );
  OA21XL U3223 ( .A0(\i_MIPS/n359 ), .A1(n3082), .B0(n5457), .Y(n5458) );
  AO21XL U3224 ( .A0(n6824), .A1(n4820), .B0(n6847), .Y(n4722) );
  OAI22X1 U3225 ( .A0(n8908), .A1(n8907), .B0(n2842), .B1(n8908), .Y(n8911) );
  OA22XL U3226 ( .A0(n3554), .A1(n547), .B0(n3512), .B1(n1466), .Y(n7339) );
  OA22XL U3227 ( .A0(n3377), .A1(n548), .B0(n3335), .B1(n1467), .Y(n7341) );
  OA22XL U3228 ( .A0(n3290), .A1(n549), .B0(n3243), .B1(n1468), .Y(n7342) );
  OA22XL U3229 ( .A0(n3553), .A1(n550), .B0(n3511), .B1(n1469), .Y(n7331) );
  OA22XL U3230 ( .A0(n3376), .A1(n551), .B0(n3334), .B1(n1470), .Y(n7333) );
  OA22XL U3231 ( .A0(n3289), .A1(n552), .B0(n3242), .B1(n1471), .Y(n7334) );
  OA22XL U3232 ( .A0(n3290), .A1(n553), .B0(n3243), .B1(n1472), .Y(n7362) );
  OA22XL U3233 ( .A0(n3468), .A1(n554), .B0(n3421), .B1(n1473), .Y(n7360) );
  OA22XL U3234 ( .A0(n3377), .A1(n555), .B0(n3335), .B1(n1474), .Y(n7361) );
  OA22XL U3235 ( .A0(n3290), .A1(n556), .B0(n3243), .B1(n1475), .Y(n7358) );
  OA22XL U3236 ( .A0(n3468), .A1(n557), .B0(n3421), .B1(n1476), .Y(n7356) );
  OA22XL U3237 ( .A0(n3377), .A1(n558), .B0(n3335), .B1(n1477), .Y(n7357) );
  OA22XL U3238 ( .A0(n3376), .A1(n559), .B0(n3334), .B1(n1478), .Y(n7337) );
  OA22XL U3239 ( .A0(n3289), .A1(n560), .B0(n3242), .B1(n1479), .Y(n7338) );
  OA22XL U3240 ( .A0(n3290), .A1(n561), .B0(n3243), .B1(n1480), .Y(n7354) );
  OA22XL U3241 ( .A0(n3468), .A1(n562), .B0(n3421), .B1(n1481), .Y(n7352) );
  OA22XL U3242 ( .A0(n3377), .A1(n563), .B0(n3335), .B1(n1482), .Y(n7353) );
  NAND4X2 U3243 ( .A(n7212), .B(n7211), .C(n7210), .D(n7209), .Y(n7837) );
  NAND2BXL U3244 ( .AN(n3576), .B(n8582), .Y(n7234) );
  AOI2BB1XL U3245 ( .A0N(n8486), .A1N(n8485), .B0(n8484), .Y(n8487) );
  INVXL U3246 ( .A(n8471), .Y(n8472) );
  NAND2XL U3247 ( .A(n2145), .B(\i_MIPS/n360 ), .Y(n5270) );
  NAND2XL U3248 ( .A(n6535), .B(n6534), .Y(n8497) );
  AOI21XL U3249 ( .A0(n5388), .A1(n8504), .B0(n5387), .Y(n2851) );
  AOI21XL U3250 ( .A0(n4970), .A1(n8506), .B0(n4969), .Y(n2852) );
  NAND2XL U3251 ( .A(n6537), .B(n5321), .Y(n5386) );
  NAND2XL U3252 ( .A(n3613), .B(n7307), .Y(n7636) );
  MXI2XL U3253 ( .A(n5481), .B(n6477), .S0(n4016), .Y(n5482) );
  NAND3XL U3254 ( .A(n8465), .B(n2833), .C(n8549), .Y(n8806) );
  NAND2BXL U3255 ( .AN(n8483), .B(n8480), .Y(n8513) );
  AOI2BB1XL U3256 ( .A0N(n4902), .A1N(n4901), .B0(n4900), .Y(n4903) );
  INVXL U3257 ( .A(n5322), .Y(n4902) );
  INVXL U3258 ( .A(n7), .Y(n8515) );
  NAND2XL U3259 ( .A(n5322), .B(n8492), .Y(n5388) );
  NAND2XL U3260 ( .A(n3094), .B(\i_MIPS/n357 ), .Y(n5456) );
  NAND2XL U3261 ( .A(n3089), .B(\i_MIPS/n357 ), .Y(n5040) );
  NAND2XL U3262 ( .A(n6129), .B(n8510), .Y(n6192) );
  NAND2XL U3263 ( .A(n4633), .B(\i_MIPS/n349 ), .Y(n8543) );
  INVX1 U3264 ( .A(n4631), .Y(n4640) );
  OAI2BB1XL U3265 ( .A0N(n4973), .A1N(n4972), .B0(n4971), .Y(n4974) );
  OAI2BB1XL U3266 ( .A0N(n5386), .A1N(n5385), .B0(n5384), .Y(n5389) );
  INVX1 U3267 ( .A(n6686), .Y(n7011) );
  OAI2BB1XL U3268 ( .A0N(n8542), .A1N(n8541), .B0(n8540), .Y(n8914) );
  INVX1 U3269 ( .A(n8531), .Y(n8532) );
  INVX3 U3270 ( .A(n8025), .Y(n8026) );
  OAI211XL U3271 ( .A0(n8505), .A1(n8504), .B0(n8503), .C0(n8502), .Y(n8508)
         );
  NAND2XL U3272 ( .A(n2816), .B(n5048), .Y(n5050) );
  NAND3BXL U3273 ( .AN(n2803), .B(n7636), .C(n7635), .Y(\i_MIPS/n470 ) );
  OA22XL U3274 ( .A0(\i_MIPS/Control_ID/n15 ), .A1(n3073), .B0(n3627), .B1(
        n4020), .Y(n7635) );
  INVXL U3275 ( .A(n6757), .Y(n6758) );
  AOI2BB1XL U3276 ( .A0N(\i_MIPS/n355 ), .A1N(n3078), .B0(n2905), .Y(n5052) );
  AND2X1 U3277 ( .A(n3069), .B(\i_MIPS/n340 ), .Y(n2874) );
  INVXL U3278 ( .A(n5321), .Y(n4898) );
  MX2XL U3279 ( .A(n5620), .B(n5619), .S0(n55), .Y(n6755) );
  INVXL U3280 ( .A(n6829), .Y(n5619) );
  MX2XL U3281 ( .A(\i_MIPS/n340 ), .B(\i_MIPS/n341 ), .S0(n3080), .Y(n6336) );
  OAI2BB1XL U3282 ( .A0N(n8469), .A1N(n7), .B0(n8468), .Y(n8475) );
  OAI221X1 U3283 ( .A0(n6332), .A1(n5815), .B0(n3068), .B1(n6475), .C0(n5814), 
        .Y(n6401) );
  OA22X2 U3284 ( .A0(n6334), .A1(n5813), .B0(n6463), .B1(n3069), .Y(n5814) );
  MXI2XL U3285 ( .A(n5962), .B(n5961), .S0(n4016), .Y(n2877) );
  OA22XL U3286 ( .A0(\i_MIPS/n362 ), .A1(n14), .B0(\i_MIPS/n361 ), .B1(n3077), 
        .Y(n5201) );
  MX2XL U3287 ( .A(n6675), .B(n6674), .S0(n55), .Y(n7000) );
  MX2XL U3288 ( .A(n5616), .B(n2985), .S0(n4016), .Y(n6759) );
  MX2XL U3289 ( .A(n5823), .B(n5822), .S0(n55), .Y(n6460) );
  AND2XL U3290 ( .A(n2863), .B(\i_MIPS/n356 ), .Y(n2844) );
  AND2XL U3291 ( .A(n3083), .B(\i_MIPS/n355 ), .Y(n2878) );
  MX2XL U3292 ( .A(n5269), .B(n5268), .S0(n4016), .Y(n6551) );
  MX2XL U3293 ( .A(n5329), .B(n5328), .S0(n4016), .Y(n6269) );
  INVXL U3294 ( .A(n6135), .Y(n5328) );
  MX2XL U3295 ( .A(n5822), .B(n5459), .S0(n55), .Y(n5684) );
  INVXL U3296 ( .A(n6463), .Y(n5459) );
  INVXL U3297 ( .A(n5746), .Y(n4916) );
  AND2XL U3298 ( .A(n3093), .B(\i_MIPS/n358 ), .Y(n2879) );
  OAI2BB1XL U3299 ( .A0N(n8550), .A1N(n8549), .B0(n8548), .Y(n8916) );
  NAND4XL U3300 ( .A(n7015), .B(n7014), .C(n7013), .D(n7012), .Y(n7016) );
  MX2XL U3301 ( .A(n7005), .B(n3071), .S0(n7003), .Y(n7015) );
  NAND2XL U3302 ( .A(n7007), .B(n7006), .Y(n7013) );
  MX2XL U3303 ( .A(n5748), .B(n6686), .S0(n4016), .Y(n5205) );
  MX2XL U3304 ( .A(n5813), .B(n5815), .S0(n4016), .Y(n5382) );
  INVXL U3305 ( .A(n6847), .Y(n4975) );
  NAND2X1 U3306 ( .A(n2983), .B(n2975), .Y(n2776) );
  CLKINVX3 U3307 ( .A(\i_MIPS/n320 ), .Y(n4014) );
  OA22XL U3308 ( .A0(n3559), .A1(n564), .B0(n3517), .B1(n1483), .Y(n7584) );
  OA22XL U3309 ( .A0(n3382), .A1(n565), .B0(n3340), .B1(n1484), .Y(n7586) );
  OA22XL U3310 ( .A0(n3295), .A1(n566), .B0(n3248), .B1(n1485), .Y(n7587) );
  OA22XL U3311 ( .A0(n3290), .A1(n567), .B0(n3243), .B1(n1486), .Y(n7350) );
  OA22XL U3312 ( .A0(n3468), .A1(n568), .B0(n3421), .B1(n1487), .Y(n7348) );
  OA22XL U3313 ( .A0(n3377), .A1(n569), .B0(n3335), .B1(n1488), .Y(n7349) );
  OA22XL U3314 ( .A0(n3555), .A1(n570), .B0(n3513), .B1(n1489), .Y(n7392) );
  OA22XL U3315 ( .A0(n3378), .A1(n571), .B0(n3336), .B1(n1490), .Y(n7394) );
  OA22XL U3316 ( .A0(n3291), .A1(n572), .B0(n3244), .B1(n1491), .Y(n7395) );
  NAND4BX1 U3317 ( .AN(n2778), .B(n7771), .C(n7770), .D(n7769), .Y(n8560) );
  OAI22XL U3318 ( .A0(n3300), .A1(n460), .B0(n3253), .B1(n1369), .Y(n2778) );
  OA22XL U3319 ( .A0(n3378), .A1(n573), .B0(n3336), .B1(n1492), .Y(n7389) );
  OA22XL U3320 ( .A0(n3555), .A1(n574), .B0(n3513), .B1(n1493), .Y(n7387) );
  OA22XL U3321 ( .A0(n3291), .A1(n575), .B0(n3244), .B1(n1494), .Y(n7390) );
  OA22XL U3322 ( .A0(n3564), .A1(n576), .B0(n3522), .B1(n1495), .Y(n7759) );
  OA22XL U3323 ( .A0(n3387), .A1(n577), .B0(n3345), .B1(n1496), .Y(n7761) );
  OA22XL U3324 ( .A0(n3300), .A1(n578), .B0(n3253), .B1(n1497), .Y(n7762) );
  OA22XL U3325 ( .A0(n3559), .A1(n579), .B0(n3517), .B1(n1498), .Y(n7575) );
  OA22XL U3326 ( .A0(n3382), .A1(n580), .B0(n3340), .B1(n1499), .Y(n7577) );
  OA22XL U3327 ( .A0(n3295), .A1(n581), .B0(n3248), .B1(n1500), .Y(n7578) );
  OA22XL U3328 ( .A0(n3558), .A1(n582), .B0(n3516), .B1(n1501), .Y(n7526) );
  OA22XL U3329 ( .A0(n3381), .A1(n583), .B0(n3339), .B1(n1502), .Y(n7528) );
  OA22XL U3330 ( .A0(n3294), .A1(n584), .B0(n3247), .B1(n1503), .Y(n7529) );
  OA22XL U3331 ( .A0(n3555), .A1(n585), .B0(n3513), .B1(n1504), .Y(n7397) );
  OA22XL U3332 ( .A0(n3378), .A1(n586), .B0(n3336), .B1(n1505), .Y(n7399) );
  OA22XL U3333 ( .A0(n3291), .A1(n587), .B0(n3244), .B1(n1506), .Y(n7400) );
  OA22XL U3334 ( .A0(n3558), .A1(n588), .B0(n3516), .B1(n1507), .Y(n7521) );
  OA22XL U3335 ( .A0(n3381), .A1(n589), .B0(n3339), .B1(n1508), .Y(n7523) );
  OA22XL U3336 ( .A0(n3294), .A1(n590), .B0(n3247), .B1(n1509), .Y(n7524) );
  OA22XL U3337 ( .A0(n3559), .A1(n591), .B0(n3517), .B1(n1510), .Y(n7565) );
  OA22XL U3338 ( .A0(n3382), .A1(n592), .B0(n3340), .B1(n1511), .Y(n7567) );
  OA22XL U3339 ( .A0(n3295), .A1(n593), .B0(n3248), .B1(n1512), .Y(n7568) );
  OA22XL U3340 ( .A0(n3558), .A1(n594), .B0(n3516), .B1(n1513), .Y(n7516) );
  OA22XL U3341 ( .A0(n3381), .A1(n595), .B0(n3339), .B1(n1514), .Y(n7518) );
  OA22XL U3342 ( .A0(n3294), .A1(n596), .B0(n3247), .B1(n1515), .Y(n7519) );
  OA22XL U3343 ( .A0(n3559), .A1(n597), .B0(n3517), .B1(n1516), .Y(n7560) );
  OA22XL U3344 ( .A0(n3382), .A1(n598), .B0(n3340), .B1(n1517), .Y(n7562) );
  OA22XL U3345 ( .A0(n3295), .A1(n599), .B0(n3248), .B1(n1518), .Y(n7563) );
  OA22XL U3346 ( .A0(n3559), .A1(n600), .B0(n3517), .B1(n1519), .Y(n7570) );
  OA22XL U3347 ( .A0(n3382), .A1(n601), .B0(n3340), .B1(n1520), .Y(n7572) );
  OA22XL U3348 ( .A0(n3295), .A1(n602), .B0(n3248), .B1(n1521), .Y(n7573) );
  NAND4BX1 U3349 ( .AN(n2779), .B(n7621), .C(n7620), .D(n7619), .Y(n8566) );
  OAI22XL U3350 ( .A0(n3296), .A1(n461), .B0(n3249), .B1(n1370), .Y(n2779) );
  OA22XL U3351 ( .A0(n3383), .A1(n603), .B0(n3341), .B1(n1522), .Y(n7611) );
  OA22XL U3352 ( .A0(n3296), .A1(n604), .B0(n3249), .B1(n1523), .Y(n7612) );
  OA22XL U3353 ( .A0(n3560), .A1(n605), .B0(n3518), .B1(n1524), .Y(n7609) );
  NAND4BX1 U3354 ( .AN(n2780), .B(n7726), .C(n7725), .D(n7724), .Y(n8594) );
  OAI22XL U3355 ( .A0(n3299), .A1(n462), .B0(n3252), .B1(n1371), .Y(n2780) );
  OA22XL U3356 ( .A0(n3386), .A1(n606), .B0(n3344), .B1(n1525), .Y(n7702) );
  OA22XL U3357 ( .A0(n3299), .A1(n607), .B0(n3252), .B1(n1526), .Y(n7703) );
  OA22XL U3358 ( .A0(n3563), .A1(n608), .B0(n3521), .B1(n1527), .Y(n7700) );
  OA22XL U3359 ( .A0(n3386), .A1(n609), .B0(n3344), .B1(n1528), .Y(n7716) );
  OA22XL U3360 ( .A0(n3299), .A1(n610), .B0(n3252), .B1(n1529), .Y(n7717) );
  OA22XL U3361 ( .A0(n3563), .A1(n611), .B0(n3521), .B1(n1530), .Y(n7714) );
  NAND4BX1 U3362 ( .AN(n2781), .B(n7698), .C(n7697), .D(n7696), .Y(n8563) );
  OA22XL U3363 ( .A0(n3564), .A1(n612), .B0(n3522), .B1(n1531), .Y(n7740) );
  OA22XL U3364 ( .A0(n3387), .A1(n613), .B0(n3345), .B1(n1532), .Y(n7742) );
  OA22XL U3365 ( .A0(n3300), .A1(n614), .B0(n3253), .B1(n1533), .Y(n7743) );
  OA22XL U3366 ( .A0(n3386), .A1(n615), .B0(n3344), .B1(n1534), .Y(n7711) );
  OA22XL U3367 ( .A0(n3299), .A1(n616), .B0(n3252), .B1(n1535), .Y(n7712) );
  OA22XL U3368 ( .A0(n3563), .A1(n617), .B0(n3521), .B1(n1536), .Y(n7709) );
  OA22XL U3369 ( .A0(n3385), .A1(n618), .B0(n3343), .B1(n1537), .Y(n7688) );
  OA22XL U3370 ( .A0(n3298), .A1(n619), .B0(n3251), .B1(n1538), .Y(n7689) );
  OA22XL U3371 ( .A0(n3562), .A1(n620), .B0(n3520), .B1(n1539), .Y(n7686) );
  OA22XL U3372 ( .A0(n3562), .A1(n621), .B0(n3520), .B1(n1540), .Y(n7677) );
  OA22XL U3373 ( .A0(n3385), .A1(n622), .B0(n3343), .B1(n1541), .Y(n7679) );
  OA22XL U3374 ( .A0(n3298), .A1(n623), .B0(n3251), .B1(n1542), .Y(n7680) );
  OA22XL U3375 ( .A0(n3562), .A1(n624), .B0(n3520), .B1(n1543), .Y(n7672) );
  OA22XL U3376 ( .A0(n3385), .A1(n625), .B0(n3343), .B1(n1544), .Y(n7674) );
  OA22XL U3377 ( .A0(n3298), .A1(n626), .B0(n3251), .B1(n1545), .Y(n7675) );
  OA22XL U3378 ( .A0(n3562), .A1(n627), .B0(n3520), .B1(n1546), .Y(n7667) );
  OA22XL U3379 ( .A0(n3385), .A1(n628), .B0(n3343), .B1(n1547), .Y(n7669) );
  OA22XL U3380 ( .A0(n3298), .A1(n629), .B0(n3251), .B1(n1548), .Y(n7670) );
  OA22XL U3381 ( .A0(n3561), .A1(n630), .B0(n3519), .B1(n1549), .Y(n7662) );
  OA22XL U3382 ( .A0(n3384), .A1(n631), .B0(n3342), .B1(n1550), .Y(n7664) );
  OA22XL U3383 ( .A0(n3297), .A1(n632), .B0(n3250), .B1(n1551), .Y(n7665) );
  OA22XL U3384 ( .A0(n3296), .A1(n633), .B0(n3249), .B1(n1552), .Y(n7602) );
  OA22XL U3385 ( .A0(n3560), .A1(n634), .B0(n3518), .B1(n1553), .Y(n7589) );
  OA22XL U3386 ( .A0(n3383), .A1(n635), .B0(n3341), .B1(n1554), .Y(n7591) );
  OA22XL U3387 ( .A0(n3296), .A1(n636), .B0(n3249), .B1(n1555), .Y(n7592) );
  OA22XL U3388 ( .A0(n3289), .A1(n637), .B0(n3242), .B1(n1556), .Y(n7300) );
  OA22XL U3389 ( .A0(n3467), .A1(n638), .B0(n3420), .B1(n1557), .Y(n7298) );
  OA22XL U3390 ( .A0(n3376), .A1(n639), .B0(n3334), .B1(n1558), .Y(n7299) );
  CLKBUFX2 U3391 ( .A(n8727), .Y(n3652) );
  CLKBUFX2 U3392 ( .A(n8727), .Y(n3653) );
  NAND2XL U3393 ( .A(n4706), .B(\i_MIPS/n341 ), .Y(n7002) );
  NAND2XL U3394 ( .A(n4624), .B(n5900), .Y(n5905) );
  NAND2XL U3395 ( .A(n4623), .B(\i_MIPS/n342 ), .Y(n5828) );
  NAND2XL U3396 ( .A(n4625), .B(\i_MIPS/n344 ), .Y(n6762) );
  NAND3BXL U3397 ( .AN(n8427), .B(n3051), .C(n8426), .Y(n8452) );
  NAND2BXL U3398 ( .AN(\D_cache/n202 ), .B(\D_cache/n316 ), .Y(\D_cache/n384 )
         );
  NAND2BXL U3399 ( .AN(n3576), .B(n8573), .Y(n7137) );
  NAND2BXL U3400 ( .AN(n3576), .B(n8572), .Y(n7161) );
  NAND2BXL U3401 ( .AN(n3576), .B(n8570), .Y(n7113) );
  NAND2BXL U3402 ( .AN(n3576), .B(n8578), .Y(n7436) );
  NAND2BXL U3403 ( .AN(n3576), .B(n8576), .Y(n8135) );
  NAND2BXL U3404 ( .AN(n3576), .B(n8577), .Y(n7460) );
  INVX1 U3405 ( .A(n7930), .Y(n7933) );
  INVX1 U3406 ( .A(n7880), .Y(n7883) );
  INVX1 U3407 ( .A(n7848), .Y(n7851) );
  NAND2XL U3408 ( .A(n3094), .B(\i_MIPS/n353 ), .Y(n5465) );
  NAND2XL U3409 ( .A(n3094), .B(\i_MIPS/n354 ), .Y(n4914) );
  INVXL U3410 ( .A(\D_cache/N48 ), .Y(n8824) );
  NAND2XL U3411 ( .A(n4723), .B(\i_MIPS/n340 ), .Y(n4729) );
  INVXL U3412 ( .A(\D_cache/N34 ), .Y(n8811) );
  INVXL U3413 ( .A(\D_cache/N38 ), .Y(n8814) );
  INVXL U3414 ( .A(\D_cache/N41 ), .Y(n8817) );
  INVXL U3415 ( .A(\D_cache/N43 ), .Y(n8819) );
  INVXL U3416 ( .A(\D_cache/N46 ), .Y(n8822) );
  INVXL U3417 ( .A(\D_cache/N50 ), .Y(n8826) );
  INVXL U3418 ( .A(\D_cache/N52 ), .Y(n8828) );
  INVXL U3419 ( .A(\D_cache/N53 ), .Y(n8829) );
  INVXL U3420 ( .A(\D_cache/N55 ), .Y(n8831) );
  INVXL U3421 ( .A(\D_cache/N37 ), .Y(n8813) );
  INVXL U3422 ( .A(\D_cache/N39 ), .Y(n8815) );
  INVXL U3423 ( .A(\D_cache/N40 ), .Y(n8816) );
  INVXL U3424 ( .A(\D_cache/N42 ), .Y(n8818) );
  INVXL U3425 ( .A(\D_cache/N44 ), .Y(n8820) );
  INVXL U3426 ( .A(\D_cache/N56 ), .Y(n8832) );
  INVXL U3427 ( .A(\D_cache/N47 ), .Y(n8823) );
  INVXL U3428 ( .A(\D_cache/N49 ), .Y(n8825) );
  INVXL U3429 ( .A(\D_cache/N51 ), .Y(n8827) );
  INVXL U3430 ( .A(\D_cache/N54 ), .Y(n8830) );
  INVXL U3431 ( .A(\D_cache/N36 ), .Y(n8812) );
  INVXL U3432 ( .A(\D_cache/N45 ), .Y(n8821) );
  INVXL U3433 ( .A(n5815), .Y(n6202) );
  OR2XL U3434 ( .A(n8807), .B(\D_cache/n247 ), .Y(n8551) );
  NAND2X1 U3435 ( .A(n2983), .B(n2976), .Y(n2782) );
  NAND2X1 U3436 ( .A(n2972), .B(n2872), .Y(n2785) );
  INVXL U3437 ( .A(n5963), .Y(n5968) );
  NAND2XL U3438 ( .A(n8471), .B(n8473), .Y(n5264) );
  INVXL U3439 ( .A(n5602), .Y(n5618) );
  NAND2XL U3440 ( .A(n8498), .B(n8502), .Y(n5394) );
  NAND2XL U3441 ( .A(n8470), .B(n8466), .Y(n5200) );
  NAND2XL U3442 ( .A(n8504), .B(n8499), .Y(n5327) );
  NAND2XL U3443 ( .A(n8522), .B(n8524), .Y(n5477) );
  NAND2XL U3444 ( .A(n6061), .B(n5474), .Y(n5478) );
  NAND2XL U3445 ( .A(n8507), .B(n8506), .Y(n4908) );
  NAND2XL U3446 ( .A(n8468), .B(n7), .Y(n6198) );
  NAND2XL U3447 ( .A(n5256), .B(n5255), .Y(n5197) );
  NAND2XL U3448 ( .A(n8549), .B(n8548), .Y(n6471) );
  NAND2XL U3449 ( .A(n6258), .B(n5270), .Y(n5261) );
  AND2XL U3450 ( .A(n8531), .B(n8533), .Y(n2876) );
  AND2XL U3451 ( .A(n8526), .B(n8528), .Y(n2875) );
  NAND2XL U3452 ( .A(n6914), .B(n6913), .Y(n6915) );
  NAND2XL U3453 ( .A(n8492), .B(n8491), .Y(n6541) );
  NAND2XL U3454 ( .A(n6690), .B(n6474), .Y(n6472) );
  NAND2XL U3455 ( .A(n8510), .B(n8509), .Y(n4978) );
  NAND2XL U3456 ( .A(n6189), .B(n6188), .Y(n6131) );
  NAND2XL U3457 ( .A(n8467), .B(n6191), .Y(n6134) );
  NAND2XL U3458 ( .A(n6127), .B(n4987), .Y(n4979) );
  NAND2XL U3459 ( .A(n5385), .B(n5384), .Y(n5324) );
  NAND2XL U3460 ( .A(n6600), .B(n15), .Y(n6607) );
  NAND2XL U3461 ( .A(n6621), .B(n6603), .Y(n6604) );
  INVXL U3462 ( .A(n6603), .Y(n6608) );
  NAND2XL U3463 ( .A(n6194), .B(n6207), .Y(n6195) );
  NAND2XL U3464 ( .A(n5905), .B(n5890), .Y(n5896) );
  INVXL U3465 ( .A(n6468), .Y(n4841) );
  INVXL U3466 ( .A(n6194), .Y(n6199) );
  NAND2XL U3467 ( .A(n6537), .B(n6552), .Y(n6538) );
  NAND2XL U3468 ( .A(n8530), .B(n5891), .Y(n5895) );
  MX2XL U3469 ( .A(\i_MIPS/n366 ), .B(\i_MIPS/n365 ), .S0(n3075), .Y(n6528) );
  MX2XL U3470 ( .A(\i_MIPS/n342 ), .B(n5900), .S0(n3075), .Y(n5825) );
  AND2XL U3471 ( .A(n3088), .B(\i_MIPS/n354 ), .Y(n2880) );
  MX2XL U3472 ( .A(n5381), .B(\i_MIPS/n368 ), .S0(n3075), .Y(n6598) );
  MX2XL U3473 ( .A(\i_MIPS/n368 ), .B(\i_MIPS/n367 ), .S0(n3075), .Y(n6527) );
  MX2XL U3474 ( .A(n5900), .B(\i_MIPS/n344 ), .S0(n3075), .Y(n6994) );
  INVXL U3475 ( .A(n6537), .Y(n6542) );
  AND2XL U3476 ( .A(n6694), .B(n6693), .Y(n6695) );
  AND2XL U3477 ( .A(n6065), .B(n6064), .Y(n6066) );
  AND2XL U3478 ( .A(n5739), .B(n5738), .Y(n5740) );
  AND2XL U3479 ( .A(n5990), .B(n5989), .Y(n5991) );
  MX2XL U3480 ( .A(DCACHE_addr[18]), .B(n8223), .S0(n3625), .Y(\i_MIPS/n449 )
         );
  MX2XL U3481 ( .A(DCACHE_addr[12]), .B(n8251), .S0(n3626), .Y(\i_MIPS/n455 )
         );
  MX2XL U3482 ( .A(DCACHE_addr[27]), .B(n8284), .S0(n3623), .Y(\i_MIPS/n440 )
         );
  MX2XL U3483 ( .A(DCACHE_addr[14]), .B(n7814), .S0(n3624), .Y(\i_MIPS/n453 )
         );
  MX2XL U3484 ( .A(DCACHE_addr[20]), .B(n8225), .S0(n3624), .Y(\i_MIPS/n447 )
         );
  MX2XL U3485 ( .A(DCACHE_addr[7]), .B(n8244), .S0(n3624), .Y(\i_MIPS/n460 )
         );
  MX2XL U3486 ( .A(DCACHE_addr[22]), .B(n8164), .S0(n3624), .Y(\i_MIPS/n445 )
         );
  MX2XL U3487 ( .A(DCACHE_addr[19]), .B(n8162), .S0(n3624), .Y(\i_MIPS/n448 )
         );
  MX2XL U3488 ( .A(DCACHE_addr[23]), .B(n8039), .S0(n3624), .Y(\i_MIPS/n444 )
         );
  OA22XL U3489 ( .A0(n3292), .A1(n1858), .B0(n3245), .B1(n924), .Y(n7418) );
  OA22XL U3490 ( .A0(n3470), .A1(n1859), .B0(n3423), .B1(n925), .Y(n7416) );
  OA22XL U3491 ( .A0(n3379), .A1(n1860), .B0(n3337), .B1(n926), .Y(n7417) );
  OA22XL U3492 ( .A0(n3292), .A1(n853), .B0(n3245), .B1(n1786), .Y(n7428) );
  OA22XL U3493 ( .A0(n3470), .A1(n854), .B0(n3423), .B1(n1787), .Y(n7426) );
  OA22XL U3494 ( .A0(n3379), .A1(n855), .B0(n3337), .B1(n1788), .Y(n7427) );
  OA22XL U3495 ( .A0(n3292), .A1(n856), .B0(n3245), .B1(n1789), .Y(n7433) );
  OA22XL U3496 ( .A0(n3470), .A1(n857), .B0(n3423), .B1(n1790), .Y(n7431) );
  OA22XL U3497 ( .A0(n3379), .A1(n858), .B0(n3337), .B1(n1791), .Y(n7432) );
  OA22XL U3498 ( .A0(n3292), .A1(n1861), .B0(n3245), .B1(n927), .Y(n7423) );
  OA22XL U3499 ( .A0(n3470), .A1(n1862), .B0(n3423), .B1(n928), .Y(n7421) );
  OA22XL U3500 ( .A0(n3379), .A1(n1863), .B0(n3337), .B1(n929), .Y(n7422) );
  OA22XL U3501 ( .A0(n3293), .A1(n859), .B0(n3246), .B1(n1792), .Y(n7500) );
  OA22XL U3502 ( .A0(n3471), .A1(n860), .B0(n3424), .B1(n1793), .Y(n7498) );
  OA22XL U3503 ( .A0(n3380), .A1(n861), .B0(n3338), .B1(n1794), .Y(n7499) );
  OA22XL U3504 ( .A0(n3293), .A1(n1864), .B0(n3246), .B1(n930), .Y(n7490) );
  OA22XL U3505 ( .A0(n3471), .A1(n1865), .B0(n3424), .B1(n931), .Y(n7488) );
  OA22XL U3506 ( .A0(n3380), .A1(n1866), .B0(n3338), .B1(n932), .Y(n7489) );
  OA22XL U3507 ( .A0(n3293), .A1(n862), .B0(n3246), .B1(n1795), .Y(n7505) );
  OA22XL U3508 ( .A0(n3471), .A1(n863), .B0(n3424), .B1(n1796), .Y(n7503) );
  OA22XL U3509 ( .A0(n3380), .A1(n864), .B0(n3338), .B1(n1797), .Y(n7504) );
  OA22XL U3510 ( .A0(n3293), .A1(n1867), .B0(n3246), .B1(n933), .Y(n7495) );
  OA22XL U3511 ( .A0(n3471), .A1(n865), .B0(n3424), .B1(n1798), .Y(n7493) );
  OA22XL U3512 ( .A0(n3380), .A1(n1868), .B0(n3338), .B1(n934), .Y(n7494) );
  OA22XL U3513 ( .A0(n3301), .A1(n1869), .B0(n3254), .B1(n935), .Y(n8102) );
  OA22XL U3514 ( .A0(n3479), .A1(n1870), .B0(n3432), .B1(n936), .Y(n8100) );
  OA22XL U3515 ( .A0(n3388), .A1(n1871), .B0(n3346), .B1(n937), .Y(n8101) );
  OA22XL U3516 ( .A0(n3301), .A1(n866), .B0(n3254), .B1(n1799), .Y(n8112) );
  OA22XL U3517 ( .A0(n3479), .A1(n867), .B0(n3432), .B1(n1800), .Y(n8110) );
  OA22XL U3518 ( .A0(n3388), .A1(n868), .B0(n3346), .B1(n1801), .Y(n8111) );
  OA22XL U3519 ( .A0(n3301), .A1(n869), .B0(n3254), .B1(n1802), .Y(n8118) );
  OA22XL U3520 ( .A0(n3479), .A1(n870), .B0(n3432), .B1(n1803), .Y(n8116) );
  OA22XL U3521 ( .A0(n3388), .A1(n871), .B0(n3346), .B1(n1804), .Y(n8117) );
  OA22XL U3522 ( .A0(n3301), .A1(n1872), .B0(n3254), .B1(n938), .Y(n8107) );
  OA22XL U3523 ( .A0(n3479), .A1(n872), .B0(n3432), .B1(n1805), .Y(n8105) );
  OA22XL U3524 ( .A0(n3388), .A1(n1873), .B0(n3346), .B1(n939), .Y(n8106) );
  OA22XL U3525 ( .A0(n3297), .A1(n873), .B0(n3250), .B1(n1806), .Y(n7650) );
  OA22XL U3526 ( .A0(n3475), .A1(n874), .B0(n3428), .B1(n1807), .Y(n7648) );
  OA22XL U3527 ( .A0(n3384), .A1(n875), .B0(n3342), .B1(n1808), .Y(n7649) );
  OA22XL U3528 ( .A0(n3297), .A1(n1874), .B0(n3250), .B1(n940), .Y(n7640) );
  OA22XL U3529 ( .A0(n3475), .A1(n1875), .B0(n3428), .B1(n941), .Y(n7638) );
  OA22XL U3530 ( .A0(n3384), .A1(n1876), .B0(n3342), .B1(n942), .Y(n7639) );
  OA22XL U3531 ( .A0(n3297), .A1(n876), .B0(n3250), .B1(n1809), .Y(n7655) );
  OA22XL U3532 ( .A0(n3475), .A1(n877), .B0(n3428), .B1(n1810), .Y(n7653) );
  OA22XL U3533 ( .A0(n3384), .A1(n878), .B0(n3342), .B1(n1811), .Y(n7654) );
  OA22XL U3534 ( .A0(n3297), .A1(n1877), .B0(n3250), .B1(n943), .Y(n7645) );
  OA22XL U3535 ( .A0(n3475), .A1(n879), .B0(n3428), .B1(n1812), .Y(n7643) );
  OA22XL U3536 ( .A0(n3384), .A1(n1878), .B0(n3342), .B1(n944), .Y(n7644) );
  OA22XL U3537 ( .A0(n3292), .A1(n1879), .B0(n3245), .B1(n945), .Y(n7442) );
  OA22XL U3538 ( .A0(n3470), .A1(n880), .B0(n3423), .B1(n1813), .Y(n7440) );
  OA22XL U3539 ( .A0(n3379), .A1(n881), .B0(n3337), .B1(n1814), .Y(n7441) );
  OA22XL U3540 ( .A0(n3293), .A1(n882), .B0(n3246), .B1(n1815), .Y(n7481) );
  OA22XL U3541 ( .A0(n3471), .A1(n883), .B0(n3424), .B1(n1816), .Y(n7479) );
  OA22XL U3542 ( .A0(n3380), .A1(n884), .B0(n3338), .B1(n1817), .Y(n7480) );
  OA22XL U3543 ( .A0(n3287), .A1(n885), .B0(n3240), .B1(n1818), .Y(n4582) );
  OA22XL U3544 ( .A0(n3464), .A1(n886), .B0(n3416), .B1(n1819), .Y(n4580) );
  OA22XL U3545 ( .A0(n3375), .A1(n887), .B0(n3332), .B1(n1820), .Y(n4581) );
  OA22XL U3546 ( .A0(n3287), .A1(n888), .B0(n3240), .B1(n1821), .Y(n4572) );
  OA22XL U3547 ( .A0(n3464), .A1(n889), .B0(n3416), .B1(n1822), .Y(n4570) );
  OA22XL U3548 ( .A0(n3375), .A1(n890), .B0(n3332), .B1(n1823), .Y(n4571) );
  OA22XL U3549 ( .A0(n3287), .A1(n891), .B0(n3240), .B1(n1824), .Y(n4577) );
  OA22XL U3550 ( .A0(n3464), .A1(n892), .B0(n3416), .B1(n1825), .Y(n4575) );
  OA22XL U3551 ( .A0(n3375), .A1(n893), .B0(n3332), .B1(n1826), .Y(n4576) );
  INVXL U3552 ( .A(\D_cache/N98 ), .Y(n8768) );
  OAI2BB1XL U3553 ( .A0N(n3051), .A1N(n8426), .B0(n8392), .Y(n8393) );
  AO21X1 U3554 ( .A0(\i_MIPS/Register/n104 ), .A1(\i_MIPS/Register/n105 ), 
        .B0(n2883), .Y(n8334) );
  AOI2BB2XL U3555 ( .B0(\i_MIPS/IF_ID[77] ), .B1(n2157), .A0N(n3595), .A1N(
        \i_MIPS/n192 ), .Y(n8219) );
  AND3X4 U3556 ( .A(n2830), .B(n2161), .C(n7827), .Y(n2904) );
  AOI22XL U3557 ( .A0(\D_cache/N134 ), .A1(n2153), .B0(n3032), .B1(
        \D_cache/N166 ), .Y(\D_cache/n190 ) );
  CLKMX2X3 U3558 ( .A(\i_MIPS/n289 ), .B(n2989), .S0(n4018), .Y(n4691) );
  INVXL U3559 ( .A(n2708), .Y(n6920) );
  OAI21X4 U3560 ( .A0(n7086), .A1(\i_MIPS/n335 ), .B0(n3622), .Y(n7828) );
  INVXL U3561 ( .A(n8200), .Y(n8198) );
  INVXL U3562 ( .A(n8215), .Y(n8213) );
  INVXL U3563 ( .A(n7959), .Y(n7957) );
  INVXL U3564 ( .A(n7972), .Y(n7971) );
  INVXL U3565 ( .A(n7990), .Y(n7988) );
  INVXL U3566 ( .A(n8030), .Y(n8028) );
  INVXL U3567 ( .A(n8073), .Y(n8072) );
  INVXL U3568 ( .A(n8093), .Y(n8092) );
  INVXL U3569 ( .A(n7835), .Y(n7826) );
  INVXL U3570 ( .A(n7857), .Y(n7855) );
  INVXL U3571 ( .A(n7876), .Y(n7874) );
  INVXL U3572 ( .A(n7888), .Y(n7886) );
  INVXL U3573 ( .A(n7904), .Y(n7902) );
  INVXL U3574 ( .A(n7924), .Y(n7922) );
  INVXL U3575 ( .A(n7939), .Y(n7937) );
  NAND2X2 U3576 ( .A(\i_MIPS/ALUin1[8] ), .B(n4667), .Y(n6191) );
  NAND2XL U3577 ( .A(\i_MIPS/ALUOp[0] ), .B(n967), .Y(n4620) );
  AOI2BB2XL U3578 ( .B0(\i_MIPS/IF_ID[71] ), .B1(n2157), .A0N(n3595), .A1N(
        \i_MIPS/n186 ), .Y(n8361) );
  AOI2BB2XL U3579 ( .B0(\D_cache/N137 ), .B1(n2153), .A0N(n23), .A1N(n8887), 
        .Y(\D_cache/n193 ) );
  NAND4X2 U3580 ( .A(n4781), .B(n4780), .C(n4779), .D(n4778), .Y(n7071) );
  XOR2XL U3581 ( .A(n7632), .B(\i_MIPS/IR_ID[17] ), .Y(n4780) );
  XOR2XL U3582 ( .A(n4774), .B(\i_MIPS/IR_ID[23] ), .Y(n4743) );
  XOR2XL U3583 ( .A(n7632), .B(\i_MIPS/IR_ID[22] ), .Y(n4741) );
  XNOR2X1 U3584 ( .A(n2996), .B(n4013), .Y(n2794) );
  NOR4X2 U3585 ( .A(n4777), .B(n4776), .C(\i_MIPS/n372 ), .D(n4775), .Y(n4778)
         );
  NAND3X2 U3586 ( .A(\D_cache/n540 ), .B(\D_cache/n541 ), .C(\D_cache/n542 ), 
        .Y(\D_cache/n536 ) );
  NAND2BX4 U3587 ( .AN(n2989), .B(n4835), .Y(n2796) );
  AO22XL U3588 ( .A0(n2159), .A1(n7794), .B0(n3073), .B1(\i_MIPS/IR_ID[31] ), 
        .Y(\i_MIPS/N86 ) );
  AO22XL U3589 ( .A0(n2159), .A1(n7796), .B0(n3073), .B1(\i_MIPS/IR_ID[30] ), 
        .Y(\i_MIPS/N85 ) );
  AO22XL U3590 ( .A0(n2159), .A1(n7795), .B0(n3073), .B1(\i_MIPS/IR_ID[29] ), 
        .Y(\i_MIPS/N84 ) );
  AO22XL U3591 ( .A0(n2160), .A1(n7838), .B0(n3073), .B1(\i_MIPS/IR_ID[28] ), 
        .Y(\i_MIPS/N83 ) );
  AO22XL U3592 ( .A0(n2160), .A1(n7837), .B0(n3073), .B1(\i_MIPS/IR_ID[27] ), 
        .Y(\i_MIPS/N82 ) );
  AO22XL U3593 ( .A0(n2160), .A1(n7797), .B0(n3073), .B1(\i_MIPS/IR_ID[26] ), 
        .Y(\i_MIPS/N81 ) );
  AO22XL U3594 ( .A0(n2161), .A1(n8074), .B0(n3073), .B1(n4015), .Y(
        \i_MIPS/N75 ) );
  AO22XL U3595 ( .A0(n2161), .A1(n8419), .B0(n3073), .B1(\i_MIPS/IR_ID[19] ), 
        .Y(\i_MIPS/N74 ) );
  AO22XL U3596 ( .A0(n2161), .A1(n8050), .B0(n3073), .B1(n7164), .Y(
        \i_MIPS/N73 ) );
  AO22XL U3597 ( .A0(n2160), .A1(n8031), .B0(n3073), .B1(n7091), .Y(
        \i_MIPS/N72 ) );
  AO22XL U3598 ( .A0(n2159), .A1(n8004), .B0(n3073), .B1(\i_MIPS/IR_ID[16] ), 
        .Y(\i_MIPS/N71 ) );
  AOI2BB2XL U3599 ( .B0(\i_MIPS/IF_ID[70] ), .B1(n2157), .A0N(n3595), .A1N(
        \i_MIPS/n185 ), .Y(n8375) );
  AOI2BB2XL U3600 ( .B0(\i_MIPS/IF_ID[68] ), .B1(n2157), .A0N(n3595), .A1N(
        \i_MIPS/n183 ), .Y(n8343) );
  AOI2BB2XL U3601 ( .B0(\i_MIPS/IF_ID[69] ), .B1(n2157), .A0N(n3595), .A1N(
        \i_MIPS/n184 ), .Y(n8390) );
  AOI2BB2XL U3602 ( .B0(\i_MIPS/IF_ID[67] ), .B1(n2157), .A0N(n3595), .A1N(
        \i_MIPS/n182 ), .Y(n8405) );
  OA22X1 U3603 ( .A0(n8422), .A1(n3599), .B0(n8420), .B1(n2158), .Y(n8423) );
  OA22XL U3604 ( .A0(n3463), .A1(n1078), .B0(n3440), .B1(n166), .Y(n4489) );
  OA22XL U3605 ( .A0(n3463), .A1(n1079), .B0(n3440), .B1(n167), .Y(n4485) );
  OA22XL U3606 ( .A0(n3462), .A1(n1080), .B0(n3441), .B1(n168), .Y(n4453) );
  OA22XL U3607 ( .A0(n3462), .A1(n1081), .B0(n3441), .B1(n169), .Y(n4457) );
  OA22XL U3608 ( .A0(n3463), .A1(n162), .B0(n3439), .B1(n1052), .Y(n4501) );
  OA22XL U3609 ( .A0(n3462), .A1(n163), .B0(n3441), .B1(n1053), .Y(n4465) );
  OA22XL U3610 ( .A0(n3463), .A1(n164), .B0(n3437), .B1(n1054), .Y(n4497) );
  OA22X4 U3611 ( .A0(n3456), .A1(n997), .B0(n3412), .B1(n109), .Y(n4408) );
  OA22X4 U3612 ( .A0(n3455), .A1(n998), .B0(n3442), .B1(n110), .Y(n4404) );
  OA22X4 U3613 ( .A0(n3454), .A1(n999), .B0(n3410), .B1(n111), .Y(n4398) );
  OA22X4 U3614 ( .A0(n3453), .A1(n1000), .B0(n3409), .B1(n112), .Y(n4394) );
  OA22X4 U3615 ( .A0(n3487), .A1(n1001), .B0(n3414), .B1(n113), .Y(n4441) );
  OA22X4 U3616 ( .A0(n3482), .A1(n1002), .B0(n3414), .B1(n114), .Y(n4445) );
  OA21XL U3617 ( .A0(\i_MIPS/ALUin1[15] ), .A1(n3092), .B0(n5040), .Y(n5041)
         );
  AOI2BB1XL U3618 ( .A0N(\i_MIPS/ALUin1[16] ), .A1N(n3092), .B0(n2880), .Y(
        n4712) );
  OA21XL U3619 ( .A0(\i_MIPS/ALUin1[19] ), .A1(n3086), .B0(n5465), .Y(n5466)
         );
  AOI2BB1XL U3620 ( .A0N(n5825), .A1N(n8), .B0(n2903), .Y(n4721) );
  INVXL U3621 ( .A(n6825), .Y(n4719) );
  OAI221XL U3622 ( .A0(\i_MIPS/ALUin1[11] ), .A1(n3091), .B0(
        \i_MIPS/ALUin1[10] ), .B1(n3086), .C0(n5039), .Y(n5320) );
  OA22XL U3623 ( .A0(\i_MIPS/ALUin1[9] ), .A1(n14), .B0(\i_MIPS/ALUin1[8] ), 
        .B1(n3078), .Y(n5039) );
  OAI221XL U3624 ( .A0(\i_MIPS/ALUin1[11] ), .A1(n3082), .B0(
        \i_MIPS/ALUin1[10] ), .B1(n3077), .C0(n4911), .Y(n5203) );
  AOI2BB1XL U3625 ( .A0N(\i_MIPS/ALUin1[12] ), .A1N(n3087), .B0(n2879), .Y(
        n4911) );
  INVX1 U3626 ( .A(\i_MIPS/ID_EX[83] ), .Y(n5483) );
  NAND2XL U3627 ( .A(\i_MIPS/ALUin1[21] ), .B(n4640), .Y(n6474) );
  NAND2XL U3628 ( .A(\i_MIPS/ALUin1[24] ), .B(n4627), .Y(n5989) );
  XOR2XL U3629 ( .A(\i_MIPS/Reg_W[3] ), .B(\i_MIPS/IR_ID[24] ), .Y(n4766) );
  XOR2XL U3630 ( .A(\i_MIPS/Reg_W[1] ), .B(\i_MIPS/IR_ID[17] ), .Y(n4803) );
  XOR2XL U3631 ( .A(\i_MIPS/Reg_W[1] ), .B(\i_MIPS/IR_ID[22] ), .Y(n4765) );
  AOI2BB1XL U3632 ( .A0N(\i_MIPS/ALUin1[16] ), .A1N(n3078), .B0(n2844), .Y(
        n4815) );
  AO21X1 U3633 ( .A0(n3090), .A1(\i_MIPS/ALU/N303 ), .B0(n5122), .Y(n6477) );
  NAND2XL U3634 ( .A(n8316), .B(ICACHE_addr[28]), .Y(n8317) );
  XOR2XL U3635 ( .A(\i_MIPS/Reg_W[2] ), .B(\i_MIPS/IR_ID[18] ), .Y(n4802) );
  NAND2XL U3636 ( .A(n2863), .B(\i_MIPS/ALUin1[1] ), .Y(n5042) );
  OAI211XL U3637 ( .A0(n7001), .A1(n7000), .B0(n6999), .C0(n6998), .Y(n7017)
         );
  OA22XL U3638 ( .A0(n6997), .A1(n6996), .B0(n6996), .B1(n6995), .Y(n6998) );
  AOI32XL U3639 ( .A0(n6993), .A1(\i_MIPS/ALUin1[30] ), .A2(n6992), .B0(n6991), 
        .B1(n6990), .Y(n6999) );
  AOI2BB1XL U3640 ( .A0N(n6994), .A1N(n8), .B0(n2899), .Y(n6997) );
  NAND2XL U3641 ( .A(\i_MIPS/ALUin1[22] ), .B(n4632), .Y(n5981) );
  NAND2XL U3642 ( .A(n3088), .B(\i_MIPS/ALUin1[7] ), .Y(n5463) );
  NAND2XL U3643 ( .A(n3094), .B(\i_MIPS/ALUin1[8] ), .Y(n5118) );
  NAND2XL U3644 ( .A(\i_MIPS/ALUin1[25] ), .B(n4626), .Y(n5474) );
  NAND2XL U3645 ( .A(n3080), .B(\i_MIPS/ALUin1[30] ), .Y(n6995) );
  NAND2XL U3646 ( .A(\i_MIPS/ALU/N303 ), .B(n4723), .Y(n8526) );
  XOR2XL U3647 ( .A(\i_MIPS/Pred_1bit/current_state ), .B(n2862), .Y(
        \i_MIPS/Pred_1bit/n2 ) );
  AND2X1 U3648 ( .A(\i_MIPS/IR_ID[21] ), .B(\i_MIPS/n229 ), .Y(n2981) );
  AND2X1 U3649 ( .A(\i_MIPS/IR_ID[16] ), .B(\i_MIPS/n314 ), .Y(n2979) );
  MX2X1 U3650 ( .A(\i_MIPS/n247 ), .B(n2884), .S0(n4018), .Y(n4723) );
  AND2X1 U3651 ( .A(\i_MIPS/IR_ID[19] ), .B(\i_MIPS/n316 ), .Y(n2974) );
  AND2X1 U3652 ( .A(\i_MIPS/IR_ID[23] ), .B(\i_MIPS/n231 ), .Y(n2975) );
  OA22XL U3653 ( .A0(\i_MIPS/Register/register[4][21] ), .A1(n3179), .B0(
        \i_MIPS/Register/register[12][21] ), .B1(n3178), .Y(n6512) );
  OA22XL U3654 ( .A0(\i_MIPS/Register/register[0][21] ), .A1(n3187), .B0(
        \i_MIPS/Register/register[8][21] ), .B1(n3184), .Y(n6511) );
  OAI211XL U3655 ( .A0(\i_MIPS/ALUin1[16] ), .A1(n3087), .B0(n4914), .C0(n4913), .Y(n5202) );
  OAI211XL U3656 ( .A0(\i_MIPS/ALUin1[15] ), .A1(n3087), .B0(n5456), .C0(n5455), .Y(n5822) );
  AOI2BB1XL U3657 ( .A0N(\i_MIPS/ALUin1[17] ), .A1N(n3078), .B0(n2878), .Y(
        n5455) );
  OA22XL U3658 ( .A0(\i_MIPS/Register/register[20][4] ), .A1(n3129), .B0(
        \i_MIPS/Register/register[28][4] ), .B1(n3126), .Y(n5353) );
  OA22XL U3659 ( .A0(\i_MIPS/Register/register[16][4] ), .A1(n3135), .B0(
        \i_MIPS/Register/register[24][4] ), .B1(n3133), .Y(n5352) );
  OA22XL U3660 ( .A0(\i_MIPS/Register/register[20][18] ), .A1(n3129), .B0(
        \i_MIPS/Register/register[28][18] ), .B1(n3127), .Y(n5777) );
  OA22XL U3661 ( .A0(\i_MIPS/Register/register[16][18] ), .A1(n3135), .B0(
        \i_MIPS/Register/register[24][18] ), .B1(n3132), .Y(n5776) );
  OA22XL U3662 ( .A0(\i_MIPS/Register/register[20][13] ), .A1(n3181), .B0(
        \i_MIPS/Register/register[28][13] ), .B1(n3178), .Y(n6449) );
  OA22XL U3663 ( .A0(\i_MIPS/Register/register[16][13] ), .A1(n3187), .B0(
        \i_MIPS/Register/register[24][13] ), .B1(n3184), .Y(n6448) );
  OA22XL U3664 ( .A0(\i_MIPS/Register/register[20][12] ), .A1(n3130), .B0(
        \i_MIPS/Register/register[28][12] ), .B1(n3126), .Y(n6293) );
  OA22XL U3665 ( .A0(\i_MIPS/Register/register[16][12] ), .A1(n3136), .B0(
        \i_MIPS/Register/register[24][12] ), .B1(n3133), .Y(n6292) );
  OA22XL U3666 ( .A0(\i_MIPS/Register/register[20][21] ), .A1(n3181), .B0(
        \i_MIPS/Register/register[28][21] ), .B1(n3178), .Y(n6521) );
  OA22XL U3667 ( .A0(\i_MIPS/Register/register[16][21] ), .A1(n3187), .B0(
        \i_MIPS/Register/register[24][21] ), .B1(n3184), .Y(n6520) );
  OA22XL U3668 ( .A0(\i_MIPS/Register/register[16][22] ), .A1(n3134), .B0(
        \i_MIPS/Register/register[24][22] ), .B1(n3132), .Y(n6741) );
  AOI2BB1XL U3669 ( .A0N(\i_MIPS/ALUin1[15] ), .A1N(n3078), .B0(n2878), .Y(
        n4985) );
  NAND2XL U3670 ( .A(n7978), .B(ICACHE_addr[13]), .Y(n7964) );
  NAND2XL U3671 ( .A(n7943), .B(ICACHE_addr[11]), .Y(n7929) );
  OR3X2 U3672 ( .A(n7312), .B(\i_MIPS/n326 ), .C(\i_MIPS/IR_ID[29] ), .Y(n7313) );
  OAI221XL U3673 ( .A0(\i_MIPS/ALUin1[12] ), .A1(n3091), .B0(
        \i_MIPS/ALUin1[11] ), .B1(n3085), .C0(n5119), .Y(n5397) );
  OA22XL U3674 ( .A0(\i_MIPS/ALUin1[10] ), .A1(n14), .B0(\i_MIPS/ALUin1[9] ), 
        .B1(n3078), .Y(n5119) );
  OAI221XL U3675 ( .A0(\i_MIPS/ALUin1[22] ), .A1(n3091), .B0(
        \i_MIPS/ALUin1[23] ), .B1(n3085), .C0(n5460), .Y(n5816) );
  OA22XL U3676 ( .A0(\i_MIPS/ALUin1[24] ), .A1(n14), .B0(\i_MIPS/ALUin1[25] ), 
        .B1(n3077), .Y(n5460) );
  OA22XL U3677 ( .A0(n3467), .A1(n448), .B0(n3415), .B1(n1362), .Y(n4541) );
  OA22XL U3678 ( .A0(n3467), .A1(n449), .B0(n3420), .B1(n1363), .Y(n7316) );
  OA22XL U3679 ( .A0(n3549), .A1(n640), .B0(n3508), .B1(n1559), .Y(n4549) );
  OA22XL U3680 ( .A0(\i_MIPS/ALUin1[7] ), .A1(n3082), .B0(\i_MIPS/ALUin1[6] ), 
        .B1(n3078), .Y(n4910) );
  OA22XL U3681 ( .A0(\i_MIPS/ALUin1[22] ), .A1(n3082), .B0(\i_MIPS/ALUin1[23] ), .B1(n3078), .Y(n4711) );
  OA22XL U3682 ( .A0(\i_MIPS/ALUin1[21] ), .A1(n14), .B0(\i_MIPS/ALUin1[22] ), 
        .B1(n3078), .Y(n6049) );
  AND2XL U3683 ( .A(n3083), .B(\i_MIPS/ALUin1[29] ), .Y(n2899) );
  AND2XL U3684 ( .A(n3079), .B(\i_MIPS/ALUin1[0] ), .Y(n2986) );
  AND2XL U3685 ( .A(n3084), .B(\i_MIPS/ALUin1[2] ), .Y(n2900) );
  OA22XL U3686 ( .A0(\i_MIPS/Register/register[4][0] ), .A1(n3179), .B0(
        \i_MIPS/Register/register[12][0] ), .B1(n2785), .Y(n5091) );
  AND2XL U3687 ( .A(n2863), .B(\i_MIPS/ALUin1[30] ), .Y(n2903) );
  MX2X1 U3688 ( .A(n1882), .B(n3034), .S0(n3626), .Y(\i_MIPS/n407 ) );
  MX2X1 U3689 ( .A(\i_MIPS/ID_EX[57] ), .B(n3021), .S0(n3626), .Y(
        \i_MIPS/n405 ) );
  NAND2XL U3690 ( .A(n7816), .B(ICACHE_addr[7]), .Y(n7817) );
  NAND2XL U3691 ( .A(n7822), .B(n10), .Y(n7823) );
  OA22XL U3692 ( .A0(\i_MIPS/Register/register[22][28] ), .A1(n3116), .B0(
        \i_MIPS/Register/register[30][28] ), .B1(n3115), .Y(n5921) );
  OA22XL U3693 ( .A0(\i_MIPS/Register/register[6][28] ), .A1(n3118), .B0(
        \i_MIPS/Register/register[14][28] ), .B1(n3115), .Y(n5912) );
  OA22XL U3694 ( .A0(\i_MIPS/Register/register[22][28] ), .A1(n3172), .B0(
        \i_MIPS/Register/register[30][28] ), .B1(n3168), .Y(n5944) );
  OA22XL U3695 ( .A0(\i_MIPS/Register/register[6][28] ), .A1(n3171), .B0(
        \i_MIPS/Register/register[14][28] ), .B1(n3168), .Y(n5935) );
  OA22XL U3696 ( .A0(\i_MIPS/Register/register[22][31] ), .A1(n3170), .B0(
        \i_MIPS/Register/register[30][31] ), .B1(n3169), .Y(n4791) );
  OA22XL U3697 ( .A0(\i_MIPS/Register/register[6][31] ), .A1(n3170), .B0(
        \i_MIPS/Register/register[14][31] ), .B1(n3167), .Y(n4782) );
  OA22XL U3698 ( .A0(\i_MIPS/Register/register[22][31] ), .A1(n3116), .B0(
        \i_MIPS/Register/register[30][31] ), .B1(n3113), .Y(n4753) );
  OA22XL U3699 ( .A0(\i_MIPS/Register/register[6][31] ), .A1(n3116), .B0(
        \i_MIPS/Register/register[14][31] ), .B1(n3113), .Y(n4744) );
  OA22XL U3700 ( .A0(\i_MIPS/Register/register[22][30] ), .A1(n3170), .B0(
        \i_MIPS/Register/register[30][30] ), .B1(n3168), .Y(n7058) );
  OA22XL U3701 ( .A0(\i_MIPS/Register/register[6][30] ), .A1(n3170), .B0(
        \i_MIPS/Register/register[14][30] ), .B1(n3169), .Y(n7049) );
  OA22XL U3702 ( .A0(\i_MIPS/Register/register[22][30] ), .A1(n3118), .B0(
        \i_MIPS/Register/register[30][30] ), .B1(n3115), .Y(n7031) );
  OA22XL U3703 ( .A0(\i_MIPS/Register/register[6][30] ), .A1(n3118), .B0(
        \i_MIPS/Register/register[14][30] ), .B1(n2782), .Y(n7022) );
  OAI221XL U3704 ( .A0(\i_MIPS/ALUin1[21] ), .A1(n3091), .B0(
        \i_MIPS/ALUin1[22] ), .B1(n3085), .C0(n5887), .Y(n5958) );
  OA22XL U3705 ( .A0(\i_MIPS/ALUin1[23] ), .A1(n14), .B0(\i_MIPS/ALUin1[24] ), 
        .B1(n3077), .Y(n5887) );
  OAI2BB2XL U3706 ( .B0(\D_cache/n298 ), .B1(n3785), .A0N(
        \D_cache/cache[7][103] ), .A1N(\D_cache/n206 ), .Y(\D_cache/n965 ) );
  OAI2BB2XL U3707 ( .B0(\D_cache/n298 ), .B1(n3805), .A0N(
        \D_cache/cache[6][103] ), .A1N(\D_cache/n207 ), .Y(\D_cache/n966 ) );
  OAI2BB2XL U3708 ( .B0(\D_cache/n298 ), .B1(n3824), .A0N(
        \D_cache/cache[5][103] ), .A1N(n3838), .Y(\D_cache/n967 ) );
  OAI2BB2XL U3709 ( .B0(\D_cache/n298 ), .B1(n3858), .A0N(
        \D_cache/cache[4][103] ), .A1N(\D_cache/n209 ), .Y(\D_cache/n968 ) );
  OAI2BB2XL U3710 ( .B0(\D_cache/n298 ), .B1(n3864), .A0N(
        \D_cache/cache[3][103] ), .A1N(n3863), .Y(\D_cache/n969 ) );
  OAI2BB2XL U3711 ( .B0(\D_cache/n298 ), .B1(n3885), .A0N(
        \D_cache/cache[2][103] ), .A1N(\D_cache/n211 ), .Y(\D_cache/n970 ) );
  OAI2BB2XL U3712 ( .B0(\D_cache/n298 ), .B1(n3905), .A0N(
        \D_cache/cache[1][103] ), .A1N(\D_cache/n212 ), .Y(\D_cache/n971 ) );
  OAI2BB2XL U3713 ( .B0(\D_cache/n298 ), .B1(n3925), .A0N(
        \D_cache/cache[0][103] ), .A1N(n3930), .Y(\D_cache/n972 ) );
  CLKBUFX3 U3714 ( .A(\i_MIPS/EX_MEM_1 ), .Y(n4022) );
  XOR2XL U3715 ( .A(n8402), .B(ICACHE_addr[0]), .Y(n8401) );
  NAND2XL U3716 ( .A(\i_MIPS/ALUin1[28] ), .B(n4704), .Y(n5890) );
  NAND2XL U3717 ( .A(\i_MIPS/ALUin1[30] ), .B(n6992), .Y(n6988) );
  XOR2XL U3718 ( .A(\i_MIPS/Reg_W[2] ), .B(\i_MIPS/IR_ID[23] ), .Y(n4768) );
  XOR2XL U3719 ( .A(\i_MIPS/Reg_W[0] ), .B(\i_MIPS/IR_ID[16] ), .Y(n4804) );
  XOR2XL U3720 ( .A(\i_MIPS/Reg_W[0] ), .B(\i_MIPS/IR_ID[21] ), .Y(n4767) );
  MXI2XL U3721 ( .A(\i_MIPS/n258 ), .B(\i_MIPS/n259 ), .S0(n3622), .Y(
        \i_MIPS/n386 ) );
  MXI2XL U3722 ( .A(\i_MIPS/n254 ), .B(\i_MIPS/n255 ), .S0(n3622), .Y(
        \i_MIPS/n382 ) );
  MXI2XL U3723 ( .A(\i_MIPS/n250 ), .B(\i_MIPS/n251 ), .S0(n3622), .Y(
        \i_MIPS/n378 ) );
  MXI2XL U3724 ( .A(n2990), .B(\i_MIPS/n221 ), .S0(n3626), .Y(\i_MIPS/n503 )
         );
  MXI2XL U3725 ( .A(\i_MIPS/n308 ), .B(\i_MIPS/n309 ), .S0(n3620), .Y(
        \i_MIPS/n436 ) );
  MXI2XL U3726 ( .A(\i_MIPS/n306 ), .B(\i_MIPS/n307 ), .S0(n3620), .Y(
        \i_MIPS/n434 ) );
  MXI2XL U3727 ( .A(\i_MIPS/n304 ), .B(\i_MIPS/n305 ), .S0(n3620), .Y(
        \i_MIPS/n432 ) );
  MXI2XL U3728 ( .A(\i_MIPS/n302 ), .B(\i_MIPS/n303 ), .S0(n3620), .Y(
        \i_MIPS/n430 ) );
  MXI2XL U3729 ( .A(\i_MIPS/n300 ), .B(\i_MIPS/n301 ), .S0(n3620), .Y(
        \i_MIPS/n428 ) );
  MXI2XL U3730 ( .A(\i_MIPS/n298 ), .B(\i_MIPS/n299 ), .S0(n3620), .Y(
        \i_MIPS/n426 ) );
  MXI2XL U3731 ( .A(\i_MIPS/n294 ), .B(\i_MIPS/n295 ), .S0(n3620), .Y(
        \i_MIPS/n422 ) );
  MXI2XL U3732 ( .A(\i_MIPS/n282 ), .B(\i_MIPS/n283 ), .S0(n3626), .Y(
        \i_MIPS/n410 ) );
  MXI2XL U3733 ( .A(\i_MIPS/n280 ), .B(\i_MIPS/n281 ), .S0(n3621), .Y(
        \i_MIPS/n408 ) );
  MXI2XL U3734 ( .A(\i_MIPS/n278 ), .B(\i_MIPS/n279 ), .S0(n3624), .Y(
        \i_MIPS/n406 ) );
  MXI2XL U3735 ( .A(\i_MIPS/n246 ), .B(\i_MIPS/n247 ), .S0(n3625), .Y(
        \i_MIPS/n374 ) );
  MXI2XL U3736 ( .A(n2989), .B(\i_MIPS/n222 ), .S0(n3622), .Y(\i_MIPS/n502 )
         );
  XOR2XL U3737 ( .A(\i_MIPS/n228 ), .B(\i_MIPS/ID_EX[111] ), .Y(n7084) );
  MXI2XL U3738 ( .A(\i_MIPS/n342 ), .B(n8299), .S0(n3622), .Y(\i_MIPS/n533 )
         );
  MXI2XL U3739 ( .A(\i_MIPS/n371 ), .B(n8262), .S0(n3622), .Y(\i_MIPS/n562 )
         );
  MXI2XL U3740 ( .A(\i_MIPS/n327 ), .B(\i_MIPS/n326 ), .S0(n3622), .Y(
        \i_MIPS/n520 ) );
  MXI2XL U3741 ( .A(\i_MIPS/n325 ), .B(\i_MIPS/n324 ), .S0(n3622), .Y(
        \i_MIPS/n519 ) );
  MXI2XL U3742 ( .A(\i_MIPS/n323 ), .B(\i_MIPS/n322 ), .S0(n3622), .Y(
        \i_MIPS/n518 ) );
  MXI2XL U3743 ( .A(n2991), .B(\i_MIPS/n223 ), .S0(n3622), .Y(\i_MIPS/n501 )
         );
  XOR2XL U3744 ( .A(\i_MIPS/ID_EX[114] ), .B(\i_MIPS/IR_ID[19] ), .Y(
        \i_MIPS/Hazard_detection/n11 ) );
  XOR2XL U3745 ( .A(\i_MIPS/ID_EX[112] ), .B(\i_MIPS/IR_ID[17] ), .Y(
        \i_MIPS/Hazard_detection/n12 ) );
  XOR2XL U3746 ( .A(\i_MIPS/ID_EX[115] ), .B(n4015), .Y(
        \i_MIPS/Hazard_detection/n13 ) );
  XOR2XL U3747 ( .A(\i_MIPS/ID_EX[114] ), .B(\i_MIPS/IR_ID[24] ), .Y(
        \i_MIPS/Hazard_detection/n8 ) );
  XOR2XL U3748 ( .A(\i_MIPS/ID_EX[112] ), .B(\i_MIPS/IR_ID[22] ), .Y(
        \i_MIPS/Hazard_detection/n9 ) );
  XOR2XL U3749 ( .A(n4013), .B(\i_MIPS/ID_EX[115] ), .Y(
        \i_MIPS/Hazard_detection/n10 ) );
  XOR2XL U3750 ( .A(\i_MIPS/n230 ), .B(\i_MIPS/ID_EX[113] ), .Y(n7085) );
  XOR2XL U3751 ( .A(\i_MIPS/n316 ), .B(\i_MIPS/ID_EX[113] ), .Y(n7083) );
  MXI2XL U3752 ( .A(\i_MIPS/n348 ), .B(n8228), .S0(n3619), .Y(\i_MIPS/n539 )
         );
  MXI2XL U3753 ( .A(\i_MIPS/n349 ), .B(n8226), .S0(n3618), .Y(\i_MIPS/n540 )
         );
  XOR2XL U3754 ( .A(\i_MIPS/n312 ), .B(\i_MIPS/ID_EX[111] ), .Y(n7082) );
  MXI2XL U3755 ( .A(n8), .B(\i_MIPS/n219 ), .S0(n3623), .Y(\i_MIPS/n505 ) );
  MXI2XL U3756 ( .A(n2993), .B(\i_MIPS/n225 ), .S0(n3623), .Y(\i_MIPS/n499 )
         );
  MXI2XL U3757 ( .A(n2994), .B(\i_MIPS/n226 ), .S0(n3623), .Y(\i_MIPS/n498 )
         );
  MXI2XL U3758 ( .A(\i_MIPS/n367 ), .B(n8385), .S0(n3619), .Y(\i_MIPS/n558 )
         );
  MXI2XL U3759 ( .A(\i_MIPS/n356 ), .B(n8254), .S0(n3621), .Y(\i_MIPS/n547 )
         );
  MXI2XL U3760 ( .A(\i_MIPS/n366 ), .B(n8370), .S0(n3619), .Y(\i_MIPS/n557 )
         );
  MXI2XL U3761 ( .A(\i_MIPS/n341 ), .B(n8312), .S0(n3623), .Y(\i_MIPS/n532 )
         );
  MXI2XL U3762 ( .A(\i_MIPS/n357 ), .B(n8252), .S0(n3618), .Y(\i_MIPS/n548 )
         );
  MXI2XL U3763 ( .A(\i_MIPS/n358 ), .B(n8250), .S0(n3618), .Y(\i_MIPS/n549 )
         );
  MXI2XL U3764 ( .A(\i_MIPS/n354 ), .B(n8256), .S0(n3617), .Y(\i_MIPS/n545 )
         );
  MXI2XL U3765 ( .A(\i_MIPS/n343 ), .B(n8282), .S0(n3619), .Y(\i_MIPS/n534 )
         );
  MXI2XL U3766 ( .A(\i_MIPS/n344 ), .B(n8458), .S0(n3620), .Y(\i_MIPS/n535 )
         );
  MXI2XL U3767 ( .A(\i_MIPS/n369 ), .B(n8400), .S0(n3619), .Y(\i_MIPS/n560 )
         );
  MXI2XL U3768 ( .A(\i_MIPS/n370 ), .B(n8239), .S0(n3619), .Y(\i_MIPS/n561 )
         );
  MXI2XL U3769 ( .A(\i_MIPS/n368 ), .B(n8338), .S0(n3619), .Y(\i_MIPS/n559 )
         );
  MXI2XL U3770 ( .A(\i_MIPS/n365 ), .B(n8356), .S0(n3617), .Y(\i_MIPS/n556 )
         );
  MXI2XL U3771 ( .A(\i_MIPS/n355 ), .B(n7976), .S0(n3617), .Y(\i_MIPS/n546 )
         );
  MXI2XL U3772 ( .A(\i_MIPS/n353 ), .B(n1086), .S0(n3617), .Y(\i_MIPS/n544 )
         );
  MXI2XL U3773 ( .A(\i_MIPS/n329 ), .B(\i_MIPS/n328 ), .S0(n3617), .Y(
        \i_MIPS/n521 ) );
  AND2X1 U3774 ( .A(\D_cache/n518 ), .B(mem_ready_D), .Y(\D_cache/n246 ) );
  NAND2XL U3775 ( .A(\i_MIPS/ALU/N303 ), .B(n4707), .Y(n4730) );
  MX2X1 U3776 ( .A(n2946), .B(n2947), .S0(n10321), .Y(\D_cache/N131 ) );
  MX4XL U3777 ( .A(\D_cache/cache[0][53] ), .B(\D_cache/cache[1][53] ), .C(
        \D_cache/cache[2][53] ), .D(\D_cache/cache[3][53] ), .S0(n2138), .S1(
        n2425), .Y(n2946) );
  MX4XL U3778 ( .A(\D_cache/cache[4][53] ), .B(\D_cache/cache[5][53] ), .C(
        \D_cache/cache[6][53] ), .D(\D_cache/cache[7][53] ), .S0(n2061), .S1(
        n2432), .Y(n2947) );
  MX2X1 U3779 ( .A(n2958), .B(n2959), .S0(n4041), .Y(\D_cache/N128 ) );
  MX4XL U3780 ( .A(\D_cache/cache[0][56] ), .B(\D_cache/cache[1][56] ), .C(
        \D_cache/cache[2][56] ), .D(\D_cache/cache[3][56] ), .S0(n2070), .S1(
        n2415), .Y(n2958) );
  MX4XL U3781 ( .A(\D_cache/cache[4][56] ), .B(\D_cache/cache[5][56] ), .C(
        \D_cache/cache[6][56] ), .D(\D_cache/cache[7][56] ), .S0(n2068), .S1(
        n2416), .Y(n2959) );
  MX2X1 U3782 ( .A(n2910), .B(n2911), .S0(DCACHE_addr[4]), .Y(\D_cache/N139 )
         );
  MX4XL U3783 ( .A(\D_cache/cache[0][45] ), .B(\D_cache/cache[1][45] ), .C(
        \D_cache/cache[2][45] ), .D(\D_cache/cache[3][45] ), .S0(n2144), .S1(
        n2229), .Y(n2910) );
  MX4XL U3784 ( .A(\D_cache/cache[4][45] ), .B(\D_cache/cache[5][45] ), .C(
        \D_cache/cache[6][45] ), .D(\D_cache/cache[7][45] ), .S0(n2061), .S1(
        n2232), .Y(n2911) );
  MX2X1 U3785 ( .A(n2964), .B(n2965), .S0(n3062), .Y(\D_cache/N126 ) );
  MX4XL U3786 ( .A(\D_cache/cache[0][58] ), .B(\D_cache/cache[1][58] ), .C(
        \D_cache/cache[2][58] ), .D(\D_cache/cache[3][58] ), .S0(n2126), .S1(
        n2434), .Y(n2964) );
  MX4XL U3787 ( .A(\D_cache/cache[4][58] ), .B(\D_cache/cache[5][58] ), .C(
        \D_cache/cache[6][58] ), .D(\D_cache/cache[7][58] ), .S0(n2114), .S1(
        n2171), .Y(n2965) );
  MX2X1 U3788 ( .A(n2908), .B(n2909), .S0(n3063), .Y(\D_cache/N141 ) );
  MX4XL U3789 ( .A(\D_cache/cache[0][43] ), .B(\D_cache/cache[1][43] ), .C(
        \D_cache/cache[2][43] ), .D(\D_cache/cache[3][43] ), .S0(n2081), .S1(
        n2231), .Y(n2908) );
  MX4XL U3790 ( .A(\D_cache/cache[4][43] ), .B(\D_cache/cache[5][43] ), .C(
        \D_cache/cache[6][43] ), .D(\D_cache/cache[7][43] ), .S0(n2080), .S1(
        n2235), .Y(n2909) );
  MX2X1 U3791 ( .A(n2936), .B(n2937), .S0(n3065), .Y(\D_cache/N143 ) );
  MX4XL U3792 ( .A(\D_cache/cache[0][41] ), .B(\D_cache/cache[1][41] ), .C(
        \D_cache/cache[2][41] ), .D(\D_cache/cache[3][41] ), .S0(n2142), .S1(
        n2283), .Y(n2936) );
  MX4XL U3793 ( .A(\D_cache/cache[4][41] ), .B(\D_cache/cache[5][41] ), .C(
        \D_cache/cache[6][41] ), .D(\D_cache/cache[7][41] ), .S0(n2141), .S1(
        n2296), .Y(n2937) );
  MX2X1 U3794 ( .A(n2920), .B(n2921), .S0(n3065), .Y(\D_cache/N137 ) );
  MX4XL U3795 ( .A(\D_cache/cache[0][47] ), .B(\D_cache/cache[1][47] ), .C(
        \D_cache/cache[2][47] ), .D(\D_cache/cache[3][47] ), .S0(n2065), .S1(
        n2294), .Y(n2920) );
  MX4XL U3796 ( .A(\D_cache/cache[4][47] ), .B(\D_cache/cache[5][47] ), .C(
        \D_cache/cache[6][47] ), .D(\D_cache/cache[7][47] ), .S0(n2070), .S1(
        n2292), .Y(n2921) );
  MX2X1 U3797 ( .A(n2924), .B(n2925), .S0(n3067), .Y(\D_cache/N122 ) );
  MX4XL U3798 ( .A(\D_cache/cache[0][62] ), .B(\D_cache/cache[1][62] ), .C(
        \D_cache/cache[2][62] ), .D(\D_cache/cache[3][62] ), .S0(n2074), .S1(
        n2172), .Y(n2924) );
  MX4XL U3799 ( .A(\D_cache/cache[4][62] ), .B(\D_cache/cache[5][62] ), .C(
        \D_cache/cache[6][62] ), .D(\D_cache/cache[7][62] ), .S0(n2073), .S1(
        n2173), .Y(n2925) );
  MX2X1 U3800 ( .A(n2938), .B(n2939), .S0(n3062), .Y(\D_cache/N144 ) );
  MX4XL U3801 ( .A(\D_cache/cache[0][40] ), .B(\D_cache/cache[1][40] ), .C(
        \D_cache/cache[2][40] ), .D(\D_cache/cache[3][40] ), .S0(n2091), .S1(
        n2221), .Y(n2938) );
  MX4XL U3802 ( .A(\D_cache/cache[4][40] ), .B(\D_cache/cache[5][40] ), .C(
        \D_cache/cache[6][40] ), .D(\D_cache/cache[7][40] ), .S0(n2063), .S1(
        n2220), .Y(n2939) );
  MX2X1 U3803 ( .A(n2916), .B(n2917), .S0(n10321), .Y(\D_cache/N138 ) );
  MX4XL U3804 ( .A(\D_cache/cache[0][46] ), .B(\D_cache/cache[1][46] ), .C(
        \D_cache/cache[2][46] ), .D(\D_cache/cache[3][46] ), .S0(n2072), .S1(
        n2230), .Y(n2916) );
  MX4XL U3805 ( .A(\D_cache/cache[4][46] ), .B(\D_cache/cache[5][46] ), .C(
        \D_cache/cache[6][46] ), .D(\D_cache/cache[7][46] ), .S0(n2096), .S1(
        n2234), .Y(n2917) );
  MX2X1 U3806 ( .A(n2954), .B(n2955), .S0(n4041), .Y(\D_cache/N150 ) );
  MX4XL U3807 ( .A(\D_cache/cache[0][34] ), .B(\D_cache/cache[1][34] ), .C(
        \D_cache/cache[2][34] ), .D(\D_cache/cache[3][34] ), .S0(n2098), .S1(
        n2314), .Y(n2954) );
  MX4XL U3808 ( .A(\D_cache/cache[4][34] ), .B(\D_cache/cache[5][34] ), .C(
        \D_cache/cache[6][34] ), .D(\D_cache/cache[7][34] ), .S0(n2095), .S1(
        n2319), .Y(n2955) );
  AND2X1 U3809 ( .A(\i_MIPS/IR_ID[21] ), .B(\i_MIPS/IR_ID[22] ), .Y(n2982) );
  AND2X1 U3810 ( .A(\i_MIPS/IR_ID[16] ), .B(\i_MIPS/IR_ID[17] ), .Y(n2980) );
  AND2X1 U3811 ( .A(\i_MIPS/IR_ID[23] ), .B(\i_MIPS/IR_ID[24] ), .Y(n2976) );
  AND2X1 U3812 ( .A(\i_MIPS/IR_ID[18] ), .B(\i_MIPS/IR_ID[19] ), .Y(n2972) );
  AND2X1 U3813 ( .A(\i_MIPS/IR_ID[22] ), .B(\i_MIPS/n228 ), .Y(n2983) );
  OA22XL U3814 ( .A0(\i_MIPS/Register/register[20][20] ), .A1(n3128), .B0(
        \i_MIPS/Register/register[28][20] ), .B1(n3125), .Y(n4885) );
  OA22XL U3815 ( .A0(\i_MIPS/Register/register[16][20] ), .A1(n3134), .B0(
        \i_MIPS/Register/register[24][20] ), .B1(n3131), .Y(n4884) );
  NAND2XL U3816 ( .A(n7916), .B(ICACHE_addr[9]), .Y(n7917) );
  NAND2XL U3817 ( .A(n7846), .B(ICACHE_addr[5]), .Y(n7847) );
  MX2X1 U3818 ( .A(n2942), .B(n2943), .S0(n4041), .Y(\D_cache/N146 ) );
  MX4XL U3819 ( .A(\D_cache/cache[0][38] ), .B(\D_cache/cache[1][38] ), .C(
        \D_cache/cache[2][38] ), .D(\D_cache/cache[3][38] ), .S0(n2087), .S1(
        n2339), .Y(n2942) );
  MX4XL U3820 ( .A(\D_cache/cache[4][38] ), .B(\D_cache/cache[5][38] ), .C(
        \D_cache/cache[6][38] ), .D(\D_cache/cache[7][38] ), .S0(n2088), .S1(
        n2346), .Y(n2943) );
  MX2X1 U3821 ( .A(n2932), .B(n2933), .S0(n3067), .Y(\D_cache/N129 ) );
  MX4XL U3822 ( .A(\D_cache/cache[0][55] ), .B(\D_cache/cache[1][55] ), .C(
        \D_cache/cache[2][55] ), .D(\D_cache/cache[3][55] ), .S0(n2103), .S1(
        n2206), .Y(n2932) );
  MX4XL U3823 ( .A(\D_cache/cache[4][55] ), .B(\D_cache/cache[5][55] ), .C(
        \D_cache/cache[6][55] ), .D(\D_cache/cache[7][55] ), .S0(n2120), .S1(
        n2209), .Y(n2933) );
  MX2X1 U3824 ( .A(n2962), .B(n2963), .S0(n3067), .Y(\D_cache/N132 ) );
  MX4XL U3825 ( .A(\D_cache/cache[0][52] ), .B(\D_cache/cache[1][52] ), .C(
        \D_cache/cache[2][52] ), .D(\D_cache/cache[3][52] ), .S0(n2119), .S1(
        n2202), .Y(n2962) );
  MX4XL U3826 ( .A(\D_cache/cache[4][52] ), .B(\D_cache/cache[5][52] ), .C(
        \D_cache/cache[6][52] ), .D(\D_cache/cache[7][52] ), .S0(n2140), .S1(
        n2203), .Y(n2963) );
  MX2X1 U3827 ( .A(n2950), .B(n2951), .S0(n3064), .Y(\D_cache/N151 ) );
  MX4XL U3828 ( .A(\D_cache/cache[0][33] ), .B(\D_cache/cache[1][33] ), .C(
        \D_cache/cache[2][33] ), .D(\D_cache/cache[3][33] ), .S0(n2100), .S1(
        n2326), .Y(n2950) );
  MX4XL U3829 ( .A(\D_cache/cache[4][33] ), .B(\D_cache/cache[5][33] ), .C(
        \D_cache/cache[6][33] ), .D(\D_cache/cache[7][33] ), .S0(n2140), .S1(
        n2334), .Y(n2951) );
  MX2X1 U3830 ( .A(n2968), .B(n2969), .S0(n10321), .Y(\D_cache/N135 ) );
  MX4XL U3831 ( .A(\D_cache/cache[0][49] ), .B(\D_cache/cache[1][49] ), .C(
        \D_cache/cache[2][49] ), .D(\D_cache/cache[3][49] ), .S0(n2117), .S1(
        n2308), .Y(n2968) );
  MX4XL U3832 ( .A(\D_cache/cache[4][49] ), .B(\D_cache/cache[5][49] ), .C(
        \D_cache/cache[6][49] ), .D(\D_cache/cache[7][49] ), .S0(n2140), .S1(
        n2316), .Y(n2969) );
  MX2X1 U3833 ( .A(n2940), .B(n2941), .S0(n2146), .Y(\D_cache/N145 ) );
  MX4XL U3834 ( .A(\D_cache/cache[0][39] ), .B(\D_cache/cache[1][39] ), .C(
        \D_cache/cache[2][39] ), .D(\D_cache/cache[3][39] ), .S0(n2125), .S1(
        n2315), .Y(n2940) );
  MX4XL U3835 ( .A(\D_cache/cache[4][39] ), .B(\D_cache/cache[5][39] ), .C(
        \D_cache/cache[6][39] ), .D(\D_cache/cache[7][39] ), .S0(n2127), .S1(
        n2321), .Y(n2941) );
  MX2X1 U3836 ( .A(n2960), .B(n2961), .S0(n3064), .Y(\D_cache/N123 ) );
  MX4XL U3837 ( .A(\D_cache/cache[0][61] ), .B(\D_cache/cache[1][61] ), .C(
        \D_cache/cache[2][61] ), .D(\D_cache/cache[3][61] ), .S0(n2117), .S1(
        n2405), .Y(n2960) );
  MX4XL U3838 ( .A(\D_cache/cache[4][61] ), .B(\D_cache/cache[5][61] ), .C(
        \D_cache/cache[6][61] ), .D(\D_cache/cache[7][61] ), .S0(n2118), .S1(
        n2406), .Y(n2961) );
  MX4XL U3839 ( .A(\D_cache/cache[0][50] ), .B(\D_cache/cache[1][50] ), .C(
        \D_cache/cache[2][50] ), .D(\D_cache/cache[3][50] ), .S0(n2138), .S1(
        n2429), .Y(n2966) );
  MX4XL U3840 ( .A(\D_cache/cache[4][50] ), .B(\D_cache/cache[5][50] ), .C(
        \D_cache/cache[6][50] ), .D(\D_cache/cache[7][50] ), .S0(
        DCACHE_addr[2]), .S1(n2428), .Y(n2967) );
  MX2X1 U3841 ( .A(n2914), .B(n2915), .S0(n3064), .Y(\D_cache/N140 ) );
  MX4XL U3842 ( .A(\D_cache/cache[0][44] ), .B(\D_cache/cache[1][44] ), .C(
        \D_cache/cache[2][44] ), .D(\D_cache/cache[3][44] ), .S0(n2089), .S1(
        n2258), .Y(n2914) );
  MX4XL U3843 ( .A(\D_cache/cache[4][44] ), .B(\D_cache/cache[5][44] ), .C(
        \D_cache/cache[6][44] ), .D(\D_cache/cache[7][44] ), .S0(n2107), .S1(
        n2256), .Y(n2915) );
  MX2X1 U3844 ( .A(n2912), .B(n2913), .S0(DCACHE_addr[4]), .Y(\D_cache/N125 )
         );
  MX4XL U3845 ( .A(\D_cache/cache[0][59] ), .B(\D_cache/cache[1][59] ), .C(
        \D_cache/cache[2][59] ), .D(\D_cache/cache[3][59] ), .S0(n2138), .S1(
        n2177), .Y(n2912) );
  MX4XL U3846 ( .A(\D_cache/cache[4][59] ), .B(\D_cache/cache[5][59] ), .C(
        \D_cache/cache[6][59] ), .D(\D_cache/cache[7][59] ), .S0(n2105), .S1(
        n2179), .Y(n2913) );
  OAI221XL U3847 ( .A0(\i_MIPS/ALUin1[24] ), .A1(n3091), .B0(
        \i_MIPS/ALUin1[25] ), .B1(n3085), .C0(n4709), .Y(n6754) );
  OA22XL U3848 ( .A0(\i_MIPS/ALUin1[26] ), .A1(n14), .B0(\i_MIPS/ALUin1[27] ), 
        .B1(n3078), .Y(n4709) );
  MX4XL U3849 ( .A(\D_cache/cache[0][32] ), .B(\D_cache/cache[1][32] ), .C(
        \D_cache/cache[2][32] ), .D(\D_cache/cache[3][32] ), .S0(n2112), .S1(
        n2439), .Y(n2928) );
  MX4XL U3850 ( .A(\D_cache/cache[4][32] ), .B(\D_cache/cache[5][32] ), .C(
        \D_cache/cache[6][32] ), .D(\D_cache/cache[7][32] ), .S0(n2097), .S1(
        n2438), .Y(n2929) );
  MX2X1 U3851 ( .A(n2918), .B(n2919), .S0(n2146), .Y(\D_cache/N147 ) );
  MX4XL U3852 ( .A(\D_cache/cache[0][37] ), .B(\D_cache/cache[1][37] ), .C(
        \D_cache/cache[2][37] ), .D(\D_cache/cache[3][37] ), .S0(n2061), .S1(
        n2272), .Y(n2918) );
  MX4XL U3853 ( .A(\D_cache/cache[4][37] ), .B(\D_cache/cache[5][37] ), .C(
        \D_cache/cache[6][37] ), .D(\D_cache/cache[7][37] ), .S0(n2062), .S1(
        n2280), .Y(n2919) );
  MX2X1 U3854 ( .A(n2922), .B(n2923), .S0(n10321), .Y(\D_cache/N136 ) );
  MX4XL U3855 ( .A(\D_cache/cache[0][48] ), .B(\D_cache/cache[1][48] ), .C(
        \D_cache/cache[2][48] ), .D(\D_cache/cache[3][48] ), .S0(n2082), .S1(
        n2348), .Y(n2922) );
  MX4XL U3856 ( .A(\D_cache/cache[4][48] ), .B(\D_cache/cache[5][48] ), .C(
        \D_cache/cache[6][48] ), .D(\D_cache/cache[7][48] ), .S0(n2114), .S1(
        n2356), .Y(n2923) );
  MX2X1 U3857 ( .A(n2934), .B(n2935), .S0(n3065), .Y(\D_cache/N142 ) );
  MX4XL U3858 ( .A(\D_cache/cache[0][42] ), .B(\D_cache/cache[1][42] ), .C(
        \D_cache/cache[2][42] ), .D(\D_cache/cache[3][42] ), .S0(n2105), .S1(
        n2278), .Y(n2934) );
  MX4XL U3859 ( .A(\D_cache/cache[4][42] ), .B(\D_cache/cache[5][42] ), .C(
        \D_cache/cache[6][42] ), .D(\D_cache/cache[7][42] ), .S0(n2102), .S1(
        n2291), .Y(n2935) );
  MX2X1 U3860 ( .A(n2952), .B(n2953), .S0(n2147), .Y(\D_cache/N127 ) );
  MX4XL U3861 ( .A(\D_cache/cache[0][57] ), .B(\D_cache/cache[1][57] ), .C(
        \D_cache/cache[2][57] ), .D(\D_cache/cache[3][57] ), .S0(n2066), .S1(
        n2338), .Y(n2952) );
  MX4XL U3862 ( .A(\D_cache/cache[4][57] ), .B(\D_cache/cache[5][57] ), .C(
        \D_cache/cache[6][57] ), .D(\D_cache/cache[7][57] ), .S0(n2114), .S1(
        n2344), .Y(n2953) );
  MX2X1 U3863 ( .A(n2956), .B(n2957), .S0(n3066), .Y(\D_cache/N149 ) );
  MX4XL U3864 ( .A(\D_cache/cache[0][35] ), .B(\D_cache/cache[1][35] ), .C(
        \D_cache/cache[2][35] ), .D(\D_cache/cache[3][35] ), .S0(n2118), .S1(
        n2236), .Y(n2956) );
  MX4XL U3865 ( .A(\D_cache/cache[4][35] ), .B(\D_cache/cache[5][35] ), .C(
        \D_cache/cache[6][35] ), .D(\D_cache/cache[7][35] ), .S0(n2108), .S1(
        n2244), .Y(n2957) );
  MX2X1 U3866 ( .A(n2970), .B(n2971), .S0(n3066), .Y(\D_cache/N133 ) );
  MX4XL U3867 ( .A(\D_cache/cache[0][51] ), .B(\D_cache/cache[1][51] ), .C(
        \D_cache/cache[2][51] ), .D(\D_cache/cache[3][51] ), .S0(n2062), .S1(
        n2357), .Y(n2970) );
  MX4XL U3868 ( .A(\D_cache/cache[4][51] ), .B(\D_cache/cache[5][51] ), .C(
        \D_cache/cache[6][51] ), .D(\D_cache/cache[7][51] ), .S0(n2081), .S1(
        n2359), .Y(n2971) );
  MX2X1 U3869 ( .A(n2926), .B(n2927), .S0(DCACHE_addr[4]), .Y(\D_cache/N130 )
         );
  MX4XL U3870 ( .A(\D_cache/cache[0][54] ), .B(\D_cache/cache[1][54] ), .C(
        \D_cache/cache[2][54] ), .D(\D_cache/cache[3][54] ), .S0(n2079), .S1(
        n2362), .Y(n2926) );
  MX4XL U3871 ( .A(\D_cache/cache[4][54] ), .B(\D_cache/cache[5][54] ), .C(
        \D_cache/cache[6][54] ), .D(\D_cache/cache[7][54] ), .S0(n2091), .S1(
        n2361), .Y(n2927) );
  MX2X1 U3872 ( .A(n2930), .B(n2931), .S0(n2147), .Y(\D_cache/N124 ) );
  MX4XL U3873 ( .A(\D_cache/cache[0][60] ), .B(\D_cache/cache[1][60] ), .C(
        \D_cache/cache[2][60] ), .D(\D_cache/cache[3][60] ), .S0(n2140), .S1(
        n2200), .Y(n2930) );
  MX4XL U3874 ( .A(\D_cache/cache[4][60] ), .B(\D_cache/cache[5][60] ), .C(
        \D_cache/cache[6][60] ), .D(\D_cache/cache[7][60] ), .S0(n2138), .S1(
        n2401), .Y(n2931) );
  MX2X1 U3875 ( .A(n2944), .B(n2945), .S0(n10321), .Y(\D_cache/N121 ) );
  MX4XL U3876 ( .A(\D_cache/cache[0][63] ), .B(\D_cache/cache[1][63] ), .C(
        \D_cache/cache[2][63] ), .D(\D_cache/cache[3][63] ), .S0(n2135), .S1(
        n2409), .Y(n2944) );
  MX4XL U3877 ( .A(\D_cache/cache[4][63] ), .B(\D_cache/cache[5][63] ), .C(
        \D_cache/cache[6][63] ), .D(\D_cache/cache[7][63] ), .S0(n2132), .S1(
        n2410), .Y(n2945) );
  MX2X1 U3878 ( .A(n2948), .B(n2949), .S0(DCACHE_addr[4]), .Y(\D_cache/N148 )
         );
  MX4XL U3879 ( .A(\D_cache/cache[0][36] ), .B(\D_cache/cache[1][36] ), .C(
        \D_cache/cache[2][36] ), .D(\D_cache/cache[3][36] ), .S0(n2087), .S1(
        n2270), .Y(n2948) );
  MX4XL U3880 ( .A(\D_cache/cache[4][36] ), .B(\D_cache/cache[5][36] ), .C(
        \D_cache/cache[6][36] ), .D(\D_cache/cache[7][36] ), .S0(n2086), .S1(
        n2268), .Y(n2949) );
  OA22XL U3881 ( .A0(\i_MIPS/Register/register[20][14] ), .A1(n3181), .B0(
        \i_MIPS/Register/register[28][14] ), .B1(n3178), .Y(n6383) );
  OA22XL U3882 ( .A0(\i_MIPS/Register/register[4][14] ), .A1(n3179), .B0(
        \i_MIPS/Register/register[12][14] ), .B1(n3178), .Y(n6374) );
  OA22XL U3883 ( .A0(\i_MIPS/Register/register[4][4] ), .A1(n3129), .B0(
        \i_MIPS/Register/register[12][4] ), .B1(n3126), .Y(n5344) );
  OA22XL U3884 ( .A0(\i_MIPS/Register/register[4][18] ), .A1(n3128), .B0(
        \i_MIPS/Register/register[12][18] ), .B1(n3127), .Y(n5768) );
  OA22XL U3885 ( .A0(\i_MIPS/Register/register[4][13] ), .A1(n3179), .B0(
        \i_MIPS/Register/register[12][13] ), .B1(n3178), .Y(n6440) );
  OA22XL U3886 ( .A0(\i_MIPS/Register/register[20][3] ), .A1(n3130), .B0(
        \i_MIPS/Register/register[28][3] ), .B1(n2787), .Y(n6571) );
  OA22XL U3887 ( .A0(\i_MIPS/Register/register[4][3] ), .A1(n3130), .B0(
        \i_MIPS/Register/register[12][3] ), .B1(n3125), .Y(n6562) );
  OA22XL U3888 ( .A0(\i_MIPS/Register/register[20][3] ), .A1(n2786), .B0(
        \i_MIPS/Register/register[28][3] ), .B1(n3178), .Y(n6592) );
  OA22XL U3889 ( .A0(\i_MIPS/Register/register[4][3] ), .A1(n2786), .B0(
        \i_MIPS/Register/register[12][3] ), .B1(n3178), .Y(n6583) );
  OA22XL U3890 ( .A0(\i_MIPS/Register/register[20][17] ), .A1(n3180), .B0(
        \i_MIPS/Register/register[28][17] ), .B1(n3177), .Y(n5726) );
  OA22XL U3891 ( .A0(\i_MIPS/Register/register[4][12] ), .A1(n3130), .B0(
        \i_MIPS/Register/register[12][12] ), .B1(n3127), .Y(n6284) );
  OA22XL U3892 ( .A0(\i_MIPS/Register/register[4][18] ), .A1(n3181), .B0(
        \i_MIPS/Register/register[12][18] ), .B1(n3177), .Y(n5789) );
  OA22XL U3893 ( .A0(\i_MIPS/Register/register[4][17] ), .A1(n3180), .B0(
        \i_MIPS/Register/register[12][17] ), .B1(n3177), .Y(n5717) );
  OA22XL U3894 ( .A0(\i_MIPS/Register/register[20][25] ), .A1(n3180), .B0(
        \i_MIPS/Register/register[28][25] ), .B1(n3176), .Y(n5528) );
  OA22XL U3895 ( .A0(\i_MIPS/Register/register[20][25] ), .A1(n3129), .B0(
        \i_MIPS/Register/register[28][25] ), .B1(n3126), .Y(n5505) );
  OA22XL U3896 ( .A0(\i_MIPS/Register/register[4][25] ), .A1(n3180), .B0(
        \i_MIPS/Register/register[12][25] ), .B1(n3176), .Y(n5519) );
  OA22XL U3897 ( .A0(\i_MIPS/Register/register[4][25] ), .A1(n3129), .B0(
        \i_MIPS/Register/register[12][25] ), .B1(n3126), .Y(n5496) );
  OA22XL U3898 ( .A0(\i_MIPS/Register/register[20][21] ), .A1(n3130), .B0(
        \i_MIPS/Register/register[28][21] ), .B1(n3126), .Y(n6498) );
  OA22XL U3899 ( .A0(\i_MIPS/Register/register[4][21] ), .A1(n3130), .B0(
        \i_MIPS/Register/register[12][21] ), .B1(n3127), .Y(n6489) );
  OA22XL U3900 ( .A0(\i_MIPS/Register/register[20][26] ), .A1(n3180), .B0(
        \i_MIPS/Register/register[28][26] ), .B1(n3177), .Y(n6115) );
  OA22XL U3901 ( .A0(\i_MIPS/Register/register[4][26] ), .A1(n3180), .B0(
        \i_MIPS/Register/register[12][26] ), .B1(n3177), .Y(n6106) );
  OA22XL U3902 ( .A0(\i_MIPS/Register/register[20][26] ), .A1(n3129), .B0(
        \i_MIPS/Register/register[28][26] ), .B1(n3127), .Y(n6092) );
  OA22XL U3903 ( .A0(\i_MIPS/Register/register[4][26] ), .A1(n3128), .B0(
        \i_MIPS/Register/register[12][26] ), .B1(n3127), .Y(n6083) );
  OA22XL U3904 ( .A0(\i_MIPS/Register/register[20][19] ), .A1(n3129), .B0(
        \i_MIPS/Register/register[28][19] ), .B1(n3126), .Y(n5643) );
  OA22XL U3905 ( .A0(\i_MIPS/Register/register[4][19] ), .A1(n3129), .B0(
        \i_MIPS/Register/register[12][19] ), .B1(n3126), .Y(n5634) );
  OA22XL U3906 ( .A0(\i_MIPS/Register/register[20][19] ), .A1(n3180), .B0(
        \i_MIPS/Register/register[28][19] ), .B1(n3176), .Y(n5666) );
  OA22XL U3907 ( .A0(\i_MIPS/Register/register[20][24] ), .A1(n3129), .B0(
        \i_MIPS/Register/register[28][24] ), .B1(n3127), .Y(n6017) );
  OA22XL U3908 ( .A0(\i_MIPS/Register/register[4][19] ), .A1(n3180), .B0(
        \i_MIPS/Register/register[12][19] ), .B1(n3176), .Y(n5657) );
  OA22XL U3909 ( .A0(\i_MIPS/Register/register[4][24] ), .A1(n3130), .B0(
        \i_MIPS/Register/register[12][24] ), .B1(n3127), .Y(n6008) );
  OA22XL U3910 ( .A0(\i_MIPS/Register/register[20][20] ), .A1(n3179), .B0(
        \i_MIPS/Register/register[28][20] ), .B1(n3176), .Y(n4862) );
  OA22XL U3911 ( .A0(\i_MIPS/Register/register[4][20] ), .A1(n3179), .B0(
        \i_MIPS/Register/register[12][20] ), .B1(n3178), .Y(n4853) );
  OA22XL U3912 ( .A0(\i_MIPS/Register/register[20][24] ), .A1(n3180), .B0(
        \i_MIPS/Register/register[28][24] ), .B1(n3177), .Y(n6040) );
  OA22XL U3913 ( .A0(\i_MIPS/Register/register[4][24] ), .A1(n3181), .B0(
        \i_MIPS/Register/register[12][24] ), .B1(n3177), .Y(n6031) );
  OA22XL U3914 ( .A0(\i_MIPS/Register/register[4][20] ), .A1(n3128), .B0(
        \i_MIPS/Register/register[12][20] ), .B1(n3125), .Y(n4876) );
  OA22XL U3915 ( .A0(\i_MIPS/Register/register[20][29] ), .A1(n3180), .B0(
        \i_MIPS/Register/register[28][29] ), .B1(n3177), .Y(n5878) );
  OA22XL U3916 ( .A0(\i_MIPS/Register/register[4][29] ), .A1(n3179), .B0(
        \i_MIPS/Register/register[12][29] ), .B1(n3177), .Y(n5869) );
  OA22XL U3917 ( .A0(\i_MIPS/Register/register[20][29] ), .A1(n3128), .B0(
        \i_MIPS/Register/register[28][29] ), .B1(n3127), .Y(n5855) );
  OA22XL U3918 ( .A0(\i_MIPS/Register/register[4][29] ), .A1(n3129), .B0(
        \i_MIPS/Register/register[12][29] ), .B1(n3127), .Y(n5846) );
  OA22XL U3919 ( .A0(\i_MIPS/Register/register[20][28] ), .A1(n2789), .B0(
        \i_MIPS/Register/register[28][28] ), .B1(n3127), .Y(n5928) );
  OA22XL U3920 ( .A0(\i_MIPS/Register/register[4][28] ), .A1(n2789), .B0(
        \i_MIPS/Register/register[12][28] ), .B1(n3127), .Y(n5919) );
  OA22XL U3921 ( .A0(\i_MIPS/Register/register[20][28] ), .A1(n3181), .B0(
        \i_MIPS/Register/register[28][28] ), .B1(n3177), .Y(n5951) );
  OA22XL U3922 ( .A0(\i_MIPS/Register/register[4][28] ), .A1(n3180), .B0(
        \i_MIPS/Register/register[12][28] ), .B1(n3177), .Y(n5942) );
  OA22XL U3923 ( .A0(\i_MIPS/Register/register[20][31] ), .A1(n3179), .B0(
        \i_MIPS/Register/register[28][31] ), .B1(n3176), .Y(n4798) );
  OA22XL U3924 ( .A0(\i_MIPS/Register/register[4][31] ), .A1(n3179), .B0(
        \i_MIPS/Register/register[12][31] ), .B1(n3178), .Y(n4789) );
  OA22XL U3925 ( .A0(\i_MIPS/Register/register[20][31] ), .A1(n3128), .B0(
        \i_MIPS/Register/register[28][31] ), .B1(n3125), .Y(n4760) );
  OA22XL U3926 ( .A0(\i_MIPS/Register/register[4][31] ), .A1(n3128), .B0(
        \i_MIPS/Register/register[12][31] ), .B1(n3125), .Y(n4751) );
  OA22XL U3927 ( .A0(\i_MIPS/Register/register[20][2] ), .A1(n3128), .B0(
        \i_MIPS/Register/register[28][2] ), .B1(n3127), .Y(n6643) );
  OA22XL U3928 ( .A0(\i_MIPS/Register/register[4][2] ), .A1(n3129), .B0(
        \i_MIPS/Register/register[12][2] ), .B1(n3125), .Y(n6634) );
  OA22XL U3929 ( .A0(\i_MIPS/Register/register[20][22] ), .A1(n3181), .B0(
        \i_MIPS/Register/register[28][22] ), .B1(n3176), .Y(n6721) );
  OA22XL U3930 ( .A0(\i_MIPS/Register/register[4][22] ), .A1(n3181), .B0(
        \i_MIPS/Register/register[12][22] ), .B1(n3178), .Y(n6712) );
  OA22XL U3931 ( .A0(\i_MIPS/Register/register[4][22] ), .A1(n3128), .B0(
        \i_MIPS/Register/register[12][22] ), .B1(n3126), .Y(n6733) );
  OA22XL U3932 ( .A0(\i_MIPS/Register/register[4][23] ), .A1(n3181), .B0(
        \i_MIPS/Register/register[12][23] ), .B1(n3176), .Y(n6865) );
  OA22XL U3933 ( .A0(\i_MIPS/Register/register[20][27] ), .A1(n3181), .B0(
        \i_MIPS/Register/register[28][27] ), .B1(n3177), .Y(n6818) );
  OA22XL U3934 ( .A0(\i_MIPS/Register/register[4][27] ), .A1(n3181), .B0(
        \i_MIPS/Register/register[12][27] ), .B1(n3176), .Y(n6809) );
  OA22XL U3935 ( .A0(\i_MIPS/Register/register[20][27] ), .A1(n3130), .B0(
        \i_MIPS/Register/register[28][27] ), .B1(n3127), .Y(n6795) );
  OA22XL U3936 ( .A0(\i_MIPS/Register/register[4][27] ), .A1(n3128), .B0(
        \i_MIPS/Register/register[12][27] ), .B1(n2787), .Y(n6786) );
  OA22XL U3937 ( .A0(\i_MIPS/Register/register[20][30] ), .A1(n3181), .B0(
        \i_MIPS/Register/register[28][30] ), .B1(n3177), .Y(n7065) );
  OA22XL U3938 ( .A0(\i_MIPS/Register/register[4][30] ), .A1(n3181), .B0(
        \i_MIPS/Register/register[12][30] ), .B1(n3178), .Y(n7056) );
  OA22XL U3939 ( .A0(\i_MIPS/Register/register[20][30] ), .A1(n3130), .B0(
        \i_MIPS/Register/register[28][30] ), .B1(n3125), .Y(n7038) );
  OA22XL U3940 ( .A0(\i_MIPS/Register/register[4][30] ), .A1(n3129), .B0(
        \i_MIPS/Register/register[12][30] ), .B1(n3125), .Y(n7029) );
  OA22XL U3941 ( .A0(\i_MIPS/Register/register[16][14] ), .A1(n3187), .B0(
        \i_MIPS/Register/register[24][14] ), .B1(n3184), .Y(n6382) );
  OA22XL U3942 ( .A0(\i_MIPS/Register/register[0][14] ), .A1(n3187), .B0(
        \i_MIPS/Register/register[8][14] ), .B1(n3184), .Y(n6373) );
  OA22XL U3943 ( .A0(\i_MIPS/Register/register[0][15] ), .A1(n3135), .B0(
        \i_MIPS/Register/register[8][15] ), .B1(n3132), .Y(n5562) );
  OA22XL U3944 ( .A0(\i_MIPS/Register/register[0][4] ), .A1(n3135), .B0(
        \i_MIPS/Register/register[8][4] ), .B1(n3132), .Y(n5343) );
  OA22XL U3945 ( .A0(\i_MIPS/Register/register[0][18] ), .A1(n3134), .B0(
        \i_MIPS/Register/register[8][18] ), .B1(n3132), .Y(n5767) );
  OA22XL U3946 ( .A0(\i_MIPS/Register/register[0][13] ), .A1(n3187), .B0(
        \i_MIPS/Register/register[8][13] ), .B1(n3184), .Y(n6439) );
  OA22XL U3947 ( .A0(\i_MIPS/Register/register[0][0] ), .A1(n2764), .B0(
        \i_MIPS/Register/register[8][0] ), .B1(n3183), .Y(n5090) );
  OA22XL U3948 ( .A0(\i_MIPS/Register/register[0][4] ), .A1(n3185), .B0(
        \i_MIPS/Register/register[8][4] ), .B1(n3182), .Y(n5364) );
  OA22XL U3949 ( .A0(\i_MIPS/Register/register[16][3] ), .A1(n3136), .B0(
        \i_MIPS/Register/register[24][3] ), .B1(n3133), .Y(n6570) );
  OA22XL U3950 ( .A0(\i_MIPS/Register/register[0][3] ), .A1(n3136), .B0(
        \i_MIPS/Register/register[8][3] ), .B1(n3133), .Y(n6561) );
  OA22XL U3951 ( .A0(\i_MIPS/Register/register[0][12] ), .A1(n3136), .B0(
        \i_MIPS/Register/register[8][12] ), .B1(n3133), .Y(n6283) );
  OA22XL U3952 ( .A0(\i_MIPS/Register/register[16][3] ), .A1(n3187), .B0(
        \i_MIPS/Register/register[24][3] ), .B1(n3184), .Y(n6591) );
  OA22XL U3953 ( .A0(\i_MIPS/Register/register[0][3] ), .A1(n3187), .B0(
        \i_MIPS/Register/register[8][3] ), .B1(n3184), .Y(n6582) );
  OA22XL U3954 ( .A0(\i_MIPS/Register/register[16][17] ), .A1(n3186), .B0(
        \i_MIPS/Register/register[24][17] ), .B1(n3183), .Y(n5725) );
  OA22XL U3955 ( .A0(\i_MIPS/Register/register[0][18] ), .A1(n3186), .B0(
        \i_MIPS/Register/register[8][18] ), .B1(n3183), .Y(n5788) );
  OA22XL U3956 ( .A0(\i_MIPS/Register/register[0][17] ), .A1(n3186), .B0(
        \i_MIPS/Register/register[8][17] ), .B1(n3183), .Y(n5716) );
  OA22XL U3957 ( .A0(\i_MIPS/Register/register[16][25] ), .A1(n3185), .B0(
        \i_MIPS/Register/register[24][25] ), .B1(n3182), .Y(n5527) );
  OA22XL U3958 ( .A0(\i_MIPS/Register/register[16][25] ), .A1(n3135), .B0(
        \i_MIPS/Register/register[24][25] ), .B1(n3131), .Y(n5504) );
  OA22XL U3959 ( .A0(\i_MIPS/Register/register[0][25] ), .A1(n3185), .B0(
        \i_MIPS/Register/register[8][25] ), .B1(n3182), .Y(n5518) );
  OA22XL U3960 ( .A0(\i_MIPS/Register/register[0][25] ), .A1(n3135), .B0(
        \i_MIPS/Register/register[8][25] ), .B1(n3133), .Y(n5495) );
  OA22XL U3961 ( .A0(\i_MIPS/Register/register[16][21] ), .A1(n3136), .B0(
        \i_MIPS/Register/register[24][21] ), .B1(n3133), .Y(n6497) );
  OA22XL U3962 ( .A0(\i_MIPS/Register/register[0][21] ), .A1(n3136), .B0(
        \i_MIPS/Register/register[8][21] ), .B1(n3133), .Y(n6488) );
  OA22XL U3963 ( .A0(\i_MIPS/Register/register[16][26] ), .A1(n3186), .B0(
        \i_MIPS/Register/register[24][26] ), .B1(n3183), .Y(n6114) );
  OA22XL U3964 ( .A0(\i_MIPS/Register/register[0][26] ), .A1(n3186), .B0(
        \i_MIPS/Register/register[8][26] ), .B1(n3183), .Y(n6105) );
  OA22XL U3965 ( .A0(\i_MIPS/Register/register[16][26] ), .A1(n3135), .B0(
        \i_MIPS/Register/register[24][26] ), .B1(n3132), .Y(n6091) );
  OA22XL U3966 ( .A0(\i_MIPS/Register/register[0][26] ), .A1(n3134), .B0(
        \i_MIPS/Register/register[8][26] ), .B1(n3132), .Y(n6082) );
  OA22XL U3967 ( .A0(\i_MIPS/Register/register[16][19] ), .A1(n3135), .B0(
        \i_MIPS/Register/register[24][19] ), .B1(n3133), .Y(n5642) );
  OA22XL U3968 ( .A0(\i_MIPS/Register/register[0][19] ), .A1(n3135), .B0(
        \i_MIPS/Register/register[8][19] ), .B1(n3132), .Y(n5633) );
  OA22XL U3969 ( .A0(\i_MIPS/Register/register[16][19] ), .A1(n3185), .B0(
        \i_MIPS/Register/register[24][19] ), .B1(n3182), .Y(n5665) );
  OA22XL U3970 ( .A0(\i_MIPS/Register/register[16][24] ), .A1(n3135), .B0(
        \i_MIPS/Register/register[24][24] ), .B1(n3132), .Y(n6016) );
  OA22XL U3971 ( .A0(\i_MIPS/Register/register[0][19] ), .A1(n3185), .B0(
        \i_MIPS/Register/register[8][19] ), .B1(n3182), .Y(n5656) );
  OA22XL U3972 ( .A0(\i_MIPS/Register/register[0][24] ), .A1(n3136), .B0(
        \i_MIPS/Register/register[8][24] ), .B1(n3132), .Y(n6007) );
  OA22XL U3973 ( .A0(\i_MIPS/Register/register[16][20] ), .A1(n3185), .B0(
        \i_MIPS/Register/register[24][20] ), .B1(n3184), .Y(n4861) );
  OA22XL U3974 ( .A0(\i_MIPS/Register/register[0][20] ), .A1(n3186), .B0(
        \i_MIPS/Register/register[8][20] ), .B1(n3183), .Y(n4852) );
  OA22XL U3975 ( .A0(\i_MIPS/Register/register[16][24] ), .A1(n3186), .B0(
        \i_MIPS/Register/register[24][24] ), .B1(n3183), .Y(n6039) );
  OA22XL U3976 ( .A0(\i_MIPS/Register/register[0][24] ), .A1(n3186), .B0(
        \i_MIPS/Register/register[8][24] ), .B1(n3183), .Y(n6030) );
  OA22XL U3977 ( .A0(\i_MIPS/Register/register[0][20] ), .A1(n3134), .B0(
        \i_MIPS/Register/register[8][20] ), .B1(n3131), .Y(n4875) );
  OA22XL U3978 ( .A0(\i_MIPS/Register/register[16][29] ), .A1(n3186), .B0(
        \i_MIPS/Register/register[24][29] ), .B1(n3183), .Y(n5877) );
  OA22XL U3979 ( .A0(\i_MIPS/Register/register[0][29] ), .A1(n3186), .B0(
        \i_MIPS/Register/register[8][29] ), .B1(n3183), .Y(n5868) );
  OA22XL U3980 ( .A0(\i_MIPS/Register/register[16][29] ), .A1(n3134), .B0(
        \i_MIPS/Register/register[24][29] ), .B1(n3132), .Y(n5854) );
  OA22XL U3981 ( .A0(\i_MIPS/Register/register[0][29] ), .A1(n3135), .B0(
        \i_MIPS/Register/register[8][29] ), .B1(n3132), .Y(n5845) );
  OA22XL U3982 ( .A0(\i_MIPS/Register/register[16][28] ), .A1(n2763), .B0(
        \i_MIPS/Register/register[24][28] ), .B1(n3132), .Y(n5927) );
  OA22XL U3983 ( .A0(\i_MIPS/Register/register[0][28] ), .A1(n2763), .B0(
        \i_MIPS/Register/register[8][28] ), .B1(n3132), .Y(n5918) );
  OA22XL U3984 ( .A0(\i_MIPS/Register/register[16][28] ), .A1(n3186), .B0(
        \i_MIPS/Register/register[24][28] ), .B1(n3183), .Y(n5950) );
  OA22XL U3985 ( .A0(\i_MIPS/Register/register[0][28] ), .A1(n3186), .B0(
        \i_MIPS/Register/register[8][28] ), .B1(n3183), .Y(n5941) );
  OA22XL U3986 ( .A0(\i_MIPS/Register/register[16][31] ), .A1(n3187), .B0(
        \i_MIPS/Register/register[24][31] ), .B1(n3183), .Y(n4797) );
  OA22XL U3987 ( .A0(\i_MIPS/Register/register[0][31] ), .A1(n3185), .B0(
        \i_MIPS/Register/register[8][31] ), .B1(n3184), .Y(n4788) );
  OA22XL U3988 ( .A0(\i_MIPS/Register/register[16][31] ), .A1(n3134), .B0(
        \i_MIPS/Register/register[24][31] ), .B1(n3131), .Y(n4759) );
  OA22XL U3989 ( .A0(\i_MIPS/Register/register[0][31] ), .A1(n3134), .B0(
        \i_MIPS/Register/register[8][31] ), .B1(n3131), .Y(n4750) );
  OA22XL U3990 ( .A0(\i_MIPS/Register/register[16][2] ), .A1(n3134), .B0(
        \i_MIPS/Register/register[24][2] ), .B1(n3132), .Y(n6642) );
  OA22XL U3991 ( .A0(\i_MIPS/Register/register[0][2] ), .A1(n3135), .B0(
        \i_MIPS/Register/register[8][2] ), .B1(n3131), .Y(n6633) );
  OA22XL U3992 ( .A0(\i_MIPS/Register/register[16][22] ), .A1(n3187), .B0(
        \i_MIPS/Register/register[24][22] ), .B1(n3183), .Y(n6720) );
  OA22XL U3993 ( .A0(\i_MIPS/Register/register[0][22] ), .A1(n3185), .B0(
        \i_MIPS/Register/register[8][22] ), .B1(n3182), .Y(n6711) );
  OA22XL U3994 ( .A0(\i_MIPS/Register/register[0][22] ), .A1(n3135), .B0(
        \i_MIPS/Register/register[8][22] ), .B1(n3131), .Y(n6732) );
  OA22XL U3995 ( .A0(\i_MIPS/Register/register[0][23] ), .A1(n3185), .B0(
        \i_MIPS/Register/register[8][23] ), .B1(n3183), .Y(n6864) );
  OA22XL U3996 ( .A0(\i_MIPS/Register/register[16][27] ), .A1(n3186), .B0(
        \i_MIPS/Register/register[24][27] ), .B1(n3182), .Y(n6817) );
  OA22XL U3997 ( .A0(\i_MIPS/Register/register[0][27] ), .A1(n3185), .B0(
        \i_MIPS/Register/register[8][27] ), .B1(n2784), .Y(n6808) );
  OA22XL U3998 ( .A0(\i_MIPS/Register/register[16][27] ), .A1(n3136), .B0(
        \i_MIPS/Register/register[24][27] ), .B1(n3131), .Y(n6794) );
  OA22XL U3999 ( .A0(\i_MIPS/Register/register[0][27] ), .A1(n3134), .B0(
        \i_MIPS/Register/register[8][27] ), .B1(n3133), .Y(n6785) );
  OA22XL U4000 ( .A0(\i_MIPS/Register/register[16][30] ), .A1(n3187), .B0(
        \i_MIPS/Register/register[24][30] ), .B1(n3182), .Y(n7064) );
  OA22XL U4001 ( .A0(\i_MIPS/Register/register[0][30] ), .A1(n3186), .B0(
        \i_MIPS/Register/register[8][30] ), .B1(n2784), .Y(n7055) );
  OA22XL U4002 ( .A0(\i_MIPS/Register/register[16][30] ), .A1(n2763), .B0(
        \i_MIPS/Register/register[24][30] ), .B1(n3132), .Y(n7037) );
  OA22XL U4003 ( .A0(\i_MIPS/Register/register[0][30] ), .A1(n3136), .B0(
        \i_MIPS/Register/register[8][30] ), .B1(n3131), .Y(n7028) );
  OA22XL U4004 ( .A0(n3471), .A1(n641), .B0(n3415), .B1(n1560), .Y(n4545) );
  OA22XL U4005 ( .A0(n3467), .A1(n450), .B0(n3420), .B1(n1364), .Y(n7320) );
  OA22XL U4006 ( .A0(n3472), .A1(n642), .B0(n3425), .B1(n1561), .Y(n7536) );
  OA22XL U4007 ( .A0(n3468), .A1(n643), .B0(n3421), .B1(n1562), .Y(n7340) );
  OA22XL U4008 ( .A0(n3467), .A1(n644), .B0(n3420), .B1(n1563), .Y(n7336) );
  OA22XL U4009 ( .A0(n3467), .A1(n645), .B0(n3420), .B1(n1564), .Y(n7332) );
  OA22XL U4010 ( .A0(n3478), .A1(n646), .B0(n3431), .B1(n1565), .Y(n7765) );
  OA22XL U4011 ( .A0(n3478), .A1(n647), .B0(n3431), .B1(n1566), .Y(n7760) );
  OA22XL U4012 ( .A0(n3472), .A1(n648), .B0(n3425), .B1(n1567), .Y(n7527) );
  OA22XL U4013 ( .A0(n3469), .A1(n649), .B0(n3422), .B1(n1568), .Y(n7398) );
  OA22XL U4014 ( .A0(n3472), .A1(n650), .B0(n3425), .B1(n1569), .Y(n7522) );
  OA22XL U4015 ( .A0(n3473), .A1(n651), .B0(n3426), .B1(n1570), .Y(n7576) );
  OA22XL U4016 ( .A0(n3472), .A1(n652), .B0(n3425), .B1(n1571), .Y(n7517) );
  OA22XL U4017 ( .A0(n3469), .A1(n653), .B0(n3422), .B1(n1572), .Y(n7393) );
  OA22XL U4018 ( .A0(n3473), .A1(n654), .B0(n3426), .B1(n1573), .Y(n7571) );
  OA22XL U4019 ( .A0(n3469), .A1(n655), .B0(n3422), .B1(n1574), .Y(n7388) );
  OA22XL U4020 ( .A0(n3473), .A1(n656), .B0(n3426), .B1(n1575), .Y(n7566) );
  OA22XL U4021 ( .A0(n3473), .A1(n657), .B0(n3426), .B1(n1576), .Y(n7561) );
  OA22XL U4022 ( .A0(n3474), .A1(n658), .B0(n3427), .B1(n1577), .Y(n7615) );
  OA22XL U4023 ( .A0(n3474), .A1(n659), .B0(n3427), .B1(n1578), .Y(n7610) );
  OA22XL U4024 ( .A0(n3477), .A1(n660), .B0(n3430), .B1(n1579), .Y(n7701) );
  OA22XL U4025 ( .A0(n3477), .A1(n661), .B0(n3430), .B1(n1580), .Y(n7715) );
  OA22XL U4026 ( .A0(n3478), .A1(n662), .B0(n3431), .B1(n1581), .Y(n7751) );
  OA22XL U4027 ( .A0(n3477), .A1(n663), .B0(n3430), .B1(n1582), .Y(n7710) );
  OA22XL U4028 ( .A0(n3476), .A1(n664), .B0(n3429), .B1(n1583), .Y(n7692) );
  OA22XL U4029 ( .A0(n3478), .A1(n665), .B0(n3431), .B1(n1584), .Y(n7741) );
  OA22XL U4030 ( .A0(n3476), .A1(n666), .B0(n3429), .B1(n1585), .Y(n7687) );
  OA22XL U4031 ( .A0(n3476), .A1(n667), .B0(n3429), .B1(n1586), .Y(n7678) );
  OA22XL U4032 ( .A0(n3476), .A1(n668), .B0(n3429), .B1(n1587), .Y(n7673) );
  OA22XL U4033 ( .A0(n3476), .A1(n669), .B0(n3429), .B1(n1588), .Y(n7668) );
  OA22XL U4034 ( .A0(n3475), .A1(n670), .B0(n3428), .B1(n1589), .Y(n7663) );
  OA22XL U4035 ( .A0(n3474), .A1(n671), .B0(n3427), .B1(n1590), .Y(n7600) );
  OA22XL U4036 ( .A0(n3474), .A1(n672), .B0(n3427), .B1(n1591), .Y(n7590) );
  OA22XL U4037 ( .A0(n3473), .A1(n673), .B0(n3426), .B1(n1592), .Y(n7585) );
  OA22XL U4038 ( .A0(n3554), .A1(n674), .B0(n3512), .B1(n1593), .Y(n7359) );
  OA22XL U4039 ( .A0(n3554), .A1(n675), .B0(n3512), .B1(n1594), .Y(n7355) );
  OA22XL U4040 ( .A0(n3554), .A1(n676), .B0(n3512), .B1(n1595), .Y(n7351) );
  OA22XL U4041 ( .A0(n3554), .A1(n677), .B0(n3512), .B1(n1596), .Y(n7347) );
  OA22XL U4042 ( .A0(n3553), .A1(n678), .B0(n3511), .B1(n1597), .Y(n7297) );
  OA22XL U4043 ( .A0(\i_MIPS/Register/register[22][12] ), .A1(n3172), .B0(
        \i_MIPS/Register/register[30][12] ), .B1(n3169), .Y(n6307) );
  OA22XL U4044 ( .A0(\i_MIPS/Register/register[22][4] ), .A1(n3116), .B0(
        \i_MIPS/Register/register[30][4] ), .B1(n3114), .Y(n5346) );
  OA22XL U4045 ( .A0(\i_MIPS/Register/register[6][4] ), .A1(n3117), .B0(
        \i_MIPS/Register/register[14][4] ), .B1(n3114), .Y(n5337) );
  OA22XL U4046 ( .A0(\i_MIPS/Register/register[22][0] ), .A1(n3116), .B0(
        \i_MIPS/Register/register[30][0] ), .B1(n3113), .Y(n5072) );
  OA22XL U4047 ( .A0(\i_MIPS/Register/register[22][18] ), .A1(n3116), .B0(
        \i_MIPS/Register/register[30][18] ), .B1(n3115), .Y(n5770) );
  OA22XL U4048 ( .A0(\i_MIPS/Register/register[6][18] ), .A1(n3117), .B0(
        \i_MIPS/Register/register[14][18] ), .B1(n3115), .Y(n5761) );
  OA22XL U4049 ( .A0(\i_MIPS/Register/register[22][13] ), .A1(n3172), .B0(
        \i_MIPS/Register/register[30][13] ), .B1(n3169), .Y(n6442) );
  OA22XL U4050 ( .A0(\i_MIPS/Register/register[6][13] ), .A1(n3172), .B0(
        \i_MIPS/Register/register[14][13] ), .B1(n3169), .Y(n6433) );
  OA22XL U4051 ( .A0(\i_MIPS/Register/register[6][0] ), .A1(n3170), .B0(
        \i_MIPS/Register/register[14][0] ), .B1(n2773), .Y(n5084) );
  OA22XL U4052 ( .A0(\i_MIPS/Register/register[6][4] ), .A1(n3171), .B0(
        \i_MIPS/Register/register[14][4] ), .B1(n3167), .Y(n5358) );
  OA22XL U4053 ( .A0(\i_MIPS/Register/register[22][3] ), .A1(n3117), .B0(
        \i_MIPS/Register/register[30][3] ), .B1(n3115), .Y(n6564) );
  OA22XL U4054 ( .A0(\i_MIPS/Register/register[6][3] ), .A1(n3117), .B0(
        \i_MIPS/Register/register[14][3] ), .B1(n3113), .Y(n6555) );
  OA22XL U4055 ( .A0(\i_MIPS/Register/register[22][3] ), .A1(n3172), .B0(
        \i_MIPS/Register/register[30][3] ), .B1(n3169), .Y(n6585) );
  OA22XL U4056 ( .A0(\i_MIPS/Register/register[6][3] ), .A1(n3172), .B0(
        \i_MIPS/Register/register[14][3] ), .B1(n3169), .Y(n6576) );
  OA22XL U4057 ( .A0(\i_MIPS/Register/register[22][17] ), .A1(n3171), .B0(
        \i_MIPS/Register/register[30][17] ), .B1(n3168), .Y(n5719) );
  OA22XL U4058 ( .A0(\i_MIPS/Register/register[6][18] ), .A1(n3172), .B0(
        \i_MIPS/Register/register[14][18] ), .B1(n3168), .Y(n5782) );
  OA22XL U4059 ( .A0(\i_MIPS/Register/register[6][17] ), .A1(n3171), .B0(
        \i_MIPS/Register/register[14][17] ), .B1(n3168), .Y(n5710) );
  OA22XL U4060 ( .A0(\i_MIPS/Register/register[22][25] ), .A1(n3171), .B0(
        \i_MIPS/Register/register[30][25] ), .B1(n3167), .Y(n5521) );
  OA22XL U4061 ( .A0(\i_MIPS/Register/register[6][25] ), .A1(n3171), .B0(
        \i_MIPS/Register/register[14][25] ), .B1(n3167), .Y(n5512) );
  OA22XL U4062 ( .A0(\i_MIPS/Register/register[22][25] ), .A1(n3118), .B0(
        \i_MIPS/Register/register[30][25] ), .B1(n3114), .Y(n5498) );
  OA22XL U4063 ( .A0(\i_MIPS/Register/register[6][25] ), .A1(n3116), .B0(
        \i_MIPS/Register/register[14][25] ), .B1(n3114), .Y(n5489) );
  OA22XL U4064 ( .A0(\i_MIPS/Register/register[22][12] ), .A1(n3117), .B0(
        \i_MIPS/Register/register[30][12] ), .B1(n3114), .Y(n6286) );
  OA22XL U4065 ( .A0(\i_MIPS/Register/register[6][12] ), .A1(n3117), .B0(
        \i_MIPS/Register/register[14][12] ), .B1(n3114), .Y(n6277) );
  OA22XL U4066 ( .A0(\i_MIPS/Register/register[22][21] ), .A1(n3117), .B0(
        \i_MIPS/Register/register[30][21] ), .B1(n3113), .Y(n6491) );
  OA22XL U4067 ( .A0(\i_MIPS/Register/register[6][21] ), .A1(n3117), .B0(
        \i_MIPS/Register/register[14][21] ), .B1(n3115), .Y(n6482) );
  OA22XL U4068 ( .A0(\i_MIPS/Register/register[22][26] ), .A1(n3171), .B0(
        \i_MIPS/Register/register[30][26] ), .B1(n3168), .Y(n6108) );
  OA22XL U4069 ( .A0(\i_MIPS/Register/register[6][26] ), .A1(n3171), .B0(
        \i_MIPS/Register/register[14][26] ), .B1(n3168), .Y(n6099) );
  OA22XL U4070 ( .A0(\i_MIPS/Register/register[22][21] ), .A1(n3172), .B0(
        \i_MIPS/Register/register[30][21] ), .B1(n3169), .Y(n6514) );
  OA22XL U4071 ( .A0(\i_MIPS/Register/register[6][21] ), .A1(n3172), .B0(
        \i_MIPS/Register/register[14][21] ), .B1(n3169), .Y(n6505) );
  OA22XL U4072 ( .A0(\i_MIPS/Register/register[22][26] ), .A1(n3116), .B0(
        \i_MIPS/Register/register[30][26] ), .B1(n3115), .Y(n6085) );
  OA22XL U4073 ( .A0(\i_MIPS/Register/register[6][26] ), .A1(n3117), .B0(
        \i_MIPS/Register/register[14][26] ), .B1(n3115), .Y(n6076) );
  OA22XL U4074 ( .A0(\i_MIPS/Register/register[22][19] ), .A1(n3118), .B0(
        \i_MIPS/Register/register[30][19] ), .B1(n3114), .Y(n5636) );
  OA22XL U4075 ( .A0(\i_MIPS/Register/register[6][19] ), .A1(n3117), .B0(
        \i_MIPS/Register/register[14][19] ), .B1(n3114), .Y(n5627) );
  OA22XL U4076 ( .A0(\i_MIPS/Register/register[22][19] ), .A1(n3171), .B0(
        \i_MIPS/Register/register[30][19] ), .B1(n3167), .Y(n5659) );
  OA22XL U4077 ( .A0(\i_MIPS/Register/register[6][19] ), .A1(n3171), .B0(
        \i_MIPS/Register/register[14][19] ), .B1(n3167), .Y(n5650) );
  OA22XL U4078 ( .A0(\i_MIPS/Register/register[22][24] ), .A1(n3118), .B0(
        \i_MIPS/Register/register[30][24] ), .B1(n3115), .Y(n6010) );
  OA22XL U4079 ( .A0(\i_MIPS/Register/register[6][24] ), .A1(n3116), .B0(
        \i_MIPS/Register/register[14][24] ), .B1(n3115), .Y(n6001) );
  OA22XL U4080 ( .A0(\i_MIPS/Register/register[22][20] ), .A1(n3170), .B0(
        \i_MIPS/Register/register[30][20] ), .B1(n3167), .Y(n4855) );
  OA22XL U4081 ( .A0(\i_MIPS/Register/register[6][20] ), .A1(n3170), .B0(
        \i_MIPS/Register/register[14][20] ), .B1(n3168), .Y(n4846) );
  OA22XL U4082 ( .A0(\i_MIPS/Register/register[22][24] ), .A1(n3171), .B0(
        \i_MIPS/Register/register[30][24] ), .B1(n3168), .Y(n6033) );
  OA22XL U4083 ( .A0(\i_MIPS/Register/register[6][24] ), .A1(n2777), .B0(
        \i_MIPS/Register/register[14][24] ), .B1(n3168), .Y(n6024) );
  OA22XL U4084 ( .A0(\i_MIPS/Register/register[6][20] ), .A1(n3116), .B0(
        \i_MIPS/Register/register[14][20] ), .B1(n3113), .Y(n4869) );
  OA22XL U4085 ( .A0(\i_MIPS/Register/register[22][20] ), .A1(n3116), .B0(
        \i_MIPS/Register/register[30][20] ), .B1(n3113), .Y(n4878) );
  OA22XL U4086 ( .A0(\i_MIPS/Register/register[22][29] ), .A1(n3171), .B0(
        \i_MIPS/Register/register[30][29] ), .B1(n3168), .Y(n5871) );
  OA22XL U4087 ( .A0(\i_MIPS/Register/register[6][29] ), .A1(n3172), .B0(
        \i_MIPS/Register/register[14][29] ), .B1(n3168), .Y(n5862) );
  OA22XL U4088 ( .A0(\i_MIPS/Register/register[22][29] ), .A1(n3118), .B0(
        \i_MIPS/Register/register[30][29] ), .B1(n3115), .Y(n5848) );
  OA22XL U4089 ( .A0(\i_MIPS/Register/register[6][29] ), .A1(n3117), .B0(
        \i_MIPS/Register/register[14][29] ), .B1(n3115), .Y(n5839) );
  OA22XL U4090 ( .A0(\i_MIPS/Register/register[22][16] ), .A1(n3118), .B0(
        \i_MIPS/Register/register[30][16] ), .B1(n2782), .Y(n6959) );
  OA22XL U4091 ( .A0(\i_MIPS/Register/register[22][2] ), .A1(n3118), .B0(
        \i_MIPS/Register/register[30][2] ), .B1(n3113), .Y(n6636) );
  OA22XL U4092 ( .A0(\i_MIPS/Register/register[6][2] ), .A1(n3118), .B0(
        \i_MIPS/Register/register[14][2] ), .B1(n3115), .Y(n6627) );
  OA22XL U4093 ( .A0(\i_MIPS/Register/register[22][22] ), .A1(n3170), .B0(
        \i_MIPS/Register/register[30][22] ), .B1(n3167), .Y(n6714) );
  OA22XL U4094 ( .A0(\i_MIPS/Register/register[6][22] ), .A1(n2777), .B0(
        \i_MIPS/Register/register[14][22] ), .B1(n3169), .Y(n6705) );
  OA22XL U4095 ( .A0(\i_MIPS/Register/register[22][22] ), .A1(n3118), .B0(
        \i_MIPS/Register/register[30][22] ), .B1(n3114), .Y(n6735) );
  OA22XL U4096 ( .A0(\i_MIPS/Register/register[6][22] ), .A1(n3118), .B0(
        \i_MIPS/Register/register[14][22] ), .B1(n3115), .Y(n6726) );
  OA22XL U4097 ( .A0(\i_MIPS/Register/register[6][23] ), .A1(n3172), .B0(
        \i_MIPS/Register/register[14][23] ), .B1(n3167), .Y(n6858) );
  OA22XL U4098 ( .A0(\i_MIPS/Register/register[22][27] ), .A1(n3172), .B0(
        \i_MIPS/Register/register[30][27] ), .B1(n3168), .Y(n6811) );
  OA22XL U4099 ( .A0(\i_MIPS/Register/register[6][27] ), .A1(n3170), .B0(
        \i_MIPS/Register/register[14][27] ), .B1(n3167), .Y(n6802) );
  OA22XL U4100 ( .A0(\i_MIPS/Register/register[22][27] ), .A1(n3118), .B0(
        \i_MIPS/Register/register[30][27] ), .B1(n3114), .Y(n6788) );
  OA22XL U4101 ( .A0(\i_MIPS/Register/register[6][27] ), .A1(n3118), .B0(
        \i_MIPS/Register/register[14][27] ), .B1(n3113), .Y(n6779) );
  AO21XL U4102 ( .A0(\i_MIPS/ID_EX[89] ), .A1(n3629), .B0(n2804), .Y(
        \i_MIPS/n496 ) );
  AO21XL U4103 ( .A0(\i_MIPS/ID_EX[90] ), .A1(n3629), .B0(n2804), .Y(
        \i_MIPS/n495 ) );
  AO21XL U4104 ( .A0(\i_MIPS/ID_EX[91] ), .A1(n3629), .B0(n2804), .Y(
        \i_MIPS/n494 ) );
  AO21XL U4105 ( .A0(\i_MIPS/ID_EX[92] ), .A1(n3629), .B0(n2804), .Y(
        \i_MIPS/n493 ) );
  AO21XL U4106 ( .A0(\i_MIPS/ID_EX[93] ), .A1(n3629), .B0(n2804), .Y(
        \i_MIPS/n492 ) );
  AO21XL U4107 ( .A0(\i_MIPS/ID_EX[94] ), .A1(n3629), .B0(n2804), .Y(
        \i_MIPS/n491 ) );
  AO21XL U4108 ( .A0(\i_MIPS/ID_EX[95] ), .A1(n3629), .B0(n2804), .Y(
        \i_MIPS/n490 ) );
  AO21XL U4109 ( .A0(\i_MIPS/ID_EX[96] ), .A1(n3629), .B0(n2804), .Y(
        \i_MIPS/n489 ) );
  AO21XL U4110 ( .A0(\i_MIPS/ID_EX[97] ), .A1(n3629), .B0(n2804), .Y(
        \i_MIPS/n488 ) );
  AO21XL U4111 ( .A0(\i_MIPS/ID_EX[98] ), .A1(n3629), .B0(n2804), .Y(
        \i_MIPS/n487 ) );
  AO21XL U4112 ( .A0(\i_MIPS/ID_EX[99] ), .A1(n3629), .B0(n2804), .Y(
        \i_MIPS/n486 ) );
  AO21XL U4113 ( .A0(\i_MIPS/ID_EX[100] ), .A1(n3629), .B0(n2804), .Y(
        \i_MIPS/n485 ) );
  AO21XL U4114 ( .A0(\i_MIPS/ID_EX[101] ), .A1(n3629), .B0(n2804), .Y(
        \i_MIPS/n484 ) );
  AO21XL U4115 ( .A0(\i_MIPS/ID_EX[102] ), .A1(n3629), .B0(n2804), .Y(
        \i_MIPS/n483 ) );
  AO21XL U4116 ( .A0(\i_MIPS/ID_EX[103] ), .A1(n3629), .B0(n2804), .Y(
        \i_MIPS/n482 ) );
  AND2XL U4117 ( .A(n3079), .B(\i_MIPS/ALU/N303 ), .Y(n2985) );
  MX2XL U4118 ( .A(\i_MIPS/ID_EX[76] ), .B(\i_MIPS/Sign_Extend_ID[3] ), .S0(
        n3623), .Y(\i_MIPS/n509 ) );
  MX2XL U4119 ( .A(n4016), .B(\i_MIPS/Sign_Extend_ID[8] ), .S0(n3623), .Y(
        \i_MIPS/n504 ) );
  MX2XL U4120 ( .A(\i_MIPS/ID_EX[77] ), .B(\i_MIPS/Sign_Extend_ID[4] ), .S0(
        n3624), .Y(\i_MIPS/n508 ) );
  MX2XL U4121 ( .A(\i_MIPS/ID_EX[52] ), .B(n7804), .S0(n3625), .Y(
        \i_MIPS/n415 ) );
  MX2XL U4122 ( .A(\i_MIPS/ID_EX[49] ), .B(n7806), .S0(n3625), .Y(
        \i_MIPS/n421 ) );
  MX2XL U4123 ( .A(n1890), .B(n8011), .S0(n3625), .Y(\i_MIPS/n417 ) );
  MX2XL U4124 ( .A(\i_MIPS/ID_EX[69] ), .B(n8265), .S0(n3625), .Y(
        \i_MIPS/n381 ) );
  MX2XL U4125 ( .A(\i_MIPS/ID_EX[67] ), .B(n8165), .S0(n3625), .Y(
        \i_MIPS/n385 ) );
  MX2XL U4126 ( .A(\i_MIPS/ID_EX[68] ), .B(n8166), .S0(n3625), .Y(
        \i_MIPS/n383 ) );
  MX2XL U4127 ( .A(\i_MIPS/EX_MEM[5] ), .B(n8257), .S0(n3625), .Y(
        \i_MIPS/n469 ) );
  MX2XL U4128 ( .A(n1889), .B(n7785), .S0(n3626), .Y(\i_MIPS/n411 ) );
  MX2XL U4129 ( .A(n1884), .B(n7782), .S0(n3626), .Y(\i_MIPS/n427 ) );
  MX2XL U4130 ( .A(n1892), .B(n2883), .S0(n3626), .Y(\i_MIPS/n530 ) );
  MX2XL U4131 ( .A(n3075), .B(\i_MIPS/Sign_Extend_ID[6] ), .S0(n3626), .Y(
        \i_MIPS/n506 ) );
  MX2XL U4132 ( .A(\i_MIPS/Reg_W[0] ), .B(\i_MIPS/EX_MEM_next[69] ), .S0(n3622), .Y(\i_MIPS/n477 ) );
  MX2XL U4133 ( .A(\i_MIPS/Reg_W[1] ), .B(\i_MIPS/EX_MEM_next[70] ), .S0(n3622), .Y(\i_MIPS/n476 ) );
  MX2XL U4134 ( .A(\i_MIPS/Reg_W[2] ), .B(\i_MIPS/EX_MEM_next[71] ), .S0(n3623), .Y(\i_MIPS/n475 ) );
  MX2XL U4135 ( .A(\i_MIPS/Reg_W[3] ), .B(n2890), .S0(n3623), .Y(\i_MIPS/n474 ) );
  MX2XL U4136 ( .A(\i_MIPS/Reg_W[4] ), .B(n2891), .S0(n3623), .Y(\i_MIPS/n473 ) );
  MX2XL U4137 ( .A(\i_MIPS/ID_EX[75] ), .B(\i_MIPS/Sign_Extend_ID[2] ), .S0(
        n3623), .Y(\i_MIPS/n510 ) );
  MX2XL U4138 ( .A(\i_MIPS/ID_EX[74] ), .B(\i_MIPS/Sign_Extend_ID[1] ), .S0(
        n3622), .Y(\i_MIPS/n511 ) );
  MX2XL U4139 ( .A(\I_cache/cache[7][128] ), .B(n8448), .S0(n3496), .Y(n9133)
         );
  MX2XL U4140 ( .A(\I_cache/cache[7][152] ), .B(n8449), .S0(n3496), .Y(n8941)
         );
  MX2XL U4141 ( .A(\I_cache/cache[6][152] ), .B(n8449), .S0(n3540), .Y(n8942)
         );
  MX2XL U4142 ( .A(\I_cache/cache[5][152] ), .B(n8449), .S0(n3405), .Y(n8943)
         );
  MX2XL U4143 ( .A(\I_cache/cache[4][152] ), .B(n8449), .S0(n3451), .Y(n8944)
         );
  MX2XL U4144 ( .A(\I_cache/cache[3][152] ), .B(n8449), .S0(n3318), .Y(n8945)
         );
  MX2XL U4145 ( .A(\I_cache/cache[2][152] ), .B(n8449), .S0(n3361), .Y(n8946)
         );
  MX2XL U4146 ( .A(\I_cache/cache[1][152] ), .B(n8449), .S0(n3228), .Y(n8947)
         );
  MX2XL U4147 ( .A(\I_cache/cache[0][152] ), .B(n8449), .S0(n3273), .Y(n8948)
         );
  MX2XL U4148 ( .A(\I_cache/cache[7][151] ), .B(n8447), .S0(n3496), .Y(n8949)
         );
  MX2XL U4149 ( .A(\I_cache/cache[6][151] ), .B(n8447), .S0(n3540), .Y(n8950)
         );
  MX2XL U4150 ( .A(\I_cache/cache[5][151] ), .B(n8447), .S0(n3405), .Y(n8951)
         );
  MX2XL U4151 ( .A(\I_cache/cache[4][151] ), .B(n8447), .S0(n3451), .Y(n8952)
         );
  MX2XL U4152 ( .A(\I_cache/cache[3][151] ), .B(n8447), .S0(n3318), .Y(n8953)
         );
  MX2XL U4153 ( .A(\I_cache/cache[2][151] ), .B(n8447), .S0(n3361), .Y(n8954)
         );
  MX2XL U4154 ( .A(\I_cache/cache[1][151] ), .B(n8447), .S0(n3228), .Y(n8955)
         );
  MX2XL U4155 ( .A(\I_cache/cache[0][151] ), .B(n8447), .S0(n3273), .Y(n8956)
         );
  MX2XL U4156 ( .A(\I_cache/cache[7][150] ), .B(n8435), .S0(n3495), .Y(n8957)
         );
  MX2XL U4157 ( .A(\I_cache/cache[6][150] ), .B(n8435), .S0(n3535), .Y(n8958)
         );
  MX2XL U4158 ( .A(\I_cache/cache[5][150] ), .B(n8435), .S0(n3407), .Y(n8959)
         );
  MX2XL U4159 ( .A(\I_cache/cache[4][150] ), .B(n8435), .S0(n3450), .Y(n8960)
         );
  MX2XL U4160 ( .A(\I_cache/cache[3][150] ), .B(n8435), .S0(n3317), .Y(n8961)
         );
  MX2XL U4161 ( .A(\I_cache/cache[2][150] ), .B(n8435), .S0(n3360), .Y(n8962)
         );
  MX2XL U4162 ( .A(\I_cache/cache[1][150] ), .B(n8435), .S0(n3227), .Y(n8963)
         );
  MX2XL U4163 ( .A(\I_cache/cache[0][150] ), .B(n8435), .S0(n3270), .Y(n8964)
         );
  MX2XL U4164 ( .A(\I_cache/cache[7][149] ), .B(n8441), .S0(n3496), .Y(n8965)
         );
  MX2XL U4165 ( .A(\I_cache/cache[6][149] ), .B(n8441), .S0(n3540), .Y(n8966)
         );
  MX2XL U4166 ( .A(\I_cache/cache[5][149] ), .B(n8441), .S0(n3405), .Y(n8967)
         );
  MX2XL U4167 ( .A(\I_cache/cache[4][149] ), .B(n8441), .S0(n3451), .Y(n8968)
         );
  MX2XL U4168 ( .A(\I_cache/cache[3][149] ), .B(n8441), .S0(n3318), .Y(n8969)
         );
  MX2XL U4169 ( .A(\I_cache/cache[2][149] ), .B(n8441), .S0(n3361), .Y(n8970)
         );
  MX2XL U4170 ( .A(\I_cache/cache[1][149] ), .B(n8441), .S0(n3228), .Y(n8971)
         );
  MX2XL U4171 ( .A(\I_cache/cache[0][149] ), .B(n8441), .S0(n3273), .Y(n8972)
         );
  MX2XL U4172 ( .A(\I_cache/cache[7][148] ), .B(n8443), .S0(n3496), .Y(n8973)
         );
  MX2XL U4173 ( .A(\I_cache/cache[6][148] ), .B(n8443), .S0(n3540), .Y(n8974)
         );
  MX2XL U4174 ( .A(\I_cache/cache[5][148] ), .B(n8443), .S0(n3405), .Y(n8975)
         );
  MX2XL U4175 ( .A(\I_cache/cache[4][148] ), .B(n8443), .S0(n3451), .Y(n8976)
         );
  MX2XL U4176 ( .A(\I_cache/cache[3][148] ), .B(n8443), .S0(n3318), .Y(n8977)
         );
  MX2XL U4177 ( .A(\I_cache/cache[2][148] ), .B(n8443), .S0(n3361), .Y(n8978)
         );
  MX2XL U4178 ( .A(\I_cache/cache[1][148] ), .B(n8443), .S0(n3228), .Y(n8979)
         );
  MX2XL U4179 ( .A(\I_cache/cache[0][148] ), .B(n8443), .S0(n3273), .Y(n8980)
         );
  MX2XL U4180 ( .A(\I_cache/cache[7][147] ), .B(n8442), .S0(n3496), .Y(n8981)
         );
  MX2XL U4181 ( .A(\I_cache/cache[6][147] ), .B(n8442), .S0(n3540), .Y(n8982)
         );
  MX2XL U4182 ( .A(\I_cache/cache[5][147] ), .B(n8442), .S0(n3405), .Y(n8983)
         );
  MX2XL U4183 ( .A(\I_cache/cache[4][147] ), .B(n8442), .S0(n3451), .Y(n8984)
         );
  MX2XL U4184 ( .A(\I_cache/cache[3][147] ), .B(n8442), .S0(n3318), .Y(n8985)
         );
  MX2XL U4185 ( .A(\I_cache/cache[2][147] ), .B(n8442), .S0(n3361), .Y(n8986)
         );
  MX2XL U4186 ( .A(\I_cache/cache[1][147] ), .B(n8442), .S0(n3228), .Y(n8987)
         );
  MX2XL U4187 ( .A(\I_cache/cache[0][147] ), .B(n8442), .S0(n3273), .Y(n8988)
         );
  MX2XL U4188 ( .A(\I_cache/cache[7][146] ), .B(n8434), .S0(n3495), .Y(n8989)
         );
  MX2XL U4189 ( .A(\I_cache/cache[6][146] ), .B(n8434), .S0(n3535), .Y(n8990)
         );
  MX2XL U4190 ( .A(\I_cache/cache[5][146] ), .B(n8434), .S0(n3405), .Y(n8991)
         );
  MX2XL U4191 ( .A(\I_cache/cache[4][146] ), .B(n8434), .S0(n3450), .Y(n8992)
         );
  MX2XL U4192 ( .A(\I_cache/cache[3][146] ), .B(n8434), .S0(n3317), .Y(n8993)
         );
  MX2XL U4193 ( .A(\I_cache/cache[2][146] ), .B(n8434), .S0(n3360), .Y(n8994)
         );
  MX2XL U4194 ( .A(\I_cache/cache[1][146] ), .B(n8434), .S0(n3227), .Y(n8995)
         );
  MX2XL U4195 ( .A(\I_cache/cache[0][146] ), .B(n8434), .S0(n3269), .Y(n8996)
         );
  MX2XL U4196 ( .A(\I_cache/cache[7][145] ), .B(n8436), .S0(n3495), .Y(n8997)
         );
  MX2XL U4197 ( .A(\I_cache/cache[6][145] ), .B(n8436), .S0(n3532), .Y(n8998)
         );
  MX2XL U4198 ( .A(\I_cache/cache[5][145] ), .B(n8436), .S0(n3398), .Y(n8999)
         );
  MX2XL U4199 ( .A(\I_cache/cache[4][145] ), .B(n8436), .S0(n3450), .Y(n9000)
         );
  MX2XL U4200 ( .A(\I_cache/cache[3][145] ), .B(n8436), .S0(n3317), .Y(n9001)
         );
  MX2XL U4201 ( .A(\I_cache/cache[2][145] ), .B(n8436), .S0(n3360), .Y(n9002)
         );
  MX2XL U4202 ( .A(\I_cache/cache[1][145] ), .B(n8436), .S0(n3227), .Y(n9003)
         );
  MX2XL U4203 ( .A(\I_cache/cache[0][145] ), .B(n8436), .S0(n3271), .Y(n9004)
         );
  MX2XL U4204 ( .A(\I_cache/cache[7][144] ), .B(n8451), .S0(n3496), .Y(n9005)
         );
  MX2XL U4205 ( .A(\I_cache/cache[6][144] ), .B(n8451), .S0(n3540), .Y(n9006)
         );
  MX2XL U4206 ( .A(\I_cache/cache[5][144] ), .B(n8451), .S0(n3405), .Y(n9007)
         );
  MX2XL U4207 ( .A(\I_cache/cache[4][144] ), .B(n8451), .S0(n3451), .Y(n9008)
         );
  MX2XL U4208 ( .A(\I_cache/cache[3][144] ), .B(n8451), .S0(n3318), .Y(n9009)
         );
  MX2XL U4209 ( .A(\I_cache/cache[2][144] ), .B(n8451), .S0(n3361), .Y(n9010)
         );
  MX2XL U4210 ( .A(\I_cache/cache[1][144] ), .B(n8451), .S0(n3228), .Y(n9011)
         );
  MX2XL U4211 ( .A(\I_cache/cache[0][144] ), .B(n8451), .S0(n3273), .Y(n9012)
         );
  MX2XL U4212 ( .A(\I_cache/cache[7][143] ), .B(n8430), .S0(n3495), .Y(n9013)
         );
  MX2XL U4213 ( .A(\I_cache/cache[6][143] ), .B(n8430), .S0(n3533), .Y(n9014)
         );
  MX2XL U4214 ( .A(\I_cache/cache[5][143] ), .B(n8430), .S0(n3399), .Y(n9015)
         );
  MX2XL U4215 ( .A(\I_cache/cache[4][143] ), .B(n8430), .S0(n3450), .Y(n9016)
         );
  MX2XL U4216 ( .A(\I_cache/cache[3][143] ), .B(n8430), .S0(n3317), .Y(n9017)
         );
  MX2XL U4217 ( .A(\I_cache/cache[2][143] ), .B(n8430), .S0(n3360), .Y(n9018)
         );
  MX2XL U4218 ( .A(\I_cache/cache[1][143] ), .B(n8430), .S0(n3227), .Y(n9019)
         );
  MX2XL U4219 ( .A(\I_cache/cache[0][143] ), .B(n8430), .S0(n3270), .Y(n9020)
         );
  MX2XL U4220 ( .A(\I_cache/cache[7][142] ), .B(n8428), .S0(n3495), .Y(n9021)
         );
  MX2XL U4221 ( .A(\I_cache/cache[6][142] ), .B(n8428), .S0(n3534), .Y(n9022)
         );
  MX2XL U4222 ( .A(\I_cache/cache[5][142] ), .B(n8428), .S0(n3407), .Y(n9023)
         );
  MX2XL U4223 ( .A(\I_cache/cache[4][142] ), .B(n8428), .S0(n3450), .Y(n9024)
         );
  MX2XL U4224 ( .A(\I_cache/cache[3][142] ), .B(n8428), .S0(n3317), .Y(n9025)
         );
  MX2XL U4225 ( .A(\I_cache/cache[2][142] ), .B(n8428), .S0(n3360), .Y(n9026)
         );
  MX2XL U4226 ( .A(\I_cache/cache[1][142] ), .B(n8428), .S0(n3227), .Y(n9027)
         );
  MX2XL U4227 ( .A(\I_cache/cache[0][142] ), .B(n8428), .S0(n3269), .Y(n9028)
         );
  MX2XL U4228 ( .A(\I_cache/cache[7][141] ), .B(n8429), .S0(n3495), .Y(n9029)
         );
  MX2XL U4229 ( .A(\I_cache/cache[6][141] ), .B(n8429), .S0(n3536), .Y(n9030)
         );
  MX2XL U4230 ( .A(\I_cache/cache[5][141] ), .B(n8429), .S0(n3403), .Y(n9031)
         );
  MX2XL U4231 ( .A(\I_cache/cache[4][141] ), .B(n8429), .S0(n3450), .Y(n9032)
         );
  MX2XL U4232 ( .A(\I_cache/cache[3][141] ), .B(n8429), .S0(n3317), .Y(n9033)
         );
  MX2XL U4233 ( .A(\I_cache/cache[2][141] ), .B(n8429), .S0(n3360), .Y(n9034)
         );
  MX2XL U4234 ( .A(\I_cache/cache[1][141] ), .B(n8429), .S0(n3227), .Y(n9035)
         );
  MX2XL U4235 ( .A(\I_cache/cache[0][141] ), .B(n8429), .S0(n3271), .Y(n9036)
         );
  MX2XL U4236 ( .A(\I_cache/cache[7][140] ), .B(n8454), .S0(n3495), .Y(n9037)
         );
  MX2XL U4237 ( .A(\I_cache/cache[6][140] ), .B(n8454), .S0(n3535), .Y(n9038)
         );
  MX2XL U4238 ( .A(\I_cache/cache[5][140] ), .B(n8454), .S0(n3402), .Y(n9039)
         );
  MX2XL U4239 ( .A(\I_cache/cache[4][140] ), .B(n8454), .S0(n3450), .Y(n9040)
         );
  MX2XL U4240 ( .A(\I_cache/cache[3][140] ), .B(n8454), .S0(n3317), .Y(n9041)
         );
  MX2XL U4241 ( .A(\I_cache/cache[2][140] ), .B(n8454), .S0(n3360), .Y(n9042)
         );
  MX2XL U4242 ( .A(\I_cache/cache[1][140] ), .B(n8454), .S0(n3227), .Y(n9043)
         );
  MX2XL U4243 ( .A(\I_cache/cache[0][140] ), .B(n8454), .S0(n3270), .Y(n9044)
         );
  MX2XL U4244 ( .A(\I_cache/cache[7][139] ), .B(n8450), .S0(n3496), .Y(n9045)
         );
  MX2XL U4245 ( .A(\I_cache/cache[6][139] ), .B(n8450), .S0(n3540), .Y(n9046)
         );
  MX2XL U4246 ( .A(\I_cache/cache[5][139] ), .B(n8450), .S0(n3405), .Y(n9047)
         );
  MX2XL U4247 ( .A(\I_cache/cache[4][139] ), .B(n8450), .S0(n3451), .Y(n9048)
         );
  MX2XL U4248 ( .A(\I_cache/cache[3][139] ), .B(n8450), .S0(n3318), .Y(n9049)
         );
  MX2XL U4249 ( .A(\I_cache/cache[2][139] ), .B(n8450), .S0(n3361), .Y(n9050)
         );
  MX2XL U4250 ( .A(\I_cache/cache[1][139] ), .B(n8450), .S0(n3228), .Y(n9051)
         );
  MX2XL U4251 ( .A(\I_cache/cache[0][139] ), .B(n8450), .S0(n3273), .Y(n9052)
         );
  MX2XL U4252 ( .A(\I_cache/cache[7][138] ), .B(n8437), .S0(n3495), .Y(n9053)
         );
  MX2XL U4253 ( .A(\I_cache/cache[6][138] ), .B(n8437), .S0(n3541), .Y(n9054)
         );
  MX2XL U4254 ( .A(\I_cache/cache[5][138] ), .B(n8437), .S0(n3404), .Y(n9055)
         );
  MX2XL U4255 ( .A(\I_cache/cache[4][138] ), .B(n8437), .S0(n3450), .Y(n9056)
         );
  MX2XL U4256 ( .A(\I_cache/cache[3][138] ), .B(n8437), .S0(n3317), .Y(n9057)
         );
  MX2XL U4257 ( .A(\I_cache/cache[2][138] ), .B(n8437), .S0(n3360), .Y(n9058)
         );
  MX2XL U4258 ( .A(\I_cache/cache[1][138] ), .B(n8437), .S0(n3227), .Y(n9059)
         );
  MX2XL U4259 ( .A(\I_cache/cache[0][138] ), .B(n8437), .S0(n3269), .Y(n9060)
         );
  MX2XL U4260 ( .A(\I_cache/cache[7][137] ), .B(n8444), .S0(n3496), .Y(n9061)
         );
  MX2XL U4261 ( .A(\I_cache/cache[6][137] ), .B(n8444), .S0(n3540), .Y(n9062)
         );
  MX2XL U4262 ( .A(\I_cache/cache[5][137] ), .B(n8444), .S0(n3405), .Y(n9063)
         );
  MX2XL U4263 ( .A(\I_cache/cache[4][137] ), .B(n8444), .S0(n3451), .Y(n9064)
         );
  MX2XL U4264 ( .A(\I_cache/cache[3][137] ), .B(n8444), .S0(n3318), .Y(n9065)
         );
  MX2XL U4265 ( .A(\I_cache/cache[2][137] ), .B(n8444), .S0(n3361), .Y(n9066)
         );
  MX2XL U4266 ( .A(\I_cache/cache[1][137] ), .B(n8444), .S0(n3228), .Y(n9067)
         );
  MX2XL U4267 ( .A(\I_cache/cache[0][137] ), .B(n8444), .S0(n3273), .Y(n9068)
         );
  MX2XL U4268 ( .A(\I_cache/cache[7][136] ), .B(n8446), .S0(n3496), .Y(n9069)
         );
  MX2XL U4269 ( .A(\I_cache/cache[6][136] ), .B(n8446), .S0(n3540), .Y(n9070)
         );
  MX2XL U4270 ( .A(\I_cache/cache[5][136] ), .B(n8446), .S0(n3405), .Y(n9071)
         );
  MX2XL U4271 ( .A(\I_cache/cache[4][136] ), .B(n8446), .S0(n3451), .Y(n9072)
         );
  MX2XL U4272 ( .A(\I_cache/cache[3][136] ), .B(n8446), .S0(n3318), .Y(n9073)
         );
  MX2XL U4273 ( .A(\I_cache/cache[2][136] ), .B(n8446), .S0(n3361), .Y(n9074)
         );
  MX2XL U4274 ( .A(\I_cache/cache[1][136] ), .B(n8446), .S0(n3228), .Y(n9075)
         );
  MX2XL U4275 ( .A(\I_cache/cache[0][136] ), .B(n8446), .S0(n3273), .Y(n9076)
         );
  MX2XL U4276 ( .A(\I_cache/cache[7][135] ), .B(n8445), .S0(n3496), .Y(n9077)
         );
  MX2XL U4277 ( .A(\I_cache/cache[6][135] ), .B(n8445), .S0(n3540), .Y(n9078)
         );
  MX2XL U4278 ( .A(\I_cache/cache[5][135] ), .B(n8445), .S0(n3405), .Y(n9079)
         );
  MX2XL U4279 ( .A(\I_cache/cache[4][135] ), .B(n8445), .S0(n3451), .Y(n9080)
         );
  MX2XL U4280 ( .A(\I_cache/cache[3][135] ), .B(n8445), .S0(n3318), .Y(n9081)
         );
  MX2XL U4281 ( .A(\I_cache/cache[2][135] ), .B(n8445), .S0(n3361), .Y(n9082)
         );
  MX2XL U4282 ( .A(\I_cache/cache[1][135] ), .B(n8445), .S0(n3228), .Y(n9083)
         );
  MX2XL U4283 ( .A(\I_cache/cache[0][135] ), .B(n8445), .S0(n3273), .Y(n9084)
         );
  MX2XL U4284 ( .A(\I_cache/cache[7][134] ), .B(n8439), .S0(n3494), .Y(n9085)
         );
  MX2XL U4285 ( .A(\I_cache/cache[6][134] ), .B(n8439), .S0(n3539), .Y(n9086)
         );
  MX2XL U4286 ( .A(\I_cache/cache[5][134] ), .B(n8439), .S0(n3404), .Y(n9087)
         );
  MX2XL U4287 ( .A(\I_cache/cache[4][134] ), .B(n8439), .S0(n3449), .Y(n9088)
         );
  MX2XL U4288 ( .A(\I_cache/cache[3][134] ), .B(n8439), .S0(n3316), .Y(n9089)
         );
  MX2XL U4289 ( .A(\I_cache/cache[2][134] ), .B(n8439), .S0(n3359), .Y(n9090)
         );
  MX2XL U4290 ( .A(\I_cache/cache[1][134] ), .B(n8439), .S0(n3226), .Y(n9091)
         );
  MX2XL U4291 ( .A(\I_cache/cache[0][134] ), .B(n8439), .S0(n3272), .Y(n9092)
         );
  MX2XL U4292 ( .A(\I_cache/cache[7][133] ), .B(n8438), .S0(n3495), .Y(n9093)
         );
  MX2XL U4293 ( .A(\I_cache/cache[6][133] ), .B(n8438), .S0(n3532), .Y(n9094)
         );
  MX2XL U4294 ( .A(\I_cache/cache[5][133] ), .B(n8438), .S0(n3401), .Y(n9095)
         );
  MX2XL U4295 ( .A(\I_cache/cache[4][133] ), .B(n8438), .S0(n3450), .Y(n9096)
         );
  MX2XL U4296 ( .A(\I_cache/cache[3][133] ), .B(n8438), .S0(n3317), .Y(n9097)
         );
  MX2XL U4297 ( .A(\I_cache/cache[2][133] ), .B(n8438), .S0(n3360), .Y(n9098)
         );
  MX2XL U4298 ( .A(\I_cache/cache[1][133] ), .B(n8438), .S0(n3227), .Y(n9099)
         );
  MX2XL U4299 ( .A(\I_cache/cache[0][133] ), .B(n8438), .S0(n3271), .Y(n9100)
         );
  MX2XL U4300 ( .A(\I_cache/cache[7][132] ), .B(n8440), .S0(n3496), .Y(n9101)
         );
  MX2XL U4301 ( .A(\I_cache/cache[6][132] ), .B(n8440), .S0(n3540), .Y(n9102)
         );
  MX2XL U4302 ( .A(\I_cache/cache[5][132] ), .B(n8440), .S0(n3405), .Y(n9103)
         );
  MX2XL U4303 ( .A(\I_cache/cache[4][132] ), .B(n8440), .S0(n3451), .Y(n9104)
         );
  MX2XL U4304 ( .A(\I_cache/cache[3][132] ), .B(n8440), .S0(n3318), .Y(n9105)
         );
  MX2XL U4305 ( .A(\I_cache/cache[2][132] ), .B(n8440), .S0(n3361), .Y(n9106)
         );
  MX2XL U4306 ( .A(\I_cache/cache[1][132] ), .B(n8440), .S0(n3228), .Y(n9107)
         );
  MX2XL U4307 ( .A(\I_cache/cache[0][132] ), .B(n8440), .S0(n3273), .Y(n9108)
         );
  MX2XL U4308 ( .A(\I_cache/cache[7][131] ), .B(n8432), .S0(n3495), .Y(n9109)
         );
  MX2XL U4309 ( .A(\I_cache/cache[6][131] ), .B(n8432), .S0(n3533), .Y(n9110)
         );
  MX2XL U4310 ( .A(\I_cache/cache[5][131] ), .B(n8432), .S0(n3405), .Y(n9111)
         );
  MX2XL U4311 ( .A(\I_cache/cache[4][131] ), .B(n8432), .S0(n3450), .Y(n9112)
         );
  MX2XL U4312 ( .A(\I_cache/cache[3][131] ), .B(n8432), .S0(n3317), .Y(n9113)
         );
  MX2XL U4313 ( .A(\I_cache/cache[2][131] ), .B(n8432), .S0(n3360), .Y(n9114)
         );
  MX2XL U4314 ( .A(\I_cache/cache[1][131] ), .B(n8432), .S0(n3227), .Y(n9115)
         );
  MX2XL U4315 ( .A(\I_cache/cache[0][131] ), .B(n8432), .S0(n3272), .Y(n9116)
         );
  MX2XL U4316 ( .A(\I_cache/cache[7][130] ), .B(n8433), .S0(n3495), .Y(n9117)
         );
  MX2XL U4317 ( .A(\I_cache/cache[6][130] ), .B(n8433), .S0(n3536), .Y(n9118)
         );
  MX2XL U4318 ( .A(\I_cache/cache[5][130] ), .B(n8433), .S0(n3401), .Y(n9119)
         );
  MX2XL U4319 ( .A(\I_cache/cache[4][130] ), .B(n8433), .S0(n3446), .Y(n9120)
         );
  MX2XL U4320 ( .A(\I_cache/cache[3][130] ), .B(n8433), .S0(n3317), .Y(n9121)
         );
  MX2XL U4321 ( .A(\I_cache/cache[2][130] ), .B(n8433), .S0(n3360), .Y(n9122)
         );
  MX2XL U4322 ( .A(\I_cache/cache[1][130] ), .B(n8433), .S0(n3226), .Y(n9123)
         );
  MX2XL U4323 ( .A(\I_cache/cache[0][130] ), .B(n8433), .S0(n3270), .Y(n9124)
         );
  MX2XL U4324 ( .A(\I_cache/cache[7][129] ), .B(n8431), .S0(n3495), .Y(n9125)
         );
  MX2XL U4325 ( .A(\I_cache/cache[6][129] ), .B(n8431), .S0(n3534), .Y(n9126)
         );
  MX2XL U4326 ( .A(\I_cache/cache[5][129] ), .B(n8431), .S0(n3398), .Y(n9127)
         );
  MX2XL U4327 ( .A(\I_cache/cache[4][129] ), .B(n8431), .S0(n3450), .Y(n9128)
         );
  MX2XL U4328 ( .A(\I_cache/cache[3][129] ), .B(n8431), .S0(n3317), .Y(n9129)
         );
  MX2XL U4329 ( .A(\I_cache/cache[2][129] ), .B(n8431), .S0(n3360), .Y(n9130)
         );
  MX2XL U4330 ( .A(\I_cache/cache[1][129] ), .B(n8431), .S0(n3227), .Y(n9131)
         );
  MX2XL U4331 ( .A(\I_cache/cache[0][129] ), .B(n8431), .S0(n3269), .Y(n9132)
         );
  MX2XL U4332 ( .A(\I_cache/cache[6][128] ), .B(n8448), .S0(n3540), .Y(n9134)
         );
  MX2XL U4333 ( .A(\I_cache/cache[5][128] ), .B(n8448), .S0(n3405), .Y(n9135)
         );
  MX2XL U4334 ( .A(\I_cache/cache[4][128] ), .B(n8448), .S0(n3451), .Y(n9136)
         );
  MX2XL U4335 ( .A(\I_cache/cache[3][128] ), .B(n8448), .S0(n3318), .Y(n9137)
         );
  MX2XL U4336 ( .A(\I_cache/cache[2][128] ), .B(n8448), .S0(n3361), .Y(n9138)
         );
  MX2XL U4337 ( .A(\I_cache/cache[1][128] ), .B(n8448), .S0(n3228), .Y(n9139)
         );
  MX2XL U4338 ( .A(\I_cache/cache[0][128] ), .B(n8448), .S0(n3273), .Y(n9140)
         );
  MX2XL U4339 ( .A(\i_MIPS/ID_EX[70] ), .B(n8283), .S0(n3623), .Y(
        \i_MIPS/n379 ) );
  MX2XL U4340 ( .A(\i_MIPS/ID_EX[71] ), .B(n2), .S0(n3623), .Y(\i_MIPS/n377 )
         );
  MX2XL U4341 ( .A(\i_MIPS/ID_EX[65] ), .B(n8037), .S0(n3623), .Y(
        \i_MIPS/n389 ) );
  MX2XL U4342 ( .A(n1887), .B(n7733), .S0(n3623), .Y(\i_MIPS/n435 ) );
  MX2XL U4343 ( .A(\i_MIPS/ID_EX[73] ), .B(\i_MIPS/Sign_Extend_ID[0] ), .S0(
        n3623), .Y(\i_MIPS/n512 ) );
  MX2XL U4344 ( .A(\i_MIPS/ID_EX[60] ), .B(n8014), .S0(n3624), .Y(
        \i_MIPS/n399 ) );
  MX2XL U4345 ( .A(\i_MIPS/ID_EX[78] ), .B(\i_MIPS/Sign_Extend_ID[5] ), .S0(
        n3624), .Y(\i_MIPS/n507 ) );
  MX2XL U4346 ( .A(\i_MIPS/EX_MEM[6] ), .B(n8235), .S0(n3624), .Y(
        \i_MIPS/n468 ) );
  MX2XL U4347 ( .A(n7802), .B(n7801), .S0(n3627), .Y(\i_MIPS/n425 ) );
  MX2XL U4348 ( .A(\I_cache/cache[7][96] ), .B(n8397), .S0(n3495), .Y(n9389)
         );
  MX2XL U4349 ( .A(\I_cache/cache[6][96] ), .B(n8397), .S0(n3532), .Y(n9390)
         );
  MX2XL U4350 ( .A(\I_cache/cache[5][96] ), .B(n8397), .S0(n3407), .Y(n9391)
         );
  MX2XL U4351 ( .A(\I_cache/cache[4][96] ), .B(n8397), .S0(n3451), .Y(n9392)
         );
  MX2XL U4352 ( .A(\I_cache/cache[3][96] ), .B(n8397), .S0(n3317), .Y(n9393)
         );
  MX2XL U4353 ( .A(\I_cache/cache[2][96] ), .B(n8397), .S0(n3360), .Y(n9394)
         );
  MX2XL U4354 ( .A(\I_cache/cache[1][96] ), .B(n8397), .S0(n3227), .Y(n9395)
         );
  MX2X1 U4355 ( .A(\I_cache/cache[0][96] ), .B(n8397), .S0(n3272), .Y(n9396)
         );
  MX2XL U4356 ( .A(\I_cache/cache[7][64] ), .B(n8398), .S0(n3492), .Y(n9645)
         );
  MX2XL U4357 ( .A(\I_cache/cache[6][64] ), .B(n8398), .S0(n3533), .Y(n9646)
         );
  MX2XL U4358 ( .A(\I_cache/cache[5][64] ), .B(n8398), .S0(n3407), .Y(n9647)
         );
  MX2XL U4359 ( .A(\I_cache/cache[4][64] ), .B(n8398), .S0(n3450), .Y(n9648)
         );
  MX2XL U4360 ( .A(\I_cache/cache[3][64] ), .B(n8398), .S0(n3317), .Y(n9649)
         );
  MX2XL U4361 ( .A(\I_cache/cache[2][64] ), .B(n8398), .S0(n3360), .Y(n9650)
         );
  MX2XL U4362 ( .A(\I_cache/cache[1][64] ), .B(n8398), .S0(n3227), .Y(n9651)
         );
  MX2X1 U4363 ( .A(\I_cache/cache[0][64] ), .B(n8398), .S0(n3272), .Y(n9652)
         );
  MX2XL U4364 ( .A(\I_cache/cache[7][32] ), .B(n8396), .S0(n3493), .Y(n9901)
         );
  MX2XL U4365 ( .A(\I_cache/cache[6][32] ), .B(n8396), .S0(n3534), .Y(n9902)
         );
  MX2XL U4366 ( .A(\I_cache/cache[5][32] ), .B(n8396), .S0(n3407), .Y(n9903)
         );
  MX2XL U4367 ( .A(\I_cache/cache[4][32] ), .B(n8396), .S0(n3451), .Y(n9904)
         );
  MX2XL U4368 ( .A(\I_cache/cache[3][32] ), .B(n8396), .S0(n3314), .Y(n9905)
         );
  MX2XL U4369 ( .A(\I_cache/cache[2][32] ), .B(n8396), .S0(n3357), .Y(n9906)
         );
  MX2XL U4370 ( .A(\I_cache/cache[1][32] ), .B(n8396), .S0(n3224), .Y(n9907)
         );
  MX2X1 U4371 ( .A(\I_cache/cache[0][32] ), .B(n8396), .S0(n3271), .Y(n9908)
         );
  MX2XL U4372 ( .A(\I_cache/cache[7][0] ), .B(n8395), .S0(n3495), .Y(n10164)
         );
  MX2XL U4373 ( .A(\I_cache/cache[6][0] ), .B(n8395), .S0(n3535), .Y(n10157)
         );
  MX2XL U4374 ( .A(\I_cache/cache[5][0] ), .B(n8395), .S0(n3407), .Y(n10158)
         );
  MX2XL U4375 ( .A(\I_cache/cache[4][0] ), .B(n8395), .S0(n3449), .Y(n10159)
         );
  MX2XL U4376 ( .A(\I_cache/cache[3][0] ), .B(n8395), .S0(n3315), .Y(n10160)
         );
  MX2X1 U4377 ( .A(\I_cache/cache[2][0] ), .B(n8395), .S0(n3358), .Y(n10161)
         );
  MX2XL U4378 ( .A(\I_cache/cache[1][0] ), .B(n8395), .S0(n3225), .Y(n10162)
         );
  MX2X1 U4379 ( .A(\I_cache/cache[0][0] ), .B(n8395), .S0(n3272), .Y(n10163)
         );
  MX2XL U4380 ( .A(n10297), .B(n8314), .S0(n3627), .Y(\i_MIPS/n438 ) );
  MX2XL U4381 ( .A(\i_MIPS/ID_EX[64] ), .B(n2441), .S0(n3627), .Y(
        \i_MIPS/n391 ) );
  MX2XL U4382 ( .A(\i_MIPS/ID_EX[63] ), .B(n7800), .S0(n3627), .Y(
        \i_MIPS/n393 ) );
  MX2XL U4383 ( .A(\i_MIPS/ID_EX[61] ), .B(n7803), .S0(n3627), .Y(
        \i_MIPS/n397 ) );
  MX2XL U4384 ( .A(n1885), .B(n25), .S0(n3627), .Y(\i_MIPS/n375 ) );
  OA22XL U4385 ( .A0(n3556), .A1(n1880), .B0(n3514), .B1(n946), .Y(n7415) );
  OA22XL U4386 ( .A0(n3556), .A1(n894), .B0(n3514), .B1(n1827), .Y(n7425) );
  OA22XL U4387 ( .A0(n3556), .A1(n895), .B0(n3514), .B1(n1828), .Y(n7430) );
  OA22XL U4388 ( .A0(n3556), .A1(n896), .B0(n3514), .B1(n1829), .Y(n7420) );
  OA22XL U4389 ( .A0(n3557), .A1(n897), .B0(n3515), .B1(n1830), .Y(n7497) );
  OA22XL U4390 ( .A0(n3557), .A1(n898), .B0(n3515), .B1(n1831), .Y(n7487) );
  OA22XL U4391 ( .A0(n3557), .A1(n899), .B0(n3515), .B1(n1832), .Y(n7502) );
  OA22XL U4392 ( .A0(n3557), .A1(n900), .B0(n3515), .B1(n1833), .Y(n7492) );
  OA22XL U4393 ( .A0(n3561), .A1(n901), .B0(n3519), .B1(n1834), .Y(n7647) );
  OA22XL U4394 ( .A0(n3561), .A1(n902), .B0(n3519), .B1(n1835), .Y(n7637) );
  OA22XL U4395 ( .A0(n3561), .A1(n903), .B0(n3519), .B1(n1836), .Y(n7652) );
  OA22XL U4396 ( .A0(n3561), .A1(n904), .B0(n3519), .B1(n1837), .Y(n7642) );
  OA22XL U4397 ( .A0(n3556), .A1(n905), .B0(n3514), .B1(n1838), .Y(n7439) );
  OA22XL U4398 ( .A0(n3557), .A1(n906), .B0(n3515), .B1(n1839), .Y(n7478) );
  OA22XL U4399 ( .A0(n3550), .A1(n907), .B0(n3509), .B1(n1840), .Y(n4579) );
  OA22XL U4400 ( .A0(n3550), .A1(n908), .B0(n3509), .B1(n1841), .Y(n4569) );
  OA22XL U4401 ( .A0(n3550), .A1(n909), .B0(n3509), .B1(n1842), .Y(n4574) );
  OA22XL U4402 ( .A0(n3565), .A1(n910), .B0(n3523), .B1(n1843), .Y(n8099) );
  OA22XL U4403 ( .A0(n3565), .A1(n911), .B0(n3523), .B1(n1844), .Y(n8109) );
  OA22XL U4404 ( .A0(n3565), .A1(n912), .B0(n3523), .B1(n1845), .Y(n8115) );
  OA22XL U4405 ( .A0(n3565), .A1(n913), .B0(n3523), .B1(n1846), .Y(n8104) );
  NOR3X1 U4406 ( .A(\i_MIPS/Reg_W[0] ), .B(\i_MIPS/Reg_W[1] ), .C(n53), .Y(
        \i_MIPS/Register/n111 ) );
  NOR3X1 U4407 ( .A(n963), .B(\i_MIPS/Reg_W[1] ), .C(n53), .Y(
        \i_MIPS/Register/n109 ) );
  NOR3X1 U4408 ( .A(n78), .B(\i_MIPS/Reg_W[0] ), .C(n53), .Y(
        \i_MIPS/Register/n107 ) );
  NOR3X1 U4409 ( .A(\i_MIPS/Reg_W[0] ), .B(\i_MIPS/Reg_W[2] ), .C(n78), .Y(
        \i_MIPS/Register/n115 ) );
  NOR3X1 U4410 ( .A(n963), .B(\i_MIPS/Reg_W[2] ), .C(n78), .Y(
        \i_MIPS/Register/n113 ) );
  NOR3X1 U4411 ( .A(\i_MIPS/Reg_W[1] ), .B(\i_MIPS/Reg_W[2] ), .C(n963), .Y(
        \i_MIPS/Register/n117 ) );
  NOR3X1 U4412 ( .A(\i_MIPS/Reg_W[1] ), .B(\i_MIPS/Reg_W[2] ), .C(
        \i_MIPS/Reg_W[0] ), .Y(\i_MIPS/Register/n119 ) );
  AO21XL U4413 ( .A0(n3051), .A1(n3537), .B0(\I_cache/cache[6][154] ), .Y(
        n8926) );
  AO21XL U4414 ( .A0(n3051), .A1(n3407), .B0(\I_cache/cache[5][154] ), .Y(
        n8927) );
  AO21XL U4415 ( .A0(n3051), .A1(n3319), .B0(\I_cache/cache[3][154] ), .Y(
        n8929) );
  AO21XL U4416 ( .A0(n3051), .A1(n3362), .B0(\I_cache/cache[2][154] ), .Y(
        n8930) );
  AO21XL U4417 ( .A0(n3051), .A1(n3229), .B0(\I_cache/cache[1][154] ), .Y(
        n8931) );
  AO21XL U4418 ( .A0(n3051), .A1(n3274), .B0(\I_cache/cache[0][154] ), .Y(
        n8932) );
  AO21XL U4419 ( .A0(n3051), .A1(n3497), .B0(\I_cache/cache[7][154] ), .Y(
        n8925) );
  AO21XL U4420 ( .A0(n3051), .A1(n3452), .B0(\I_cache/cache[4][154] ), .Y(
        n8928) );
  NAND4XL U4421 ( .A(n4728), .B(n5048), .C(n4727), .D(n4726), .Y(n6983) );
  INVX3 U4422 ( .A(n3628), .Y(n3618) );
  INVX3 U4423 ( .A(n3628), .Y(n3619) );
  INVX3 U4424 ( .A(n3628), .Y(n3620) );
  INVX3 U4425 ( .A(n3628), .Y(n3621) );
  INVX3 U4426 ( .A(n3628), .Y(n3617) );
  INVX3 U4427 ( .A(n3630), .Y(n3627) );
  CLKBUFX3 U4428 ( .A(n3630), .Y(n3628) );
  CLKBUFX3 U4429 ( .A(n3630), .Y(n3629) );
  CLKBUFX3 U4430 ( .A(n3783), .Y(n3794) );
  CLKBUFX3 U4431 ( .A(n3783), .Y(n3795) );
  CLKBUFX3 U4432 ( .A(n3783), .Y(n3796) );
  CLKBUFX3 U4433 ( .A(n3792), .Y(n3802) );
  CLKBUFX3 U4434 ( .A(n3783), .Y(n3801) );
  CLKBUFX3 U4435 ( .A(n3783), .Y(n3799) );
  CLKBUFX3 U4436 ( .A(n3793), .Y(n3798) );
  CLKBUFX3 U4437 ( .A(n3783), .Y(n3800) );
  CLKBUFX3 U4438 ( .A(n3783), .Y(n3797) );
  CLKBUFX3 U4439 ( .A(n3793), .Y(n3784) );
  CLKBUFX3 U4440 ( .A(\D_cache/n206 ), .Y(n3785) );
  CLKBUFX3 U4441 ( .A(\D_cache/n206 ), .Y(n3786) );
  CLKBUFX3 U4442 ( .A(n3783), .Y(n3787) );
  CLKBUFX3 U4443 ( .A(n3783), .Y(n3788) );
  CLKBUFX3 U4444 ( .A(n3783), .Y(n3789) );
  CLKBUFX3 U4445 ( .A(n3783), .Y(n3790) );
  CLKBUFX3 U4446 ( .A(\D_cache/n206 ), .Y(n3793) );
  CLKBUFX3 U4447 ( .A(\D_cache/n206 ), .Y(n3791) );
  CLKBUFX3 U4448 ( .A(\D_cache/n206 ), .Y(n3792) );
  CLKBUFX3 U4449 ( .A(n8552), .Y(n3616) );
  CLKBUFX3 U4450 ( .A(n8333), .Y(n3582) );
  CLKBUFX3 U4451 ( .A(n8333), .Y(n3583) );
  CLKBUFX3 U4452 ( .A(n3803), .Y(n3814) );
  CLKBUFX3 U4453 ( .A(n3842), .Y(n3832) );
  CLKBUFX3 U4454 ( .A(n3843), .Y(n3854) );
  CLKBUFX3 U4455 ( .A(n3882), .Y(n3873) );
  CLKBUFX3 U4456 ( .A(n3883), .Y(n3894) );
  CLKBUFX3 U4457 ( .A(n3903), .Y(n3915) );
  CLKBUFX3 U4458 ( .A(n3924), .Y(n3936) );
  CLKBUFX3 U4459 ( .A(n3803), .Y(n3815) );
  CLKBUFX3 U4460 ( .A(n3842), .Y(n3833) );
  CLKBUFX3 U4461 ( .A(n3843), .Y(n3855) );
  CLKBUFX3 U4462 ( .A(n3882), .Y(n3874) );
  CLKBUFX3 U4463 ( .A(n3883), .Y(n3895) );
  CLKBUFX3 U4464 ( .A(n3903), .Y(n3916) );
  CLKBUFX3 U4465 ( .A(n3924), .Y(n3937) );
  CLKBUFX3 U4466 ( .A(n3803), .Y(n3816) );
  CLKBUFX3 U4467 ( .A(n3841), .Y(n3834) );
  CLKBUFX3 U4468 ( .A(n3843), .Y(n3856) );
  CLKBUFX3 U4469 ( .A(n3882), .Y(n3875) );
  CLKBUFX3 U4470 ( .A(n3883), .Y(n3896) );
  CLKBUFX3 U4471 ( .A(n3903), .Y(n3917) );
  CLKBUFX3 U4472 ( .A(n3924), .Y(n3938) );
  CLKBUFX3 U4473 ( .A(n3812), .Y(n3822) );
  CLKBUFX3 U4474 ( .A(n3823), .Y(n3839) );
  CLKBUFX3 U4475 ( .A(\D_cache/n209 ), .Y(n3862) );
  CLKBUFX3 U4476 ( .A(n3863), .Y(n3881) );
  CLKBUFX3 U4477 ( .A(n3892), .Y(n3902) );
  CLKBUFX3 U4478 ( .A(n3913), .Y(n3923) );
  CLKBUFX3 U4479 ( .A(\D_cache/n213 ), .Y(n3944) );
  CLKBUFX3 U4480 ( .A(n3803), .Y(n3821) );
  CLKBUFX3 U4481 ( .A(n3823), .Y(n3838) );
  CLKBUFX3 U4482 ( .A(n3843), .Y(n3861) );
  CLKBUFX3 U4483 ( .A(\D_cache/n210 ), .Y(n3880) );
  CLKBUFX3 U4484 ( .A(n3883), .Y(n3901) );
  CLKBUFX3 U4485 ( .A(n3903), .Y(n3922) );
  CLKBUFX3 U4486 ( .A(n3924), .Y(n3943) );
  CLKBUFX3 U4487 ( .A(n3803), .Y(n3819) );
  CLKBUFX3 U4488 ( .A(n3840), .Y(n3837) );
  CLKBUFX3 U4489 ( .A(n3843), .Y(n3859) );
  CLKBUFX3 U4490 ( .A(n3863), .Y(n3878) );
  CLKBUFX3 U4491 ( .A(n3883), .Y(n3899) );
  CLKBUFX3 U4492 ( .A(n3903), .Y(n3920) );
  CLKBUFX3 U4493 ( .A(n3924), .Y(n3941) );
  CLKBUFX3 U4494 ( .A(n3813), .Y(n3818) );
  CLKBUFX3 U4495 ( .A(n3840), .Y(n3836) );
  CLKBUFX3 U4496 ( .A(\D_cache/n209 ), .Y(n3858) );
  CLKBUFX3 U4497 ( .A(n3863), .Y(n3877) );
  CLKBUFX3 U4498 ( .A(n3893), .Y(n3898) );
  CLKBUFX3 U4499 ( .A(n3914), .Y(n3919) );
  CLKBUFX3 U4500 ( .A(\D_cache/n213 ), .Y(n3940) );
  CLKBUFX3 U4501 ( .A(n3803), .Y(n3820) );
  CLKBUFX3 U4502 ( .A(n3843), .Y(n3860) );
  CLKBUFX3 U4503 ( .A(n3863), .Y(n3879) );
  CLKBUFX3 U4504 ( .A(n3883), .Y(n3900) );
  CLKBUFX3 U4505 ( .A(n3903), .Y(n3921) );
  CLKBUFX3 U4506 ( .A(n3924), .Y(n3942) );
  CLKBUFX3 U4507 ( .A(n3803), .Y(n3817) );
  CLKBUFX3 U4508 ( .A(n3841), .Y(n3835) );
  CLKBUFX3 U4509 ( .A(n3843), .Y(n3857) );
  CLKBUFX3 U4510 ( .A(n3863), .Y(n3876) );
  CLKBUFX3 U4511 ( .A(n3883), .Y(n3897) );
  CLKBUFX3 U4512 ( .A(n3903), .Y(n3918) );
  CLKBUFX3 U4513 ( .A(n3924), .Y(n3939) );
  CLKBUFX3 U4514 ( .A(n3813), .Y(n3804) );
  CLKBUFX3 U4515 ( .A(n3893), .Y(n3884) );
  CLKBUFX3 U4516 ( .A(n3914), .Y(n3904) );
  CLKBUFX3 U4517 ( .A(\D_cache/n207 ), .Y(n3805) );
  CLKBUFX3 U4518 ( .A(n3823), .Y(n3824) );
  CLKBUFX3 U4519 ( .A(n3863), .Y(n3864) );
  CLKBUFX3 U4520 ( .A(\D_cache/n211 ), .Y(n3885) );
  CLKBUFX3 U4521 ( .A(\D_cache/n212 ), .Y(n3905) );
  CLKBUFX3 U4522 ( .A(\D_cache/n213 ), .Y(n3925) );
  CLKBUFX3 U4523 ( .A(\D_cache/n207 ), .Y(n3806) );
  CLKBUFX3 U4524 ( .A(n3823), .Y(n3825) );
  CLKBUFX3 U4525 ( .A(n3853), .Y(n3844) );
  CLKBUFX3 U4526 ( .A(n3863), .Y(n3865) );
  CLKBUFX3 U4527 ( .A(\D_cache/n211 ), .Y(n3886) );
  CLKBUFX3 U4528 ( .A(\D_cache/n212 ), .Y(n3906) );
  CLKBUFX3 U4529 ( .A(\D_cache/n213 ), .Y(n3926) );
  CLKBUFX3 U4530 ( .A(n3803), .Y(n3807) );
  CLKBUFX3 U4531 ( .A(n3823), .Y(n3826) );
  CLKBUFX3 U4532 ( .A(n3852), .Y(n3845) );
  CLKBUFX3 U4533 ( .A(n3883), .Y(n3887) );
  CLKBUFX3 U4534 ( .A(n3903), .Y(n3907) );
  CLKBUFX3 U4535 ( .A(n3924), .Y(n3927) );
  CLKBUFX3 U4536 ( .A(n3803), .Y(n3808) );
  CLKBUFX3 U4537 ( .A(n3823), .Y(n3827) );
  CLKBUFX3 U4538 ( .A(n3843), .Y(n3846) );
  CLKBUFX3 U4539 ( .A(n3883), .Y(n3888) );
  CLKBUFX3 U4540 ( .A(n3903), .Y(n3908) );
  CLKBUFX3 U4541 ( .A(n3924), .Y(n3928) );
  CLKBUFX3 U4542 ( .A(n3803), .Y(n3809) );
  CLKBUFX3 U4543 ( .A(n3823), .Y(n3828) );
  CLKBUFX3 U4544 ( .A(n3843), .Y(n3847) );
  CLKBUFX3 U4545 ( .A(n3863), .Y(n3866) );
  CLKBUFX3 U4546 ( .A(n3883), .Y(n3889) );
  CLKBUFX3 U4547 ( .A(n3903), .Y(n3909) );
  CLKBUFX3 U4548 ( .A(n3924), .Y(n3929) );
  CLKBUFX3 U4549 ( .A(n3803), .Y(n3810) );
  CLKBUFX3 U4550 ( .A(n3843), .Y(n3848) );
  CLKBUFX3 U4551 ( .A(n3863), .Y(n3867) );
  CLKBUFX3 U4552 ( .A(n3883), .Y(n3890) );
  CLKBUFX3 U4553 ( .A(n3903), .Y(n3910) );
  CLKBUFX3 U4554 ( .A(\D_cache/n213 ), .Y(n3930) );
  CLKBUFX3 U4555 ( .A(\D_cache/n207 ), .Y(n3813) );
  CLKBUFX3 U4556 ( .A(n3823), .Y(n3831) );
  CLKBUFX3 U4557 ( .A(\D_cache/n209 ), .Y(n3853) );
  CLKBUFX3 U4558 ( .A(n3863), .Y(n3872) );
  CLKBUFX3 U4559 ( .A(\D_cache/n211 ), .Y(n3893) );
  CLKBUFX3 U4560 ( .A(\D_cache/n212 ), .Y(n3914) );
  CLKBUFX3 U4561 ( .A(n3924), .Y(n3935) );
  CLKBUFX3 U4562 ( .A(n3823), .Y(n3830) );
  CLKBUFX3 U4563 ( .A(n3843), .Y(n3851) );
  CLKBUFX3 U4564 ( .A(n3863), .Y(n3870) );
  CLKBUFX3 U4565 ( .A(n3924), .Y(n3933) );
  CLKBUFX3 U4566 ( .A(n3843), .Y(n3850) );
  CLKBUFX3 U4567 ( .A(n3863), .Y(n3869) );
  CLKBUFX3 U4568 ( .A(n3903), .Y(n3912) );
  CLKBUFX3 U4569 ( .A(n3924), .Y(n3932) );
  CLKBUFX3 U4570 ( .A(\D_cache/n207 ), .Y(n3811) );
  CLKBUFX3 U4571 ( .A(n3823), .Y(n3829) );
  CLKBUFX3 U4572 ( .A(n3843), .Y(n3849) );
  CLKBUFX3 U4573 ( .A(n3863), .Y(n3868) );
  CLKBUFX3 U4574 ( .A(\D_cache/n211 ), .Y(n3891) );
  CLKBUFX3 U4575 ( .A(\D_cache/n212 ), .Y(n3911) );
  CLKBUFX3 U4576 ( .A(n3924), .Y(n3931) );
  CLKBUFX3 U4577 ( .A(\D_cache/n207 ), .Y(n3812) );
  CLKBUFX3 U4578 ( .A(\D_cache/n209 ), .Y(n3852) );
  CLKBUFX3 U4579 ( .A(n3863), .Y(n3871) );
  CLKBUFX3 U4580 ( .A(\D_cache/n211 ), .Y(n3892) );
  CLKBUFX3 U4581 ( .A(\D_cache/n212 ), .Y(n3913) );
  CLKBUFX3 U4582 ( .A(n3924), .Y(n3934) );
  INVX3 U4583 ( .A(n3546), .Y(n3532) );
  INVX3 U4584 ( .A(n3543), .Y(n3535) );
  INVX3 U4585 ( .A(n3551), .Y(n3538) );
  INVX3 U4586 ( .A(n3551), .Y(n3537) );
  INVX3 U4587 ( .A(n3542), .Y(n3536) );
  INVX3 U4588 ( .A(n3545), .Y(n3533) );
  INVX3 U4589 ( .A(n3544), .Y(n3534) );
  INVX3 U4590 ( .A(n3328), .Y(n3310) );
  INVX3 U4591 ( .A(n3325), .Y(n3313) );
  INVX3 U4592 ( .A(n3323), .Y(n3315) );
  INVX3 U4593 ( .A(n3324), .Y(n3314) );
  INVX3 U4594 ( .A(n3327), .Y(n3311) );
  INVX3 U4595 ( .A(n3321), .Y(n3317) );
  INVX3 U4596 ( .A(n3326), .Y(n3312) );
  CLKINVX1 U4597 ( .A(n6845), .Y(n6476) );
  CLKBUFX3 U4598 ( .A(n3572), .Y(n3542) );
  CLKBUFX3 U4599 ( .A(n3571), .Y(n3546) );
  CLKBUFX3 U4600 ( .A(n3571), .Y(n3545) );
  CLKBUFX3 U4601 ( .A(n3571), .Y(n3544) );
  CLKBUFX3 U4602 ( .A(n3571), .Y(n3543) );
  CLKBUFX3 U4603 ( .A(n3352), .Y(n3324) );
  CLKBUFX3 U4604 ( .A(n3329), .Y(n3320) );
  CLKBUFX3 U4605 ( .A(n3352), .Y(n3322) );
  CLKBUFX3 U4606 ( .A(n3351), .Y(n3328) );
  CLKBUFX3 U4607 ( .A(n3351), .Y(n3327) );
  CLKBUFX3 U4608 ( .A(n3351), .Y(n3326) );
  CLKBUFX3 U4609 ( .A(n3351), .Y(n3325) );
  CLKBUFX3 U4610 ( .A(n3352), .Y(n3323) );
  CLKBUFX3 U4611 ( .A(n3566), .Y(n3550) );
  CLKBUFX3 U4612 ( .A(n3569), .Y(n3554) );
  CLKBUFX3 U4613 ( .A(n3568), .Y(n3555) );
  CLKBUFX3 U4614 ( .A(n3567), .Y(n3559) );
  CLKBUFX3 U4615 ( .A(n3567), .Y(n3558) );
  CLKBUFX3 U4616 ( .A(n3350), .Y(n3332) );
  CLKBUFX3 U4617 ( .A(n3350), .Y(n3335) );
  CLKBUFX3 U4618 ( .A(n3349), .Y(n3336) );
  CLKBUFX3 U4619 ( .A(n3348), .Y(n3340) );
  CLKBUFX3 U4620 ( .A(n3348), .Y(n3339) );
  CLKBUFX3 U4621 ( .A(n8457), .Y(n3613) );
  CLKBUFX3 U4622 ( .A(n8457), .Y(n3612) );
  CLKBUFX3 U4623 ( .A(n3569), .Y(n3553) );
  CLKBUFX3 U4624 ( .A(n3568), .Y(n3556) );
  CLKBUFX3 U4625 ( .A(n3566), .Y(n3564) );
  CLKBUFX3 U4626 ( .A(n3566), .Y(n3563) );
  CLKBUFX3 U4627 ( .A(n3566), .Y(n3562) );
  CLKBUFX3 U4628 ( .A(n3567), .Y(n3561) );
  CLKBUFX3 U4629 ( .A(n3567), .Y(n3560) );
  CLKBUFX3 U4630 ( .A(n3568), .Y(n3557) );
  CLKBUFX3 U4631 ( .A(n3350), .Y(n3334) );
  CLKBUFX3 U4632 ( .A(n3349), .Y(n3337) );
  CLKBUFX3 U4633 ( .A(n3347), .Y(n3345) );
  CLKBUFX3 U4634 ( .A(n3347), .Y(n3344) );
  CLKBUFX3 U4635 ( .A(n3347), .Y(n3343) );
  CLKBUFX3 U4636 ( .A(n3348), .Y(n3342) );
  CLKBUFX3 U4637 ( .A(n3348), .Y(n3341) );
  CLKBUFX3 U4638 ( .A(n3349), .Y(n3338) );
  CLKBUFX3 U4639 ( .A(n3566), .Y(n3565) );
  CLKBUFX3 U4640 ( .A(n3347), .Y(n3346) );
  CLKBUFX3 U4641 ( .A(n2764), .Y(n3186) );
  CLKBUFX3 U4642 ( .A(n2764), .Y(n3187) );
  CLKBUFX3 U4643 ( .A(n2763), .Y(n3136) );
  CLKBUFX3 U4644 ( .A(n2764), .Y(n3185) );
  CLKBUFX3 U4645 ( .A(n2763), .Y(n3135) );
  CLKBUFX3 U4646 ( .A(n2763), .Y(n3134) );
  CLKBUFX3 U4647 ( .A(n3586), .Y(n3588) );
  CLKBUFX3 U4648 ( .A(n3586), .Y(n3590) );
  CLKBUFX3 U4649 ( .A(n3586), .Y(n3587) );
  CLKBUFX3 U4650 ( .A(n3586), .Y(n3591) );
  CLKBUFX3 U4651 ( .A(n3586), .Y(n3589) );
  INVX3 U4652 ( .A(n2808), .Y(n3977) );
  INVX3 U4653 ( .A(n2808), .Y(n3978) );
  CLKBUFX3 U4654 ( .A(n3569), .Y(n3552) );
  CLKBUFX3 U4655 ( .A(n3570), .Y(n3551) );
  CLKBUFX3 U4656 ( .A(n3350), .Y(n3333) );
  INVX3 U4657 ( .A(n3956), .Y(n3949) );
  INVX3 U4658 ( .A(n3956), .Y(n3947) );
  INVX3 U4659 ( .A(n3956), .Y(n3951) );
  INVX3 U4660 ( .A(n3956), .Y(n3952) );
  INVX3 U4661 ( .A(n3956), .Y(n3950) );
  INVX3 U4662 ( .A(n3970), .Y(n3953) );
  INVX3 U4663 ( .A(n3971), .Y(n3948) );
  INVX3 U4664 ( .A(n3970), .Y(n3946) );
  INVX3 U4665 ( .A(n3970), .Y(n3945) );
  INVX3 U4666 ( .A(n3955), .Y(n3954) );
  CLKBUFX3 U4667 ( .A(n8453), .Y(n3604) );
  CLKBUFX3 U4668 ( .A(n8453), .Y(n3605) );
  CLKBUFX3 U4669 ( .A(n8453), .Y(n3606) );
  CLKBUFX3 U4670 ( .A(n8453), .Y(n3607) );
  CLKBUFX3 U4671 ( .A(n8453), .Y(n3608) );
  CLKBUFX3 U4672 ( .A(n8453), .Y(n3609) );
  INVX3 U4673 ( .A(n3454), .Y(n3451) );
  INVX3 U4674 ( .A(n3479), .Y(n3443) );
  INVX3 U4675 ( .A(n3371), .Y(n3353) );
  INVX3 U4676 ( .A(n3284), .Y(n3265) );
  INVX3 U4677 ( .A(n3278), .Y(n3271) );
  INVX3 U4678 ( .A(n3460), .Y(n3445) );
  INVX3 U4679 ( .A(n3368), .Y(n3356) );
  INVX3 U4680 ( .A(n3281), .Y(n3268) );
  INVX3 U4681 ( .A(n3457), .Y(n3448) );
  INVX3 U4682 ( .A(n3366), .Y(n3358) );
  INVX3 U4683 ( .A(n3456), .Y(n3449) );
  INVX3 U4684 ( .A(n3458), .Y(n3447) );
  INVX3 U4685 ( .A(n3367), .Y(n3357) );
  INVX3 U4686 ( .A(n3459), .Y(n3446) );
  INVX3 U4687 ( .A(n3370), .Y(n3354) );
  INVX3 U4688 ( .A(n3283), .Y(n3266) );
  INVX3 U4689 ( .A(n3455), .Y(n3450) );
  INVX3 U4690 ( .A(n3364), .Y(n3360) );
  INVX3 U4691 ( .A(n3453), .Y(n3452) );
  INVX3 U4692 ( .A(n3461), .Y(n3444) );
  INVX3 U4693 ( .A(n3369), .Y(n3355) );
  INVX3 U4694 ( .A(n3282), .Y(n3267) );
  INVX3 U4695 ( .A(n3410), .Y(n3405) );
  INVX3 U4696 ( .A(n3505), .Y(n3488) );
  INVX3 U4697 ( .A(n3418), .Y(n3398) );
  INVX3 U4698 ( .A(n3236), .Y(n3220) );
  INVX3 U4699 ( .A(n3502), .Y(n3491) );
  INVX3 U4700 ( .A(n3233), .Y(n3223) );
  INVX3 U4701 ( .A(n3500), .Y(n3493) );
  INVX3 U4702 ( .A(n3418), .Y(n3403) );
  INVX3 U4703 ( .A(n3232), .Y(n3225) );
  INVX3 U4704 ( .A(n3418), .Y(n3404) );
  INVX3 U4705 ( .A(n3501), .Y(n3492) );
  INVX3 U4706 ( .A(n3411), .Y(n3402) );
  INVX3 U4707 ( .A(n3412), .Y(n3401) );
  INVX3 U4708 ( .A(n3504), .Y(n3489) );
  INVX3 U4709 ( .A(n3414), .Y(n3399) );
  INVX3 U4710 ( .A(n3235), .Y(n3221) );
  INVX3 U4711 ( .A(n3498), .Y(n3495) );
  INVX3 U4712 ( .A(n3409), .Y(n3406) );
  INVX3 U4713 ( .A(n3231), .Y(n3227) );
  INVX3 U4714 ( .A(n3503), .Y(n3490) );
  INVX3 U4715 ( .A(n3413), .Y(n3400) );
  INVX3 U4716 ( .A(n3234), .Y(n3222) );
  INVX3 U4717 ( .A(n3408), .Y(n3407) );
  CLKBUFX3 U4718 ( .A(\D_cache/n206 ), .Y(n3783) );
  CLKBUFX3 U4719 ( .A(n3863), .Y(n3882) );
  CLKBUFX3 U4720 ( .A(n3823), .Y(n3842) );
  CLKBUFX3 U4721 ( .A(n3823), .Y(n3840) );
  CLKBUFX3 U4722 ( .A(n3823), .Y(n3841) );
  CLKBUFX3 U4723 ( .A(n4361), .Y(n4359) );
  CLKBUFX3 U4724 ( .A(n4361), .Y(n4358) );
  CLKBUFX3 U4725 ( .A(n4361), .Y(n4357) );
  CLKBUFX3 U4726 ( .A(n4361), .Y(n4356) );
  CLKBUFX3 U4727 ( .A(n4361), .Y(n4355) );
  CLKBUFX3 U4728 ( .A(n4361), .Y(n4354) );
  CLKBUFX3 U4729 ( .A(n4361), .Y(n4353) );
  CLKBUFX3 U4730 ( .A(n4361), .Y(n4352) );
  CLKBUFX3 U4731 ( .A(n4361), .Y(n4351) );
  CLKBUFX3 U4732 ( .A(n4361), .Y(n4350) );
  CLKBUFX3 U4733 ( .A(n4361), .Y(n4349) );
  CLKBUFX3 U4734 ( .A(n4360), .Y(n4348) );
  CLKBUFX3 U4735 ( .A(n4361), .Y(n4347) );
  CLKBUFX3 U4736 ( .A(n4366), .Y(n4346) );
  CLKBUFX3 U4737 ( .A(n4362), .Y(n4345) );
  CLKBUFX3 U4738 ( .A(n4370), .Y(n4344) );
  CLKBUFX3 U4739 ( .A(n4373), .Y(n4343) );
  CLKBUFX3 U4740 ( .A(n4371), .Y(n4342) );
  CLKBUFX3 U4741 ( .A(n4379), .Y(n4341) );
  CLKBUFX3 U4742 ( .A(n4360), .Y(n4340) );
  CLKBUFX3 U4743 ( .A(n4361), .Y(n4339) );
  CLKBUFX3 U4744 ( .A(n4386), .Y(n4338) );
  CLKBUFX3 U4745 ( .A(n4364), .Y(n4337) );
  CLKBUFX3 U4746 ( .A(n4362), .Y(n4336) );
  CLKBUFX3 U4747 ( .A(n4362), .Y(n4335) );
  CLKBUFX3 U4748 ( .A(n4362), .Y(n4334) );
  CLKBUFX3 U4749 ( .A(n4362), .Y(n4333) );
  CLKBUFX3 U4750 ( .A(n4362), .Y(n4332) );
  CLKBUFX3 U4751 ( .A(n4362), .Y(n4331) );
  CLKBUFX3 U4752 ( .A(n4362), .Y(n4330) );
  CLKBUFX3 U4753 ( .A(n4362), .Y(n4329) );
  CLKBUFX3 U4754 ( .A(n4362), .Y(n4328) );
  CLKBUFX3 U4755 ( .A(n4362), .Y(n4327) );
  CLKBUFX3 U4756 ( .A(n4362), .Y(n4326) );
  CLKBUFX3 U4757 ( .A(n4362), .Y(n4325) );
  CLKBUFX3 U4758 ( .A(n4363), .Y(n4324) );
  CLKBUFX3 U4759 ( .A(n4363), .Y(n4323) );
  CLKBUFX3 U4760 ( .A(n4363), .Y(n4322) );
  CLKBUFX3 U4761 ( .A(n4363), .Y(n4321) );
  CLKBUFX3 U4762 ( .A(n4363), .Y(n4320) );
  CLKBUFX3 U4763 ( .A(n4363), .Y(n4319) );
  CLKBUFX3 U4764 ( .A(n4363), .Y(n4318) );
  CLKBUFX3 U4765 ( .A(n4363), .Y(n4317) );
  CLKBUFX3 U4766 ( .A(n4363), .Y(n4316) );
  CLKBUFX3 U4767 ( .A(n4363), .Y(n4315) );
  CLKBUFX3 U4768 ( .A(n4363), .Y(n4314) );
  CLKBUFX3 U4769 ( .A(n4363), .Y(n4313) );
  CLKBUFX3 U4770 ( .A(n4364), .Y(n4312) );
  CLKBUFX3 U4771 ( .A(n4364), .Y(n4311) );
  CLKBUFX3 U4772 ( .A(n4364), .Y(n4310) );
  CLKBUFX3 U4773 ( .A(n4364), .Y(n4309) );
  CLKBUFX3 U4774 ( .A(n4364), .Y(n4308) );
  CLKBUFX3 U4775 ( .A(n4364), .Y(n4307) );
  CLKBUFX3 U4776 ( .A(n4364), .Y(n4306) );
  CLKBUFX3 U4777 ( .A(n4364), .Y(n4305) );
  CLKBUFX3 U4778 ( .A(n4364), .Y(n4304) );
  CLKBUFX3 U4779 ( .A(n4364), .Y(n4303) );
  CLKBUFX3 U4780 ( .A(n4364), .Y(n4302) );
  CLKBUFX3 U4781 ( .A(n4364), .Y(n4301) );
  CLKBUFX3 U4782 ( .A(n4365), .Y(n4300) );
  CLKBUFX3 U4783 ( .A(n4365), .Y(n4299) );
  CLKBUFX3 U4784 ( .A(n4365), .Y(n4298) );
  CLKBUFX3 U4785 ( .A(n4365), .Y(n4297) );
  CLKBUFX3 U4786 ( .A(n4365), .Y(n4296) );
  CLKBUFX3 U4787 ( .A(n4365), .Y(n4295) );
  CLKBUFX3 U4788 ( .A(n4365), .Y(n4294) );
  CLKBUFX3 U4789 ( .A(n4365), .Y(n4293) );
  CLKBUFX3 U4790 ( .A(n4365), .Y(n4292) );
  CLKBUFX3 U4791 ( .A(n4365), .Y(n4291) );
  CLKBUFX3 U4792 ( .A(n4365), .Y(n4290) );
  CLKBUFX3 U4793 ( .A(n4365), .Y(n4289) );
  CLKBUFX3 U4794 ( .A(n4366), .Y(n4288) );
  CLKBUFX3 U4795 ( .A(n4366), .Y(n4287) );
  CLKBUFX3 U4796 ( .A(n4366), .Y(n4286) );
  CLKBUFX3 U4797 ( .A(n4366), .Y(n4285) );
  CLKBUFX3 U4798 ( .A(n4366), .Y(n4284) );
  CLKBUFX3 U4799 ( .A(n4366), .Y(n4283) );
  CLKBUFX3 U4800 ( .A(n4366), .Y(n4282) );
  CLKBUFX3 U4801 ( .A(n4366), .Y(n4281) );
  CLKBUFX3 U4802 ( .A(n4366), .Y(n4280) );
  CLKBUFX3 U4803 ( .A(n4366), .Y(n4279) );
  CLKBUFX3 U4804 ( .A(n4366), .Y(n4278) );
  CLKBUFX3 U4805 ( .A(n4366), .Y(n4277) );
  CLKBUFX3 U4806 ( .A(n4367), .Y(n4276) );
  CLKBUFX3 U4807 ( .A(n4367), .Y(n4275) );
  CLKBUFX3 U4808 ( .A(n4367), .Y(n4274) );
  CLKBUFX3 U4809 ( .A(n4367), .Y(n4273) );
  CLKBUFX3 U4810 ( .A(n4367), .Y(n4272) );
  CLKBUFX3 U4811 ( .A(n4367), .Y(n4271) );
  CLKBUFX3 U4812 ( .A(n4367), .Y(n4270) );
  CLKBUFX3 U4813 ( .A(n4367), .Y(n4269) );
  CLKBUFX3 U4814 ( .A(n4367), .Y(n4268) );
  CLKBUFX3 U4815 ( .A(n4367), .Y(n4267) );
  CLKBUFX3 U4816 ( .A(n4367), .Y(n4266) );
  CLKBUFX3 U4817 ( .A(n4367), .Y(n4265) );
  CLKBUFX3 U4818 ( .A(n4368), .Y(n4264) );
  CLKBUFX3 U4819 ( .A(n4368), .Y(n4263) );
  CLKBUFX3 U4820 ( .A(n4368), .Y(n4262) );
  CLKBUFX3 U4821 ( .A(n4368), .Y(n4261) );
  CLKBUFX3 U4822 ( .A(n4368), .Y(n4260) );
  CLKBUFX3 U4823 ( .A(n4368), .Y(n4259) );
  CLKBUFX3 U4824 ( .A(n4368), .Y(n4258) );
  CLKBUFX3 U4825 ( .A(n4377), .Y(n4153) );
  CLKBUFX3 U4826 ( .A(n4377), .Y(n4152) );
  CLKBUFX3 U4827 ( .A(n4377), .Y(n4151) );
  CLKBUFX3 U4828 ( .A(n4377), .Y(n4150) );
  CLKBUFX3 U4829 ( .A(n4377), .Y(n4149) );
  CLKBUFX3 U4830 ( .A(n4377), .Y(n4148) );
  CLKBUFX3 U4831 ( .A(n4377), .Y(n4147) );
  CLKBUFX3 U4832 ( .A(n4377), .Y(n4146) );
  CLKBUFX3 U4833 ( .A(n4377), .Y(n4145) );
  CLKBUFX3 U4834 ( .A(n4378), .Y(n4144) );
  CLKBUFX3 U4835 ( .A(n4378), .Y(n4143) );
  CLKBUFX3 U4836 ( .A(n4378), .Y(n4142) );
  CLKBUFX3 U4837 ( .A(n4378), .Y(n4141) );
  CLKBUFX3 U4838 ( .A(n4378), .Y(n4140) );
  CLKBUFX3 U4839 ( .A(n4378), .Y(n4139) );
  CLKBUFX3 U4840 ( .A(n4378), .Y(n4138) );
  CLKBUFX3 U4841 ( .A(n4378), .Y(n4137) );
  CLKBUFX3 U4842 ( .A(n4378), .Y(n4136) );
  CLKBUFX3 U4843 ( .A(n4378), .Y(n4135) );
  CLKBUFX3 U4844 ( .A(n4378), .Y(n4134) );
  CLKBUFX3 U4845 ( .A(n4378), .Y(n4133) );
  CLKBUFX3 U4846 ( .A(n4379), .Y(n4132) );
  CLKBUFX3 U4847 ( .A(n4379), .Y(n4131) );
  CLKBUFX3 U4848 ( .A(n4379), .Y(n4130) );
  CLKBUFX3 U4849 ( .A(n4379), .Y(n4129) );
  CLKBUFX3 U4850 ( .A(n4379), .Y(n4128) );
  CLKBUFX3 U4851 ( .A(n4379), .Y(n4127) );
  CLKBUFX3 U4852 ( .A(n4379), .Y(n4126) );
  CLKBUFX3 U4853 ( .A(n4379), .Y(n4125) );
  CLKBUFX3 U4854 ( .A(n4379), .Y(n4124) );
  CLKBUFX3 U4855 ( .A(n4379), .Y(n4123) );
  CLKBUFX3 U4856 ( .A(n4379), .Y(n4122) );
  CLKBUFX3 U4857 ( .A(n4379), .Y(n4121) );
  CLKBUFX3 U4858 ( .A(n4380), .Y(n4120) );
  CLKBUFX3 U4859 ( .A(n4380), .Y(n4119) );
  CLKBUFX3 U4860 ( .A(n4380), .Y(n4118) );
  CLKBUFX3 U4861 ( .A(n4380), .Y(n4117) );
  CLKBUFX3 U4862 ( .A(n4380), .Y(n4116) );
  CLKBUFX3 U4863 ( .A(n4380), .Y(n4115) );
  CLKBUFX3 U4864 ( .A(n4380), .Y(n4114) );
  CLKBUFX3 U4865 ( .A(n4380), .Y(n4113) );
  CLKBUFX3 U4866 ( .A(n4380), .Y(n4112) );
  CLKBUFX3 U4867 ( .A(n4380), .Y(n4111) );
  CLKBUFX3 U4868 ( .A(n4380), .Y(n4110) );
  CLKBUFX3 U4869 ( .A(n4380), .Y(n4109) );
  CLKBUFX3 U4870 ( .A(n4381), .Y(n4108) );
  CLKBUFX3 U4871 ( .A(n4381), .Y(n4107) );
  CLKBUFX3 U4872 ( .A(n4381), .Y(n4106) );
  CLKBUFX3 U4873 ( .A(n4381), .Y(n4105) );
  CLKBUFX3 U4874 ( .A(n4381), .Y(n4104) );
  CLKBUFX3 U4875 ( .A(n4381), .Y(n4103) );
  CLKBUFX3 U4876 ( .A(n4381), .Y(n4102) );
  CLKBUFX3 U4877 ( .A(n4381), .Y(n4101) );
  CLKBUFX3 U4878 ( .A(n4381), .Y(n4100) );
  CLKBUFX3 U4879 ( .A(n4381), .Y(n4099) );
  CLKBUFX3 U4880 ( .A(n4381), .Y(n4098) );
  CLKBUFX3 U4881 ( .A(n4381), .Y(n4097) );
  CLKBUFX3 U4882 ( .A(n4382), .Y(n4096) );
  CLKBUFX3 U4883 ( .A(n4382), .Y(n4095) );
  CLKBUFX3 U4884 ( .A(n4382), .Y(n4094) );
  CLKBUFX3 U4885 ( .A(n4382), .Y(n4093) );
  CLKBUFX3 U4886 ( .A(n4382), .Y(n4092) );
  CLKBUFX3 U4887 ( .A(n4382), .Y(n4091) );
  CLKBUFX3 U4888 ( .A(n4382), .Y(n4090) );
  CLKBUFX3 U4889 ( .A(n4382), .Y(n4089) );
  CLKBUFX3 U4890 ( .A(n4382), .Y(n4088) );
  CLKBUFX3 U4891 ( .A(n4382), .Y(n4087) );
  CLKBUFX3 U4892 ( .A(n4382), .Y(n4086) );
  CLKBUFX3 U4893 ( .A(n4382), .Y(n4085) );
  CLKBUFX3 U4894 ( .A(n4383), .Y(n4084) );
  CLKBUFX3 U4895 ( .A(n4383), .Y(n4083) );
  CLKBUFX3 U4896 ( .A(n4383), .Y(n4082) );
  CLKBUFX3 U4897 ( .A(n4383), .Y(n4081) );
  CLKBUFX3 U4898 ( .A(n4383), .Y(n4080) );
  CLKBUFX3 U4899 ( .A(n4383), .Y(n4079) );
  CLKBUFX3 U4900 ( .A(n4383), .Y(n4078) );
  CLKBUFX3 U4901 ( .A(n4383), .Y(n4077) );
  CLKBUFX3 U4902 ( .A(n4383), .Y(n4076) );
  CLKBUFX3 U4903 ( .A(n4383), .Y(n4075) );
  CLKBUFX3 U4904 ( .A(n4383), .Y(n4074) );
  CLKBUFX3 U4905 ( .A(n4383), .Y(n4073) );
  CLKBUFX3 U4906 ( .A(n4368), .Y(n4257) );
  CLKBUFX3 U4907 ( .A(n4368), .Y(n4256) );
  CLKBUFX3 U4908 ( .A(n4368), .Y(n4255) );
  CLKBUFX3 U4909 ( .A(n4368), .Y(n4254) );
  CLKBUFX3 U4910 ( .A(n4368), .Y(n4253) );
  CLKBUFX3 U4911 ( .A(n4369), .Y(n4252) );
  CLKBUFX3 U4912 ( .A(n4369), .Y(n4251) );
  CLKBUFX3 U4913 ( .A(n4369), .Y(n4250) );
  CLKBUFX3 U4914 ( .A(n4369), .Y(n4249) );
  CLKBUFX3 U4915 ( .A(n4369), .Y(n4248) );
  CLKBUFX3 U4916 ( .A(n4369), .Y(n4247) );
  CLKBUFX3 U4917 ( .A(n4369), .Y(n4246) );
  CLKBUFX3 U4918 ( .A(n4369), .Y(n4245) );
  CLKBUFX3 U4919 ( .A(n4369), .Y(n4244) );
  CLKBUFX3 U4920 ( .A(n4369), .Y(n4243) );
  CLKBUFX3 U4921 ( .A(n4369), .Y(n4242) );
  CLKBUFX3 U4922 ( .A(n4369), .Y(n4241) );
  CLKBUFX3 U4923 ( .A(n4370), .Y(n4240) );
  CLKBUFX3 U4924 ( .A(n4370), .Y(n4239) );
  CLKBUFX3 U4925 ( .A(n4370), .Y(n4238) );
  CLKBUFX3 U4926 ( .A(n4370), .Y(n4237) );
  CLKBUFX3 U4927 ( .A(n4370), .Y(n4236) );
  CLKBUFX3 U4928 ( .A(n4370), .Y(n4235) );
  CLKBUFX3 U4929 ( .A(n4370), .Y(n4234) );
  CLKBUFX3 U4930 ( .A(n4370), .Y(n4233) );
  CLKBUFX3 U4931 ( .A(n4370), .Y(n4232) );
  CLKBUFX3 U4932 ( .A(n4370), .Y(n4231) );
  CLKBUFX3 U4933 ( .A(n4370), .Y(n4230) );
  CLKBUFX3 U4934 ( .A(n4370), .Y(n4229) );
  CLKBUFX3 U4935 ( .A(n4371), .Y(n4228) );
  CLKBUFX3 U4936 ( .A(n4371), .Y(n4227) );
  CLKBUFX3 U4937 ( .A(n4371), .Y(n4226) );
  CLKBUFX3 U4938 ( .A(n4371), .Y(n4225) );
  CLKBUFX3 U4939 ( .A(n4371), .Y(n4224) );
  CLKBUFX3 U4940 ( .A(n4371), .Y(n4223) );
  CLKBUFX3 U4941 ( .A(n4371), .Y(n4222) );
  CLKBUFX3 U4942 ( .A(n4371), .Y(n4221) );
  CLKBUFX3 U4943 ( .A(n4371), .Y(n4220) );
  CLKBUFX3 U4944 ( .A(n4371), .Y(n4219) );
  CLKBUFX3 U4945 ( .A(n4371), .Y(n4218) );
  CLKBUFX3 U4946 ( .A(n4371), .Y(n4217) );
  CLKBUFX3 U4947 ( .A(n4372), .Y(n4216) );
  CLKBUFX3 U4948 ( .A(n4372), .Y(n4215) );
  CLKBUFX3 U4949 ( .A(n4372), .Y(n4214) );
  CLKBUFX3 U4950 ( .A(n4372), .Y(n4213) );
  CLKBUFX3 U4951 ( .A(n4372), .Y(n4212) );
  CLKBUFX3 U4952 ( .A(n4372), .Y(n4211) );
  CLKBUFX3 U4953 ( .A(n4372), .Y(n4210) );
  CLKBUFX3 U4954 ( .A(n4372), .Y(n4209) );
  CLKBUFX3 U4955 ( .A(n4372), .Y(n4208) );
  CLKBUFX3 U4956 ( .A(n4372), .Y(n4207) );
  CLKBUFX3 U4957 ( .A(n4372), .Y(n4206) );
  CLKBUFX3 U4958 ( .A(n4372), .Y(n4205) );
  CLKBUFX3 U4959 ( .A(n4373), .Y(n4204) );
  CLKBUFX3 U4960 ( .A(n4373), .Y(n4203) );
  CLKBUFX3 U4961 ( .A(n4373), .Y(n4202) );
  CLKBUFX3 U4962 ( .A(n4373), .Y(n4201) );
  CLKBUFX3 U4963 ( .A(n4373), .Y(n4200) );
  CLKBUFX3 U4964 ( .A(n4373), .Y(n4199) );
  CLKBUFX3 U4965 ( .A(n4373), .Y(n4198) );
  CLKBUFX3 U4966 ( .A(n4373), .Y(n4197) );
  CLKBUFX3 U4967 ( .A(n4373), .Y(n4196) );
  CLKBUFX3 U4968 ( .A(n4373), .Y(n4195) );
  CLKBUFX3 U4969 ( .A(n4373), .Y(n4194) );
  CLKBUFX3 U4970 ( .A(n4373), .Y(n4193) );
  CLKBUFX3 U4971 ( .A(n4374), .Y(n4192) );
  CLKBUFX3 U4972 ( .A(n4374), .Y(n4191) );
  CLKBUFX3 U4973 ( .A(n4374), .Y(n4190) );
  CLKBUFX3 U4974 ( .A(n4374), .Y(n4189) );
  CLKBUFX3 U4975 ( .A(n4374), .Y(n4188) );
  CLKBUFX3 U4976 ( .A(n4374), .Y(n4187) );
  CLKBUFX3 U4977 ( .A(n4374), .Y(n4186) );
  CLKBUFX3 U4978 ( .A(n4374), .Y(n4185) );
  CLKBUFX3 U4979 ( .A(n4374), .Y(n4184) );
  CLKBUFX3 U4980 ( .A(n4374), .Y(n4183) );
  CLKBUFX3 U4981 ( .A(n4374), .Y(n4182) );
  CLKBUFX3 U4982 ( .A(n4374), .Y(n4181) );
  CLKBUFX3 U4983 ( .A(n4375), .Y(n4180) );
  CLKBUFX3 U4984 ( .A(n4375), .Y(n4179) );
  CLKBUFX3 U4985 ( .A(n4375), .Y(n4178) );
  CLKBUFX3 U4986 ( .A(n4375), .Y(n4177) );
  CLKBUFX3 U4987 ( .A(n4375), .Y(n4176) );
  CLKBUFX3 U4988 ( .A(n4375), .Y(n4175) );
  CLKBUFX3 U4989 ( .A(n4375), .Y(n4174) );
  CLKBUFX3 U4990 ( .A(n4375), .Y(n4173) );
  CLKBUFX3 U4991 ( .A(n4375), .Y(n4172) );
  CLKBUFX3 U4992 ( .A(n4375), .Y(n4171) );
  CLKBUFX3 U4993 ( .A(n4375), .Y(n4170) );
  CLKBUFX3 U4994 ( .A(n4375), .Y(n4169) );
  CLKBUFX3 U4995 ( .A(n4376), .Y(n4168) );
  CLKBUFX3 U4996 ( .A(n4376), .Y(n4167) );
  CLKBUFX3 U4997 ( .A(n4376), .Y(n4166) );
  CLKBUFX3 U4998 ( .A(n4376), .Y(n4165) );
  CLKBUFX3 U4999 ( .A(n4376), .Y(n4164) );
  CLKBUFX3 U5000 ( .A(n4376), .Y(n4163) );
  CLKBUFX3 U5001 ( .A(n4376), .Y(n4162) );
  CLKBUFX3 U5002 ( .A(n4376), .Y(n4161) );
  CLKBUFX3 U5003 ( .A(n4376), .Y(n4160) );
  CLKBUFX3 U5004 ( .A(n4376), .Y(n4159) );
  CLKBUFX3 U5005 ( .A(n4376), .Y(n4158) );
  CLKBUFX3 U5006 ( .A(n4376), .Y(n4157) );
  CLKBUFX3 U5007 ( .A(n4377), .Y(n4156) );
  CLKBUFX3 U5008 ( .A(n4377), .Y(n4155) );
  CLKBUFX3 U5009 ( .A(n4377), .Y(n4154) );
  CLKBUFX3 U5010 ( .A(n4361), .Y(n4360) );
  CLKBUFX3 U5011 ( .A(n3687), .Y(n3038) );
  NAND2X1 U5012 ( .A(n6848), .B(n4909), .Y(n6918) );
  NAND2X1 U5013 ( .A(n4983), .B(n4016), .Y(n5614) );
  OAI221XL U5014 ( .A0(n3106), .A1(n5540), .B0(n2823), .B1(n3098), .C0(n3097), 
        .Y(n5541) );
  CLKINVX1 U5015 ( .A(n4820), .Y(n6832) );
  NAND2X1 U5016 ( .A(n4016), .B(n6905), .Y(n5888) );
  CLKINVX1 U5017 ( .A(n6908), .Y(n6774) );
  CLKINVX1 U5018 ( .A(n5192), .Y(n4595) );
  NAND2BX1 U5019 ( .AN(n5190), .B(n5191), .Y(n6129) );
  CLKINVX1 U5020 ( .A(n6996), .Y(n6620) );
  NAND2X1 U5021 ( .A(n7948), .B(n7947), .Y(n7951) );
  AND2X2 U5022 ( .A(n2824), .B(n4912), .Y(n2805) );
  CLKINVX1 U5023 ( .A(n6831), .Y(n5551) );
  NAND2X1 U5024 ( .A(n8349), .B(n8350), .Y(n7872) );
  CLKINVX1 U5025 ( .A(n4824), .Y(n5673) );
  CLKINVX1 U5026 ( .A(n6546), .Y(n5617) );
  AND2X2 U5027 ( .A(n8207), .B(n7910), .Y(n2807) );
  CLKINVX1 U5028 ( .A(n6464), .Y(n6407) );
  CLKINVX1 U5029 ( .A(n6685), .Y(n6341) );
  AO22X1 U5030 ( .A0(n6337), .A1(n5611), .B0(n5610), .B1(n5609), .Y(n5613) );
  CLKINVX1 U5031 ( .A(n5186), .Y(n4685) );
  CLKBUFX3 U5032 ( .A(n3309), .Y(n3279) );
  CLKBUFX3 U5033 ( .A(n3394), .Y(n3367) );
  CLKBUFX3 U5034 ( .A(n3309), .Y(n3280) );
  CLKBUFX3 U5035 ( .A(n3285), .Y(n3275) );
  CLKBUFX3 U5036 ( .A(n3395), .Y(n3363) );
  CLKBUFX3 U5037 ( .A(n3485), .Y(n3455) );
  CLKBUFX3 U5038 ( .A(n3484), .Y(n3456) );
  CLKBUFX3 U5039 ( .A(n3394), .Y(n3365) );
  CLKBUFX3 U5040 ( .A(n3307), .Y(n3284) );
  CLKBUFX3 U5041 ( .A(n3393), .Y(n3371) );
  CLKBUFX3 U5042 ( .A(n3307), .Y(n3283) );
  CLKBUFX3 U5043 ( .A(n3393), .Y(n3370) );
  CLKBUFX3 U5044 ( .A(n3307), .Y(n3282) );
  CLKBUFX3 U5045 ( .A(n3393), .Y(n3369) );
  CLKBUFX3 U5046 ( .A(n3307), .Y(n3281) );
  CLKBUFX3 U5047 ( .A(n3393), .Y(n3368) );
  CLKBUFX3 U5048 ( .A(n3484), .Y(n3457) );
  CLKBUFX3 U5049 ( .A(n3309), .Y(n3278) );
  CLKBUFX3 U5050 ( .A(n3394), .Y(n3366) );
  CLKBUFX3 U5051 ( .A(n3484), .Y(n3458) );
  CLKBUFX3 U5052 ( .A(n3484), .Y(n3459) );
  CLKBUFX3 U5053 ( .A(n3529), .Y(n3501) );
  CLKBUFX3 U5054 ( .A(n3262), .Y(n3230) );
  CLKBUFX3 U5055 ( .A(n3529), .Y(n3499) );
  CLKBUFX3 U5056 ( .A(n3260), .Y(n3236) );
  CLKBUFX3 U5057 ( .A(n3528), .Y(n3505) );
  CLKBUFX3 U5058 ( .A(n3437), .Y(n3414) );
  CLKBUFX3 U5059 ( .A(n3260), .Y(n3235) );
  CLKBUFX3 U5060 ( .A(n3528), .Y(n3504) );
  CLKBUFX3 U5061 ( .A(n3260), .Y(n3234) );
  CLKBUFX3 U5062 ( .A(n3528), .Y(n3503) );
  CLKBUFX3 U5063 ( .A(n3260), .Y(n3233) );
  CLKBUFX3 U5064 ( .A(n3528), .Y(n3502) );
  CLKBUFX3 U5065 ( .A(n3261), .Y(n3232) );
  CLKBUFX3 U5066 ( .A(n3529), .Y(n3500) );
  CLKBUFX3 U5067 ( .A(n3438), .Y(n3411) );
  CLKBUFX3 U5068 ( .A(n3438), .Y(n3412) );
  CLKBUFX3 U5069 ( .A(n2156), .Y(n3374) );
  CLKBUFX3 U5070 ( .A(n3481), .Y(n3472) );
  CLKBUFX3 U5071 ( .A(n3392), .Y(n3375) );
  CLKBUFX3 U5072 ( .A(n3306), .Y(n3287) );
  CLKBUFX3 U5073 ( .A(n3305), .Y(n3290) );
  CLKBUFX3 U5074 ( .A(n3392), .Y(n3377) );
  CLKBUFX3 U5075 ( .A(n3392), .Y(n3376) );
  CLKBUFX3 U5076 ( .A(n3304), .Y(n3291) );
  CLKBUFX3 U5077 ( .A(n3391), .Y(n3378) );
  CLKBUFX3 U5078 ( .A(n3303), .Y(n3295) );
  CLKBUFX3 U5079 ( .A(n3390), .Y(n3382) );
  CLKBUFX3 U5080 ( .A(n3303), .Y(n3294) );
  CLKBUFX3 U5081 ( .A(n3390), .Y(n3381) );
  CLKBUFX3 U5082 ( .A(n3441), .Y(n3415) );
  CLKBUFX3 U5083 ( .A(n3264), .Y(n3239) );
  CLKBUFX3 U5084 ( .A(n3530), .Y(n3508) );
  CLKBUFX3 U5085 ( .A(n3434), .Y(n3425) );
  CLKBUFX3 U5086 ( .A(n3527), .Y(n3509) );
  CLKBUFX3 U5087 ( .A(n3436), .Y(n3416) );
  CLKBUFX3 U5088 ( .A(n3255), .Y(n3240) );
  CLKBUFX3 U5089 ( .A(n3436), .Y(n3421) );
  CLKBUFX3 U5090 ( .A(n3258), .Y(n3243) );
  CLKBUFX3 U5091 ( .A(n3527), .Y(n3512) );
  CLKBUFX3 U5092 ( .A(n3436), .Y(n3420) );
  CLKBUFX3 U5093 ( .A(n3258), .Y(n3242) );
  CLKBUFX3 U5094 ( .A(n3527), .Y(n3511) );
  CLKBUFX3 U5095 ( .A(n3435), .Y(n3422) );
  CLKBUFX3 U5096 ( .A(n3434), .Y(n3426) );
  CLKBUFX3 U5097 ( .A(n3256), .Y(n3248) );
  CLKBUFX3 U5098 ( .A(n3256), .Y(n3247) );
  CLKBUFX3 U5099 ( .A(n3525), .Y(n3516) );
  CLKBUFX3 U5100 ( .A(n3972), .Y(n3957) );
  AO22X1 U5101 ( .A0(n2821), .A1(n3101), .B0(n3111), .B1(n6536), .Y(n6539) );
  AO22X1 U5102 ( .A0(n6912), .A1(n3100), .B0(n3111), .B1(n6911), .Y(n6916) );
  INVX3 U5103 ( .A(n2863), .Y(n3082) );
  CLKBUFX3 U5104 ( .A(n3657), .Y(n3658) );
  CLKBUFX3 U5105 ( .A(n3648), .Y(n3649) );
  CLKINVX1 U5106 ( .A(n8687), .Y(n8713) );
  CLKBUFX3 U5107 ( .A(n3682), .Y(n3683) );
  CLKINVX1 U5108 ( .A(n6268), .Y(n5908) );
  CLKINVX1 U5109 ( .A(n8683), .Y(n8427) );
  CLKINVX1 U5110 ( .A(n5319), .Y(n6272) );
  CLKBUFX3 U5111 ( .A(n8735), .Y(n3016) );
  CLKBUFX3 U5112 ( .A(n3973), .Y(n3955) );
  CLKBUFX3 U5113 ( .A(n3483), .Y(n3464) );
  CLKBUFX3 U5114 ( .A(n3483), .Y(n3468) );
  CLKBUFX3 U5115 ( .A(n3483), .Y(n3467) );
  CLKBUFX3 U5116 ( .A(n3305), .Y(n3289) );
  CLKBUFX3 U5117 ( .A(n3304), .Y(n3292) );
  CLKBUFX3 U5118 ( .A(n3391), .Y(n3379) );
  CLKBUFX3 U5119 ( .A(n3480), .Y(n3478) );
  CLKBUFX3 U5120 ( .A(n3302), .Y(n3300) );
  CLKBUFX3 U5121 ( .A(n3389), .Y(n3387) );
  CLKBUFX3 U5122 ( .A(n3480), .Y(n3477) );
  CLKBUFX3 U5123 ( .A(n3302), .Y(n3299) );
  CLKBUFX3 U5124 ( .A(n3389), .Y(n3386) );
  CLKBUFX3 U5125 ( .A(n3480), .Y(n3476) );
  CLKBUFX3 U5126 ( .A(n3302), .Y(n3298) );
  CLKBUFX3 U5127 ( .A(n3389), .Y(n3385) );
  CLKBUFX3 U5128 ( .A(n3303), .Y(n3297) );
  CLKBUFX3 U5129 ( .A(n3390), .Y(n3384) );
  CLKBUFX3 U5130 ( .A(n3303), .Y(n3296) );
  CLKBUFX3 U5131 ( .A(n3390), .Y(n3383) );
  CLKBUFX3 U5132 ( .A(n3304), .Y(n3293) );
  CLKBUFX3 U5133 ( .A(n3391), .Y(n3380) );
  CLKBUFX3 U5134 ( .A(n3527), .Y(n3510) );
  CLKBUFX3 U5135 ( .A(n3435), .Y(n3423) );
  CLKBUFX3 U5136 ( .A(n3433), .Y(n3431) );
  CLKBUFX3 U5137 ( .A(n3255), .Y(n3253) );
  CLKBUFX3 U5138 ( .A(n3524), .Y(n3522) );
  CLKBUFX3 U5139 ( .A(n3433), .Y(n3430) );
  CLKBUFX3 U5140 ( .A(n3524), .Y(n3521) );
  CLKBUFX3 U5141 ( .A(n3255), .Y(n3252) );
  CLKBUFX3 U5142 ( .A(n3433), .Y(n3429) );
  CLKBUFX3 U5143 ( .A(n3255), .Y(n3251) );
  CLKBUFX3 U5144 ( .A(n3524), .Y(n3520) );
  CLKBUFX3 U5145 ( .A(n3434), .Y(n3428) );
  CLKBUFX3 U5146 ( .A(n3256), .Y(n3250) );
  CLKBUFX3 U5147 ( .A(n3434), .Y(n3427) );
  CLKBUFX3 U5148 ( .A(n3256), .Y(n3249) );
  CLKBUFX3 U5149 ( .A(n3435), .Y(n3424) );
  CLKINVX1 U5150 ( .A(n8337), .Y(n8339) );
  CLKBUFX3 U5151 ( .A(n2792), .Y(n3174) );
  CLKBUFX3 U5152 ( .A(n2792), .Y(n3175) );
  CLKBUFX3 U5153 ( .A(n2792), .Y(n3173) );
  CLKBUFX3 U5154 ( .A(n2791), .Y(n3123) );
  CLKBUFX3 U5155 ( .A(n2791), .Y(n3122) );
  CLKBUFX3 U5156 ( .A(n2791), .Y(n3124) );
  CLKBUFX3 U5157 ( .A(n2790), .Y(n3119) );
  CLKBUFX3 U5158 ( .A(n2790), .Y(n3120) );
  CLKBUFX3 U5159 ( .A(n3480), .Y(n3479) );
  CLKBUFX3 U5160 ( .A(n3302), .Y(n3301) );
  CLKBUFX3 U5161 ( .A(n3389), .Y(n3388) );
  CLKINVX1 U5162 ( .A(n6206), .Y(n6209) );
  CLKBUFX3 U5163 ( .A(n3433), .Y(n3432) );
  CLKBUFX3 U5164 ( .A(n3255), .Y(n3254) );
  CLKBUFX3 U5165 ( .A(n3524), .Y(n3523) );
  CLKBUFX3 U5166 ( .A(n2773), .Y(n3168) );
  CLKBUFX3 U5167 ( .A(n2784), .Y(n3183) );
  CLKBUFX3 U5168 ( .A(n2785), .Y(n3177) );
  CLKBUFX3 U5169 ( .A(n2782), .Y(n3115) );
  CLKBUFX3 U5170 ( .A(n2782), .Y(n3113) );
  CLKBUFX3 U5171 ( .A(n2773), .Y(n3169) );
  CLKBUFX3 U5172 ( .A(n2784), .Y(n3184) );
  CLKBUFX3 U5173 ( .A(n2785), .Y(n3178) );
  CLKBUFX3 U5174 ( .A(n2788), .Y(n3133) );
  CLKBUFX3 U5175 ( .A(n2773), .Y(n3167) );
  CLKBUFX3 U5176 ( .A(n2782), .Y(n3114) );
  CLKBUFX3 U5177 ( .A(n2784), .Y(n3182) );
  CLKBUFX3 U5178 ( .A(n2785), .Y(n3176) );
  CLKBUFX3 U5179 ( .A(n2787), .Y(n3126) );
  CLKBUFX3 U5180 ( .A(n2788), .Y(n3131) );
  CLKBUFX3 U5181 ( .A(n2787), .Y(n3125) );
  CLKBUFX3 U5182 ( .A(n2788), .Y(n3132) );
  CLKBUFX3 U5183 ( .A(n2787), .Y(n3127) );
  CLKBUFX3 U5184 ( .A(n2776), .Y(n3116) );
  CLKBUFX3 U5185 ( .A(n2777), .Y(n3170) );
  CLKBUFX3 U5186 ( .A(n2777), .Y(n3172) );
  CLKBUFX3 U5187 ( .A(n2776), .Y(n3117) );
  CLKBUFX3 U5188 ( .A(n2786), .Y(n3179) );
  CLKBUFX3 U5189 ( .A(n2789), .Y(n3130) );
  CLKBUFX3 U5190 ( .A(n2777), .Y(n3171) );
  CLKBUFX3 U5191 ( .A(n2786), .Y(n3180) );
  CLKBUFX3 U5192 ( .A(n2789), .Y(n3129) );
  CLKBUFX3 U5193 ( .A(n2789), .Y(n3128) );
  CLKBUFX3 U5194 ( .A(n8715), .Y(n3634) );
  CLKINVX1 U5195 ( .A(n6989), .Y(n6991) );
  CLKBUFX3 U5196 ( .A(n186), .Y(n3159) );
  CLKBUFX3 U5197 ( .A(n191), .Y(n3211) );
  CLKBUFX3 U5198 ( .A(n190), .Y(n3205) );
  CLKBUFX3 U5199 ( .A(n189), .Y(n3198) );
  CLKBUFX3 U5200 ( .A(n188), .Y(n3192) );
  CLKBUFX3 U5201 ( .A(n186), .Y(n3160) );
  CLKBUFX3 U5202 ( .A(n183), .Y(n3153) );
  CLKBUFX3 U5203 ( .A(n185), .Y(n3147) );
  CLKBUFX3 U5204 ( .A(n181), .Y(n3141) );
  CLKBUFX3 U5205 ( .A(n189), .Y(n3200) );
  CLKBUFX3 U5206 ( .A(n188), .Y(n3194) );
  CLKBUFX3 U5207 ( .A(n191), .Y(n3213) );
  CLKBUFX3 U5208 ( .A(n191), .Y(n3212) );
  CLKBUFX3 U5209 ( .A(n190), .Y(n3206) );
  CLKBUFX3 U5210 ( .A(n189), .Y(n3199) );
  CLKBUFX3 U5211 ( .A(n188), .Y(n3193) );
  CLKBUFX3 U5212 ( .A(n190), .Y(n3204) );
  CLKBUFX3 U5213 ( .A(n186), .Y(n3161) );
  CLKBUFX3 U5214 ( .A(n183), .Y(n3154) );
  CLKBUFX3 U5215 ( .A(n185), .Y(n3148) );
  CLKBUFX3 U5216 ( .A(n181), .Y(n3142) );
  CLKBUFX3 U5217 ( .A(n183), .Y(n3152) );
  CLKBUFX3 U5218 ( .A(n185), .Y(n3146) );
  CLKBUFX3 U5219 ( .A(n181), .Y(n3140) );
  CLKBUFX3 U5220 ( .A(n2775), .Y(n3207) );
  CLKBUFX3 U5221 ( .A(n2775), .Y(n3208) );
  CLKBUFX3 U5222 ( .A(n179), .Y(n3201) );
  CLKBUFX3 U5223 ( .A(n187), .Y(n3188) );
  CLKBUFX3 U5224 ( .A(n2774), .Y(n3155) );
  CLKBUFX3 U5225 ( .A(n182), .Y(n3149) );
  CLKBUFX3 U5226 ( .A(n184), .Y(n3143) );
  CLKBUFX3 U5227 ( .A(n180), .Y(n3137) );
  CLKBUFX3 U5228 ( .A(n179), .Y(n3203) );
  CLKBUFX3 U5229 ( .A(n192), .Y(n3196) );
  CLKBUFX3 U5230 ( .A(n187), .Y(n3190) );
  CLKBUFX3 U5231 ( .A(n3208), .Y(n3210) );
  CLKBUFX3 U5232 ( .A(n3208), .Y(n3209) );
  CLKBUFX3 U5233 ( .A(n3157), .Y(n3156) );
  CLKBUFX3 U5234 ( .A(n192), .Y(n3197) );
  CLKBUFX3 U5235 ( .A(n3188), .Y(n3191) );
  CLKBUFX3 U5236 ( .A(n179), .Y(n3202) );
  CLKBUFX3 U5237 ( .A(n192), .Y(n3195) );
  CLKBUFX3 U5238 ( .A(n3188), .Y(n3189) );
  CLKBUFX3 U5239 ( .A(n3157), .Y(n3158) );
  CLKBUFX3 U5240 ( .A(n182), .Y(n3151) );
  CLKBUFX3 U5241 ( .A(n184), .Y(n3145) );
  CLKBUFX3 U5242 ( .A(n180), .Y(n3139) );
  CLKBUFX3 U5243 ( .A(n8452), .Y(n3601) );
  CLKBUFX3 U5244 ( .A(n8452), .Y(n3600) );
  NAND2X1 U5245 ( .A(n3585), .B(n3688), .Y(n8333) );
  CLKBUFX3 U5246 ( .A(n3976), .Y(n3956) );
  CLKBUFX3 U5247 ( .A(n3483), .Y(n3466) );
  CLKBUFX3 U5248 ( .A(n3305), .Y(n3288) );
  CLKBUFX3 U5249 ( .A(n3466), .Y(n3465) );
  CLKBUFX3 U5250 ( .A(n3436), .Y(n3419) );
  CLKBUFX3 U5251 ( .A(n3436), .Y(n3418) );
  CLKBUFX3 U5252 ( .A(n3418), .Y(n3417) );
  CLKBUFX3 U5253 ( .A(n3259), .Y(n3241) );
  CLKBUFX3 U5254 ( .A(n3971), .Y(n3958) );
  CLKBUFX3 U5255 ( .A(n3971), .Y(n3959) );
  CLKBUFX3 U5256 ( .A(n3971), .Y(n3960) );
  CLKBUFX3 U5257 ( .A(n3971), .Y(n3961) );
  CLKBUFX3 U5258 ( .A(n3971), .Y(n3962) );
  CLKBUFX3 U5259 ( .A(n3970), .Y(n3963) );
  CLKBUFX3 U5260 ( .A(n3970), .Y(n3964) );
  CLKBUFX3 U5261 ( .A(n3970), .Y(n3965) );
  CLKBUFX3 U5262 ( .A(n3976), .Y(n3966) );
  CLKBUFX3 U5263 ( .A(n3976), .Y(n3967) );
  CLKBUFX3 U5264 ( .A(n3970), .Y(n3968) );
  CLKBUFX3 U5265 ( .A(n3970), .Y(n3969) );
  CLKBUFX3 U5266 ( .A(n8453), .Y(n3603) );
  CLKBUFX3 U5267 ( .A(n8453), .Y(n3602) );
  CLKBUFX3 U5268 ( .A(n44), .Y(n3761) );
  CLKBUFX3 U5269 ( .A(n43), .Y(n3758) );
  CLKBUFX3 U5270 ( .A(n42), .Y(n3755) );
  CLKBUFX3 U5271 ( .A(n41), .Y(n3752) );
  CLKBUFX3 U5272 ( .A(n40), .Y(n3749) );
  CLKBUFX3 U5273 ( .A(n39), .Y(n3746) );
  CLKBUFX3 U5274 ( .A(n38), .Y(n3743) );
  CLKBUFX3 U5275 ( .A(n37), .Y(n3740) );
  CLKBUFX3 U5276 ( .A(n36), .Y(n3737) );
  CLKBUFX3 U5277 ( .A(n35), .Y(n3734) );
  CLKBUFX3 U5278 ( .A(n34), .Y(n3731) );
  CLKBUFX3 U5279 ( .A(n33), .Y(n3728) );
  CLKBUFX3 U5280 ( .A(n32), .Y(n3725) );
  CLKBUFX3 U5281 ( .A(n31), .Y(n3722) );
  CLKBUFX3 U5282 ( .A(n30), .Y(n3719) );
  CLKBUFX3 U5283 ( .A(n29), .Y(n3716) );
  CLKBUFX3 U5284 ( .A(n28), .Y(n3713) );
  CLKBUFX3 U5285 ( .A(\i_MIPS/Register/n118 ), .Y(n3710) );
  CLKBUFX3 U5286 ( .A(\i_MIPS/Register/n116 ), .Y(n3707) );
  CLKBUFX3 U5287 ( .A(\i_MIPS/Register/n114 ), .Y(n3704) );
  CLKBUFX3 U5288 ( .A(\i_MIPS/Register/n112 ), .Y(n3701) );
  CLKBUFX3 U5289 ( .A(\i_MIPS/Register/n110 ), .Y(n3698) );
  CLKBUFX3 U5290 ( .A(\i_MIPS/Register/n108 ), .Y(n3695) );
  CLKBUFX3 U5291 ( .A(\i_MIPS/Register/n106 ), .Y(n3692) );
  CLKBUFX3 U5292 ( .A(n44), .Y(n3759) );
  CLKBUFX3 U5293 ( .A(n44), .Y(n3760) );
  CLKBUFX3 U5294 ( .A(n43), .Y(n3756) );
  CLKBUFX3 U5295 ( .A(n43), .Y(n3757) );
  CLKBUFX3 U5296 ( .A(n42), .Y(n3753) );
  CLKBUFX3 U5297 ( .A(n42), .Y(n3754) );
  CLKBUFX3 U5298 ( .A(n41), .Y(n3750) );
  CLKBUFX3 U5299 ( .A(n41), .Y(n3751) );
  CLKBUFX3 U5300 ( .A(n40), .Y(n3747) );
  CLKBUFX3 U5301 ( .A(n40), .Y(n3748) );
  CLKBUFX3 U5302 ( .A(n39), .Y(n3744) );
  CLKBUFX3 U5303 ( .A(n39), .Y(n3745) );
  CLKBUFX3 U5304 ( .A(n38), .Y(n3741) );
  CLKBUFX3 U5305 ( .A(n38), .Y(n3742) );
  CLKBUFX3 U5306 ( .A(n37), .Y(n3738) );
  CLKBUFX3 U5307 ( .A(n37), .Y(n3739) );
  CLKBUFX3 U5308 ( .A(n36), .Y(n3735) );
  CLKBUFX3 U5309 ( .A(n36), .Y(n3736) );
  CLKBUFX3 U5310 ( .A(n35), .Y(n3732) );
  CLKBUFX3 U5311 ( .A(n35), .Y(n3733) );
  CLKBUFX3 U5312 ( .A(n34), .Y(n3729) );
  CLKBUFX3 U5313 ( .A(n34), .Y(n3730) );
  CLKBUFX3 U5314 ( .A(n33), .Y(n3726) );
  CLKBUFX3 U5315 ( .A(n33), .Y(n3727) );
  CLKBUFX3 U5316 ( .A(n32), .Y(n3723) );
  CLKBUFX3 U5317 ( .A(n32), .Y(n3724) );
  CLKBUFX3 U5318 ( .A(n31), .Y(n3720) );
  CLKBUFX3 U5319 ( .A(n31), .Y(n3721) );
  CLKBUFX3 U5320 ( .A(n30), .Y(n3717) );
  CLKBUFX3 U5321 ( .A(n30), .Y(n3718) );
  CLKBUFX3 U5322 ( .A(n29), .Y(n3714) );
  CLKBUFX3 U5323 ( .A(n29), .Y(n3715) );
  CLKBUFX3 U5324 ( .A(n28), .Y(n3711) );
  CLKBUFX3 U5325 ( .A(n28), .Y(n3712) );
  CLKBUFX3 U5326 ( .A(\i_MIPS/Register/n118 ), .Y(n3708) );
  CLKBUFX3 U5327 ( .A(\i_MIPS/Register/n118 ), .Y(n3709) );
  CLKBUFX3 U5328 ( .A(\i_MIPS/Register/n116 ), .Y(n3705) );
  CLKBUFX3 U5329 ( .A(\i_MIPS/Register/n116 ), .Y(n3706) );
  CLKBUFX3 U5330 ( .A(\i_MIPS/Register/n114 ), .Y(n3702) );
  CLKBUFX3 U5331 ( .A(\i_MIPS/Register/n114 ), .Y(n3703) );
  CLKBUFX3 U5332 ( .A(\i_MIPS/Register/n112 ), .Y(n3699) );
  CLKBUFX3 U5333 ( .A(\i_MIPS/Register/n112 ), .Y(n3700) );
  CLKBUFX3 U5334 ( .A(\i_MIPS/Register/n110 ), .Y(n3696) );
  CLKBUFX3 U5335 ( .A(\i_MIPS/Register/n110 ), .Y(n3697) );
  CLKBUFX3 U5336 ( .A(\i_MIPS/Register/n108 ), .Y(n3693) );
  CLKBUFX3 U5337 ( .A(\i_MIPS/Register/n108 ), .Y(n3694) );
  CLKBUFX3 U5338 ( .A(\i_MIPS/Register/n106 ), .Y(n3690) );
  CLKBUFX3 U5339 ( .A(\i_MIPS/Register/n106 ), .Y(n3691) );
  CLKBUFX3 U5340 ( .A(n51), .Y(n3782) );
  CLKBUFX3 U5341 ( .A(n50), .Y(n3779) );
  CLKBUFX3 U5342 ( .A(n49), .Y(n3776) );
  CLKBUFX3 U5343 ( .A(n48), .Y(n3773) );
  CLKBUFX3 U5344 ( .A(n47), .Y(n3770) );
  CLKBUFX3 U5345 ( .A(n46), .Y(n3767) );
  CLKBUFX3 U5346 ( .A(n45), .Y(n3764) );
  CLKBUFX3 U5347 ( .A(n51), .Y(n3781) );
  CLKBUFX3 U5348 ( .A(n50), .Y(n3778) );
  CLKBUFX3 U5349 ( .A(n49), .Y(n3775) );
  CLKBUFX3 U5350 ( .A(n48), .Y(n3772) );
  CLKBUFX3 U5351 ( .A(n47), .Y(n3769) );
  CLKBUFX3 U5352 ( .A(n46), .Y(n3766) );
  CLKBUFX3 U5353 ( .A(n45), .Y(n3763) );
  CLKBUFX3 U5354 ( .A(n51), .Y(n3780) );
  CLKBUFX3 U5355 ( .A(n50), .Y(n3777) );
  CLKBUFX3 U5356 ( .A(n49), .Y(n3774) );
  CLKBUFX3 U5357 ( .A(n48), .Y(n3771) );
  CLKBUFX3 U5358 ( .A(n47), .Y(n3768) );
  CLKBUFX3 U5359 ( .A(n46), .Y(n3765) );
  CLKBUFX3 U5360 ( .A(n45), .Y(n3762) );
  INVX3 U5361 ( .A(n2883), .Y(n3688) );
  INVX3 U5362 ( .A(n2883), .Y(n3689) );
  CLKBUFX3 U5363 ( .A(\D_cache/n211 ), .Y(n3883) );
  CLKBUFX3 U5364 ( .A(\D_cache/n207 ), .Y(n3803) );
  CLKBUFX3 U5365 ( .A(\D_cache/n209 ), .Y(n3843) );
  CLKBUFX3 U5366 ( .A(\D_cache/n208 ), .Y(n3823) );
  CLKBUFX3 U5367 ( .A(\D_cache/n212 ), .Y(n3903) );
  CLKBUFX3 U5368 ( .A(\D_cache/n213 ), .Y(n3924) );
  CLKBUFX3 U5369 ( .A(\D_cache/n210 ), .Y(n3863) );
  CLKBUFX3 U5370 ( .A(n4384), .Y(n4072) );
  CLKBUFX3 U5371 ( .A(n4384), .Y(n4071) );
  CLKBUFX3 U5372 ( .A(n4384), .Y(n4070) );
  CLKBUFX3 U5373 ( .A(n4384), .Y(n4069) );
  CLKBUFX3 U5374 ( .A(n4384), .Y(n4065) );
  CLKBUFX3 U5375 ( .A(n4384), .Y(n4064) );
  CLKBUFX3 U5376 ( .A(n4384), .Y(n4063) );
  CLKBUFX3 U5377 ( .A(n4384), .Y(n4061) );
  CLKBUFX3 U5378 ( .A(n4385), .Y(n4060) );
  CLKBUFX3 U5379 ( .A(n4385), .Y(n4059) );
  CLKBUFX3 U5380 ( .A(n4385), .Y(n4058) );
  CLKBUFX3 U5381 ( .A(n4385), .Y(n4057) );
  CLKBUFX3 U5382 ( .A(n4385), .Y(n4056) );
  CLKBUFX3 U5383 ( .A(n4385), .Y(n4055) );
  CLKBUFX3 U5384 ( .A(n4385), .Y(n4050) );
  CLKBUFX3 U5385 ( .A(n4385), .Y(n4049) );
  CLKBUFX3 U5386 ( .A(n4386), .Y(n4048) );
  CLKBUFX3 U5387 ( .A(n4386), .Y(n4046) );
  CLKBUFX3 U5388 ( .A(rst_n), .Y(n4045) );
  CLKBUFX3 U5389 ( .A(n4386), .Y(n4044) );
  CLKBUFX3 U5390 ( .A(n4386), .Y(n4043) );
  CLKBUFX3 U5391 ( .A(n4372), .Y(n4042) );
  CLKBUFX3 U5392 ( .A(n4384), .Y(n4066) );
  CLKBUFX3 U5393 ( .A(n4360), .Y(n4047) );
  CLKBUFX3 U5394 ( .A(n4384), .Y(n4062) );
  CLKBUFX3 U5395 ( .A(n4385), .Y(n4052) );
  CLKBUFX3 U5396 ( .A(n4385), .Y(n4051) );
  CLKBUFX3 U5397 ( .A(n4384), .Y(n4068) );
  CLKBUFX3 U5398 ( .A(n4384), .Y(n4067) );
  CLKBUFX3 U5399 ( .A(n4385), .Y(n4053) );
  CLKBUFX3 U5400 ( .A(n4385), .Y(n4054) );
  CLKBUFX3 U5401 ( .A(n4386), .Y(n4361) );
  CLKBUFX3 U5402 ( .A(n4367), .Y(n4362) );
  CLKBUFX3 U5403 ( .A(rst_n), .Y(n4363) );
  CLKBUFX3 U5404 ( .A(n4372), .Y(n4364) );
  CLKBUFX3 U5405 ( .A(n4376), .Y(n4365) );
  CLKBUFX3 U5406 ( .A(n4364), .Y(n4366) );
  CLKBUFX3 U5407 ( .A(n4369), .Y(n4367) );
  CLKBUFX3 U5408 ( .A(n4386), .Y(n4378) );
  CLKBUFX3 U5409 ( .A(n4365), .Y(n4379) );
  CLKBUFX3 U5410 ( .A(n4386), .Y(n4380) );
  CLKBUFX3 U5411 ( .A(n4386), .Y(n4381) );
  CLKBUFX3 U5412 ( .A(n4368), .Y(n4382) );
  CLKBUFX3 U5413 ( .A(n4386), .Y(n4383) );
  CLKBUFX3 U5414 ( .A(n4386), .Y(n4368) );
  CLKBUFX3 U5415 ( .A(rst_n), .Y(n4369) );
  CLKBUFX3 U5416 ( .A(n4377), .Y(n4370) );
  CLKBUFX3 U5417 ( .A(n4375), .Y(n4371) );
  CLKBUFX3 U5418 ( .A(rst_n), .Y(n4372) );
  CLKBUFX3 U5419 ( .A(n4363), .Y(n4373) );
  CLKBUFX3 U5420 ( .A(n4386), .Y(n4374) );
  CLKBUFX3 U5421 ( .A(rst_n), .Y(n4375) );
  CLKBUFX3 U5422 ( .A(rst_n), .Y(n4376) );
  CLKBUFX3 U5423 ( .A(n4369), .Y(n4377) );
  CLKBUFX3 U5424 ( .A(n3661), .Y(n3025) );
  CLKBUFX3 U5425 ( .A(n3650), .Y(n3651) );
  CLKBUFX3 U5426 ( .A(n3680), .Y(n3681) );
  CLKINVX1 U5427 ( .A(n5613), .Y(n5615) );
  XNOR2X4 U5428 ( .A(n7661), .B(n25), .Y(n7787) );
  OAI221XL U5429 ( .A0(n3106), .A1(n6190), .B0(n6130), .B1(n3098), .C0(n3097), 
        .Y(n6133) );
  OAI221XL U5430 ( .A0(n3106), .A1(n5389), .B0(n2851), .B1(n3098), .C0(n3097), 
        .Y(n5393) );
  OAI221XL U5431 ( .A0(n3107), .A1(n4973), .B0(n4904), .B1(n3099), .C0(n3097), 
        .Y(n4907) );
  CLKINVX1 U5432 ( .A(n6462), .Y(n6465) );
  CLKMX2X2 U5433 ( .A(n7005), .B(n3071), .S0(n5957), .Y(n6000) );
  AOI222XL U5434 ( .A0(n2877), .A1(n6680), .B0(n5968), .B1(n7006), .C0(n5967), 
        .C1(n6990), .Y(n5998) );
  NAND2X1 U5435 ( .A(n6614), .B(n5970), .Y(n5548) );
  OAI221XL U5436 ( .A0(n5904), .A1(n5331), .B0(n5902), .B1(n6824), .C0(n4817), 
        .Y(n4845) );
  AOI222XL U5437 ( .A0(n4841), .A1(n6993), .B0(n2805), .B1(n6267), .C0(n6476), 
        .C1(n5973), .Y(n4842) );
  AOI222XL U5438 ( .A0(n6683), .A1(n6682), .B0(n6681), .B1(n6990), .C0(n6680), 
        .C1(n6679), .Y(n6702) );
  CLKMX2X2 U5439 ( .A(n7005), .B(n3071), .S0(n6904), .Y(n6928) );
  CLKMX2X2 U5440 ( .A(n7005), .B(n3071), .S0(n6622), .Y(n6623) );
  AOI222X1 U5441 ( .A0(n6620), .A1(n6619), .B0(n2817), .B1(n6618), .C0(n6617), 
        .C1(n6616), .Y(n6624) );
  CLKINVX1 U5442 ( .A(n4592), .Y(n4594) );
  NAND2X1 U5443 ( .A(n8221), .B(n8211), .Y(n7947) );
  NAND2X1 U5444 ( .A(n8543), .B(n8548), .Y(n5978) );
  NAND2X1 U5445 ( .A(n5971), .B(n5970), .Y(n6137) );
  CLKINVX1 U5446 ( .A(n8275), .Y(n8282) );
  AND2X2 U5447 ( .A(n6614), .B(n5480), .Y(n2809) );
  NAND2X1 U5448 ( .A(n7986), .B(n7985), .Y(n8021) );
  AOI2BB1X1 U5449 ( .A0N(n2855), .A1N(n2814), .B0(n8351), .Y(n8353) );
  CLKINVX1 U5450 ( .A(n8350), .Y(n8351) );
  AOI2BB1X1 U5451 ( .A0N(n2857), .A1N(n2827), .B0(n7884), .Y(n7885) );
  CLKINVX1 U5452 ( .A(n7894), .Y(n7884) );
  AOI2BB1X1 U5453 ( .A0N(n2858), .A1N(n7935), .B0(n7934), .Y(n7936) );
  CLKINVX1 U5454 ( .A(n7948), .Y(n7934) );
  CLKINVX1 U5455 ( .A(n8022), .Y(n7999) );
  NAND2X1 U5456 ( .A(n7899), .B(n7898), .Y(n7910) );
  NAND2X1 U5457 ( .A(n6690), .B(n6694), .Y(n5984) );
  CLKINVX1 U5458 ( .A(n7979), .Y(n7984) );
  NAND2X1 U5459 ( .A(n7968), .B(n7967), .Y(n7980) );
  NAND2X1 U5460 ( .A(n7956), .B(n7955), .Y(n7981) );
  NAND2X1 U5461 ( .A(n7933), .B(n7932), .Y(n7948) );
  NAND2X1 U5462 ( .A(n7883), .B(n7882), .Y(n7894) );
  NAND2BX1 U5463 ( .AN(n8553), .B(n8682), .Y(n8685) );
  AOI2BB1X1 U5464 ( .A0N(n2854), .A1N(n7853), .B0(n7852), .Y(n7854) );
  CLKINVX1 U5465 ( .A(n7865), .Y(n7852) );
  CLKINVX1 U5466 ( .A(n8207), .Y(n8208) );
  CLKINVX1 U5467 ( .A(n8206), .Y(n8210) );
  AOI2BB1X1 U5468 ( .A0N(n2856), .A1N(n2806), .B0(n7969), .Y(n7970) );
  CLKINVX1 U5469 ( .A(n7980), .Y(n7969) );
  NAND2BX1 U5470 ( .AN(n5979), .B(n2833), .Y(n4603) );
  CLKINVX1 U5471 ( .A(n8464), .Y(n8716) );
  OAI21XL U5472 ( .A0(n8806), .A1(n8919), .B0(n8918), .Y(n8920) );
  OAI21XL U5473 ( .A0(n8912), .A1(n8911), .B0(n8910), .Y(n8921) );
  OAI22XL U5474 ( .A0(n8917), .A1(n8916), .B0(n2833), .B1(n8917), .Y(n8918) );
  NAND2X1 U5475 ( .A(n4893), .B(n5970), .Y(n6677) );
  CLKMX2X2 U5476 ( .A(n6333), .B(n6619), .S0(n4016), .Y(n4893) );
  CLKINVX1 U5477 ( .A(n6913), .Y(n6904) );
  AOI21X1 U5478 ( .A0(n8481), .A1(n8482), .B0(n8483), .Y(n8484) );
  CLKINVX1 U5479 ( .A(n5964), .Y(n4983) );
  CLKBUFX2 U5480 ( .A(n8741), .Y(n3679) );
  CLKINVX1 U5481 ( .A(n4833), .Y(n4816) );
  CLKINVX1 U5482 ( .A(n5739), .Y(n5749) );
  CLKINVX1 U5483 ( .A(n8497), .Y(n6602) );
  CLKINVX1 U5484 ( .A(n6834), .Y(n8544) );
  OAI211X1 U5485 ( .A0(n4637), .A1(n4641), .B0(n5990), .C0(n6837), .Y(n4638)
         );
  AO21X1 U5486 ( .A0(n4832), .A1(n4831), .B0(n5755), .Y(n5604) );
  CLKINVX1 U5487 ( .A(n4679), .Y(n4684) );
  CLKINVX1 U5488 ( .A(n8211), .Y(n8217) );
  CLKINVX1 U5489 ( .A(n6678), .Y(n6681) );
  CLKINVX1 U5490 ( .A(n7985), .Y(n7983) );
  CLKINVX1 U5491 ( .A(n7955), .Y(n7945) );
  CLKINVX1 U5492 ( .A(n6394), .Y(n6262) );
  NOR2X4 U5493 ( .A(n5600), .B(n5599), .Y(n5808) );
  NAND2BX1 U5494 ( .AN(n2163), .B(n8652), .Y(n7366) );
  CLKINVX1 U5495 ( .A(n6192), .Y(n6130) );
  NAND2BX1 U5496 ( .AN(n7900), .B(n7910), .Y(n7901) );
  AOI2BB1X1 U5497 ( .A0N(n7897), .A1N(n7911), .B0(n7913), .Y(n7900) );
  CLKINVX1 U5498 ( .A(n6059), .Y(n5475) );
  CLKINVX1 U5499 ( .A(n4970), .Y(n4904) );
  NOR2X4 U5500 ( .A(n6671), .B(n6670), .Y(n6750) );
  NOR2X1 U5501 ( .A(n7921), .B(n7920), .Y(n7935) );
  CLKINVX1 U5502 ( .A(n7947), .Y(n7920) );
  CLKINVX1 U5503 ( .A(n7954), .Y(n7919) );
  AND2X2 U5504 ( .A(n4725), .B(n4728), .Y(n2816) );
  AOI21X1 U5505 ( .A0(n5754), .A1(n6336), .B0(n5753), .Y(n2817) );
  CLKINVX1 U5506 ( .A(n6759), .Y(n5612) );
  CLKINVX1 U5507 ( .A(n5601), .Y(n5603) );
  AND2X2 U5508 ( .A(n4710), .B(n5049), .Y(n2819) );
  CLKINVX1 U5509 ( .A(n8470), .Y(n8474) );
  AND2X2 U5510 ( .A(n6339), .B(n5549), .Y(n2825) );
  NAND2BX1 U5511 ( .AN(n8496), .B(n8497), .Y(n8500) );
  CLKINVX1 U5512 ( .A(n7825), .Y(n7853) );
  NAND2BX1 U5513 ( .AN(n7824), .B(n7864), .Y(n7825) );
  AOI2BB1X1 U5514 ( .A0N(n7873), .A1N(n7872), .B0(n7868), .Y(n7824) );
  CLKINVX1 U5515 ( .A(n8535), .Y(n8536) );
  AO21X1 U5516 ( .A0(n5267), .A1(n6337), .B0(n2874), .Y(n6756) );
  AO21X1 U5517 ( .A0(n5551), .A1(n5970), .B0(n4983), .Y(n6828) );
  AO21X1 U5518 ( .A0(n5899), .A1(n6337), .B0(n2874), .Y(n6270) );
  AO22X1 U5519 ( .A0(n5116), .A1(n5970), .B0(n5115), .B1(n5480), .Y(n5123) );
  CLKINVX1 U5520 ( .A(n8518), .Y(n8519) );
  CLKINVX1 U5521 ( .A(n8514), .Y(n8476) );
  BUFX8 U5522 ( .A(n3581), .Y(n3578) );
  CLKBUFX3 U5523 ( .A(\D_cache/n455 ), .Y(n3997) );
  CLKINVX1 U5524 ( .A(n3071), .Y(n6405) );
  AO22X1 U5525 ( .A0(n4904), .A1(n3100), .B0(n3111), .B1(n4973), .Y(n4906) );
  CLKBUFX3 U5526 ( .A(n2864), .Y(n3079) );
  CLKBUFX3 U5527 ( .A(n2864), .Y(n3080) );
  CLKMX2X2 U5528 ( .A(n3072), .B(n2865), .S0(n5270), .Y(n5271) );
  CLKMX2X2 U5529 ( .A(n3072), .B(n2865), .S0(n6189), .Y(n6139) );
  CLKMX2X2 U5530 ( .A(n3072), .B(n2865), .S0(n5385), .Y(n5332) );
  AO22X1 U5531 ( .A0(n6602), .A1(n3100), .B0(n3110), .B1(n6601), .Y(n6605) );
  CLKMX2X2 U5532 ( .A(n3071), .B(n7005), .S0(n6762), .Y(n6753) );
  CLKINVX1 U5533 ( .A(n5811), .Y(n5812) );
  AO22X1 U5534 ( .A0(n6130), .A1(n3102), .B0(n3108), .B1(n6190), .Y(n6132) );
  AO22X1 U5535 ( .A0(n2820), .A1(n3101), .B0(n3108), .B1(n6193), .Y(n6196) );
  AO22X1 U5536 ( .A0(n2851), .A1(n3103), .B0(n3110), .B1(n5389), .Y(n5392) );
  AO22X1 U5537 ( .A0(n2852), .A1(n3103), .B0(n3109), .B1(n4974), .Y(n4980) );
  INVX3 U5538 ( .A(n2907), .Y(n3087) );
  CLKINVX1 U5539 ( .A(n6547), .Y(n6548) );
  INVX3 U5540 ( .A(n3090), .Y(n3085) );
  CLKINVX1 U5541 ( .A(n8806), .Y(n8913) );
  AO22X1 U5542 ( .A0(n2847), .A1(n3102), .B0(n3109), .B1(n6063), .Y(n6068) );
  AOI222XL U5543 ( .A0(n6205), .A1(n6614), .B0(n2881), .B1(n6204), .C0(n6617), 
        .C1(n6203), .Y(n6211) );
  CLKBUFX3 U5544 ( .A(n3440), .Y(n3437) );
  CLKBUFX3 U5545 ( .A(n3440), .Y(n3439) );
  CLKBUFX3 U5546 ( .A(n3486), .Y(n3485) );
  CLKBUFX3 U5547 ( .A(n3263), .Y(n3262) );
  CLKBUFX3 U5548 ( .A(n3396), .Y(n3395) );
  CLKBUFX3 U5549 ( .A(n3487), .Y(n3481) );
  CLKBUFX3 U5550 ( .A(n3487), .Y(n3482) );
  CLKBUFX3 U5551 ( .A(n3264), .Y(n3257) );
  CLKBUFX3 U5552 ( .A(n3531), .Y(n3526) );
  CLKBUFX3 U5553 ( .A(n3531), .Y(n3525) );
  CLKINVX1 U5554 ( .A(n6984), .Y(n3105) );
  CLKBUFX3 U5555 ( .A(n2767), .Y(n3574) );
  CLKBUFX3 U5556 ( .A(n2767), .Y(n3575) );
  CLKBUFX3 U5557 ( .A(n6983), .Y(n3095) );
  CLKBUFX3 U5558 ( .A(n27), .Y(n3656) );
  CLKBUFX3 U5559 ( .A(n27), .Y(n3655) );
  CLKBUFX3 U5560 ( .A(n3669), .Y(n3670) );
  OA22X2 U5561 ( .A0(n8715), .A1(n8822), .B0(n1625), .B1(n3977), .Y(
        \D_cache/n235 ) );
  OA22X2 U5562 ( .A0(n8715), .A1(n8828), .B0(n1622), .B1(n3977), .Y(
        \D_cache/n241 ) );
  OA22X2 U5563 ( .A0(n8715), .A1(n8830), .B0(n1624), .B1(n3977), .Y(
        \D_cache/n243 ) );
  OA22X2 U5564 ( .A0(n3634), .A1(n8831), .B0(n1623), .B1(n3977), .Y(
        \D_cache/n244 ) );
  OA22X2 U5565 ( .A0(n3634), .A1(n8811), .B0(n1092), .B1(n3978), .Y(
        \D_cache/n223 ) );
  OA22X2 U5566 ( .A0(n3634), .A1(n8814), .B0(n1089), .B1(n3978), .Y(
        \D_cache/n227 ) );
  OA22X2 U5567 ( .A0(n3634), .A1(n8815), .B0(n1090), .B1(n3978), .Y(
        \D_cache/n228 ) );
  OA22X2 U5568 ( .A0(n3634), .A1(n8817), .B0(n1091), .B1(n3978), .Y(
        \D_cache/n230 ) );
  OA22X2 U5569 ( .A0(n3634), .A1(n8818), .B0(n1088), .B1(n3978), .Y(
        \D_cache/n231 ) );
  OA22X2 U5570 ( .A0(n3634), .A1(n8819), .B0(n1087), .B1(n3978), .Y(
        \D_cache/n232 ) );
  OA22X2 U5571 ( .A0(n3634), .A1(n8823), .B0(n1070), .B1(n3977), .Y(
        \D_cache/n236 ) );
  OA22X2 U5572 ( .A0(n3634), .A1(n8825), .B0(n1071), .B1(n3977), .Y(
        \D_cache/n238 ) );
  OA22X2 U5573 ( .A0(n3634), .A1(n8829), .B0(n1626), .B1(n3977), .Y(
        \D_cache/n242 ) );
  OA22X1 U5574 ( .A0(n6334), .A1(n5266), .B0(n6829), .B1(n3069), .Y(n4717) );
  AND2X2 U5575 ( .A(n7798), .B(n7838), .Y(n2829) );
  NAND3BX1 U5576 ( .AN(n7838), .B(n2830), .C(n7837), .Y(n7841) );
  CLKINVX1 U5577 ( .A(n8551), .Y(n8715) );
  CLKBUFX3 U5578 ( .A(n8729), .Y(n3659) );
  CLKINVX1 U5579 ( .A(n7837), .Y(n7827) );
  NAND2X1 U5580 ( .A(n4966), .B(n5970), .Y(n6826) );
  CLKMX2X2 U5581 ( .A(n6330), .B(n6333), .S0(n4016), .Y(n6054) );
  CLKINVX1 U5582 ( .A(n8258), .Y(n8262) );
  NAND2BX1 U5583 ( .AN(n2163), .B(n8676), .Y(n7188) );
  NAND2BX1 U5584 ( .AN(n2163), .B(n8679), .Y(n7260) );
  NAND2BX1 U5585 ( .AN(n2163), .B(n8681), .Y(n7304) );
  NAND2BX1 U5586 ( .AN(n2163), .B(n8680), .Y(n7284) );
  NAND2BX1 U5587 ( .AN(n2163), .B(n8678), .Y(n7236) );
  NAND2BX1 U5588 ( .AN(n2163), .B(n8677), .Y(n7212) );
  CLKINVX1 U5589 ( .A(n6336), .Y(n5204) );
  CLKINVX1 U5590 ( .A(n7636), .Y(n8455) );
  CLKINVX1 U5591 ( .A(n6552), .Y(n6553) );
  CLKINVX1 U5592 ( .A(n5124), .Y(n5111) );
  CLKINVX1 U5593 ( .A(n6694), .Y(n6672) );
  CLKINVX1 U5594 ( .A(n6065), .Y(n6046) );
  CLKBUFX3 U5595 ( .A(n3677), .Y(n3678) );
  CLKBUFX3 U5596 ( .A(\D_cache/n246 ), .Y(n3979) );
  CLKBUFX3 U5597 ( .A(\D_cache/n246 ), .Y(n3980) );
  CLKBUFX3 U5598 ( .A(n3980), .Y(n3981) );
  CLKBUFX3 U5599 ( .A(\D_cache/n246 ), .Y(n3982) );
  CLKBUFX3 U5600 ( .A(\D_cache/n246 ), .Y(n3983) );
  CLKBUFX3 U5601 ( .A(\D_cache/n246 ), .Y(n3984) );
  CLKBUFX3 U5602 ( .A(\D_cache/n246 ), .Y(n3985) );
  CLKBUFX3 U5603 ( .A(\D_cache/n319 ), .Y(n3989) );
  CLKBUFX3 U5604 ( .A(\D_cache/n454 ), .Y(n3995) );
  CLKBUFX3 U5605 ( .A(\D_cache/n250 ), .Y(n3986) );
  CLKBUFX3 U5606 ( .A(\D_cache/n387 ), .Y(n3992) );
  CLKINVX1 U5607 ( .A(n5832), .Y(n5834) );
  CLKINVX1 U5608 ( .A(n6615), .Y(n6616) );
  CLKBUFX3 U5609 ( .A(n7046), .Y(n3162) );
  CLKBUFX3 U5610 ( .A(n3164), .Y(n3166) );
  CLKINVX1 U5611 ( .A(n7000), .Y(n6676) );
  CLKBUFX3 U5612 ( .A(n2786), .Y(n3181) );
  CLKBUFX3 U5613 ( .A(n2776), .Y(n3118) );
  CLKINVX1 U5614 ( .A(n6528), .Y(n6530) );
  NAND2X1 U5615 ( .A(n5970), .B(n1082), .Y(n5965) );
  CLKBUFX3 U5616 ( .A(n5966), .Y(n3068) );
  NAND2X1 U5617 ( .A(n55), .B(n5970), .Y(n5966) );
  NAND2BX1 U5618 ( .AN(n2163), .B(n8674), .Y(n7438) );
  NAND2BX1 U5619 ( .AN(n2163), .B(n8672), .Y(n8137) );
  NAND2BX1 U5620 ( .AN(n2163), .B(n8673), .Y(n7462) );
  CLKINVX1 U5621 ( .A(n7312), .Y(n7308) );
  CLKINVX1 U5622 ( .A(\i_MIPS/Control_ID/n10 ), .Y(n7075) );
  CLKINVX1 U5623 ( .A(n8419), .Y(n8422) );
  CLKINVX1 U5624 ( .A(n8050), .Y(n8052) );
  CLKINVX1 U5625 ( .A(n8031), .Y(n8032) );
  CLKINVX1 U5626 ( .A(n8004), .Y(n8005) );
  CLKINVX1 U5627 ( .A(n8153), .Y(n8154) );
  CLKINVX1 U5628 ( .A(n8094), .Y(n8095) );
  CLKBUFX3 U5629 ( .A(n8334), .Y(n3585) );
  CLKBUFX3 U5630 ( .A(n3976), .Y(n3970) );
  CLKBUFX3 U5631 ( .A(n8334), .Y(n3584) );
  CLKBUFX3 U5632 ( .A(n4386), .Y(n4384) );
  CLKBUFX3 U5633 ( .A(n4386), .Y(n4385) );
  AOI2BB1X1 U5634 ( .A0N(n5900), .A1N(n3092), .B0(n2895), .Y(n5114) );
  OAI221X1 U5635 ( .A0(\i_MIPS/n342 ), .A1(n3091), .B0(n5900), .B1(n3086), 
        .C0(n4895), .Y(n5748) );
  AOI2BB1X1 U5636 ( .A0N(\i_MIPS/n344 ), .A1N(n3092), .B0(n2897), .Y(n4813) );
  CLKINVX1 U5637 ( .A(n6598), .Y(n6599) );
  OAI221X1 U5638 ( .A0(\i_MIPS/n350 ), .A1(n3091), .B0(\i_MIPS/n351 ), .B1(
        n3086), .C0(n4915), .Y(n5746) );
  OAI221X1 U5639 ( .A0(\i_MIPS/n363 ), .A1(n14), .B0(\i_MIPS/n362 ), .B1(n3077), .C0(n5464), .Y(n6475) );
  OAI221X1 U5640 ( .A0(\i_MIPS/n352 ), .A1(n3091), .B0(\i_MIPS/n353 ), .B1(
        n3085), .C0(n5052), .Y(n6135) );
  OAI221X1 U5641 ( .A0(\i_MIPS/n361 ), .A1(n3091), .B0(\i_MIPS/n360 ), .B1(
        n3085), .C0(n5458), .Y(n6463) );
  OAI221X1 U5642 ( .A0(\i_MIPS/n348 ), .A1(n3091), .B0(\i_MIPS/n349 ), .B1(
        n3087), .C0(n4812), .Y(n6123) );
  OA22X1 U5643 ( .A0(\i_MIPS/n350 ), .A1(n3082), .B0(\i_MIPS/n351 ), .B1(n3078), .Y(n4812) );
  OAI221X1 U5644 ( .A0(\i_MIPS/n348 ), .A1(n3082), .B0(\i_MIPS/n349 ), .B1(
        n3077), .C0(n4894), .Y(n5747) );
  AOI2BB1X1 U5645 ( .A0N(\i_MIPS/n347 ), .A1N(n3087), .B0(n2894), .Y(n4894) );
  OAI221X1 U5646 ( .A0(\i_MIPS/n366 ), .A1(n14), .B0(\i_MIPS/n365 ), .B1(n3077), .C0(n4892), .Y(n6333) );
  OAI222XL U5647 ( .A0(n3585), .A1(n199), .B0(n3667), .B1(n3582), .C0(n3689), 
        .C1(\i_MIPS/n186 ), .Y(n8798) );
  NAND2X1 U5648 ( .A(n2834), .B(n5483), .Y(n6402) );
  NAND4BX1 U5649 ( .AN(n6810), .B(n6809), .C(n6808), .D(n6807), .Y(n6821) );
  NAND4BX1 U5650 ( .AN(n6819), .B(n6818), .C(n6817), .D(n6816), .Y(n6820) );
  NAND4BX1 U5651 ( .AN(n5870), .B(n5869), .C(n5868), .D(n5867), .Y(n5881) );
  NAND4BX1 U5652 ( .AN(n5879), .B(n5878), .C(n5877), .D(n5876), .Y(n5880) );
  CLKMX2X2 U5653 ( .A(n6118), .B(n6117), .S0(n4015), .Y(n6119) );
  NAND4BX1 U5654 ( .AN(n6107), .B(n6106), .C(n6105), .D(n6104), .Y(n6118) );
  NAND4BX1 U5655 ( .AN(n6116), .B(n6115), .C(n6114), .D(n6113), .Y(n6117) );
  CLKMX2X2 U5656 ( .A(n6043), .B(n6042), .S0(n4014), .Y(n6044) );
  NAND4BX1 U5657 ( .AN(n6032), .B(n6031), .C(n6030), .D(n6029), .Y(n6043) );
  NAND4BX1 U5658 ( .AN(n6041), .B(n6040), .C(n6039), .D(n6038), .Y(n6042) );
  NAND4BX1 U5659 ( .AN(n5943), .B(n5942), .C(n5941), .D(n5940), .Y(n5954) );
  NAND4BX1 U5660 ( .AN(n5952), .B(n5951), .C(n5950), .D(n5949), .Y(n5953) );
  CLKMX2X2 U5661 ( .A(n5669), .B(n5668), .S0(n4014), .Y(n5670) );
  NAND4BX1 U5662 ( .AN(n5658), .B(n5657), .C(n5656), .D(n5655), .Y(n5669) );
  NAND4BX1 U5663 ( .AN(n5667), .B(n5666), .C(n5665), .D(n5664), .Y(n5668) );
  NAND4BX1 U5664 ( .AN(n5240), .B(n5239), .C(n5238), .D(n5237), .Y(n5251) );
  NAND4BX1 U5665 ( .AN(n5249), .B(n5248), .C(n5247), .D(n5246), .Y(n5250) );
  CLKMX2X2 U5666 ( .A(n5446), .B(n5445), .S0(n4014), .Y(n5447) );
  NAND4BX1 U5667 ( .AN(n5435), .B(n5434), .C(n5433), .D(n5432), .Y(n5446) );
  NAND4BX1 U5668 ( .AN(n5444), .B(n5443), .C(n5442), .D(n5441), .Y(n5445) );
  NAND4BX1 U5669 ( .AN(n6787), .B(n6786), .C(n6785), .D(n6784), .Y(n6798) );
  NAND4BX1 U5670 ( .AN(n6796), .B(n6795), .C(n6794), .D(n6793), .Y(n6797) );
  NAND4BX1 U5671 ( .AN(n5847), .B(n5846), .C(n5845), .D(n5844), .Y(n5858) );
  NAND4BX1 U5672 ( .AN(n5856), .B(n5855), .C(n5854), .D(n5853), .Y(n5857) );
  CLKMX2X2 U5673 ( .A(n6020), .B(n6019), .S0(n4013), .Y(n6023) );
  NAND4BX1 U5674 ( .AN(n6009), .B(n6008), .C(n6007), .D(n6006), .Y(n6020) );
  NAND4BX1 U5675 ( .AN(n6018), .B(n6017), .C(n6016), .D(n6015), .Y(n6019) );
  CLKMX2X2 U5676 ( .A(n6095), .B(n6094), .S0(n4012), .Y(n6098) );
  NAND4BX1 U5677 ( .AN(n6084), .B(n6083), .C(n6082), .D(n6081), .Y(n6095) );
  NAND4BX1 U5678 ( .AN(n6093), .B(n6092), .C(n6091), .D(n6090), .Y(n6094) );
  CLKMX2X2 U5679 ( .A(n6646), .B(n6645), .S0(n4012), .Y(n6647) );
  NAND4BX1 U5680 ( .AN(n6635), .B(n6634), .C(n6633), .D(n6632), .Y(n6646) );
  NAND4BX1 U5681 ( .AN(n6644), .B(n6643), .C(n6642), .D(n6641), .Y(n6645) );
  CLKMX2X2 U5682 ( .A(n5508), .B(n5507), .S0(n4013), .Y(n5511) );
  NAND4BX1 U5683 ( .AN(n5497), .B(n5496), .C(n5495), .D(n5494), .Y(n5508) );
  NAND4BX1 U5684 ( .AN(n5506), .B(n5505), .C(n5504), .D(n5503), .Y(n5507) );
  NAND4BX1 U5685 ( .AN(n5920), .B(n5919), .C(n5918), .D(n5917), .Y(n5931) );
  NAND4BX1 U5686 ( .AN(n5929), .B(n5928), .C(n5927), .D(n5926), .Y(n5930) );
  CLKMX2X2 U5687 ( .A(n6501), .B(n6500), .S0(n4013), .Y(n6504) );
  NAND4BX1 U5688 ( .AN(n6490), .B(n6489), .C(n6488), .D(n6487), .Y(n6501) );
  NAND4BX1 U5689 ( .AN(n6499), .B(n6498), .C(n6497), .D(n6496), .Y(n6500) );
  CLKMX2X2 U5690 ( .A(n5646), .B(n5645), .S0(n4013), .Y(n5649) );
  NAND4BX1 U5691 ( .AN(n5635), .B(n5634), .C(n5633), .D(n5632), .Y(n5646) );
  NAND4BX1 U5692 ( .AN(n5644), .B(n5643), .C(n5642), .D(n5641), .Y(n5645) );
  CLKMX2X2 U5693 ( .A(n6233), .B(n6232), .S0(n4012), .Y(n6234) );
  NAND4BX1 U5694 ( .AN(n6222), .B(n6221), .C(n6220), .D(n6219), .Y(n6233) );
  NAND4BX1 U5695 ( .AN(n6231), .B(n6230), .C(n6229), .D(n6228), .Y(n6232) );
  CLKMX2X2 U5696 ( .A(n6431), .B(n6430), .S0(n4012), .Y(n6432) );
  NAND4BX1 U5697 ( .AN(n6420), .B(n6419), .C(n6418), .D(n6417), .Y(n6431) );
  NAND4BX1 U5698 ( .AN(n6429), .B(n6428), .C(n6427), .D(n6426), .Y(n6430) );
  CLKMX2X2 U5699 ( .A(n6365), .B(n6364), .S0(n4012), .Y(n6366) );
  NAND4BX1 U5700 ( .AN(n6354), .B(n6353), .C(n6352), .D(n6351), .Y(n6365) );
  NAND4BX1 U5701 ( .AN(n6363), .B(n6362), .C(n6361), .D(n6360), .Y(n6364) );
  CLKMX2X2 U5702 ( .A(n5295), .B(n5294), .S0(n4012), .Y(n5296) );
  NAND4BX1 U5703 ( .AN(n5284), .B(n5283), .C(n5282), .D(n5281), .Y(n5295) );
  NAND4BX1 U5704 ( .AN(n5293), .B(n5292), .C(n5291), .D(n5290), .Y(n5294) );
  CLKMX2X2 U5705 ( .A(n5230), .B(n5229), .S0(n4013), .Y(n5231) );
  NAND4BX1 U5706 ( .AN(n5219), .B(n5218), .C(n5217), .D(n5216), .Y(n5230) );
  NAND4BX1 U5707 ( .AN(n5228), .B(n5227), .C(n5226), .D(n5225), .Y(n5229) );
  CLKMX2X2 U5708 ( .A(n5425), .B(n5424), .S0(n4012), .Y(n5426) );
  NAND4BX1 U5709 ( .AN(n5414), .B(n5413), .C(n5412), .D(n5411), .Y(n5425) );
  NAND4BX1 U5710 ( .AN(n5423), .B(n5422), .C(n5421), .D(n5420), .Y(n5424) );
  CLKMX2X2 U5711 ( .A(n5012), .B(n5011), .S0(n4013), .Y(n5013) );
  NAND4BX1 U5712 ( .AN(n5001), .B(n5000), .C(n4999), .D(n4998), .Y(n5012) );
  NAND4BX1 U5713 ( .AN(n5010), .B(n5009), .C(n5008), .D(n5007), .Y(n5011) );
  CLKMX2X2 U5714 ( .A(n4942), .B(n4941), .S0(n4013), .Y(n4943) );
  NAND4BX1 U5715 ( .AN(n4931), .B(n4930), .C(n4929), .D(n4928), .Y(n4942) );
  NAND4BX1 U5716 ( .AN(n4940), .B(n4939), .C(n4938), .D(n4937), .Y(n4941) );
  CLKMX2X2 U5717 ( .A(n5154), .B(n5153), .S0(n4013), .Y(n5155) );
  NAND4BX1 U5718 ( .AN(n5143), .B(n5142), .C(n5141), .D(n5140), .Y(n5154) );
  NAND4BX1 U5719 ( .AN(n5152), .B(n5151), .C(n5150), .D(n5149), .Y(n5153) );
  CLKMX2X2 U5720 ( .A(n6667), .B(n6666), .S0(n4015), .Y(n6668) );
  NAND4BX1 U5721 ( .AN(n6656), .B(n6655), .C(n6654), .D(n6653), .Y(n6667) );
  NAND4BX1 U5722 ( .AN(n6665), .B(n6664), .C(n6663), .D(n6662), .Y(n6666) );
  CLKMX2X2 U5723 ( .A(n6595), .B(n6594), .S0(n4015), .Y(n6596) );
  NAND4BX1 U5724 ( .AN(n6584), .B(n6583), .C(n6582), .D(n6581), .Y(n6595) );
  NAND4BX1 U5725 ( .AN(n6593), .B(n6592), .C(n6591), .D(n6590), .Y(n6594) );
  CLKMX2X2 U5726 ( .A(n5531), .B(n5530), .S0(n4014), .Y(n5532) );
  NAND4BX1 U5727 ( .AN(n5520), .B(n5519), .C(n5518), .D(n5517), .Y(n5531) );
  NAND4BX1 U5728 ( .AN(n5529), .B(n5528), .C(n5527), .D(n5526), .Y(n5530) );
  NAND4BX1 U5729 ( .AN(n4854), .B(n4853), .C(n4852), .D(n4851), .Y(n4865) );
  NAND4BX1 U5730 ( .AN(n4863), .B(n4862), .C(n4861), .D(n4860), .Y(n4864) );
  CLKMX2X2 U5731 ( .A(n6877), .B(n6876), .S0(\i_MIPS/IR_ID[20] ), .Y(n6880) );
  NAND4BX1 U5732 ( .AN(n6866), .B(n6865), .C(n6864), .D(n6863), .Y(n6877) );
  NAND4BX1 U5733 ( .AN(n6875), .B(n6874), .C(n6873), .D(n6872), .Y(n6876) );
  CLKMX2X2 U5734 ( .A(n6724), .B(n6723), .S0(\i_MIPS/IR_ID[20] ), .Y(n6725) );
  NAND4BX1 U5735 ( .AN(n6713), .B(n6712), .C(n6711), .D(n6710), .Y(n6724) );
  NAND4BX1 U5736 ( .AN(n6722), .B(n6721), .C(n6720), .D(n6719), .Y(n6723) );
  CLKMX2X2 U5737 ( .A(n6254), .B(n6253), .S0(n4014), .Y(n6255) );
  NAND4BX1 U5738 ( .AN(n6243), .B(n6242), .C(n6241), .D(n6240), .Y(n6254) );
  CLKMX2X2 U5739 ( .A(n6386), .B(n6385), .S0(n4015), .Y(n6387) );
  NAND4BX1 U5740 ( .AN(n6375), .B(n6374), .C(n6373), .D(n6372), .Y(n6386) );
  NAND4BX1 U5741 ( .AN(n6384), .B(n6383), .C(n6382), .D(n6381), .Y(n6385) );
  NAND4BX1 U5742 ( .AN(n5022), .B(n5021), .C(n5020), .D(n5019), .Y(n5033) );
  NAND4BX1 U5743 ( .AN(n5031), .B(n5030), .C(n5029), .D(n5028), .Y(n5032) );
  CLKMX2X2 U5744 ( .A(n5801), .B(n5800), .S0(n4014), .Y(n5802) );
  NAND4BX1 U5745 ( .AN(n5790), .B(n5789), .C(n5788), .D(n5787), .Y(n5801) );
  NAND4BX1 U5746 ( .AN(n5799), .B(n5798), .C(n5797), .D(n5796), .Y(n5800) );
  CLKMX2X2 U5747 ( .A(n5729), .B(n5728), .S0(n4014), .Y(n5730) );
  NAND4BX1 U5748 ( .AN(n5718), .B(n5717), .C(n5716), .D(n5715), .Y(n5729) );
  NAND4BX1 U5749 ( .AN(n5727), .B(n5726), .C(n5725), .D(n5724), .Y(n5728) );
  CLKMX2X2 U5750 ( .A(n6164), .B(n6163), .S0(n4012), .Y(n6165) );
  NAND4BX1 U5751 ( .AN(n6153), .B(n6152), .C(n6151), .D(n6150), .Y(n6164) );
  NAND4BX1 U5752 ( .AN(n6162), .B(n6161), .C(n6160), .D(n6159), .Y(n6163) );
  OA22X1 U5753 ( .A0(n3304), .A1(n1598), .B0(n3239), .B1(n177), .Y(n4535) );
  OA22X1 U5754 ( .A0(n3374), .A1(n1599), .B0(n3331), .B1(n178), .Y(n4534) );
  OAI221XL U5755 ( .A0(\i_MIPS/n349 ), .A1(n3091), .B0(\i_MIPS/n350 ), .B1(
        n3086), .C0(n4986), .Y(n5265) );
  OAI222XL U5756 ( .A0(n3585), .A1(n61), .B0(n3677), .B1(n3582), .C0(n3689), 
        .C1(\i_MIPS/n187 ), .Y(n8797) );
  NAND2X1 U5757 ( .A(n5484), .B(n5483), .Y(n6056) );
  OAI222XL U5758 ( .A0(n3584), .A1(n58), .B0(n3650), .B1(n3583), .C0(n3688), 
        .C1(\i_MIPS/n193 ), .Y(n8791) );
  OAI222XL U5759 ( .A0(n3584), .A1(n62), .B0(n3647), .B1(n3583), .C0(n3688), 
        .C1(\i_MIPS/n195 ), .Y(n8789) );
  AOI2BB1X1 U5760 ( .A0N(\i_MIPS/n346 ), .A1N(n3087), .B0(n2896), .Y(n4967) );
  NAND2X1 U5761 ( .A(n6763), .B(n6762), .Y(n6769) );
  OA22X1 U5762 ( .A0(\i_MIPS/n353 ), .A1(n14), .B0(\i_MIPS/n354 ), .B1(n3078), 
        .Y(n5112) );
  OAI222XL U5763 ( .A0(n3070), .A1(n4730), .B0(n4729), .B1(n3071), .C0(n2875), 
        .C1(n3096), .Y(n4731) );
  OAI222XL U5764 ( .A0(n6460), .A1(n7001), .B0(n5904), .B1(n6403), .C0(n5827), 
        .C1(n6996), .Y(n5830) );
  AOI211X1 U5765 ( .A0(n5826), .A1(n8), .B0(n2896), .C0(n2895), .Y(n5827) );
  CLKINVX1 U5766 ( .A(n5825), .Y(n5826) );
  OAI222XL U5767 ( .A0(n7001), .A1(n6907), .B0(n6138), .B1(n6544), .C0(n6137), 
        .C1(n6136), .Y(n6140) );
  OA22X1 U5768 ( .A0(n6840), .A1(n3107), .B0(n3099), .B1(n6839), .Y(n6843) );
  OAI222XL U5769 ( .A0(n5904), .A1(n6270), .B0(n5903), .B1(n6996), .C0(n5902), 
        .C1(n7001), .Y(n5907) );
  AOI211X1 U5770 ( .A0(n5901), .A1(n8), .B0(n2897), .C0(n2894), .Y(n5903) );
  CLKINVX1 U5771 ( .A(n6994), .Y(n5901) );
  NOR4X1 U5772 ( .A(n8516), .B(n8515), .C(n8514), .D(n8513), .Y(n8904) );
  NAND4X1 U5773 ( .A(n4552), .B(n4551), .C(n4550), .D(n4549), .Y(n8651) );
  OA22X1 U5774 ( .A0(n3287), .A1(n472), .B0(n3239), .B1(n1387), .Y(n4552) );
  OA22X1 U5775 ( .A0(n3471), .A1(n473), .B0(n3415), .B1(n1388), .Y(n4550) );
  OA22X1 U5776 ( .A0(n3374), .A1(n474), .B0(n3331), .B1(n1389), .Y(n4551) );
  NAND4X1 U5777 ( .A(n4562), .B(n4561), .C(n4560), .D(n4559), .Y(n8555) );
  OA22X1 U5778 ( .A0(n3287), .A1(n475), .B0(n3240), .B1(n1390), .Y(n4562) );
  OA22X1 U5779 ( .A0(n3464), .A1(n476), .B0(n3416), .B1(n1391), .Y(n4560) );
  OA22X1 U5780 ( .A0(n3375), .A1(n477), .B0(n3332), .B1(n1392), .Y(n4561) );
  NAND4X1 U5781 ( .A(n4567), .B(n4566), .C(n4565), .D(n4564), .Y(n8587) );
  OA22X1 U5782 ( .A0(n3287), .A1(n478), .B0(n3240), .B1(n1393), .Y(n4567) );
  OA22X1 U5783 ( .A0(n3464), .A1(n479), .B0(n3416), .B1(n1394), .Y(n4565) );
  OA22X1 U5784 ( .A0(n3375), .A1(n480), .B0(n3332), .B1(n1395), .Y(n4566) );
  NAND4X1 U5785 ( .A(n4557), .B(n4556), .C(n4555), .D(n4554), .Y(n8619) );
  OA22X1 U5786 ( .A0(n3287), .A1(n481), .B0(n3240), .B1(n1396), .Y(n4557) );
  OA22X1 U5787 ( .A0(n3464), .A1(n482), .B0(n3416), .B1(n1397), .Y(n4555) );
  OA22X1 U5788 ( .A0(n3375), .A1(n483), .B0(n3332), .B1(n1398), .Y(n4556) );
  NAND4X1 U5789 ( .A(n7370), .B(n7369), .C(n7368), .D(n7367), .Y(n8650) );
  OA22X1 U5790 ( .A0(n3290), .A1(n679), .B0(n3243), .B1(n1600), .Y(n7370) );
  OA22X1 U5791 ( .A0(n3468), .A1(n684), .B0(n3421), .B1(n1601), .Y(n7368) );
  OA22X1 U5792 ( .A0(n3377), .A1(n680), .B0(n3335), .B1(n1602), .Y(n7369) );
  NAND4X1 U5793 ( .A(n7378), .B(n7377), .C(n7376), .D(n7375), .Y(n8554) );
  OA22X1 U5794 ( .A0(n3291), .A1(n681), .B0(n3244), .B1(n1603), .Y(n7378) );
  OA22X1 U5795 ( .A0(n3469), .A1(n685), .B0(n3422), .B1(n1604), .Y(n7376) );
  OA22X1 U5796 ( .A0(n3378), .A1(n686), .B0(n3336), .B1(n1605), .Y(n7377) );
  NAND4X1 U5797 ( .A(n7382), .B(n7381), .C(n7380), .D(n7379), .Y(n8586) );
  OA22X1 U5798 ( .A0(n3291), .A1(n682), .B0(n3244), .B1(n1606), .Y(n7382) );
  OA22X1 U5799 ( .A0(n3469), .A1(n687), .B0(n3422), .B1(n1607), .Y(n7380) );
  OA22X1 U5800 ( .A0(n3378), .A1(n688), .B0(n3336), .B1(n1608), .Y(n7381) );
  NAND4X1 U5801 ( .A(n7374), .B(n7373), .C(n7372), .D(n7371), .Y(n8618) );
  OA22X1 U5802 ( .A0(n3291), .A1(n683), .B0(n3244), .B1(n1609), .Y(n7374) );
  OA22X1 U5803 ( .A0(n3469), .A1(n689), .B0(n3422), .B1(n1610), .Y(n7372) );
  OA22X1 U5804 ( .A0(n3378), .A1(n690), .B0(n3336), .B1(n1611), .Y(n7373) );
  NAND4X1 U5805 ( .A(n4543), .B(n4542), .C(n4541), .D(n4540), .Y(n8653) );
  OA22X1 U5806 ( .A0(n3374), .A1(n434), .B0(n3331), .B1(n1349), .Y(n4542) );
  OA22X1 U5807 ( .A0(n3287), .A1(n435), .B0(n3239), .B1(n1350), .Y(n4543) );
  NAND4X1 U5808 ( .A(n7322), .B(n7321), .C(n7320), .D(n7319), .Y(n8557) );
  OA22X1 U5809 ( .A0(n3553), .A1(n436), .B0(n3511), .B1(n1351), .Y(n7319) );
  OA22X1 U5810 ( .A0(n3376), .A1(n437), .B0(n3334), .B1(n1352), .Y(n7321) );
  OA22X1 U5811 ( .A0(n3289), .A1(n438), .B0(n3242), .B1(n1353), .Y(n7322) );
  NAND4X1 U5812 ( .A(n7326), .B(n7325), .C(n7324), .D(n7323), .Y(n8589) );
  OA22X1 U5813 ( .A0(n3553), .A1(n439), .B0(n3511), .B1(n1354), .Y(n7323) );
  OA22X1 U5814 ( .A0(n3376), .A1(n440), .B0(n3334), .B1(n1355), .Y(n7325) );
  OA22X1 U5815 ( .A0(n3289), .A1(n441), .B0(n3242), .B1(n1356), .Y(n7326) );
  NAND4X1 U5816 ( .A(n7318), .B(n7317), .C(n7316), .D(n7315), .Y(n8621) );
  OA22X1 U5817 ( .A0(n3553), .A1(n442), .B0(n3511), .B1(n1357), .Y(n7315) );
  OA22X1 U5818 ( .A0(n3376), .A1(n443), .B0(n3334), .B1(n1358), .Y(n7317) );
  OA22X1 U5819 ( .A0(n3289), .A1(n444), .B0(n3242), .B1(n1359), .Y(n7318) );
  AOI2BB1X1 U5820 ( .A0N(n6527), .A1N(n8), .B0(n2900), .Y(n5127) );
  NAND2X1 U5821 ( .A(n4672), .B(\i_MIPS/n365 ), .Y(n8506) );
  NAND2X1 U5822 ( .A(n4640), .B(\i_MIPS/n350 ), .Y(n8548) );
  NAND2X1 U5823 ( .A(n4660), .B(\i_MIPS/n352 ), .Y(n5621) );
  NAND2X1 U5824 ( .A(n4626), .B(\i_MIPS/n346 ), .Y(n8522) );
  NAND2X1 U5825 ( .A(n4631), .B(\i_MIPS/n350 ), .Y(n6690) );
  NAND2X1 U5826 ( .A(n4647), .B(\i_MIPS/n356 ), .Y(n8488) );
  AOI211X1 U5827 ( .A0(n6905), .A1(n6054), .B0(n5207), .C0(n5206), .Y(n5208)
         );
  NAND2X1 U5828 ( .A(n4674), .B(\i_MIPS/n365 ), .Y(n4972) );
  NAND2X1 U5829 ( .A(n4657), .B(\i_MIPS/n354 ), .Y(n5734) );
  NAND4X1 U5830 ( .A(n7548), .B(n7547), .C(n7546), .D(n7545), .Y(n8569) );
  OA22X1 U5831 ( .A0(n3294), .A1(n484), .B0(n3247), .B1(n1399), .Y(n7548) );
  OA22X1 U5832 ( .A0(n3381), .A1(n485), .B0(n3339), .B1(n1400), .Y(n7547) );
  OA22X1 U5833 ( .A0(n3558), .A1(n486), .B0(n3516), .B1(n1401), .Y(n7545) );
  NAND4X1 U5834 ( .A(n7543), .B(n7542), .C(n7541), .D(n7540), .Y(n8633) );
  OA22X1 U5835 ( .A0(n3558), .A1(n445), .B0(n3516), .B1(n1360), .Y(n7540) );
  OA22X1 U5836 ( .A0(n3381), .A1(n1374), .B0(n3339), .B1(n451), .Y(n7542) );
  OA22X1 U5837 ( .A0(n3294), .A1(n1375), .B0(n3247), .B1(n452), .Y(n7543) );
  NAND4X1 U5838 ( .A(n7538), .B(n7537), .C(n7536), .D(n7535), .Y(n8665) );
  OA22X1 U5839 ( .A0(n3558), .A1(n1376), .B0(n3516), .B1(n453), .Y(n7535) );
  OA22X1 U5840 ( .A0(n3381), .A1(n1377), .B0(n3339), .B1(n454), .Y(n7537) );
  OA22X1 U5841 ( .A0(n3294), .A1(n1378), .B0(n3247), .B1(n455), .Y(n7538) );
  NAND2X1 U5842 ( .A(n4645), .B(\i_MIPS/n357 ), .Y(n8485) );
  NAND2X1 U5843 ( .A(n4691), .B(\i_MIPS/n361 ), .Y(n5256) );
  NAND2X1 U5844 ( .A(n8482), .B(n8480), .Y(n6266) );
  NAND2X1 U5845 ( .A(n6391), .B(n6390), .Y(n6263) );
  AO22X1 U5846 ( .A0(n6262), .A1(n3101), .B0(n3108), .B1(n6392), .Y(n6264) );
  XNOR2X1 U5847 ( .A(\D_cache/N39 ), .B(DCACHE_addr[22]), .Y(\D_cache/n542 )
         );
  XNOR2X1 U5848 ( .A(\D_cache/N34 ), .B(DCACHE_addr[27]), .Y(\D_cache/n541 )
         );
  NAND3X1 U5849 ( .A(\D_cache/n554 ), .B(\D_cache/n555 ), .C(\D_cache/n556 ), 
        .Y(\D_cache/n550 ) );
  XNOR2X1 U5850 ( .A(\D_cache/N41 ), .B(DCACHE_addr[20]), .Y(\D_cache/n556 )
         );
  XNOR2X1 U5851 ( .A(\D_cache/N38 ), .B(DCACHE_addr[23]), .Y(\D_cache/n540 )
         );
  OAI221XL U5852 ( .A0(\i_MIPS/n340 ), .A1(n7005), .B0(n4723), .B1(n7005), 
        .C0(n4722), .Y(n4732) );
  CLKINVX1 U5853 ( .A(n5823), .Y(n5467) );
  CLKINVX1 U5854 ( .A(n6200), .Y(n5468) );
  OAI221XL U5855 ( .A0(n3070), .A1(n5821), .B0(n2876), .B1(n3096), .C0(n5820), 
        .Y(n5831) );
  AOI222X1 U5856 ( .A0(n5819), .A1(n6682), .B0(n5818), .B1(n7006), .C0(n5817), 
        .C1(n6477), .Y(n5820) );
  CLKINVX1 U5857 ( .A(n5816), .Y(n5818) );
  CLKINVX1 U5858 ( .A(n6401), .Y(n5819) );
  AND3X2 U5859 ( .A(n5974), .B(n3076), .C(n6682), .Y(n5995) );
  OAI222XL U5860 ( .A0(n3070), .A1(n5989), .B0(n6056), .B1(n6137), .C0(n6906), 
        .C1(n6908), .Y(n5996) );
  AND2X2 U5861 ( .A(n2813), .B(n6619), .Y(n6070) );
  OAI222XL U5862 ( .A0(n3070), .A1(n6064), .B0(n6057), .B1(n6056), .C0(n6055), 
        .C1(n6908), .Y(n6071) );
  AO22X1 U5863 ( .A0(n6832), .A1(n6685), .B0(n6684), .B1(n6993), .Y(n6700) );
  AND2X2 U5864 ( .A(n2805), .B(n6686), .Y(n6699) );
  NAND2X1 U5865 ( .A(n6339), .B(n6335), .Y(n6326) );
  NAND2X1 U5866 ( .A(n6404), .B(n6400), .Y(n6396) );
  AOI2BB2X1 U5867 ( .B0(\D_cache/N144 ), .B1(n2153), .A0N(n24), .A1N(n8894), 
        .Y(\D_cache/n169 ) );
  AOI2BB2X1 U5868 ( .B0(\D_cache/N138 ), .B1(n2153), .A0N(n3040), .A1N(n8888), 
        .Y(\D_cache/n194 ) );
  AOI2BB2X1 U5869 ( .B0(\D_cache/N136 ), .B1(n2153), .A0N(n24), .A1N(n8886), 
        .Y(\D_cache/n192 ) );
  AOI222XL U5870 ( .A0(n6680), .A1(n6053), .B0(n6052), .B1(n7006), .C0(n6051), 
        .C1(n6990), .Y(n6073) );
  NAND2X1 U5871 ( .A(n4704), .B(n5900), .Y(n8530) );
  NAND2X1 U5872 ( .A(n4673), .B(\i_MIPS/n364 ), .Y(n4987) );
  NAND2X1 U5873 ( .A(n6992), .B(\i_MIPS/n341 ), .Y(n8525) );
  XOR2X1 U5874 ( .A(n7958), .B(n7811), .Y(n5599) );
  NAND2X1 U5875 ( .A(n4643), .B(\i_MIPS/n353 ), .Y(n4827) );
  NAND2X1 U5876 ( .A(n4703), .B(\i_MIPS/n344 ), .Y(n8518) );
  CLKINVX1 U5877 ( .A(n6128), .Y(n5188) );
  NAND2X1 U5878 ( .A(n4705), .B(\i_MIPS/n342 ), .Y(n8531) );
  NAND2X1 U5879 ( .A(n6468), .B(n4833), .Y(n4838) );
  AO22X1 U5880 ( .A0(n2848), .A1(n3100), .B0(n3110), .B1(n4834), .Y(n4839) );
  NAND3BX1 U5881 ( .AN(n8460), .B(n2841), .C(n8533), .Y(n8912) );
  NAND2X1 U5882 ( .A(n8535), .B(n8537), .Y(n5606) );
  NAND2X1 U5883 ( .A(n5549), .B(n5545), .Y(n5543) );
  NAND2X1 U5884 ( .A(n8488), .B(n8477), .Y(n5542) );
  AO22X1 U5885 ( .A0(n2823), .A1(n3102), .B0(n3110), .B1(n5540), .Y(n5544) );
  XOR2X1 U5886 ( .A(n8046), .B(n8051), .Y(n8047) );
  AOI21X1 U5887 ( .A0(n8062), .A1(n8045), .B0(n8044), .Y(n8046) );
  NAND4X1 U5888 ( .A(n6345), .B(n6344), .C(n6343), .D(n6342), .Y(n8251) );
  OA22X1 U5889 ( .A0(n7008), .A1(n6402), .B0(n6335), .B1(n3070), .Y(n6344) );
  OA22X1 U5890 ( .A0(n2796), .A1(n6989), .B0(n6544), .B1(n6338), .Y(n6343) );
  AOI2BB1X1 U5891 ( .A0N(n6341), .A1N(n6550), .B0(n6340), .Y(n6342) );
  OAI221XL U5892 ( .A0(n6755), .A1(n7001), .B0(n6754), .B1(n6996), .C0(n6753), 
        .Y(n6778) );
  AOI222X1 U5893 ( .A0(n6689), .A1(n6993), .B0(n2805), .B1(n6477), .C0(n6476), 
        .C1(n6475), .Y(n6478) );
  AND2X2 U5894 ( .A(n6548), .B(n6614), .Y(n2835) );
  OAI22XL U5895 ( .A0(n6551), .A1(n6550), .B0(n6549), .B1(n6996), .Y(n2836) );
  MXI2X1 U5896 ( .A(n7005), .B(n3071), .S0(n6553), .Y(n2837) );
  OAI221XL U5897 ( .A0(n7001), .A1(n5684), .B0(n6996), .B1(n5816), .C0(n5461), 
        .Y(n5488) );
  AOI222X1 U5898 ( .A0(n6060), .A1(n6993), .B0(n2813), .B1(n5815), .C0(n6205), 
        .C1(n5756), .Y(n5485) );
  XNOR2X1 U5899 ( .A(n2703), .B(\D_cache/N56 ), .Y(\D_cache/n538 ) );
  NAND2X1 U5900 ( .A(n6909), .B(n8539), .Y(n6924) );
  NAND2X1 U5901 ( .A(n6834), .B(n8545), .Y(n6853) );
  AND2X2 U5902 ( .A(n4826), .B(n8537), .Y(n2838) );
  NAND2BX1 U5903 ( .AN(n3000), .B(n8625), .Y(n7757) );
  NAND2BX2 U5904 ( .AN(n2163), .B(n8657), .Y(n7758) );
  NAND2BX1 U5905 ( .AN(n3001), .B(n8593), .Y(n7755) );
  NAND2BX1 U5906 ( .AN(n3000), .B(n8631), .Y(n7582) );
  NAND2BX1 U5907 ( .AN(n2163), .B(n8663), .Y(n7583) );
  NAND2BX1 U5908 ( .AN(n3001), .B(n8599), .Y(n7580) );
  NAND2BX1 U5909 ( .AN(n3000), .B(n8623), .Y(n7409) );
  NAND2BX1 U5910 ( .AN(n2163), .B(n8655), .Y(n7410) );
  NAND2BX1 U5911 ( .AN(n3000), .B(n8622), .Y(n7345) );
  NAND2BX1 U5912 ( .AN(n3001), .B(n8590), .Y(n7343) );
  NAND2BX1 U5913 ( .AN(n2163), .B(n8654), .Y(n7346) );
  NAND2BX1 U5914 ( .AN(n3000), .B(n8629), .Y(n7606) );
  NAND2BX1 U5915 ( .AN(n3001), .B(n8597), .Y(n7604) );
  NAND2BX1 U5916 ( .AN(n3000), .B(n8620), .Y(n7365) );
  NAND2BX1 U5917 ( .AN(n3001), .B(n8588), .Y(n7363) );
  NAND2BX1 U5918 ( .AN(n3576), .B(n8556), .Y(n7364) );
  NAND2BX1 U5919 ( .AN(n3001), .B(n8594), .Y(n7728) );
  AOI2BB1X1 U5920 ( .A0N(n8495), .A1N(n8494), .B0(n8496), .Y(n8501) );
  OA22X1 U5921 ( .A0(n5546), .A1(n6402), .B0(n3070), .B1(n5545), .Y(n5554) );
  OA22X1 U5922 ( .A0(n6847), .A1(n5548), .B0(n6544), .B1(n5547), .Y(n5553) );
  AOI2BB1X1 U5923 ( .A0N(n5551), .A1N(n6550), .B0(n5550), .Y(n5552) );
  OA22X1 U5924 ( .A0(n2796), .A1(n6270), .B0(n6544), .B1(n6269), .Y(n6274) );
  AOI2BB1X1 U5925 ( .A0N(n6272), .A1N(n6550), .B0(n6271), .Y(n6273) );
  OA22X1 U5926 ( .A0(n6402), .A1(n6401), .B0(n3070), .B1(n6400), .Y(n6410) );
  OA22X1 U5927 ( .A0(n2796), .A1(n6403), .B0(n2831), .B1(n6544), .Y(n6409) );
  AOI2BB1X1 U5928 ( .A0N(n6407), .A1N(n6550), .B0(n6406), .Y(n6408) );
  CLKINVX1 U5929 ( .A(n8321), .Y(n8303) );
  AOI211X1 U5930 ( .A0(n6905), .A1(n5898), .B0(n5333), .C0(n5332), .Y(n5334)
         );
  OAI222XL U5931 ( .A0(n3070), .A1(n5890), .B0(n5899), .B1(n7010), .C0(n5888), 
        .C1(n5958), .Y(n5911) );
  AOI211X1 U5932 ( .A0(n5908), .A1(n6682), .B0(n5907), .C0(n5906), .Y(n5909)
         );
  AOI211X1 U5933 ( .A0(n6905), .A1(n6141), .B0(n6140), .C0(n6139), .Y(n6142)
         );
  AOI211X1 U5934 ( .A0(n6905), .A1(n6773), .B0(n5272), .C0(n5271), .Y(n5273)
         );
  AOI221X1 U5935 ( .A0(n4980), .A1(n4979), .B0(n4978), .B1(n4977), .C0(n4976), 
        .Y(n4991) );
  OAI222XL U5936 ( .A0(n3070), .A1(n6127), .B0(n6826), .B1(n6402), .C0(n5551), 
        .C1(n5548), .Y(n4992) );
  NAND2X1 U5937 ( .A(n3076), .B(n5483), .Y(n6849) );
  NAND2X1 U5938 ( .A(n5205), .B(n5970), .Y(n6057) );
  NAND2X1 U5939 ( .A(n4630), .B(\i_MIPS/n345 ), .Y(n8517) );
  NAND2X1 U5940 ( .A(n6693), .B(n6841), .Y(n4641) );
  NAND2X1 U5941 ( .A(n5469), .B(n8524), .Y(n8462) );
  NOR2X4 U5942 ( .A(n4463), .B(n4462), .Y(n4530) );
  NOR2X4 U5943 ( .A(n4495), .B(n4494), .Y(n4529) );
  AOI2BB1X1 U5944 ( .A0N(n5194), .A1N(n5193), .B0(n5192), .Y(n5195) );
  CLKINVX1 U5945 ( .A(n6129), .Y(n5194) );
  OA22X1 U5946 ( .A0(n3372), .A1(n145), .B0(n3329), .B1(n1036), .Y(n4474) );
  OA22X1 U5947 ( .A0(n3372), .A1(n146), .B0(n3329), .B1(n1037), .Y(n4470) );
  OA22X1 U5948 ( .A0(n3285), .A1(n147), .B0(n3237), .B1(n1038), .Y(n4471) );
  OA22X1 U5949 ( .A0(n3547), .A1(n148), .B0(n3506), .B1(n1039), .Y(n4464) );
  OA22X1 U5950 ( .A0(n3372), .A1(n149), .B0(n3329), .B1(n1040), .Y(n4466) );
  OA22X1 U5951 ( .A0(n3285), .A1(n150), .B0(n3237), .B1(n1041), .Y(n4467) );
  OA22X1 U5952 ( .A0(n3373), .A1(n151), .B0(n3330), .B1(n1042), .Y(n4502) );
  OA22X1 U5953 ( .A0(n3286), .A1(n152), .B0(n3238), .B1(n1043), .Y(n4503) );
  OA22X1 U5954 ( .A0(n3373), .A1(n153), .B0(n3330), .B1(n1044), .Y(n4498) );
  OA22X1 U5955 ( .A0(n3286), .A1(n154), .B0(n3238), .B1(n1045), .Y(n4499) );
  CLKINVX1 U5956 ( .A(n7043), .Y(n3023) );
  NAND2X1 U5957 ( .A(n8465), .B(n8549), .Y(n5979) );
  NAND4X2 U5958 ( .A(n4455), .B(n4454), .C(n4453), .D(n4452), .Y(n8705) );
  NAND4X2 U5959 ( .A(n4459), .B(n4458), .C(n4457), .D(n4456), .Y(n8710) );
  NAND2X1 U5960 ( .A(n5738), .B(n5602), .Y(n4666) );
  OA22X1 U5961 ( .A0(n3372), .A1(n156), .B0(n3329), .B1(n1047), .Y(n4478) );
  OA22X1 U5962 ( .A0(n3463), .A1(n157), .B0(n3442), .B1(n1048), .Y(n4509) );
  NAND2X1 U5963 ( .A(n8510), .B(n6191), .Y(n5193) );
  AOI2BB1X1 U5964 ( .A0N(n6598), .A1N(n8), .B0(n5043), .Y(n5046) );
  NAND2X1 U5965 ( .A(n6468), .B(n6474), .Y(n5985) );
  CLKINVX1 U5966 ( .A(n5474), .Y(n6060) );
  NAND2BX2 U5967 ( .AN(n3576), .B(n8557), .Y(n7328) );
  AOI2BB2X2 U5968 ( .B0(\D_cache/N146 ), .B1(n2153), .A0N(n24), .A1N(n8896), 
        .Y(\D_cache/n171 ) );
  OA22X1 U5969 ( .A0(n3374), .A1(n158), .B0(n3331), .B1(n1049), .Y(n4518) );
  OA22X1 U5970 ( .A0(n3373), .A1(n159), .B0(n3330), .B1(n1050), .Y(n4506) );
  OA22X1 U5971 ( .A0(n3286), .A1(n160), .B0(n3238), .B1(n1051), .Y(n4507) );
  CLKINVX1 U5972 ( .A(n4723), .Y(n4707) );
  CLKMX2X2 U5973 ( .A(n5780), .B(n5779), .S0(n4013), .Y(n5781) );
  NAND4BX1 U5974 ( .AN(n5769), .B(n5768), .C(n5767), .D(n5766), .Y(n5780) );
  AOI222X1 U5975 ( .A0(n2809), .A1(n6477), .B0(n5394), .B1(n5393), .C0(n5392), 
        .C1(n5391), .Y(n5404) );
  CLKINVX1 U5976 ( .A(n4673), .Y(n4686) );
  CLKINVX1 U5977 ( .A(n4691), .Y(n4688) );
  CLKINVX1 U5978 ( .A(n4653), .Y(n4651) );
  CLKINVX1 U5979 ( .A(n4654), .Y(n4645) );
  CLKINVX1 U5980 ( .A(n4646), .Y(n4647) );
  AND2X2 U5981 ( .A(n8528), .B(n8459), .Y(n2841) );
  CLKINVX1 U5982 ( .A(n6191), .Y(n8516) );
  CLKINVX1 U5983 ( .A(n8541), .Y(n5047) );
  CLKINVX1 U5984 ( .A(n7632), .Y(\i_MIPS/EX_MEM_next[70] ) );
  AO21X1 U5985 ( .A0(n8546), .A1(n8545), .B0(n8544), .Y(n8917) );
  OAI22XL U5986 ( .A0(n8915), .A1(n8914), .B0(n2838), .B1(n8915), .Y(n8919) );
  AO21X1 U5987 ( .A0(n8538), .A1(n8537), .B0(n8536), .Y(n8915) );
  AO21X1 U5988 ( .A0(n2845), .A1(n8524), .B0(n8523), .Y(n8907) );
  AO21X1 U5989 ( .A0(n8534), .A1(n8533), .B0(n8532), .Y(n8805) );
  AO21X1 U5990 ( .A0(n8529), .A1(n8528), .B0(n8527), .Y(n8909) );
  CLKINVX1 U5991 ( .A(n8477), .Y(n8486) );
  AOI21X1 U5992 ( .A0(n6982), .A1(n8525), .B0(n4607), .Y(n2843) );
  CLKMX2X2 U5993 ( .A(n5708), .B(n5707), .S0(n4013), .Y(n5709) );
  NAND4BX1 U5994 ( .AN(n5697), .B(n5696), .C(n5695), .D(n5694), .Y(n5708) );
  CLKINVX1 U5995 ( .A(n5989), .Y(n5471) );
  AND2X2 U5996 ( .A(n4627), .B(\i_MIPS/n347 ), .Y(n2845) );
  NAND2BX1 U5997 ( .AN(n4618), .B(n2885), .Y(n4612) );
  AOI21X1 U5998 ( .A0(n6839), .A1(n6834), .B0(n5983), .Y(n2846) );
  INVX3 U5999 ( .A(n4891), .Y(n8224) );
  OAI222X1 U6000 ( .A0(n4890), .A1(n3166), .B0(n4889), .B1(n2761), .C0(n8744), 
        .C1(n3163), .Y(n4891) );
  CLKMX2X2 U6001 ( .A(n4888), .B(n4887), .S0(n4013), .Y(n4889) );
  NAND4BX1 U6002 ( .AN(n4877), .B(n4876), .C(n4875), .D(n4874), .Y(n4888) );
  CLKMX2X2 U6003 ( .A(n5202), .B(n4916), .S0(n4016), .Y(n6338) );
  CLKMX2X2 U6004 ( .A(n6900), .B(n6899), .S0(n4012), .Y(n6901) );
  NAND4BX1 U6005 ( .AN(n6889), .B(n6888), .C(n6887), .D(n6886), .Y(n6900) );
  CLKMX2X2 U6006 ( .A(n6745), .B(n6744), .S0(n4012), .Y(n6746) );
  NAND4BX1 U6007 ( .AN(n6734), .B(n6733), .C(n6732), .D(n6731), .Y(n6745) );
  CLKMX2X2 U6008 ( .A(n5320), .B(n5329), .S0(n4016), .Y(n6138) );
  CLKMX2X2 U6009 ( .A(n1617), .B(\D_cache/n189 ), .S0(n4023), .Y(n5647) );
  OAI221X1 U6010 ( .A0(n8765), .A1(n7044), .B0(n8752), .B1(n7043), .C0(n5509), 
        .Y(n5510) );
  CLKMX2X2 U6011 ( .A(n1089), .B(\D_cache/n182 ), .S0(n4023), .Y(n5509) );
  CLKINVX1 U6012 ( .A(n5891), .Y(n8460) );
  CLKMX2X2 U6013 ( .A(n6969), .B(n6968), .S0(n4012), .Y(n6970) );
  NAND4BX1 U6014 ( .AN(n6958), .B(n6957), .C(n6956), .D(n6955), .Y(n6969) );
  CLKMX2X2 U6015 ( .A(n4963), .B(n4962), .S0(n4015), .Y(n4964) );
  NAND4BX1 U6016 ( .AN(n4952), .B(n4951), .C(n4950), .D(n4949), .Y(n4963) );
  NAND4BX1 U6017 ( .AN(n4961), .B(n4960), .C(n4959), .D(n4958), .Y(n4962) );
  CLKMX2X2 U6018 ( .A(n5175), .B(n5174), .S0(n4015), .Y(n5176) );
  NAND4BX1 U6019 ( .AN(n5164), .B(n5163), .C(n5162), .D(n5161), .Y(n5175) );
  NAND4BX1 U6020 ( .AN(n5173), .B(n5172), .C(n5171), .D(n5170), .Y(n5174) );
  NAND2X1 U6021 ( .A(n4729), .B(n4730), .Y(n4737) );
  NOR2X1 U6022 ( .A(n2891), .B(n2890), .Y(\i_MIPS/forward_unit/n32 ) );
  OAI2BB1X4 U6023 ( .A0N(n6986), .A1N(n7002), .B0(n6988), .Y(n4708) );
  AO21X2 U6024 ( .A0(n3580), .A1(n8025), .B0(n2859), .Y(n8061) );
  OAI2BB1X1 U6025 ( .A0N(n5257), .A1N(n5256), .B0(n5255), .Y(n5260) );
  CLKMX2X2 U6026 ( .A(n6574), .B(n6573), .S0(n4012), .Y(n6575) );
  NAND4BX1 U6027 ( .AN(n6563), .B(n6562), .C(n6561), .D(n6560), .Y(n6574) );
  NAND4BX1 U6028 ( .AN(n6572), .B(n6571), .C(n6570), .D(n6569), .Y(n6573) );
  CLKMX2X2 U6029 ( .A(n1619), .B(\D_cache/n184 ), .S0(n4022), .Y(n6878) );
  AOI2BB2X2 U6030 ( .B0(\D_cache/N129 ), .B1(n2153), .A0N(n24), .A1N(n8879), 
        .Y(\D_cache/n184 ) );
  CLKMX2X2 U6031 ( .A(n1090), .B(\D_cache/n183 ), .S0(n4022), .Y(n6021) );
  CLKMX2X3 U6032 ( .A(n1084), .B(\D_cache/n180 ), .S0(n4023), .Y(n6799) );
  OAI221X1 U6033 ( .A0(n8764), .A1(n7044), .B0(n8751), .B1(n7043), .C0(n6096), 
        .Y(n6097) );
  CLKMX2X2 U6034 ( .A(n1618), .B(\D_cache/n181 ), .S0(n4022), .Y(n6096) );
  OAI221XL U6035 ( .A0(n8760), .A1(n7044), .B0(n8747), .B1(n7043), .C0(n7042), 
        .Y(n7045) );
  CLKMX2X2 U6036 ( .A(n1616), .B(\D_cache/n176 ), .S0(n4021), .Y(n7042) );
  AOI2BB2X1 U6037 ( .B0(\D_cache/N122 ), .B1(n2153), .A0N(n23), .A1N(n8872), 
        .Y(\D_cache/n176 ) );
  CLKINVX1 U6038 ( .A(n6477), .Y(n5117) );
  AND2X2 U6039 ( .A(n3075), .B(n8), .Y(n2863) );
  AND4X1 U6040 ( .A(\D_cache/n218 ), .B(\D_cache/N30 ), .C(n3957), .D(
        \D_cache/n520 ), .Y(n2866) );
  CLKINVX1 U6041 ( .A(n8526), .Y(n8527) );
  CLKMX2X2 U6042 ( .A(n6452), .B(n6451), .S0(n4014), .Y(n6453) );
  NAND4BX1 U6043 ( .AN(n6441), .B(n6440), .C(n6439), .D(n6438), .Y(n6452) );
  CLKMX2X2 U6044 ( .A(n5356), .B(n5355), .S0(n4013), .Y(n5357) );
  NAND4BX1 U6045 ( .AN(n5345), .B(n5344), .C(n5343), .D(n5342), .Y(n5356) );
  CLKMX2X2 U6046 ( .A(n5082), .B(n5081), .S0(n4013), .Y(n5083) );
  NAND4BX1 U6047 ( .AN(n5071), .B(n5070), .C(n5069), .D(n5068), .Y(n5082) );
  CLKINVX1 U6048 ( .A(n8601), .Y(n7555) );
  CLKMX2X2 U6049 ( .A(n6317), .B(n6316), .S0(n4015), .Y(n6318) );
  NAND4BX1 U6050 ( .AN(n6306), .B(n6305), .C(n6304), .D(n6303), .Y(n6317) );
  OAI222XL U6051 ( .A0(n6550), .A1(n6269), .B0(n2796), .B1(n5331), .C0(n6610), 
        .C1(n5330), .Y(n5333) );
  CLKMX2X2 U6052 ( .A(n6185), .B(n6184), .S0(n4014), .Y(n6186) );
  CLKBUFX3 U6053 ( .A(n7048), .Y(n3165) );
  CLKMX2X2 U6054 ( .A(n5316), .B(n5315), .S0(n4014), .Y(n5317) );
  CLKMX2X2 U6055 ( .A(n6524), .B(n6523), .S0(n4014), .Y(n6525) );
  CLKINVX1 U6056 ( .A(\D_cache/n214 ), .Y(n3975) );
  CLKBUFX3 U6057 ( .A(n2156), .Y(n3396) );
  CLKBUFX3 U6058 ( .A(n2798), .Y(n3486) );
  CLKBUFX3 U6059 ( .A(n2797), .Y(n3308) );
  CLKBUFX3 U6060 ( .A(n8114), .Y(n3442) );
  CLKBUFX3 U6061 ( .A(n2798), .Y(n3487) );
  CLKBUFX3 U6062 ( .A(n2797), .Y(n3309) );
  CLKBUFX3 U6063 ( .A(n2156), .Y(n3397) );
  CLKBUFX3 U6064 ( .A(n2800), .Y(n3530) );
  CLKBUFX3 U6065 ( .A(n2800), .Y(n3531) );
  OAI221X1 U6066 ( .A0(\i_MIPS/n362 ), .A1(n3091), .B0(\i_MIPS/n361 ), .B1(
        n3086), .C0(n4818), .Y(n5960) );
  OA22X1 U6067 ( .A0(\i_MIPS/n360 ), .A1(n3082), .B0(\i_MIPS/n359 ), .B1(n3078), .Y(n4818) );
  OAI221X1 U6068 ( .A0(\i_MIPS/n364 ), .A1(n14), .B0(\i_MIPS/n363 ), .B1(n3077), .C0(n4840), .Y(n5973) );
  OAI221X1 U6069 ( .A0(\i_MIPS/n361 ), .A1(n14), .B0(\i_MIPS/n360 ), .B1(n3077), .C0(n4714), .Y(n6836) );
  OA22X2 U6070 ( .A0(n3634), .A1(n8827), .B0(n3037), .B1(n3977), .Y(
        \D_cache/n240 ) );
  OA22X2 U6071 ( .A0(n8715), .A1(n8826), .B0(n1621), .B1(n3977), .Y(
        \D_cache/n239 ) );
  OA22X2 U6072 ( .A0(n3634), .A1(n8810), .B0(n1616), .B1(n3978), .Y(
        \D_cache/n222 ) );
  OA22X2 U6073 ( .A0(n3634), .A1(n2751), .B0(n8722), .B1(n3978), .Y(
        \D_cache/n224 ) );
  OA22X2 U6074 ( .A0(n3634), .A1(n8812), .B0(n1084), .B1(n3978), .Y(
        \D_cache/n225 ) );
  OA22X2 U6075 ( .A0(n3634), .A1(n8813), .B0(n1618), .B1(n3978), .Y(
        \D_cache/n226 ) );
  OA22X2 U6076 ( .A0(n3634), .A1(n8816), .B0(n1619), .B1(n3978), .Y(
        \D_cache/n229 ) );
  OA22X2 U6077 ( .A0(n3634), .A1(n8820), .B0(n1617), .B1(n3977), .Y(
        \D_cache/n233 ) );
  OA22X2 U6078 ( .A0(n8715), .A1(n8821), .B0(n1620), .B1(n3977), .Y(
        \D_cache/n234 ) );
  OA22X2 U6079 ( .A0(n3634), .A1(n8824), .B0(n1085), .B1(n3977), .Y(
        \D_cache/n237 ) );
  OA22X2 U6080 ( .A0(n3634), .A1(n8832), .B0(n2703), .B1(n3977), .Y(
        \D_cache/n245 ) );
  OAI221X1 U6081 ( .A0(n5381), .A1(n3091), .B0(\i_MIPS/n368 ), .B1(n3085), 
        .C0(n5380), .Y(n5813) );
  OAI221X1 U6082 ( .A0(\i_MIPS/n367 ), .A1(n3092), .B0(\i_MIPS/n366 ), .B1(
        n3087), .C0(n4715), .Y(n5266) );
  OA22X1 U6083 ( .A0(\i_MIPS/n365 ), .A1(n3082), .B0(\i_MIPS/n364 ), .B1(n3078), .Y(n4715) );
  OA21X2 U6084 ( .A0(n3949), .A1(\D_cache/n216 ), .B0(\D_cache/n217 ), .Y(
        \D_cache/n215 ) );
  OAI21XL U6085 ( .A0(\D_cache/n218 ), .A1(n8807), .B0(\D_cache/N31 ), .Y(
        \D_cache/n217 ) );
  OAI222XL U6086 ( .A0(n3584), .A1(n59), .B0(n3648), .B1(n3583), .C0(n3688), 
        .C1(\i_MIPS/n194 ), .Y(n8790) );
  NAND2X1 U6087 ( .A(n55), .B(n3076), .Y(n6332) );
  OAI222XL U6088 ( .A0(n3584), .A1(n60), .B0(n3680), .B1(n3583), .C0(n3688), 
        .C1(\i_MIPS/n191 ), .Y(n8793) );
  OAI221XL U6089 ( .A0(n3068), .A1(n5462), .B0(n3069), .B1(n5481), .C0(n5964), 
        .Y(n6200) );
  OAI221XL U6090 ( .A0(\i_MIPS/n370 ), .A1(n3091), .B0(n5381), .B1(n3086), 
        .C0(n4819), .Y(n5972) );
  OAI221XL U6091 ( .A0(\i_MIPS/n360 ), .A1(n3091), .B0(\i_MIPS/n359 ), .B1(
        n3085), .C0(n5745), .Y(n6331) );
  NAND4X1 U6092 ( .A(n4392), .B(n4391), .C(n4390), .D(n4389), .Y(n8392) );
  OA22X1 U6093 ( .A0(n3304), .A1(n172), .B0(n3258), .B1(n1402), .Y(n4392) );
  OA22X1 U6094 ( .A0(n3483), .A1(n173), .B0(n3408), .B1(n1403), .Y(n4390) );
  OA22X1 U6095 ( .A0(n3392), .A1(n174), .B0(n3350), .B1(n1404), .Y(n4391) );
  OAI222XL U6096 ( .A0(n3585), .A1(n64), .B0(n3661), .B1(n3582), .C0(n3689), 
        .C1(\i_MIPS/n198 ), .Y(n8786) );
  OAI222XL U6097 ( .A0(n3584), .A1(n200), .B0(n3663), .B1(n3583), .C0(n3689), 
        .C1(\i_MIPS/n182 ), .Y(n8802) );
  OAI222XL U6098 ( .A0(n3584), .A1(n196), .B0(n3687), .B1(n3583), .C0(n3689), 
        .C1(\i_MIPS/n188 ), .Y(n8796) );
  OAI222XL U6099 ( .A0(n3585), .A1(n63), .B0(n3658), .B1(n3582), .C0(n3689), 
        .C1(\i_MIPS/n196 ), .Y(n8788) );
  NAND4X1 U6100 ( .A(n7168), .B(n7167), .C(n7166), .D(n7165), .Y(n8676) );
  OA22X1 U6101 ( .A0(n3288), .A1(n695), .B0(n3259), .B1(n1628), .Y(n7168) );
  OA22X1 U6102 ( .A0(n3465), .A1(n696), .B0(n3417), .B1(n1629), .Y(n7166) );
  OA22X1 U6103 ( .A0(n3388), .A1(n697), .B0(n3333), .B1(n1630), .Y(n7167) );
  NAND4X1 U6104 ( .A(n7183), .B(n7182), .C(n7181), .D(n7180), .Y(n8612) );
  OA22X1 U6105 ( .A0(n3287), .A1(n698), .B0(n3259), .B1(n1631), .Y(n7183) );
  OA22X1 U6106 ( .A0(n3465), .A1(n699), .B0(n3417), .B1(n1632), .Y(n7181) );
  OA22X1 U6107 ( .A0(n3375), .A1(n700), .B0(n3333), .B1(n1633), .Y(n7182) );
  NAND4X1 U6108 ( .A(n7173), .B(n7172), .C(n7171), .D(n7170), .Y(n8644) );
  OA22X1 U6109 ( .A0(n3291), .A1(n701), .B0(n3259), .B1(n1634), .Y(n7173) );
  OA22X1 U6110 ( .A0(n3465), .A1(n702), .B0(n3417), .B1(n1635), .Y(n7171) );
  OA22X1 U6111 ( .A0(n3377), .A1(n703), .B0(n3333), .B1(n1636), .Y(n7172) );
  NAND4X1 U6112 ( .A(n7178), .B(n7177), .C(n7176), .D(n7175), .Y(n8580) );
  OA22X1 U6113 ( .A0(n3297), .A1(n704), .B0(n3259), .B1(n1637), .Y(n7178) );
  OA22X1 U6114 ( .A0(n3465), .A1(n705), .B0(n3417), .B1(n1638), .Y(n7176) );
  OA22X1 U6115 ( .A0(n3375), .A1(n706), .B0(n3333), .B1(n1639), .Y(n7177) );
  NAND4X1 U6116 ( .A(n7240), .B(n7239), .C(n7238), .D(n7237), .Y(n8679) );
  OA22X1 U6117 ( .A0(n3288), .A1(n707), .B0(n3244), .B1(n1640), .Y(n7240) );
  OA22X1 U6118 ( .A0(n3466), .A1(n708), .B0(n3418), .B1(n1641), .Y(n7238) );
  OA22X1 U6119 ( .A0(n3383), .A1(n709), .B0(n3333), .B1(n1642), .Y(n7239) );
  NAND4X1 U6120 ( .A(n7250), .B(n7249), .C(n7248), .D(n7247), .Y(n8583) );
  OA22X1 U6121 ( .A0(n3288), .A1(n710), .B0(n3259), .B1(n1643), .Y(n7250) );
  OA22X1 U6122 ( .A0(n3466), .A1(n711), .B0(n3418), .B1(n1644), .Y(n7248) );
  OA22X1 U6123 ( .A0(n3378), .A1(n712), .B0(n3333), .B1(n1645), .Y(n7249) );
  NAND4X1 U6124 ( .A(n7255), .B(n7254), .C(n7253), .D(n7252), .Y(n8615) );
  OA22X1 U6125 ( .A0(n3288), .A1(n713), .B0(n3259), .B1(n1646), .Y(n7255) );
  OA22X1 U6126 ( .A0(n3466), .A1(n714), .B0(n3418), .B1(n1647), .Y(n7253) );
  OA22X1 U6127 ( .A0(n3384), .A1(n715), .B0(n3333), .B1(n1648), .Y(n7254) );
  NAND4X1 U6128 ( .A(n7245), .B(n7244), .C(n7243), .D(n7242), .Y(n8647) );
  OA22X1 U6129 ( .A0(n3288), .A1(n716), .B0(n3259), .B1(n1649), .Y(n7245) );
  OA22X1 U6130 ( .A0(n3466), .A1(n717), .B0(n3418), .B1(n1650), .Y(n7243) );
  OA22X1 U6131 ( .A0(n3388), .A1(n718), .B0(n3333), .B1(n1651), .Y(n7244) );
  NAND4X1 U6132 ( .A(n7288), .B(n7287), .C(n7286), .D(n7285), .Y(n8681) );
  OA22X1 U6133 ( .A0(n3288), .A1(n719), .B0(n3244), .B1(n1652), .Y(n7288) );
  OA22X1 U6134 ( .A0(n3466), .A1(n720), .B0(n3419), .B1(n1653), .Y(n7286) );
  OA22X1 U6135 ( .A0(n3384), .A1(n721), .B0(n3333), .B1(n1654), .Y(n7287) );
  NAND4X1 U6136 ( .A(n7296), .B(n7295), .C(n7294), .D(n7293), .Y(n8585) );
  OA22X1 U6137 ( .A0(n3288), .A1(n722), .B0(n3244), .B1(n1655), .Y(n7296) );
  OA22X1 U6138 ( .A0(n3465), .A1(n723), .B0(n3419), .B1(n1656), .Y(n7294) );
  OA22X1 U6139 ( .A0(n3376), .A1(n724), .B0(n3333), .B1(n1657), .Y(n7295) );
  NAND4X1 U6140 ( .A(n7300), .B(n7299), .C(n7298), .D(n7297), .Y(n8617) );
  NAND4X1 U6141 ( .A(n7292), .B(n7291), .C(n7290), .D(n7289), .Y(n8649) );
  OA22X1 U6142 ( .A0(n3288), .A1(n725), .B0(n3244), .B1(n1658), .Y(n7292) );
  OA22X1 U6143 ( .A0(n3466), .A1(n726), .B0(n3419), .B1(n1659), .Y(n7290) );
  OA22X1 U6144 ( .A0(n3387), .A1(n727), .B0(n3333), .B1(n1660), .Y(n7291) );
  NAND4X1 U6145 ( .A(n7264), .B(n7263), .C(n7262), .D(n7261), .Y(n8680) );
  OA22X1 U6146 ( .A0(n3288), .A1(n728), .B0(n3240), .B1(n1661), .Y(n7264) );
  OA22X1 U6147 ( .A0(n3466), .A1(n729), .B0(n3418), .B1(n1662), .Y(n7262) );
  OA22X1 U6148 ( .A0(n3378), .A1(n730), .B0(n3332), .B1(n1663), .Y(n7263) );
  NAND4X1 U6149 ( .A(n7274), .B(n7273), .C(n7272), .D(n7271), .Y(n8584) );
  OA22X1 U6150 ( .A0(n3288), .A1(n731), .B0(n3250), .B1(n1664), .Y(n7274) );
  OA22X1 U6151 ( .A0(n3466), .A1(n732), .B0(n3419), .B1(n1665), .Y(n7272) );
  OA22X1 U6152 ( .A0(n3379), .A1(n733), .B0(n3333), .B1(n1666), .Y(n7273) );
  NAND4X1 U6153 ( .A(n7279), .B(n7278), .C(n7277), .D(n7276), .Y(n8616) );
  OA22X1 U6154 ( .A0(n3288), .A1(n734), .B0(n3244), .B1(n1667), .Y(n7279) );
  OA22X1 U6155 ( .A0(n3466), .A1(n735), .B0(n3419), .B1(n1668), .Y(n7277) );
  OA22X1 U6156 ( .A0(n3375), .A1(n736), .B0(n3333), .B1(n1669), .Y(n7278) );
  NAND4X1 U6157 ( .A(n7269), .B(n7268), .C(n7267), .D(n7266), .Y(n8648) );
  OA22X1 U6158 ( .A0(n3300), .A1(n737), .B0(n3244), .B1(n1670), .Y(n7269) );
  OA22X1 U6159 ( .A0(n3466), .A1(n738), .B0(n3419), .B1(n1671), .Y(n7267) );
  OA22X1 U6160 ( .A0(n3377), .A1(n739), .B0(n3333), .B1(n1672), .Y(n7268) );
  NAND4X1 U6161 ( .A(n7216), .B(n7215), .C(n7214), .D(n7213), .Y(n8678) );
  OA22X1 U6162 ( .A0(n3289), .A1(n740), .B0(n3259), .B1(n1673), .Y(n7216) );
  OA22X1 U6163 ( .A0(n3466), .A1(n741), .B0(n3419), .B1(n1674), .Y(n7214) );
  OA22X1 U6164 ( .A0(n3387), .A1(n742), .B0(n3333), .B1(n1675), .Y(n7215) );
  NAND4X1 U6165 ( .A(n7231), .B(n7230), .C(n7229), .D(n7228), .Y(n8614) );
  OA22X1 U6166 ( .A0(n3288), .A1(n743), .B0(n3250), .B1(n1676), .Y(n7231) );
  OA22X1 U6167 ( .A0(n3466), .A1(n744), .B0(n3418), .B1(n1677), .Y(n7229) );
  OA22X1 U6168 ( .A0(n3383), .A1(n745), .B0(n3338), .B1(n1678), .Y(n7230) );
  NAND4X1 U6169 ( .A(n7221), .B(n7220), .C(n7219), .D(n7218), .Y(n8646) );
  OA22X1 U6170 ( .A0(n3292), .A1(n746), .B0(n3259), .B1(n1679), .Y(n7221) );
  OA22X1 U6171 ( .A0(n3466), .A1(n747), .B0(n3419), .B1(n1680), .Y(n7219) );
  OA22X1 U6172 ( .A0(n3375), .A1(n748), .B0(n3333), .B1(n1681), .Y(n7220) );
  NAND4X1 U6173 ( .A(n7226), .B(n7225), .C(n7224), .D(n7223), .Y(n8582) );
  OA22X1 U6174 ( .A0(n3297), .A1(n749), .B0(n3259), .B1(n1682), .Y(n7226) );
  OA22X1 U6175 ( .A0(n3466), .A1(n750), .B0(n3419), .B1(n1683), .Y(n7224) );
  OA22X1 U6176 ( .A0(n3376), .A1(n751), .B0(n3333), .B1(n1684), .Y(n7225) );
  NAND4X1 U6177 ( .A(n7192), .B(n7191), .C(n7190), .D(n7189), .Y(n8677) );
  OA22X1 U6178 ( .A0(n3288), .A1(n752), .B0(n3241), .B1(n1685), .Y(n7192) );
  OA22X1 U6179 ( .A0(n3465), .A1(n753), .B0(n3417), .B1(n1686), .Y(n7190) );
  OA22X1 U6180 ( .A0(n3383), .A1(n754), .B0(n3332), .B1(n1687), .Y(n7191) );
  NAND4X1 U6181 ( .A(n7207), .B(n7206), .C(n7205), .D(n7204), .Y(n8613) );
  OA22X1 U6182 ( .A0(n3298), .A1(n755), .B0(n3259), .B1(n1688), .Y(n7207) );
  OA22X1 U6183 ( .A0(n3466), .A1(n756), .B0(n3419), .B1(n1689), .Y(n7205) );
  OA22X1 U6184 ( .A0(n3380), .A1(n757), .B0(n3333), .B1(n1690), .Y(n7206) );
  NAND4X1 U6185 ( .A(n7197), .B(n7196), .C(n7195), .D(n7194), .Y(n8645) );
  OA22X1 U6186 ( .A0(n3287), .A1(n758), .B0(n3259), .B1(n1691), .Y(n7197) );
  OA22X1 U6187 ( .A0(n3466), .A1(n759), .B0(n3419), .B1(n1692), .Y(n7195) );
  OA22X1 U6188 ( .A0(n3388), .A1(n760), .B0(n3333), .B1(n1693), .Y(n7196) );
  NAND4X1 U6189 ( .A(n7202), .B(n7201), .C(n7200), .D(n7199), .Y(n8581) );
  OA22X1 U6190 ( .A0(n3301), .A1(n761), .B0(n3259), .B1(n1694), .Y(n7202) );
  OA22X1 U6191 ( .A0(n3466), .A1(n762), .B0(n3419), .B1(n1695), .Y(n7200) );
  OA22X1 U6192 ( .A0(n3383), .A1(n763), .B0(n3333), .B1(n1696), .Y(n7201) );
  NAND4X1 U6193 ( .A(n7418), .B(n7417), .C(n7416), .D(n7415), .Y(n8674) );
  NAND4X1 U6194 ( .A(n7428), .B(n7427), .C(n7426), .D(n7425), .Y(n8578) );
  NAND4X1 U6195 ( .A(n7433), .B(n7432), .C(n7431), .D(n7430), .Y(n8610) );
  NAND4X1 U6196 ( .A(n7423), .B(n7422), .C(n7421), .D(n7420), .Y(n8642) );
  NAND4X1 U6197 ( .A(n7500), .B(n7499), .C(n7498), .D(n7497), .Y(n8574) );
  NAND4X1 U6198 ( .A(n7490), .B(n7489), .C(n7488), .D(n7487), .Y(n8670) );
  NAND4X1 U6199 ( .A(n7505), .B(n7504), .C(n7503), .D(n7502), .Y(n8606) );
  NAND4X1 U6200 ( .A(n7495), .B(n7494), .C(n7493), .D(n7492), .Y(n8638) );
  NAND4X1 U6201 ( .A(n7134), .B(n7133), .C(n7132), .D(n7131), .Y(n8605) );
  OA22X1 U6202 ( .A0(n3288), .A1(n764), .B0(n3241), .B1(n1697), .Y(n7134) );
  OA22X1 U6203 ( .A0(n3464), .A1(n765), .B0(n3419), .B1(n1698), .Y(n7132) );
  OA22X1 U6204 ( .A0(n3380), .A1(n766), .B0(n3345), .B1(n1699), .Y(n7133) );
  NAND4X1 U6205 ( .A(n7124), .B(n7123), .C(n7122), .D(n7121), .Y(n8637) );
  OA22X1 U6206 ( .A0(n3288), .A1(n767), .B0(n3241), .B1(n1700), .Y(n7124) );
  OA22X1 U6207 ( .A0(n3464), .A1(n768), .B0(n3419), .B1(n1701), .Y(n7122) );
  OA22X1 U6208 ( .A0(n3376), .A1(n769), .B0(n3332), .B1(n1702), .Y(n7123) );
  NAND4X1 U6209 ( .A(n7129), .B(n7128), .C(n7127), .D(n7126), .Y(n8573) );
  OA22X1 U6210 ( .A0(n3301), .A1(n770), .B0(n3241), .B1(n1703), .Y(n7129) );
  OA22X1 U6211 ( .A0(n3466), .A1(n771), .B0(n3417), .B1(n1704), .Y(n7127) );
  OA22X1 U6212 ( .A0(n3392), .A1(n772), .B0(n3338), .B1(n1705), .Y(n7128) );
  NAND4X1 U6213 ( .A(n7119), .B(n7118), .C(n7117), .D(n7116), .Y(n8669) );
  OA22X1 U6214 ( .A0(n3287), .A1(n1848), .B0(n3241), .B1(n914), .Y(n7119) );
  OA22X1 U6215 ( .A0(n3469), .A1(n773), .B0(n3419), .B1(n1706), .Y(n7117) );
  OA22X1 U6216 ( .A0(n3391), .A1(n1849), .B0(n3346), .B1(n915), .Y(n7118) );
  NAND4X1 U6217 ( .A(n7650), .B(n7649), .C(n7648), .D(n7647), .Y(n8579) );
  NAND4X1 U6218 ( .A(n7640), .B(n7639), .C(n7638), .D(n7637), .Y(n8675) );
  NAND4X1 U6219 ( .A(n7655), .B(n7654), .C(n7653), .D(n7652), .Y(n8611) );
  NAND4X1 U6220 ( .A(n7645), .B(n7644), .C(n7643), .D(n7642), .Y(n8643) );
  NAND4X1 U6221 ( .A(n7442), .B(n7441), .C(n7440), .D(n7439), .Y(n8673) );
  NAND4X1 U6222 ( .A(n7452), .B(n7451), .C(n7450), .D(n7449), .Y(n8577) );
  OA22X1 U6223 ( .A0(n3288), .A1(n774), .B0(n3241), .B1(n1707), .Y(n7452) );
  OA22X1 U6224 ( .A0(n3469), .A1(n775), .B0(n3418), .B1(n1708), .Y(n7450) );
  OA22X1 U6225 ( .A0(n3379), .A1(n776), .B0(n3338), .B1(n1709), .Y(n7451) );
  NAND4X1 U6226 ( .A(n7457), .B(n7456), .C(n7455), .D(n7454), .Y(n8609) );
  OA22X1 U6227 ( .A0(n3291), .A1(n777), .B0(n3241), .B1(n1710), .Y(n7457) );
  OA22X1 U6228 ( .A0(n3469), .A1(n778), .B0(n3419), .B1(n1711), .Y(n7455) );
  OA22X1 U6229 ( .A0(n3380), .A1(n779), .B0(n3333), .B1(n1712), .Y(n7456) );
  NAND4X1 U6230 ( .A(n7447), .B(n7446), .C(n7445), .D(n7444), .Y(n8641) );
  OA22X1 U6231 ( .A0(n3293), .A1(n1850), .B0(n3241), .B1(n916), .Y(n7447) );
  OA22X1 U6232 ( .A0(n3464), .A1(n780), .B0(n3418), .B1(n1713), .Y(n7445) );
  OA22X1 U6233 ( .A0(n3375), .A1(n781), .B0(n3343), .B1(n1714), .Y(n7446) );
  NAND4X1 U6234 ( .A(n7476), .B(n7475), .C(n7474), .D(n7473), .Y(n8575) );
  OA22X1 U6235 ( .A0(n3288), .A1(n782), .B0(n3241), .B1(n1715), .Y(n7476) );
  OA22X1 U6236 ( .A0(n3469), .A1(n783), .B0(n3419), .B1(n1716), .Y(n7474) );
  OA22X1 U6237 ( .A0(n3386), .A1(n784), .B0(n3332), .B1(n1717), .Y(n7475) );
  NAND4X1 U6238 ( .A(n7466), .B(n7465), .C(n7464), .D(n7463), .Y(n8671) );
  OA22X1 U6239 ( .A0(n3293), .A1(n1851), .B0(n3241), .B1(n917), .Y(n7466) );
  OA22X1 U6240 ( .A0(n3465), .A1(n785), .B0(n3418), .B1(n1718), .Y(n7464) );
  OA22X1 U6241 ( .A0(n3377), .A1(n1852), .B0(n3332), .B1(n918), .Y(n7465) );
  NAND4X1 U6242 ( .A(n7481), .B(n7480), .C(n7479), .D(n7478), .Y(n8607) );
  NAND4X1 U6243 ( .A(n7471), .B(n7470), .C(n7469), .D(n7468), .Y(n8639) );
  OA22X1 U6244 ( .A0(n3287), .A1(n1853), .B0(n3241), .B1(n919), .Y(n7471) );
  OA22X1 U6245 ( .A0(n3469), .A1(n786), .B0(n3418), .B1(n1719), .Y(n7469) );
  OA22X1 U6246 ( .A0(n3375), .A1(n787), .B0(n3349), .B1(n1720), .Y(n7470) );
  NAND4X1 U6247 ( .A(n7158), .B(n7157), .C(n7156), .D(n7155), .Y(n8604) );
  OA22X1 U6248 ( .A0(n3288), .A1(n788), .B0(n3241), .B1(n1721), .Y(n7158) );
  OA22X1 U6249 ( .A0(n3465), .A1(n789), .B0(n3417), .B1(n1722), .Y(n7156) );
  OA22X1 U6250 ( .A0(n3389), .A1(n790), .B0(n3332), .B1(n1723), .Y(n7157) );
  NAND4X1 U6251 ( .A(n7148), .B(n7147), .C(n7146), .D(n7145), .Y(n8636) );
  OA22X1 U6252 ( .A0(n3288), .A1(n791), .B0(n3241), .B1(n1724), .Y(n7148) );
  OA22X1 U6253 ( .A0(n3469), .A1(n792), .B0(n3419), .B1(n1725), .Y(n7146) );
  OA22X1 U6254 ( .A0(n3375), .A1(n793), .B0(n3338), .B1(n1726), .Y(n7147) );
  NAND4X1 U6255 ( .A(n7153), .B(n7152), .C(n7151), .D(n7150), .Y(n8572) );
  OA22X1 U6256 ( .A0(n3300), .A1(n794), .B0(n3241), .B1(n1727), .Y(n7153) );
  OA22X1 U6257 ( .A0(n3469), .A1(n795), .B0(n3419), .B1(n1728), .Y(n7151) );
  OA22X1 U6258 ( .A0(n3387), .A1(n796), .B0(n3332), .B1(n1729), .Y(n7152) );
  NAND4X1 U6259 ( .A(n7143), .B(n7142), .C(n7141), .D(n7140), .Y(n8668) );
  OA22X1 U6260 ( .A0(n3293), .A1(n1854), .B0(n3241), .B1(n920), .Y(n7143) );
  OA22X1 U6261 ( .A0(n3464), .A1(n797), .B0(n3418), .B1(n1730), .Y(n7141) );
  OA22X1 U6262 ( .A0(n3380), .A1(n1855), .B0(n3334), .B1(n921), .Y(n7142) );
  NAND4X1 U6263 ( .A(n4582), .B(n4581), .C(n4580), .D(n4579), .Y(n8571) );
  NAND4X1 U6264 ( .A(n4572), .B(n4571), .C(n4570), .D(n4569), .Y(n8667) );
  NAND4X1 U6265 ( .A(n4587), .B(n4586), .C(n4585), .D(n4584), .Y(n8603) );
  OA22X1 U6266 ( .A0(n3288), .A1(n798), .B0(n3241), .B1(n1731), .Y(n4587) );
  OA22X1 U6267 ( .A0(n3469), .A1(n799), .B0(n3418), .B1(n1732), .Y(n4585) );
  OA22X1 U6268 ( .A0(n3384), .A1(n800), .B0(n3346), .B1(n1733), .Y(n4586) );
  NAND4X1 U6269 ( .A(n4577), .B(n4576), .C(n4575), .D(n4574), .Y(n8635) );
  NAND4X1 U6270 ( .A(n7110), .B(n7109), .C(n7108), .D(n7107), .Y(n8602) );
  OA22X1 U6271 ( .A0(n3293), .A1(n801), .B0(n3241), .B1(n1734), .Y(n7110) );
  OA22X1 U6272 ( .A0(n3466), .A1(n802), .B0(n3418), .B1(n1735), .Y(n7108) );
  OA22X1 U6273 ( .A0(n3384), .A1(n803), .B0(n3337), .B1(n1736), .Y(n7109) );
  NAND4X1 U6274 ( .A(n7100), .B(n7099), .C(n7098), .D(n7097), .Y(n8634) );
  OA22X1 U6275 ( .A0(n3288), .A1(n804), .B0(n3241), .B1(n1737), .Y(n7100) );
  OA22X1 U6276 ( .A0(n3466), .A1(n805), .B0(n3419), .B1(n1738), .Y(n7098) );
  OA22X1 U6277 ( .A0(n3380), .A1(n806), .B0(n3336), .B1(n1739), .Y(n7099) );
  NAND4X1 U6278 ( .A(n7105), .B(n7104), .C(n7103), .D(n7102), .Y(n8570) );
  OA22X1 U6279 ( .A0(n3298), .A1(n807), .B0(n3241), .B1(n1740), .Y(n7105) );
  OA22X1 U6280 ( .A0(n3464), .A1(n808), .B0(n3418), .B1(n1741), .Y(n7103) );
  OA22X1 U6281 ( .A0(n3385), .A1(n809), .B0(n3338), .B1(n1742), .Y(n7104) );
  NAND4X1 U6282 ( .A(n7095), .B(n7094), .C(n7093), .D(n7092), .Y(n8666) );
  OA22X1 U6283 ( .A0(n3287), .A1(n1856), .B0(n3241), .B1(n922), .Y(n7095) );
  OA22X1 U6284 ( .A0(n3469), .A1(n810), .B0(n3419), .B1(n1743), .Y(n7093) );
  OA22X1 U6285 ( .A0(n3375), .A1(n1857), .B0(n3345), .B1(n923), .Y(n7094) );
  NAND4X1 U6286 ( .A(n7350), .B(n7349), .C(n7348), .D(n7347), .Y(n8652) );
  NAND4X1 U6287 ( .A(n7358), .B(n7357), .C(n7356), .D(n7355), .Y(n8556) );
  NAND4X1 U6288 ( .A(n7362), .B(n7361), .C(n7360), .D(n7359), .Y(n8588) );
  NAND4X1 U6289 ( .A(n7354), .B(n7353), .C(n7352), .D(n7351), .Y(n8620) );
  NAND4X1 U6290 ( .A(n7338), .B(n7337), .C(n7336), .D(n7335), .Y(n8558) );
  NAND4X1 U6291 ( .A(n4547), .B(n4546), .C(n4545), .D(n4544), .Y(n8654) );
  OA22X1 U6292 ( .A0(n3374), .A1(n487), .B0(n3331), .B1(n1405), .Y(n4546) );
  OA22X1 U6293 ( .A0(n3287), .A1(n488), .B0(n3239), .B1(n1406), .Y(n4547) );
  NAND4X1 U6294 ( .A(n7342), .B(n7341), .C(n7340), .D(n7339), .Y(n8590) );
  NAND4X1 U6295 ( .A(n7334), .B(n7333), .C(n7332), .D(n7331), .Y(n8622) );
  NAND4X1 U6296 ( .A(n7400), .B(n7399), .C(n7398), .D(n7397), .Y(n8559) );
  NAND4X1 U6297 ( .A(n7390), .B(n7389), .C(n7388), .D(n7387), .Y(n8655) );
  NAND4X1 U6298 ( .A(n7405), .B(n7404), .C(n7403), .D(n7402), .Y(n8591) );
  OA22X1 U6299 ( .A0(n3556), .A1(n489), .B0(n3514), .B1(n1407), .Y(n7402) );
  OA22X1 U6300 ( .A0(n3379), .A1(n490), .B0(n3337), .B1(n1408), .Y(n7404) );
  OA22X1 U6301 ( .A0(n3292), .A1(n491), .B0(n3245), .B1(n1409), .Y(n7405) );
  NAND4X1 U6302 ( .A(n7395), .B(n7394), .C(n7393), .D(n7392), .Y(n8623) );
  OA22X1 U6303 ( .A0(n3564), .A1(n492), .B0(n3522), .B1(n1410), .Y(n7769) );
  OA22X1 U6304 ( .A0(n3387), .A1(n493), .B0(n3345), .B1(n1411), .Y(n7771) );
  NAND4X1 U6305 ( .A(n7776), .B(n7775), .C(n7774), .D(n7773), .Y(n8592) );
  OA22X1 U6306 ( .A0(n3565), .A1(n494), .B0(n3523), .B1(n1412), .Y(n7773) );
  OA22X1 U6307 ( .A0(n3388), .A1(n495), .B0(n3346), .B1(n1413), .Y(n7775) );
  OA22X1 U6308 ( .A0(n3301), .A1(n496), .B0(n3254), .B1(n1414), .Y(n7776) );
  NAND4X1 U6309 ( .A(n7762), .B(n7761), .C(n7760), .D(n7759), .Y(n8656) );
  NAND4X1 U6310 ( .A(n7767), .B(n7766), .C(n7765), .D(n7764), .Y(n8624) );
  OA22X1 U6311 ( .A0(n3564), .A1(n497), .B0(n3522), .B1(n1415), .Y(n7764) );
  OA22X1 U6312 ( .A0(n3387), .A1(n498), .B0(n3345), .B1(n1416), .Y(n7766) );
  OA22X1 U6313 ( .A0(n3300), .A1(n499), .B0(n3253), .B1(n1417), .Y(n7767) );
  NAND4X1 U6314 ( .A(n7748), .B(n7747), .C(n7746), .D(n7745), .Y(n8561) );
  NAND4X1 U6315 ( .A(n7753), .B(n7752), .C(n7751), .D(n7750), .Y(n8593) );
  NAND4X1 U6316 ( .A(n7738), .B(n7737), .C(n7736), .D(n7735), .Y(n8657) );
  NAND4X1 U6317 ( .A(n7743), .B(n7742), .C(n7741), .D(n7740), .Y(n8625) );
  NAND4X1 U6318 ( .A(n7722), .B(n7721), .C(n7720), .D(n7719), .Y(n8562) );
  OA22X1 U6319 ( .A0(n3386), .A1(n500), .B0(n3344), .B1(n1418), .Y(n7721) );
  OA22X1 U6320 ( .A0(n3563), .A1(n501), .B0(n3521), .B1(n1419), .Y(n7719) );
  OA22X1 U6321 ( .A0(n3299), .A1(n502), .B0(n3252), .B1(n1420), .Y(n7722) );
  OA22X1 U6322 ( .A0(n3386), .A1(n503), .B0(n3344), .B1(n1421), .Y(n7726) );
  OA22X1 U6323 ( .A0(n3563), .A1(n504), .B0(n3521), .B1(n1422), .Y(n7724) );
  NAND4X1 U6324 ( .A(n7712), .B(n7711), .C(n7710), .D(n7709), .Y(n8658) );
  NAND4X1 U6325 ( .A(n7717), .B(n7716), .C(n7715), .D(n7714), .Y(n8626) );
  OA22X1 U6326 ( .A0(n3385), .A1(n505), .B0(n3343), .B1(n1423), .Y(n7698) );
  OA22X1 U6327 ( .A0(n3562), .A1(n506), .B0(n3520), .B1(n1424), .Y(n7696) );
  NAND4X1 U6328 ( .A(n7703), .B(n7702), .C(n7701), .D(n7700), .Y(n8595) );
  NAND4X1 U6329 ( .A(n7689), .B(n7688), .C(n7687), .D(n7686), .Y(n8659) );
  NAND4X1 U6330 ( .A(n7694), .B(n7693), .C(n7692), .D(n7691), .Y(n8627) );
  OA22X1 U6331 ( .A0(n3385), .A1(n507), .B0(n3343), .B1(n1425), .Y(n7693) );
  OA22X1 U6332 ( .A0(n3298), .A1(n508), .B0(n3251), .B1(n1426), .Y(n7694) );
  OA22X1 U6333 ( .A0(n3562), .A1(n509), .B0(n3520), .B1(n1427), .Y(n7691) );
  NAND4X1 U6334 ( .A(n7675), .B(n7674), .C(n7673), .D(n7672), .Y(n8564) );
  NAND4X1 U6335 ( .A(n7680), .B(n7679), .C(n7678), .D(n7677), .Y(n8596) );
  NAND4X1 U6336 ( .A(n7665), .B(n7664), .C(n7663), .D(n7662), .Y(n8660) );
  NAND4X1 U6337 ( .A(n7670), .B(n7669), .C(n7668), .D(n7667), .Y(n8628) );
  NAND4X1 U6338 ( .A(n7597), .B(n7596), .C(n7595), .D(n7594), .Y(n8565) );
  NAND4X1 U6339 ( .A(n7602), .B(n7601), .C(n7600), .D(n7599), .Y(n8597) );
  NAND4X1 U6340 ( .A(n7587), .B(n7586), .C(n7585), .D(n7584), .Y(n8661) );
  NAND4X1 U6341 ( .A(n7592), .B(n7591), .C(n7590), .D(n7589), .Y(n8629) );
  OA22X1 U6342 ( .A0(n3383), .A1(n510), .B0(n3341), .B1(n1428), .Y(n7621) );
  OA22X1 U6343 ( .A0(n3560), .A1(n511), .B0(n3518), .B1(n1429), .Y(n7619) );
  NAND4X1 U6344 ( .A(n7626), .B(n7625), .C(n7624), .D(n7623), .Y(n8598) );
  OA22X1 U6345 ( .A0(n3384), .A1(n512), .B0(n3342), .B1(n1430), .Y(n7625) );
  OA22X1 U6346 ( .A0(n3561), .A1(n513), .B0(n3519), .B1(n1431), .Y(n7623) );
  OA22X1 U6347 ( .A0(n3297), .A1(n514), .B0(n3250), .B1(n1432), .Y(n7626) );
  NAND4X1 U6348 ( .A(n7612), .B(n7611), .C(n7610), .D(n7609), .Y(n8662) );
  NAND4X1 U6349 ( .A(n7617), .B(n7616), .C(n7615), .D(n7614), .Y(n8630) );
  OA22X1 U6350 ( .A0(n3383), .A1(n515), .B0(n3341), .B1(n1433), .Y(n7616) );
  OA22X1 U6351 ( .A0(n3560), .A1(n516), .B0(n3518), .B1(n1434), .Y(n7614) );
  OA22X1 U6352 ( .A0(n3296), .A1(n517), .B0(n3249), .B1(n1435), .Y(n7617) );
  NAND4X1 U6353 ( .A(n7573), .B(n7572), .C(n7571), .D(n7570), .Y(n8567) );
  NAND4X1 U6354 ( .A(n7578), .B(n7577), .C(n7576), .D(n7575), .Y(n8599) );
  NAND4X1 U6355 ( .A(n7563), .B(n7562), .C(n7561), .D(n7560), .Y(n8663) );
  NAND4X1 U6356 ( .A(n7568), .B(n7567), .C(n7566), .D(n7565), .Y(n8631) );
  NAND4X1 U6357 ( .A(n7524), .B(n7523), .C(n7522), .D(n7521), .Y(n8568) );
  NAND4X1 U6358 ( .A(n7529), .B(n7528), .C(n7527), .D(n7526), .Y(n8600) );
  NAND4X1 U6359 ( .A(n7514), .B(n7513), .C(n7512), .D(n7511), .Y(n8664) );
  OA22X1 U6360 ( .A0(n3557), .A1(n518), .B0(n3515), .B1(n1436), .Y(n7511) );
  OA22X1 U6361 ( .A0(n3380), .A1(n519), .B0(n3338), .B1(n1437), .Y(n7513) );
  OA22X1 U6362 ( .A0(n3293), .A1(n520), .B0(n3246), .B1(n1438), .Y(n7514) );
  NAND4X1 U6363 ( .A(n7519), .B(n7518), .C(n7517), .D(n7516), .Y(n8632) );
  NAND2X1 U6364 ( .A(n2986), .B(n4017), .Y(n6907) );
  OAI222XL U6365 ( .A0(n3585), .A1(n198), .B0(n3682), .B1(n3582), .C0(n3689), 
        .C1(\i_MIPS/n190 ), .Y(n8794) );
  OAI222XL U6366 ( .A0(n3584), .A1(n57), .B0(n3664), .B1(n3583), .C0(n3688), 
        .C1(\i_MIPS/n189 ), .Y(n8795) );
  OAI222XL U6367 ( .A0(n3584), .A1(n201), .B0(n3669), .B1(n3583), .C0(n3688), 
        .C1(\i_MIPS/n183 ), .Y(n8801) );
  OAI222XL U6368 ( .A0(n3584), .A1(n203), .B0(n3660), .B1(n3583), .C0(n3689), 
        .C1(\i_MIPS/n203 ), .Y(n8781) );
  OAI222XL U6369 ( .A0(n3584), .A1(n202), .B0(n3017), .B1(n3583), .C0(n3689), 
        .C1(\i_MIPS/n202 ), .Y(n8782) );
  OAI222XL U6370 ( .A0(n3584), .A1(n204), .B0(n8744), .B1(n3582), .C0(n3689), 
        .C1(\i_MIPS/n200 ), .Y(n8784) );
  OAI222XL U6371 ( .A0(n3585), .A1(n65), .B0(n27), .B1(n8333), .C0(n3688), 
        .C1(\i_MIPS/n197 ), .Y(n8787) );
  OAI222XL U6372 ( .A0(n3584), .A1(n197), .B0(n3668), .B1(n3583), .C0(n3689), 
        .C1(\i_MIPS/n184 ), .Y(n8800) );
  NAND2X1 U6373 ( .A(n2985), .B(n1082), .Y(n6847) );
  NAND2X1 U6374 ( .A(n4628), .B(\i_MIPS/n346 ), .Y(n6061) );
  NAND2X1 U6375 ( .A(n4636), .B(\i_MIPS/n348 ), .Y(n6837) );
  NOR4X1 U6376 ( .A(n6179), .B(n6178), .C(n6177), .D(n6176), .Y(n6180) );
  AO22X1 U6377 ( .A0(n3194), .A1(n196), .B0(n3190), .B1(n1093), .Y(n6179) );
  AO22X1 U6378 ( .A0(n3200), .A1(n210), .B0(n3196), .B1(n1094), .Y(n6178) );
  AO22X1 U6379 ( .A0(n3204), .A1(n211), .B0(n3203), .B1(n1095), .Y(n6177) );
  NOR4X1 U6380 ( .A(n6170), .B(n6169), .C(n6168), .D(n6167), .Y(n6171) );
  AO22X1 U6381 ( .A0(n3194), .A1(n1107), .B0(n3190), .B1(n222), .Y(n6170) );
  AO22X1 U6382 ( .A0(n3200), .A1(n212), .B0(n3196), .B1(n1096), .Y(n6169) );
  AO22X1 U6383 ( .A0(n190), .A1(n213), .B0(n3203), .B1(n1097), .Y(n6168) );
  NOR4X1 U6384 ( .A(n5310), .B(n5309), .C(n5308), .D(n5307), .Y(n5311) );
  AO22X1 U6385 ( .A0(n3192), .A1(n60), .B0(n3188), .B1(n1137), .Y(n5310) );
  AO22X1 U6386 ( .A0(n3198), .A1(n249), .B0(n192), .B1(n1138), .Y(n5309) );
  AO22X1 U6387 ( .A0(n3205), .A1(n1109), .B0(n3201), .B1(n224), .Y(n5308) );
  NOR4X1 U6388 ( .A(n5301), .B(n5300), .C(n5299), .D(n5298), .Y(n5302) );
  AO22X1 U6389 ( .A0(n3192), .A1(n250), .B0(n3188), .B1(n1139), .Y(n5301) );
  AO22X1 U6390 ( .A0(n3198), .A1(n251), .B0(n192), .B1(n1140), .Y(n5300) );
  AO22X1 U6391 ( .A0(n3205), .A1(n1110), .B0(n3201), .B1(n225), .Y(n5299) );
  NOR4X1 U6392 ( .A(n6311), .B(n6310), .C(n6309), .D(n6308), .Y(n6312) );
  AO22X1 U6393 ( .A0(n3194), .A1(n209), .B0(n3190), .B1(n1113), .Y(n6311) );
  AO22X1 U6394 ( .A0(n3200), .A1(n229), .B0(n3196), .B1(n1114), .Y(n6310) );
  AO22X1 U6395 ( .A0(n190), .A1(n230), .B0(n3203), .B1(n1115), .Y(n6309) );
  NOR4X1 U6396 ( .A(n6302), .B(n6301), .C(n6300), .D(n6299), .Y(n6303) );
  AO22X1 U6397 ( .A0(n3194), .A1(n231), .B0(n3190), .B1(n1116), .Y(n6302) );
  AO22X1 U6398 ( .A0(n3200), .A1(n232), .B0(n3196), .B1(n1117), .Y(n6301) );
  AO22X1 U6399 ( .A0(n190), .A1(n233), .B0(n3203), .B1(n1118), .Y(n6300) );
  NOR4X1 U6400 ( .A(n6290), .B(n6289), .C(n6288), .D(n6287), .Y(n6291) );
  AO22X1 U6401 ( .A0(n3141), .A1(n209), .B0(n3138), .B1(n1113), .Y(n6290) );
  AO22X1 U6402 ( .A0(n3147), .A1(n229), .B0(n3144), .B1(n1114), .Y(n6289) );
  AO22X1 U6403 ( .A0(n3153), .A1(n230), .B0(n3150), .B1(n1115), .Y(n6288) );
  NOR4X1 U6404 ( .A(n6281), .B(n6280), .C(n6279), .D(n6278), .Y(n6282) );
  AO22X1 U6405 ( .A0(n3141), .A1(n231), .B0(n3138), .B1(n1116), .Y(n6281) );
  AO22X1 U6406 ( .A0(n3147), .A1(n232), .B0(n3144), .B1(n1117), .Y(n6280) );
  AO22X1 U6407 ( .A0(n3153), .A1(n233), .B0(n3150), .B1(n1118), .Y(n6279) );
  NOR4X1 U6408 ( .A(n6446), .B(n6445), .C(n6444), .D(n6443), .Y(n6447) );
  AO22X1 U6409 ( .A0(n3194), .A1(n58), .B0(n3190), .B1(n1098), .Y(n6446) );
  AO22X1 U6410 ( .A0(n3200), .A1(n214), .B0(n3196), .B1(n1099), .Y(n6445) );
  AO22X1 U6411 ( .A0(n190), .A1(n215), .B0(n3203), .B1(n1100), .Y(n6444) );
  NOR4X1 U6412 ( .A(n6437), .B(n6436), .C(n6435), .D(n6434), .Y(n6438) );
  AO22X1 U6413 ( .A0(n3194), .A1(n1108), .B0(n3190), .B1(n223), .Y(n6437) );
  AO22X1 U6414 ( .A0(n3200), .A1(n216), .B0(n3196), .B1(n1101), .Y(n6436) );
  AO22X1 U6415 ( .A0(n190), .A1(n217), .B0(n3203), .B1(n1102), .Y(n6435) );
  NOR4X1 U6416 ( .A(n5350), .B(n5349), .C(n5348), .D(n5347), .Y(n5351) );
  AO22X1 U6417 ( .A0(n3141), .A1(n197), .B0(n3137), .B1(n1131), .Y(n5350) );
  AO22X1 U6418 ( .A0(n3147), .A1(n244), .B0(n3143), .B1(n1132), .Y(n5349) );
  AO22X1 U6419 ( .A0(n3153), .A1(n245), .B0(n3149), .B1(n1133), .Y(n5348) );
  NOR4X1 U6420 ( .A(n5341), .B(n5340), .C(n5339), .D(n5338), .Y(n5342) );
  AO22X1 U6421 ( .A0(n3141), .A1(n246), .B0(n3137), .B1(n1134), .Y(n5341) );
  AO22X1 U6422 ( .A0(n3147), .A1(n247), .B0(n3143), .B1(n1135), .Y(n5340) );
  AO22X1 U6423 ( .A0(n3153), .A1(n248), .B0(n3149), .B1(n1136), .Y(n5339) );
  NOR4X1 U6424 ( .A(n5076), .B(n5075), .C(n5074), .D(n5073), .Y(n5077) );
  AO22X1 U6425 ( .A0(n3140), .A1(n70), .B0(n180), .B1(n1171), .Y(n5076) );
  AO22X1 U6426 ( .A0(n3146), .A1(n277), .B0(n184), .B1(n1172), .Y(n5075) );
  AO22X1 U6427 ( .A0(n3152), .A1(n278), .B0(n182), .B1(n1173), .Y(n5074) );
  NOR4X1 U6428 ( .A(n5067), .B(n5066), .C(n5065), .D(n5064), .Y(n5068) );
  AO22X1 U6429 ( .A0(n3140), .A1(n279), .B0(n180), .B1(n1174), .Y(n5067) );
  AO22X1 U6430 ( .A0(n3146), .A1(n280), .B0(n184), .B1(n1175), .Y(n5066) );
  AO22X1 U6431 ( .A0(n3152), .A1(n281), .B0(n182), .B1(n1176), .Y(n5065) );
  NOR4X1 U6432 ( .A(n6158), .B(n6157), .C(n6156), .D(n6155), .Y(n6159) );
  AO22X1 U6433 ( .A0(n3141), .A1(n196), .B0(n3138), .B1(n1093), .Y(n6158) );
  AO22X1 U6434 ( .A0(n3147), .A1(n210), .B0(n3144), .B1(n1094), .Y(n6157) );
  AO22X1 U6435 ( .A0(n3153), .A1(n211), .B0(n3150), .B1(n1095), .Y(n6156) );
  NOR4X1 U6436 ( .A(n6149), .B(n6148), .C(n6147), .D(n6146), .Y(n6150) );
  AO22X1 U6437 ( .A0(n3141), .A1(n1107), .B0(n3138), .B1(n222), .Y(n6149) );
  AO22X1 U6438 ( .A0(n3147), .A1(n212), .B0(n3144), .B1(n1096), .Y(n6148) );
  AO22X1 U6439 ( .A0(n3153), .A1(n213), .B0(n3150), .B1(n1097), .Y(n6147) );
  NOR4X1 U6440 ( .A(n6227), .B(n6226), .C(n6225), .D(n6224), .Y(n6228) );
  AO22X1 U6441 ( .A0(n3141), .A1(n57), .B0(n3138), .B1(n1119), .Y(n6227) );
  AO22X1 U6442 ( .A0(n3147), .A1(n234), .B0(n3144), .B1(n1120), .Y(n6226) );
  AO22X1 U6443 ( .A0(n3153), .A1(n235), .B0(n3150), .B1(n1121), .Y(n6225) );
  NOR4X1 U6444 ( .A(n6218), .B(n6217), .C(n6216), .D(n6215), .Y(n6219) );
  AO22X1 U6445 ( .A0(n3142), .A1(n236), .B0(n3138), .B1(n1122), .Y(n6218) );
  AO22X1 U6446 ( .A0(n3148), .A1(n237), .B0(n3144), .B1(n1123), .Y(n6217) );
  AO22X1 U6447 ( .A0(n3154), .A1(n238), .B0(n3150), .B1(n1124), .Y(n6216) );
  NOR4X1 U6448 ( .A(n6248), .B(n6247), .C(n6246), .D(n6245), .Y(n6249) );
  AO22X1 U6449 ( .A0(n3194), .A1(n57), .B0(n3190), .B1(n1119), .Y(n6248) );
  AO22X1 U6450 ( .A0(n3200), .A1(n234), .B0(n3196), .B1(n1120), .Y(n6247) );
  AO22X1 U6451 ( .A0(n3204), .A1(n235), .B0(n3203), .B1(n1121), .Y(n6246) );
  NOR4X1 U6452 ( .A(n6239), .B(n6238), .C(n6237), .D(n6236), .Y(n6240) );
  AO22X1 U6453 ( .A0(n3194), .A1(n236), .B0(n3190), .B1(n1122), .Y(n6239) );
  AO22X1 U6454 ( .A0(n3200), .A1(n237), .B0(n3196), .B1(n1123), .Y(n6238) );
  AO22X1 U6455 ( .A0(n3205), .A1(n238), .B0(n3203), .B1(n1124), .Y(n6237) );
  NOR4X1 U6456 ( .A(n6425), .B(n6424), .C(n6423), .D(n6422), .Y(n6426) );
  AO22X1 U6457 ( .A0(n3141), .A1(n58), .B0(n3138), .B1(n1098), .Y(n6425) );
  AO22X1 U6458 ( .A0(n3147), .A1(n214), .B0(n3144), .B1(n1099), .Y(n6424) );
  AO22X1 U6459 ( .A0(n3153), .A1(n215), .B0(n3150), .B1(n1100), .Y(n6423) );
  NOR4X1 U6460 ( .A(n6416), .B(n6415), .C(n6414), .D(n6413), .Y(n6417) );
  AO22X1 U6461 ( .A0(n3142), .A1(n1108), .B0(n3138), .B1(n223), .Y(n6416) );
  AO22X1 U6462 ( .A0(n3148), .A1(n216), .B0(n3144), .B1(n1101), .Y(n6415) );
  AO22X1 U6463 ( .A0(n3154), .A1(n217), .B0(n3150), .B1(n1102), .Y(n6414) );
  NOR4X1 U6464 ( .A(n6380), .B(n6379), .C(n6378), .D(n6377), .Y(n6381) );
  AO22X1 U6465 ( .A0(n3194), .A1(n59), .B0(n3190), .B1(n1125), .Y(n6380) );
  AO22X1 U6466 ( .A0(n3200), .A1(n239), .B0(n3196), .B1(n1126), .Y(n6379) );
  AO22X1 U6467 ( .A0(n190), .A1(n240), .B0(n3203), .B1(n1127), .Y(n6378) );
  NOR4X1 U6468 ( .A(n6371), .B(n6370), .C(n6369), .D(n6368), .Y(n6372) );
  AO22X1 U6469 ( .A0(n3194), .A1(n241), .B0(n3190), .B1(n1128), .Y(n6371) );
  AO22X1 U6470 ( .A0(n3200), .A1(n242), .B0(n3196), .B1(n1129), .Y(n6370) );
  AO22X1 U6471 ( .A0(n190), .A1(n243), .B0(n3203), .B1(n1130), .Y(n6369) );
  NOR4X1 U6472 ( .A(n6359), .B(n6358), .C(n6357), .D(n6356), .Y(n6360) );
  AO22X1 U6473 ( .A0(n3141), .A1(n59), .B0(n3138), .B1(n1125), .Y(n6359) );
  AO22X1 U6474 ( .A0(n3147), .A1(n239), .B0(n3144), .B1(n1126), .Y(n6358) );
  AO22X1 U6475 ( .A0(n3153), .A1(n240), .B0(n3150), .B1(n1127), .Y(n6357) );
  NOR4X1 U6476 ( .A(n6350), .B(n6349), .C(n6348), .D(n6347), .Y(n6351) );
  AO22X1 U6477 ( .A0(n3142), .A1(n241), .B0(n3138), .B1(n1128), .Y(n6350) );
  AO22X1 U6478 ( .A0(n3148), .A1(n242), .B0(n3144), .B1(n1129), .Y(n6349) );
  AO22X1 U6479 ( .A0(n3154), .A1(n243), .B0(n3150), .B1(n1130), .Y(n6348) );
  NOR4X1 U6480 ( .A(n6518), .B(n6517), .C(n6516), .D(n6515), .Y(n6519) );
  AO22X1 U6481 ( .A0(n3193), .A1(n205), .B0(n3191), .B1(n1201), .Y(n6518) );
  AO22X1 U6482 ( .A0(n3199), .A1(n302), .B0(n3197), .B1(n1202), .Y(n6517) );
  AO22X1 U6483 ( .A0(n3206), .A1(n303), .B0(n179), .B1(n1203), .Y(n6516) );
  NOR4X1 U6484 ( .A(n6509), .B(n6508), .C(n6507), .D(n6506), .Y(n6510) );
  AO22X1 U6485 ( .A0(n3193), .A1(n304), .B0(n3191), .B1(n1204), .Y(n6509) );
  AO22X1 U6486 ( .A0(n3199), .A1(n305), .B0(n3197), .B1(n1205), .Y(n6508) );
  AO22X1 U6487 ( .A0(n3206), .A1(n306), .B0(n3202), .B1(n1206), .Y(n6507) );
  NOR4X1 U6488 ( .A(n5371), .B(n5370), .C(n5369), .D(n5368), .Y(n5372) );
  AO22X1 U6489 ( .A0(n3192), .A1(n197), .B0(n3188), .B1(n1131), .Y(n5371) );
  AO22X1 U6490 ( .A0(n3198), .A1(n244), .B0(n192), .B1(n1132), .Y(n5370) );
  AO22X1 U6491 ( .A0(n3205), .A1(n245), .B0(n3201), .B1(n1133), .Y(n5369) );
  NOR4X1 U6492 ( .A(n5362), .B(n5361), .C(n5360), .D(n5359), .Y(n5363) );
  AO22X1 U6493 ( .A0(n3192), .A1(n246), .B0(n3188), .B1(n1134), .Y(n5362) );
  AO22X1 U6494 ( .A0(n3198), .A1(n247), .B0(n192), .B1(n1135), .Y(n5361) );
  AO22X1 U6495 ( .A0(n3205), .A1(n248), .B0(n3201), .B1(n1136), .Y(n5360) );
  NOR4X1 U6496 ( .A(n5289), .B(n5288), .C(n5287), .D(n5286), .Y(n5290) );
  AO22X1 U6497 ( .A0(n3141), .A1(n60), .B0(n3137), .B1(n1137), .Y(n5289) );
  AO22X1 U6498 ( .A0(n3147), .A1(n249), .B0(n3143), .B1(n1138), .Y(n5288) );
  AO22X1 U6499 ( .A0(n3153), .A1(n1109), .B0(n3149), .B1(n224), .Y(n5287) );
  NOR4X1 U6500 ( .A(n5280), .B(n5279), .C(n5278), .D(n5277), .Y(n5281) );
  AO22X1 U6501 ( .A0(n3141), .A1(n250), .B0(n3137), .B1(n1139), .Y(n5280) );
  AO22X1 U6502 ( .A0(n3147), .A1(n251), .B0(n3143), .B1(n1140), .Y(n5279) );
  AO22X1 U6503 ( .A0(n3153), .A1(n1110), .B0(n3149), .B1(n225), .Y(n5278) );
  NOR4X1 U6504 ( .A(n5245), .B(n5244), .C(n5243), .D(n5242), .Y(n5246) );
  AO22X1 U6505 ( .A0(n3192), .A1(n198), .B0(n3188), .B1(n1141), .Y(n5245) );
  AO22X1 U6506 ( .A0(n3198), .A1(n252), .B0(n192), .B1(n1142), .Y(n5244) );
  AO22X1 U6507 ( .A0(n3205), .A1(n253), .B0(n3201), .B1(n1143), .Y(n5243) );
  NOR4X1 U6508 ( .A(n5236), .B(n5235), .C(n5234), .D(n5233), .Y(n5237) );
  AO22X1 U6509 ( .A0(n3192), .A1(n254), .B0(n3188), .B1(n1144), .Y(n5236) );
  AO22X1 U6510 ( .A0(n3198), .A1(n255), .B0(n192), .B1(n1145), .Y(n5235) );
  AO22X1 U6511 ( .A0(n3205), .A1(n256), .B0(n3201), .B1(n1146), .Y(n5234) );
  NOR4X1 U6512 ( .A(n5224), .B(n5223), .C(n5222), .D(n5221), .Y(n5225) );
  AO22X1 U6513 ( .A0(n3141), .A1(n198), .B0(n3137), .B1(n1141), .Y(n5224) );
  AO22X1 U6514 ( .A0(n3147), .A1(n252), .B0(n3143), .B1(n1142), .Y(n5223) );
  AO22X1 U6515 ( .A0(n3153), .A1(n253), .B0(n3149), .B1(n1143), .Y(n5222) );
  NOR4X1 U6516 ( .A(n5215), .B(n5214), .C(n5213), .D(n5212), .Y(n5216) );
  AO22X1 U6517 ( .A0(n3141), .A1(n254), .B0(n3137), .B1(n1144), .Y(n5215) );
  AO22X1 U6518 ( .A0(n3147), .A1(n255), .B0(n3143), .B1(n1145), .Y(n5214) );
  AO22X1 U6519 ( .A0(n3153), .A1(n256), .B0(n3149), .B1(n1146), .Y(n5213) );
  NOR4X1 U6520 ( .A(n5440), .B(n5439), .C(n5438), .D(n5437), .Y(n5441) );
  AO22X1 U6521 ( .A0(n3192), .A1(n207), .B0(n3188), .B1(n1147), .Y(n5440) );
  AO22X1 U6522 ( .A0(n3198), .A1(n257), .B0(n3197), .B1(n1148), .Y(n5439) );
  AO22X1 U6523 ( .A0(n3205), .A1(n258), .B0(n3201), .B1(n1149), .Y(n5438) );
  NOR4X1 U6524 ( .A(n5431), .B(n5430), .C(n5429), .D(n5428), .Y(n5432) );
  AO22X1 U6525 ( .A0(n3192), .A1(n259), .B0(n3188), .B1(n1150), .Y(n5431) );
  AO22X1 U6526 ( .A0(n3198), .A1(n260), .B0(n3195), .B1(n1151), .Y(n5430) );
  AO22X1 U6527 ( .A0(n3205), .A1(n261), .B0(n3201), .B1(n1152), .Y(n5429) );
  NOR4X1 U6528 ( .A(n5419), .B(n5418), .C(n5417), .D(n5416), .Y(n5420) );
  AO22X1 U6529 ( .A0(n3141), .A1(n207), .B0(n3137), .B1(n1147), .Y(n5419) );
  AO22X1 U6530 ( .A0(n3147), .A1(n257), .B0(n3143), .B1(n1148), .Y(n5418) );
  AO22X1 U6531 ( .A0(n3153), .A1(n258), .B0(n3149), .B1(n1149), .Y(n5417) );
  NOR4X1 U6532 ( .A(n5410), .B(n5409), .C(n5408), .D(n5407), .Y(n5411) );
  AO22X1 U6533 ( .A0(n3141), .A1(n259), .B0(n3137), .B1(n1150), .Y(n5410) );
  AO22X1 U6534 ( .A0(n3147), .A1(n260), .B0(n3143), .B1(n1151), .Y(n5409) );
  AO22X1 U6535 ( .A0(n3153), .A1(n261), .B0(n3149), .B1(n1152), .Y(n5408) );
  NOR4X1 U6536 ( .A(n5027), .B(n5026), .C(n5025), .D(n5024), .Y(n5028) );
  AO22X1 U6537 ( .A0(n188), .A1(n61), .B0(n3190), .B1(n1153), .Y(n5027) );
  AO22X1 U6538 ( .A0(n189), .A1(n262), .B0(n3195), .B1(n1154), .Y(n5026) );
  AO22X1 U6539 ( .A0(n3204), .A1(n263), .B0(n3203), .B1(n1155), .Y(n5025) );
  NOR4X1 U6540 ( .A(n5018), .B(n5017), .C(n5016), .D(n5015), .Y(n5019) );
  AO22X1 U6541 ( .A0(n188), .A1(n264), .B0(n3190), .B1(n1156), .Y(n5018) );
  AO22X1 U6542 ( .A0(n189), .A1(n265), .B0(n3197), .B1(n1157), .Y(n5017) );
  AO22X1 U6543 ( .A0(n3204), .A1(n266), .B0(n3203), .B1(n1158), .Y(n5016) );
  NOR4X1 U6544 ( .A(n5006), .B(n5005), .C(n5004), .D(n5003), .Y(n5007) );
  AO22X1 U6545 ( .A0(n3140), .A1(n61), .B0(n180), .B1(n1153), .Y(n5006) );
  AO22X1 U6546 ( .A0(n3146), .A1(n262), .B0(n184), .B1(n1154), .Y(n5005) );
  AO22X1 U6547 ( .A0(n3152), .A1(n263), .B0(n182), .B1(n1155), .Y(n5004) );
  NOR4X1 U6548 ( .A(n4997), .B(n4996), .C(n4995), .D(n4994), .Y(n4998) );
  AO22X1 U6549 ( .A0(n3140), .A1(n264), .B0(n180), .B1(n1156), .Y(n4997) );
  AO22X1 U6550 ( .A0(n3146), .A1(n265), .B0(n184), .B1(n1157), .Y(n4996) );
  AO22X1 U6551 ( .A0(n3152), .A1(n266), .B0(n182), .B1(n1158), .Y(n4995) );
  NOR4X1 U6552 ( .A(n4957), .B(n4956), .C(n4955), .D(n4954), .Y(n4958) );
  AO22X1 U6553 ( .A0(n188), .A1(n199), .B0(n3190), .B1(n1159), .Y(n4957) );
  AO22X1 U6554 ( .A0(n189), .A1(n267), .B0(n3196), .B1(n1160), .Y(n4956) );
  AO22X1 U6555 ( .A0(n3204), .A1(n268), .B0(n3202), .B1(n1161), .Y(n4955) );
  NOR4X1 U6556 ( .A(n4948), .B(n4947), .C(n4946), .D(n4945), .Y(n4949) );
  AO22X1 U6557 ( .A0(n188), .A1(n269), .B0(n3190), .B1(n1162), .Y(n4948) );
  AO22X1 U6558 ( .A0(n189), .A1(n270), .B0(n3197), .B1(n1163), .Y(n4947) );
  AO22X1 U6559 ( .A0(n3204), .A1(n271), .B0(n3201), .B1(n1164), .Y(n4946) );
  NOR4X1 U6560 ( .A(n4936), .B(n4935), .C(n4934), .D(n4933), .Y(n4937) );
  AO22X1 U6561 ( .A0(n3140), .A1(n199), .B0(n180), .B1(n1159), .Y(n4936) );
  AO22X1 U6562 ( .A0(n3146), .A1(n267), .B0(n184), .B1(n1160), .Y(n4935) );
  AO22X1 U6563 ( .A0(n3152), .A1(n268), .B0(n182), .B1(n1161), .Y(n4934) );
  NOR4X1 U6564 ( .A(n4927), .B(n4926), .C(n4925), .D(n4924), .Y(n4928) );
  AO22X1 U6565 ( .A0(n3140), .A1(n269), .B0(n180), .B1(n1162), .Y(n4927) );
  AO22X1 U6566 ( .A0(n3146), .A1(n270), .B0(n184), .B1(n1163), .Y(n4926) );
  AO22X1 U6567 ( .A0(n3152), .A1(n271), .B0(n182), .B1(n1164), .Y(n4925) );
  NOR4X1 U6568 ( .A(n5169), .B(n5168), .C(n5167), .D(n5166), .Y(n5170) );
  AO22X1 U6569 ( .A0(n188), .A1(n206), .B0(n3190), .B1(n1165), .Y(n5169) );
  AO22X1 U6570 ( .A0(n189), .A1(n272), .B0(n3196), .B1(n1166), .Y(n5168) );
  AO22X1 U6571 ( .A0(n3204), .A1(n273), .B0(n3201), .B1(n1167), .Y(n5167) );
  NOR4X1 U6572 ( .A(n5160), .B(n5159), .C(n5158), .D(n5157), .Y(n5161) );
  AO22X1 U6573 ( .A0(n188), .A1(n274), .B0(n3190), .B1(n1168), .Y(n5160) );
  AO22X1 U6574 ( .A0(n189), .A1(n275), .B0(n3196), .B1(n1169), .Y(n5159) );
  AO22X1 U6575 ( .A0(n3204), .A1(n276), .B0(n3201), .B1(n1170), .Y(n5158) );
  NOR4X1 U6576 ( .A(n5148), .B(n5147), .C(n5146), .D(n5145), .Y(n5149) );
  AO22X1 U6577 ( .A0(n3140), .A1(n206), .B0(n3138), .B1(n1165), .Y(n5148) );
  AO22X1 U6578 ( .A0(n3146), .A1(n272), .B0(n3144), .B1(n1166), .Y(n5147) );
  AO22X1 U6579 ( .A0(n3152), .A1(n273), .B0(n3150), .B1(n1167), .Y(n5146) );
  NOR4X1 U6580 ( .A(n5139), .B(n5138), .C(n5137), .D(n5136), .Y(n5140) );
  AO22X1 U6581 ( .A0(n3140), .A1(n274), .B0(n180), .B1(n1168), .Y(n5139) );
  AO22X1 U6582 ( .A0(n3146), .A1(n275), .B0(n184), .B1(n1169), .Y(n5138) );
  AO22X1 U6583 ( .A0(n3152), .A1(n276), .B0(n182), .B1(n1170), .Y(n5137) );
  AO22X1 U6584 ( .A0(n188), .A1(n70), .B0(n3190), .B1(n1171), .Y(n5097) );
  AO22X1 U6585 ( .A0(n189), .A1(n277), .B0(n3195), .B1(n1172), .Y(n5096) );
  AO22X1 U6586 ( .A0(n3204), .A1(n278), .B0(n179), .B1(n1173), .Y(n5095) );
  NOR4X1 U6587 ( .A(n5088), .B(n5087), .C(n5086), .D(n5085), .Y(n5089) );
  AO22X1 U6588 ( .A0(n188), .A1(n279), .B0(n3190), .B1(n1174), .Y(n5088) );
  AO22X1 U6589 ( .A0(n189), .A1(n280), .B0(n3196), .B1(n1175), .Y(n5087) );
  AO22X1 U6590 ( .A0(n3204), .A1(n281), .B0(n3202), .B1(n1176), .Y(n5086) );
  NOR4X1 U6591 ( .A(n6661), .B(n6660), .C(n6659), .D(n6658), .Y(n6662) );
  AO22X1 U6592 ( .A0(n3192), .A1(n200), .B0(n3191), .B1(n1177), .Y(n6661) );
  AO22X1 U6593 ( .A0(n3198), .A1(n282), .B0(n3197), .B1(n1178), .Y(n6660) );
  AO22X1 U6594 ( .A0(n3206), .A1(n283), .B0(n3202), .B1(n1179), .Y(n6659) );
  NOR4X1 U6595 ( .A(n6652), .B(n6651), .C(n6650), .D(n6649), .Y(n6653) );
  AO22X1 U6596 ( .A0(n3192), .A1(n284), .B0(n3191), .B1(n1180), .Y(n6652) );
  AO22X1 U6597 ( .A0(n3198), .A1(n285), .B0(n3197), .B1(n1181), .Y(n6651) );
  AO22X1 U6598 ( .A0(n3206), .A1(n286), .B0(n179), .B1(n1182), .Y(n6650) );
  NOR4X1 U6599 ( .A(n6640), .B(n6639), .C(n6638), .D(n6637), .Y(n6641) );
  AO22X1 U6600 ( .A0(n3142), .A1(n200), .B0(n3139), .B1(n1177), .Y(n6640) );
  AO22X1 U6601 ( .A0(n3148), .A1(n282), .B0(n3145), .B1(n1178), .Y(n6639) );
  AO22X1 U6602 ( .A0(n3154), .A1(n283), .B0(n3151), .B1(n1179), .Y(n6638) );
  NOR4X1 U6603 ( .A(n6631), .B(n6630), .C(n6629), .D(n6628), .Y(n6632) );
  AO22X1 U6604 ( .A0(n3142), .A1(n284), .B0(n3139), .B1(n1180), .Y(n6631) );
  AO22X1 U6605 ( .A0(n3148), .A1(n285), .B0(n3145), .B1(n1181), .Y(n6630) );
  AO22X1 U6606 ( .A0(n3154), .A1(n286), .B0(n3151), .B1(n1182), .Y(n6629) );
  NOR4X1 U6607 ( .A(n6589), .B(n6588), .C(n6587), .D(n6586), .Y(n6590) );
  AO22X1 U6608 ( .A0(n3194), .A1(n201), .B0(n3191), .B1(n1183), .Y(n6589) );
  AO22X1 U6609 ( .A0(n3200), .A1(n287), .B0(n3197), .B1(n1184), .Y(n6588) );
  AO22X1 U6610 ( .A0(n3206), .A1(n288), .B0(n179), .B1(n1185), .Y(n6587) );
  NOR4X1 U6611 ( .A(n6580), .B(n6579), .C(n6578), .D(n6577), .Y(n6581) );
  AO22X1 U6612 ( .A0(n3192), .A1(n289), .B0(n3191), .B1(n1186), .Y(n6580) );
  AO22X1 U6613 ( .A0(n3198), .A1(n290), .B0(n3197), .B1(n1187), .Y(n6579) );
  AO22X1 U6614 ( .A0(n3206), .A1(n291), .B0(n179), .B1(n1188), .Y(n6578) );
  NOR4X1 U6615 ( .A(n6568), .B(n6567), .C(n6566), .D(n6565), .Y(n6569) );
  AO22X1 U6616 ( .A0(n3142), .A1(n201), .B0(n3139), .B1(n1183), .Y(n6568) );
  AO22X1 U6617 ( .A0(n3148), .A1(n287), .B0(n3145), .B1(n1184), .Y(n6567) );
  AO22X1 U6618 ( .A0(n3154), .A1(n288), .B0(n3151), .B1(n1185), .Y(n6566) );
  NOR4X1 U6619 ( .A(n6559), .B(n6558), .C(n6557), .D(n6556), .Y(n6560) );
  AO22X1 U6620 ( .A0(n3142), .A1(n289), .B0(n3139), .B1(n1186), .Y(n6559) );
  AO22X1 U6621 ( .A0(n3148), .A1(n290), .B0(n3145), .B1(n1187), .Y(n6558) );
  AO22X1 U6622 ( .A0(n3154), .A1(n291), .B0(n3151), .B1(n1188), .Y(n6557) );
  NOR4X1 U6623 ( .A(n6963), .B(n6962), .C(n6961), .D(n6960), .Y(n6964) );
  AO22X1 U6624 ( .A0(n3142), .A1(n63), .B0(n3137), .B1(n1219), .Y(n6963) );
  AO22X1 U6625 ( .A0(n3148), .A1(n317), .B0(n3143), .B1(n1220), .Y(n6962) );
  AO22X1 U6626 ( .A0(n3154), .A1(n318), .B0(n3149), .B1(n1221), .Y(n6961) );
  NOR4X1 U6627 ( .A(n6954), .B(n6953), .C(n6952), .D(n6951), .Y(n6955) );
  AO22X1 U6628 ( .A0(n3142), .A1(n319), .B0(n3137), .B1(n1222), .Y(n6954) );
  AO22X1 U6629 ( .A0(n3148), .A1(n320), .B0(n3143), .B1(n1223), .Y(n6953) );
  AO22X1 U6630 ( .A0(n3154), .A1(n321), .B0(n3149), .B1(n1224), .Y(n6952) );
  NOR4X1 U6631 ( .A(n5795), .B(n5794), .C(n5793), .D(n5792), .Y(n5796) );
  AO22X1 U6632 ( .A0(n3193), .A1(n64), .B0(n3189), .B1(n1279), .Y(n5795) );
  AO22X1 U6633 ( .A0(n3199), .A1(n367), .B0(n3195), .B1(n1280), .Y(n5794) );
  AO22X1 U6634 ( .A0(n190), .A1(n368), .B0(n3202), .B1(n1281), .Y(n5793) );
  NOR4X1 U6635 ( .A(n5786), .B(n5785), .C(n5784), .D(n5783), .Y(n5787) );
  AO22X1 U6636 ( .A0(n3193), .A1(n369), .B0(n3189), .B1(n1282), .Y(n5786) );
  AO22X1 U6637 ( .A0(n3199), .A1(n370), .B0(n3195), .B1(n1283), .Y(n5785) );
  AO22X1 U6638 ( .A0(n3206), .A1(n371), .B0(n3202), .B1(n1284), .Y(n5784) );
  NOR4X1 U6639 ( .A(n5723), .B(n5722), .C(n5721), .D(n5720), .Y(n5724) );
  AO22X1 U6640 ( .A0(n3193), .A1(n65), .B0(n3189), .B1(n1285), .Y(n5723) );
  AO22X1 U6641 ( .A0(n3199), .A1(n372), .B0(n3195), .B1(n1286), .Y(n5722) );
  AO22X1 U6642 ( .A0(n3206), .A1(n373), .B0(n3202), .B1(n1287), .Y(n5721) );
  NOR4X1 U6643 ( .A(n5714), .B(n5713), .C(n5712), .D(n5711), .Y(n5715) );
  AO22X1 U6644 ( .A0(n3193), .A1(n374), .B0(n3189), .B1(n1288), .Y(n5714) );
  AO22X1 U6645 ( .A0(n3199), .A1(n375), .B0(n3195), .B1(n1289), .Y(n5713) );
  AO22X1 U6646 ( .A0(n3206), .A1(n376), .B0(n3202), .B1(n1290), .Y(n5712) );
  NOR4X1 U6647 ( .A(n5525), .B(n5524), .C(n5523), .D(n5522), .Y(n5526) );
  AO22X1 U6648 ( .A0(n3192), .A1(n193), .B0(n3188), .B1(n1189), .Y(n5525) );
  AO22X1 U6649 ( .A0(n3198), .A1(n292), .B0(n3197), .B1(n1190), .Y(n5524) );
  AO22X1 U6650 ( .A0(n3205), .A1(n293), .B0(n3201), .B1(n1191), .Y(n5523) );
  NOR4X1 U6651 ( .A(n5516), .B(n5515), .C(n5514), .D(n5513), .Y(n5517) );
  AO22X1 U6652 ( .A0(n3192), .A1(n294), .B0(n3188), .B1(n1192), .Y(n5516) );
  AO22X1 U6653 ( .A0(n3198), .A1(n295), .B0(n3195), .B1(n1193), .Y(n5515) );
  AO22X1 U6654 ( .A0(n3205), .A1(n296), .B0(n3201), .B1(n1194), .Y(n5514) );
  NOR4X1 U6655 ( .A(n5502), .B(n5501), .C(n5500), .D(n5499), .Y(n5503) );
  AO22X1 U6656 ( .A0(n3141), .A1(n193), .B0(n3137), .B1(n1189), .Y(n5502) );
  AO22X1 U6657 ( .A0(n3147), .A1(n292), .B0(n3143), .B1(n1190), .Y(n5501) );
  AO22X1 U6658 ( .A0(n3153), .A1(n293), .B0(n3149), .B1(n1191), .Y(n5500) );
  NOR4X1 U6659 ( .A(n5493), .B(n5492), .C(n5491), .D(n5490), .Y(n5494) );
  AO22X1 U6660 ( .A0(n3141), .A1(n294), .B0(n3137), .B1(n1192), .Y(n5493) );
  AO22X1 U6661 ( .A0(n3147), .A1(n295), .B0(n3143), .B1(n1193), .Y(n5492) );
  AO22X1 U6662 ( .A0(n3153), .A1(n296), .B0(n3149), .B1(n1194), .Y(n5491) );
  NOR4X1 U6663 ( .A(n5590), .B(n5589), .C(n5588), .D(n5587), .Y(n5591) );
  AO22X1 U6664 ( .A0(n3192), .A1(n62), .B0(n3188), .B1(n1195), .Y(n5590) );
  AO22X1 U6665 ( .A0(n3198), .A1(n297), .B0(n192), .B1(n1196), .Y(n5589) );
  AO22X1 U6666 ( .A0(n3205), .A1(n298), .B0(n3201), .B1(n1197), .Y(n5588) );
  NOR4X1 U6667 ( .A(n5581), .B(n5580), .C(n5579), .D(n5578), .Y(n5582) );
  AO22X1 U6668 ( .A0(n3192), .A1(n299), .B0(n3188), .B1(n1198), .Y(n5581) );
  AO22X1 U6669 ( .A0(n3198), .A1(n300), .B0(n3196), .B1(n1199), .Y(n5580) );
  AO22X1 U6670 ( .A0(n3205), .A1(n301), .B0(n3201), .B1(n1200), .Y(n5579) );
  NOR4X1 U6671 ( .A(n5569), .B(n5568), .C(n5567), .D(n5566), .Y(n5570) );
  AO22X1 U6672 ( .A0(n3141), .A1(n62), .B0(n3137), .B1(n1195), .Y(n5569) );
  AO22X1 U6673 ( .A0(n3147), .A1(n297), .B0(n3143), .B1(n1196), .Y(n5568) );
  AO22X1 U6674 ( .A0(n3153), .A1(n298), .B0(n3149), .B1(n1197), .Y(n5567) );
  NOR4X1 U6675 ( .A(n5560), .B(n5559), .C(n5558), .D(n5557), .Y(n5561) );
  AO22X1 U6676 ( .A0(n3141), .A1(n299), .B0(n3137), .B1(n1198), .Y(n5560) );
  AO22X1 U6677 ( .A0(n3147), .A1(n300), .B0(n3143), .B1(n1199), .Y(n5559) );
  AO22X1 U6678 ( .A0(n3153), .A1(n301), .B0(n3149), .B1(n1200), .Y(n5558) );
  NOR4X1 U6679 ( .A(n6495), .B(n6494), .C(n6493), .D(n6492), .Y(n6496) );
  AO22X1 U6680 ( .A0(n3142), .A1(n205), .B0(n3139), .B1(n1201), .Y(n6495) );
  AO22X1 U6681 ( .A0(n3148), .A1(n302), .B0(n3145), .B1(n1202), .Y(n6494) );
  AO22X1 U6682 ( .A0(n3154), .A1(n303), .B0(n3151), .B1(n1203), .Y(n6493) );
  NOR4X1 U6683 ( .A(n6486), .B(n6485), .C(n6484), .D(n6483), .Y(n6487) );
  AO22X1 U6684 ( .A0(n3142), .A1(n304), .B0(n3139), .B1(n1204), .Y(n6486) );
  AO22X1 U6685 ( .A0(n3148), .A1(n305), .B0(n3145), .B1(n1205), .Y(n6485) );
  AO22X1 U6686 ( .A0(n3154), .A1(n306), .B0(n3151), .B1(n1206), .Y(n6484) );
  NOR4X1 U6687 ( .A(n6718), .B(n6717), .C(n6716), .D(n6715), .Y(n6719) );
  AO22X1 U6688 ( .A0(n3193), .A1(n202), .B0(n3191), .B1(n1261), .Y(n6718) );
  AO22X1 U6689 ( .A0(n3199), .A1(n352), .B0(n3197), .B1(n1262), .Y(n6717) );
  AO22X1 U6690 ( .A0(n3206), .A1(n353), .B0(n3202), .B1(n1263), .Y(n6716) );
  NOR4X1 U6691 ( .A(n6709), .B(n6708), .C(n6707), .D(n6706), .Y(n6710) );
  AO22X1 U6692 ( .A0(n3194), .A1(n354), .B0(n3191), .B1(n1264), .Y(n6709) );
  AO22X1 U6693 ( .A0(n3200), .A1(n355), .B0(n3197), .B1(n1265), .Y(n6708) );
  AO22X1 U6694 ( .A0(n3206), .A1(n356), .B0(n3201), .B1(n1266), .Y(n6707) );
  NOR4X1 U6695 ( .A(n6037), .B(n6036), .C(n6035), .D(n6034), .Y(n6038) );
  AO22X1 U6696 ( .A0(n3193), .A1(n208), .B0(n3189), .B1(n1207), .Y(n6037) );
  AO22X1 U6697 ( .A0(n3199), .A1(n307), .B0(n3195), .B1(n1208), .Y(n6036) );
  AO22X1 U6698 ( .A0(n190), .A1(n308), .B0(n3202), .B1(n1209), .Y(n6035) );
  NOR4X1 U6699 ( .A(n6028), .B(n6027), .C(n6026), .D(n6025), .Y(n6029) );
  AO22X1 U6700 ( .A0(n3193), .A1(n309), .B0(n3189), .B1(n1210), .Y(n6028) );
  AO22X1 U6701 ( .A0(n3199), .A1(n310), .B0(n3195), .B1(n1211), .Y(n6027) );
  AO22X1 U6702 ( .A0(n3206), .A1(n311), .B0(n3202), .B1(n1212), .Y(n6026) );
  NOR4X1 U6703 ( .A(n6014), .B(n6013), .C(n6012), .D(n6011), .Y(n6015) );
  AO22X1 U6704 ( .A0(n3140), .A1(n208), .B0(n3139), .B1(n1207), .Y(n6014) );
  AO22X1 U6705 ( .A0(n3146), .A1(n307), .B0(n3145), .B1(n1208), .Y(n6013) );
  AO22X1 U6706 ( .A0(n3152), .A1(n308), .B0(n3151), .B1(n1209), .Y(n6012) );
  NOR4X1 U6707 ( .A(n6005), .B(n6004), .C(n6003), .D(n6002), .Y(n6006) );
  AO22X1 U6708 ( .A0(n3140), .A1(n309), .B0(n3139), .B1(n1210), .Y(n6005) );
  AO22X1 U6709 ( .A0(n3146), .A1(n310), .B0(n3145), .B1(n1211), .Y(n6004) );
  AO22X1 U6710 ( .A0(n3152), .A1(n311), .B0(n3151), .B1(n1212), .Y(n6003) );
  NOR4X1 U6711 ( .A(n6112), .B(n6111), .C(n6110), .D(n6109), .Y(n6113) );
  AO22X1 U6712 ( .A0(n3194), .A1(n71), .B0(n3190), .B1(n1213), .Y(n6112) );
  AO22X1 U6713 ( .A0(n3200), .A1(n312), .B0(n3196), .B1(n1214), .Y(n6111) );
  AO22X1 U6714 ( .A0(n190), .A1(n313), .B0(n3203), .B1(n1215), .Y(n6110) );
  NOR4X1 U6715 ( .A(n6103), .B(n6102), .C(n6101), .D(n6100), .Y(n6104) );
  AO22X1 U6716 ( .A0(n3194), .A1(n314), .B0(n3190), .B1(n1216), .Y(n6103) );
  AO22X1 U6717 ( .A0(n3200), .A1(n315), .B0(n3196), .B1(n1217), .Y(n6102) );
  AO22X1 U6718 ( .A0(n190), .A1(n316), .B0(n3203), .B1(n1218), .Y(n6101) );
  NOR4X1 U6719 ( .A(n6089), .B(n6088), .C(n6087), .D(n6086), .Y(n6090) );
  AO22X1 U6720 ( .A0(n3141), .A1(n71), .B0(n3138), .B1(n1213), .Y(n6089) );
  AO22X1 U6721 ( .A0(n3147), .A1(n312), .B0(n3144), .B1(n1214), .Y(n6088) );
  AO22X1 U6722 ( .A0(n3153), .A1(n313), .B0(n3150), .B1(n1215), .Y(n6087) );
  NOR4X1 U6723 ( .A(n6080), .B(n6079), .C(n6078), .D(n6077), .Y(n6081) );
  AO22X1 U6724 ( .A0(n3142), .A1(n314), .B0(n3138), .B1(n1216), .Y(n6080) );
  AO22X1 U6725 ( .A0(n3148), .A1(n315), .B0(n3144), .B1(n1217), .Y(n6079) );
  AO22X1 U6726 ( .A0(n3154), .A1(n316), .B0(n3150), .B1(n1218), .Y(n6078) );
  NOR4X1 U6727 ( .A(n6871), .B(n6870), .C(n6869), .D(n6868), .Y(n6872) );
  AO22X1 U6728 ( .A0(n3194), .A1(n203), .B0(n3191), .B1(n1267), .Y(n6871) );
  AO22X1 U6729 ( .A0(n3200), .A1(n357), .B0(n3197), .B1(n1268), .Y(n6870) );
  AO22X1 U6730 ( .A0(n3206), .A1(n358), .B0(n3201), .B1(n1269), .Y(n6869) );
  NOR4X1 U6731 ( .A(n6862), .B(n6861), .C(n6860), .D(n6859), .Y(n6863) );
  AO22X1 U6732 ( .A0(n3192), .A1(n359), .B0(n3191), .B1(n1270), .Y(n6862) );
  AO22X1 U6733 ( .A0(n3198), .A1(n360), .B0(n3197), .B1(n1271), .Y(n6861) );
  AO22X1 U6734 ( .A0(n3206), .A1(n361), .B0(n3203), .B1(n1272), .Y(n6860) );
  NOR4X1 U6735 ( .A(n6942), .B(n6941), .C(n6940), .D(n6939), .Y(n6943) );
  AO22X1 U6736 ( .A0(n3193), .A1(n63), .B0(n3188), .B1(n1219), .Y(n6942) );
  AO22X1 U6737 ( .A0(n3199), .A1(n317), .B0(n3196), .B1(n1220), .Y(n6941) );
  AO22X1 U6738 ( .A0(n3205), .A1(n318), .B0(n179), .B1(n1221), .Y(n6940) );
  NOR4X1 U6739 ( .A(n6933), .B(n6932), .C(n6931), .D(n6930), .Y(n6934) );
  AO22X1 U6740 ( .A0(n3193), .A1(n319), .B0(n3188), .B1(n1222), .Y(n6933) );
  AO22X1 U6741 ( .A0(n3199), .A1(n320), .B0(n3197), .B1(n1223), .Y(n6932) );
  AO22X1 U6742 ( .A0(n3205), .A1(n321), .B0(n179), .B1(n1224), .Y(n6931) );
  NOR4X1 U6743 ( .A(n5663), .B(n5662), .C(n5661), .D(n5660), .Y(n5664) );
  AO22X1 U6744 ( .A0(n3193), .A1(n194), .B0(n3189), .B1(n1225), .Y(n5663) );
  AO22X1 U6745 ( .A0(n3199), .A1(n322), .B0(n3195), .B1(n1226), .Y(n5662) );
  AO22X1 U6746 ( .A0(n3206), .A1(n323), .B0(n3202), .B1(n1227), .Y(n5661) );
  NOR4X1 U6747 ( .A(n5654), .B(n5653), .C(n5652), .D(n5651), .Y(n5655) );
  AO22X1 U6748 ( .A0(n3193), .A1(n324), .B0(n3189), .B1(n1228), .Y(n5654) );
  AO22X1 U6749 ( .A0(n3199), .A1(n325), .B0(n3195), .B1(n1229), .Y(n5653) );
  AO22X1 U6750 ( .A0(n3206), .A1(n326), .B0(n3202), .B1(n1230), .Y(n5652) );
  NOR4X1 U6751 ( .A(n5640), .B(n5639), .C(n5638), .D(n5637), .Y(n5641) );
  AO22X1 U6752 ( .A0(n3140), .A1(n194), .B0(n3139), .B1(n1225), .Y(n5640) );
  AO22X1 U6753 ( .A0(n3146), .A1(n322), .B0(n3145), .B1(n1226), .Y(n5639) );
  AO22X1 U6754 ( .A0(n3152), .A1(n323), .B0(n3151), .B1(n1227), .Y(n5638) );
  NOR4X1 U6755 ( .A(n5631), .B(n5630), .C(n5629), .D(n5628), .Y(n5632) );
  AO22X1 U6756 ( .A0(n3140), .A1(n324), .B0(n3138), .B1(n1228), .Y(n5631) );
  AO22X1 U6757 ( .A0(n3146), .A1(n325), .B0(n3144), .B1(n1229), .Y(n5630) );
  AO22X1 U6758 ( .A0(n3152), .A1(n326), .B0(n3150), .B1(n1230), .Y(n5629) );
  NOR4X1 U6759 ( .A(n6815), .B(n6814), .C(n6813), .D(n6812), .Y(n6816) );
  AO22X1 U6760 ( .A0(n188), .A1(n195), .B0(n3191), .B1(n1231), .Y(n6815) );
  AO22X1 U6761 ( .A0(n189), .A1(n327), .B0(n3197), .B1(n1232), .Y(n6814) );
  AO22X1 U6762 ( .A0(n3206), .A1(n328), .B0(n3203), .B1(n1233), .Y(n6813) );
  NOR4X1 U6763 ( .A(n6806), .B(n6805), .C(n6804), .D(n6803), .Y(n6807) );
  AO22X1 U6764 ( .A0(n188), .A1(n329), .B0(n3191), .B1(n1234), .Y(n6806) );
  AO22X1 U6765 ( .A0(n189), .A1(n330), .B0(n3197), .B1(n1235), .Y(n6805) );
  AO22X1 U6766 ( .A0(n3206), .A1(n331), .B0(n3202), .B1(n1236), .Y(n6804) );
  NOR4X1 U6767 ( .A(n6792), .B(n6791), .C(n6790), .D(n6789), .Y(n6793) );
  AO22X1 U6768 ( .A0(n3142), .A1(n195), .B0(n3139), .B1(n1231), .Y(n6792) );
  AO22X1 U6769 ( .A0(n3148), .A1(n327), .B0(n3145), .B1(n1232), .Y(n6791) );
  AO22X1 U6770 ( .A0(n3154), .A1(n328), .B0(n3151), .B1(n1233), .Y(n6790) );
  NOR4X1 U6771 ( .A(n6783), .B(n6782), .C(n6781), .D(n6780), .Y(n6784) );
  AO22X1 U6772 ( .A0(n3142), .A1(n329), .B0(n3139), .B1(n1234), .Y(n6783) );
  AO22X1 U6773 ( .A0(n3148), .A1(n330), .B0(n3145), .B1(n1235), .Y(n6782) );
  AO22X1 U6774 ( .A0(n3154), .A1(n331), .B0(n3151), .B1(n1236), .Y(n6781) );
  NOR4X1 U6775 ( .A(n5875), .B(n5874), .C(n5873), .D(n5872), .Y(n5876) );
  AO22X1 U6776 ( .A0(n3193), .A1(n69), .B0(n3189), .B1(n1237), .Y(n5875) );
  AO22X1 U6777 ( .A0(n3199), .A1(n332), .B0(n3195), .B1(n1238), .Y(n5874) );
  AO22X1 U6778 ( .A0(n3204), .A1(n333), .B0(n3202), .B1(n1239), .Y(n5873) );
  NOR4X1 U6779 ( .A(n5866), .B(n5865), .C(n5864), .D(n5863), .Y(n5867) );
  AO22X1 U6780 ( .A0(n3193), .A1(n334), .B0(n3189), .B1(n1240), .Y(n5866) );
  AO22X1 U6781 ( .A0(n3199), .A1(n335), .B0(n3195), .B1(n1241), .Y(n5865) );
  AO22X1 U6782 ( .A0(n3205), .A1(n336), .B0(n3202), .B1(n1242), .Y(n5864) );
  NOR4X1 U6783 ( .A(n5852), .B(n5851), .C(n5850), .D(n5849), .Y(n5853) );
  AO22X1 U6784 ( .A0(n3140), .A1(n69), .B0(n3139), .B1(n1237), .Y(n5852) );
  AO22X1 U6785 ( .A0(n3146), .A1(n332), .B0(n3145), .B1(n1238), .Y(n5851) );
  AO22X1 U6786 ( .A0(n3152), .A1(n333), .B0(n3151), .B1(n1239), .Y(n5850) );
  NOR4X1 U6787 ( .A(n5843), .B(n5842), .C(n5841), .D(n5840), .Y(n5844) );
  AO22X1 U6788 ( .A0(n3142), .A1(n334), .B0(n3137), .B1(n1240), .Y(n5843) );
  AO22X1 U6789 ( .A0(n3148), .A1(n335), .B0(n3143), .B1(n1241), .Y(n5842) );
  AO22X1 U6790 ( .A0(n3154), .A1(n336), .B0(n3149), .B1(n1242), .Y(n5841) );
  NOR4X1 U6791 ( .A(n4859), .B(n4858), .C(n4857), .D(n4856), .Y(n4860) );
  AO22X1 U6792 ( .A0(n188), .A1(n204), .B0(n3190), .B1(n1273), .Y(n4859) );
  AO22X1 U6793 ( .A0(n189), .A1(n362), .B0(n192), .B1(n1274), .Y(n4858) );
  AO22X1 U6794 ( .A0(n3204), .A1(n363), .B0(n3202), .B1(n1275), .Y(n4857) );
  NOR4X1 U6795 ( .A(n4850), .B(n4849), .C(n4848), .D(n4847), .Y(n4851) );
  AO22X1 U6796 ( .A0(n3193), .A1(n364), .B0(n3190), .B1(n1276), .Y(n4850) );
  AO22X1 U6797 ( .A0(n3199), .A1(n365), .B0(n192), .B1(n1277), .Y(n4849) );
  AO22X1 U6798 ( .A0(n3204), .A1(n366), .B0(n179), .B1(n1278), .Y(n4848) );
  NOR4X1 U6799 ( .A(n5948), .B(n5947), .C(n5946), .D(n5945), .Y(n5949) );
  AO22X1 U6800 ( .A0(n3193), .A1(n67), .B0(n3189), .B1(n1243), .Y(n5948) );
  AO22X1 U6801 ( .A0(n3199), .A1(n337), .B0(n3195), .B1(n1244), .Y(n5947) );
  AO22X1 U6802 ( .A0(n3206), .A1(n338), .B0(n3202), .B1(n1245), .Y(n5946) );
  NOR4X1 U6803 ( .A(n5939), .B(n5938), .C(n5937), .D(n5936), .Y(n5940) );
  AO22X1 U6804 ( .A0(n3193), .A1(n339), .B0(n3189), .B1(n1246), .Y(n5939) );
  AO22X1 U6805 ( .A0(n3199), .A1(n340), .B0(n3195), .B1(n1247), .Y(n5938) );
  AO22X1 U6806 ( .A0(n3204), .A1(n341), .B0(n3202), .B1(n1248), .Y(n5937) );
  NOR4X1 U6807 ( .A(n5925), .B(n5924), .C(n5923), .D(n5922), .Y(n5926) );
  AO22X1 U6808 ( .A0(n181), .A1(n67), .B0(n3138), .B1(n1243), .Y(n5925) );
  AO22X1 U6809 ( .A0(n185), .A1(n337), .B0(n3144), .B1(n1244), .Y(n5924) );
  AO22X1 U6810 ( .A0(n183), .A1(n338), .B0(n3150), .B1(n1245), .Y(n5923) );
  NOR4X1 U6811 ( .A(n5916), .B(n5915), .C(n5914), .D(n5913), .Y(n5917) );
  AO22X1 U6812 ( .A0(n181), .A1(n339), .B0(n3139), .B1(n1246), .Y(n5916) );
  AO22X1 U6813 ( .A0(n185), .A1(n340), .B0(n3145), .B1(n1247), .Y(n5915) );
  AO22X1 U6814 ( .A0(n183), .A1(n341), .B0(n3151), .B1(n1248), .Y(n5914) );
  NOR4X1 U6815 ( .A(n4795), .B(n4794), .C(n4793), .D(n4792), .Y(n4796) );
  AO22X1 U6816 ( .A0(n3194), .A1(n66), .B0(n3189), .B1(n1249), .Y(n4795) );
  AO22X1 U6817 ( .A0(n3200), .A1(n342), .B0(n192), .B1(n1250), .Y(n4794) );
  AO22X1 U6818 ( .A0(n3204), .A1(n343), .B0(n3202), .B1(n1251), .Y(n4793) );
  NOR4X1 U6819 ( .A(n4786), .B(n4785), .C(n4784), .D(n4783), .Y(n4787) );
  AO22X1 U6820 ( .A0(n3192), .A1(n344), .B0(n3189), .B1(n1252), .Y(n4786) );
  AO22X1 U6821 ( .A0(n3198), .A1(n345), .B0(n192), .B1(n1253), .Y(n4785) );
  AO22X1 U6822 ( .A0(n3204), .A1(n346), .B0(n179), .B1(n1254), .Y(n4784) );
  NOR4X1 U6823 ( .A(n7062), .B(n7061), .C(n7060), .D(n7059), .Y(n7063) );
  AO22X1 U6824 ( .A0(n3193), .A1(n68), .B0(n3188), .B1(n1255), .Y(n7062) );
  AO22X1 U6825 ( .A0(n3199), .A1(n347), .B0(n3195), .B1(n1256), .Y(n7061) );
  AO22X1 U6826 ( .A0(n3205), .A1(n348), .B0(n179), .B1(n1257), .Y(n7060) );
  NOR4X1 U6827 ( .A(n7053), .B(n7052), .C(n7051), .D(n7050), .Y(n7054) );
  AO22X1 U6828 ( .A0(n3193), .A1(n349), .B0(n3188), .B1(n1258), .Y(n7053) );
  AO22X1 U6829 ( .A0(n3199), .A1(n350), .B0(n3196), .B1(n1259), .Y(n7052) );
  AO22X1 U6830 ( .A0(n3205), .A1(n351), .B0(n179), .B1(n1260), .Y(n7051) );
  NOR4X1 U6831 ( .A(n4757), .B(n4756), .C(n4755), .D(n4754), .Y(n4758) );
  AO22X1 U6832 ( .A0(n3140), .A1(n66), .B0(n3137), .B1(n1249), .Y(n4757) );
  AO22X1 U6833 ( .A0(n3146), .A1(n342), .B0(n3143), .B1(n1250), .Y(n4756) );
  AO22X1 U6834 ( .A0(n3152), .A1(n343), .B0(n3149), .B1(n1251), .Y(n4755) );
  NOR4X1 U6835 ( .A(n4748), .B(n4747), .C(n4746), .D(n4745), .Y(n4749) );
  AO22X1 U6836 ( .A0(n3140), .A1(n344), .B0(n3139), .B1(n1252), .Y(n4748) );
  AO22X1 U6837 ( .A0(n3146), .A1(n345), .B0(n3145), .B1(n1253), .Y(n4747) );
  AO22X1 U6838 ( .A0(n3152), .A1(n346), .B0(n3151), .B1(n1254), .Y(n4746) );
  NOR4X1 U6839 ( .A(n7035), .B(n7034), .C(n7033), .D(n7032), .Y(n7036) );
  AO22X1 U6840 ( .A0(n3142), .A1(n68), .B0(n180), .B1(n1255), .Y(n7035) );
  AO22X1 U6841 ( .A0(n3148), .A1(n347), .B0(n184), .B1(n1256), .Y(n7034) );
  AO22X1 U6842 ( .A0(n3154), .A1(n348), .B0(n182), .B1(n1257), .Y(n7033) );
  NOR4X1 U6843 ( .A(n7026), .B(n7025), .C(n7024), .D(n7023), .Y(n7027) );
  AO22X1 U6844 ( .A0(n3142), .A1(n349), .B0(n180), .B1(n1258), .Y(n7026) );
  AO22X1 U6845 ( .A0(n3148), .A1(n350), .B0(n184), .B1(n1259), .Y(n7025) );
  AO22X1 U6846 ( .A0(n3154), .A1(n351), .B0(n182), .B1(n1260), .Y(n7024) );
  NOR4X1 U6847 ( .A(n6739), .B(n6738), .C(n6737), .D(n6736), .Y(n6740) );
  AO22X1 U6848 ( .A0(n3142), .A1(n202), .B0(n3139), .B1(n1261), .Y(n6739) );
  AO22X1 U6849 ( .A0(n3148), .A1(n352), .B0(n3145), .B1(n1262), .Y(n6738) );
  AO22X1 U6850 ( .A0(n3154), .A1(n353), .B0(n3151), .B1(n1263), .Y(n6737) );
  NOR4X1 U6851 ( .A(n6730), .B(n6729), .C(n6728), .D(n6727), .Y(n6731) );
  AO22X1 U6852 ( .A0(n3142), .A1(n354), .B0(n3139), .B1(n1264), .Y(n6730) );
  AO22X1 U6853 ( .A0(n3148), .A1(n355), .B0(n3145), .B1(n1265), .Y(n6729) );
  AO22X1 U6854 ( .A0(n3154), .A1(n356), .B0(n3151), .B1(n1266), .Y(n6728) );
  NOR4X1 U6855 ( .A(n6894), .B(n6893), .C(n6892), .D(n6891), .Y(n6895) );
  AO22X1 U6856 ( .A0(n3142), .A1(n203), .B0(n3139), .B1(n1267), .Y(n6894) );
  AO22X1 U6857 ( .A0(n3148), .A1(n357), .B0(n3145), .B1(n1268), .Y(n6893) );
  AO22X1 U6858 ( .A0(n3154), .A1(n358), .B0(n3151), .B1(n1269), .Y(n6892) );
  NOR4X1 U6859 ( .A(n6885), .B(n6884), .C(n6883), .D(n6882), .Y(n6886) );
  AO22X1 U6860 ( .A0(n3142), .A1(n359), .B0(n3139), .B1(n1270), .Y(n6885) );
  AO22X1 U6861 ( .A0(n3148), .A1(n360), .B0(n3145), .B1(n1271), .Y(n6884) );
  AO22X1 U6862 ( .A0(n3154), .A1(n361), .B0(n3151), .B1(n1272), .Y(n6883) );
  NOR4X1 U6863 ( .A(n4882), .B(n4881), .C(n4880), .D(n4879), .Y(n4883) );
  AO22X1 U6864 ( .A0(n3140), .A1(n204), .B0(n180), .B1(n1273), .Y(n4882) );
  AO22X1 U6865 ( .A0(n3146), .A1(n362), .B0(n184), .B1(n1274), .Y(n4881) );
  AO22X1 U6866 ( .A0(n3152), .A1(n363), .B0(n182), .B1(n1275), .Y(n4880) );
  NOR4X1 U6867 ( .A(n4873), .B(n4872), .C(n4871), .D(n4870), .Y(n4874) );
  AO22X1 U6868 ( .A0(n3140), .A1(n364), .B0(n180), .B1(n1276), .Y(n4873) );
  AO22X1 U6869 ( .A0(n3146), .A1(n365), .B0(n184), .B1(n1277), .Y(n4872) );
  AO22X1 U6870 ( .A0(n3152), .A1(n366), .B0(n182), .B1(n1278), .Y(n4871) );
  NOR4X1 U6871 ( .A(n5774), .B(n5773), .C(n5772), .D(n5771), .Y(n5775) );
  AO22X1 U6872 ( .A0(n3140), .A1(n64), .B0(n3139), .B1(n1279), .Y(n5774) );
  AO22X1 U6873 ( .A0(n3146), .A1(n367), .B0(n3145), .B1(n1280), .Y(n5773) );
  AO22X1 U6874 ( .A0(n3152), .A1(n368), .B0(n3151), .B1(n1281), .Y(n5772) );
  NOR4X1 U6875 ( .A(n5765), .B(n5764), .C(n5763), .D(n5762), .Y(n5766) );
  AO22X1 U6876 ( .A0(n3140), .A1(n369), .B0(n3138), .B1(n1282), .Y(n5765) );
  AO22X1 U6877 ( .A0(n3146), .A1(n370), .B0(n3144), .B1(n1283), .Y(n5764) );
  AO22X1 U6878 ( .A0(n3152), .A1(n371), .B0(n3150), .B1(n1284), .Y(n5763) );
  NOR4X1 U6879 ( .A(n5702), .B(n5701), .C(n5700), .D(n5699), .Y(n5703) );
  AO22X1 U6880 ( .A0(n3140), .A1(n65), .B0(n3139), .B1(n1285), .Y(n5702) );
  AO22X1 U6881 ( .A0(n3146), .A1(n372), .B0(n3145), .B1(n1286), .Y(n5701) );
  AO22X1 U6882 ( .A0(n3152), .A1(n373), .B0(n3151), .B1(n1287), .Y(n5700) );
  NOR4X1 U6883 ( .A(n5693), .B(n5692), .C(n5691), .D(n5690), .Y(n5694) );
  AO22X1 U6884 ( .A0(n3140), .A1(n374), .B0(n3138), .B1(n1288), .Y(n5693) );
  AO22X1 U6885 ( .A0(n3146), .A1(n375), .B0(n3144), .B1(n1289), .Y(n5692) );
  AO22X1 U6886 ( .A0(n3152), .A1(n376), .B0(n3150), .B1(n1290), .Y(n5691) );
  NAND2X2 U6887 ( .A(n3010), .B(\D_cache/n315 ), .Y(\D_cache/n250 ) );
  NAND2X2 U6888 ( .A(n3010), .B(\D_cache/n451 ), .Y(\D_cache/n387 ) );
  NAND2X1 U6889 ( .A(n4635), .B(\i_MIPS/n347 ), .Y(n5990) );
  CLKINVX1 U6890 ( .A(n8340), .Y(n8336) );
  NAND2X2 U6891 ( .A(n3076), .B(n4017), .Y(n6334) );
  AND2X2 U6892 ( .A(\i_MIPS/n318 ), .B(\i_MIPS/n316 ), .Y(n2870) );
  AND2X2 U6893 ( .A(\i_MIPS/n230 ), .B(\i_MIPS/n231 ), .Y(n2871) );
  AND2X2 U6894 ( .A(\i_MIPS/n314 ), .B(\i_MIPS/n312 ), .Y(n2872) );
  AND2X2 U6895 ( .A(\i_MIPS/n228 ), .B(\i_MIPS/n229 ), .Y(n2873) );
  NAND3BX1 U6896 ( .AN(n2987), .B(n5457), .C(n5120), .Y(n5396) );
  OA22X1 U6897 ( .A0(\i_MIPS/n355 ), .A1(n3092), .B0(\i_MIPS/n356 ), .B1(n3087), .Y(n5120) );
  NAND3BX1 U6898 ( .AN(n2905), .B(n5744), .C(n5743), .Y(n6673) );
  OA22X1 U6899 ( .A0(\i_MIPS/n356 ), .A1(n3092), .B0(\i_MIPS/n355 ), .B1(n3087), .Y(n5743) );
  CLKINVX1 U6900 ( .A(n8372), .Y(n8368) );
  CLKINVX1 U6901 ( .A(n8387), .Y(n8383) );
  CLKINVX1 U6902 ( .A(n8358), .Y(n8354) );
  CLKINVX1 U6903 ( .A(\D_cache/N63 ), .Y(n8752) );
  CLKINVX1 U6904 ( .A(\D_cache/N69 ), .Y(n8758) );
  CLKINVX1 U6905 ( .A(\D_cache/N57 ), .Y(n8746) );
  CLKINVX1 U6906 ( .A(\D_cache/N60 ), .Y(n8749) );
  CLKINVX1 U6907 ( .A(\D_cache/N95 ), .Y(n8765) );
  CLKINVX1 U6908 ( .A(\D_cache/N101 ), .Y(n8771) );
  CLKINVX1 U6909 ( .A(\D_cache/N89 ), .Y(n8759) );
  CLKINVX1 U6910 ( .A(\D_cache/N92 ), .Y(n8762) );
  CLKINVX1 U6911 ( .A(\D_cache/N166 ), .Y(n8884) );
  NAND2BX1 U6912 ( .AN(n3000), .B(n8645), .Y(n7211) );
  NAND2BX1 U6913 ( .AN(n3001), .B(n8613), .Y(n7209) );
  CLKINVX1 U6914 ( .A(\D_cache/N67 ), .Y(n8756) );
  CLKINVX1 U6915 ( .A(\D_cache/N64 ), .Y(n8753) );
  CLKINVX1 U6916 ( .A(\D_cache/N62 ), .Y(n8751) );
  CLKINVX1 U6917 ( .A(\D_cache/N65 ), .Y(n8754) );
  CLKINVX1 U6918 ( .A(\D_cache/N61 ), .Y(n8750) );
  CLKINVX1 U6919 ( .A(\D_cache/N59 ), .Y(n8748) );
  CLKINVX1 U6920 ( .A(\D_cache/N58 ), .Y(n8747) );
  CLKINVX1 U6921 ( .A(\D_cache/N68 ), .Y(n8757) );
  CLKINVX1 U6922 ( .A(\D_cache/N99 ), .Y(n8769) );
  CLKINVX1 U6923 ( .A(\D_cache/N96 ), .Y(n8766) );
  CLKINVX1 U6924 ( .A(\D_cache/N94 ), .Y(n8764) );
  CLKINVX1 U6925 ( .A(\D_cache/N93 ), .Y(n8763) );
  CLKINVX1 U6926 ( .A(\D_cache/N91 ), .Y(n8761) );
  CLKINVX1 U6927 ( .A(\D_cache/N90 ), .Y(n8760) );
  CLKINVX1 U6928 ( .A(\D_cache/N100 ), .Y(n8770) );
  NAND2BX1 U6929 ( .AN(n3000), .B(n8646), .Y(n7235) );
  NAND2BX1 U6930 ( .AN(n3001), .B(n8614), .Y(n7233) );
  NAND2X1 U6931 ( .A(n5828), .B(n5821), .Y(n5832) );
  CLKINVX1 U6932 ( .A(\i_MIPS/Control_ID/n12 ), .Y(n7307) );
  CLKINVX1 U6933 ( .A(n7842), .Y(n8278) );
  NAND2X1 U6934 ( .A(n5382), .B(n5970), .Y(n6461) );
  CLKMX2X2 U6935 ( .A(n5972), .B(n2986), .S0(n4016), .Y(n5898) );
  NAND2BX1 U6936 ( .AN(n3000), .B(n8644), .Y(n7187) );
  NAND2BX1 U6937 ( .AN(n3001), .B(n8612), .Y(n7185) );
  NAND4X1 U6938 ( .A(n7260), .B(n7259), .C(n7258), .D(n7257), .Y(n7795) );
  NAND2BX1 U6939 ( .AN(n3000), .B(n8647), .Y(n7259) );
  NAND2BX1 U6940 ( .AN(n3001), .B(n8615), .Y(n7257) );
  NAND2BX1 U6941 ( .AN(n3576), .B(n8583), .Y(n7258) );
  NAND4X1 U6942 ( .A(n7304), .B(n7303), .C(n7302), .D(n7301), .Y(n7794) );
  NAND2BX1 U6943 ( .AN(n3000), .B(n8649), .Y(n7303) );
  NAND2BX1 U6944 ( .AN(n3001), .B(n8617), .Y(n7301) );
  NAND2BX1 U6945 ( .AN(n3576), .B(n8585), .Y(n7302) );
  NAND4X1 U6946 ( .A(n7284), .B(n7283), .C(n7282), .D(n7281), .Y(n7796) );
  NAND2BX1 U6947 ( .AN(n3000), .B(n8648), .Y(n7283) );
  NAND2BX1 U6948 ( .AN(n3001), .B(n8616), .Y(n7281) );
  NAND2BX1 U6949 ( .AN(n3576), .B(n8584), .Y(n7282) );
  CLKINVX1 U6950 ( .A(n6474), .Y(n6689) );
  CLKINVX1 U6951 ( .A(n5681), .Y(n5733) );
  CLKINVX1 U6952 ( .A(n5738), .Y(n5755) );
  CLKINVX1 U6953 ( .A(n6914), .Y(n6917) );
  CLKINVX1 U6954 ( .A(\D_cache/N31 ), .Y(n8809) );
  CLKINVX1 U6955 ( .A(n5958), .Y(n5959) );
  CLKINVX1 U6956 ( .A(n6613), .Y(n4919) );
  CLKINVX1 U6957 ( .A(n6763), .Y(n6771) );
  CLKINVX1 U6958 ( .A(\D_cache/N77 ), .Y(n8840) );
  CLKINVX1 U6959 ( .A(\D_cache/N80 ), .Y(n8843) );
  CLKINVX1 U6960 ( .A(\D_cache/N79 ), .Y(n8842) );
  CLKINVX1 U6961 ( .A(\D_cache/N75 ), .Y(n8838) );
  CLKINVX1 U6962 ( .A(\D_cache/N78 ), .Y(n8841) );
  CLKINVX1 U6963 ( .A(\D_cache/N74 ), .Y(n8837) );
  CLKINVX1 U6964 ( .A(\D_cache/N85 ), .Y(n8848) );
  CLKINVX1 U6965 ( .A(\D_cache/N72 ), .Y(n8835) );
  CLKINVX1 U6966 ( .A(\D_cache/N71 ), .Y(n8834) );
  CLKINVX1 U6967 ( .A(\D_cache/N70 ), .Y(n8833) );
  CLKINVX1 U6968 ( .A(\D_cache/N76 ), .Y(n8839) );
  CLKINVX1 U6969 ( .A(\D_cache/N81 ), .Y(n8844) );
  CLKINVX1 U6970 ( .A(\D_cache/N86 ), .Y(n8849) );
  CLKINVX1 U6971 ( .A(\D_cache/N109 ), .Y(n8859) );
  CLKINVX1 U6972 ( .A(\D_cache/N117 ), .Y(n8867) );
  CLKINVX1 U6973 ( .A(\D_cache/N113 ), .Y(n8863) );
  CLKINVX1 U6974 ( .A(\D_cache/N118 ), .Y(n8868) );
  CLKINVX1 U6975 ( .A(\D_cache/N107 ), .Y(n8857) );
  CLKINVX1 U6976 ( .A(\D_cache/N102 ), .Y(n8852) );
  CLKINVX1 U6977 ( .A(\D_cache/N108 ), .Y(n8858) );
  CLKINVX1 U6978 ( .A(\D_cache/N172 ), .Y(n8890) );
  CLKINVX1 U6979 ( .A(\D_cache/N169 ), .Y(n8887) );
  CLKINVX1 U6980 ( .A(\D_cache/N154 ), .Y(n8872) );
  CLKINVX1 U6981 ( .A(\D_cache/N162 ), .Y(n8880) );
  CLKINVX1 U6982 ( .A(\D_cache/N156 ), .Y(n8874) );
  CLKINVX1 U6983 ( .A(\D_cache/N182 ), .Y(n8900) );
  CLKINVX1 U6984 ( .A(\D_cache/N155 ), .Y(n8873) );
  CLKINVX1 U6985 ( .A(\D_cache/N153 ), .Y(n8871) );
  CLKINVX1 U6986 ( .A(\D_cache/N105 ), .Y(n8855) );
  CLKINVX1 U6987 ( .A(\D_cache/N73 ), .Y(n8836) );
  CLKMX2X2 U6988 ( .A(n6757), .B(n5620), .S0(n4016), .Y(n6825) );
  CLKINVX1 U6989 ( .A(n6693), .Y(n6684) );
  OAI222XL U6990 ( .A0(n3585), .A1(n205), .B0(n3685), .B1(n3582), .C0(n3689), 
        .C1(\i_MIPS/n201 ), .Y(n8783) );
  MXI2X1 U6991 ( .A(n5397), .B(n5121), .S0(n4016), .Y(n2881) );
  CLKINVX1 U6992 ( .A(\D_cache/N33 ), .Y(n8810) );
  CLKINVX1 U6993 ( .A(n5042), .Y(n5043) );
  INVX3 U6994 ( .A(n3076), .Y(n5970) );
  AO22X1 U6995 ( .A0(n3211), .A1(n218), .B0(n3207), .B1(n1103), .Y(n6176) );
  AO22X1 U6996 ( .A0(n3211), .A1(n219), .B0(n3207), .B1(n1104), .Y(n6167) );
  AO22X1 U6997 ( .A0(n3211), .A1(n1111), .B0(n3208), .B1(n226), .Y(n5307) );
  AO22X1 U6998 ( .A0(n3211), .A1(n1112), .B0(n3208), .B1(n227), .Y(n5298) );
  AO22X1 U6999 ( .A0(n3213), .A1(n377), .B0(n3207), .B1(n1291), .Y(n6308) );
  AO22X1 U7000 ( .A0(n3211), .A1(n378), .B0(n3207), .B1(n1292), .Y(n6299) );
  AO22X1 U7001 ( .A0(n3160), .A1(n377), .B0(n3157), .B1(n1291), .Y(n6287) );
  AO22X1 U7002 ( .A0(n3160), .A1(n378), .B0(n3157), .B1(n1292), .Y(n6278) );
  AO22X1 U7003 ( .A0(n3211), .A1(n220), .B0(n3207), .B1(n1105), .Y(n6443) );
  AO22X1 U7004 ( .A0(n3213), .A1(n221), .B0(n3207), .B1(n1106), .Y(n6434) );
  AO22X1 U7005 ( .A0(n3160), .A1(n383), .B0(n3155), .B1(n1297), .Y(n5347) );
  AO22X1 U7006 ( .A0(n3160), .A1(n384), .B0(n3155), .B1(n1298), .Y(n5338) );
  AO22X1 U7007 ( .A0(n3159), .A1(n228), .B0(n3155), .B1(n1348), .Y(n5073) );
  AO22X1 U7008 ( .A0(n3159), .A1(n395), .B0(n3155), .B1(n1309), .Y(n5064) );
  AO22X1 U7009 ( .A0(n3160), .A1(n218), .B0(n3157), .B1(n1103), .Y(n6155) );
  AO22X1 U7010 ( .A0(n3160), .A1(n219), .B0(n3157), .B1(n1104), .Y(n6146) );
  AO22X1 U7011 ( .A0(n3160), .A1(n379), .B0(n3157), .B1(n1293), .Y(n6224) );
  AO22X1 U7012 ( .A0(n3161), .A1(n380), .B0(n3157), .B1(n1294), .Y(n6215) );
  AO22X1 U7013 ( .A0(n191), .A1(n379), .B0(n3207), .B1(n1293), .Y(n6245) );
  AO22X1 U7014 ( .A0(n3213), .A1(n380), .B0(n3207), .B1(n1294), .Y(n6236) );
  AO22X1 U7015 ( .A0(n3160), .A1(n220), .B0(n3157), .B1(n1105), .Y(n6422) );
  AO22X1 U7016 ( .A0(n3161), .A1(n221), .B0(n3157), .B1(n1106), .Y(n6413) );
  AO22X1 U7017 ( .A0(n3213), .A1(n381), .B0(n3207), .B1(n1295), .Y(n6377) );
  AO22X1 U7018 ( .A0(n3212), .A1(n382), .B0(n3207), .B1(n1296), .Y(n6368) );
  AO22X1 U7019 ( .A0(n3160), .A1(n381), .B0(n3157), .B1(n1295), .Y(n6356) );
  AO22X1 U7020 ( .A0(n3161), .A1(n382), .B0(n3157), .B1(n1296), .Y(n6347) );
  AO22X1 U7021 ( .A0(n3213), .A1(n404), .B0(n3210), .B1(n1318), .Y(n6515) );
  AO22X1 U7022 ( .A0(n3213), .A1(n405), .B0(n3210), .B1(n1319), .Y(n6506) );
  AO22X1 U7023 ( .A0(n3211), .A1(n383), .B0(n3208), .B1(n1297), .Y(n5368) );
  AO22X1 U7024 ( .A0(n3211), .A1(n384), .B0(n3208), .B1(n1298), .Y(n5359) );
  AO22X1 U7025 ( .A0(n3160), .A1(n1111), .B0(n3155), .B1(n226), .Y(n5286) );
  AO22X1 U7026 ( .A0(n3160), .A1(n1112), .B0(n3155), .B1(n227), .Y(n5277) );
  AO22X1 U7027 ( .A0(n3211), .A1(n385), .B0(n3208), .B1(n1299), .Y(n5242) );
  AO22X1 U7028 ( .A0(n3211), .A1(n386), .B0(n3208), .B1(n1300), .Y(n5233) );
  AO22X1 U7029 ( .A0(n3160), .A1(n385), .B0(n3155), .B1(n1299), .Y(n5221) );
  AO22X1 U7030 ( .A0(n3160), .A1(n386), .B0(n3155), .B1(n1300), .Y(n5212) );
  AO22X1 U7031 ( .A0(n3211), .A1(n387), .B0(n3208), .B1(n1301), .Y(n5437) );
  AO22X1 U7032 ( .A0(n3211), .A1(n388), .B0(n3208), .B1(n1302), .Y(n5428) );
  AO22X1 U7033 ( .A0(n3160), .A1(n387), .B0(n3155), .B1(n1301), .Y(n5416) );
  AO22X1 U7034 ( .A0(n3160), .A1(n388), .B0(n3155), .B1(n1302), .Y(n5407) );
  AO22X1 U7035 ( .A0(n191), .A1(n389), .B0(n3207), .B1(n1303), .Y(n5024) );
  AO22X1 U7036 ( .A0(n191), .A1(n390), .B0(n3207), .B1(n1304), .Y(n5015) );
  AO22X1 U7037 ( .A0(n3159), .A1(n389), .B0(n3155), .B1(n1303), .Y(n5003) );
  AO22X1 U7038 ( .A0(n3159), .A1(n390), .B0(n3155), .B1(n1304), .Y(n4994) );
  AO22X1 U7039 ( .A0(n3213), .A1(n391), .B0(n3207), .B1(n1305), .Y(n4954) );
  AO22X1 U7040 ( .A0(n191), .A1(n392), .B0(n3207), .B1(n1306), .Y(n4945) );
  AO22X1 U7041 ( .A0(n3159), .A1(n391), .B0(n3155), .B1(n1305), .Y(n4933) );
  AO22X1 U7042 ( .A0(n3159), .A1(n392), .B0(n3155), .B1(n1306), .Y(n4924) );
  AO22X1 U7043 ( .A0(n191), .A1(n393), .B0(n3207), .B1(n1307), .Y(n5166) );
  AO22X1 U7044 ( .A0(n191), .A1(n394), .B0(n3207), .B1(n1308), .Y(n5157) );
  AO22X1 U7045 ( .A0(n3159), .A1(n393), .B0(n3155), .B1(n1307), .Y(n5145) );
  AO22X1 U7046 ( .A0(n3159), .A1(n394), .B0(n3155), .B1(n1308), .Y(n5136) );
  AO22X1 U7047 ( .A0(n191), .A1(n395), .B0(n3207), .B1(n1309), .Y(n5085) );
  AO22X1 U7048 ( .A0(n3213), .A1(n396), .B0(n3210), .B1(n1310), .Y(n6658) );
  AO22X1 U7049 ( .A0(n3213), .A1(n397), .B0(n3210), .B1(n1311), .Y(n6649) );
  AO22X1 U7050 ( .A0(n3161), .A1(n396), .B0(n3158), .B1(n1310), .Y(n6637) );
  AO22X1 U7051 ( .A0(n3161), .A1(n397), .B0(n3158), .B1(n1311), .Y(n6628) );
  AO22X1 U7052 ( .A0(n3213), .A1(n398), .B0(n3210), .B1(n1312), .Y(n6586) );
  AO22X1 U7053 ( .A0(n3213), .A1(n399), .B0(n3210), .B1(n1313), .Y(n6577) );
  AO22X1 U7054 ( .A0(n3161), .A1(n398), .B0(n3158), .B1(n1312), .Y(n6565) );
  AO22X1 U7055 ( .A0(n3161), .A1(n399), .B0(n3158), .B1(n1313), .Y(n6556) );
  AO22X1 U7056 ( .A0(n3161), .A1(n410), .B0(n3157), .B1(n1324), .Y(n6960) );
  AO22X1 U7057 ( .A0(n3161), .A1(n411), .B0(n3157), .B1(n1325), .Y(n6951) );
  AO22X1 U7058 ( .A0(n3212), .A1(n430), .B0(n3209), .B1(n1344), .Y(n5792) );
  AO22X1 U7059 ( .A0(n3212), .A1(n431), .B0(n3209), .B1(n1345), .Y(n5783) );
  AO22X1 U7060 ( .A0(n3212), .A1(n432), .B0(n3209), .B1(n1346), .Y(n5720) );
  AO22X1 U7061 ( .A0(n3212), .A1(n433), .B0(n3209), .B1(n1347), .Y(n5711) );
  AO22X1 U7062 ( .A0(n3211), .A1(n400), .B0(n3208), .B1(n1314), .Y(n5522) );
  AO22X1 U7063 ( .A0(n3211), .A1(n401), .B0(n3208), .B1(n1315), .Y(n5513) );
  AO22X1 U7064 ( .A0(n3160), .A1(n400), .B0(n3155), .B1(n1314), .Y(n5499) );
  AO22X1 U7065 ( .A0(n3160), .A1(n401), .B0(n3155), .B1(n1315), .Y(n5490) );
  AO22X1 U7066 ( .A0(n3211), .A1(n402), .B0(n3208), .B1(n1316), .Y(n5587) );
  AO22X1 U7067 ( .A0(n3211), .A1(n403), .B0(n3208), .B1(n1317), .Y(n5578) );
  AO22X1 U7068 ( .A0(n3160), .A1(n402), .B0(n3155), .B1(n1316), .Y(n5566) );
  AO22X1 U7069 ( .A0(n3160), .A1(n403), .B0(n3155), .B1(n1317), .Y(n5557) );
  AO22X1 U7070 ( .A0(n3161), .A1(n404), .B0(n3158), .B1(n1318), .Y(n6492) );
  AO22X1 U7071 ( .A0(n3161), .A1(n405), .B0(n3158), .B1(n1319), .Y(n6483) );
  AO22X1 U7072 ( .A0(n3213), .A1(n424), .B0(n3210), .B1(n1338), .Y(n6715) );
  AO22X1 U7073 ( .A0(n3213), .A1(n425), .B0(n3210), .B1(n1339), .Y(n6706) );
  AO22X1 U7074 ( .A0(n3212), .A1(n406), .B0(n3209), .B1(n1320), .Y(n6034) );
  AO22X1 U7075 ( .A0(n3212), .A1(n407), .B0(n3209), .B1(n1321), .Y(n6025) );
  AO22X1 U7076 ( .A0(n3159), .A1(n406), .B0(n3156), .B1(n1320), .Y(n6011) );
  AO22X1 U7077 ( .A0(n3159), .A1(n407), .B0(n3156), .B1(n1321), .Y(n6002) );
  AO22X1 U7078 ( .A0(n3212), .A1(n408), .B0(n3209), .B1(n1322), .Y(n6109) );
  AO22X1 U7079 ( .A0(n3211), .A1(n409), .B0(n3209), .B1(n1323), .Y(n6100) );
  AO22X1 U7080 ( .A0(n3160), .A1(n408), .B0(n3157), .B1(n1322), .Y(n6086) );
  AO22X1 U7081 ( .A0(n3161), .A1(n409), .B0(n3157), .B1(n1323), .Y(n6077) );
  AO22X1 U7082 ( .A0(n3213), .A1(n426), .B0(n3210), .B1(n1340), .Y(n6868) );
  AO22X1 U7083 ( .A0(n3213), .A1(n427), .B0(n3210), .B1(n1341), .Y(n6859) );
  AO22X1 U7084 ( .A0(n3212), .A1(n410), .B0(n3208), .B1(n1324), .Y(n6939) );
  AO22X1 U7085 ( .A0(n3212), .A1(n411), .B0(n3208), .B1(n1325), .Y(n6930) );
  AO22X1 U7086 ( .A0(n3212), .A1(n412), .B0(n3209), .B1(n1326), .Y(n5660) );
  AO22X1 U7087 ( .A0(n3212), .A1(n413), .B0(n3209), .B1(n1327), .Y(n5651) );
  AO22X1 U7088 ( .A0(n3159), .A1(n412), .B0(n3156), .B1(n1326), .Y(n5637) );
  AO22X1 U7089 ( .A0(n3159), .A1(n413), .B0(n3156), .B1(n1327), .Y(n5628) );
  AO22X1 U7090 ( .A0(n3213), .A1(n414), .B0(n3210), .B1(n1328), .Y(n6812) );
  AO22X1 U7091 ( .A0(n3213), .A1(n415), .B0(n3210), .B1(n1329), .Y(n6803) );
  AO22X1 U7092 ( .A0(n3161), .A1(n414), .B0(n3158), .B1(n1328), .Y(n6789) );
  AO22X1 U7093 ( .A0(n3161), .A1(n415), .B0(n3158), .B1(n1329), .Y(n6780) );
  AO22X1 U7094 ( .A0(n3212), .A1(n416), .B0(n3209), .B1(n1330), .Y(n5872) );
  AO22X1 U7095 ( .A0(n3212), .A1(n417), .B0(n3209), .B1(n1331), .Y(n5863) );
  AO22X1 U7096 ( .A0(n3159), .A1(n416), .B0(n3156), .B1(n1330), .Y(n5849) );
  AO22X1 U7097 ( .A0(n3161), .A1(n417), .B0(n3156), .B1(n1331), .Y(n5840) );
  AO22X1 U7098 ( .A0(n191), .A1(n428), .B0(n3207), .B1(n1342), .Y(n4856) );
  AO22X1 U7099 ( .A0(n191), .A1(n429), .B0(n3207), .B1(n1343), .Y(n4847) );
  AO22X1 U7100 ( .A0(n3212), .A1(n418), .B0(n3209), .B1(n1332), .Y(n5945) );
  AO22X1 U7101 ( .A0(n3212), .A1(n419), .B0(n3209), .B1(n1333), .Y(n5936) );
  AO22X1 U7102 ( .A0(n186), .A1(n418), .B0(n3156), .B1(n1332), .Y(n5922) );
  AO22X1 U7103 ( .A0(n186), .A1(n419), .B0(n3156), .B1(n1333), .Y(n5913) );
  AO22X1 U7104 ( .A0(n191), .A1(n420), .B0(n3207), .B1(n1334), .Y(n4792) );
  AO22X1 U7105 ( .A0(n3211), .A1(n421), .B0(n3207), .B1(n1335), .Y(n4783) );
  AO22X1 U7106 ( .A0(n3212), .A1(n422), .B0(n3208), .B1(n1336), .Y(n7059) );
  AO22X1 U7107 ( .A0(n3212), .A1(n423), .B0(n3208), .B1(n1337), .Y(n7050) );
  AO22X1 U7108 ( .A0(n3159), .A1(n420), .B0(n3156), .B1(n1334), .Y(n4754) );
  AO22X1 U7109 ( .A0(n3159), .A1(n421), .B0(n3156), .B1(n1335), .Y(n4745) );
  AO22X1 U7110 ( .A0(n3161), .A1(n422), .B0(n3157), .B1(n1336), .Y(n7032) );
  AO22X1 U7111 ( .A0(n3161), .A1(n423), .B0(n3157), .B1(n1337), .Y(n7023) );
  AO22X1 U7112 ( .A0(n3161), .A1(n424), .B0(n3158), .B1(n1338), .Y(n6736) );
  AO22X1 U7113 ( .A0(n3161), .A1(n425), .B0(n3158), .B1(n1339), .Y(n6727) );
  AO22X1 U7114 ( .A0(n3161), .A1(n426), .B0(n3158), .B1(n1340), .Y(n6891) );
  AO22X1 U7115 ( .A0(n3161), .A1(n427), .B0(n3158), .B1(n1341), .Y(n6882) );
  AO22X1 U7116 ( .A0(n3159), .A1(n428), .B0(n3155), .B1(n1342), .Y(n4879) );
  AO22X1 U7117 ( .A0(n3159), .A1(n429), .B0(n3155), .B1(n1343), .Y(n4870) );
  AO22X1 U7118 ( .A0(n3159), .A1(n430), .B0(n3156), .B1(n1344), .Y(n5771) );
  AO22X1 U7119 ( .A0(n3159), .A1(n431), .B0(n3156), .B1(n1345), .Y(n5762) );
  AO22X1 U7120 ( .A0(n3159), .A1(n432), .B0(n3156), .B1(n1346), .Y(n5699) );
  AO22X1 U7121 ( .A0(n3159), .A1(n433), .B0(n3156), .B1(n1347), .Y(n5690) );
  CLKINVX1 U7122 ( .A(\i_MIPS/forward_unit/n10 ), .Y(n4764) );
  CLKINVX1 U7123 ( .A(\D_cache/n214 ), .Y(n3974) );
  CLKBUFX3 U7124 ( .A(n1082), .Y(n4017) );
  CLKBUFX3 U7125 ( .A(n8410), .Y(n3586) );
  OA21X2 U7126 ( .A0(n3949), .A1(n8772), .B0(n8808), .Y(\D_cache/n205 ) );
  NOR3X1 U7127 ( .A(n78), .B(n963), .C(n53), .Y(\i_MIPS/Register/n105 ) );
  NAND3BX1 U7128 ( .AN(n7305), .B(n7308), .C(\i_MIPS/n324 ), .Y(
        \i_MIPS/Control_ID/n10 ) );
  NAND4X1 U7129 ( .A(n8102), .B(n8101), .C(n8100), .D(n8099), .Y(n8672) );
  NAND4X1 U7130 ( .A(n8112), .B(n8111), .C(n8110), .D(n8109), .Y(n8576) );
  NAND4X1 U7131 ( .A(n8118), .B(n8117), .C(n8116), .D(n8115), .Y(n8608) );
  NAND4X1 U7132 ( .A(n8107), .B(n8106), .C(n8105), .D(n8104), .Y(n8640) );
  NAND2X1 U7133 ( .A(\i_MIPS/n322 ), .B(\i_MIPS/n332 ), .Y(n7312) );
  NAND4X1 U7134 ( .A(n7510), .B(n7509), .C(n7508), .D(n7507), .Y(n8074) );
  NAND2BX1 U7135 ( .AN(n3000), .B(n8638), .Y(n7509) );
  NAND2BX1 U7136 ( .AN(n3001), .B(n8606), .Y(n7507) );
  NAND2BX1 U7137 ( .AN(n2163), .B(n8670), .Y(n7510) );
  NAND4X1 U7138 ( .A(n7139), .B(n7138), .C(n7137), .D(n7136), .Y(n8419) );
  NAND2BX1 U7139 ( .AN(n2163), .B(n8669), .Y(n7139) );
  NAND4X1 U7140 ( .A(n7163), .B(n7162), .C(n7161), .D(n7160), .Y(n8050) );
  NAND2BX1 U7141 ( .AN(n2163), .B(n8668), .Y(n7163) );
  NAND4X1 U7142 ( .A(n7090), .B(n7089), .C(n7088), .D(n7087), .Y(n8031) );
  NAND2BX1 U7143 ( .AN(n3000), .B(n8635), .Y(n7089) );
  NAND2BX1 U7144 ( .AN(n3001), .B(n8603), .Y(n7087) );
  NAND2BX1 U7145 ( .AN(n2163), .B(n8667), .Y(n7090) );
  NAND4X1 U7146 ( .A(n7115), .B(n7114), .C(n7113), .D(n7112), .Y(n8004) );
  NAND2BX1 U7147 ( .AN(n2163), .B(n8666), .Y(n7115) );
  NAND4X1 U7148 ( .A(n7438), .B(n7437), .C(n7436), .D(n7435), .Y(n8179) );
  NAND2BX1 U7149 ( .AN(n3000), .B(n8642), .Y(n7437) );
  NAND4X1 U7150 ( .A(n8137), .B(n8136), .C(n8135), .D(n8134), .Y(n8456) );
  NAND2BX1 U7151 ( .AN(n3000), .B(n8640), .Y(n8136) );
  NAND4X1 U7152 ( .A(n7660), .B(n7659), .C(n7658), .D(n7657), .Y(n8201) );
  NAND2BX1 U7153 ( .AN(n3000), .B(n8643), .Y(n7659) );
  NAND2BX1 U7154 ( .AN(n3001), .B(n8611), .Y(n7657) );
  NAND2BX1 U7155 ( .AN(n2163), .B(n8675), .Y(n7660) );
  NAND4X1 U7156 ( .A(n7462), .B(n7461), .C(n7460), .D(n7459), .Y(n8153) );
  NAND2BX1 U7157 ( .AN(n3000), .B(n8641), .Y(n7461) );
  NAND4X1 U7158 ( .A(n7486), .B(n7485), .C(n7484), .D(n7483), .Y(n8094) );
  NAND2BX1 U7159 ( .AN(n3000), .B(n8639), .Y(n7485) );
  NAND2BX1 U7160 ( .AN(n3001), .B(n8607), .Y(n7483) );
  NAND2BX1 U7161 ( .AN(n2163), .B(n8671), .Y(n7486) );
  AND2X2 U7162 ( .A(n4536), .B(n3051), .Y(n8453) );
  OAI21XL U7163 ( .A0(n8392), .A1(n4537), .B0(n4538), .Y(n4536) );
  NAND2BX1 U7164 ( .AN(n3001), .B(n8605), .Y(n7136) );
  NAND2BX1 U7165 ( .AN(n3001), .B(n8604), .Y(n7160) );
  NAND2BX1 U7166 ( .AN(n3001), .B(n8602), .Y(n7112) );
  CLKINVX1 U7167 ( .A(n3051), .Y(n8682) );
  AND2X2 U7168 ( .A(n7306), .B(n2995), .Y(n2882) );
  AND2X2 U7169 ( .A(n2882), .B(\i_MIPS/n332 ), .Y(n2883) );
  CLKINVX1 U7170 ( .A(\D_cache/n214 ), .Y(n3976) );
  NAND2X1 U7171 ( .A(\i_MIPS/Register/n119 ), .B(\i_MIPS/Register/n104 ), .Y(
        \i_MIPS/Register/n118 ) );
  NAND2X1 U7172 ( .A(\i_MIPS/Register/n117 ), .B(\i_MIPS/Register/n104 ), .Y(
        \i_MIPS/Register/n116 ) );
  NAND2X1 U7173 ( .A(\i_MIPS/Register/n115 ), .B(\i_MIPS/Register/n104 ), .Y(
        \i_MIPS/Register/n114 ) );
  NAND2X1 U7174 ( .A(\i_MIPS/Register/n113 ), .B(\i_MIPS/Register/n104 ), .Y(
        \i_MIPS/Register/n112 ) );
  NAND2X1 U7175 ( .A(\i_MIPS/Register/n111 ), .B(\i_MIPS/Register/n104 ), .Y(
        \i_MIPS/Register/n110 ) );
  NAND2X1 U7176 ( .A(\i_MIPS/Register/n109 ), .B(\i_MIPS/Register/n104 ), .Y(
        \i_MIPS/Register/n108 ) );
  NAND2X1 U7177 ( .A(\i_MIPS/Register/n107 ), .B(\i_MIPS/Register/n104 ), .Y(
        \i_MIPS/Register/n106 ) );
  NAND2X1 U7178 ( .A(\i_MIPS/Control_ID/n15 ), .B(\i_MIPS/Control_ID/n10 ), 
        .Y(\i_MIPS/control_out[7] ) );
  CLKBUFX3 U7179 ( .A(n4376), .Y(n4386) );
  AOI2BB2X2 U7180 ( .B0(\D_cache/N121 ), .B1(n3945), .A0N(n3947), .A1N(
        \D_cache/n386 ), .Y(\D_cache/n385 ) );
  AOI222XL U7181 ( .A0(\D_cache/N121 ), .A1(\D_cache/n387 ), .B0(
        \D_cache/n388 ), .B1(n10324), .C0(mem_rdata_D[95]), .C1(n3982), .Y(
        \D_cache/n386 ) );
  AOI2BB2X2 U7182 ( .B0(\D_cache/N122 ), .B1(n3945), .A0N(n3947), .A1N(
        \D_cache/n390 ), .Y(\D_cache/n389 ) );
  AOI222XL U7183 ( .A0(\D_cache/N122 ), .A1(n3992), .B0(n3994), .B1(n10325), 
        .C0(mem_rdata_D[94]), .C1(n3982), .Y(\D_cache/n390 ) );
  AOI2BB2X2 U7184 ( .B0(\D_cache/N123 ), .B1(n3946), .A0N(n3947), .A1N(
        \D_cache/n392 ), .Y(\D_cache/n391 ) );
  AOI222XL U7185 ( .A0(\D_cache/N123 ), .A1(n3992), .B0(n3993), .B1(n10326), 
        .C0(mem_rdata_D[93]), .C1(n3982), .Y(\D_cache/n392 ) );
  AOI2BB2X2 U7186 ( .B0(\D_cache/N124 ), .B1(n3945), .A0N(n3947), .A1N(
        \D_cache/n394 ), .Y(\D_cache/n393 ) );
  AOI222XL U7187 ( .A0(\D_cache/N124 ), .A1(n3992), .B0(n3994), .B1(n10327), 
        .C0(mem_rdata_D[92]), .C1(n3982), .Y(\D_cache/n394 ) );
  AOI2BB2X2 U7188 ( .B0(\D_cache/N125 ), .B1(n3946), .A0N(n3948), .A1N(
        \D_cache/n396 ), .Y(\D_cache/n395 ) );
  AOI222XL U7189 ( .A0(\D_cache/N125 ), .A1(n3992), .B0(n3993), .B1(n10328), 
        .C0(mem_rdata_D[91]), .C1(n3982), .Y(\D_cache/n396 ) );
  AOI2BB2X2 U7190 ( .B0(\D_cache/N126 ), .B1(n3946), .A0N(n3947), .A1N(
        \D_cache/n398 ), .Y(\D_cache/n397 ) );
  AOI222XL U7191 ( .A0(\D_cache/N126 ), .A1(n3992), .B0(n3994), .B1(n10329), 
        .C0(mem_rdata_D[90]), .C1(n3982), .Y(\D_cache/n398 ) );
  AOI2BB2X2 U7192 ( .B0(\D_cache/N127 ), .B1(n3945), .A0N(n3947), .A1N(
        \D_cache/n400 ), .Y(\D_cache/n399 ) );
  AOI222XL U7193 ( .A0(\D_cache/N127 ), .A1(n3992), .B0(n3994), .B1(n10330), 
        .C0(mem_rdata_D[89]), .C1(n3982), .Y(\D_cache/n400 ) );
  AOI2BB2X2 U7194 ( .B0(\D_cache/N128 ), .B1(n3945), .A0N(n3949), .A1N(
        \D_cache/n402 ), .Y(\D_cache/n401 ) );
  AOI222XL U7195 ( .A0(\D_cache/N128 ), .A1(n3992), .B0(n3994), .B1(n10331), 
        .C0(mem_rdata_D[88]), .C1(n3982), .Y(\D_cache/n402 ) );
  AOI2BB2X2 U7196 ( .B0(\D_cache/N129 ), .B1(n3947), .A0N(n3949), .A1N(
        \D_cache/n404 ), .Y(\D_cache/n403 ) );
  AOI222XL U7197 ( .A0(\D_cache/N129 ), .A1(n3992), .B0(n3994), .B1(n10332), 
        .C0(mem_rdata_D[87]), .C1(n3982), .Y(\D_cache/n404 ) );
  AOI2BB2X2 U7198 ( .B0(\D_cache/N130 ), .B1(n3947), .A0N(n3949), .A1N(
        \D_cache/n406 ), .Y(\D_cache/n405 ) );
  AOI222XL U7199 ( .A0(\D_cache/N130 ), .A1(n3992), .B0(n3994), .B1(n10333), 
        .C0(mem_rdata_D[86]), .C1(n3982), .Y(\D_cache/n406 ) );
  AOI2BB2X2 U7200 ( .B0(\D_cache/N131 ), .B1(n3946), .A0N(n3948), .A1N(
        \D_cache/n408 ), .Y(\D_cache/n407 ) );
  AOI222XL U7201 ( .A0(\D_cache/N131 ), .A1(n3992), .B0(n3994), .B1(n10334), 
        .C0(mem_rdata_D[85]), .C1(n3983), .Y(\D_cache/n408 ) );
  AOI2BB2X2 U7202 ( .B0(\D_cache/N132 ), .B1(n3947), .A0N(n3949), .A1N(
        \D_cache/n410 ), .Y(\D_cache/n409 ) );
  AOI222XL U7203 ( .A0(\D_cache/N132 ), .A1(n3992), .B0(n3994), .B1(n10335), 
        .C0(mem_rdata_D[84]), .C1(n3983), .Y(\D_cache/n410 ) );
  AOI2BB2X2 U7204 ( .B0(\D_cache/N133 ), .B1(n3947), .A0N(n3949), .A1N(
        \D_cache/n412 ), .Y(\D_cache/n411 ) );
  AOI222XL U7205 ( .A0(\D_cache/N133 ), .A1(n3992), .B0(n3994), .B1(n10336), 
        .C0(mem_rdata_D[83]), .C1(n3983), .Y(\D_cache/n412 ) );
  AOI2BB2X2 U7206 ( .B0(\D_cache/N134 ), .B1(n3946), .A0N(n3949), .A1N(
        \D_cache/n414 ), .Y(\D_cache/n413 ) );
  AOI222XL U7207 ( .A0(\D_cache/N134 ), .A1(n3992), .B0(n3994), .B1(n10337), 
        .C0(mem_rdata_D[82]), .C1(n3983), .Y(\D_cache/n414 ) );
  AOI2BB2X2 U7208 ( .B0(\D_cache/N135 ), .B1(n3946), .A0N(n3948), .A1N(
        \D_cache/n416 ), .Y(\D_cache/n415 ) );
  AOI222XL U7209 ( .A0(\D_cache/N135 ), .A1(n3992), .B0(n3994), .B1(n10338), 
        .C0(mem_rdata_D[81]), .C1(n3983), .Y(\D_cache/n416 ) );
  AOI2BB2X2 U7210 ( .B0(\D_cache/N136 ), .B1(n3945), .A0N(n3949), .A1N(
        \D_cache/n418 ), .Y(\D_cache/n417 ) );
  AOI222XL U7211 ( .A0(\D_cache/N136 ), .A1(n3992), .B0(n3994), .B1(n10339), 
        .C0(mem_rdata_D[80]), .C1(n3983), .Y(\D_cache/n418 ) );
  AOI2BB2X2 U7212 ( .B0(\D_cache/N137 ), .B1(n3946), .A0N(n3949), .A1N(
        \D_cache/n420 ), .Y(\D_cache/n419 ) );
  AOI222XL U7213 ( .A0(\D_cache/N137 ), .A1(n3992), .B0(n3994), .B1(n10340), 
        .C0(mem_rdata_D[79]), .C1(n3983), .Y(\D_cache/n420 ) );
  AOI2BB2X2 U7214 ( .B0(\D_cache/N138 ), .B1(n3947), .A0N(n3948), .A1N(
        \D_cache/n422 ), .Y(\D_cache/n421 ) );
  AOI222XL U7215 ( .A0(\D_cache/N138 ), .A1(n3992), .B0(n3994), .B1(n10341), 
        .C0(mem_rdata_D[78]), .C1(n3983), .Y(\D_cache/n422 ) );
  AOI2BB2X2 U7216 ( .B0(\D_cache/N139 ), .B1(n3947), .A0N(n3949), .A1N(
        \D_cache/n424 ), .Y(\D_cache/n423 ) );
  AOI222XL U7217 ( .A0(\D_cache/N139 ), .A1(n3992), .B0(n3994), .B1(n10342), 
        .C0(mem_rdata_D[77]), .C1(n3983), .Y(\D_cache/n424 ) );
  AOI2BB2X2 U7218 ( .B0(\D_cache/N140 ), .B1(n3946), .A0N(n3948), .A1N(
        \D_cache/n426 ), .Y(\D_cache/n425 ) );
  AOI222XL U7219 ( .A0(\D_cache/N140 ), .A1(n3992), .B0(n3993), .B1(n10343), 
        .C0(mem_rdata_D[76]), .C1(n3983), .Y(\D_cache/n426 ) );
  AOI2BB2X2 U7220 ( .B0(\D_cache/N141 ), .B1(n3947), .A0N(n3948), .A1N(
        \D_cache/n428 ), .Y(\D_cache/n427 ) );
  AOI222XL U7221 ( .A0(\D_cache/N141 ), .A1(\D_cache/n387 ), .B0(n3993), .B1(
        n10344), .C0(mem_rdata_D[75]), .C1(n3983), .Y(\D_cache/n428 ) );
  AOI2BB2X2 U7222 ( .B0(\D_cache/N142 ), .B1(n3945), .A0N(n3948), .A1N(
        \D_cache/n430 ), .Y(\D_cache/n429 ) );
  AOI222XL U7223 ( .A0(\D_cache/N142 ), .A1(\D_cache/n387 ), .B0(n3993), .B1(
        n10345), .C0(mem_rdata_D[74]), .C1(n3983), .Y(\D_cache/n430 ) );
  AOI2BB2X2 U7224 ( .B0(\D_cache/N143 ), .B1(n3945), .A0N(n3948), .A1N(
        \D_cache/n432 ), .Y(\D_cache/n431 ) );
  AOI222XL U7225 ( .A0(\D_cache/N143 ), .A1(\D_cache/n387 ), .B0(n3993), .B1(
        n10346), .C0(mem_rdata_D[73]), .C1(n3983), .Y(\D_cache/n432 ) );
  AOI2BB2X2 U7226 ( .B0(\D_cache/N144 ), .B1(n3945), .A0N(n3948), .A1N(
        \D_cache/n434 ), .Y(\D_cache/n433 ) );
  AOI222XL U7227 ( .A0(\D_cache/N144 ), .A1(\D_cache/n387 ), .B0(n3993), .B1(
        n10347), .C0(mem_rdata_D[72]), .C1(n3983), .Y(\D_cache/n434 ) );
  AOI2BB2X2 U7228 ( .B0(\D_cache/N145 ), .B1(n3947), .A0N(n3948), .A1N(
        \D_cache/n436 ), .Y(\D_cache/n435 ) );
  AOI222XL U7229 ( .A0(\D_cache/N145 ), .A1(n3992), .B0(n3993), .B1(n10348), 
        .C0(mem_rdata_D[71]), .C1(n3983), .Y(\D_cache/n436 ) );
  AOI2BB2X2 U7230 ( .B0(\D_cache/N146 ), .B1(n3945), .A0N(n3948), .A1N(
        \D_cache/n438 ), .Y(\D_cache/n437 ) );
  AOI222XL U7231 ( .A0(\D_cache/N146 ), .A1(\D_cache/n387 ), .B0(n3993), .B1(
        n10349), .C0(mem_rdata_D[70]), .C1(n3984), .Y(\D_cache/n438 ) );
  AOI2BB2X2 U7232 ( .B0(\D_cache/N147 ), .B1(n3946), .A0N(n3948), .A1N(
        \D_cache/n440 ), .Y(\D_cache/n439 ) );
  AOI222XL U7233 ( .A0(\D_cache/N147 ), .A1(\D_cache/n387 ), .B0(n3993), .B1(
        n10350), .C0(mem_rdata_D[69]), .C1(n3984), .Y(\D_cache/n440 ) );
  AOI2BB2X2 U7234 ( .B0(\D_cache/N148 ), .B1(n3946), .A0N(n3948), .A1N(
        \D_cache/n442 ), .Y(\D_cache/n441 ) );
  AOI222XL U7235 ( .A0(\D_cache/N148 ), .A1(\D_cache/n387 ), .B0(n3993), .B1(
        n10351), .C0(mem_rdata_D[68]), .C1(n3984), .Y(\D_cache/n442 ) );
  AOI2BB2X2 U7236 ( .B0(\D_cache/N149 ), .B1(n3945), .A0N(n3948), .A1N(
        \D_cache/n444 ), .Y(\D_cache/n443 ) );
  AOI222XL U7237 ( .A0(\D_cache/N149 ), .A1(\D_cache/n387 ), .B0(n3993), .B1(
        n10352), .C0(mem_rdata_D[67]), .C1(n3984), .Y(\D_cache/n444 ) );
  AOI2BB2X2 U7238 ( .B0(\D_cache/N150 ), .B1(n3946), .A0N(n3948), .A1N(
        \D_cache/n446 ), .Y(\D_cache/n445 ) );
  AOI222XL U7239 ( .A0(\D_cache/N150 ), .A1(\D_cache/n387 ), .B0(n3993), .B1(
        n10353), .C0(mem_rdata_D[66]), .C1(n3984), .Y(\D_cache/n446 ) );
  AOI2BB2X2 U7240 ( .B0(\D_cache/N151 ), .B1(n3946), .A0N(n3948), .A1N(
        \D_cache/n448 ), .Y(\D_cache/n447 ) );
  AOI222XL U7241 ( .A0(\D_cache/N151 ), .A1(\D_cache/n387 ), .B0(n3993), .B1(
        n10354), .C0(mem_rdata_D[65]), .C1(n3984), .Y(\D_cache/n448 ) );
  AOI2BB2X2 U7242 ( .B0(\D_cache/N152 ), .B1(n3945), .A0N(n3948), .A1N(
        \D_cache/n450 ), .Y(\D_cache/n449 ) );
  AOI222XL U7243 ( .A0(\D_cache/N152 ), .A1(\D_cache/n387 ), .B0(n3993), .B1(
        n10355), .C0(mem_rdata_D[64]), .C1(n3984), .Y(\D_cache/n450 ) );
  OA22X2 U7244 ( .A0(n8759), .A1(n3967), .B0(n3950), .B1(\D_cache/n318 ), .Y(
        \D_cache/n317 ) );
  AOI222XL U7245 ( .A0(\D_cache/N89 ), .A1(\D_cache/n319 ), .B0(\D_cache/n320 ), .B1(n10324), .C0(mem_rdata_D[63]), .C1(n3983), .Y(\D_cache/n318 ) );
  OA22X2 U7246 ( .A0(n8760), .A1(n3966), .B0(n3949), .B1(\D_cache/n322 ), .Y(
        \D_cache/n321 ) );
  AOI222XL U7247 ( .A0(\D_cache/N90 ), .A1(\D_cache/n319 ), .B0(n3990), .B1(
        n10325), .C0(mem_rdata_D[62]), .C1(n3983), .Y(\D_cache/n322 ) );
  OA22X2 U7248 ( .A0(n8761), .A1(n3961), .B0(n3949), .B1(\D_cache/n324 ), .Y(
        \D_cache/n323 ) );
  AOI222XL U7249 ( .A0(\D_cache/N91 ), .A1(n3989), .B0(n3991), .B1(n10326), 
        .C0(mem_rdata_D[61]), .C1(n3984), .Y(\D_cache/n324 ) );
  OA22X2 U7250 ( .A0(n8762), .A1(n3961), .B0(n3950), .B1(\D_cache/n326 ), .Y(
        \D_cache/n325 ) );
  AOI222XL U7251 ( .A0(\D_cache/N92 ), .A1(n3989), .B0(n3990), .B1(n10327), 
        .C0(mem_rdata_D[60]), .C1(n3984), .Y(\D_cache/n326 ) );
  OA22X2 U7252 ( .A0(n8763), .A1(n3961), .B0(n3950), .B1(\D_cache/n328 ), .Y(
        \D_cache/n327 ) );
  AOI222XL U7253 ( .A0(\D_cache/N93 ), .A1(n3989), .B0(n3991), .B1(n10328), 
        .C0(mem_rdata_D[59]), .C1(n3979), .Y(\D_cache/n328 ) );
  OA22X2 U7254 ( .A0(n8764), .A1(n3961), .B0(n3949), .B1(\D_cache/n330 ), .Y(
        \D_cache/n329 ) );
  AOI222XL U7255 ( .A0(\D_cache/N94 ), .A1(n3989), .B0(n3990), .B1(n10329), 
        .C0(mem_rdata_D[58]), .C1(n3979), .Y(\D_cache/n330 ) );
  OA22X2 U7256 ( .A0(n8765), .A1(n3961), .B0(n3952), .B1(\D_cache/n332 ), .Y(
        \D_cache/n331 ) );
  AOI222XL U7257 ( .A0(\D_cache/N95 ), .A1(n3989), .B0(n3991), .B1(n10330), 
        .C0(mem_rdata_D[57]), .C1(n3984), .Y(\D_cache/n332 ) );
  OA22X2 U7258 ( .A0(n8766), .A1(n3961), .B0(n3949), .B1(\D_cache/n334 ), .Y(
        \D_cache/n333 ) );
  AOI222XL U7259 ( .A0(\D_cache/N96 ), .A1(n3989), .B0(n3991), .B1(n10331), 
        .C0(mem_rdata_D[56]), .C1(n3982), .Y(\D_cache/n334 ) );
  OA22X2 U7260 ( .A0(n8767), .A1(n3962), .B0(n3949), .B1(\D_cache/n336 ), .Y(
        \D_cache/n335 ) );
  AOI222XL U7261 ( .A0(\D_cache/N97 ), .A1(n3989), .B0(n3991), .B1(n10332), 
        .C0(mem_rdata_D[55]), .C1(n3983), .Y(\D_cache/n336 ) );
  OA22X2 U7262 ( .A0(n8768), .A1(n3962), .B0(n3950), .B1(\D_cache/n338 ), .Y(
        \D_cache/n337 ) );
  AOI222XL U7263 ( .A0(\D_cache/N98 ), .A1(n3989), .B0(n3991), .B1(n10333), 
        .C0(mem_rdata_D[54]), .C1(n3979), .Y(\D_cache/n338 ) );
  OA22X2 U7264 ( .A0(n8769), .A1(n3962), .B0(n3949), .B1(\D_cache/n340 ), .Y(
        \D_cache/n339 ) );
  AOI222XL U7265 ( .A0(\D_cache/N99 ), .A1(n3989), .B0(n3991), .B1(n10334), 
        .C0(mem_rdata_D[53]), .C1(n3984), .Y(\D_cache/n340 ) );
  OA22X2 U7266 ( .A0(n8770), .A1(n3962), .B0(n3950), .B1(\D_cache/n342 ), .Y(
        \D_cache/n341 ) );
  AOI222XL U7267 ( .A0(\D_cache/N100 ), .A1(n3989), .B0(n3991), .B1(n10335), 
        .C0(mem_rdata_D[52]), .C1(n3982), .Y(\D_cache/n342 ) );
  OA22X2 U7268 ( .A0(n8771), .A1(n3962), .B0(n3950), .B1(\D_cache/n344 ), .Y(
        \D_cache/n343 ) );
  AOI222XL U7269 ( .A0(\D_cache/N101 ), .A1(n3989), .B0(n3991), .B1(n10336), 
        .C0(mem_rdata_D[51]), .C1(n3981), .Y(\D_cache/n344 ) );
  OA22X2 U7270 ( .A0(n8852), .A1(n3962), .B0(n3949), .B1(\D_cache/n346 ), .Y(
        \D_cache/n345 ) );
  AOI222XL U7271 ( .A0(\D_cache/N102 ), .A1(n3989), .B0(n3991), .B1(n10337), 
        .C0(mem_rdata_D[50]), .C1(n3981), .Y(\D_cache/n346 ) );
  OA22X2 U7272 ( .A0(n8853), .A1(n3963), .B0(n3950), .B1(\D_cache/n348 ), .Y(
        \D_cache/n347 ) );
  AOI222XL U7273 ( .A0(\D_cache/N103 ), .A1(n3989), .B0(n3991), .B1(n10338), 
        .C0(mem_rdata_D[49]), .C1(n3981), .Y(\D_cache/n348 ) );
  OA22X2 U7274 ( .A0(n8854), .A1(n3963), .B0(n3952), .B1(\D_cache/n350 ), .Y(
        \D_cache/n349 ) );
  AOI222XL U7275 ( .A0(\D_cache/N104 ), .A1(n3989), .B0(n3991), .B1(n10339), 
        .C0(mem_rdata_D[48]), .C1(n3981), .Y(\D_cache/n350 ) );
  OA22X2 U7276 ( .A0(n8855), .A1(n3963), .B0(n3952), .B1(\D_cache/n352 ), .Y(
        \D_cache/n351 ) );
  AOI222XL U7277 ( .A0(\D_cache/N105 ), .A1(n3989), .B0(n3991), .B1(n10340), 
        .C0(mem_rdata_D[47]), .C1(n3981), .Y(\D_cache/n352 ) );
  OA22X2 U7278 ( .A0(n8856), .A1(n3963), .B0(n3952), .B1(\D_cache/n354 ), .Y(
        \D_cache/n353 ) );
  AOI222XL U7279 ( .A0(\D_cache/N106 ), .A1(n3989), .B0(n3991), .B1(n10341), 
        .C0(mem_rdata_D[46]), .C1(n3981), .Y(\D_cache/n354 ) );
  OA22X2 U7280 ( .A0(n8857), .A1(n3963), .B0(n3952), .B1(\D_cache/n356 ), .Y(
        \D_cache/n355 ) );
  AOI222XL U7281 ( .A0(\D_cache/N107 ), .A1(n3989), .B0(n3991), .B1(n10342), 
        .C0(mem_rdata_D[45]), .C1(n3981), .Y(\D_cache/n356 ) );
  OA22X2 U7282 ( .A0(n8858), .A1(n3964), .B0(n3952), .B1(\D_cache/n358 ), .Y(
        \D_cache/n357 ) );
  AOI222XL U7283 ( .A0(\D_cache/N108 ), .A1(n3989), .B0(n3990), .B1(n10343), 
        .C0(mem_rdata_D[44]), .C1(n3981), .Y(\D_cache/n358 ) );
  OA22X2 U7284 ( .A0(n8859), .A1(n3964), .B0(n3952), .B1(\D_cache/n360 ), .Y(
        \D_cache/n359 ) );
  AOI222XL U7285 ( .A0(\D_cache/N109 ), .A1(n3989), .B0(n3990), .B1(n10344), 
        .C0(mem_rdata_D[43]), .C1(n3981), .Y(\D_cache/n360 ) );
  OA22X2 U7286 ( .A0(n8860), .A1(n3964), .B0(n3952), .B1(\D_cache/n362 ), .Y(
        \D_cache/n361 ) );
  AOI222XL U7287 ( .A0(\D_cache/N110 ), .A1(n3989), .B0(n3990), .B1(n10345), 
        .C0(mem_rdata_D[42]), .C1(n3981), .Y(\D_cache/n362 ) );
  OA22X2 U7288 ( .A0(n8861), .A1(n3964), .B0(n3952), .B1(\D_cache/n364 ), .Y(
        \D_cache/n363 ) );
  AOI222XL U7289 ( .A0(\D_cache/N111 ), .A1(\D_cache/n319 ), .B0(n3990), .B1(
        n10346), .C0(mem_rdata_D[41]), .C1(n3981), .Y(\D_cache/n364 ) );
  OA22X2 U7290 ( .A0(n8862), .A1(n3964), .B0(n3952), .B1(\D_cache/n366 ), .Y(
        \D_cache/n365 ) );
  AOI222XL U7291 ( .A0(\D_cache/N112 ), .A1(\D_cache/n319 ), .B0(n3990), .B1(
        n10347), .C0(mem_rdata_D[40]), .C1(n3981), .Y(\D_cache/n366 ) );
  OA22X2 U7292 ( .A0(n8863), .A1(n3964), .B0(n3952), .B1(\D_cache/n368 ), .Y(
        \D_cache/n367 ) );
  AOI222XL U7293 ( .A0(\D_cache/N113 ), .A1(\D_cache/n319 ), .B0(n3990), .B1(
        n10348), .C0(mem_rdata_D[39]), .C1(n3981), .Y(\D_cache/n368 ) );
  OA22X2 U7294 ( .A0(n8864), .A1(n3965), .B0(n3952), .B1(\D_cache/n370 ), .Y(
        \D_cache/n369 ) );
  AOI222XL U7295 ( .A0(\D_cache/N114 ), .A1(\D_cache/n319 ), .B0(n3990), .B1(
        n10349), .C0(mem_rdata_D[38]), .C1(n3981), .Y(\D_cache/n370 ) );
  OA22X2 U7296 ( .A0(n8865), .A1(n3965), .B0(n3952), .B1(\D_cache/n372 ), .Y(
        \D_cache/n371 ) );
  AOI222XL U7297 ( .A0(\D_cache/N115 ), .A1(\D_cache/n319 ), .B0(n3990), .B1(
        n10350), .C0(mem_rdata_D[37]), .C1(n3981), .Y(\D_cache/n372 ) );
  OA22X2 U7298 ( .A0(n8866), .A1(n3965), .B0(n3952), .B1(\D_cache/n374 ), .Y(
        \D_cache/n373 ) );
  AOI222XL U7299 ( .A0(\D_cache/N116 ), .A1(\D_cache/n319 ), .B0(n3990), .B1(
        n10351), .C0(mem_rdata_D[36]), .C1(n3982), .Y(\D_cache/n374 ) );
  OA22X2 U7300 ( .A0(n8867), .A1(n3965), .B0(n3953), .B1(\D_cache/n376 ), .Y(
        \D_cache/n375 ) );
  AOI222XL U7301 ( .A0(\D_cache/N117 ), .A1(\D_cache/n319 ), .B0(n3990), .B1(
        n10352), .C0(mem_rdata_D[35]), .C1(n3982), .Y(\D_cache/n376 ) );
  OA22X2 U7302 ( .A0(n8868), .A1(n3965), .B0(n3953), .B1(\D_cache/n378 ), .Y(
        \D_cache/n377 ) );
  AOI222XL U7303 ( .A0(\D_cache/N118 ), .A1(\D_cache/n319 ), .B0(n3990), .B1(
        n10353), .C0(mem_rdata_D[34]), .C1(n3982), .Y(\D_cache/n378 ) );
  OA22X2 U7304 ( .A0(n8869), .A1(n3965), .B0(n3953), .B1(\D_cache/n380 ), .Y(
        \D_cache/n379 ) );
  AOI222XL U7305 ( .A0(\D_cache/N119 ), .A1(\D_cache/n319 ), .B0(n3990), .B1(
        n10354), .C0(mem_rdata_D[33]), .C1(n3982), .Y(\D_cache/n380 ) );
  OA22X2 U7306 ( .A0(n8870), .A1(n3966), .B0(n3953), .B1(\D_cache/n382 ), .Y(
        \D_cache/n381 ) );
  AOI222XL U7307 ( .A0(\D_cache/N120 ), .A1(\D_cache/n319 ), .B0(n3990), .B1(
        n10355), .C0(mem_rdata_D[32]), .C1(n3982), .Y(\D_cache/n382 ) );
  OA22X2 U7308 ( .A0(n8871), .A1(n3966), .B0(n3953), .B1(\D_cache/n453 ), .Y(
        \D_cache/n452 ) );
  AOI222XL U7309 ( .A0(\D_cache/N153 ), .A1(\D_cache/n454 ), .B0(n3997), .B1(
        n10324), .C0(mem_rdata_D[127]), .C1(n3984), .Y(\D_cache/n453 ) );
  OA22X2 U7310 ( .A0(n8872), .A1(n3966), .B0(n3953), .B1(\D_cache/n457 ), .Y(
        \D_cache/n456 ) );
  AOI222XL U7311 ( .A0(\D_cache/N154 ), .A1(\D_cache/n454 ), .B0(n3997), .B1(
        n10325), .C0(mem_rdata_D[126]), .C1(n3984), .Y(\D_cache/n457 ) );
  OA22X2 U7312 ( .A0(n8873), .A1(n3966), .B0(n3953), .B1(\D_cache/n459 ), .Y(
        \D_cache/n458 ) );
  AOI222XL U7313 ( .A0(\D_cache/N155 ), .A1(n3995), .B0(n3997), .B1(n10326), 
        .C0(mem_rdata_D[125]), .C1(n3984), .Y(\D_cache/n459 ) );
  OA22X2 U7314 ( .A0(n8874), .A1(n3966), .B0(n3953), .B1(\D_cache/n461 ), .Y(
        \D_cache/n460 ) );
  AOI222XL U7315 ( .A0(\D_cache/N156 ), .A1(n3995), .B0(n3997), .B1(n10327), 
        .C0(mem_rdata_D[124]), .C1(n3984), .Y(\D_cache/n461 ) );
  OA22X2 U7316 ( .A0(n8875), .A1(n3966), .B0(n3953), .B1(\D_cache/n463 ), .Y(
        \D_cache/n462 ) );
  AOI222XL U7317 ( .A0(\D_cache/N157 ), .A1(n3995), .B0(n3997), .B1(n10328), 
        .C0(mem_rdata_D[123]), .C1(n3984), .Y(\D_cache/n463 ) );
  OA22X2 U7318 ( .A0(n8876), .A1(n3967), .B0(n3953), .B1(\D_cache/n465 ), .Y(
        \D_cache/n464 ) );
  AOI222XL U7319 ( .A0(\D_cache/N158 ), .A1(n3995), .B0(n3997), .B1(n10329), 
        .C0(mem_rdata_D[122]), .C1(n3984), .Y(\D_cache/n465 ) );
  OA22X2 U7320 ( .A0(n8877), .A1(n3967), .B0(n3953), .B1(\D_cache/n467 ), .Y(
        \D_cache/n466 ) );
  AOI222XL U7321 ( .A0(\D_cache/N159 ), .A1(n3995), .B0(n3997), .B1(n10330), 
        .C0(mem_rdata_D[121]), .C1(n3984), .Y(\D_cache/n467 ) );
  OA22X2 U7322 ( .A0(n8878), .A1(n3967), .B0(n3953), .B1(\D_cache/n469 ), .Y(
        \D_cache/n468 ) );
  AOI222XL U7323 ( .A0(\D_cache/N160 ), .A1(n3995), .B0(n3997), .B1(n10331), 
        .C0(mem_rdata_D[120]), .C1(n3984), .Y(\D_cache/n469 ) );
  OA22X2 U7324 ( .A0(n8879), .A1(n3967), .B0(n3953), .B1(\D_cache/n471 ), .Y(
        \D_cache/n470 ) );
  AOI222XL U7325 ( .A0(\D_cache/N161 ), .A1(n3995), .B0(n3997), .B1(n10332), 
        .C0(mem_rdata_D[119]), .C1(n3985), .Y(\D_cache/n471 ) );
  OA22X2 U7326 ( .A0(n8880), .A1(n3967), .B0(n3953), .B1(\D_cache/n473 ), .Y(
        \D_cache/n472 ) );
  AOI222XL U7327 ( .A0(\D_cache/N162 ), .A1(n3995), .B0(n3997), .B1(n10333), 
        .C0(mem_rdata_D[118]), .C1(n3985), .Y(\D_cache/n473 ) );
  OA22X2 U7328 ( .A0(n8881), .A1(n3967), .B0(n3953), .B1(\D_cache/n475 ), .Y(
        \D_cache/n474 ) );
  AOI222XL U7329 ( .A0(\D_cache/N163 ), .A1(n3995), .B0(n3997), .B1(n10334), 
        .C0(mem_rdata_D[117]), .C1(n3985), .Y(\D_cache/n475 ) );
  OA22X2 U7330 ( .A0(n8882), .A1(n3969), .B0(n3953), .B1(\D_cache/n477 ), .Y(
        \D_cache/n476 ) );
  AOI222XL U7331 ( .A0(\D_cache/N164 ), .A1(n3995), .B0(n3997), .B1(n10335), 
        .C0(mem_rdata_D[116]), .C1(n3985), .Y(\D_cache/n477 ) );
  OA22X2 U7332 ( .A0(n8883), .A1(n3966), .B0(n3953), .B1(\D_cache/n479 ), .Y(
        \D_cache/n478 ) );
  AOI222XL U7333 ( .A0(\D_cache/N165 ), .A1(n3995), .B0(n3997), .B1(n10336), 
        .C0(mem_rdata_D[115]), .C1(n3985), .Y(\D_cache/n479 ) );
  OA22X2 U7334 ( .A0(n8884), .A1(n3967), .B0(n3953), .B1(\D_cache/n481 ), .Y(
        \D_cache/n480 ) );
  AOI222XL U7335 ( .A0(\D_cache/N166 ), .A1(n3995), .B0(n3997), .B1(n10337), 
        .C0(mem_rdata_D[114]), .C1(n3985), .Y(\D_cache/n481 ) );
  OA22X2 U7336 ( .A0(n8885), .A1(n3965), .B0(n3954), .B1(\D_cache/n483 ), .Y(
        \D_cache/n482 ) );
  AOI222XL U7337 ( .A0(\D_cache/N167 ), .A1(n3995), .B0(n3997), .B1(n10338), 
        .C0(mem_rdata_D[113]), .C1(n3985), .Y(\D_cache/n483 ) );
  OA22X2 U7338 ( .A0(n8886), .A1(n3964), .B0(n3954), .B1(\D_cache/n485 ), .Y(
        \D_cache/n484 ) );
  AOI222XL U7339 ( .A0(\D_cache/N168 ), .A1(n3995), .B0(n3997), .B1(n10339), 
        .C0(mem_rdata_D[112]), .C1(n3985), .Y(\D_cache/n485 ) );
  OA22X2 U7340 ( .A0(n8887), .A1(n3969), .B0(n3954), .B1(\D_cache/n487 ), .Y(
        \D_cache/n486 ) );
  AOI222XL U7341 ( .A0(\D_cache/N169 ), .A1(n3995), .B0(n3997), .B1(n10340), 
        .C0(mem_rdata_D[111]), .C1(n3985), .Y(\D_cache/n487 ) );
  OA22X2 U7342 ( .A0(n8888), .A1(n3968), .B0(n3954), .B1(\D_cache/n489 ), .Y(
        \D_cache/n488 ) );
  AOI222XL U7343 ( .A0(\D_cache/N170 ), .A1(n3995), .B0(n3997), .B1(n10341), 
        .C0(mem_rdata_D[110]), .C1(n3985), .Y(\D_cache/n489 ) );
  OA22X2 U7344 ( .A0(n8889), .A1(n3968), .B0(n3954), .B1(\D_cache/n491 ), .Y(
        \D_cache/n490 ) );
  AOI222XL U7345 ( .A0(\D_cache/N171 ), .A1(n3995), .B0(n3997), .B1(n10342), 
        .C0(mem_rdata_D[109]), .C1(n3985), .Y(\D_cache/n491 ) );
  OA22X2 U7346 ( .A0(n8890), .A1(n3968), .B0(n3954), .B1(\D_cache/n493 ), .Y(
        \D_cache/n492 ) );
  AOI222XL U7347 ( .A0(\D_cache/N172 ), .A1(n3995), .B0(n3996), .B1(n10343), 
        .C0(mem_rdata_D[108]), .C1(n3985), .Y(\D_cache/n493 ) );
  OA22X2 U7348 ( .A0(n8891), .A1(n3968), .B0(n3954), .B1(\D_cache/n495 ), .Y(
        \D_cache/n494 ) );
  AOI222XL U7349 ( .A0(\D_cache/N173 ), .A1(n3995), .B0(n3996), .B1(n10344), 
        .C0(mem_rdata_D[107]), .C1(n3985), .Y(\D_cache/n495 ) );
  OA22X2 U7350 ( .A0(n8892), .A1(n3968), .B0(n3954), .B1(\D_cache/n497 ), .Y(
        \D_cache/n496 ) );
  AOI222XL U7351 ( .A0(\D_cache/N174 ), .A1(n3995), .B0(n3996), .B1(n10345), 
        .C0(mem_rdata_D[106]), .C1(n3985), .Y(\D_cache/n497 ) );
  OA22X2 U7352 ( .A0(n8893), .A1(n3968), .B0(n3954), .B1(\D_cache/n499 ), .Y(
        \D_cache/n498 ) );
  AOI222XL U7353 ( .A0(\D_cache/N175 ), .A1(\D_cache/n454 ), .B0(n3996), .B1(
        n10346), .C0(mem_rdata_D[105]), .C1(n3985), .Y(\D_cache/n499 ) );
  OA22X2 U7354 ( .A0(n8894), .A1(n3969), .B0(n3954), .B1(\D_cache/n501 ), .Y(
        \D_cache/n500 ) );
  AOI222XL U7355 ( .A0(\D_cache/N176 ), .A1(\D_cache/n454 ), .B0(n3996), .B1(
        n10347), .C0(mem_rdata_D[104]), .C1(n3985), .Y(\D_cache/n501 ) );
  OA22X2 U7356 ( .A0(n8895), .A1(n3969), .B0(n3954), .B1(\D_cache/n503 ), .Y(
        \D_cache/n502 ) );
  AOI222XL U7357 ( .A0(\D_cache/N177 ), .A1(\D_cache/n454 ), .B0(n3996), .B1(
        n10348), .C0(mem_rdata_D[103]), .C1(n3985), .Y(\D_cache/n503 ) );
  OA22X2 U7358 ( .A0(n8896), .A1(n3969), .B0(n3954), .B1(\D_cache/n505 ), .Y(
        \D_cache/n504 ) );
  AOI222XL U7359 ( .A0(\D_cache/N178 ), .A1(\D_cache/n454 ), .B0(n3996), .B1(
        n10349), .C0(mem_rdata_D[102]), .C1(n3985), .Y(\D_cache/n505 ) );
  OA22X2 U7360 ( .A0(n8897), .A1(n3969), .B0(n3954), .B1(\D_cache/n507 ), .Y(
        \D_cache/n506 ) );
  AOI222XL U7361 ( .A0(\D_cache/N179 ), .A1(\D_cache/n454 ), .B0(n3996), .B1(
        n10350), .C0(mem_rdata_D[101]), .C1(n3982), .Y(\D_cache/n507 ) );
  OA22X2 U7362 ( .A0(n8898), .A1(n3969), .B0(n3954), .B1(\D_cache/n509 ), .Y(
        \D_cache/n508 ) );
  AOI222XL U7363 ( .A0(\D_cache/N180 ), .A1(\D_cache/n454 ), .B0(n3996), .B1(
        n10351), .C0(mem_rdata_D[100]), .C1(n3983), .Y(\D_cache/n509 ) );
  OA22X2 U7364 ( .A0(n8899), .A1(n3969), .B0(n3954), .B1(\D_cache/n511 ), .Y(
        \D_cache/n510 ) );
  AOI222XL U7365 ( .A0(\D_cache/N181 ), .A1(\D_cache/n454 ), .B0(n3996), .B1(
        n10352), .C0(mem_rdata_D[99]), .C1(n3985), .Y(\D_cache/n511 ) );
  OA22X2 U7366 ( .A0(n8900), .A1(n3968), .B0(n3954), .B1(\D_cache/n513 ), .Y(
        \D_cache/n512 ) );
  AOI222XL U7367 ( .A0(\D_cache/N182 ), .A1(\D_cache/n454 ), .B0(n3996), .B1(
        n10353), .C0(mem_rdata_D[98]), .C1(n3982), .Y(\D_cache/n513 ) );
  OA22X2 U7368 ( .A0(n8901), .A1(n3969), .B0(n3954), .B1(\D_cache/n515 ), .Y(
        \D_cache/n514 ) );
  AOI222XL U7369 ( .A0(\D_cache/N183 ), .A1(\D_cache/n454 ), .B0(n3996), .B1(
        n10354), .C0(mem_rdata_D[97]), .C1(n3983), .Y(\D_cache/n515 ) );
  OA22X2 U7370 ( .A0(n8902), .A1(n3966), .B0(n3950), .B1(\D_cache/n517 ), .Y(
        \D_cache/n516 ) );
  AOI222XL U7371 ( .A0(\D_cache/N184 ), .A1(\D_cache/n454 ), .B0(n3996), .B1(
        n10355), .C0(mem_rdata_D[96]), .C1(n3985), .Y(\D_cache/n517 ) );
  OA22X2 U7372 ( .A0(n8746), .A1(n3959), .B0(n3952), .B1(\D_cache/n249 ), .Y(
        \D_cache/n248 ) );
  AOI222XL U7373 ( .A0(\D_cache/N57 ), .A1(\D_cache/n250 ), .B0(n10324), .B1(
        n3987), .C0(mem_rdata_D[31]), .C1(n3979), .Y(\D_cache/n249 ) );
  OA22X2 U7374 ( .A0(n8747), .A1(n3958), .B0(n3952), .B1(\D_cache/n253 ), .Y(
        \D_cache/n252 ) );
  AOI222XL U7375 ( .A0(\D_cache/N58 ), .A1(n3986), .B0(n10325), .B1(n3988), 
        .C0(mem_rdata_D[30]), .C1(n3979), .Y(\D_cache/n253 ) );
  OA22X2 U7376 ( .A0(n8748), .A1(n3960), .B0(n3952), .B1(\D_cache/n255 ), .Y(
        \D_cache/n254 ) );
  AOI222XL U7377 ( .A0(\D_cache/N59 ), .A1(n3986), .B0(n10326), .B1(
        \D_cache/n251 ), .C0(mem_rdata_D[29]), .C1(n3979), .Y(\D_cache/n255 )
         );
  OA22X2 U7378 ( .A0(n8749), .A1(n3956), .B0(n3952), .B1(\D_cache/n257 ), .Y(
        \D_cache/n256 ) );
  AOI222XL U7379 ( .A0(\D_cache/N60 ), .A1(\D_cache/n250 ), .B0(n10327), .B1(
        n3987), .C0(mem_rdata_D[28]), .C1(n3979), .Y(\D_cache/n257 ) );
  OA22X2 U7380 ( .A0(n8750), .A1(n3959), .B0(n3951), .B1(\D_cache/n259 ), .Y(
        \D_cache/n258 ) );
  AOI222XL U7381 ( .A0(\D_cache/N61 ), .A1(n3986), .B0(n10328), .B1(n3988), 
        .C0(mem_rdata_D[27]), .C1(n3979), .Y(\D_cache/n259 ) );
  OA22X2 U7382 ( .A0(n8751), .A1(n3958), .B0(n3951), .B1(\D_cache/n261 ), .Y(
        \D_cache/n260 ) );
  AOI222XL U7383 ( .A0(\D_cache/N62 ), .A1(n3986), .B0(n10329), .B1(n3987), 
        .C0(mem_rdata_D[26]), .C1(n3979), .Y(\D_cache/n261 ) );
  OA22X2 U7384 ( .A0(n8752), .A1(n3967), .B0(n3951), .B1(\D_cache/n263 ), .Y(
        \D_cache/n262 ) );
  AOI222XL U7385 ( .A0(\D_cache/N63 ), .A1(n3986), .B0(n10330), .B1(n3988), 
        .C0(mem_rdata_D[25]), .C1(n3979), .Y(\D_cache/n263 ) );
  OA22X2 U7386 ( .A0(n8753), .A1(n3963), .B0(n3951), .B1(\D_cache/n265 ), .Y(
        \D_cache/n264 ) );
  AOI222XL U7387 ( .A0(\D_cache/N64 ), .A1(n3986), .B0(n10331), .B1(n3987), 
        .C0(mem_rdata_D[24]), .C1(n3979), .Y(\D_cache/n265 ) );
  OA22X2 U7388 ( .A0(n8754), .A1(n3957), .B0(n3951), .B1(\D_cache/n267 ), .Y(
        \D_cache/n266 ) );
  AOI222XL U7389 ( .A0(\D_cache/N65 ), .A1(n3986), .B0(n10332), .B1(n3988), 
        .C0(mem_rdata_D[23]), .C1(n3979), .Y(\D_cache/n267 ) );
  OA22X2 U7390 ( .A0(n8755), .A1(n3958), .B0(n3951), .B1(\D_cache/n269 ), .Y(
        \D_cache/n268 ) );
  AOI222XL U7391 ( .A0(\D_cache/N66 ), .A1(n3986), .B0(n10333), .B1(n3988), 
        .C0(mem_rdata_D[22]), .C1(n3979), .Y(\D_cache/n269 ) );
  OA22X2 U7392 ( .A0(n8756), .A1(n3958), .B0(n3951), .B1(\D_cache/n271 ), .Y(
        \D_cache/n270 ) );
  AOI222XL U7393 ( .A0(\D_cache/N67 ), .A1(n3986), .B0(n10334), .B1(n3988), 
        .C0(mem_rdata_D[21]), .C1(n3979), .Y(\D_cache/n271 ) );
  OA22X2 U7394 ( .A0(n8757), .A1(n3958), .B0(n3951), .B1(\D_cache/n273 ), .Y(
        \D_cache/n272 ) );
  AOI222XL U7395 ( .A0(\D_cache/N68 ), .A1(n3986), .B0(n10335), .B1(n3988), 
        .C0(mem_rdata_D[20]), .C1(n3979), .Y(\D_cache/n273 ) );
  OA22X2 U7396 ( .A0(n8758), .A1(n3958), .B0(n3951), .B1(\D_cache/n275 ), .Y(
        \D_cache/n274 ) );
  AOI222XL U7397 ( .A0(\D_cache/N69 ), .A1(n3986), .B0(n10336), .B1(n3988), 
        .C0(mem_rdata_D[19]), .C1(n3979), .Y(\D_cache/n275 ) );
  OA22X2 U7398 ( .A0(n8833), .A1(n3958), .B0(n3951), .B1(\D_cache/n277 ), .Y(
        \D_cache/n276 ) );
  AOI222XL U7399 ( .A0(\D_cache/N70 ), .A1(n3986), .B0(n10337), .B1(n3988), 
        .C0(mem_rdata_D[18]), .C1(n3979), .Y(\D_cache/n277 ) );
  OA22X2 U7400 ( .A0(n8834), .A1(n3958), .B0(n3951), .B1(\D_cache/n279 ), .Y(
        \D_cache/n278 ) );
  AOI222XL U7401 ( .A0(\D_cache/N71 ), .A1(n3986), .B0(n10338), .B1(n3988), 
        .C0(mem_rdata_D[17]), .C1(n3980), .Y(\D_cache/n279 ) );
  OA22X2 U7402 ( .A0(n8835), .A1(n3959), .B0(n3951), .B1(\D_cache/n281 ), .Y(
        \D_cache/n280 ) );
  AOI222XL U7403 ( .A0(\D_cache/N72 ), .A1(n3986), .B0(n10339), .B1(n3988), 
        .C0(mem_rdata_D[16]), .C1(n3980), .Y(\D_cache/n281 ) );
  OA22X2 U7404 ( .A0(n8836), .A1(n3959), .B0(n3951), .B1(\D_cache/n283 ), .Y(
        \D_cache/n282 ) );
  AOI222XL U7405 ( .A0(\D_cache/N73 ), .A1(n3986), .B0(n10340), .B1(n3988), 
        .C0(mem_rdata_D[15]), .C1(n3980), .Y(\D_cache/n283 ) );
  OA22X2 U7406 ( .A0(n8837), .A1(n3959), .B0(n3951), .B1(\D_cache/n285 ), .Y(
        \D_cache/n284 ) );
  AOI222XL U7407 ( .A0(\D_cache/N74 ), .A1(n3986), .B0(n10341), .B1(n3988), 
        .C0(mem_rdata_D[14]), .C1(n3980), .Y(\D_cache/n285 ) );
  OA22X2 U7408 ( .A0(n8838), .A1(n3959), .B0(n3951), .B1(\D_cache/n287 ), .Y(
        \D_cache/n286 ) );
  AOI222XL U7409 ( .A0(\D_cache/N75 ), .A1(n3986), .B0(n10342), .B1(n3988), 
        .C0(mem_rdata_D[13]), .C1(n3980), .Y(\D_cache/n287 ) );
  OA22X2 U7410 ( .A0(n8839), .A1(n3959), .B0(n3951), .B1(\D_cache/n289 ), .Y(
        \D_cache/n288 ) );
  AOI222XL U7411 ( .A0(\D_cache/N76 ), .A1(n3986), .B0(n10343), .B1(n3988), 
        .C0(mem_rdata_D[12]), .C1(n3980), .Y(\D_cache/n289 ) );
  OA22X2 U7412 ( .A0(n8840), .A1(n3959), .B0(n3951), .B1(\D_cache/n291 ), .Y(
        \D_cache/n290 ) );
  AOI222XL U7413 ( .A0(\D_cache/N77 ), .A1(n3986), .B0(n10344), .B1(n3987), 
        .C0(mem_rdata_D[11]), .C1(n3980), .Y(\D_cache/n291 ) );
  OA22X2 U7414 ( .A0(n8841), .A1(n3960), .B0(n3951), .B1(\D_cache/n293 ), .Y(
        \D_cache/n292 ) );
  AOI222XL U7415 ( .A0(\D_cache/N78 ), .A1(n3986), .B0(n10345), .B1(n3987), 
        .C0(mem_rdata_D[10]), .C1(n3980), .Y(\D_cache/n293 ) );
  OA22X2 U7416 ( .A0(n8842), .A1(n3960), .B0(n3950), .B1(\D_cache/n295 ), .Y(
        \D_cache/n294 ) );
  AOI222XL U7417 ( .A0(\D_cache/N79 ), .A1(\D_cache/n250 ), .B0(n10346), .B1(
        n3987), .C0(mem_rdata_D[9]), .C1(n3980), .Y(\D_cache/n295 ) );
  OA22X2 U7418 ( .A0(n8843), .A1(n3960), .B0(n3950), .B1(\D_cache/n297 ), .Y(
        \D_cache/n296 ) );
  AOI222XL U7419 ( .A0(\D_cache/N80 ), .A1(\D_cache/n250 ), .B0(n10347), .B1(
        n3987), .C0(mem_rdata_D[8]), .C1(n3980), .Y(\D_cache/n297 ) );
  OA22X2 U7420 ( .A0(n8844), .A1(n3960), .B0(n3950), .B1(\D_cache/n299 ), .Y(
        \D_cache/n298 ) );
  AOI222XL U7421 ( .A0(\D_cache/N81 ), .A1(\D_cache/n250 ), .B0(n10348), .B1(
        n3987), .C0(mem_rdata_D[7]), .C1(n3980), .Y(\D_cache/n299 ) );
  OA22X2 U7422 ( .A0(n8845), .A1(n3963), .B0(n3950), .B1(\D_cache/n301 ), .Y(
        \D_cache/n300 ) );
  AOI222XL U7423 ( .A0(\D_cache/N82 ), .A1(\D_cache/n250 ), .B0(n10349), .B1(
        n3987), .C0(mem_rdata_D[6]), .C1(n3980), .Y(\D_cache/n301 ) );
  OA22X2 U7424 ( .A0(n8846), .A1(n3960), .B0(n3950), .B1(\D_cache/n303 ), .Y(
        \D_cache/n302 ) );
  AOI222XL U7425 ( .A0(\D_cache/N83 ), .A1(\D_cache/n250 ), .B0(n10350), .B1(
        n3987), .C0(mem_rdata_D[5]), .C1(n3980), .Y(\D_cache/n303 ) );
  OA22X2 U7426 ( .A0(n8847), .A1(n3960), .B0(n3950), .B1(\D_cache/n305 ), .Y(
        \D_cache/n304 ) );
  AOI222XL U7427 ( .A0(\D_cache/N84 ), .A1(\D_cache/n250 ), .B0(n10351), .B1(
        n3987), .C0(mem_rdata_D[4]), .C1(n3980), .Y(\D_cache/n305 ) );
  OA22X2 U7428 ( .A0(n8848), .A1(n3967), .B0(n3950), .B1(\D_cache/n307 ), .Y(
        \D_cache/n306 ) );
  AOI222XL U7429 ( .A0(\D_cache/N85 ), .A1(\D_cache/n250 ), .B0(n10352), .B1(
        n3987), .C0(mem_rdata_D[3]), .C1(n3980), .Y(\D_cache/n307 ) );
  OA22X2 U7430 ( .A0(n8849), .A1(n3966), .B0(n3950), .B1(\D_cache/n309 ), .Y(
        \D_cache/n308 ) );
  AOI222XL U7431 ( .A0(\D_cache/N86 ), .A1(\D_cache/n250 ), .B0(n10353), .B1(
        n3987), .C0(mem_rdata_D[2]), .C1(n3979), .Y(\D_cache/n309 ) );
  OA22X2 U7432 ( .A0(n8850), .A1(n3966), .B0(n3950), .B1(\D_cache/n311 ), .Y(
        \D_cache/n310 ) );
  AOI222XL U7433 ( .A0(\D_cache/N87 ), .A1(\D_cache/n250 ), .B0(n10354), .B1(
        n3987), .C0(mem_rdata_D[1]), .C1(n3982), .Y(\D_cache/n311 ) );
  OA22X2 U7434 ( .A0(n8851), .A1(n3967), .B0(n3950), .B1(\D_cache/n313 ), .Y(
        \D_cache/n312 ) );
  AOI222XL U7435 ( .A0(\D_cache/N88 ), .A1(\D_cache/n250 ), .B0(n10355), .B1(
        n3987), .C0(mem_rdata_D[0]), .C1(n3984), .Y(\D_cache/n313 ) );
  NOR2BX1 U7436 ( .AN(n10322), .B(n10323), .Y(\D_cache/n201 ) );
  NOR2BX1 U7437 ( .AN(n10323), .B(n10322), .Y(\D_cache/n203 ) );
  AOI2BB2X1 U7438 ( .B0(\D_cache/N145 ), .B1(n2153), .A0N(n24), .A1N(n8895), 
        .Y(\D_cache/n170 ) );
  CLKINVX1 U7439 ( .A(n7081), .Y(n7078) );
  NOR2X1 U7440 ( .A(n10323), .B(n10322), .Y(\D_cache/n202 ) );
  XOR2X1 U7441 ( .A(n7994), .B(ICACHE_addr[15]), .Y(n7996) );
  XOR2X1 U7442 ( .A(n7963), .B(ICACHE_addr[13]), .Y(n7965) );
  XOR2X1 U7443 ( .A(n7928), .B(ICACHE_addr[11]), .Y(n7930) );
  XOR2X1 U7444 ( .A(n7929), .B(ICACHE_addr[12]), .Y(n7944) );
  NAND2X1 U7445 ( .A(\i_MIPS/ALUin1[21] ), .B(n4631), .Y(n8549) );
  NOR4X1 U7446 ( .A(n4768), .B(n4767), .C(n4766), .D(n4765), .Y(n4769) );
  AND2X2 U7447 ( .A(\i_MIPS/EX_MEM_0 ), .B(n4764), .Y(n4770) );
  NAND4X1 U7448 ( .A(n4808), .B(n4807), .C(n4806), .D(n4805), .Y(n7069) );
  XOR2X1 U7449 ( .A(\i_MIPS/n320 ), .B(\i_MIPS/Reg_W[4] ), .Y(n4807) );
  XOR2X1 U7450 ( .A(\i_MIPS/n318 ), .B(\i_MIPS/Reg_W[3] ), .Y(n4808) );
  NOR4X1 U7451 ( .A(\i_MIPS/forward_unit/n10 ), .B(n4804), .C(n4803), .D(n4802), .Y(n4805) );
  NAND2X1 U7452 ( .A(\i_MIPS/ALUin1[13] ), .B(n4653), .Y(n6389) );
  NAND2X1 U7453 ( .A(\i_MIPS/ALUin1[12] ), .B(n4652), .Y(n8480) );
  NAND2X1 U7454 ( .A(\i_MIPS/ALUin1[10] ), .B(n4691), .Y(n8466) );
  OAI2BB2XL U7455 ( .B0(n3666), .B1(n3780), .A0N(
        \i_MIPS/Register/register[0][6] ), .A1N(n3782), .Y(
        \i_MIPS/Register/n1114 ) );
  OAI2BB2XL U7456 ( .B0(n3666), .B1(n3777), .A0N(
        \i_MIPS/Register/register[1][6] ), .A1N(n3779), .Y(
        \i_MIPS/Register/n1082 ) );
  OAI2BB2XL U7457 ( .B0(n3666), .B1(n3774), .A0N(
        \i_MIPS/Register/register[2][6] ), .A1N(n3776), .Y(
        \i_MIPS/Register/n1050 ) );
  OAI2BB2XL U7458 ( .B0(n3666), .B1(n3771), .A0N(
        \i_MIPS/Register/register[3][6] ), .A1N(n3773), .Y(
        \i_MIPS/Register/n1018 ) );
  OAI2BB2XL U7459 ( .B0(n3666), .B1(n3768), .A0N(
        \i_MIPS/Register/register[4][6] ), .A1N(n3770), .Y(
        \i_MIPS/Register/n986 ) );
  OAI2BB2XL U7460 ( .B0(n3666), .B1(n3765), .A0N(
        \i_MIPS/Register/register[5][6] ), .A1N(n3767), .Y(
        \i_MIPS/Register/n954 ) );
  OAI2BB2XL U7461 ( .B0(n3666), .B1(n3762), .A0N(
        \i_MIPS/Register/register[6][6] ), .A1N(n3764), .Y(
        \i_MIPS/Register/n922 ) );
  OAI2BB2XL U7462 ( .B0(n3666), .B1(n3726), .A0N(
        \i_MIPS/Register/register[18][6] ), .A1N(n3728), .Y(
        \i_MIPS/Register/n538 ) );
  OAI2BB2XL U7463 ( .B0(n3666), .B1(n3723), .A0N(
        \i_MIPS/Register/register[19][6] ), .A1N(n3725), .Y(
        \i_MIPS/Register/n506 ) );
  OAI2BB2XL U7464 ( .B0(n3666), .B1(n3720), .A0N(
        \i_MIPS/Register/register[20][6] ), .A1N(n3722), .Y(
        \i_MIPS/Register/n474 ) );
  OAI2BB2XL U7465 ( .B0(n3666), .B1(n3717), .A0N(
        \i_MIPS/Register/register[21][6] ), .A1N(n3719), .Y(
        \i_MIPS/Register/n442 ) );
  OAI2BB2XL U7466 ( .B0(n3666), .B1(n3714), .A0N(
        \i_MIPS/Register/register[22][6] ), .A1N(n3716), .Y(
        \i_MIPS/Register/n410 ) );
  OAI2BB2XL U7467 ( .B0(n3666), .B1(n3711), .A0N(
        \i_MIPS/Register/register[23][6] ), .A1N(n3713), .Y(
        \i_MIPS/Register/n378 ) );
  OAI2BB2XL U7468 ( .B0(n3666), .B1(n3708), .A0N(
        \i_MIPS/Register/register[24][6] ), .A1N(n3710), .Y(
        \i_MIPS/Register/n346 ) );
  OAI2BB2XL U7469 ( .B0(n3666), .B1(n3705), .A0N(
        \i_MIPS/Register/register[25][6] ), .A1N(n3707), .Y(
        \i_MIPS/Register/n314 ) );
  OAI2BB2XL U7470 ( .B0(n3666), .B1(n3702), .A0N(
        \i_MIPS/Register/register[26][6] ), .A1N(n3704), .Y(
        \i_MIPS/Register/n282 ) );
  OAI2BB2XL U7471 ( .B0(n3666), .B1(n3699), .A0N(
        \i_MIPS/Register/register[27][6] ), .A1N(n3701), .Y(
        \i_MIPS/Register/n250 ) );
  OAI2BB2XL U7472 ( .B0(n3666), .B1(n3696), .A0N(
        \i_MIPS/Register/register[28][6] ), .A1N(n3698), .Y(
        \i_MIPS/Register/n218 ) );
  OAI2BB2XL U7473 ( .B0(n3666), .B1(n3693), .A0N(
        \i_MIPS/Register/register[29][6] ), .A1N(n3695), .Y(
        \i_MIPS/Register/n186 ) );
  NAND2X1 U7474 ( .A(\i_MIPS/ALUin1[20] ), .B(n4642), .Y(n8465) );
  NAND2X1 U7475 ( .A(\i_MIPS/ALUin1[29] ), .B(n4623), .Y(n8533) );
  NAND2X1 U7476 ( .A(\i_MIPS/ALUin1[25] ), .B(n4628), .Y(n8524) );
  NAND2X1 U7477 ( .A(\i_MIPS/ALUin1[23] ), .B(n4636), .Y(n8545) );
  NAND2X1 U7478 ( .A(\i_MIPS/ALUin1[12] ), .B(n4662), .Y(n6390) );
  NAND2X1 U7479 ( .A(\i_MIPS/ALUin1[27] ), .B(n4625), .Y(n8520) );
  NAND2X1 U7480 ( .A(\i_MIPS/ALUin1[20] ), .B(n4639), .Y(n6468) );
  OAI2BB2XL U7481 ( .B0(n3639), .B1(n3781), .A0N(
        \i_MIPS/Register/register[0][30] ), .A1N(n3780), .Y(
        \i_MIPS/Register/n1138 ) );
  OAI2BB2XL U7482 ( .B0(n3644), .B1(n3780), .A0N(
        \i_MIPS/Register/register[0][27] ), .A1N(n3782), .Y(
        \i_MIPS/Register/n1135 ) );
  OAI2BB2XL U7483 ( .B0(n3675), .B1(n3781), .A0N(
        \i_MIPS/Register/register[0][25] ), .A1N(n3782), .Y(
        \i_MIPS/Register/n1133 ) );
  OAI2BB2XL U7484 ( .B0(n3684), .B1(n3781), .A0N(
        \i_MIPS/Register/register[0][21] ), .A1N(n3781), .Y(
        \i_MIPS/Register/n1129 ) );
  OAI2BB2XL U7485 ( .B0(n3635), .B1(n3781), .A0N(
        \i_MIPS/Register/register[0][19] ), .A1N(n3782), .Y(
        \i_MIPS/Register/n1127 ) );
  OAI2BB2XL U7486 ( .B0(n3641), .B1(n3778), .A0N(
        \i_MIPS/Register/register[1][29] ), .A1N(n3779), .Y(
        \i_MIPS/Register/n1105 ) );
  OAI2BB2XL U7487 ( .B0(n3639), .B1(n3775), .A0N(
        \i_MIPS/Register/register[2][30] ), .A1N(n3774), .Y(
        \i_MIPS/Register/n1074 ) );
  OAI2BB2XL U7488 ( .B0(n3644), .B1(n3774), .A0N(
        \i_MIPS/Register/register[2][27] ), .A1N(n3776), .Y(
        \i_MIPS/Register/n1071 ) );
  OAI2BB2XL U7489 ( .B0(n3675), .B1(n3775), .A0N(
        \i_MIPS/Register/register[2][25] ), .A1N(n3776), .Y(
        \i_MIPS/Register/n1069 ) );
  OAI2BB2XL U7490 ( .B0(n3684), .B1(n3775), .A0N(
        \i_MIPS/Register/register[2][21] ), .A1N(n3775), .Y(
        \i_MIPS/Register/n1065 ) );
  OAI2BB2XL U7491 ( .B0(n3635), .B1(n3775), .A0N(
        \i_MIPS/Register/register[2][19] ), .A1N(n3776), .Y(
        \i_MIPS/Register/n1063 ) );
  OAI2BB2XL U7492 ( .B0(n3641), .B1(n3772), .A0N(
        \i_MIPS/Register/register[3][29] ), .A1N(n3773), .Y(
        \i_MIPS/Register/n1041 ) );
  OAI2BB2XL U7493 ( .B0(n3639), .B1(n3769), .A0N(
        \i_MIPS/Register/register[4][30] ), .A1N(n3769), .Y(
        \i_MIPS/Register/n1010 ) );
  OAI2BB2XL U7494 ( .B0(n3644), .B1(n3768), .A0N(
        \i_MIPS/Register/register[4][27] ), .A1N(n3770), .Y(
        \i_MIPS/Register/n1007 ) );
  OAI2BB2XL U7495 ( .B0(n3675), .B1(n3769), .A0N(
        \i_MIPS/Register/register[4][25] ), .A1N(n3770), .Y(
        \i_MIPS/Register/n1005 ) );
  OAI2BB2XL U7496 ( .B0(n3684), .B1(n3769), .A0N(
        \i_MIPS/Register/register[4][21] ), .A1N(n3769), .Y(
        \i_MIPS/Register/n1001 ) );
  OAI2BB2XL U7497 ( .B0(n3635), .B1(n3769), .A0N(
        \i_MIPS/Register/register[4][19] ), .A1N(n3770), .Y(
        \i_MIPS/Register/n999 ) );
  OAI2BB2XL U7498 ( .B0(n3641), .B1(n3766), .A0N(
        \i_MIPS/Register/register[5][29] ), .A1N(n3767), .Y(
        \i_MIPS/Register/n977 ) );
  OAI2BB2XL U7499 ( .B0(n3639), .B1(n3763), .A0N(
        \i_MIPS/Register/register[6][30] ), .A1N(n3762), .Y(
        \i_MIPS/Register/n946 ) );
  OAI2BB2XL U7500 ( .B0(n3644), .B1(n3762), .A0N(
        \i_MIPS/Register/register[6][27] ), .A1N(n3764), .Y(
        \i_MIPS/Register/n943 ) );
  OAI2BB2XL U7501 ( .B0(n3675), .B1(n3763), .A0N(
        \i_MIPS/Register/register[6][25] ), .A1N(n3764), .Y(
        \i_MIPS/Register/n941 ) );
  OAI2BB2XL U7502 ( .B0(n3684), .B1(n3763), .A0N(
        \i_MIPS/Register/register[6][21] ), .A1N(n3763), .Y(
        \i_MIPS/Register/n937 ) );
  OAI2BB2XL U7503 ( .B0(n3635), .B1(n3763), .A0N(
        \i_MIPS/Register/register[6][19] ), .A1N(n3764), .Y(
        \i_MIPS/Register/n935 ) );
  OAI2BB2XL U7504 ( .B0(n3639), .B1(n3760), .A0N(
        \i_MIPS/Register/register[7][30] ), .A1N(n3759), .Y(
        \i_MIPS/Register/n914 ) );
  OAI2BB2XL U7505 ( .B0(n3641), .B1(n44), .A0N(
        \i_MIPS/Register/register[7][29] ), .A1N(n3761), .Y(
        \i_MIPS/Register/n913 ) );
  OAI2BB2XL U7506 ( .B0(n3644), .B1(n44), .A0N(
        \i_MIPS/Register/register[7][27] ), .A1N(n3761), .Y(
        \i_MIPS/Register/n911 ) );
  OAI2BB2XL U7507 ( .B0(n3675), .B1(n44), .A0N(
        \i_MIPS/Register/register[7][25] ), .A1N(n3761), .Y(
        \i_MIPS/Register/n909 ) );
  OAI2BB2XL U7508 ( .B0(n3684), .B1(n3760), .A0N(
        \i_MIPS/Register/register[7][21] ), .A1N(n3761), .Y(
        \i_MIPS/Register/n905 ) );
  OAI2BB2XL U7509 ( .B0(n3635), .B1(n3760), .A0N(
        \i_MIPS/Register/register[7][19] ), .A1N(n3759), .Y(
        \i_MIPS/Register/n903 ) );
  OAI2BB2XL U7510 ( .B0(n3639), .B1(n3753), .A0N(
        \i_MIPS/Register/register[9][30] ), .A1N(n3753), .Y(
        \i_MIPS/Register/n850 ) );
  OAI2BB2XL U7511 ( .B0(n3641), .B1(n3754), .A0N(
        \i_MIPS/Register/register[9][29] ), .A1N(n3755), .Y(
        \i_MIPS/Register/n849 ) );
  OAI2BB2XL U7512 ( .B0(n3644), .B1(n3753), .A0N(
        \i_MIPS/Register/register[9][27] ), .A1N(n3755), .Y(
        \i_MIPS/Register/n847 ) );
  OAI2BB2XL U7513 ( .B0(n3675), .B1(n42), .A0N(
        \i_MIPS/Register/register[9][25] ), .A1N(n3755), .Y(
        \i_MIPS/Register/n845 ) );
  OAI2BB2XL U7514 ( .B0(n3684), .B1(n3754), .A0N(
        \i_MIPS/Register/register[9][21] ), .A1N(n3753), .Y(
        \i_MIPS/Register/n841 ) );
  OAI2BB2XL U7515 ( .B0(n3635), .B1(n3754), .A0N(
        \i_MIPS/Register/register[9][19] ), .A1N(n3755), .Y(
        \i_MIPS/Register/n839 ) );
  OAI2BB2XL U7516 ( .B0(n3639), .B1(n3747), .A0N(
        \i_MIPS/Register/register[11][30] ), .A1N(n3747), .Y(
        \i_MIPS/Register/n786 ) );
  OAI2BB2XL U7517 ( .B0(n3641), .B1(n3748), .A0N(
        \i_MIPS/Register/register[11][29] ), .A1N(n3749), .Y(
        \i_MIPS/Register/n785 ) );
  OAI2BB2XL U7518 ( .B0(n3644), .B1(n3747), .A0N(
        \i_MIPS/Register/register[11][27] ), .A1N(n3749), .Y(
        \i_MIPS/Register/n783 ) );
  OAI2BB2XL U7519 ( .B0(n3675), .B1(n40), .A0N(
        \i_MIPS/Register/register[11][25] ), .A1N(n3749), .Y(
        \i_MIPS/Register/n781 ) );
  OAI2BB2XL U7520 ( .B0(n3684), .B1(n3748), .A0N(
        \i_MIPS/Register/register[11][21] ), .A1N(n3747), .Y(
        \i_MIPS/Register/n777 ) );
  OAI2BB2XL U7521 ( .B0(n3635), .B1(n3748), .A0N(
        \i_MIPS/Register/register[11][19] ), .A1N(n3749), .Y(
        \i_MIPS/Register/n775 ) );
  OAI2BB2XL U7522 ( .B0(n3641), .B1(n3744), .A0N(
        \i_MIPS/Register/register[12][29] ), .A1N(n3746), .Y(
        \i_MIPS/Register/n753 ) );
  OAI2BB2XL U7523 ( .B0(n3639), .B1(n3741), .A0N(
        \i_MIPS/Register/register[13][30] ), .A1N(n3741), .Y(
        \i_MIPS/Register/n722 ) );
  OAI2BB2XL U7524 ( .B0(n3644), .B1(n3742), .A0N(
        \i_MIPS/Register/register[13][27] ), .A1N(n3743), .Y(
        \i_MIPS/Register/n719 ) );
  OAI2BB2XL U7525 ( .B0(n3675), .B1(n3741), .A0N(
        \i_MIPS/Register/register[13][25] ), .A1N(n3743), .Y(
        \i_MIPS/Register/n717 ) );
  OAI2BB2XL U7526 ( .B0(n3684), .B1(n3742), .A0N(
        \i_MIPS/Register/register[13][21] ), .A1N(n3741), .Y(
        \i_MIPS/Register/n713 ) );
  OAI2BB2XL U7527 ( .B0(n3635), .B1(n3742), .A0N(
        \i_MIPS/Register/register[13][19] ), .A1N(n3743), .Y(
        \i_MIPS/Register/n711 ) );
  OAI2BB2XL U7528 ( .B0(n3639), .B1(n3738), .A0N(
        \i_MIPS/Register/register[14][30] ), .A1N(n3739), .Y(
        \i_MIPS/Register/n690 ) );
  OAI2BB2XL U7529 ( .B0(n3644), .B1(n3739), .A0N(
        \i_MIPS/Register/register[14][27] ), .A1N(n3740), .Y(
        \i_MIPS/Register/n687 ) );
  OAI2BB2XL U7530 ( .B0(n3675), .B1(n3738), .A0N(
        \i_MIPS/Register/register[14][25] ), .A1N(n3740), .Y(
        \i_MIPS/Register/n685 ) );
  OAI2BB2XL U7531 ( .B0(n3684), .B1(n3739), .A0N(
        \i_MIPS/Register/register[14][21] ), .A1N(n3738), .Y(
        \i_MIPS/Register/n681 ) );
  OAI2BB2XL U7532 ( .B0(n3635), .B1(n3739), .A0N(
        \i_MIPS/Register/register[14][19] ), .A1N(n3740), .Y(
        \i_MIPS/Register/n679 ) );
  OAI2BB2XL U7533 ( .B0(n3641), .B1(n3735), .A0N(
        \i_MIPS/Register/register[15][29] ), .A1N(n3737), .Y(
        \i_MIPS/Register/n657 ) );
  OAI2BB2XL U7534 ( .B0(n3639), .B1(n3733), .A0N(
        \i_MIPS/Register/register[16][30] ), .A1N(n3733), .Y(
        \i_MIPS/Register/n626 ) );
  OAI2BB2XL U7535 ( .B0(n3644), .B1(n3732), .A0N(
        \i_MIPS/Register/register[16][27] ), .A1N(n3734), .Y(
        \i_MIPS/Register/n623 ) );
  OAI2BB2XL U7536 ( .B0(n3675), .B1(n3733), .A0N(
        \i_MIPS/Register/register[16][25] ), .A1N(n3734), .Y(
        \i_MIPS/Register/n621 ) );
  OAI2BB2XL U7537 ( .B0(n3684), .B1(n3733), .A0N(
        \i_MIPS/Register/register[16][21] ), .A1N(n3733), .Y(
        \i_MIPS/Register/n617 ) );
  OAI2BB2XL U7538 ( .B0(n3635), .B1(n3733), .A0N(
        \i_MIPS/Register/register[16][19] ), .A1N(n3734), .Y(
        \i_MIPS/Register/n615 ) );
  OAI2BB2XL U7539 ( .B0(n3641), .B1(n3730), .A0N(
        \i_MIPS/Register/register[17][29] ), .A1N(n3731), .Y(
        \i_MIPS/Register/n593 ) );
  OAI2BB2XL U7540 ( .B0(n3639), .B1(n3727), .A0N(
        \i_MIPS/Register/register[18][30] ), .A1N(n3727), .Y(
        \i_MIPS/Register/n562 ) );
  OAI2BB2XL U7541 ( .B0(n3641), .B1(n33), .A0N(
        \i_MIPS/Register/register[18][29] ), .A1N(n3728), .Y(
        \i_MIPS/Register/n561 ) );
  OAI2BB2XL U7542 ( .B0(n3644), .B1(n33), .A0N(
        \i_MIPS/Register/register[18][27] ), .A1N(n3728), .Y(
        \i_MIPS/Register/n559 ) );
  OAI2BB2XL U7543 ( .B0(n3675), .B1(n33), .A0N(
        \i_MIPS/Register/register[18][25] ), .A1N(n3728), .Y(
        \i_MIPS/Register/n557 ) );
  OAI2BB2XL U7544 ( .B0(n3684), .B1(n3727), .A0N(
        \i_MIPS/Register/register[18][21] ), .A1N(n3728), .Y(
        \i_MIPS/Register/n553 ) );
  OAI2BB2XL U7545 ( .B0(n3635), .B1(n3727), .A0N(
        \i_MIPS/Register/register[18][19] ), .A1N(n3726), .Y(
        \i_MIPS/Register/n551 ) );
  OAI2BB2XL U7546 ( .B0(n3639), .B1(n3721), .A0N(
        \i_MIPS/Register/register[20][30] ), .A1N(n3721), .Y(
        \i_MIPS/Register/n498 ) );
  OAI2BB2XL U7547 ( .B0(n3641), .B1(n31), .A0N(
        \i_MIPS/Register/register[20][29] ), .A1N(n3722), .Y(
        \i_MIPS/Register/n497 ) );
  OAI2BB2XL U7548 ( .B0(n3644), .B1(n31), .A0N(
        \i_MIPS/Register/register[20][27] ), .A1N(n3722), .Y(
        \i_MIPS/Register/n495 ) );
  OAI2BB2XL U7549 ( .B0(n3675), .B1(n31), .A0N(
        \i_MIPS/Register/register[20][25] ), .A1N(n3722), .Y(
        \i_MIPS/Register/n493 ) );
  OAI2BB2XL U7550 ( .B0(n3684), .B1(n3721), .A0N(
        \i_MIPS/Register/register[20][21] ), .A1N(n3722), .Y(
        \i_MIPS/Register/n489 ) );
  OAI2BB2XL U7551 ( .B0(n3635), .B1(n3721), .A0N(
        \i_MIPS/Register/register[20][19] ), .A1N(n3720), .Y(
        \i_MIPS/Register/n487 ) );
  OAI2BB2XL U7552 ( .B0(n3639), .B1(n3715), .A0N(
        \i_MIPS/Register/register[22][30] ), .A1N(n3715), .Y(
        \i_MIPS/Register/n434 ) );
  OAI2BB2XL U7553 ( .B0(n3641), .B1(n29), .A0N(
        \i_MIPS/Register/register[22][29] ), .A1N(n3716), .Y(
        \i_MIPS/Register/n433 ) );
  OAI2BB2XL U7554 ( .B0(n3644), .B1(n29), .A0N(
        \i_MIPS/Register/register[22][27] ), .A1N(n3716), .Y(
        \i_MIPS/Register/n431 ) );
  OAI2BB2XL U7555 ( .B0(n3675), .B1(n29), .A0N(
        \i_MIPS/Register/register[22][25] ), .A1N(n3716), .Y(
        \i_MIPS/Register/n429 ) );
  OAI2BB2XL U7556 ( .B0(n3684), .B1(n3715), .A0N(
        \i_MIPS/Register/register[22][21] ), .A1N(n3716), .Y(
        \i_MIPS/Register/n425 ) );
  OAI2BB2XL U7557 ( .B0(n3635), .B1(n3715), .A0N(
        \i_MIPS/Register/register[22][19] ), .A1N(n3714), .Y(
        \i_MIPS/Register/n423 ) );
  OAI2BB2XL U7558 ( .B0(n3639), .B1(n3709), .A0N(
        \i_MIPS/Register/register[24][30] ), .A1N(n3709), .Y(
        \i_MIPS/Register/n370 ) );
  OAI2BB2XL U7559 ( .B0(n3641), .B1(\i_MIPS/Register/n118 ), .A0N(
        \i_MIPS/Register/register[24][29] ), .A1N(n3710), .Y(
        \i_MIPS/Register/n369 ) );
  OAI2BB2XL U7560 ( .B0(n3644), .B1(\i_MIPS/Register/n118 ), .A0N(
        \i_MIPS/Register/register[24][27] ), .A1N(n3710), .Y(
        \i_MIPS/Register/n367 ) );
  OAI2BB2XL U7561 ( .B0(n3675), .B1(\i_MIPS/Register/n118 ), .A0N(
        \i_MIPS/Register/register[24][25] ), .A1N(n3710), .Y(
        \i_MIPS/Register/n365 ) );
  OAI2BB2XL U7562 ( .B0(n3684), .B1(n3709), .A0N(
        \i_MIPS/Register/register[24][21] ), .A1N(n3710), .Y(
        \i_MIPS/Register/n361 ) );
  OAI2BB2XL U7563 ( .B0(n3635), .B1(n3709), .A0N(
        \i_MIPS/Register/register[24][19] ), .A1N(n3708), .Y(
        \i_MIPS/Register/n359 ) );
  OAI2BB2XL U7564 ( .B0(n3639), .B1(n3703), .A0N(
        \i_MIPS/Register/register[26][30] ), .A1N(n3702), .Y(
        \i_MIPS/Register/n306 ) );
  OAI2BB2XL U7565 ( .B0(n3641), .B1(\i_MIPS/Register/n114 ), .A0N(
        \i_MIPS/Register/register[26][29] ), .A1N(n3704), .Y(
        \i_MIPS/Register/n305 ) );
  OAI2BB2XL U7566 ( .B0(n3644), .B1(\i_MIPS/Register/n114 ), .A0N(
        \i_MIPS/Register/register[26][27] ), .A1N(n3704), .Y(
        \i_MIPS/Register/n303 ) );
  OAI2BB2XL U7567 ( .B0(n3675), .B1(\i_MIPS/Register/n114 ), .A0N(
        \i_MIPS/Register/register[26][25] ), .A1N(n3704), .Y(
        \i_MIPS/Register/n301 ) );
  OAI2BB2XL U7568 ( .B0(n3684), .B1(n3703), .A0N(
        \i_MIPS/Register/register[26][21] ), .A1N(n3704), .Y(
        \i_MIPS/Register/n297 ) );
  OAI2BB2XL U7569 ( .B0(n3635), .B1(n3703), .A0N(
        \i_MIPS/Register/register[26][19] ), .A1N(n3702), .Y(
        \i_MIPS/Register/n295 ) );
  OAI2BB2XL U7570 ( .B0(n3639), .B1(n3697), .A0N(
        \i_MIPS/Register/register[28][30] ), .A1N(n3697), .Y(
        \i_MIPS/Register/n242 ) );
  OAI2BB2XL U7571 ( .B0(n3641), .B1(\i_MIPS/Register/n110 ), .A0N(
        \i_MIPS/Register/register[28][29] ), .A1N(n3698), .Y(
        \i_MIPS/Register/n241 ) );
  OAI2BB2XL U7572 ( .B0(n3644), .B1(\i_MIPS/Register/n110 ), .A0N(
        \i_MIPS/Register/register[28][27] ), .A1N(n3698), .Y(
        \i_MIPS/Register/n239 ) );
  OAI2BB2XL U7573 ( .B0(n3675), .B1(\i_MIPS/Register/n110 ), .A0N(
        \i_MIPS/Register/register[28][25] ), .A1N(n3698), .Y(
        \i_MIPS/Register/n237 ) );
  OAI2BB2XL U7574 ( .B0(n3684), .B1(n3697), .A0N(
        \i_MIPS/Register/register[28][21] ), .A1N(n3698), .Y(
        \i_MIPS/Register/n233 ) );
  OAI2BB2XL U7575 ( .B0(n3635), .B1(n3697), .A0N(
        \i_MIPS/Register/register[28][19] ), .A1N(n3696), .Y(
        \i_MIPS/Register/n231 ) );
  OAI2BB2XL U7576 ( .B0(n3641), .B1(n3690), .A0N(
        \i_MIPS/Register/register[30][29] ), .A1N(n3692), .Y(
        \i_MIPS/Register/n177 ) );
  AOI222XL U7577 ( .A0(n4835), .A1(\i_MIPS/ALU/N303 ), .B0(n6680), .B1(n4719), 
        .C0(n4718), .C1(n6682), .Y(n4720) );
  OAI2BB2XL U7578 ( .B0(n3665), .B1(n3774), .A0N(
        \i_MIPS/Register/register[2][9] ), .A1N(n3776), .Y(
        \i_MIPS/Register/n1053 ) );
  OAI2BB2XL U7579 ( .B0(n3665), .B1(n3765), .A0N(
        \i_MIPS/Register/register[5][9] ), .A1N(n3767), .Y(
        \i_MIPS/Register/n957 ) );
  OAI2BB2XL U7580 ( .B0(n3665), .B1(n3759), .A0N(
        \i_MIPS/Register/register[7][9] ), .A1N(n3761), .Y(
        \i_MIPS/Register/n893 ) );
  OAI2BB2XL U7581 ( .B0(n3665), .B1(n3756), .A0N(
        \i_MIPS/Register/register[8][9] ), .A1N(n3758), .Y(
        \i_MIPS/Register/n861 ) );
  OAI2BB2XL U7582 ( .B0(n3665), .B1(n3753), .A0N(
        \i_MIPS/Register/register[9][9] ), .A1N(n3755), .Y(
        \i_MIPS/Register/n829 ) );
  OAI2BB2XL U7583 ( .B0(n3665), .B1(n3750), .A0N(
        \i_MIPS/Register/register[10][9] ), .A1N(n3752), .Y(
        \i_MIPS/Register/n797 ) );
  OAI2BB2XL U7584 ( .B0(n3665), .B1(n3747), .A0N(
        \i_MIPS/Register/register[11][9] ), .A1N(n3749), .Y(
        \i_MIPS/Register/n765 ) );
  OAI2BB2XL U7585 ( .B0(n3665), .B1(n3738), .A0N(
        \i_MIPS/Register/register[14][9] ), .A1N(n3740), .Y(
        \i_MIPS/Register/n669 ) );
  OAI2BB2XL U7586 ( .B0(n3665), .B1(n3729), .A0N(
        \i_MIPS/Register/register[17][9] ), .A1N(n3731), .Y(
        \i_MIPS/Register/n573 ) );
  OAI2BB2XL U7587 ( .B0(n3665), .B1(n3726), .A0N(
        \i_MIPS/Register/register[18][9] ), .A1N(n3728), .Y(
        \i_MIPS/Register/n541 ) );
  OAI2BB2XL U7588 ( .B0(n3665), .B1(n3723), .A0N(
        \i_MIPS/Register/register[19][9] ), .A1N(n3725), .Y(
        \i_MIPS/Register/n509 ) );
  OAI2BB2XL U7589 ( .B0(n3665), .B1(n3720), .A0N(
        \i_MIPS/Register/register[20][9] ), .A1N(n3722), .Y(
        \i_MIPS/Register/n477 ) );
  OAI2BB2XL U7590 ( .B0(n3665), .B1(n3717), .A0N(
        \i_MIPS/Register/register[21][9] ), .A1N(n3719), .Y(
        \i_MIPS/Register/n445 ) );
  OAI2BB2XL U7591 ( .B0(n3665), .B1(n3714), .A0N(
        \i_MIPS/Register/register[22][9] ), .A1N(n3716), .Y(
        \i_MIPS/Register/n413 ) );
  OAI2BB2XL U7592 ( .B0(n3665), .B1(n3711), .A0N(
        \i_MIPS/Register/register[23][9] ), .A1N(n3713), .Y(
        \i_MIPS/Register/n381 ) );
  OAI2BB2XL U7593 ( .B0(n3665), .B1(n3708), .A0N(
        \i_MIPS/Register/register[24][9] ), .A1N(n3710), .Y(
        \i_MIPS/Register/n349 ) );
  OAI2BB2XL U7594 ( .B0(n3665), .B1(n3705), .A0N(
        \i_MIPS/Register/register[25][9] ), .A1N(n3707), .Y(
        \i_MIPS/Register/n317 ) );
  OAI2BB2XL U7595 ( .B0(n3665), .B1(n3702), .A0N(
        \i_MIPS/Register/register[26][9] ), .A1N(n3704), .Y(
        \i_MIPS/Register/n285 ) );
  OAI2BB2XL U7596 ( .B0(n3665), .B1(n3699), .A0N(
        \i_MIPS/Register/register[27][9] ), .A1N(n3701), .Y(
        \i_MIPS/Register/n253 ) );
  OAI2BB2XL U7597 ( .B0(n3665), .B1(n3696), .A0N(
        \i_MIPS/Register/register[28][9] ), .A1N(n3698), .Y(
        \i_MIPS/Register/n221 ) );
  OAI2BB2XL U7598 ( .B0(n3665), .B1(n3693), .A0N(
        \i_MIPS/Register/register[29][9] ), .A1N(n3695), .Y(
        \i_MIPS/Register/n189 ) );
  OAI2BB2XL U7599 ( .B0(n3665), .B1(n3690), .A0N(
        \i_MIPS/Register/register[30][9] ), .A1N(n3692), .Y(
        \i_MIPS/Register/n157 ) );
  XOR2X1 U7600 ( .A(\i_MIPS/IR_ID[18] ), .B(\i_MIPS/EX_MEM_next[71] ), .Y(
        n4777) );
  XOR2X1 U7601 ( .A(n4015), .B(n2891), .Y(n4776) );
  NOR4X1 U7602 ( .A(n4739), .B(n4738), .C(\i_MIPS/forward_unit/n15 ), .D(
        \i_MIPS/n372 ), .Y(n4740) );
  XOR2X1 U7603 ( .A(n4013), .B(n2891), .Y(n4739) );
  XOR2X1 U7604 ( .A(\i_MIPS/IR_ID[24] ), .B(n2890), .Y(n4738) );
  OAI2BB2XL U7605 ( .B0(n3642), .B1(n51), .A0N(
        \i_MIPS/Register/register[0][29] ), .A1N(n3782), .Y(
        \i_MIPS/Register/n1137 ) );
  OAI2BB2XL U7606 ( .B0(n3640), .B1(n50), .A0N(
        \i_MIPS/Register/register[1][30] ), .A1N(n3778), .Y(
        \i_MIPS/Register/n1106 ) );
  OAI2BB2XL U7607 ( .B0(n3645), .B1(n3778), .A0N(
        \i_MIPS/Register/register[1][27] ), .A1N(n3779), .Y(
        \i_MIPS/Register/n1103 ) );
  OAI2BB2XL U7608 ( .B0(n3676), .B1(n50), .A0N(
        \i_MIPS/Register/register[1][25] ), .A1N(n3779), .Y(
        \i_MIPS/Register/n1101 ) );
  OAI2BB2XL U7609 ( .B0(n3685), .B1(n3778), .A0N(
        \i_MIPS/Register/register[1][21] ), .A1N(n3778), .Y(
        \i_MIPS/Register/n1097 ) );
  OAI2BB2XL U7610 ( .B0(n3636), .B1(n3778), .A0N(
        \i_MIPS/Register/register[1][19] ), .A1N(n3777), .Y(
        \i_MIPS/Register/n1095 ) );
  OAI2BB2XL U7611 ( .B0(n3642), .B1(n49), .A0N(
        \i_MIPS/Register/register[2][29] ), .A1N(n3776), .Y(
        \i_MIPS/Register/n1073 ) );
  OAI2BB2XL U7612 ( .B0(n3640), .B1(n48), .A0N(
        \i_MIPS/Register/register[3][30] ), .A1N(n3772), .Y(
        \i_MIPS/Register/n1042 ) );
  OAI2BB2XL U7613 ( .B0(n3645), .B1(n3771), .A0N(
        \i_MIPS/Register/register[3][27] ), .A1N(n3773), .Y(
        \i_MIPS/Register/n1039 ) );
  OAI2BB2XL U7614 ( .B0(n3676), .B1(n3772), .A0N(
        \i_MIPS/Register/register[3][25] ), .A1N(n3773), .Y(
        \i_MIPS/Register/n1037 ) );
  OAI2BB2XL U7615 ( .B0(n3685), .B1(n3772), .A0N(
        \i_MIPS/Register/register[3][21] ), .A1N(n3773), .Y(
        \i_MIPS/Register/n1033 ) );
  OAI2BB2XL U7616 ( .B0(n3636), .B1(n3772), .A0N(
        \i_MIPS/Register/register[3][19] ), .A1N(n3772), .Y(
        \i_MIPS/Register/n1031 ) );
  OAI2BB2XL U7617 ( .B0(n3642), .B1(n47), .A0N(
        \i_MIPS/Register/register[4][29] ), .A1N(n3770), .Y(
        \i_MIPS/Register/n1009 ) );
  OAI2BB2XL U7618 ( .B0(n3640), .B1(n46), .A0N(
        \i_MIPS/Register/register[5][30] ), .A1N(n3766), .Y(
        \i_MIPS/Register/n978 ) );
  OAI2BB2XL U7619 ( .B0(n3645), .B1(n3766), .A0N(
        \i_MIPS/Register/register[5][27] ), .A1N(n3767), .Y(
        \i_MIPS/Register/n975 ) );
  OAI2BB2XL U7620 ( .B0(n3676), .B1(n46), .A0N(
        \i_MIPS/Register/register[5][25] ), .A1N(n3767), .Y(
        \i_MIPS/Register/n973 ) );
  OAI2BB2XL U7621 ( .B0(n3685), .B1(n3766), .A0N(
        \i_MIPS/Register/register[5][21] ), .A1N(n3766), .Y(
        \i_MIPS/Register/n969 ) );
  OAI2BB2XL U7622 ( .B0(n3636), .B1(n3766), .A0N(
        \i_MIPS/Register/register[5][19] ), .A1N(n3765), .Y(
        \i_MIPS/Register/n967 ) );
  OAI2BB2XL U7623 ( .B0(n3642), .B1(n45), .A0N(
        \i_MIPS/Register/register[6][29] ), .A1N(n3764), .Y(
        \i_MIPS/Register/n945 ) );
  OAI2BB2XL U7624 ( .B0(n3640), .B1(n43), .A0N(
        \i_MIPS/Register/register[8][30] ), .A1N(n3756), .Y(
        \i_MIPS/Register/n882 ) );
  OAI2BB2XL U7625 ( .B0(n3642), .B1(n43), .A0N(
        \i_MIPS/Register/register[8][29] ), .A1N(n3758), .Y(
        \i_MIPS/Register/n881 ) );
  OAI2BB2XL U7626 ( .B0(n3645), .B1(n43), .A0N(
        \i_MIPS/Register/register[8][27] ), .A1N(n3758), .Y(
        \i_MIPS/Register/n879 ) );
  OAI2BB2XL U7627 ( .B0(n3676), .B1(n43), .A0N(
        \i_MIPS/Register/register[8][25] ), .A1N(n3758), .Y(
        \i_MIPS/Register/n877 ) );
  OAI2BB2XL U7628 ( .B0(n3685), .B1(n3757), .A0N(
        \i_MIPS/Register/register[8][21] ), .A1N(n3757), .Y(
        \i_MIPS/Register/n873 ) );
  OAI2BB2XL U7629 ( .B0(n3636), .B1(n3757), .A0N(
        \i_MIPS/Register/register[8][19] ), .A1N(n3758), .Y(
        \i_MIPS/Register/n871 ) );
  OAI2BB2XL U7630 ( .B0(n3640), .B1(n41), .A0N(
        \i_MIPS/Register/register[10][30] ), .A1N(n3751), .Y(
        \i_MIPS/Register/n818 ) );
  OAI2BB2XL U7631 ( .B0(n3642), .B1(n41), .A0N(
        \i_MIPS/Register/register[10][29] ), .A1N(n3752), .Y(
        \i_MIPS/Register/n817 ) );
  OAI2BB2XL U7632 ( .B0(n3645), .B1(n3751), .A0N(
        \i_MIPS/Register/register[10][27] ), .A1N(n3752), .Y(
        \i_MIPS/Register/n815 ) );
  OAI2BB2XL U7633 ( .B0(n3676), .B1(n3750), .A0N(
        \i_MIPS/Register/register[10][25] ), .A1N(n3752), .Y(
        \i_MIPS/Register/n813 ) );
  OAI2BB2XL U7634 ( .B0(n3685), .B1(n3751), .A0N(
        \i_MIPS/Register/register[10][21] ), .A1N(n3752), .Y(
        \i_MIPS/Register/n809 ) );
  OAI2BB2XL U7635 ( .B0(n3636), .B1(n3751), .A0N(
        \i_MIPS/Register/register[10][19] ), .A1N(n3750), .Y(
        \i_MIPS/Register/n807 ) );
  OAI2BB2XL U7636 ( .B0(n3640), .B1(n39), .A0N(
        \i_MIPS/Register/register[12][30] ), .A1N(n3745), .Y(
        \i_MIPS/Register/n754 ) );
  OAI2BB2XL U7637 ( .B0(n3645), .B1(n3744), .A0N(
        \i_MIPS/Register/register[12][27] ), .A1N(n3746), .Y(
        \i_MIPS/Register/n751 ) );
  OAI2BB2XL U7638 ( .B0(n3676), .B1(n39), .A0N(
        \i_MIPS/Register/register[12][25] ), .A1N(n3746), .Y(
        \i_MIPS/Register/n749 ) );
  OAI2BB2XL U7639 ( .B0(n3685), .B1(n3745), .A0N(
        \i_MIPS/Register/register[12][21] ), .A1N(n3746), .Y(
        \i_MIPS/Register/n745 ) );
  OAI2BB2XL U7640 ( .B0(n3636), .B1(n3745), .A0N(
        \i_MIPS/Register/register[12][19] ), .A1N(n3744), .Y(
        \i_MIPS/Register/n743 ) );
  OAI2BB2XL U7641 ( .B0(n3642), .B1(n38), .A0N(
        \i_MIPS/Register/register[13][29] ), .A1N(n3743), .Y(
        \i_MIPS/Register/n721 ) );
  OAI2BB2XL U7642 ( .B0(n3642), .B1(n37), .A0N(
        \i_MIPS/Register/register[14][29] ), .A1N(n3740), .Y(
        \i_MIPS/Register/n689 ) );
  OAI2BB2XL U7643 ( .B0(n3640), .B1(n36), .A0N(
        \i_MIPS/Register/register[15][30] ), .A1N(n3735), .Y(
        \i_MIPS/Register/n658 ) );
  OAI2BB2XL U7644 ( .B0(n3645), .B1(n3735), .A0N(
        \i_MIPS/Register/register[15][27] ), .A1N(n3737), .Y(
        \i_MIPS/Register/n655 ) );
  OAI2BB2XL U7645 ( .B0(n3676), .B1(n36), .A0N(
        \i_MIPS/Register/register[15][25] ), .A1N(n3737), .Y(
        \i_MIPS/Register/n653 ) );
  OAI2BB2XL U7646 ( .B0(n3685), .B1(n3736), .A0N(
        \i_MIPS/Register/register[15][21] ), .A1N(n3735), .Y(
        \i_MIPS/Register/n649 ) );
  OAI2BB2XL U7647 ( .B0(n3636), .B1(n3736), .A0N(
        \i_MIPS/Register/register[15][19] ), .A1N(n3736), .Y(
        \i_MIPS/Register/n647 ) );
  OAI2BB2XL U7648 ( .B0(n3642), .B1(n35), .A0N(
        \i_MIPS/Register/register[16][29] ), .A1N(n3734), .Y(
        \i_MIPS/Register/n625 ) );
  OAI2BB2XL U7649 ( .B0(n3640), .B1(n34), .A0N(
        \i_MIPS/Register/register[17][30] ), .A1N(n3729), .Y(
        \i_MIPS/Register/n594 ) );
  OAI2BB2XL U7650 ( .B0(n3645), .B1(n3730), .A0N(
        \i_MIPS/Register/register[17][27] ), .A1N(n3731), .Y(
        \i_MIPS/Register/n591 ) );
  OAI2BB2XL U7651 ( .B0(n3676), .B1(n34), .A0N(
        \i_MIPS/Register/register[17][25] ), .A1N(n3731), .Y(
        \i_MIPS/Register/n589 ) );
  OAI2BB2XL U7652 ( .B0(n3685), .B1(n3730), .A0N(
        \i_MIPS/Register/register[17][21] ), .A1N(n3730), .Y(
        \i_MIPS/Register/n585 ) );
  OAI2BB2XL U7653 ( .B0(n3636), .B1(n3730), .A0N(
        \i_MIPS/Register/register[17][19] ), .A1N(n3729), .Y(
        \i_MIPS/Register/n583 ) );
  OAI2BB2XL U7654 ( .B0(n3640), .B1(n32), .A0N(
        \i_MIPS/Register/register[19][30] ), .A1N(n3723), .Y(
        \i_MIPS/Register/n530 ) );
  OAI2BB2XL U7655 ( .B0(n3642), .B1(n32), .A0N(
        \i_MIPS/Register/register[19][29] ), .A1N(n3725), .Y(
        \i_MIPS/Register/n529 ) );
  OAI2BB2XL U7656 ( .B0(n3645), .B1(n32), .A0N(
        \i_MIPS/Register/register[19][27] ), .A1N(n3725), .Y(
        \i_MIPS/Register/n527 ) );
  OAI2BB2XL U7657 ( .B0(n3676), .B1(n32), .A0N(
        \i_MIPS/Register/register[19][25] ), .A1N(n3725), .Y(
        \i_MIPS/Register/n525 ) );
  OAI2BB2XL U7658 ( .B0(n3685), .B1(n3724), .A0N(
        \i_MIPS/Register/register[19][21] ), .A1N(n3725), .Y(
        \i_MIPS/Register/n521 ) );
  OAI2BB2XL U7659 ( .B0(n3636), .B1(n3724), .A0N(
        \i_MIPS/Register/register[19][19] ), .A1N(n3724), .Y(
        \i_MIPS/Register/n519 ) );
  OAI2BB2XL U7660 ( .B0(n3640), .B1(n30), .A0N(
        \i_MIPS/Register/register[21][30] ), .A1N(n3717), .Y(
        \i_MIPS/Register/n466 ) );
  OAI2BB2XL U7661 ( .B0(n3642), .B1(n30), .A0N(
        \i_MIPS/Register/register[21][29] ), .A1N(n3719), .Y(
        \i_MIPS/Register/n465 ) );
  OAI2BB2XL U7662 ( .B0(n3645), .B1(n30), .A0N(
        \i_MIPS/Register/register[21][27] ), .A1N(n3719), .Y(
        \i_MIPS/Register/n463 ) );
  OAI2BB2XL U7663 ( .B0(n3676), .B1(n30), .A0N(
        \i_MIPS/Register/register[21][25] ), .A1N(n3719), .Y(
        \i_MIPS/Register/n461 ) );
  OAI2BB2XL U7664 ( .B0(n3685), .B1(n3718), .A0N(
        \i_MIPS/Register/register[21][21] ), .A1N(n3719), .Y(
        \i_MIPS/Register/n457 ) );
  OAI2BB2XL U7665 ( .B0(n3636), .B1(n3718), .A0N(
        \i_MIPS/Register/register[21][19] ), .A1N(n3718), .Y(
        \i_MIPS/Register/n455 ) );
  OAI2BB2XL U7666 ( .B0(n3640), .B1(n28), .A0N(
        \i_MIPS/Register/register[23][30] ), .A1N(n3711), .Y(
        \i_MIPS/Register/n402 ) );
  OAI2BB2XL U7667 ( .B0(n3641), .B1(n3712), .A0N(
        \i_MIPS/Register/register[23][29] ), .A1N(n3713), .Y(
        \i_MIPS/Register/n401 ) );
  OAI2BB2XL U7668 ( .B0(n3645), .B1(n28), .A0N(
        \i_MIPS/Register/register[23][27] ), .A1N(n3713), .Y(
        \i_MIPS/Register/n399 ) );
  OAI2BB2XL U7669 ( .B0(n3676), .B1(n28), .A0N(
        \i_MIPS/Register/register[23][25] ), .A1N(n3713), .Y(
        \i_MIPS/Register/n397 ) );
  OAI2BB2XL U7670 ( .B0(n3685), .B1(n3712), .A0N(
        \i_MIPS/Register/register[23][21] ), .A1N(n3713), .Y(
        \i_MIPS/Register/n393 ) );
  OAI2BB2XL U7671 ( .B0(n3636), .B1(n3712), .A0N(
        \i_MIPS/Register/register[23][19] ), .A1N(n3712), .Y(
        \i_MIPS/Register/n391 ) );
  OAI2BB2XL U7672 ( .B0(n3639), .B1(n3706), .A0N(
        \i_MIPS/Register/register[25][30] ), .A1N(n3706), .Y(
        \i_MIPS/Register/n338 ) );
  OAI2BB2XL U7673 ( .B0(n3641), .B1(\i_MIPS/Register/n116 ), .A0N(
        \i_MIPS/Register/register[25][29] ), .A1N(n3707), .Y(
        \i_MIPS/Register/n337 ) );
  OAI2BB2XL U7674 ( .B0(n3644), .B1(\i_MIPS/Register/n116 ), .A0N(
        \i_MIPS/Register/register[25][27] ), .A1N(n3707), .Y(
        \i_MIPS/Register/n335 ) );
  OAI2BB2XL U7675 ( .B0(n3675), .B1(\i_MIPS/Register/n116 ), .A0N(
        \i_MIPS/Register/register[25][25] ), .A1N(n3707), .Y(
        \i_MIPS/Register/n333 ) );
  OAI2BB2XL U7676 ( .B0(n3684), .B1(n3706), .A0N(
        \i_MIPS/Register/register[25][21] ), .A1N(n3707), .Y(
        \i_MIPS/Register/n329 ) );
  OAI2BB2XL U7677 ( .B0(n3635), .B1(n3706), .A0N(
        \i_MIPS/Register/register[25][19] ), .A1N(n3705), .Y(
        \i_MIPS/Register/n327 ) );
  OAI2BB2XL U7678 ( .B0(n3639), .B1(n3700), .A0N(
        \i_MIPS/Register/register[27][30] ), .A1N(n3700), .Y(
        \i_MIPS/Register/n274 ) );
  OAI2BB2XL U7679 ( .B0(n3642), .B1(\i_MIPS/Register/n112 ), .A0N(
        \i_MIPS/Register/register[27][29] ), .A1N(n3701), .Y(
        \i_MIPS/Register/n273 ) );
  OAI2BB2XL U7680 ( .B0(n3644), .B1(\i_MIPS/Register/n112 ), .A0N(
        \i_MIPS/Register/register[27][27] ), .A1N(n3701), .Y(
        \i_MIPS/Register/n271 ) );
  OAI2BB2XL U7681 ( .B0(n3675), .B1(\i_MIPS/Register/n112 ), .A0N(
        \i_MIPS/Register/register[27][25] ), .A1N(n3701), .Y(
        \i_MIPS/Register/n269 ) );
  OAI2BB2XL U7682 ( .B0(n3684), .B1(n3700), .A0N(
        \i_MIPS/Register/register[27][21] ), .A1N(n3701), .Y(
        \i_MIPS/Register/n265 ) );
  OAI2BB2XL U7683 ( .B0(n3635), .B1(n3700), .A0N(
        \i_MIPS/Register/register[27][19] ), .A1N(n3699), .Y(
        \i_MIPS/Register/n263 ) );
  OAI2BB2XL U7684 ( .B0(n3640), .B1(\i_MIPS/Register/n108 ), .A0N(
        \i_MIPS/Register/register[29][30] ), .A1N(n3694), .Y(
        \i_MIPS/Register/n210 ) );
  OAI2BB2XL U7685 ( .B0(n3641), .B1(n3694), .A0N(
        \i_MIPS/Register/register[29][29] ), .A1N(n3695), .Y(
        \i_MIPS/Register/n209 ) );
  OAI2BB2XL U7686 ( .B0(n3645), .B1(\i_MIPS/Register/n108 ), .A0N(
        \i_MIPS/Register/register[29][27] ), .A1N(n3695), .Y(
        \i_MIPS/Register/n207 ) );
  OAI2BB2XL U7687 ( .B0(n3676), .B1(\i_MIPS/Register/n108 ), .A0N(
        \i_MIPS/Register/register[29][25] ), .A1N(n3695), .Y(
        \i_MIPS/Register/n205 ) );
  OAI2BB2XL U7688 ( .B0(n3685), .B1(n3694), .A0N(
        \i_MIPS/Register/register[29][21] ), .A1N(n3694), .Y(
        \i_MIPS/Register/n201 ) );
  OAI2BB2XL U7689 ( .B0(n3636), .B1(n3694), .A0N(
        \i_MIPS/Register/register[29][19] ), .A1N(n3693), .Y(
        \i_MIPS/Register/n199 ) );
  OAI2BB2XL U7690 ( .B0(n3639), .B1(n3691), .A0N(
        \i_MIPS/Register/register[30][30] ), .A1N(n3690), .Y(
        \i_MIPS/Register/n178 ) );
  OAI2BB2XL U7691 ( .B0(n3644), .B1(n3690), .A0N(
        \i_MIPS/Register/register[30][27] ), .A1N(n3692), .Y(
        \i_MIPS/Register/n175 ) );
  OAI2BB2XL U7692 ( .B0(n3675), .B1(\i_MIPS/Register/n106 ), .A0N(
        \i_MIPS/Register/register[30][25] ), .A1N(n3692), .Y(
        \i_MIPS/Register/n173 ) );
  OAI2BB2XL U7693 ( .B0(n3684), .B1(n3691), .A0N(
        \i_MIPS/Register/register[30][21] ), .A1N(n3690), .Y(
        \i_MIPS/Register/n169 ) );
  OAI2BB2XL U7694 ( .B0(n3635), .B1(n3691), .A0N(
        \i_MIPS/Register/register[30][19] ), .A1N(n3692), .Y(
        \i_MIPS/Register/n167 ) );
  OAI2BB2XL U7695 ( .B0(n3671), .B1(n3756), .A0N(
        \i_MIPS/Register/register[8][26] ), .A1N(n3758), .Y(
        \i_MIPS/Register/n878 ) );
  OAI2BB2XL U7696 ( .B0(n3674), .B1(n3757), .A0N(
        \i_MIPS/Register/register[8][24] ), .A1N(n3758), .Y(
        \i_MIPS/Register/n876 ) );
  OAI2BB2XL U7697 ( .B0(n3671), .B1(n3750), .A0N(
        \i_MIPS/Register/register[10][26] ), .A1N(n3752), .Y(
        \i_MIPS/Register/n814 ) );
  OAI2BB2XL U7698 ( .B0(n3673), .B1(n3751), .A0N(
        \i_MIPS/Register/register[10][24] ), .A1N(n3752), .Y(
        \i_MIPS/Register/n812 ) );
  OAI2BB2XL U7699 ( .B0(n3671), .B1(n3745), .A0N(
        \i_MIPS/Register/register[12][26] ), .A1N(n3746), .Y(
        \i_MIPS/Register/n750 ) );
  OAI2BB2XL U7700 ( .B0(n3674), .B1(n3745), .A0N(
        \i_MIPS/Register/register[12][24] ), .A1N(n3746), .Y(
        \i_MIPS/Register/n748 ) );
  OAI2BB2XL U7701 ( .B0(n3671), .B1(n3736), .A0N(
        \i_MIPS/Register/register[15][26] ), .A1N(n3737), .Y(
        \i_MIPS/Register/n654 ) );
  OAI2BB2XL U7702 ( .B0(n3673), .B1(n3736), .A0N(
        \i_MIPS/Register/register[15][24] ), .A1N(n3737), .Y(
        \i_MIPS/Register/n652 ) );
  OAI2BB2XL U7703 ( .B0(n3671), .B1(n3729), .A0N(
        \i_MIPS/Register/register[17][26] ), .A1N(n3731), .Y(
        \i_MIPS/Register/n590 ) );
  OAI2BB2XL U7704 ( .B0(n3673), .B1(n3730), .A0N(
        \i_MIPS/Register/register[17][24] ), .A1N(n3731), .Y(
        \i_MIPS/Register/n588 ) );
  OAI2BB2XL U7705 ( .B0(n3671), .B1(n3724), .A0N(
        \i_MIPS/Register/register[19][26] ), .A1N(n3725), .Y(
        \i_MIPS/Register/n526 ) );
  OAI2BB2XL U7706 ( .B0(n3674), .B1(n3724), .A0N(
        \i_MIPS/Register/register[19][24] ), .A1N(n3725), .Y(
        \i_MIPS/Register/n524 ) );
  OAI2BB2XL U7707 ( .B0(n3671), .B1(n3718), .A0N(
        \i_MIPS/Register/register[21][26] ), .A1N(n3719), .Y(
        \i_MIPS/Register/n462 ) );
  OAI2BB2XL U7708 ( .B0(n3673), .B1(n3718), .A0N(
        \i_MIPS/Register/register[21][24] ), .A1N(n3719), .Y(
        \i_MIPS/Register/n460 ) );
  OAI2BB2XL U7709 ( .B0(n3671), .B1(n28), .A0N(
        \i_MIPS/Register/register[23][26] ), .A1N(n3713), .Y(
        \i_MIPS/Register/n398 ) );
  OAI2BB2XL U7710 ( .B0(n3674), .B1(n3712), .A0N(
        \i_MIPS/Register/register[23][24] ), .A1N(n3713), .Y(
        \i_MIPS/Register/n396 ) );
  OAI2BB2XL U7711 ( .B0(n3671), .B1(\i_MIPS/Register/n116 ), .A0N(
        \i_MIPS/Register/register[25][26] ), .A1N(n3707), .Y(
        \i_MIPS/Register/n334 ) );
  OAI2BB2XL U7712 ( .B0(n3673), .B1(n3706), .A0N(
        \i_MIPS/Register/register[25][24] ), .A1N(n3707), .Y(
        \i_MIPS/Register/n332 ) );
  OAI2BB2XL U7713 ( .B0(n3671), .B1(\i_MIPS/Register/n112 ), .A0N(
        \i_MIPS/Register/register[27][26] ), .A1N(n3701), .Y(
        \i_MIPS/Register/n270 ) );
  OAI2BB2XL U7714 ( .B0(n3674), .B1(n3700), .A0N(
        \i_MIPS/Register/register[27][24] ), .A1N(n3701), .Y(
        \i_MIPS/Register/n268 ) );
  OAI2BB2XL U7715 ( .B0(n3671), .B1(\i_MIPS/Register/n108 ), .A0N(
        \i_MIPS/Register/register[29][26] ), .A1N(n3695), .Y(
        \i_MIPS/Register/n206 ) );
  OAI2BB2XL U7716 ( .B0(n3673), .B1(n3694), .A0N(
        \i_MIPS/Register/register[29][24] ), .A1N(n3695), .Y(
        \i_MIPS/Register/n204 ) );
  OAI2BB2XL U7717 ( .B0(n3671), .B1(\i_MIPS/Register/n106 ), .A0N(
        \i_MIPS/Register/register[30][26] ), .A1N(n3692), .Y(
        \i_MIPS/Register/n174 ) );
  OAI2BB2XL U7718 ( .B0(n3673), .B1(n3691), .A0N(
        \i_MIPS/Register/register[30][24] ), .A1N(n3692), .Y(
        \i_MIPS/Register/n172 ) );
  OAI2BB2XL U7719 ( .B0(n3672), .B1(n44), .A0N(
        \i_MIPS/Register/register[7][26] ), .A1N(n3761), .Y(
        \i_MIPS/Register/n910 ) );
  OAI2BB2XL U7720 ( .B0(n3673), .B1(n3760), .A0N(
        \i_MIPS/Register/register[7][24] ), .A1N(n3761), .Y(
        \i_MIPS/Register/n908 ) );
  OAI2BB2XL U7721 ( .B0(n3672), .B1(n42), .A0N(
        \i_MIPS/Register/register[9][26] ), .A1N(n3755), .Y(
        \i_MIPS/Register/n846 ) );
  OAI2BB2XL U7722 ( .B0(n3674), .B1(n3754), .A0N(
        \i_MIPS/Register/register[9][24] ), .A1N(n3755), .Y(
        \i_MIPS/Register/n844 ) );
  OAI2BB2XL U7723 ( .B0(n3672), .B1(n40), .A0N(
        \i_MIPS/Register/register[11][26] ), .A1N(n3749), .Y(
        \i_MIPS/Register/n782 ) );
  OAI2BB2XL U7724 ( .B0(n3673), .B1(n3748), .A0N(
        \i_MIPS/Register/register[11][24] ), .A1N(n3749), .Y(
        \i_MIPS/Register/n780 ) );
  OAI2BB2XL U7725 ( .B0(n3672), .B1(n38), .A0N(
        \i_MIPS/Register/register[13][26] ), .A1N(n3743), .Y(
        \i_MIPS/Register/n718 ) );
  OAI2BB2XL U7726 ( .B0(n3674), .B1(n3742), .A0N(
        \i_MIPS/Register/register[13][24] ), .A1N(n3743), .Y(
        \i_MIPS/Register/n716 ) );
  OAI2BB2XL U7727 ( .B0(n3672), .B1(n37), .A0N(
        \i_MIPS/Register/register[14][26] ), .A1N(n3740), .Y(
        \i_MIPS/Register/n686 ) );
  OAI2BB2XL U7728 ( .B0(n3673), .B1(n3739), .A0N(
        \i_MIPS/Register/register[14][24] ), .A1N(n3740), .Y(
        \i_MIPS/Register/n684 ) );
  OAI2BB2XL U7729 ( .B0(n3672), .B1(n35), .A0N(
        \i_MIPS/Register/register[16][26] ), .A1N(n3734), .Y(
        \i_MIPS/Register/n622 ) );
  OAI2BB2XL U7730 ( .B0(n3673), .B1(n3733), .A0N(
        \i_MIPS/Register/register[16][24] ), .A1N(n3734), .Y(
        \i_MIPS/Register/n620 ) );
  OAI2BB2XL U7731 ( .B0(n3672), .B1(n33), .A0N(
        \i_MIPS/Register/register[18][26] ), .A1N(n3728), .Y(
        \i_MIPS/Register/n558 ) );
  OAI2BB2XL U7732 ( .B0(n3674), .B1(n3727), .A0N(
        \i_MIPS/Register/register[18][24] ), .A1N(n3728), .Y(
        \i_MIPS/Register/n556 ) );
  OAI2BB2XL U7733 ( .B0(n3672), .B1(n31), .A0N(
        \i_MIPS/Register/register[20][26] ), .A1N(n3722), .Y(
        \i_MIPS/Register/n494 ) );
  OAI2BB2XL U7734 ( .B0(n3673), .B1(n3721), .A0N(
        \i_MIPS/Register/register[20][24] ), .A1N(n3722), .Y(
        \i_MIPS/Register/n492 ) );
  OAI2BB2XL U7735 ( .B0(n3672), .B1(n29), .A0N(
        \i_MIPS/Register/register[22][26] ), .A1N(n3716), .Y(
        \i_MIPS/Register/n430 ) );
  OAI2BB2XL U7736 ( .B0(n3674), .B1(n3715), .A0N(
        \i_MIPS/Register/register[22][24] ), .A1N(n3716), .Y(
        \i_MIPS/Register/n428 ) );
  OAI2BB2XL U7737 ( .B0(n3672), .B1(\i_MIPS/Register/n118 ), .A0N(
        \i_MIPS/Register/register[24][26] ), .A1N(n3710), .Y(
        \i_MIPS/Register/n366 ) );
  OAI2BB2XL U7738 ( .B0(n3673), .B1(n3709), .A0N(
        \i_MIPS/Register/register[24][24] ), .A1N(n3710), .Y(
        \i_MIPS/Register/n364 ) );
  OAI2BB2XL U7739 ( .B0(n3672), .B1(\i_MIPS/Register/n114 ), .A0N(
        \i_MIPS/Register/register[26][26] ), .A1N(n3704), .Y(
        \i_MIPS/Register/n302 ) );
  OAI2BB2XL U7740 ( .B0(n3674), .B1(n3703), .A0N(
        \i_MIPS/Register/register[26][24] ), .A1N(n3704), .Y(
        \i_MIPS/Register/n300 ) );
  OAI2BB2XL U7741 ( .B0(n3671), .B1(\i_MIPS/Register/n110 ), .A0N(
        \i_MIPS/Register/register[28][26] ), .A1N(n3698), .Y(
        \i_MIPS/Register/n238 ) );
  OAI2BB2XL U7742 ( .B0(n3674), .B1(n3697), .A0N(
        \i_MIPS/Register/register[28][24] ), .A1N(n3698), .Y(
        \i_MIPS/Register/n236 ) );
  MXI3X1 U7743 ( .A(n6531), .B(n6530), .C(n6529), .S0(\i_MIPS/ID_EX[80] ), 
        .S1(n4016), .Y(n6545) );
  CLKINVX1 U7744 ( .A(n6527), .Y(n6531) );
  NOR4BX1 U7745 ( .AN(n5058), .B(n5057), .C(n5056), .D(n5055), .Y(n5059) );
  AND3X2 U7746 ( .A(n5054), .B(\i_MIPS/ID_EX[83] ), .C(n2708), .Y(n5055) );
  AOI2BB1X1 U7747 ( .A0N(n6905), .A1N(n6204), .B0(n6907), .Y(n5056) );
  MXI2X1 U7748 ( .A(\i_MIPS/ID_EX[52] ), .B(\i_MIPS/ID_EX[84] ), .S0(n4019), 
        .Y(n4692) );
  MXI2X1 U7749 ( .A(\i_MIPS/ID_EX[62] ), .B(\i_MIPS/ID_EX[94] ), .S0(n4018), 
        .Y(n4631) );
  MXI2X1 U7750 ( .A(\i_MIPS/ID_EX[67] ), .B(\i_MIPS/ID_EX[99] ), .S0(n4018), 
        .Y(n4629) );
  MXI2X1 U7751 ( .A(\i_MIPS/ID_EX[65] ), .B(\i_MIPS/ID_EX[97] ), .S0(n4018), 
        .Y(n4635) );
  MXI2X1 U7752 ( .A(\i_MIPS/ID_EX[63] ), .B(\i_MIPS/ID_EX[95] ), .S0(n4018), 
        .Y(n4632) );
  MXI2X1 U7753 ( .A(\i_MIPS/ID_EX[69] ), .B(\i_MIPS/ID_EX[101] ), .S0(n4018), 
        .Y(n4624) );
  MXI2X1 U7754 ( .A(\i_MIPS/ID_EX[66] ), .B(\i_MIPS/ID_EX[98] ), .S0(n4018), 
        .Y(n4628) );
  MXI2X1 U7755 ( .A(\i_MIPS/ID_EX[70] ), .B(\i_MIPS/ID_EX[102] ), .S0(n4018), 
        .Y(n4623) );
  MXI2X1 U7756 ( .A(\i_MIPS/ID_EX[64] ), .B(\i_MIPS/ID_EX[96] ), .S0(n4018), 
        .Y(n4636) );
  MXI2X1 U7757 ( .A(\i_MIPS/ID_EX[68] ), .B(\i_MIPS/ID_EX[100] ), .S0(n4018), 
        .Y(n4625) );
  MXI2X1 U7758 ( .A(\i_MIPS/ID_EX[61] ), .B(\i_MIPS/ID_EX[93] ), .S0(n4018), 
        .Y(n4642) );
  MXI2X1 U7759 ( .A(\i_MIPS/ID_EX[71] ), .B(\i_MIPS/ID_EX[103] ), .S0(n4018), 
        .Y(n4706) );
  NAND2X1 U7760 ( .A(\i_MIPS/ALUin1[30] ), .B(n4706), .Y(n8459) );
  OAI2BB2XL U7761 ( .B0(n3667), .B1(n3759), .A0N(
        \i_MIPS/Register/register[7][6] ), .A1N(n3761), .Y(
        \i_MIPS/Register/n890 ) );
  OAI2BB2XL U7762 ( .B0(n3667), .B1(n3756), .A0N(
        \i_MIPS/Register/register[8][6] ), .A1N(n3758), .Y(
        \i_MIPS/Register/n858 ) );
  OAI2BB2XL U7763 ( .B0(n3667), .B1(n3753), .A0N(
        \i_MIPS/Register/register[9][6] ), .A1N(n3755), .Y(
        \i_MIPS/Register/n826 ) );
  OAI2BB2XL U7764 ( .B0(n3667), .B1(n3750), .A0N(
        \i_MIPS/Register/register[10][6] ), .A1N(n3752), .Y(
        \i_MIPS/Register/n794 ) );
  OAI2BB2XL U7765 ( .B0(n3667), .B1(n3747), .A0N(
        \i_MIPS/Register/register[11][6] ), .A1N(n3749), .Y(
        \i_MIPS/Register/n762 ) );
  OAI2BB2XL U7766 ( .B0(n3667), .B1(n3744), .A0N(
        \i_MIPS/Register/register[12][6] ), .A1N(n3746), .Y(
        \i_MIPS/Register/n730 ) );
  OAI2BB2XL U7767 ( .B0(n3667), .B1(n3741), .A0N(
        \i_MIPS/Register/register[13][6] ), .A1N(n3743), .Y(
        \i_MIPS/Register/n698 ) );
  OAI2BB2XL U7768 ( .B0(n3667), .B1(n3738), .A0N(
        \i_MIPS/Register/register[14][6] ), .A1N(n3740), .Y(
        \i_MIPS/Register/n666 ) );
  OAI2BB2XL U7769 ( .B0(n3667), .B1(n3735), .A0N(
        \i_MIPS/Register/register[15][6] ), .A1N(n3737), .Y(
        \i_MIPS/Register/n634 ) );
  OAI2BB2XL U7770 ( .B0(n3667), .B1(n3732), .A0N(
        \i_MIPS/Register/register[16][6] ), .A1N(n3734), .Y(
        \i_MIPS/Register/n602 ) );
  OAI2BB2XL U7771 ( .B0(n3667), .B1(n3729), .A0N(
        \i_MIPS/Register/register[17][6] ), .A1N(n3731), .Y(
        \i_MIPS/Register/n570 ) );
  OAI2BB2XL U7772 ( .B0(n3667), .B1(n3690), .A0N(
        \i_MIPS/Register/register[30][6] ), .A1N(n3692), .Y(
        \i_MIPS/Register/n154 ) );
  NAND2X1 U7773 ( .A(\i_MIPS/ALUin1[19] ), .B(n4644), .Y(n5602) );
  NOR4X4 U7774 ( .A(\D_cache/n536 ), .B(\D_cache/n537 ), .C(\D_cache/n538 ), 
        .D(\D_cache/n539 ), .Y(\D_cache/n526 ) );
  MXI2X1 U7775 ( .A(\i_MIPS/EX_MEM[6] ), .B(DCACHE_rdata[1]), .S0(n4022), .Y(
        n8732) );
  NAND3X2 U7776 ( .A(ICACHE_addr[8]), .B(ICACHE_addr[7]), .C(n7816), .Y(n7892)
         );
  NAND3X2 U7777 ( .A(ICACHE_addr[10]), .B(ICACHE_addr[9]), .C(n7916), .Y(n7928) );
  OAI2BB2XL U7778 ( .B0(n3650), .B1(n3781), .A0N(
        \i_MIPS/Register/register[0][13] ), .A1N(n3782), .Y(
        \i_MIPS/Register/n1121 ) );
  OAI2BB2XL U7779 ( .B0(n3650), .B1(n3778), .A0N(
        \i_MIPS/Register/register[1][13] ), .A1N(n3779), .Y(
        \i_MIPS/Register/n1089 ) );
  OAI2BB2XL U7780 ( .B0(n3650), .B1(n3775), .A0N(
        \i_MIPS/Register/register[2][13] ), .A1N(n3776), .Y(
        \i_MIPS/Register/n1057 ) );
  OAI2BB2XL U7781 ( .B0(n3650), .B1(n3769), .A0N(
        \i_MIPS/Register/register[4][13] ), .A1N(n3770), .Y(
        \i_MIPS/Register/n993 ) );
  OAI2BB2XL U7782 ( .B0(n3650), .B1(n3763), .A0N(
        \i_MIPS/Register/register[6][13] ), .A1N(n3764), .Y(
        \i_MIPS/Register/n929 ) );
  OAI2BB2XL U7783 ( .B0(n3647), .B1(n3781), .A0N(
        \i_MIPS/Register/register[0][15] ), .A1N(n3782), .Y(
        \i_MIPS/Register/n1123 ) );
  OAI2BB2XL U7784 ( .B0(n3647), .B1(n3778), .A0N(
        \i_MIPS/Register/register[1][15] ), .A1N(n3779), .Y(
        \i_MIPS/Register/n1091 ) );
  OAI2BB2XL U7785 ( .B0(n3647), .B1(n3775), .A0N(
        \i_MIPS/Register/register[2][15] ), .A1N(n3776), .Y(
        \i_MIPS/Register/n1059 ) );
  OAI2BB2XL U7786 ( .B0(n3647), .B1(n3772), .A0N(
        \i_MIPS/Register/register[3][15] ), .A1N(n3771), .Y(
        \i_MIPS/Register/n1027 ) );
  OAI2BB2XL U7787 ( .B0(n3647), .B1(n3769), .A0N(
        \i_MIPS/Register/register[4][15] ), .A1N(n3768), .Y(
        \i_MIPS/Register/n995 ) );
  OAI2BB2XL U7788 ( .B0(n3647), .B1(n3766), .A0N(
        \i_MIPS/Register/register[5][15] ), .A1N(n3767), .Y(
        \i_MIPS/Register/n963 ) );
  OAI2BB2XL U7789 ( .B0(n3647), .B1(n3763), .A0N(
        \i_MIPS/Register/register[6][15] ), .A1N(n3762), .Y(
        \i_MIPS/Register/n931 ) );
  OAI2BB2XL U7790 ( .B0(n3647), .B1(n3727), .A0N(
        \i_MIPS/Register/register[18][15] ), .A1N(n3728), .Y(
        \i_MIPS/Register/n547 ) );
  OAI2BB2XL U7791 ( .B0(n3647), .B1(n3724), .A0N(
        \i_MIPS/Register/register[19][15] ), .A1N(n3723), .Y(
        \i_MIPS/Register/n515 ) );
  OAI2BB2XL U7792 ( .B0(n3647), .B1(n3721), .A0N(
        \i_MIPS/Register/register[20][15] ), .A1N(n3722), .Y(
        \i_MIPS/Register/n483 ) );
  OAI2BB2XL U7793 ( .B0(n3647), .B1(n3718), .A0N(
        \i_MIPS/Register/register[21][15] ), .A1N(n3717), .Y(
        \i_MIPS/Register/n451 ) );
  OAI2BB2XL U7794 ( .B0(n3647), .B1(n3715), .A0N(
        \i_MIPS/Register/register[22][15] ), .A1N(n3716), .Y(
        \i_MIPS/Register/n419 ) );
  OAI2BB2XL U7795 ( .B0(n3647), .B1(n3712), .A0N(
        \i_MIPS/Register/register[23][15] ), .A1N(n3711), .Y(
        \i_MIPS/Register/n387 ) );
  OAI2BB2XL U7796 ( .B0(n3647), .B1(n3709), .A0N(
        \i_MIPS/Register/register[24][15] ), .A1N(n3710), .Y(
        \i_MIPS/Register/n355 ) );
  OAI2BB2XL U7797 ( .B0(n3647), .B1(n3706), .A0N(
        \i_MIPS/Register/register[25][15] ), .A1N(n3707), .Y(
        \i_MIPS/Register/n323 ) );
  OAI2BB2XL U7798 ( .B0(n3647), .B1(n3703), .A0N(
        \i_MIPS/Register/register[26][15] ), .A1N(n3704), .Y(
        \i_MIPS/Register/n291 ) );
  OAI2BB2XL U7799 ( .B0(n3647), .B1(n3700), .A0N(
        \i_MIPS/Register/register[27][15] ), .A1N(n3701), .Y(
        \i_MIPS/Register/n259 ) );
  OAI2BB2XL U7800 ( .B0(n3647), .B1(n3697), .A0N(
        \i_MIPS/Register/register[28][15] ), .A1N(n3698), .Y(
        \i_MIPS/Register/n227 ) );
  OAI2BB2XL U7801 ( .B0(n3647), .B1(n3694), .A0N(
        \i_MIPS/Register/register[29][15] ), .A1N(n3695), .Y(
        \i_MIPS/Register/n195 ) );
  INVX1 U7802 ( .A(n8315), .Y(n8316) );
  OAI2BB2XL U7803 ( .B0(\i_MIPS/n232 ), .B1(n12), .A0N(n2160), .A1N(n8201), 
        .Y(\i_MIPS/N80 ) );
  OAI2BB2XL U7804 ( .B0(\i_MIPS/n231 ), .B1(n8457), .A0N(n2159), .A1N(n8179), 
        .Y(\i_MIPS/N79 ) );
  OAI2BB2XL U7805 ( .B0(\i_MIPS/n230 ), .B1(n3615), .A0N(n2159), .A1N(n8153), 
        .Y(\i_MIPS/N78 ) );
  OAI2BB2XL U7806 ( .B0(\i_MIPS/n229 ), .B1(n3611), .A0N(n2161), .A1N(n8456), 
        .Y(\i_MIPS/N77 ) );
  OAI2BB2XL U7807 ( .B0(\i_MIPS/n228 ), .B1(n3611), .A0N(n2159), .A1N(n8094), 
        .Y(\i_MIPS/N76 ) );
  OAI2BB2XL U7808 ( .B0(\i_MIPS/n227 ), .B1(n13), .A0N(n2159), .A1N(n3577), 
        .Y(\i_MIPS/N70 ) );
  OAI2BB2XL U7809 ( .B0(\i_MIPS/n226 ), .B1(n3614), .A0N(n2161), .A1N(n7985), 
        .Y(\i_MIPS/N69 ) );
  OAI2BB2XL U7810 ( .B0(\i_MIPS/n225 ), .B1(n3614), .A0N(n2160), .A1N(n7967), 
        .Y(\i_MIPS/N68 ) );
  OAI2BB2XL U7811 ( .B0(\i_MIPS/n224 ), .B1(n12), .A0N(n2160), .A1N(n7955), 
        .Y(\i_MIPS/N67 ) );
  OAI2BB2XL U7812 ( .B0(\i_MIPS/n223 ), .B1(n3614), .A0N(n2159), .A1N(n7932), 
        .Y(\i_MIPS/N66 ) );
  OAI2BB2XL U7813 ( .B0(\i_MIPS/n222 ), .B1(n3614), .A0N(n2161), .A1N(n8211), 
        .Y(\i_MIPS/N65 ) );
  OAI2BB2XL U7814 ( .B0(\i_MIPS/n221 ), .B1(n13), .A0N(n2161), .A1N(n7908), 
        .Y(\i_MIPS/N64 ) );
  OAI2BB2XL U7815 ( .B0(\i_MIPS/n220 ), .B1(n12), .A0N(n2160), .A1N(n7898), 
        .Y(\i_MIPS/N63 ) );
  OAI2BB2XL U7816 ( .B0(\i_MIPS/n219 ), .B1(n12), .A0N(n2161), .A1N(n7882), 
        .Y(\i_MIPS/N62 ) );
  OAI2BB2XL U7817 ( .B0(\i_MIPS/n218 ), .B1(n3614), .A0N(n2159), .A1N(n7862), 
        .Y(\i_MIPS/N61 ) );
  OAI2BB2XL U7818 ( .B0(\i_MIPS/n217 ), .B1(n3615), .A0N(n2161), .A1N(n7850), 
        .Y(\i_MIPS/N60 ) );
  OAI2BB2XL U7819 ( .B0(\i_MIPS/n216 ), .B1(n8457), .A0N(n2160), .A1N(n8352), 
        .Y(\i_MIPS/N59 ) );
  OAI2BB2XL U7820 ( .B0(\i_MIPS/n215 ), .B1(n3615), .A0N(n2161), .A1N(n8367), 
        .Y(\i_MIPS/N58 ) );
  OAI2BB2XL U7821 ( .B0(\i_MIPS/n213 ), .B1(n3612), .A0N(n2159), .A1N(n8335), 
        .Y(\i_MIPS/N56 ) );
  OAI2BB2XL U7822 ( .B0(\i_MIPS/n233 ), .B1(n3614), .A0N(n8278), .A1N(n2161), 
        .Y(\i_MIPS/N87 ) );
  OAI2BB2XL U7823 ( .B0(\i_MIPS/n182 ), .B1(n3613), .A0N(n2160), .A1N(
        \i_MIPS/PC/n4 ), .Y(\i_MIPS/N25 ) );
  OAI2BB2XL U7824 ( .B0(\i_MIPS/n183 ), .B1(n3612), .A0N(n2161), .A1N(n8336), 
        .Y(\i_MIPS/N26 ) );
  OAI2BB2XL U7825 ( .B0(\i_MIPS/n184 ), .B1(n3612), .A0N(n8383), .A1N(n2160), 
        .Y(\i_MIPS/N27 ) );
  OAI2BB2XL U7826 ( .B0(\i_MIPS/n185 ), .B1(n12), .A0N(n8368), .A1N(n2160), 
        .Y(\i_MIPS/N28 ) );
  OAI2BB2XL U7827 ( .B0(\i_MIPS/n186 ), .B1(n3610), .A0N(n8354), .A1N(n2161), 
        .Y(\i_MIPS/N29 ) );
  OAI2BB2XL U7828 ( .B0(\i_MIPS/n187 ), .B1(n3612), .A0N(n7851), .A1N(n2161), 
        .Y(\i_MIPS/N30 ) );
  OAI2BB2XL U7829 ( .B0(\i_MIPS/n188 ), .B1(n12), .A0N(n7863), .A1N(n2160), 
        .Y(\i_MIPS/N31 ) );
  OAI2BB2XL U7830 ( .B0(\i_MIPS/n189 ), .B1(n3610), .A0N(n7883), .A1N(n2161), 
        .Y(\i_MIPS/N32 ) );
  OAI2BB2XL U7831 ( .B0(\i_MIPS/n190 ), .B1(n3611), .A0N(n7899), .A1N(n2159), 
        .Y(\i_MIPS/N33 ) );
  OAI2BB2XL U7832 ( .B0(\i_MIPS/n191 ), .B1(n12), .A0N(n7909), .A1N(n2160), 
        .Y(\i_MIPS/N34 ) );
  OAI2BB2XL U7833 ( .B0(\i_MIPS/n192 ), .B1(n12), .A0N(n8221), .A1N(n2160), 
        .Y(\i_MIPS/N35 ) );
  OAI2BB2XL U7834 ( .B0(\i_MIPS/n193 ), .B1(n8457), .A0N(n7933), .A1N(n2159), 
        .Y(\i_MIPS/N36 ) );
  OAI2BB2XL U7835 ( .B0(\i_MIPS/n194 ), .B1(n3613), .A0N(n7956), .A1N(n2159), 
        .Y(\i_MIPS/N37 ) );
  OAI2BB2XL U7836 ( .B0(\i_MIPS/n195 ), .B1(n3610), .A0N(n7968), .A1N(n2159), 
        .Y(\i_MIPS/N38 ) );
  OAI2BB2XL U7837 ( .B0(\i_MIPS/n196 ), .B1(n8457), .A0N(n7986), .A1N(n2159), 
        .Y(\i_MIPS/N39 ) );
  OAI2BB2XL U7838 ( .B0(\i_MIPS/n197 ), .B1(n3612), .A0N(n7998), .A1N(n2161), 
        .Y(\i_MIPS/N40 ) );
  OAI2BB2XL U7839 ( .B0(\i_MIPS/n198 ), .B1(n3615), .A0N(n8026), .A1N(n2160), 
        .Y(\i_MIPS/N41 ) );
  OAI2BB2XL U7840 ( .B0(\i_MIPS/n199 ), .B1(n3610), .A0N(n8043), .A1N(n2160), 
        .Y(\i_MIPS/N42 ) );
  OAI2BB2XL U7841 ( .B0(\i_MIPS/n200 ), .B1(n3613), .A0N(n8066), .A1N(n2159), 
        .Y(\i_MIPS/N43 ) );
  OAI2BB2XL U7842 ( .B0(\i_MIPS/n201 ), .B1(n3615), .A0N(n8413), .A1N(n2161), 
        .Y(\i_MIPS/N44 ) );
  OAI2BB2XL U7843 ( .B0(\i_MIPS/n202 ), .B1(n3615), .A0N(n8091), .A1N(n2161), 
        .Y(\i_MIPS/N45 ) );
  OAI2BB2XL U7844 ( .B0(\i_MIPS/n203 ), .B1(n3613), .A0N(n8124), .A1N(n2160), 
        .Y(\i_MIPS/N46 ) );
  OAI2BB2XL U7845 ( .B0(\i_MIPS/n204 ), .B1(n3611), .A0N(n8148), .A1N(n2160), 
        .Y(\i_MIPS/N47 ) );
  OAI2BB2XL U7846 ( .B0(\i_MIPS/n205 ), .B1(n3610), .A0N(n8171), .A1N(n2159), 
        .Y(\i_MIPS/N48 ) );
  OAI2BB2XL U7847 ( .B0(\i_MIPS/n206 ), .B1(n3612), .A0N(n8197), .A1N(n2161), 
        .Y(\i_MIPS/N49 ) );
  OAI2BB2XL U7848 ( .B0(\i_MIPS/n208 ), .B1(n3615), .A0N(n8293), .A1N(n2159), 
        .Y(\i_MIPS/N51 ) );
  OAI2BB2XL U7849 ( .B0(\i_MIPS/n209 ), .B1(n13), .A0N(n8302), .A1N(n2159), 
        .Y(\i_MIPS/N52 ) );
  OAI2BB2XL U7850 ( .B0(\i_MIPS/n210 ), .B1(n3615), .A0N(n8325), .A1N(n2159), 
        .Y(\i_MIPS/N53 ) );
  OAI2BB2XL U7851 ( .B0(\i_MIPS/n236 ), .B1(n3611), .A0N(n8399), .A1N(n2160), 
        .Y(\i_MIPS/N90 ) );
  CLKINVX1 U7852 ( .A(n8401), .Y(n8399) );
  OAI2BB2XL U7853 ( .B0(\i_MIPS/n237 ), .B1(n3610), .A0N(n2160), .A1N(n8337), 
        .Y(\i_MIPS/N91 ) );
  OAI2BB2XL U7854 ( .B0(\i_MIPS/n238 ), .B1(n3612), .A0N(n2160), .A1N(n8384), 
        .Y(\i_MIPS/N92 ) );
  CLKINVX1 U7855 ( .A(n8386), .Y(n8384) );
  OAI2BB2XL U7856 ( .B0(\i_MIPS/n239 ), .B1(n3610), .A0N(n2161), .A1N(n8369), 
        .Y(\i_MIPS/N93 ) );
  CLKINVX1 U7857 ( .A(n8371), .Y(n8369) );
  OAI2BB2XL U7858 ( .B0(\i_MIPS/n240 ), .B1(n3613), .A0N(n2161), .A1N(n8355), 
        .Y(\i_MIPS/N94 ) );
  CLKINVX1 U7859 ( .A(n8357), .Y(n8355) );
  OAI2BB2XL U7860 ( .B0(\i_MIPS/n241 ), .B1(n3612), .A0N(n2159), .A1N(n7826), 
        .Y(\i_MIPS/N95 ) );
  OAI2BB2XL U7861 ( .B0(\i_MIPS/n242 ), .B1(n13), .A0N(n2159), .A1N(n7855), 
        .Y(\i_MIPS/N96 ) );
  OAI2BB2XL U7862 ( .B0(\i_MIPS/n243 ), .B1(n8457), .A0N(n2160), .A1N(n7874), 
        .Y(\i_MIPS/N97 ) );
  OAI2BB2XL U7863 ( .B0(\i_MIPS/n244 ), .B1(n3613), .A0N(n2160), .A1N(n7886), 
        .Y(\i_MIPS/N98 ) );
  OAI2BB2XL U7864 ( .B0(\i_MIPS/n245 ), .B1(n13), .A0N(n2160), .A1N(n7902), 
        .Y(\i_MIPS/N99 ) );
  OAI2BB2XL U7865 ( .B0(\i_MIPS/n159 ), .B1(n8457), .A0N(n2161), .A1N(n8213), 
        .Y(\i_MIPS/N100 ) );
  OAI2BB2XL U7866 ( .B0(\i_MIPS/n160 ), .B1(n3611), .A0N(n2161), .A1N(n7922), 
        .Y(\i_MIPS/N101 ) );
  OAI2BB2XL U7867 ( .B0(\i_MIPS/n161 ), .B1(n3614), .A0N(n2161), .A1N(n7937), 
        .Y(\i_MIPS/N102 ) );
  OAI2BB2XL U7868 ( .B0(\i_MIPS/n162 ), .B1(n13), .A0N(n2159), .A1N(n7957), 
        .Y(\i_MIPS/N103 ) );
  OAI2BB2XL U7869 ( .B0(\i_MIPS/n163 ), .B1(n8457), .A0N(n2159), .A1N(n7971), 
        .Y(\i_MIPS/N104 ) );
  OAI2BB2XL U7870 ( .B0(\i_MIPS/n164 ), .B1(n3613), .A0N(n2159), .A1N(n7988), 
        .Y(\i_MIPS/N105 ) );
  OAI2BB2XL U7871 ( .B0(\i_MIPS/n166 ), .B1(n12), .A0N(n2160), .A1N(n8028), 
        .Y(\i_MIPS/N107 ) );
  OAI2BB2XL U7872 ( .B0(\i_MIPS/n168 ), .B1(n13), .A0N(n2159), .A1N(n8414), 
        .Y(\i_MIPS/N109 ) );
  CLKINVX1 U7873 ( .A(n8418), .Y(n8414) );
  OAI2BB2XL U7874 ( .B0(\i_MIPS/n170 ), .B1(n3614), .A0N(n2161), .A1N(n8092), 
        .Y(\i_MIPS/N111 ) );
  OAI2BB2XL U7875 ( .B0(\i_MIPS/n174 ), .B1(n3613), .A0N(n2160), .A1N(n8198), 
        .Y(\i_MIPS/N115 ) );
  OAI2BB2XL U7876 ( .B0(n3025), .B1(n3781), .A0N(
        \i_MIPS/Register/register[0][18] ), .A1N(n3782), .Y(
        \i_MIPS/Register/n1126 ) );
  OAI2BB2XL U7877 ( .B0(n3038), .B1(n3780), .A0N(
        \i_MIPS/Register/register[0][8] ), .A1N(n3782), .Y(
        \i_MIPS/Register/n1116 ) );
  OAI2BB2XL U7878 ( .B0(n3663), .B1(n3780), .A0N(
        \i_MIPS/Register/register[0][2] ), .A1N(n3780), .Y(
        \i_MIPS/Register/n1110 ) );
  OAI2BB2XL U7879 ( .B0(n3025), .B1(n3778), .A0N(
        \i_MIPS/Register/register[1][18] ), .A1N(n3779), .Y(
        \i_MIPS/Register/n1094 ) );
  OAI2BB2XL U7880 ( .B0(n3038), .B1(n3777), .A0N(
        \i_MIPS/Register/register[1][8] ), .A1N(n3779), .Y(
        \i_MIPS/Register/n1084 ) );
  OAI2BB2XL U7881 ( .B0(n3663), .B1(n3777), .A0N(
        \i_MIPS/Register/register[1][2] ), .A1N(n3778), .Y(
        \i_MIPS/Register/n1078 ) );
  OAI2BB2XL U7882 ( .B0(n3025), .B1(n3775), .A0N(
        \i_MIPS/Register/register[2][18] ), .A1N(n3774), .Y(
        \i_MIPS/Register/n1062 ) );
  OAI2BB2XL U7883 ( .B0(n3038), .B1(n3774), .A0N(
        \i_MIPS/Register/register[2][8] ), .A1N(n3776), .Y(
        \i_MIPS/Register/n1052 ) );
  OAI2BB2XL U7884 ( .B0(n3663), .B1(n3774), .A0N(
        \i_MIPS/Register/register[2][2] ), .A1N(n3774), .Y(
        \i_MIPS/Register/n1046 ) );
  OAI2BB2XL U7885 ( .B0(n3661), .B1(n3772), .A0N(
        \i_MIPS/Register/register[3][18] ), .A1N(n3773), .Y(
        \i_MIPS/Register/n1030 ) );
  OAI2BB2XL U7886 ( .B0(n3687), .B1(n3771), .A0N(
        \i_MIPS/Register/register[3][8] ), .A1N(n3773), .Y(
        \i_MIPS/Register/n1020 ) );
  OAI2BB2XL U7887 ( .B0(n3663), .B1(n3771), .A0N(
        \i_MIPS/Register/register[3][2] ), .A1N(n3772), .Y(
        \i_MIPS/Register/n1014 ) );
  OAI2BB2XL U7888 ( .B0(n3025), .B1(n3760), .A0N(
        \i_MIPS/Register/register[7][18] ), .A1N(n3760), .Y(
        \i_MIPS/Register/n902 ) );
  OAI2BB2XL U7889 ( .B0(n3038), .B1(n3759), .A0N(
        \i_MIPS/Register/register[7][8] ), .A1N(n3761), .Y(
        \i_MIPS/Register/n892 ) );
  OAI2BB2XL U7890 ( .B0(n3663), .B1(n3759), .A0N(
        \i_MIPS/Register/register[7][2] ), .A1N(n3760), .Y(
        \i_MIPS/Register/n886 ) );
  OAI2BB2XL U7891 ( .B0(n3661), .B1(n3757), .A0N(
        \i_MIPS/Register/register[8][18] ), .A1N(n3757), .Y(
        \i_MIPS/Register/n870 ) );
  OAI2BB2XL U7892 ( .B0(n3687), .B1(n3756), .A0N(
        \i_MIPS/Register/register[8][8] ), .A1N(n3758), .Y(
        \i_MIPS/Register/n860 ) );
  OAI2BB2XL U7893 ( .B0(n3663), .B1(n3756), .A0N(
        \i_MIPS/Register/register[8][2] ), .A1N(n3756), .Y(
        \i_MIPS/Register/n854 ) );
  OAI2BB2XL U7894 ( .B0(n3025), .B1(n3754), .A0N(
        \i_MIPS/Register/register[9][18] ), .A1N(n3754), .Y(
        \i_MIPS/Register/n838 ) );
  OAI2BB2XL U7895 ( .B0(n3038), .B1(n3753), .A0N(
        \i_MIPS/Register/register[9][8] ), .A1N(n3755), .Y(
        \i_MIPS/Register/n828 ) );
  OAI2BB2XL U7896 ( .B0(n3663), .B1(n3753), .A0N(
        \i_MIPS/Register/register[9][2] ), .A1N(n3753), .Y(
        \i_MIPS/Register/n822 ) );
  OAI2BB2XL U7897 ( .B0(n3661), .B1(n3751), .A0N(
        \i_MIPS/Register/register[10][18] ), .A1N(n3751), .Y(
        \i_MIPS/Register/n806 ) );
  OAI2BB2XL U7898 ( .B0(n3687), .B1(n3750), .A0N(
        \i_MIPS/Register/register[10][8] ), .A1N(n3752), .Y(
        \i_MIPS/Register/n796 ) );
  OAI2BB2XL U7899 ( .B0(n3663), .B1(n3750), .A0N(
        \i_MIPS/Register/register[10][2] ), .A1N(n3750), .Y(
        \i_MIPS/Register/n790 ) );
  OAI2BB2XL U7900 ( .B0(n3025), .B1(n3748), .A0N(
        \i_MIPS/Register/register[11][18] ), .A1N(n3748), .Y(
        \i_MIPS/Register/n774 ) );
  OAI2BB2XL U7901 ( .B0(n3038), .B1(n3747), .A0N(
        \i_MIPS/Register/register[11][8] ), .A1N(n3749), .Y(
        \i_MIPS/Register/n764 ) );
  OAI2BB2XL U7902 ( .B0(n3663), .B1(n3747), .A0N(
        \i_MIPS/Register/register[11][2] ), .A1N(n3747), .Y(
        \i_MIPS/Register/n758 ) );
  OAI2BB2XL U7903 ( .B0(n3661), .B1(n3745), .A0N(
        \i_MIPS/Register/register[12][18] ), .A1N(n3745), .Y(
        \i_MIPS/Register/n742 ) );
  OAI2BB2XL U7904 ( .B0(n3687), .B1(n3744), .A0N(
        \i_MIPS/Register/register[12][8] ), .A1N(n3746), .Y(
        \i_MIPS/Register/n732 ) );
  OAI2BB2XL U7905 ( .B0(n3663), .B1(n3744), .A0N(
        \i_MIPS/Register/register[12][2] ), .A1N(n3744), .Y(
        \i_MIPS/Register/n726 ) );
  OAI2BB2XL U7906 ( .B0(n3025), .B1(n3742), .A0N(
        \i_MIPS/Register/register[13][18] ), .A1N(n3742), .Y(
        \i_MIPS/Register/n710 ) );
  OAI2BB2XL U7907 ( .B0(n3038), .B1(n3741), .A0N(
        \i_MIPS/Register/register[13][8] ), .A1N(n3743), .Y(
        \i_MIPS/Register/n700 ) );
  OAI2BB2XL U7908 ( .B0(n3663), .B1(n3741), .A0N(
        \i_MIPS/Register/register[13][2] ), .A1N(n3741), .Y(
        \i_MIPS/Register/n694 ) );
  OAI2BB2XL U7909 ( .B0(n3025), .B1(n3739), .A0N(
        \i_MIPS/Register/register[14][18] ), .A1N(n3740), .Y(
        \i_MIPS/Register/n678 ) );
  OAI2BB2XL U7910 ( .B0(n3038), .B1(n3738), .A0N(
        \i_MIPS/Register/register[14][8] ), .A1N(n3740), .Y(
        \i_MIPS/Register/n668 ) );
  OAI2BB2XL U7911 ( .B0(n3663), .B1(n3738), .A0N(
        \i_MIPS/Register/register[14][2] ), .A1N(n3738), .Y(
        \i_MIPS/Register/n662 ) );
  OAI2BB2XL U7912 ( .B0(n3661), .B1(n3736), .A0N(
        \i_MIPS/Register/register[15][18] ), .A1N(n3737), .Y(
        \i_MIPS/Register/n646 ) );
  OAI2BB2XL U7913 ( .B0(n3687), .B1(n3735), .A0N(
        \i_MIPS/Register/register[15][8] ), .A1N(n3737), .Y(
        \i_MIPS/Register/n636 ) );
  OAI2BB2XL U7914 ( .B0(n3663), .B1(n3735), .A0N(
        \i_MIPS/Register/register[15][2] ), .A1N(n3735), .Y(
        \i_MIPS/Register/n630 ) );
  OAI2BB2XL U7915 ( .B0(n3025), .B1(n3733), .A0N(
        \i_MIPS/Register/register[16][18] ), .A1N(n3734), .Y(
        \i_MIPS/Register/n614 ) );
  OAI2BB2XL U7916 ( .B0(n3038), .B1(n3732), .A0N(
        \i_MIPS/Register/register[16][8] ), .A1N(n3734), .Y(
        \i_MIPS/Register/n604 ) );
  OAI2BB2XL U7917 ( .B0(n3663), .B1(n3732), .A0N(
        \i_MIPS/Register/register[16][2] ), .A1N(n3733), .Y(
        \i_MIPS/Register/n598 ) );
  OAI2BB2XL U7918 ( .B0(n3661), .B1(n3730), .A0N(
        \i_MIPS/Register/register[17][18] ), .A1N(n3731), .Y(
        \i_MIPS/Register/n582 ) );
  OAI2BB2XL U7919 ( .B0(n3687), .B1(n3729), .A0N(
        \i_MIPS/Register/register[17][8] ), .A1N(n3731), .Y(
        \i_MIPS/Register/n572 ) );
  OAI2BB2XL U7920 ( .B0(n3663), .B1(n3729), .A0N(
        \i_MIPS/Register/register[17][2] ), .A1N(n3729), .Y(
        \i_MIPS/Register/n566 ) );
  OAI2BB2XL U7921 ( .B0(n3025), .B1(n3727), .A0N(
        \i_MIPS/Register/register[18][18] ), .A1N(n3726), .Y(
        \i_MIPS/Register/n550 ) );
  OAI2BB2XL U7922 ( .B0(n3038), .B1(n3726), .A0N(
        \i_MIPS/Register/register[18][8] ), .A1N(n3728), .Y(
        \i_MIPS/Register/n540 ) );
  OAI2BB2XL U7923 ( .B0(n3663), .B1(n3726), .A0N(
        \i_MIPS/Register/register[18][2] ), .A1N(n3727), .Y(
        \i_MIPS/Register/n534 ) );
  OAI2BB2XL U7924 ( .B0(n3661), .B1(n3724), .A0N(
        \i_MIPS/Register/register[19][18] ), .A1N(n3725), .Y(
        \i_MIPS/Register/n518 ) );
  OAI2BB2XL U7925 ( .B0(n3687), .B1(n3723), .A0N(
        \i_MIPS/Register/register[19][8] ), .A1N(n3725), .Y(
        \i_MIPS/Register/n508 ) );
  OAI2BB2XL U7926 ( .B0(n3663), .B1(n3723), .A0N(
        \i_MIPS/Register/register[19][2] ), .A1N(n3724), .Y(
        \i_MIPS/Register/n502 ) );
  OAI2BB2XL U7927 ( .B0(n3025), .B1(n3721), .A0N(
        \i_MIPS/Register/register[20][18] ), .A1N(n3720), .Y(
        \i_MIPS/Register/n486 ) );
  OAI2BB2XL U7928 ( .B0(n3038), .B1(n3720), .A0N(
        \i_MIPS/Register/register[20][8] ), .A1N(n3722), .Y(
        \i_MIPS/Register/n476 ) );
  OAI2BB2XL U7929 ( .B0(n3663), .B1(n3720), .A0N(
        \i_MIPS/Register/register[20][2] ), .A1N(n3721), .Y(
        \i_MIPS/Register/n470 ) );
  OAI2BB2XL U7930 ( .B0(n3661), .B1(n3718), .A0N(
        \i_MIPS/Register/register[21][18] ), .A1N(n3719), .Y(
        \i_MIPS/Register/n454 ) );
  OAI2BB2XL U7931 ( .B0(n3687), .B1(n3717), .A0N(
        \i_MIPS/Register/register[21][8] ), .A1N(n3719), .Y(
        \i_MIPS/Register/n444 ) );
  OAI2BB2XL U7932 ( .B0(n3663), .B1(n3717), .A0N(
        \i_MIPS/Register/register[21][2] ), .A1N(n3718), .Y(
        \i_MIPS/Register/n438 ) );
  OAI2BB2XL U7933 ( .B0(n3025), .B1(n3715), .A0N(
        \i_MIPS/Register/register[22][18] ), .A1N(n3714), .Y(
        \i_MIPS/Register/n422 ) );
  OAI2BB2XL U7934 ( .B0(n3038), .B1(n3714), .A0N(
        \i_MIPS/Register/register[22][8] ), .A1N(n3716), .Y(
        \i_MIPS/Register/n412 ) );
  OAI2BB2XL U7935 ( .B0(n3663), .B1(n3714), .A0N(
        \i_MIPS/Register/register[22][2] ), .A1N(n3715), .Y(
        \i_MIPS/Register/n406 ) );
  OAI2BB2XL U7936 ( .B0(n3661), .B1(n3712), .A0N(
        \i_MIPS/Register/register[23][18] ), .A1N(n3713), .Y(
        \i_MIPS/Register/n390 ) );
  OAI2BB2XL U7937 ( .B0(n3687), .B1(n3711), .A0N(
        \i_MIPS/Register/register[23][8] ), .A1N(n3713), .Y(
        \i_MIPS/Register/n380 ) );
  OAI2BB2XL U7938 ( .B0(n3663), .B1(n3711), .A0N(
        \i_MIPS/Register/register[23][2] ), .A1N(n3711), .Y(
        \i_MIPS/Register/n374 ) );
  OAI2BB2XL U7939 ( .B0(n3025), .B1(n3709), .A0N(
        \i_MIPS/Register/register[24][18] ), .A1N(n3708), .Y(
        \i_MIPS/Register/n358 ) );
  OAI2BB2XL U7940 ( .B0(n3038), .B1(n3708), .A0N(
        \i_MIPS/Register/register[24][8] ), .A1N(n3710), .Y(
        \i_MIPS/Register/n348 ) );
  OAI2BB2XL U7941 ( .B0(n3663), .B1(n3708), .A0N(
        \i_MIPS/Register/register[24][2] ), .A1N(n3709), .Y(
        \i_MIPS/Register/n342 ) );
  OAI2BB2XL U7942 ( .B0(n3025), .B1(n3706), .A0N(
        \i_MIPS/Register/register[25][18] ), .A1N(n3705), .Y(
        \i_MIPS/Register/n326 ) );
  OAI2BB2XL U7943 ( .B0(n3038), .B1(n3705), .A0N(
        \i_MIPS/Register/register[25][8] ), .A1N(n3707), .Y(
        \i_MIPS/Register/n316 ) );
  OAI2BB2XL U7944 ( .B0(n3663), .B1(n3705), .A0N(
        \i_MIPS/Register/register[25][2] ), .A1N(n3706), .Y(
        \i_MIPS/Register/n310 ) );
  OAI2BB2XL U7945 ( .B0(n3025), .B1(n3703), .A0N(
        \i_MIPS/Register/register[26][18] ), .A1N(n3702), .Y(
        \i_MIPS/Register/n294 ) );
  OAI2BB2XL U7946 ( .B0(n3038), .B1(n3702), .A0N(
        \i_MIPS/Register/register[26][8] ), .A1N(n3704), .Y(
        \i_MIPS/Register/n284 ) );
  OAI2BB2XL U7947 ( .B0(n3663), .B1(n3702), .A0N(
        \i_MIPS/Register/register[26][2] ), .A1N(n3703), .Y(
        \i_MIPS/Register/n278 ) );
  OAI2BB2XL U7948 ( .B0(n3025), .B1(n3700), .A0N(
        \i_MIPS/Register/register[27][18] ), .A1N(n3699), .Y(
        \i_MIPS/Register/n262 ) );
  OAI2BB2XL U7949 ( .B0(n3038), .B1(n3699), .A0N(
        \i_MIPS/Register/register[27][8] ), .A1N(n3701), .Y(
        \i_MIPS/Register/n252 ) );
  OAI2BB2XL U7950 ( .B0(n3663), .B1(n3699), .A0N(
        \i_MIPS/Register/register[27][2] ), .A1N(n3700), .Y(
        \i_MIPS/Register/n246 ) );
  OAI2BB2XL U7951 ( .B0(n3025), .B1(n3697), .A0N(
        \i_MIPS/Register/register[28][18] ), .A1N(n3696), .Y(
        \i_MIPS/Register/n230 ) );
  OAI2BB2XL U7952 ( .B0(n3038), .B1(n3696), .A0N(
        \i_MIPS/Register/register[28][8] ), .A1N(n3698), .Y(
        \i_MIPS/Register/n220 ) );
  OAI2BB2XL U7953 ( .B0(n3663), .B1(n3696), .A0N(
        \i_MIPS/Register/register[28][2] ), .A1N(n3697), .Y(
        \i_MIPS/Register/n214 ) );
  OAI2BB2XL U7954 ( .B0(n3025), .B1(n3694), .A0N(
        \i_MIPS/Register/register[29][18] ), .A1N(n3695), .Y(
        \i_MIPS/Register/n198 ) );
  OAI2BB2XL U7955 ( .B0(n3038), .B1(n3693), .A0N(
        \i_MIPS/Register/register[29][8] ), .A1N(n3695), .Y(
        \i_MIPS/Register/n188 ) );
  OAI2BB2XL U7956 ( .B0(n3663), .B1(n3693), .A0N(
        \i_MIPS/Register/register[29][2] ), .A1N(n3694), .Y(
        \i_MIPS/Register/n182 ) );
  OAI2BB2XL U7957 ( .B0(n3025), .B1(n3691), .A0N(
        \i_MIPS/Register/register[30][18] ), .A1N(n3692), .Y(
        \i_MIPS/Register/n166 ) );
  OAI2BB2XL U7958 ( .B0(n3038), .B1(n3690), .A0N(
        \i_MIPS/Register/register[30][8] ), .A1N(n3692), .Y(
        \i_MIPS/Register/n156 ) );
  OAI2BB2XL U7959 ( .B0(n3663), .B1(n3690), .A0N(
        \i_MIPS/Register/register[30][2] ), .A1N(n3690), .Y(
        \i_MIPS/Register/n150 ) );
  XNOR2X1 U7960 ( .A(\D_cache/N50 ), .B(n10315), .Y(\D_cache/n534 ) );
  XNOR2X1 U7961 ( .A(\D_cache/N52 ), .B(DCACHE_addr[9]), .Y(\D_cache/n535 ) );
  OAI2BB2XL U7962 ( .B0(n3651), .B1(n3772), .A0N(
        \i_MIPS/Register/register[3][13] ), .A1N(n3773), .Y(
        \i_MIPS/Register/n1025 ) );
  OAI2BB2XL U7963 ( .B0(n3681), .B1(n3771), .A0N(
        \i_MIPS/Register/register[3][11] ), .A1N(n3773), .Y(
        \i_MIPS/Register/n1023 ) );
  OAI2BB2XL U7964 ( .B0(n3651), .B1(n3766), .A0N(
        \i_MIPS/Register/register[5][13] ), .A1N(n3767), .Y(
        \i_MIPS/Register/n961 ) );
  OAI2BB2XL U7965 ( .B0(n3681), .B1(n3765), .A0N(
        \i_MIPS/Register/register[5][11] ), .A1N(n3767), .Y(
        \i_MIPS/Register/n959 ) );
  OAI2BB2XL U7966 ( .B0(n3650), .B1(n3760), .A0N(
        \i_MIPS/Register/register[7][13] ), .A1N(n3761), .Y(
        \i_MIPS/Register/n897 ) );
  OAI2BB2XL U7967 ( .B0(n3680), .B1(n3759), .A0N(
        \i_MIPS/Register/register[7][11] ), .A1N(n3761), .Y(
        \i_MIPS/Register/n895 ) );
  OAI2BB2XL U7968 ( .B0(n3019), .B1(n3757), .A0N(
        \i_MIPS/Register/register[8][13] ), .A1N(n3758), .Y(
        \i_MIPS/Register/n865 ) );
  OAI2BB2XL U7969 ( .B0(n3680), .B1(n3756), .A0N(
        \i_MIPS/Register/register[8][11] ), .A1N(n3758), .Y(
        \i_MIPS/Register/n863 ) );
  OAI2BB2XL U7970 ( .B0(n3019), .B1(n3754), .A0N(
        \i_MIPS/Register/register[9][13] ), .A1N(n3755), .Y(
        \i_MIPS/Register/n833 ) );
  OAI2BB2XL U7971 ( .B0(n3680), .B1(n3753), .A0N(
        \i_MIPS/Register/register[9][11] ), .A1N(n3755), .Y(
        \i_MIPS/Register/n831 ) );
  OAI2BB2XL U7972 ( .B0(n3019), .B1(n3751), .A0N(
        \i_MIPS/Register/register[10][13] ), .A1N(n3752), .Y(
        \i_MIPS/Register/n801 ) );
  OAI2BB2XL U7973 ( .B0(n3680), .B1(n3750), .A0N(
        \i_MIPS/Register/register[10][11] ), .A1N(n3752), .Y(
        \i_MIPS/Register/n799 ) );
  OAI2BB2XL U7974 ( .B0(n3019), .B1(n3748), .A0N(
        \i_MIPS/Register/register[11][13] ), .A1N(n3749), .Y(
        \i_MIPS/Register/n769 ) );
  OAI2BB2XL U7975 ( .B0(n3680), .B1(n3747), .A0N(
        \i_MIPS/Register/register[11][11] ), .A1N(n3749), .Y(
        \i_MIPS/Register/n767 ) );
  OAI2BB2XL U7976 ( .B0(n3019), .B1(n3745), .A0N(
        \i_MIPS/Register/register[12][13] ), .A1N(n3746), .Y(
        \i_MIPS/Register/n737 ) );
  OAI2BB2XL U7977 ( .B0(n3680), .B1(n3744), .A0N(
        \i_MIPS/Register/register[12][11] ), .A1N(n3746), .Y(
        \i_MIPS/Register/n735 ) );
  OAI2BB2XL U7978 ( .B0(n3019), .B1(n3742), .A0N(
        \i_MIPS/Register/register[13][13] ), .A1N(n3743), .Y(
        \i_MIPS/Register/n705 ) );
  OAI2BB2XL U7979 ( .B0(n3680), .B1(n3741), .A0N(
        \i_MIPS/Register/register[13][11] ), .A1N(n3743), .Y(
        \i_MIPS/Register/n703 ) );
  OAI2BB2XL U7980 ( .B0(n3650), .B1(n3739), .A0N(
        \i_MIPS/Register/register[14][13] ), .A1N(n3740), .Y(
        \i_MIPS/Register/n673 ) );
  OAI2BB2XL U7981 ( .B0(n3681), .B1(n3738), .A0N(
        \i_MIPS/Register/register[14][11] ), .A1N(n3740), .Y(
        \i_MIPS/Register/n671 ) );
  OAI2BB2XL U7982 ( .B0(n3650), .B1(n3736), .A0N(
        \i_MIPS/Register/register[15][13] ), .A1N(n3737), .Y(
        \i_MIPS/Register/n641 ) );
  OAI2BB2XL U7983 ( .B0(n3681), .B1(n3735), .A0N(
        \i_MIPS/Register/register[15][11] ), .A1N(n3737), .Y(
        \i_MIPS/Register/n639 ) );
  OAI2BB2XL U7984 ( .B0(n3650), .B1(n3733), .A0N(
        \i_MIPS/Register/register[16][13] ), .A1N(n3734), .Y(
        \i_MIPS/Register/n609 ) );
  OAI2BB2XL U7985 ( .B0(n3681), .B1(n3732), .A0N(
        \i_MIPS/Register/register[16][11] ), .A1N(n3734), .Y(
        \i_MIPS/Register/n607 ) );
  OAI2BB2XL U7986 ( .B0(n3650), .B1(n3730), .A0N(
        \i_MIPS/Register/register[17][13] ), .A1N(n3731), .Y(
        \i_MIPS/Register/n577 ) );
  OAI2BB2XL U7987 ( .B0(n3681), .B1(n3729), .A0N(
        \i_MIPS/Register/register[17][11] ), .A1N(n3731), .Y(
        \i_MIPS/Register/n575 ) );
  OAI2BB2XL U7988 ( .B0(n3651), .B1(n3727), .A0N(
        \i_MIPS/Register/register[18][13] ), .A1N(n3728), .Y(
        \i_MIPS/Register/n545 ) );
  OAI2BB2XL U7989 ( .B0(n3681), .B1(n3726), .A0N(
        \i_MIPS/Register/register[18][11] ), .A1N(n3728), .Y(
        \i_MIPS/Register/n543 ) );
  OAI2BB2XL U7990 ( .B0(n3651), .B1(n3724), .A0N(
        \i_MIPS/Register/register[19][13] ), .A1N(n3725), .Y(
        \i_MIPS/Register/n513 ) );
  OAI2BB2XL U7991 ( .B0(n3681), .B1(n3723), .A0N(
        \i_MIPS/Register/register[19][11] ), .A1N(n3725), .Y(
        \i_MIPS/Register/n511 ) );
  OAI2BB2XL U7992 ( .B0(n3651), .B1(n3721), .A0N(
        \i_MIPS/Register/register[20][13] ), .A1N(n3722), .Y(
        \i_MIPS/Register/n481 ) );
  OAI2BB2XL U7993 ( .B0(n3681), .B1(n3720), .A0N(
        \i_MIPS/Register/register[20][11] ), .A1N(n3722), .Y(
        \i_MIPS/Register/n479 ) );
  OAI2BB2XL U7994 ( .B0(n3651), .B1(n3718), .A0N(
        \i_MIPS/Register/register[21][13] ), .A1N(n3719), .Y(
        \i_MIPS/Register/n449 ) );
  OAI2BB2XL U7995 ( .B0(n3681), .B1(n3717), .A0N(
        \i_MIPS/Register/register[21][11] ), .A1N(n3719), .Y(
        \i_MIPS/Register/n447 ) );
  OAI2BB2XL U7996 ( .B0(n3651), .B1(n3715), .A0N(
        \i_MIPS/Register/register[22][13] ), .A1N(n3716), .Y(
        \i_MIPS/Register/n417 ) );
  OAI2BB2XL U7997 ( .B0(n3681), .B1(n3714), .A0N(
        \i_MIPS/Register/register[22][11] ), .A1N(n3716), .Y(
        \i_MIPS/Register/n415 ) );
  OAI2BB2XL U7998 ( .B0(n3651), .B1(n3712), .A0N(
        \i_MIPS/Register/register[23][13] ), .A1N(n3713), .Y(
        \i_MIPS/Register/n385 ) );
  OAI2BB2XL U7999 ( .B0(n3681), .B1(n3711), .A0N(
        \i_MIPS/Register/register[23][11] ), .A1N(n3713), .Y(
        \i_MIPS/Register/n383 ) );
  OAI2BB2XL U8000 ( .B0(n3651), .B1(n3709), .A0N(
        \i_MIPS/Register/register[24][13] ), .A1N(n3710), .Y(
        \i_MIPS/Register/n353 ) );
  OAI2BB2XL U8001 ( .B0(n3681), .B1(n3708), .A0N(
        \i_MIPS/Register/register[24][11] ), .A1N(n3710), .Y(
        \i_MIPS/Register/n351 ) );
  OAI2BB2XL U8002 ( .B0(n3651), .B1(n3706), .A0N(
        \i_MIPS/Register/register[25][13] ), .A1N(n3707), .Y(
        \i_MIPS/Register/n321 ) );
  OAI2BB2XL U8003 ( .B0(n3681), .B1(n3705), .A0N(
        \i_MIPS/Register/register[25][11] ), .A1N(n3707), .Y(
        \i_MIPS/Register/n319 ) );
  OAI2BB2XL U8004 ( .B0(n3651), .B1(n3703), .A0N(
        \i_MIPS/Register/register[26][13] ), .A1N(n3704), .Y(
        \i_MIPS/Register/n289 ) );
  OAI2BB2XL U8005 ( .B0(n3681), .B1(n3702), .A0N(
        \i_MIPS/Register/register[26][11] ), .A1N(n3704), .Y(
        \i_MIPS/Register/n287 ) );
  OAI2BB2XL U8006 ( .B0(n3651), .B1(n3700), .A0N(
        \i_MIPS/Register/register[27][13] ), .A1N(n3701), .Y(
        \i_MIPS/Register/n257 ) );
  OAI2BB2XL U8007 ( .B0(n3681), .B1(n3699), .A0N(
        \i_MIPS/Register/register[27][11] ), .A1N(n3701), .Y(
        \i_MIPS/Register/n255 ) );
  OAI2BB2XL U8008 ( .B0(n3651), .B1(n3697), .A0N(
        \i_MIPS/Register/register[28][13] ), .A1N(n3698), .Y(
        \i_MIPS/Register/n225 ) );
  OAI2BB2XL U8009 ( .B0(n3681), .B1(n3696), .A0N(
        \i_MIPS/Register/register[28][11] ), .A1N(n3698), .Y(
        \i_MIPS/Register/n223 ) );
  OAI2BB2XL U8010 ( .B0(n3651), .B1(n3694), .A0N(
        \i_MIPS/Register/register[29][13] ), .A1N(n3695), .Y(
        \i_MIPS/Register/n193 ) );
  OAI2BB2XL U8011 ( .B0(n3681), .B1(n3693), .A0N(
        \i_MIPS/Register/register[29][11] ), .A1N(n3695), .Y(
        \i_MIPS/Register/n191 ) );
  OAI2BB2XL U8012 ( .B0(n3650), .B1(n3691), .A0N(
        \i_MIPS/Register/register[30][13] ), .A1N(n3692), .Y(
        \i_MIPS/Register/n161 ) );
  OAI2BB2XL U8013 ( .B0(n3681), .B1(n3690), .A0N(
        \i_MIPS/Register/register[30][11] ), .A1N(n3692), .Y(
        \i_MIPS/Register/n159 ) );
  NAND3X4 U8014 ( .A(ICACHE_addr[22]), .B(ICACHE_addr[21]), .C(n8142), .Y(
        n8168) );
  MXI2X1 U8015 ( .A(\i_MIPS/ID_EX[111] ), .B(\i_MIPS/ID_EX[84] ), .S0(
        \i_MIPS/ID_EX_5 ), .Y(n7608) );
  OAI2BB2XL U8016 ( .B0(\D_cache/n395 ), .B1(n3789), .A0N(
        \D_cache/cache[7][59] ), .A1N(n3800), .Y(\D_cache/n1317 ) );
  OAI2BB2XL U8017 ( .B0(\D_cache/n395 ), .B1(n3809), .A0N(
        \D_cache/cache[6][59] ), .A1N(n3820), .Y(\D_cache/n1318 ) );
  OAI2BB2XL U8018 ( .B0(\D_cache/n395 ), .B1(n3828), .A0N(
        \D_cache/cache[5][59] ), .A1N(n3838), .Y(\D_cache/n1319 ) );
  OAI2BB2XL U8019 ( .B0(\D_cache/n395 ), .B1(n3847), .A0N(
        \D_cache/cache[4][59] ), .A1N(n3860), .Y(\D_cache/n1320 ) );
  OAI2BB2XL U8020 ( .B0(\D_cache/n395 ), .B1(n3866), .A0N(
        \D_cache/cache[3][59] ), .A1N(n3879), .Y(\D_cache/n1321 ) );
  OAI2BB2XL U8021 ( .B0(\D_cache/n395 ), .B1(n3889), .A0N(
        \D_cache/cache[2][59] ), .A1N(n3900), .Y(\D_cache/n1322 ) );
  OAI2BB2XL U8022 ( .B0(\D_cache/n395 ), .B1(n3909), .A0N(
        \D_cache/cache[1][59] ), .A1N(n3921), .Y(\D_cache/n1323 ) );
  OAI2BB2XL U8023 ( .B0(\D_cache/n395 ), .B1(n3929), .A0N(
        \D_cache/cache[0][59] ), .A1N(n3942), .Y(\D_cache/n1324 ) );
  OAI2BB2XL U8024 ( .B0(\D_cache/n423 ), .B1(n3791), .A0N(
        \D_cache/cache[7][45] ), .A1N(n3799), .Y(\D_cache/n1429 ) );
  OAI2BB2XL U8025 ( .B0(\D_cache/n423 ), .B1(n3811), .A0N(
        \D_cache/cache[6][45] ), .A1N(n3819), .Y(\D_cache/n1430 ) );
  OAI2BB2XL U8026 ( .B0(\D_cache/n423 ), .B1(n3829), .A0N(
        \D_cache/cache[5][45] ), .A1N(n3837), .Y(\D_cache/n1431 ) );
  OAI2BB2XL U8027 ( .B0(\D_cache/n423 ), .B1(n3849), .A0N(
        \D_cache/cache[4][45] ), .A1N(n3859), .Y(\D_cache/n1432 ) );
  OAI2BB2XL U8028 ( .B0(\D_cache/n423 ), .B1(n3868), .A0N(
        \D_cache/cache[3][45] ), .A1N(n3878), .Y(\D_cache/n1433 ) );
  OAI2BB2XL U8029 ( .B0(\D_cache/n423 ), .B1(n3891), .A0N(
        \D_cache/cache[2][45] ), .A1N(n3899), .Y(\D_cache/n1434 ) );
  OAI2BB2XL U8030 ( .B0(\D_cache/n423 ), .B1(n3911), .A0N(
        \D_cache/cache[1][45] ), .A1N(n3920), .Y(\D_cache/n1435 ) );
  OAI2BB2XL U8031 ( .B0(\D_cache/n423 ), .B1(n3931), .A0N(
        \D_cache/cache[0][45] ), .A1N(n3941), .Y(\D_cache/n1436 ) );
  OAI2BB2XL U8032 ( .B0(\D_cache/n427 ), .B1(n3794), .A0N(
        \D_cache/cache[7][43] ), .A1N(n3799), .Y(\D_cache/n1445 ) );
  OAI2BB2XL U8033 ( .B0(\D_cache/n427 ), .B1(n3814), .A0N(
        \D_cache/cache[6][43] ), .A1N(n3819), .Y(\D_cache/n1446 ) );
  OAI2BB2XL U8034 ( .B0(\D_cache/n427 ), .B1(n3832), .A0N(
        \D_cache/cache[5][43] ), .A1N(n3837), .Y(\D_cache/n1447 ) );
  OAI2BB2XL U8035 ( .B0(\D_cache/n427 ), .B1(n3854), .A0N(
        \D_cache/cache[4][43] ), .A1N(n3859), .Y(\D_cache/n1448 ) );
  OAI2BB2XL U8036 ( .B0(\D_cache/n427 ), .B1(n3873), .A0N(
        \D_cache/cache[3][43] ), .A1N(n3878), .Y(\D_cache/n1449 ) );
  OAI2BB2XL U8037 ( .B0(\D_cache/n427 ), .B1(n3894), .A0N(
        \D_cache/cache[2][43] ), .A1N(n3899), .Y(\D_cache/n1450 ) );
  OAI2BB2XL U8038 ( .B0(\D_cache/n427 ), .B1(n3915), .A0N(
        \D_cache/cache[1][43] ), .A1N(n3920), .Y(\D_cache/n1451 ) );
  OAI2BB2XL U8039 ( .B0(\D_cache/n427 ), .B1(n3936), .A0N(
        \D_cache/cache[0][43] ), .A1N(n3941), .Y(\D_cache/n1452 ) );
  OAI2BB2XL U8040 ( .B0(\D_cache/n389 ), .B1(n3789), .A0N(
        \D_cache/cache[7][62] ), .A1N(n3800), .Y(\D_cache/n1293 ) );
  OAI2BB2XL U8041 ( .B0(\D_cache/n389 ), .B1(n3809), .A0N(
        \D_cache/cache[6][62] ), .A1N(n3820), .Y(\D_cache/n1294 ) );
  OAI2BB2XL U8042 ( .B0(\D_cache/n389 ), .B1(n3828), .A0N(
        \D_cache/cache[5][62] ), .A1N(n3829), .Y(\D_cache/n1295 ) );
  OAI2BB2XL U8043 ( .B0(\D_cache/n389 ), .B1(n3847), .A0N(
        \D_cache/cache[4][62] ), .A1N(n3860), .Y(\D_cache/n1296 ) );
  OAI2BB2XL U8044 ( .B0(\D_cache/n389 ), .B1(n3866), .A0N(
        \D_cache/cache[3][62] ), .A1N(n3879), .Y(\D_cache/n1297 ) );
  OAI2BB2XL U8045 ( .B0(\D_cache/n389 ), .B1(n3889), .A0N(
        \D_cache/cache[2][62] ), .A1N(n3900), .Y(\D_cache/n1298 ) );
  OAI2BB2XL U8046 ( .B0(\D_cache/n389 ), .B1(n3909), .A0N(
        \D_cache/cache[1][62] ), .A1N(n3921), .Y(\D_cache/n1299 ) );
  OAI2BB2XL U8047 ( .B0(\D_cache/n389 ), .B1(n3929), .A0N(
        \D_cache/cache[0][62] ), .A1N(n3942), .Y(\D_cache/n1300 ) );
  OAI2BB2XL U8048 ( .B0(\D_cache/n393 ), .B1(n3789), .A0N(
        \D_cache/cache[7][60] ), .A1N(n3800), .Y(\D_cache/n1309 ) );
  OAI2BB2XL U8049 ( .B0(\D_cache/n393 ), .B1(n3809), .A0N(
        \D_cache/cache[6][60] ), .A1N(n3820), .Y(\D_cache/n1310 ) );
  OAI2BB2XL U8050 ( .B0(\D_cache/n393 ), .B1(n3828), .A0N(
        \D_cache/cache[5][60] ), .A1N(n3828), .Y(\D_cache/n1311 ) );
  OAI2BB2XL U8051 ( .B0(\D_cache/n393 ), .B1(n3847), .A0N(
        \D_cache/cache[4][60] ), .A1N(n3860), .Y(\D_cache/n1312 ) );
  OAI2BB2XL U8052 ( .B0(\D_cache/n393 ), .B1(n3866), .A0N(
        \D_cache/cache[3][60] ), .A1N(n3879), .Y(\D_cache/n1313 ) );
  OAI2BB2XL U8053 ( .B0(\D_cache/n393 ), .B1(n3889), .A0N(
        \D_cache/cache[2][60] ), .A1N(n3900), .Y(\D_cache/n1314 ) );
  OAI2BB2XL U8054 ( .B0(\D_cache/n393 ), .B1(n3909), .A0N(
        \D_cache/cache[1][60] ), .A1N(n3921), .Y(\D_cache/n1315 ) );
  OAI2BB2XL U8055 ( .B0(\D_cache/n393 ), .B1(n3929), .A0N(
        \D_cache/cache[0][60] ), .A1N(n3942), .Y(\D_cache/n1316 ) );
  OAI2BB2XL U8056 ( .B0(\D_cache/n403 ), .B1(n3789), .A0N(
        \D_cache/cache[7][55] ), .A1N(n3800), .Y(\D_cache/n1349 ) );
  OAI2BB2XL U8057 ( .B0(\D_cache/n403 ), .B1(n3809), .A0N(
        \D_cache/cache[6][55] ), .A1N(n3820), .Y(\D_cache/n1350 ) );
  OAI2BB2XL U8058 ( .B0(\D_cache/n403 ), .B1(n3828), .A0N(
        \D_cache/cache[5][55] ), .A1N(n3839), .Y(\D_cache/n1351 ) );
  OAI2BB2XL U8059 ( .B0(\D_cache/n403 ), .B1(n3847), .A0N(
        \D_cache/cache[4][55] ), .A1N(n3860), .Y(\D_cache/n1352 ) );
  OAI2BB2XL U8060 ( .B0(\D_cache/n403 ), .B1(n3866), .A0N(
        \D_cache/cache[3][55] ), .A1N(n3879), .Y(\D_cache/n1353 ) );
  OAI2BB2XL U8061 ( .B0(\D_cache/n403 ), .B1(n3889), .A0N(
        \D_cache/cache[2][55] ), .A1N(n3900), .Y(\D_cache/n1354 ) );
  OAI2BB2XL U8062 ( .B0(\D_cache/n403 ), .B1(n3909), .A0N(
        \D_cache/cache[1][55] ), .A1N(n3921), .Y(\D_cache/n1355 ) );
  OAI2BB2XL U8063 ( .B0(\D_cache/n403 ), .B1(n3929), .A0N(
        \D_cache/cache[0][55] ), .A1N(n3942), .Y(\D_cache/n1356 ) );
  OAI2BB2XL U8064 ( .B0(\D_cache/n405 ), .B1(n3790), .A0N(
        \D_cache/cache[7][54] ), .A1N(n3800), .Y(\D_cache/n1357 ) );
  OAI2BB2XL U8065 ( .B0(\D_cache/n405 ), .B1(n3810), .A0N(
        \D_cache/cache[6][54] ), .A1N(n3820), .Y(\D_cache/n1358 ) );
  OAI2BB2XL U8066 ( .B0(\D_cache/n405 ), .B1(n3829), .A0N(
        \D_cache/cache[5][54] ), .A1N(n3839), .Y(\D_cache/n1359 ) );
  OAI2BB2XL U8067 ( .B0(\D_cache/n405 ), .B1(n3848), .A0N(
        \D_cache/cache[4][54] ), .A1N(n3860), .Y(\D_cache/n1360 ) );
  OAI2BB2XL U8068 ( .B0(\D_cache/n405 ), .B1(n3867), .A0N(
        \D_cache/cache[3][54] ), .A1N(n3879), .Y(\D_cache/n1361 ) );
  OAI2BB2XL U8069 ( .B0(\D_cache/n405 ), .B1(n3890), .A0N(
        \D_cache/cache[2][54] ), .A1N(n3900), .Y(\D_cache/n1362 ) );
  OAI2BB2XL U8070 ( .B0(\D_cache/n405 ), .B1(n3910), .A0N(
        \D_cache/cache[1][54] ), .A1N(n3921), .Y(\D_cache/n1363 ) );
  OAI2BB2XL U8071 ( .B0(\D_cache/n405 ), .B1(n3930), .A0N(
        \D_cache/cache[0][54] ), .A1N(n3942), .Y(\D_cache/n1364 ) );
  OAI2BB2XL U8072 ( .B0(\D_cache/n417 ), .B1(n3790), .A0N(
        \D_cache/cache[7][48] ), .A1N(n3800), .Y(\D_cache/n1405 ) );
  OAI2BB2XL U8073 ( .B0(\D_cache/n417 ), .B1(n3810), .A0N(
        \D_cache/cache[6][48] ), .A1N(n3820), .Y(\D_cache/n1406 ) );
  OAI2BB2XL U8074 ( .B0(\D_cache/n417 ), .B1(n3828), .A0N(
        \D_cache/cache[5][48] ), .A1N(n3825), .Y(\D_cache/n1407 ) );
  OAI2BB2XL U8075 ( .B0(\D_cache/n417 ), .B1(n3848), .A0N(
        \D_cache/cache[4][48] ), .A1N(n3860), .Y(\D_cache/n1408 ) );
  OAI2BB2XL U8076 ( .B0(\D_cache/n417 ), .B1(n3867), .A0N(
        \D_cache/cache[3][48] ), .A1N(n3879), .Y(\D_cache/n1409 ) );
  OAI2BB2XL U8077 ( .B0(\D_cache/n417 ), .B1(n3890), .A0N(
        \D_cache/cache[2][48] ), .A1N(n3900), .Y(\D_cache/n1410 ) );
  OAI2BB2XL U8078 ( .B0(\D_cache/n417 ), .B1(n3910), .A0N(
        \D_cache/cache[1][48] ), .A1N(n3921), .Y(\D_cache/n1411 ) );
  OAI2BB2XL U8079 ( .B0(\D_cache/n417 ), .B1(n3930), .A0N(
        \D_cache/cache[0][48] ), .A1N(n3942), .Y(\D_cache/n1412 ) );
  OAI2BB2XL U8080 ( .B0(\D_cache/n419 ), .B1(n3790), .A0N(
        \D_cache/cache[7][47] ), .A1N(n3800), .Y(\D_cache/n1413 ) );
  OAI2BB2XL U8081 ( .B0(\D_cache/n419 ), .B1(n3810), .A0N(
        \D_cache/cache[6][47] ), .A1N(n3820), .Y(\D_cache/n1414 ) );
  OAI2BB2XL U8082 ( .B0(\D_cache/n419 ), .B1(n3827), .A0N(
        \D_cache/cache[5][47] ), .A1N(n3827), .Y(\D_cache/n1415 ) );
  OAI2BB2XL U8083 ( .B0(\D_cache/n419 ), .B1(n3848), .A0N(
        \D_cache/cache[4][47] ), .A1N(n3860), .Y(\D_cache/n1416 ) );
  OAI2BB2XL U8084 ( .B0(\D_cache/n419 ), .B1(n3867), .A0N(
        \D_cache/cache[3][47] ), .A1N(n3879), .Y(\D_cache/n1417 ) );
  OAI2BB2XL U8085 ( .B0(\D_cache/n419 ), .B1(n3890), .A0N(
        \D_cache/cache[2][47] ), .A1N(n3900), .Y(\D_cache/n1418 ) );
  OAI2BB2XL U8086 ( .B0(\D_cache/n419 ), .B1(n3910), .A0N(
        \D_cache/cache[1][47] ), .A1N(n3921), .Y(\D_cache/n1419 ) );
  OAI2BB2XL U8087 ( .B0(\D_cache/n419 ), .B1(n3930), .A0N(
        \D_cache/cache[0][47] ), .A1N(n3942), .Y(\D_cache/n1420 ) );
  OAI2BB2XL U8088 ( .B0(\D_cache/n421 ), .B1(n3791), .A0N(
        \D_cache/cache[7][46] ), .A1N(n3799), .Y(\D_cache/n1421 ) );
  OAI2BB2XL U8089 ( .B0(\D_cache/n421 ), .B1(n3811), .A0N(
        \D_cache/cache[6][46] ), .A1N(n3819), .Y(\D_cache/n1422 ) );
  OAI2BB2XL U8090 ( .B0(\D_cache/n421 ), .B1(n3829), .A0N(
        \D_cache/cache[5][46] ), .A1N(n3837), .Y(\D_cache/n1423 ) );
  OAI2BB2XL U8091 ( .B0(\D_cache/n421 ), .B1(n3849), .A0N(
        \D_cache/cache[4][46] ), .A1N(n3859), .Y(\D_cache/n1424 ) );
  OAI2BB2XL U8092 ( .B0(\D_cache/n421 ), .B1(n3868), .A0N(
        \D_cache/cache[3][46] ), .A1N(n3878), .Y(\D_cache/n1425 ) );
  OAI2BB2XL U8093 ( .B0(\D_cache/n421 ), .B1(n3891), .A0N(
        \D_cache/cache[2][46] ), .A1N(n3899), .Y(\D_cache/n1426 ) );
  OAI2BB2XL U8094 ( .B0(\D_cache/n421 ), .B1(n3911), .A0N(
        \D_cache/cache[1][46] ), .A1N(n3920), .Y(\D_cache/n1427 ) );
  OAI2BB2XL U8095 ( .B0(\D_cache/n421 ), .B1(n3931), .A0N(
        \D_cache/cache[0][46] ), .A1N(n3941), .Y(\D_cache/n1428 ) );
  OAI2BB2XL U8096 ( .B0(\D_cache/n425 ), .B1(n3791), .A0N(
        \D_cache/cache[7][44] ), .A1N(n3799), .Y(\D_cache/n1437 ) );
  OAI2BB2XL U8097 ( .B0(\D_cache/n425 ), .B1(n3811), .A0N(
        \D_cache/cache[6][44] ), .A1N(n3819), .Y(\D_cache/n1438 ) );
  OAI2BB2XL U8098 ( .B0(\D_cache/n425 ), .B1(n3829), .A0N(
        \D_cache/cache[5][44] ), .A1N(n3837), .Y(\D_cache/n1439 ) );
  OAI2BB2XL U8099 ( .B0(\D_cache/n425 ), .B1(n3849), .A0N(
        \D_cache/cache[4][44] ), .A1N(n3859), .Y(\D_cache/n1440 ) );
  OAI2BB2XL U8100 ( .B0(\D_cache/n425 ), .B1(n3868), .A0N(
        \D_cache/cache[3][44] ), .A1N(n3878), .Y(\D_cache/n1441 ) );
  OAI2BB2XL U8101 ( .B0(\D_cache/n425 ), .B1(n3891), .A0N(
        \D_cache/cache[2][44] ), .A1N(n3899), .Y(\D_cache/n1442 ) );
  OAI2BB2XL U8102 ( .B0(\D_cache/n425 ), .B1(n3911), .A0N(
        \D_cache/cache[1][44] ), .A1N(n3920), .Y(\D_cache/n1443 ) );
  OAI2BB2XL U8103 ( .B0(\D_cache/n425 ), .B1(n3931), .A0N(
        \D_cache/cache[0][44] ), .A1N(n3941), .Y(\D_cache/n1444 ) );
  OAI2BB2XL U8104 ( .B0(\D_cache/n429 ), .B1(n3793), .A0N(
        \D_cache/cache[7][42] ), .A1N(n3799), .Y(\D_cache/n1453 ) );
  OAI2BB2XL U8105 ( .B0(\D_cache/n429 ), .B1(n3813), .A0N(
        \D_cache/cache[6][42] ), .A1N(n3819), .Y(\D_cache/n1454 ) );
  OAI2BB2XL U8106 ( .B0(\D_cache/n429 ), .B1(n3831), .A0N(
        \D_cache/cache[5][42] ), .A1N(n3837), .Y(\D_cache/n1455 ) );
  OAI2BB2XL U8107 ( .B0(\D_cache/n429 ), .B1(n3853), .A0N(
        \D_cache/cache[4][42] ), .A1N(n3859), .Y(\D_cache/n1456 ) );
  OAI2BB2XL U8108 ( .B0(\D_cache/n429 ), .B1(n3872), .A0N(
        \D_cache/cache[3][42] ), .A1N(n3878), .Y(\D_cache/n1457 ) );
  OAI2BB2XL U8109 ( .B0(\D_cache/n429 ), .B1(n3893), .A0N(
        \D_cache/cache[2][42] ), .A1N(n3899), .Y(\D_cache/n1458 ) );
  OAI2BB2XL U8110 ( .B0(\D_cache/n429 ), .B1(n3914), .A0N(
        \D_cache/cache[1][42] ), .A1N(n3920), .Y(\D_cache/n1459 ) );
  OAI2BB2XL U8111 ( .B0(\D_cache/n429 ), .B1(n3935), .A0N(
        \D_cache/cache[0][42] ), .A1N(n3941), .Y(\D_cache/n1460 ) );
  OAI2BB2XL U8112 ( .B0(\D_cache/n431 ), .B1(n3794), .A0N(
        \D_cache/cache[7][41] ), .A1N(n3799), .Y(\D_cache/n1461 ) );
  OAI2BB2XL U8113 ( .B0(\D_cache/n431 ), .B1(n3814), .A0N(
        \D_cache/cache[6][41] ), .A1N(n3819), .Y(\D_cache/n1462 ) );
  OAI2BB2XL U8114 ( .B0(\D_cache/n431 ), .B1(n3832), .A0N(
        \D_cache/cache[5][41] ), .A1N(n3837), .Y(\D_cache/n1463 ) );
  OAI2BB2XL U8115 ( .B0(\D_cache/n431 ), .B1(n3854), .A0N(
        \D_cache/cache[4][41] ), .A1N(n3859), .Y(\D_cache/n1464 ) );
  OAI2BB2XL U8116 ( .B0(\D_cache/n431 ), .B1(n3873), .A0N(
        \D_cache/cache[3][41] ), .A1N(n3878), .Y(\D_cache/n1465 ) );
  OAI2BB2XL U8117 ( .B0(\D_cache/n431 ), .B1(n3894), .A0N(
        \D_cache/cache[2][41] ), .A1N(n3899), .Y(\D_cache/n1466 ) );
  OAI2BB2XL U8118 ( .B0(\D_cache/n431 ), .B1(n3915), .A0N(
        \D_cache/cache[1][41] ), .A1N(n3920), .Y(\D_cache/n1467 ) );
  OAI2BB2XL U8119 ( .B0(\D_cache/n431 ), .B1(n3936), .A0N(
        \D_cache/cache[0][41] ), .A1N(n3941), .Y(\D_cache/n1468 ) );
  OAI2BB2XL U8120 ( .B0(\D_cache/n433 ), .B1(n3794), .A0N(
        \D_cache/cache[7][40] ), .A1N(n3799), .Y(\D_cache/n1469 ) );
  OAI2BB2XL U8121 ( .B0(\D_cache/n433 ), .B1(n3814), .A0N(
        \D_cache/cache[6][40] ), .A1N(n3819), .Y(\D_cache/n1470 ) );
  OAI2BB2XL U8122 ( .B0(\D_cache/n433 ), .B1(n3832), .A0N(
        \D_cache/cache[5][40] ), .A1N(n3837), .Y(\D_cache/n1471 ) );
  OAI2BB2XL U8123 ( .B0(\D_cache/n433 ), .B1(n3854), .A0N(
        \D_cache/cache[4][40] ), .A1N(n3859), .Y(\D_cache/n1472 ) );
  OAI2BB2XL U8124 ( .B0(\D_cache/n433 ), .B1(n3873), .A0N(
        \D_cache/cache[3][40] ), .A1N(n3878), .Y(\D_cache/n1473 ) );
  OAI2BB2XL U8125 ( .B0(\D_cache/n433 ), .B1(n3894), .A0N(
        \D_cache/cache[2][40] ), .A1N(n3899), .Y(\D_cache/n1474 ) );
  OAI2BB2XL U8126 ( .B0(\D_cache/n433 ), .B1(n3915), .A0N(
        \D_cache/cache[1][40] ), .A1N(n3920), .Y(\D_cache/n1475 ) );
  OAI2BB2XL U8127 ( .B0(\D_cache/n433 ), .B1(n3936), .A0N(
        \D_cache/cache[0][40] ), .A1N(n3941), .Y(\D_cache/n1476 ) );
  OAI2BB2XL U8128 ( .B0(\D_cache/n435 ), .B1(n3794), .A0N(
        \D_cache/cache[7][39] ), .A1N(n3799), .Y(\D_cache/n1477 ) );
  OAI2BB2XL U8129 ( .B0(\D_cache/n435 ), .B1(n3814), .A0N(
        \D_cache/cache[6][39] ), .A1N(n3819), .Y(\D_cache/n1478 ) );
  OAI2BB2XL U8130 ( .B0(\D_cache/n435 ), .B1(n3832), .A0N(
        \D_cache/cache[5][39] ), .A1N(n3837), .Y(\D_cache/n1479 ) );
  OAI2BB2XL U8131 ( .B0(\D_cache/n435 ), .B1(n3854), .A0N(
        \D_cache/cache[4][39] ), .A1N(n3859), .Y(\D_cache/n1480 ) );
  OAI2BB2XL U8132 ( .B0(\D_cache/n435 ), .B1(n3873), .A0N(
        \D_cache/cache[3][39] ), .A1N(n3878), .Y(\D_cache/n1481 ) );
  OAI2BB2XL U8133 ( .B0(\D_cache/n435 ), .B1(n3894), .A0N(
        \D_cache/cache[2][39] ), .A1N(n3899), .Y(\D_cache/n1482 ) );
  OAI2BB2XL U8134 ( .B0(\D_cache/n435 ), .B1(n3915), .A0N(
        \D_cache/cache[1][39] ), .A1N(n3920), .Y(\D_cache/n1483 ) );
  OAI2BB2XL U8135 ( .B0(\D_cache/n435 ), .B1(n3936), .A0N(
        \D_cache/cache[0][39] ), .A1N(n3941), .Y(\D_cache/n1484 ) );
  OAI2BB2XL U8136 ( .B0(\D_cache/n437 ), .B1(n3793), .A0N(
        \D_cache/cache[7][38] ), .A1N(n3799), .Y(\D_cache/n1485 ) );
  OAI2BB2XL U8137 ( .B0(\D_cache/n437 ), .B1(n3813), .A0N(
        \D_cache/cache[6][38] ), .A1N(n3819), .Y(\D_cache/n1486 ) );
  OAI2BB2XL U8138 ( .B0(\D_cache/n437 ), .B1(n3831), .A0N(
        \D_cache/cache[5][38] ), .A1N(n3837), .Y(\D_cache/n1487 ) );
  OAI2BB2XL U8139 ( .B0(\D_cache/n437 ), .B1(n3853), .A0N(
        \D_cache/cache[4][38] ), .A1N(n3859), .Y(\D_cache/n1488 ) );
  OAI2BB2XL U8140 ( .B0(\D_cache/n437 ), .B1(n3872), .A0N(
        \D_cache/cache[3][38] ), .A1N(n3878), .Y(\D_cache/n1489 ) );
  OAI2BB2XL U8141 ( .B0(\D_cache/n437 ), .B1(n3893), .A0N(
        \D_cache/cache[2][38] ), .A1N(n3899), .Y(\D_cache/n1490 ) );
  OAI2BB2XL U8142 ( .B0(\D_cache/n437 ), .B1(n3914), .A0N(
        \D_cache/cache[1][38] ), .A1N(n3920), .Y(\D_cache/n1491 ) );
  OAI2BB2XL U8143 ( .B0(\D_cache/n437 ), .B1(n3935), .A0N(
        \D_cache/cache[0][38] ), .A1N(n3941), .Y(\D_cache/n1492 ) );
  OAI2BB2XL U8144 ( .B0(\D_cache/n439 ), .B1(n3793), .A0N(
        \D_cache/cache[7][37] ), .A1N(n3799), .Y(\D_cache/n1493 ) );
  OAI2BB2XL U8145 ( .B0(\D_cache/n439 ), .B1(n3813), .A0N(
        \D_cache/cache[6][37] ), .A1N(n3819), .Y(\D_cache/n1494 ) );
  OAI2BB2XL U8146 ( .B0(\D_cache/n439 ), .B1(n3831), .A0N(
        \D_cache/cache[5][37] ), .A1N(n3837), .Y(\D_cache/n1495 ) );
  OAI2BB2XL U8147 ( .B0(\D_cache/n439 ), .B1(n3853), .A0N(
        \D_cache/cache[4][37] ), .A1N(n3859), .Y(\D_cache/n1496 ) );
  OAI2BB2XL U8148 ( .B0(\D_cache/n439 ), .B1(n3872), .A0N(
        \D_cache/cache[3][37] ), .A1N(n3878), .Y(\D_cache/n1497 ) );
  OAI2BB2XL U8149 ( .B0(\D_cache/n439 ), .B1(n3893), .A0N(
        \D_cache/cache[2][37] ), .A1N(n3899), .Y(\D_cache/n1498 ) );
  OAI2BB2XL U8150 ( .B0(\D_cache/n439 ), .B1(n3914), .A0N(
        \D_cache/cache[1][37] ), .A1N(n3920), .Y(\D_cache/n1499 ) );
  OAI2BB2XL U8151 ( .B0(\D_cache/n439 ), .B1(n3935), .A0N(
        \D_cache/cache[0][37] ), .A1N(n3941), .Y(\D_cache/n1500 ) );
  OAI2BB2XL U8152 ( .B0(\D_cache/n449 ), .B1(n3793), .A0N(
        \D_cache/cache[7][32] ), .A1N(n3799), .Y(\D_cache/n1533 ) );
  OAI2BB2XL U8153 ( .B0(\D_cache/n449 ), .B1(n3813), .A0N(
        \D_cache/cache[6][32] ), .A1N(n3819), .Y(\D_cache/n1534 ) );
  OAI2BB2XL U8154 ( .B0(\D_cache/n449 ), .B1(n3831), .A0N(
        \D_cache/cache[5][32] ), .A1N(n3837), .Y(\D_cache/n1535 ) );
  OAI2BB2XL U8155 ( .B0(\D_cache/n449 ), .B1(n3853), .A0N(
        \D_cache/cache[4][32] ), .A1N(n3859), .Y(\D_cache/n1536 ) );
  OAI2BB2XL U8156 ( .B0(\D_cache/n449 ), .B1(n3872), .A0N(
        \D_cache/cache[3][32] ), .A1N(n3878), .Y(\D_cache/n1537 ) );
  OAI2BB2XL U8157 ( .B0(\D_cache/n449 ), .B1(n3893), .A0N(
        \D_cache/cache[2][32] ), .A1N(n3899), .Y(\D_cache/n1538 ) );
  OAI2BB2XL U8158 ( .B0(\D_cache/n449 ), .B1(n3914), .A0N(
        \D_cache/cache[1][32] ), .A1N(n3920), .Y(\D_cache/n1539 ) );
  OAI2BB2XL U8159 ( .B0(\D_cache/n449 ), .B1(n3935), .A0N(
        \D_cache/cache[0][32] ), .A1N(n3941), .Y(\D_cache/n1540 ) );
  OAI2BB2XL U8160 ( .B0(\D_cache/n385 ), .B1(n3788), .A0N(
        \D_cache/cache[7][63] ), .A1N(n3800), .Y(\D_cache/n1285 ) );
  OAI2BB2XL U8161 ( .B0(\D_cache/n385 ), .B1(n3808), .A0N(
        \D_cache/cache[6][63] ), .A1N(n3820), .Y(\D_cache/n1286 ) );
  OAI2BB2XL U8162 ( .B0(\D_cache/n385 ), .B1(n3827), .A0N(
        \D_cache/cache[5][63] ), .A1N(n3831), .Y(\D_cache/n1287 ) );
  OAI2BB2XL U8163 ( .B0(\D_cache/n385 ), .B1(n3846), .A0N(
        \D_cache/cache[4][63] ), .A1N(n3860), .Y(\D_cache/n1288 ) );
  OAI2BB2XL U8164 ( .B0(\D_cache/n385 ), .B1(n3880), .A0N(
        \D_cache/cache[3][63] ), .A1N(n3879), .Y(\D_cache/n1289 ) );
  OAI2BB2XL U8165 ( .B0(\D_cache/n385 ), .B1(n3888), .A0N(
        \D_cache/cache[2][63] ), .A1N(n3900), .Y(\D_cache/n1290 ) );
  OAI2BB2XL U8166 ( .B0(\D_cache/n385 ), .B1(n3908), .A0N(
        \D_cache/cache[1][63] ), .A1N(n3921), .Y(\D_cache/n1291 ) );
  OAI2BB2XL U8167 ( .B0(\D_cache/n385 ), .B1(n3928), .A0N(
        \D_cache/cache[0][63] ), .A1N(n3942), .Y(\D_cache/n1292 ) );
  OAI2BB2XL U8168 ( .B0(\D_cache/n391 ), .B1(n3789), .A0N(
        \D_cache/cache[7][61] ), .A1N(n3800), .Y(\D_cache/n1301 ) );
  OAI2BB2XL U8169 ( .B0(\D_cache/n391 ), .B1(n3809), .A0N(
        \D_cache/cache[6][61] ), .A1N(n3820), .Y(\D_cache/n1302 ) );
  OAI2BB2XL U8170 ( .B0(\D_cache/n391 ), .B1(n3828), .A0N(
        \D_cache/cache[5][61] ), .A1N(n3826), .Y(\D_cache/n1303 ) );
  OAI2BB2XL U8171 ( .B0(\D_cache/n391 ), .B1(n3847), .A0N(
        \D_cache/cache[4][61] ), .A1N(n3860), .Y(\D_cache/n1304 ) );
  OAI2BB2XL U8172 ( .B0(\D_cache/n391 ), .B1(n3866), .A0N(
        \D_cache/cache[3][61] ), .A1N(n3879), .Y(\D_cache/n1305 ) );
  OAI2BB2XL U8173 ( .B0(\D_cache/n391 ), .B1(n3889), .A0N(
        \D_cache/cache[2][61] ), .A1N(n3900), .Y(\D_cache/n1306 ) );
  OAI2BB2XL U8174 ( .B0(\D_cache/n391 ), .B1(n3909), .A0N(
        \D_cache/cache[1][61] ), .A1N(n3921), .Y(\D_cache/n1307 ) );
  OAI2BB2XL U8175 ( .B0(\D_cache/n391 ), .B1(n3929), .A0N(
        \D_cache/cache[0][61] ), .A1N(n3942), .Y(\D_cache/n1308 ) );
  OAI2BB2XL U8176 ( .B0(\D_cache/n399 ), .B1(n3789), .A0N(
        \D_cache/cache[7][57] ), .A1N(n3800), .Y(\D_cache/n1333 ) );
  OAI2BB2XL U8177 ( .B0(\D_cache/n399 ), .B1(n3809), .A0N(
        \D_cache/cache[6][57] ), .A1N(n3820), .Y(\D_cache/n1334 ) );
  OAI2BB2XL U8178 ( .B0(\D_cache/n399 ), .B1(n3828), .A0N(
        \D_cache/cache[5][57] ), .A1N(n3830), .Y(\D_cache/n1335 ) );
  OAI2BB2XL U8179 ( .B0(\D_cache/n399 ), .B1(n3847), .A0N(
        \D_cache/cache[4][57] ), .A1N(n3860), .Y(\D_cache/n1336 ) );
  OAI2BB2XL U8180 ( .B0(\D_cache/n399 ), .B1(n3866), .A0N(
        \D_cache/cache[3][57] ), .A1N(n3879), .Y(\D_cache/n1337 ) );
  OAI2BB2XL U8181 ( .B0(\D_cache/n399 ), .B1(n3889), .A0N(
        \D_cache/cache[2][57] ), .A1N(n3900), .Y(\D_cache/n1338 ) );
  OAI2BB2XL U8182 ( .B0(\D_cache/n399 ), .B1(n3909), .A0N(
        \D_cache/cache[1][57] ), .A1N(n3921), .Y(\D_cache/n1339 ) );
  OAI2BB2XL U8183 ( .B0(\D_cache/n399 ), .B1(n3929), .A0N(
        \D_cache/cache[0][57] ), .A1N(n3942), .Y(\D_cache/n1340 ) );
  OAI2BB2XL U8184 ( .B0(\D_cache/n401 ), .B1(n3789), .A0N(
        \D_cache/cache[7][56] ), .A1N(n3800), .Y(\D_cache/n1341 ) );
  OAI2BB2XL U8185 ( .B0(\D_cache/n401 ), .B1(n3809), .A0N(
        \D_cache/cache[6][56] ), .A1N(n3820), .Y(\D_cache/n1342 ) );
  OAI2BB2XL U8186 ( .B0(\D_cache/n401 ), .B1(n3828), .A0N(
        \D_cache/cache[5][56] ), .A1N(n3824), .Y(\D_cache/n1343 ) );
  OAI2BB2XL U8187 ( .B0(\D_cache/n401 ), .B1(n3847), .A0N(
        \D_cache/cache[4][56] ), .A1N(n3860), .Y(\D_cache/n1344 ) );
  OAI2BB2XL U8188 ( .B0(\D_cache/n401 ), .B1(n3866), .A0N(
        \D_cache/cache[3][56] ), .A1N(n3879), .Y(\D_cache/n1345 ) );
  OAI2BB2XL U8189 ( .B0(\D_cache/n401 ), .B1(n3889), .A0N(
        \D_cache/cache[2][56] ), .A1N(n3900), .Y(\D_cache/n1346 ) );
  OAI2BB2XL U8190 ( .B0(\D_cache/n401 ), .B1(n3909), .A0N(
        \D_cache/cache[1][56] ), .A1N(n3921), .Y(\D_cache/n1347 ) );
  OAI2BB2XL U8191 ( .B0(\D_cache/n401 ), .B1(n3929), .A0N(
        \D_cache/cache[0][56] ), .A1N(n3942), .Y(\D_cache/n1348 ) );
  OAI2BB2XL U8192 ( .B0(\D_cache/n407 ), .B1(n3790), .A0N(
        \D_cache/cache[7][53] ), .A1N(n3800), .Y(\D_cache/n1365 ) );
  OAI2BB2XL U8193 ( .B0(\D_cache/n407 ), .B1(n3810), .A0N(
        \D_cache/cache[6][53] ), .A1N(n3820), .Y(\D_cache/n1366 ) );
  OAI2BB2XL U8194 ( .B0(\D_cache/n407 ), .B1(n3831), .A0N(
        \D_cache/cache[5][53] ), .A1N(n3832), .Y(\D_cache/n1367 ) );
  OAI2BB2XL U8195 ( .B0(\D_cache/n407 ), .B1(n3848), .A0N(
        \D_cache/cache[4][53] ), .A1N(n3860), .Y(\D_cache/n1368 ) );
  OAI2BB2XL U8196 ( .B0(\D_cache/n407 ), .B1(n3867), .A0N(
        \D_cache/cache[3][53] ), .A1N(n3879), .Y(\D_cache/n1369 ) );
  OAI2BB2XL U8197 ( .B0(\D_cache/n407 ), .B1(n3890), .A0N(
        \D_cache/cache[2][53] ), .A1N(n3900), .Y(\D_cache/n1370 ) );
  OAI2BB2XL U8198 ( .B0(\D_cache/n407 ), .B1(n3910), .A0N(
        \D_cache/cache[1][53] ), .A1N(n3921), .Y(\D_cache/n1371 ) );
  OAI2BB2XL U8199 ( .B0(\D_cache/n407 ), .B1(n3930), .A0N(
        \D_cache/cache[0][53] ), .A1N(n3942), .Y(\D_cache/n1372 ) );
  OAI2BB2XL U8200 ( .B0(\D_cache/n409 ), .B1(n3790), .A0N(
        \D_cache/cache[7][52] ), .A1N(n3800), .Y(\D_cache/n1373 ) );
  OAI2BB2XL U8201 ( .B0(\D_cache/n409 ), .B1(n3810), .A0N(
        \D_cache/cache[6][52] ), .A1N(n3820), .Y(\D_cache/n1374 ) );
  OAI2BB2XL U8202 ( .B0(\D_cache/n409 ), .B1(n3825), .A0N(
        \D_cache/cache[5][52] ), .A1N(n3838), .Y(\D_cache/n1375 ) );
  OAI2BB2XL U8203 ( .B0(\D_cache/n409 ), .B1(n3848), .A0N(
        \D_cache/cache[4][52] ), .A1N(n3860), .Y(\D_cache/n1376 ) );
  OAI2BB2XL U8204 ( .B0(\D_cache/n409 ), .B1(n3867), .A0N(
        \D_cache/cache[3][52] ), .A1N(n3879), .Y(\D_cache/n1377 ) );
  OAI2BB2XL U8205 ( .B0(\D_cache/n409 ), .B1(n3890), .A0N(
        \D_cache/cache[2][52] ), .A1N(n3900), .Y(\D_cache/n1378 ) );
  OAI2BB2XL U8206 ( .B0(\D_cache/n409 ), .B1(n3910), .A0N(
        \D_cache/cache[1][52] ), .A1N(n3921), .Y(\D_cache/n1379 ) );
  OAI2BB2XL U8207 ( .B0(\D_cache/n409 ), .B1(n3930), .A0N(
        \D_cache/cache[0][52] ), .A1N(n3942), .Y(\D_cache/n1380 ) );
  OAI2BB2XL U8208 ( .B0(\D_cache/n441 ), .B1(n3794), .A0N(
        \D_cache/cache[7][36] ), .A1N(n3799), .Y(\D_cache/n1501 ) );
  OAI2BB2XL U8209 ( .B0(\D_cache/n441 ), .B1(n3814), .A0N(
        \D_cache/cache[6][36] ), .A1N(n3819), .Y(\D_cache/n1502 ) );
  OAI2BB2XL U8210 ( .B0(\D_cache/n441 ), .B1(n3832), .A0N(
        \D_cache/cache[5][36] ), .A1N(n3837), .Y(\D_cache/n1503 ) );
  OAI2BB2XL U8211 ( .B0(\D_cache/n441 ), .B1(n3854), .A0N(
        \D_cache/cache[4][36] ), .A1N(n3859), .Y(\D_cache/n1504 ) );
  OAI2BB2XL U8212 ( .B0(\D_cache/n441 ), .B1(n3873), .A0N(
        \D_cache/cache[3][36] ), .A1N(n3878), .Y(\D_cache/n1505 ) );
  OAI2BB2XL U8213 ( .B0(\D_cache/n441 ), .B1(n3894), .A0N(
        \D_cache/cache[2][36] ), .A1N(n3899), .Y(\D_cache/n1506 ) );
  OAI2BB2XL U8214 ( .B0(\D_cache/n441 ), .B1(n3915), .A0N(
        \D_cache/cache[1][36] ), .A1N(n3920), .Y(\D_cache/n1507 ) );
  OAI2BB2XL U8215 ( .B0(\D_cache/n441 ), .B1(n3936), .A0N(
        \D_cache/cache[0][36] ), .A1N(n3941), .Y(\D_cache/n1508 ) );
  OAI2BB2XL U8216 ( .B0(\D_cache/n443 ), .B1(n3794), .A0N(
        \D_cache/cache[7][35] ), .A1N(n3799), .Y(\D_cache/n1509 ) );
  OAI2BB2XL U8217 ( .B0(\D_cache/n443 ), .B1(n3814), .A0N(
        \D_cache/cache[6][35] ), .A1N(n3819), .Y(\D_cache/n1510 ) );
  OAI2BB2XL U8218 ( .B0(\D_cache/n443 ), .B1(n3832), .A0N(
        \D_cache/cache[5][35] ), .A1N(n3837), .Y(\D_cache/n1511 ) );
  OAI2BB2XL U8219 ( .B0(\D_cache/n443 ), .B1(n3854), .A0N(
        \D_cache/cache[4][35] ), .A1N(n3859), .Y(\D_cache/n1512 ) );
  OAI2BB2XL U8220 ( .B0(\D_cache/n443 ), .B1(n3873), .A0N(
        \D_cache/cache[3][35] ), .A1N(n3878), .Y(\D_cache/n1513 ) );
  OAI2BB2XL U8221 ( .B0(\D_cache/n443 ), .B1(n3894), .A0N(
        \D_cache/cache[2][35] ), .A1N(n3899), .Y(\D_cache/n1514 ) );
  OAI2BB2XL U8222 ( .B0(\D_cache/n443 ), .B1(n3915), .A0N(
        \D_cache/cache[1][35] ), .A1N(n3920), .Y(\D_cache/n1515 ) );
  OAI2BB2XL U8223 ( .B0(\D_cache/n443 ), .B1(n3936), .A0N(
        \D_cache/cache[0][35] ), .A1N(n3941), .Y(\D_cache/n1516 ) );
  OAI2BB2XL U8224 ( .B0(\D_cache/n445 ), .B1(n3794), .A0N(
        \D_cache/cache[7][34] ), .A1N(n3799), .Y(\D_cache/n1517 ) );
  OAI2BB2XL U8225 ( .B0(\D_cache/n445 ), .B1(n3814), .A0N(
        \D_cache/cache[6][34] ), .A1N(n3819), .Y(\D_cache/n1518 ) );
  OAI2BB2XL U8226 ( .B0(\D_cache/n445 ), .B1(n3832), .A0N(
        \D_cache/cache[5][34] ), .A1N(n3837), .Y(\D_cache/n1519 ) );
  OAI2BB2XL U8227 ( .B0(\D_cache/n445 ), .B1(n3854), .A0N(
        \D_cache/cache[4][34] ), .A1N(n3859), .Y(\D_cache/n1520 ) );
  OAI2BB2XL U8228 ( .B0(\D_cache/n445 ), .B1(n3873), .A0N(
        \D_cache/cache[3][34] ), .A1N(n3878), .Y(\D_cache/n1521 ) );
  OAI2BB2XL U8229 ( .B0(\D_cache/n445 ), .B1(n3894), .A0N(
        \D_cache/cache[2][34] ), .A1N(n3899), .Y(\D_cache/n1522 ) );
  OAI2BB2XL U8230 ( .B0(\D_cache/n445 ), .B1(n3915), .A0N(
        \D_cache/cache[1][34] ), .A1N(n3920), .Y(\D_cache/n1523 ) );
  OAI2BB2XL U8231 ( .B0(\D_cache/n445 ), .B1(n3936), .A0N(
        \D_cache/cache[0][34] ), .A1N(n3941), .Y(\D_cache/n1524 ) );
  OAI2BB2XL U8232 ( .B0(\D_cache/n447 ), .B1(n3794), .A0N(
        \D_cache/cache[7][33] ), .A1N(n3799), .Y(\D_cache/n1525 ) );
  OAI2BB2XL U8233 ( .B0(\D_cache/n447 ), .B1(n3814), .A0N(
        \D_cache/cache[6][33] ), .A1N(n3819), .Y(\D_cache/n1526 ) );
  OAI2BB2XL U8234 ( .B0(\D_cache/n447 ), .B1(n3832), .A0N(
        \D_cache/cache[5][33] ), .A1N(n3837), .Y(\D_cache/n1527 ) );
  OAI2BB2XL U8235 ( .B0(\D_cache/n447 ), .B1(n3854), .A0N(
        \D_cache/cache[4][33] ), .A1N(n3859), .Y(\D_cache/n1528 ) );
  OAI2BB2XL U8236 ( .B0(\D_cache/n447 ), .B1(n3873), .A0N(
        \D_cache/cache[3][33] ), .A1N(n3878), .Y(\D_cache/n1529 ) );
  OAI2BB2XL U8237 ( .B0(\D_cache/n447 ), .B1(n3894), .A0N(
        \D_cache/cache[2][33] ), .A1N(n3899), .Y(\D_cache/n1530 ) );
  OAI2BB2XL U8238 ( .B0(\D_cache/n447 ), .B1(n3915), .A0N(
        \D_cache/cache[1][33] ), .A1N(n3920), .Y(\D_cache/n1531 ) );
  OAI2BB2XL U8239 ( .B0(\D_cache/n447 ), .B1(n3936), .A0N(
        \D_cache/cache[0][33] ), .A1N(n3941), .Y(\D_cache/n1532 ) );
  OAI2BB2XL U8240 ( .B0(\D_cache/n397 ), .B1(n3789), .A0N(
        \D_cache/cache[7][58] ), .A1N(n3800), .Y(\D_cache/n1325 ) );
  OAI2BB2XL U8241 ( .B0(\D_cache/n397 ), .B1(n3809), .A0N(
        \D_cache/cache[6][58] ), .A1N(n3820), .Y(\D_cache/n1326 ) );
  OAI2BB2XL U8242 ( .B0(\D_cache/n397 ), .B1(n3828), .A0N(
        \D_cache/cache[5][58] ), .A1N(n3829), .Y(\D_cache/n1327 ) );
  OAI2BB2XL U8243 ( .B0(\D_cache/n397 ), .B1(n3847), .A0N(
        \D_cache/cache[4][58] ), .A1N(n3860), .Y(\D_cache/n1328 ) );
  OAI2BB2XL U8244 ( .B0(\D_cache/n397 ), .B1(n3866), .A0N(
        \D_cache/cache[3][58] ), .A1N(n3879), .Y(\D_cache/n1329 ) );
  OAI2BB2XL U8245 ( .B0(\D_cache/n397 ), .B1(n3889), .A0N(
        \D_cache/cache[2][58] ), .A1N(n3900), .Y(\D_cache/n1330 ) );
  OAI2BB2XL U8246 ( .B0(\D_cache/n397 ), .B1(n3909), .A0N(
        \D_cache/cache[1][58] ), .A1N(n3921), .Y(\D_cache/n1331 ) );
  OAI2BB2XL U8247 ( .B0(\D_cache/n397 ), .B1(n3929), .A0N(
        \D_cache/cache[0][58] ), .A1N(n3942), .Y(\D_cache/n1332 ) );
  OAI2BB2XL U8248 ( .B0(\D_cache/n413 ), .B1(n3790), .A0N(
        \D_cache/cache[7][50] ), .A1N(n3800), .Y(\D_cache/n1389 ) );
  OAI2BB2XL U8249 ( .B0(\D_cache/n413 ), .B1(n3810), .A0N(
        \D_cache/cache[6][50] ), .A1N(n3820), .Y(\D_cache/n1390 ) );
  OAI2BB2XL U8250 ( .B0(\D_cache/n413 ), .B1(n3826), .A0N(
        \D_cache/cache[5][50] ), .A1N(n3828), .Y(\D_cache/n1391 ) );
  OAI2BB2XL U8251 ( .B0(\D_cache/n413 ), .B1(n3848), .A0N(
        \D_cache/cache[4][50] ), .A1N(n3860), .Y(\D_cache/n1392 ) );
  OAI2BB2XL U8252 ( .B0(\D_cache/n413 ), .B1(n3867), .A0N(
        \D_cache/cache[3][50] ), .A1N(n3879), .Y(\D_cache/n1393 ) );
  OAI2BB2XL U8253 ( .B0(\D_cache/n413 ), .B1(n3890), .A0N(
        \D_cache/cache[2][50] ), .A1N(n3900), .Y(\D_cache/n1394 ) );
  OAI2BB2XL U8254 ( .B0(\D_cache/n413 ), .B1(n3910), .A0N(
        \D_cache/cache[1][50] ), .A1N(n3921), .Y(\D_cache/n1395 ) );
  OAI2BB2XL U8255 ( .B0(\D_cache/n413 ), .B1(n3930), .A0N(
        \D_cache/cache[0][50] ), .A1N(n3942), .Y(\D_cache/n1396 ) );
  OAI2BB2XL U8256 ( .B0(\D_cache/n415 ), .B1(n3790), .A0N(
        \D_cache/cache[7][49] ), .A1N(n3800), .Y(\D_cache/n1397 ) );
  OAI2BB2XL U8257 ( .B0(\D_cache/n415 ), .B1(n3810), .A0N(
        \D_cache/cache[6][49] ), .A1N(n3820), .Y(\D_cache/n1398 ) );
  OAI2BB2XL U8258 ( .B0(\D_cache/n415 ), .B1(n3829), .A0N(
        \D_cache/cache[5][49] ), .A1N(n3825), .Y(\D_cache/n1399 ) );
  OAI2BB2XL U8259 ( .B0(\D_cache/n415 ), .B1(n3848), .A0N(
        \D_cache/cache[4][49] ), .A1N(n3860), .Y(\D_cache/n1400 ) );
  OAI2BB2XL U8260 ( .B0(\D_cache/n415 ), .B1(n3867), .A0N(
        \D_cache/cache[3][49] ), .A1N(n3879), .Y(\D_cache/n1401 ) );
  OAI2BB2XL U8261 ( .B0(\D_cache/n415 ), .B1(n3890), .A0N(
        \D_cache/cache[2][49] ), .A1N(n3900), .Y(\D_cache/n1402 ) );
  OAI2BB2XL U8262 ( .B0(\D_cache/n415 ), .B1(n3910), .A0N(
        \D_cache/cache[1][49] ), .A1N(n3921), .Y(\D_cache/n1403 ) );
  OAI2BB2XL U8263 ( .B0(\D_cache/n415 ), .B1(n3930), .A0N(
        \D_cache/cache[0][49] ), .A1N(n3942), .Y(\D_cache/n1404 ) );
  OAI2BB2XL U8264 ( .B0(\D_cache/n411 ), .B1(n3790), .A0N(
        \D_cache/cache[7][51] ), .A1N(n3800), .Y(\D_cache/n1381 ) );
  OAI2BB2XL U8265 ( .B0(\D_cache/n411 ), .B1(n3810), .A0N(
        \D_cache/cache[6][51] ), .A1N(n3820), .Y(\D_cache/n1382 ) );
  OAI2BB2XL U8266 ( .B0(\D_cache/n411 ), .B1(n3828), .A0N(
        \D_cache/cache[5][51] ), .A1N(n3839), .Y(\D_cache/n1383 ) );
  OAI2BB2XL U8267 ( .B0(\D_cache/n411 ), .B1(n3848), .A0N(
        \D_cache/cache[4][51] ), .A1N(n3860), .Y(\D_cache/n1384 ) );
  OAI2BB2XL U8268 ( .B0(\D_cache/n411 ), .B1(n3867), .A0N(
        \D_cache/cache[3][51] ), .A1N(n3879), .Y(\D_cache/n1385 ) );
  OAI2BB2XL U8269 ( .B0(\D_cache/n411 ), .B1(n3890), .A0N(
        \D_cache/cache[2][51] ), .A1N(n3900), .Y(\D_cache/n1386 ) );
  OAI2BB2XL U8270 ( .B0(\D_cache/n411 ), .B1(n3910), .A0N(
        \D_cache/cache[1][51] ), .A1N(n3921), .Y(\D_cache/n1387 ) );
  OAI2BB2XL U8271 ( .B0(\D_cache/n411 ), .B1(n3930), .A0N(
        \D_cache/cache[0][51] ), .A1N(n3942), .Y(\D_cache/n1388 ) );
  AO21X1 U8272 ( .A0(\i_MIPS/ID_EX[80] ), .A1(\i_MIPS/ALU/N303 ), .B0(n5122), 
        .Y(n5462) );
  NAND3X4 U8273 ( .A(ICACHE_addr[16]), .B(ICACHE_addr[15]), .C(n8016), .Y(
        n8040) );
  OAI2BB2XL U8274 ( .B0(\D_cache/n248 ), .B1(n3790), .A0N(
        \D_cache/cache[7][127] ), .A1N(n3796), .Y(\D_cache/n773 ) );
  OAI2BB2XL U8275 ( .B0(\D_cache/n248 ), .B1(n3810), .A0N(
        \D_cache/cache[6][127] ), .A1N(n3816), .Y(\D_cache/n774 ) );
  OAI2BB2XL U8276 ( .B0(\D_cache/n248 ), .B1(n3827), .A0N(
        \D_cache/cache[5][127] ), .A1N(n3834), .Y(\D_cache/n775 ) );
  OAI2BB2XL U8277 ( .B0(\D_cache/n248 ), .B1(n3848), .A0N(
        \D_cache/cache[4][127] ), .A1N(n3856), .Y(\D_cache/n776 ) );
  OAI2BB2XL U8278 ( .B0(\D_cache/n248 ), .B1(n3867), .A0N(
        \D_cache/cache[3][127] ), .A1N(n3875), .Y(\D_cache/n777 ) );
  OAI2BB2XL U8279 ( .B0(\D_cache/n248 ), .B1(n3890), .A0N(
        \D_cache/cache[2][127] ), .A1N(n3896), .Y(\D_cache/n778 ) );
  OAI2BB2XL U8280 ( .B0(\D_cache/n248 ), .B1(n3910), .A0N(
        \D_cache/cache[1][127] ), .A1N(n3917), .Y(\D_cache/n779 ) );
  OAI2BB2XL U8281 ( .B0(\D_cache/n248 ), .B1(n3930), .A0N(
        \D_cache/cache[0][127] ), .A1N(n3938), .Y(\D_cache/n780 ) );
  OAI2BB2XL U8282 ( .B0(\D_cache/n252 ), .B1(n3789), .A0N(
        \D_cache/cache[7][126] ), .A1N(n3796), .Y(\D_cache/n781 ) );
  OAI2BB2XL U8283 ( .B0(\D_cache/n252 ), .B1(n3809), .A0N(
        \D_cache/cache[6][126] ), .A1N(n3816), .Y(\D_cache/n782 ) );
  OAI2BB2XL U8284 ( .B0(\D_cache/n252 ), .B1(n3828), .A0N(
        \D_cache/cache[5][126] ), .A1N(n3834), .Y(\D_cache/n783 ) );
  OAI2BB2XL U8285 ( .B0(\D_cache/n252 ), .B1(n3847), .A0N(
        \D_cache/cache[4][126] ), .A1N(n3856), .Y(\D_cache/n784 ) );
  OAI2BB2XL U8286 ( .B0(\D_cache/n252 ), .B1(n3866), .A0N(
        \D_cache/cache[3][126] ), .A1N(n3875), .Y(\D_cache/n785 ) );
  OAI2BB2XL U8287 ( .B0(\D_cache/n252 ), .B1(n3889), .A0N(
        \D_cache/cache[2][126] ), .A1N(n3896), .Y(\D_cache/n786 ) );
  OAI2BB2XL U8288 ( .B0(\D_cache/n252 ), .B1(n3909), .A0N(
        \D_cache/cache[1][126] ), .A1N(n3917), .Y(\D_cache/n787 ) );
  OAI2BB2XL U8289 ( .B0(\D_cache/n252 ), .B1(n3929), .A0N(
        \D_cache/cache[0][126] ), .A1N(n3938), .Y(\D_cache/n788 ) );
  OAI2BB2XL U8290 ( .B0(\D_cache/n254 ), .B1(n3789), .A0N(
        \D_cache/cache[7][125] ), .A1N(n3795), .Y(\D_cache/n789 ) );
  OAI2BB2XL U8291 ( .B0(\D_cache/n254 ), .B1(n3809), .A0N(
        \D_cache/cache[6][125] ), .A1N(n3815), .Y(\D_cache/n790 ) );
  OAI2BB2XL U8292 ( .B0(\D_cache/n254 ), .B1(n3828), .A0N(
        \D_cache/cache[5][125] ), .A1N(n3833), .Y(\D_cache/n791 ) );
  OAI2BB2XL U8293 ( .B0(\D_cache/n254 ), .B1(n3847), .A0N(
        \D_cache/cache[4][125] ), .A1N(n3855), .Y(\D_cache/n792 ) );
  OAI2BB2XL U8294 ( .B0(\D_cache/n254 ), .B1(n3866), .A0N(
        \D_cache/cache[3][125] ), .A1N(n3874), .Y(\D_cache/n793 ) );
  OAI2BB2XL U8295 ( .B0(\D_cache/n254 ), .B1(n3889), .A0N(
        \D_cache/cache[2][125] ), .A1N(n3895), .Y(\D_cache/n794 ) );
  OAI2BB2XL U8296 ( .B0(\D_cache/n254 ), .B1(n3909), .A0N(
        \D_cache/cache[1][125] ), .A1N(n3916), .Y(\D_cache/n795 ) );
  OAI2BB2XL U8297 ( .B0(\D_cache/n254 ), .B1(n3929), .A0N(
        \D_cache/cache[0][125] ), .A1N(n3937), .Y(\D_cache/n796 ) );
  OAI2BB2XL U8298 ( .B0(\D_cache/n256 ), .B1(n3789), .A0N(
        \D_cache/cache[7][124] ), .A1N(n3795), .Y(\D_cache/n797 ) );
  OAI2BB2XL U8299 ( .B0(\D_cache/n256 ), .B1(n3809), .A0N(
        \D_cache/cache[6][124] ), .A1N(n3815), .Y(\D_cache/n798 ) );
  OAI2BB2XL U8300 ( .B0(\D_cache/n256 ), .B1(n3828), .A0N(
        \D_cache/cache[5][124] ), .A1N(n3833), .Y(\D_cache/n799 ) );
  OAI2BB2XL U8301 ( .B0(\D_cache/n256 ), .B1(n3847), .A0N(
        \D_cache/cache[4][124] ), .A1N(n3855), .Y(\D_cache/n800 ) );
  OAI2BB2XL U8302 ( .B0(\D_cache/n256 ), .B1(n3866), .A0N(
        \D_cache/cache[3][124] ), .A1N(n3874), .Y(\D_cache/n801 ) );
  OAI2BB2XL U8303 ( .B0(\D_cache/n256 ), .B1(n3889), .A0N(
        \D_cache/cache[2][124] ), .A1N(n3895), .Y(\D_cache/n802 ) );
  OAI2BB2XL U8304 ( .B0(\D_cache/n256 ), .B1(n3909), .A0N(
        \D_cache/cache[1][124] ), .A1N(n3916), .Y(\D_cache/n803 ) );
  OAI2BB2XL U8305 ( .B0(\D_cache/n256 ), .B1(n3929), .A0N(
        \D_cache/cache[0][124] ), .A1N(n3937), .Y(\D_cache/n804 ) );
  OAI2BB2XL U8306 ( .B0(\D_cache/n258 ), .B1(n3789), .A0N(
        \D_cache/cache[7][123] ), .A1N(n3794), .Y(\D_cache/n805 ) );
  OAI2BB2XL U8307 ( .B0(\D_cache/n258 ), .B1(n3809), .A0N(
        \D_cache/cache[6][123] ), .A1N(n3814), .Y(\D_cache/n806 ) );
  OAI2BB2XL U8308 ( .B0(\D_cache/n258 ), .B1(n3828), .A0N(
        \D_cache/cache[5][123] ), .A1N(n3832), .Y(\D_cache/n807 ) );
  OAI2BB2XL U8309 ( .B0(\D_cache/n258 ), .B1(n3847), .A0N(
        \D_cache/cache[4][123] ), .A1N(n3854), .Y(\D_cache/n808 ) );
  OAI2BB2XL U8310 ( .B0(\D_cache/n258 ), .B1(n3866), .A0N(
        \D_cache/cache[3][123] ), .A1N(n3873), .Y(\D_cache/n809 ) );
  OAI2BB2XL U8311 ( .B0(\D_cache/n258 ), .B1(n3889), .A0N(
        \D_cache/cache[2][123] ), .A1N(n3894), .Y(\D_cache/n810 ) );
  OAI2BB2XL U8312 ( .B0(\D_cache/n258 ), .B1(n3909), .A0N(
        \D_cache/cache[1][123] ), .A1N(n3915), .Y(\D_cache/n811 ) );
  OAI2BB2XL U8313 ( .B0(\D_cache/n258 ), .B1(n3929), .A0N(
        \D_cache/cache[0][123] ), .A1N(n3936), .Y(\D_cache/n812 ) );
  OAI2BB2XL U8314 ( .B0(\D_cache/n260 ), .B1(n3788), .A0N(
        \D_cache/cache[7][122] ), .A1N(n3795), .Y(\D_cache/n813 ) );
  OAI2BB2XL U8315 ( .B0(\D_cache/n260 ), .B1(n3808), .A0N(
        \D_cache/cache[6][122] ), .A1N(n3815), .Y(\D_cache/n814 ) );
  OAI2BB2XL U8316 ( .B0(\D_cache/n260 ), .B1(n3827), .A0N(
        \D_cache/cache[5][122] ), .A1N(n3833), .Y(\D_cache/n815 ) );
  OAI2BB2XL U8317 ( .B0(\D_cache/n260 ), .B1(n3846), .A0N(
        \D_cache/cache[4][122] ), .A1N(n3855), .Y(\D_cache/n816 ) );
  OAI2BB2XL U8318 ( .B0(\D_cache/n260 ), .B1(n3880), .A0N(
        \D_cache/cache[3][122] ), .A1N(n3874), .Y(\D_cache/n817 ) );
  OAI2BB2XL U8319 ( .B0(\D_cache/n260 ), .B1(n3888), .A0N(
        \D_cache/cache[2][122] ), .A1N(n3895), .Y(\D_cache/n818 ) );
  OAI2BB2XL U8320 ( .B0(\D_cache/n260 ), .B1(n3908), .A0N(
        \D_cache/cache[1][122] ), .A1N(n3916), .Y(\D_cache/n819 ) );
  OAI2BB2XL U8321 ( .B0(\D_cache/n260 ), .B1(n3928), .A0N(
        \D_cache/cache[0][122] ), .A1N(n3937), .Y(\D_cache/n820 ) );
  OAI2BB2XL U8322 ( .B0(\D_cache/n262 ), .B1(n3788), .A0N(
        \D_cache/cache[7][121] ), .A1N(n3795), .Y(\D_cache/n821 ) );
  OAI2BB2XL U8323 ( .B0(\D_cache/n262 ), .B1(n3808), .A0N(
        \D_cache/cache[6][121] ), .A1N(n3815), .Y(\D_cache/n822 ) );
  OAI2BB2XL U8324 ( .B0(\D_cache/n262 ), .B1(n3827), .A0N(
        \D_cache/cache[5][121] ), .A1N(n3833), .Y(\D_cache/n823 ) );
  OAI2BB2XL U8325 ( .B0(\D_cache/n262 ), .B1(n3846), .A0N(
        \D_cache/cache[4][121] ), .A1N(n3855), .Y(\D_cache/n824 ) );
  OAI2BB2XL U8326 ( .B0(\D_cache/n262 ), .B1(n3880), .A0N(
        \D_cache/cache[3][121] ), .A1N(n3874), .Y(\D_cache/n825 ) );
  OAI2BB2XL U8327 ( .B0(\D_cache/n262 ), .B1(n3888), .A0N(
        \D_cache/cache[2][121] ), .A1N(n3895), .Y(\D_cache/n826 ) );
  OAI2BB2XL U8328 ( .B0(\D_cache/n262 ), .B1(n3908), .A0N(
        \D_cache/cache[1][121] ), .A1N(n3916), .Y(\D_cache/n827 ) );
  OAI2BB2XL U8329 ( .B0(\D_cache/n262 ), .B1(n3928), .A0N(
        \D_cache/cache[0][121] ), .A1N(n3937), .Y(\D_cache/n828 ) );
  OAI2BB2XL U8330 ( .B0(\D_cache/n264 ), .B1(n3788), .A0N(
        \D_cache/cache[7][120] ), .A1N(n3795), .Y(\D_cache/n829 ) );
  OAI2BB2XL U8331 ( .B0(\D_cache/n264 ), .B1(n3808), .A0N(
        \D_cache/cache[6][120] ), .A1N(n3815), .Y(\D_cache/n830 ) );
  OAI2BB2XL U8332 ( .B0(\D_cache/n264 ), .B1(n3827), .A0N(
        \D_cache/cache[5][120] ), .A1N(n3833), .Y(\D_cache/n831 ) );
  OAI2BB2XL U8333 ( .B0(\D_cache/n264 ), .B1(n3846), .A0N(
        \D_cache/cache[4][120] ), .A1N(n3855), .Y(\D_cache/n832 ) );
  OAI2BB2XL U8334 ( .B0(\D_cache/n264 ), .B1(n3866), .A0N(
        \D_cache/cache[3][120] ), .A1N(n3874), .Y(\D_cache/n833 ) );
  OAI2BB2XL U8335 ( .B0(\D_cache/n264 ), .B1(n3888), .A0N(
        \D_cache/cache[2][120] ), .A1N(n3895), .Y(\D_cache/n834 ) );
  OAI2BB2XL U8336 ( .B0(\D_cache/n264 ), .B1(n3908), .A0N(
        \D_cache/cache[1][120] ), .A1N(n3916), .Y(\D_cache/n835 ) );
  OAI2BB2XL U8337 ( .B0(\D_cache/n264 ), .B1(n3928), .A0N(
        \D_cache/cache[0][120] ), .A1N(n3937), .Y(\D_cache/n836 ) );
  OAI2BB2XL U8338 ( .B0(\D_cache/n266 ), .B1(n3788), .A0N(
        \D_cache/cache[7][119] ), .A1N(n3795), .Y(\D_cache/n837 ) );
  OAI2BB2XL U8339 ( .B0(\D_cache/n266 ), .B1(n3808), .A0N(
        \D_cache/cache[6][119] ), .A1N(n3815), .Y(\D_cache/n838 ) );
  OAI2BB2XL U8340 ( .B0(\D_cache/n266 ), .B1(n3827), .A0N(
        \D_cache/cache[5][119] ), .A1N(n3833), .Y(\D_cache/n839 ) );
  OAI2BB2XL U8341 ( .B0(\D_cache/n266 ), .B1(n3846), .A0N(
        \D_cache/cache[4][119] ), .A1N(n3855), .Y(\D_cache/n840 ) );
  OAI2BB2XL U8342 ( .B0(\D_cache/n266 ), .B1(n3868), .A0N(
        \D_cache/cache[3][119] ), .A1N(n3874), .Y(\D_cache/n841 ) );
  OAI2BB2XL U8343 ( .B0(\D_cache/n266 ), .B1(n3888), .A0N(
        \D_cache/cache[2][119] ), .A1N(n3895), .Y(\D_cache/n842 ) );
  OAI2BB2XL U8344 ( .B0(\D_cache/n266 ), .B1(n3908), .A0N(
        \D_cache/cache[1][119] ), .A1N(n3916), .Y(\D_cache/n843 ) );
  OAI2BB2XL U8345 ( .B0(\D_cache/n266 ), .B1(n3928), .A0N(
        \D_cache/cache[0][119] ), .A1N(n3937), .Y(\D_cache/n844 ) );
  OAI2BB2XL U8346 ( .B0(\D_cache/n268 ), .B1(n3787), .A0N(
        \D_cache/cache[7][118] ), .A1N(n3795), .Y(\D_cache/n845 ) );
  OAI2BB2XL U8347 ( .B0(\D_cache/n268 ), .B1(n3807), .A0N(
        \D_cache/cache[6][118] ), .A1N(n3815), .Y(\D_cache/n846 ) );
  OAI2BB2XL U8348 ( .B0(\D_cache/n268 ), .B1(n3826), .A0N(
        \D_cache/cache[5][118] ), .A1N(n3833), .Y(\D_cache/n847 ) );
  OAI2BB2XL U8349 ( .B0(\D_cache/n268 ), .B1(n3845), .A0N(
        \D_cache/cache[4][118] ), .A1N(n3855), .Y(\D_cache/n848 ) );
  OAI2BB2XL U8350 ( .B0(\D_cache/n268 ), .B1(n3865), .A0N(
        \D_cache/cache[3][118] ), .A1N(n3874), .Y(\D_cache/n849 ) );
  OAI2BB2XL U8351 ( .B0(\D_cache/n268 ), .B1(n3887), .A0N(
        \D_cache/cache[2][118] ), .A1N(n3895), .Y(\D_cache/n850 ) );
  OAI2BB2XL U8352 ( .B0(\D_cache/n268 ), .B1(n3907), .A0N(
        \D_cache/cache[1][118] ), .A1N(n3916), .Y(\D_cache/n851 ) );
  OAI2BB2XL U8353 ( .B0(\D_cache/n268 ), .B1(n3927), .A0N(
        \D_cache/cache[0][118] ), .A1N(n3937), .Y(\D_cache/n852 ) );
  OAI2BB2XL U8354 ( .B0(\D_cache/n270 ), .B1(n3787), .A0N(
        \D_cache/cache[7][117] ), .A1N(n3795), .Y(\D_cache/n853 ) );
  OAI2BB2XL U8355 ( .B0(\D_cache/n270 ), .B1(n3807), .A0N(
        \D_cache/cache[6][117] ), .A1N(n3815), .Y(\D_cache/n854 ) );
  OAI2BB2XL U8356 ( .B0(\D_cache/n270 ), .B1(n3826), .A0N(
        \D_cache/cache[5][117] ), .A1N(n3833), .Y(\D_cache/n855 ) );
  OAI2BB2XL U8357 ( .B0(\D_cache/n270 ), .B1(n3845), .A0N(
        \D_cache/cache[4][117] ), .A1N(n3855), .Y(\D_cache/n856 ) );
  OAI2BB2XL U8358 ( .B0(\D_cache/n270 ), .B1(n3865), .A0N(
        \D_cache/cache[3][117] ), .A1N(n3874), .Y(\D_cache/n857 ) );
  OAI2BB2XL U8359 ( .B0(\D_cache/n270 ), .B1(n3887), .A0N(
        \D_cache/cache[2][117] ), .A1N(n3895), .Y(\D_cache/n858 ) );
  OAI2BB2XL U8360 ( .B0(\D_cache/n270 ), .B1(n3907), .A0N(
        \D_cache/cache[1][117] ), .A1N(n3916), .Y(\D_cache/n859 ) );
  OAI2BB2XL U8361 ( .B0(\D_cache/n270 ), .B1(n3927), .A0N(
        \D_cache/cache[0][117] ), .A1N(n3937), .Y(\D_cache/n860 ) );
  OAI2BB2XL U8362 ( .B0(\D_cache/n272 ), .B1(n3787), .A0N(
        \D_cache/cache[7][116] ), .A1N(n3795), .Y(\D_cache/n861 ) );
  OAI2BB2XL U8363 ( .B0(\D_cache/n272 ), .B1(n3807), .A0N(
        \D_cache/cache[6][116] ), .A1N(n3815), .Y(\D_cache/n862 ) );
  OAI2BB2XL U8364 ( .B0(\D_cache/n272 ), .B1(n3826), .A0N(
        \D_cache/cache[5][116] ), .A1N(n3833), .Y(\D_cache/n863 ) );
  OAI2BB2XL U8365 ( .B0(\D_cache/n272 ), .B1(n3845), .A0N(
        \D_cache/cache[4][116] ), .A1N(n3855), .Y(\D_cache/n864 ) );
  OAI2BB2XL U8366 ( .B0(\D_cache/n272 ), .B1(n3866), .A0N(
        \D_cache/cache[3][116] ), .A1N(n3874), .Y(\D_cache/n865 ) );
  OAI2BB2XL U8367 ( .B0(\D_cache/n272 ), .B1(n3887), .A0N(
        \D_cache/cache[2][116] ), .A1N(n3895), .Y(\D_cache/n866 ) );
  OAI2BB2XL U8368 ( .B0(\D_cache/n272 ), .B1(n3907), .A0N(
        \D_cache/cache[1][116] ), .A1N(n3916), .Y(\D_cache/n867 ) );
  OAI2BB2XL U8369 ( .B0(\D_cache/n272 ), .B1(n3927), .A0N(
        \D_cache/cache[0][116] ), .A1N(n3937), .Y(\D_cache/n868 ) );
  OAI2BB2XL U8370 ( .B0(\D_cache/n274 ), .B1(n3787), .A0N(
        \D_cache/cache[7][115] ), .A1N(n3796), .Y(\D_cache/n869 ) );
  OAI2BB2XL U8371 ( .B0(\D_cache/n274 ), .B1(n3807), .A0N(
        \D_cache/cache[6][115] ), .A1N(n3816), .Y(\D_cache/n870 ) );
  OAI2BB2XL U8372 ( .B0(\D_cache/n274 ), .B1(n3826), .A0N(
        \D_cache/cache[5][115] ), .A1N(n3834), .Y(\D_cache/n871 ) );
  OAI2BB2XL U8373 ( .B0(\D_cache/n274 ), .B1(n3845), .A0N(
        \D_cache/cache[4][115] ), .A1N(n3856), .Y(\D_cache/n872 ) );
  OAI2BB2XL U8374 ( .B0(\D_cache/n274 ), .B1(n3868), .A0N(
        \D_cache/cache[3][115] ), .A1N(n3875), .Y(\D_cache/n873 ) );
  OAI2BB2XL U8375 ( .B0(\D_cache/n274 ), .B1(n3887), .A0N(
        \D_cache/cache[2][115] ), .A1N(n3896), .Y(\D_cache/n874 ) );
  OAI2BB2XL U8376 ( .B0(\D_cache/n274 ), .B1(n3907), .A0N(
        \D_cache/cache[1][115] ), .A1N(n3917), .Y(\D_cache/n875 ) );
  OAI2BB2XL U8377 ( .B0(\D_cache/n274 ), .B1(n3927), .A0N(
        \D_cache/cache[0][115] ), .A1N(n3938), .Y(\D_cache/n876 ) );
  OAI2BB2XL U8378 ( .B0(\D_cache/n276 ), .B1(n3786), .A0N(
        \D_cache/cache[7][114] ), .A1N(n3796), .Y(\D_cache/n877 ) );
  OAI2BB2XL U8379 ( .B0(\D_cache/n276 ), .B1(n3806), .A0N(
        \D_cache/cache[6][114] ), .A1N(n3816), .Y(\D_cache/n878 ) );
  OAI2BB2XL U8380 ( .B0(\D_cache/n276 ), .B1(n3825), .A0N(
        \D_cache/cache[5][114] ), .A1N(n3834), .Y(\D_cache/n879 ) );
  OAI2BB2XL U8381 ( .B0(\D_cache/n276 ), .B1(n3844), .A0N(
        \D_cache/cache[4][114] ), .A1N(n3856), .Y(\D_cache/n880 ) );
  OAI2BB2XL U8382 ( .B0(\D_cache/n276 ), .B1(n3865), .A0N(
        \D_cache/cache[3][114] ), .A1N(n3875), .Y(\D_cache/n881 ) );
  OAI2BB2XL U8383 ( .B0(\D_cache/n276 ), .B1(n3886), .A0N(
        \D_cache/cache[2][114] ), .A1N(n3896), .Y(\D_cache/n882 ) );
  OAI2BB2XL U8384 ( .B0(\D_cache/n276 ), .B1(n3906), .A0N(
        \D_cache/cache[1][114] ), .A1N(n3917), .Y(\D_cache/n883 ) );
  OAI2BB2XL U8385 ( .B0(\D_cache/n276 ), .B1(n3926), .A0N(
        \D_cache/cache[0][114] ), .A1N(n3938), .Y(\D_cache/n884 ) );
  OAI2BB2XL U8386 ( .B0(\D_cache/n278 ), .B1(n3786), .A0N(
        \D_cache/cache[7][113] ), .A1N(n3796), .Y(\D_cache/n885 ) );
  OAI2BB2XL U8387 ( .B0(\D_cache/n278 ), .B1(n3806), .A0N(
        \D_cache/cache[6][113] ), .A1N(n3816), .Y(\D_cache/n886 ) );
  OAI2BB2XL U8388 ( .B0(\D_cache/n278 ), .B1(n3825), .A0N(
        \D_cache/cache[5][113] ), .A1N(n3834), .Y(\D_cache/n887 ) );
  OAI2BB2XL U8389 ( .B0(\D_cache/n278 ), .B1(n3844), .A0N(
        \D_cache/cache[4][113] ), .A1N(n3856), .Y(\D_cache/n888 ) );
  OAI2BB2XL U8390 ( .B0(\D_cache/n278 ), .B1(n3865), .A0N(
        \D_cache/cache[3][113] ), .A1N(n3875), .Y(\D_cache/n889 ) );
  OAI2BB2XL U8391 ( .B0(\D_cache/n278 ), .B1(n3886), .A0N(
        \D_cache/cache[2][113] ), .A1N(n3896), .Y(\D_cache/n890 ) );
  OAI2BB2XL U8392 ( .B0(\D_cache/n278 ), .B1(n3906), .A0N(
        \D_cache/cache[1][113] ), .A1N(n3917), .Y(\D_cache/n891 ) );
  OAI2BB2XL U8393 ( .B0(\D_cache/n278 ), .B1(n3926), .A0N(
        \D_cache/cache[0][113] ), .A1N(n3938), .Y(\D_cache/n892 ) );
  OAI2BB2XL U8394 ( .B0(\D_cache/n280 ), .B1(n3786), .A0N(
        \D_cache/cache[7][112] ), .A1N(n3796), .Y(\D_cache/n893 ) );
  OAI2BB2XL U8395 ( .B0(\D_cache/n280 ), .B1(n3806), .A0N(
        \D_cache/cache[6][112] ), .A1N(n3816), .Y(\D_cache/n894 ) );
  OAI2BB2XL U8396 ( .B0(\D_cache/n280 ), .B1(n3825), .A0N(
        \D_cache/cache[5][112] ), .A1N(n3834), .Y(\D_cache/n895 ) );
  OAI2BB2XL U8397 ( .B0(\D_cache/n280 ), .B1(n3844), .A0N(
        \D_cache/cache[4][112] ), .A1N(n3856), .Y(\D_cache/n896 ) );
  OAI2BB2XL U8398 ( .B0(\D_cache/n280 ), .B1(n3865), .A0N(
        \D_cache/cache[3][112] ), .A1N(n3875), .Y(\D_cache/n897 ) );
  OAI2BB2XL U8399 ( .B0(\D_cache/n280 ), .B1(n3886), .A0N(
        \D_cache/cache[2][112] ), .A1N(n3896), .Y(\D_cache/n898 ) );
  OAI2BB2XL U8400 ( .B0(\D_cache/n280 ), .B1(n3906), .A0N(
        \D_cache/cache[1][112] ), .A1N(n3917), .Y(\D_cache/n899 ) );
  OAI2BB2XL U8401 ( .B0(\D_cache/n280 ), .B1(n3926), .A0N(
        \D_cache/cache[0][112] ), .A1N(n3938), .Y(\D_cache/n900 ) );
  OAI2BB2XL U8402 ( .B0(\D_cache/n282 ), .B1(n3786), .A0N(
        \D_cache/cache[7][111] ), .A1N(n3796), .Y(\D_cache/n901 ) );
  OAI2BB2XL U8403 ( .B0(\D_cache/n282 ), .B1(n3806), .A0N(
        \D_cache/cache[6][111] ), .A1N(n3816), .Y(\D_cache/n902 ) );
  OAI2BB2XL U8404 ( .B0(\D_cache/n282 ), .B1(n3825), .A0N(
        \D_cache/cache[5][111] ), .A1N(n3834), .Y(\D_cache/n903 ) );
  OAI2BB2XL U8405 ( .B0(\D_cache/n282 ), .B1(n3844), .A0N(
        \D_cache/cache[4][111] ), .A1N(n3856), .Y(\D_cache/n904 ) );
  OAI2BB2XL U8406 ( .B0(\D_cache/n282 ), .B1(n3865), .A0N(
        \D_cache/cache[3][111] ), .A1N(n3875), .Y(\D_cache/n905 ) );
  OAI2BB2XL U8407 ( .B0(\D_cache/n282 ), .B1(n3886), .A0N(
        \D_cache/cache[2][111] ), .A1N(n3896), .Y(\D_cache/n906 ) );
  OAI2BB2XL U8408 ( .B0(\D_cache/n282 ), .B1(n3906), .A0N(
        \D_cache/cache[1][111] ), .A1N(n3917), .Y(\D_cache/n907 ) );
  OAI2BB2XL U8409 ( .B0(\D_cache/n282 ), .B1(n3926), .A0N(
        \D_cache/cache[0][111] ), .A1N(n3938), .Y(\D_cache/n908 ) );
  OAI2BB2XL U8410 ( .B0(\D_cache/n284 ), .B1(n3785), .A0N(
        \D_cache/cache[7][110] ), .A1N(n3796), .Y(\D_cache/n909 ) );
  OAI2BB2XL U8411 ( .B0(\D_cache/n284 ), .B1(n3805), .A0N(
        \D_cache/cache[6][110] ), .A1N(n3816), .Y(\D_cache/n910 ) );
  OAI2BB2XL U8412 ( .B0(\D_cache/n284 ), .B1(n3824), .A0N(
        \D_cache/cache[5][110] ), .A1N(n3834), .Y(\D_cache/n911 ) );
  OAI2BB2XL U8413 ( .B0(\D_cache/n284 ), .B1(n3862), .A0N(
        \D_cache/cache[4][110] ), .A1N(n3856), .Y(\D_cache/n912 ) );
  OAI2BB2XL U8414 ( .B0(\D_cache/n284 ), .B1(n3864), .A0N(
        \D_cache/cache[3][110] ), .A1N(n3875), .Y(\D_cache/n913 ) );
  OAI2BB2XL U8415 ( .B0(\D_cache/n284 ), .B1(n3885), .A0N(
        \D_cache/cache[2][110] ), .A1N(n3896), .Y(\D_cache/n914 ) );
  OAI2BB2XL U8416 ( .B0(\D_cache/n284 ), .B1(n3905), .A0N(
        \D_cache/cache[1][110] ), .A1N(n3917), .Y(\D_cache/n915 ) );
  OAI2BB2XL U8417 ( .B0(\D_cache/n284 ), .B1(n3925), .A0N(
        \D_cache/cache[0][110] ), .A1N(n3938), .Y(\D_cache/n916 ) );
  OAI2BB2XL U8418 ( .B0(\D_cache/n286 ), .B1(n3785), .A0N(
        \D_cache/cache[7][109] ), .A1N(n3796), .Y(\D_cache/n917 ) );
  OAI2BB2XL U8419 ( .B0(\D_cache/n286 ), .B1(n3805), .A0N(
        \D_cache/cache[6][109] ), .A1N(n3816), .Y(\D_cache/n918 ) );
  OAI2BB2XL U8420 ( .B0(\D_cache/n286 ), .B1(n3824), .A0N(
        \D_cache/cache[5][109] ), .A1N(n3834), .Y(\D_cache/n919 ) );
  OAI2BB2XL U8421 ( .B0(\D_cache/n286 ), .B1(n3858), .A0N(
        \D_cache/cache[4][109] ), .A1N(n3856), .Y(\D_cache/n920 ) );
  OAI2BB2XL U8422 ( .B0(\D_cache/n286 ), .B1(n3864), .A0N(
        \D_cache/cache[3][109] ), .A1N(n3875), .Y(\D_cache/n921 ) );
  OAI2BB2XL U8423 ( .B0(\D_cache/n286 ), .B1(n3885), .A0N(
        \D_cache/cache[2][109] ), .A1N(n3896), .Y(\D_cache/n922 ) );
  OAI2BB2XL U8424 ( .B0(\D_cache/n286 ), .B1(n3905), .A0N(
        \D_cache/cache[1][109] ), .A1N(n3917), .Y(\D_cache/n923 ) );
  OAI2BB2XL U8425 ( .B0(\D_cache/n286 ), .B1(n3925), .A0N(
        \D_cache/cache[0][109] ), .A1N(n3938), .Y(\D_cache/n924 ) );
  OAI2BB2XL U8426 ( .B0(\D_cache/n288 ), .B1(n3785), .A0N(
        \D_cache/cache[7][108] ), .A1N(n3797), .Y(\D_cache/n925 ) );
  OAI2BB2XL U8427 ( .B0(\D_cache/n288 ), .B1(n3805), .A0N(
        \D_cache/cache[6][108] ), .A1N(n3817), .Y(\D_cache/n926 ) );
  OAI2BB2XL U8428 ( .B0(\D_cache/n288 ), .B1(n3824), .A0N(
        \D_cache/cache[5][108] ), .A1N(n3835), .Y(\D_cache/n927 ) );
  OAI2BB2XL U8429 ( .B0(\D_cache/n288 ), .B1(n3862), .A0N(
        \D_cache/cache[4][108] ), .A1N(n3857), .Y(\D_cache/n928 ) );
  OAI2BB2XL U8430 ( .B0(\D_cache/n288 ), .B1(n3864), .A0N(
        \D_cache/cache[3][108] ), .A1N(n3876), .Y(\D_cache/n929 ) );
  OAI2BB2XL U8431 ( .B0(\D_cache/n288 ), .B1(n3885), .A0N(
        \D_cache/cache[2][108] ), .A1N(n3897), .Y(\D_cache/n930 ) );
  OAI2BB2XL U8432 ( .B0(\D_cache/n288 ), .B1(n3905), .A0N(
        \D_cache/cache[1][108] ), .A1N(n3918), .Y(\D_cache/n931 ) );
  OAI2BB2XL U8433 ( .B0(\D_cache/n288 ), .B1(n3925), .A0N(
        \D_cache/cache[0][108] ), .A1N(n3939), .Y(\D_cache/n932 ) );
  OAI2BB2XL U8434 ( .B0(\D_cache/n290 ), .B1(n3785), .A0N(
        \D_cache/cache[7][107] ), .A1N(n3797), .Y(\D_cache/n933 ) );
  OAI2BB2XL U8435 ( .B0(\D_cache/n290 ), .B1(n3805), .A0N(
        \D_cache/cache[6][107] ), .A1N(n3817), .Y(\D_cache/n934 ) );
  OAI2BB2XL U8436 ( .B0(\D_cache/n290 ), .B1(n3824), .A0N(
        \D_cache/cache[5][107] ), .A1N(n3835), .Y(\D_cache/n935 ) );
  OAI2BB2XL U8437 ( .B0(\D_cache/n290 ), .B1(n3858), .A0N(
        \D_cache/cache[4][107] ), .A1N(n3857), .Y(\D_cache/n936 ) );
  OAI2BB2XL U8438 ( .B0(\D_cache/n290 ), .B1(n3864), .A0N(
        \D_cache/cache[3][107] ), .A1N(n3876), .Y(\D_cache/n937 ) );
  OAI2BB2XL U8439 ( .B0(\D_cache/n290 ), .B1(n3885), .A0N(
        \D_cache/cache[2][107] ), .A1N(n3897), .Y(\D_cache/n938 ) );
  OAI2BB2XL U8440 ( .B0(\D_cache/n290 ), .B1(n3905), .A0N(
        \D_cache/cache[1][107] ), .A1N(n3918), .Y(\D_cache/n939 ) );
  OAI2BB2XL U8441 ( .B0(\D_cache/n290 ), .B1(n3925), .A0N(
        \D_cache/cache[0][107] ), .A1N(n3939), .Y(\D_cache/n940 ) );
  OAI2BB2XL U8442 ( .B0(\D_cache/n292 ), .B1(n3784), .A0N(
        \D_cache/cache[7][106] ), .A1N(n3797), .Y(\D_cache/n941 ) );
  OAI2BB2XL U8443 ( .B0(\D_cache/n292 ), .B1(n3804), .A0N(
        \D_cache/cache[6][106] ), .A1N(n3817), .Y(\D_cache/n942 ) );
  OAI2BB2XL U8444 ( .B0(\D_cache/n292 ), .B1(n3824), .A0N(
        \D_cache/cache[5][106] ), .A1N(n3835), .Y(\D_cache/n943 ) );
  OAI2BB2XL U8445 ( .B0(\D_cache/n292 ), .B1(n3853), .A0N(
        \D_cache/cache[4][106] ), .A1N(n3857), .Y(\D_cache/n944 ) );
  OAI2BB2XL U8446 ( .B0(\D_cache/n292 ), .B1(n3867), .A0N(
        \D_cache/cache[3][106] ), .A1N(n3876), .Y(\D_cache/n945 ) );
  OAI2BB2XL U8447 ( .B0(\D_cache/n292 ), .B1(n3884), .A0N(
        \D_cache/cache[2][106] ), .A1N(n3897), .Y(\D_cache/n946 ) );
  OAI2BB2XL U8448 ( .B0(\D_cache/n292 ), .B1(n3904), .A0N(
        \D_cache/cache[1][106] ), .A1N(n3918), .Y(\D_cache/n947 ) );
  OAI2BB2XL U8449 ( .B0(\D_cache/n292 ), .B1(n3925), .A0N(
        \D_cache/cache[0][106] ), .A1N(n3939), .Y(\D_cache/n948 ) );
  OAI2BB2XL U8450 ( .B0(\D_cache/n294 ), .B1(n3784), .A0N(
        \D_cache/cache[7][105] ), .A1N(n3797), .Y(\D_cache/n949 ) );
  OAI2BB2XL U8451 ( .B0(\D_cache/n294 ), .B1(n3804), .A0N(
        \D_cache/cache[6][105] ), .A1N(n3817), .Y(\D_cache/n950 ) );
  OAI2BB2XL U8452 ( .B0(\D_cache/n294 ), .B1(n3824), .A0N(
        \D_cache/cache[5][105] ), .A1N(n3835), .Y(\D_cache/n951 ) );
  OAI2BB2XL U8453 ( .B0(\D_cache/n294 ), .B1(n3852), .A0N(
        \D_cache/cache[4][105] ), .A1N(n3857), .Y(\D_cache/n952 ) );
  OAI2BB2XL U8454 ( .B0(\D_cache/n294 ), .B1(n3872), .A0N(
        \D_cache/cache[3][105] ), .A1N(n3876), .Y(\D_cache/n953 ) );
  OAI2BB2XL U8455 ( .B0(\D_cache/n294 ), .B1(n3884), .A0N(
        \D_cache/cache[2][105] ), .A1N(n3897), .Y(\D_cache/n954 ) );
  OAI2BB2XL U8456 ( .B0(\D_cache/n294 ), .B1(n3904), .A0N(
        \D_cache/cache[1][105] ), .A1N(n3918), .Y(\D_cache/n955 ) );
  OAI2BB2XL U8457 ( .B0(\D_cache/n294 ), .B1(n3925), .A0N(
        \D_cache/cache[0][105] ), .A1N(n3939), .Y(\D_cache/n956 ) );
  OAI2BB2XL U8458 ( .B0(\D_cache/n296 ), .B1(n3784), .A0N(
        \D_cache/cache[7][104] ), .A1N(n3797), .Y(\D_cache/n957 ) );
  OAI2BB2XL U8459 ( .B0(\D_cache/n296 ), .B1(n3804), .A0N(
        \D_cache/cache[6][104] ), .A1N(n3817), .Y(\D_cache/n958 ) );
  OAI2BB2XL U8460 ( .B0(\D_cache/n296 ), .B1(n3830), .A0N(
        \D_cache/cache[5][104] ), .A1N(n3835), .Y(\D_cache/n959 ) );
  OAI2BB2XL U8461 ( .B0(\D_cache/n296 ), .B1(n3853), .A0N(
        \D_cache/cache[4][104] ), .A1N(n3857), .Y(\D_cache/n960 ) );
  OAI2BB2XL U8462 ( .B0(\D_cache/n296 ), .B1(n3870), .A0N(
        \D_cache/cache[3][104] ), .A1N(n3876), .Y(\D_cache/n961 ) );
  OAI2BB2XL U8463 ( .B0(\D_cache/n296 ), .B1(n3884), .A0N(
        \D_cache/cache[2][104] ), .A1N(n3897), .Y(\D_cache/n962 ) );
  OAI2BB2XL U8464 ( .B0(\D_cache/n296 ), .B1(n3904), .A0N(
        \D_cache/cache[1][104] ), .A1N(n3918), .Y(\D_cache/n963 ) );
  OAI2BB2XL U8465 ( .B0(\D_cache/n296 ), .B1(n3925), .A0N(
        \D_cache/cache[0][104] ), .A1N(n3939), .Y(\D_cache/n964 ) );
  OAI2BB2XL U8466 ( .B0(\D_cache/n300 ), .B1(n3784), .A0N(
        \D_cache/cache[7][102] ), .A1N(n3802), .Y(\D_cache/n973 ) );
  OAI2BB2XL U8467 ( .B0(\D_cache/n300 ), .B1(n3804), .A0N(
        \D_cache/cache[6][102] ), .A1N(n3822), .Y(\D_cache/n974 ) );
  OAI2BB2XL U8468 ( .B0(\D_cache/n300 ), .B1(n3829), .A0N(
        \D_cache/cache[5][102] ), .A1N(n3839), .Y(\D_cache/n975 ) );
  OAI2BB2XL U8469 ( .B0(\D_cache/n300 ), .B1(n3852), .A0N(
        \D_cache/cache[4][102] ), .A1N(n3862), .Y(\D_cache/n976 ) );
  OAI2BB2XL U8470 ( .B0(\D_cache/n300 ), .B1(n3869), .A0N(
        \D_cache/cache[3][102] ), .A1N(n3881), .Y(\D_cache/n977 ) );
  OAI2BB2XL U8471 ( .B0(\D_cache/n300 ), .B1(n3884), .A0N(
        \D_cache/cache[2][102] ), .A1N(n3902), .Y(\D_cache/n978 ) );
  OAI2BB2XL U8472 ( .B0(\D_cache/n300 ), .B1(n3904), .A0N(
        \D_cache/cache[1][102] ), .A1N(n3923), .Y(\D_cache/n979 ) );
  OAI2BB2XL U8473 ( .B0(\D_cache/n300 ), .B1(n3925), .A0N(
        \D_cache/cache[0][102] ), .A1N(n3944), .Y(\D_cache/n980 ) );
  OAI2BB2XL U8474 ( .B0(\D_cache/n302 ), .B1(n3784), .A0N(
        \D_cache/cache[7][101] ), .A1N(n3802), .Y(\D_cache/n981 ) );
  OAI2BB2XL U8475 ( .B0(\D_cache/n302 ), .B1(n3804), .A0N(
        \D_cache/cache[6][101] ), .A1N(n3822), .Y(\D_cache/n982 ) );
  OAI2BB2XL U8476 ( .B0(\D_cache/n302 ), .B1(n3824), .A0N(
        \D_cache/cache[5][101] ), .A1N(n3839), .Y(\D_cache/n983 ) );
  OAI2BB2XL U8477 ( .B0(\D_cache/n302 ), .B1(n3853), .A0N(
        \D_cache/cache[4][101] ), .A1N(n3862), .Y(\D_cache/n984 ) );
  OAI2BB2XL U8478 ( .B0(\D_cache/n302 ), .B1(n3871), .A0N(
        \D_cache/cache[3][101] ), .A1N(n3881), .Y(\D_cache/n985 ) );
  OAI2BB2XL U8479 ( .B0(\D_cache/n302 ), .B1(n3884), .A0N(
        \D_cache/cache[2][101] ), .A1N(n3902), .Y(\D_cache/n986 ) );
  OAI2BB2XL U8480 ( .B0(\D_cache/n302 ), .B1(n3904), .A0N(
        \D_cache/cache[1][101] ), .A1N(n3923), .Y(\D_cache/n987 ) );
  OAI2BB2XL U8481 ( .B0(\D_cache/n302 ), .B1(n3925), .A0N(
        \D_cache/cache[0][101] ), .A1N(n3944), .Y(\D_cache/n988 ) );
  OAI2BB2XL U8482 ( .B0(\D_cache/n304 ), .B1(n3784), .A0N(
        \D_cache/cache[7][100] ), .A1N(n3802), .Y(\D_cache/n989 ) );
  OAI2BB2XL U8483 ( .B0(\D_cache/n304 ), .B1(n3804), .A0N(
        \D_cache/cache[6][100] ), .A1N(n3822), .Y(\D_cache/n990 ) );
  OAI2BB2XL U8484 ( .B0(\D_cache/n304 ), .B1(n3830), .A0N(
        \D_cache/cache[5][100] ), .A1N(n3839), .Y(\D_cache/n991 ) );
  OAI2BB2XL U8485 ( .B0(\D_cache/n304 ), .B1(n3852), .A0N(
        \D_cache/cache[4][100] ), .A1N(n3862), .Y(\D_cache/n992 ) );
  OAI2BB2XL U8486 ( .B0(\D_cache/n304 ), .B1(n3864), .A0N(
        \D_cache/cache[3][100] ), .A1N(n3881), .Y(\D_cache/n993 ) );
  OAI2BB2XL U8487 ( .B0(\D_cache/n304 ), .B1(n3884), .A0N(
        \D_cache/cache[2][100] ), .A1N(n3902), .Y(\D_cache/n994 ) );
  OAI2BB2XL U8488 ( .B0(\D_cache/n304 ), .B1(n3904), .A0N(
        \D_cache/cache[1][100] ), .A1N(n3923), .Y(\D_cache/n995 ) );
  OAI2BB2XL U8489 ( .B0(\D_cache/n304 ), .B1(n3925), .A0N(
        \D_cache/cache[0][100] ), .A1N(n3944), .Y(\D_cache/n996 ) );
  OAI2BB2XL U8490 ( .B0(\D_cache/n306 ), .B1(n3784), .A0N(
        \D_cache/cache[7][99] ), .A1N(n3802), .Y(\D_cache/n997 ) );
  OAI2BB2XL U8491 ( .B0(\D_cache/n306 ), .B1(n3804), .A0N(
        \D_cache/cache[6][99] ), .A1N(n3822), .Y(\D_cache/n998 ) );
  OAI2BB2XL U8492 ( .B0(\D_cache/n306 ), .B1(n3828), .A0N(
        \D_cache/cache[5][99] ), .A1N(n3839), .Y(\D_cache/n999 ) );
  OAI2BB2XL U8493 ( .B0(\D_cache/n306 ), .B1(n3853), .A0N(
        \D_cache/cache[4][99] ), .A1N(n3862), .Y(\D_cache/n1000 ) );
  OAI2BB2XL U8494 ( .B0(\D_cache/n306 ), .B1(n3866), .A0N(
        \D_cache/cache[3][99] ), .A1N(n3881), .Y(\D_cache/n1001 ) );
  OAI2BB2XL U8495 ( .B0(\D_cache/n306 ), .B1(n3884), .A0N(
        \D_cache/cache[2][99] ), .A1N(n3902), .Y(\D_cache/n1002 ) );
  OAI2BB2XL U8496 ( .B0(\D_cache/n306 ), .B1(n3904), .A0N(
        \D_cache/cache[1][99] ), .A1N(n3923), .Y(\D_cache/n1003 ) );
  OAI2BB2XL U8497 ( .B0(\D_cache/n306 ), .B1(n3925), .A0N(
        \D_cache/cache[0][99] ), .A1N(n3944), .Y(\D_cache/n1004 ) );
  OAI2BB2XL U8498 ( .B0(\D_cache/n308 ), .B1(n3784), .A0N(
        \D_cache/cache[7][98] ), .A1N(n3802), .Y(\D_cache/n1005 ) );
  OAI2BB2XL U8499 ( .B0(\D_cache/n308 ), .B1(n3804), .A0N(
        \D_cache/cache[6][98] ), .A1N(n3822), .Y(\D_cache/n1006 ) );
  OAI2BB2XL U8500 ( .B0(\D_cache/n308 ), .B1(n3824), .A0N(
        \D_cache/cache[5][98] ), .A1N(n3839), .Y(\D_cache/n1007 ) );
  OAI2BB2XL U8501 ( .B0(\D_cache/n308 ), .B1(n3852), .A0N(
        \D_cache/cache[4][98] ), .A1N(n3862), .Y(\D_cache/n1008 ) );
  OAI2BB2XL U8502 ( .B0(\D_cache/n308 ), .B1(n3868), .A0N(
        \D_cache/cache[3][98] ), .A1N(n3881), .Y(\D_cache/n1009 ) );
  OAI2BB2XL U8503 ( .B0(\D_cache/n308 ), .B1(n3884), .A0N(
        \D_cache/cache[2][98] ), .A1N(n3902), .Y(\D_cache/n1010 ) );
  OAI2BB2XL U8504 ( .B0(\D_cache/n308 ), .B1(n3904), .A0N(
        \D_cache/cache[1][98] ), .A1N(n3923), .Y(\D_cache/n1011 ) );
  OAI2BB2XL U8505 ( .B0(\D_cache/n308 ), .B1(n3944), .A0N(
        \D_cache/cache[0][98] ), .A1N(n3944), .Y(\D_cache/n1012 ) );
  OAI2BB2XL U8506 ( .B0(\D_cache/n310 ), .B1(n3784), .A0N(
        \D_cache/cache[7][97] ), .A1N(n3802), .Y(\D_cache/n1013 ) );
  OAI2BB2XL U8507 ( .B0(\D_cache/n310 ), .B1(n3804), .A0N(
        \D_cache/cache[6][97] ), .A1N(n3822), .Y(\D_cache/n1014 ) );
  OAI2BB2XL U8508 ( .B0(\D_cache/n310 ), .B1(n3830), .A0N(
        \D_cache/cache[5][97] ), .A1N(n3839), .Y(\D_cache/n1015 ) );
  OAI2BB2XL U8509 ( .B0(\D_cache/n310 ), .B1(n3853), .A0N(
        \D_cache/cache[4][97] ), .A1N(n3862), .Y(\D_cache/n1016 ) );
  OAI2BB2XL U8510 ( .B0(\D_cache/n310 ), .B1(n3867), .A0N(
        \D_cache/cache[3][97] ), .A1N(n3881), .Y(\D_cache/n1017 ) );
  OAI2BB2XL U8511 ( .B0(\D_cache/n310 ), .B1(n3884), .A0N(
        \D_cache/cache[2][97] ), .A1N(n3902), .Y(\D_cache/n1018 ) );
  OAI2BB2XL U8512 ( .B0(\D_cache/n310 ), .B1(n3904), .A0N(
        \D_cache/cache[1][97] ), .A1N(n3923), .Y(\D_cache/n1019 ) );
  OAI2BB2XL U8513 ( .B0(\D_cache/n310 ), .B1(n3925), .A0N(
        \D_cache/cache[0][97] ), .A1N(n3944), .Y(\D_cache/n1020 ) );
  OAI2BB2XL U8514 ( .B0(\D_cache/n312 ), .B1(n3784), .A0N(
        \D_cache/cache[7][96] ), .A1N(n3802), .Y(\D_cache/n1021 ) );
  OAI2BB2XL U8515 ( .B0(\D_cache/n312 ), .B1(n3804), .A0N(
        \D_cache/cache[6][96] ), .A1N(n3822), .Y(\D_cache/n1022 ) );
  OAI2BB2XL U8516 ( .B0(\D_cache/n312 ), .B1(n3825), .A0N(
        \D_cache/cache[5][96] ), .A1N(n3839), .Y(\D_cache/n1023 ) );
  OAI2BB2XL U8517 ( .B0(\D_cache/n312 ), .B1(n3852), .A0N(
        \D_cache/cache[4][96] ), .A1N(n3862), .Y(\D_cache/n1024 ) );
  OAI2BB2XL U8518 ( .B0(\D_cache/n312 ), .B1(n3872), .A0N(
        \D_cache/cache[3][96] ), .A1N(n3881), .Y(\D_cache/n1025 ) );
  OAI2BB2XL U8519 ( .B0(\D_cache/n312 ), .B1(n3884), .A0N(
        \D_cache/cache[2][96] ), .A1N(n3902), .Y(\D_cache/n1026 ) );
  OAI2BB2XL U8520 ( .B0(\D_cache/n312 ), .B1(n3904), .A0N(
        \D_cache/cache[1][96] ), .A1N(n3923), .Y(\D_cache/n1027 ) );
  OAI2BB2XL U8521 ( .B0(\D_cache/n312 ), .B1(n3944), .A0N(
        \D_cache/cache[0][96] ), .A1N(n3944), .Y(\D_cache/n1028 ) );
  OAI2BB2XL U8522 ( .B0(\D_cache/n317 ), .B1(n3784), .A0N(
        \D_cache/cache[7][95] ), .A1N(n3802), .Y(\D_cache/n1029 ) );
  OAI2BB2XL U8523 ( .B0(\D_cache/n317 ), .B1(n3804), .A0N(
        \D_cache/cache[6][95] ), .A1N(n3822), .Y(\D_cache/n1030 ) );
  OAI2BB2XL U8524 ( .B0(\D_cache/n317 ), .B1(n3824), .A0N(
        \D_cache/cache[5][95] ), .A1N(n3839), .Y(\D_cache/n1031 ) );
  OAI2BB2XL U8525 ( .B0(\D_cache/n317 ), .B1(n3853), .A0N(
        \D_cache/cache[4][95] ), .A1N(n3862), .Y(\D_cache/n1032 ) );
  OAI2BB2XL U8526 ( .B0(\D_cache/n317 ), .B1(n3870), .A0N(
        \D_cache/cache[3][95] ), .A1N(n3881), .Y(\D_cache/n1033 ) );
  OAI2BB2XL U8527 ( .B0(\D_cache/n317 ), .B1(n3884), .A0N(
        \D_cache/cache[2][95] ), .A1N(n3902), .Y(\D_cache/n1034 ) );
  OAI2BB2XL U8528 ( .B0(\D_cache/n317 ), .B1(n3904), .A0N(
        \D_cache/cache[1][95] ), .A1N(n3923), .Y(\D_cache/n1035 ) );
  OAI2BB2XL U8529 ( .B0(\D_cache/n317 ), .B1(n3926), .A0N(
        \D_cache/cache[0][95] ), .A1N(n3944), .Y(\D_cache/n1036 ) );
  OAI2BB2XL U8530 ( .B0(\D_cache/n321 ), .B1(n3785), .A0N(
        \D_cache/cache[7][94] ), .A1N(n3802), .Y(\D_cache/n1037 ) );
  OAI2BB2XL U8531 ( .B0(\D_cache/n321 ), .B1(n3805), .A0N(
        \D_cache/cache[6][94] ), .A1N(n3822), .Y(\D_cache/n1038 ) );
  OAI2BB2XL U8532 ( .B0(\D_cache/n321 ), .B1(n3824), .A0N(
        \D_cache/cache[5][94] ), .A1N(n3839), .Y(\D_cache/n1039 ) );
  OAI2BB2XL U8533 ( .B0(\D_cache/n321 ), .B1(n3862), .A0N(
        \D_cache/cache[4][94] ), .A1N(n3862), .Y(\D_cache/n1040 ) );
  OAI2BB2XL U8534 ( .B0(\D_cache/n321 ), .B1(n3864), .A0N(
        \D_cache/cache[3][94] ), .A1N(n3881), .Y(\D_cache/n1041 ) );
  OAI2BB2XL U8535 ( .B0(\D_cache/n321 ), .B1(n3885), .A0N(
        \D_cache/cache[2][94] ), .A1N(n3902), .Y(\D_cache/n1042 ) );
  OAI2BB2XL U8536 ( .B0(\D_cache/n321 ), .B1(n3905), .A0N(
        \D_cache/cache[1][94] ), .A1N(n3923), .Y(\D_cache/n1043 ) );
  OAI2BB2XL U8537 ( .B0(\D_cache/n321 ), .B1(n3925), .A0N(
        \D_cache/cache[0][94] ), .A1N(n3944), .Y(\D_cache/n1044 ) );
  OAI2BB2XL U8538 ( .B0(\D_cache/n323 ), .B1(n3785), .A0N(
        \D_cache/cache[7][93] ), .A1N(n3802), .Y(\D_cache/n1045 ) );
  OAI2BB2XL U8539 ( .B0(\D_cache/n323 ), .B1(n3805), .A0N(
        \D_cache/cache[6][93] ), .A1N(n3822), .Y(\D_cache/n1046 ) );
  OAI2BB2XL U8540 ( .B0(\D_cache/n323 ), .B1(n3824), .A0N(
        \D_cache/cache[5][93] ), .A1N(n3839), .Y(\D_cache/n1047 ) );
  OAI2BB2XL U8541 ( .B0(\D_cache/n323 ), .B1(n3849), .A0N(
        \D_cache/cache[4][93] ), .A1N(n3862), .Y(\D_cache/n1048 ) );
  OAI2BB2XL U8542 ( .B0(\D_cache/n323 ), .B1(n3864), .A0N(
        \D_cache/cache[3][93] ), .A1N(n3881), .Y(\D_cache/n1049 ) );
  OAI2BB2XL U8543 ( .B0(\D_cache/n323 ), .B1(n3885), .A0N(
        \D_cache/cache[2][93] ), .A1N(n3902), .Y(\D_cache/n1050 ) );
  OAI2BB2XL U8544 ( .B0(\D_cache/n323 ), .B1(n3905), .A0N(
        \D_cache/cache[1][93] ), .A1N(n3923), .Y(\D_cache/n1051 ) );
  OAI2BB2XL U8545 ( .B0(\D_cache/n323 ), .B1(n3925), .A0N(
        \D_cache/cache[0][93] ), .A1N(n3944), .Y(\D_cache/n1052 ) );
  OAI2BB2XL U8546 ( .B0(\D_cache/n325 ), .B1(n3785), .A0N(
        \D_cache/cache[7][92] ), .A1N(n3802), .Y(\D_cache/n1053 ) );
  OAI2BB2XL U8547 ( .B0(\D_cache/n325 ), .B1(n3805), .A0N(
        \D_cache/cache[6][92] ), .A1N(n3822), .Y(\D_cache/n1054 ) );
  OAI2BB2XL U8548 ( .B0(\D_cache/n325 ), .B1(n3824), .A0N(
        \D_cache/cache[5][92] ), .A1N(n3839), .Y(\D_cache/n1055 ) );
  OAI2BB2XL U8549 ( .B0(\D_cache/n325 ), .B1(n3847), .A0N(
        \D_cache/cache[4][92] ), .A1N(n3862), .Y(\D_cache/n1056 ) );
  OAI2BB2XL U8550 ( .B0(\D_cache/n325 ), .B1(n3864), .A0N(
        \D_cache/cache[3][92] ), .A1N(n3881), .Y(\D_cache/n1057 ) );
  OAI2BB2XL U8551 ( .B0(\D_cache/n325 ), .B1(n3885), .A0N(
        \D_cache/cache[2][92] ), .A1N(n3902), .Y(\D_cache/n1058 ) );
  OAI2BB2XL U8552 ( .B0(\D_cache/n325 ), .B1(n3905), .A0N(
        \D_cache/cache[1][92] ), .A1N(n3923), .Y(\D_cache/n1059 ) );
  OAI2BB2XL U8553 ( .B0(\D_cache/n325 ), .B1(n3925), .A0N(
        \D_cache/cache[0][92] ), .A1N(n3944), .Y(\D_cache/n1060 ) );
  OAI2BB2XL U8554 ( .B0(\D_cache/n327 ), .B1(n3785), .A0N(
        \D_cache/cache[7][91] ), .A1N(n3802), .Y(\D_cache/n1061 ) );
  OAI2BB2XL U8555 ( .B0(\D_cache/n327 ), .B1(n3805), .A0N(
        \D_cache/cache[6][91] ), .A1N(n3822), .Y(\D_cache/n1062 ) );
  OAI2BB2XL U8556 ( .B0(\D_cache/n327 ), .B1(n3824), .A0N(
        \D_cache/cache[5][91] ), .A1N(n3839), .Y(\D_cache/n1063 ) );
  OAI2BB2XL U8557 ( .B0(\D_cache/n327 ), .B1(n3848), .A0N(
        \D_cache/cache[4][91] ), .A1N(n3862), .Y(\D_cache/n1064 ) );
  OAI2BB2XL U8558 ( .B0(\D_cache/n327 ), .B1(n3864), .A0N(
        \D_cache/cache[3][91] ), .A1N(n3881), .Y(\D_cache/n1065 ) );
  OAI2BB2XL U8559 ( .B0(\D_cache/n327 ), .B1(n3885), .A0N(
        \D_cache/cache[2][91] ), .A1N(n3902), .Y(\D_cache/n1066 ) );
  OAI2BB2XL U8560 ( .B0(\D_cache/n327 ), .B1(n3905), .A0N(
        \D_cache/cache[1][91] ), .A1N(n3923), .Y(\D_cache/n1067 ) );
  OAI2BB2XL U8561 ( .B0(\D_cache/n327 ), .B1(n3925), .A0N(
        \D_cache/cache[0][91] ), .A1N(n3944), .Y(\D_cache/n1068 ) );
  OAI2BB2XL U8562 ( .B0(\D_cache/n329 ), .B1(n3791), .A0N(
        \D_cache/cache[7][90] ), .A1N(n3802), .Y(\D_cache/n1069 ) );
  OAI2BB2XL U8563 ( .B0(\D_cache/n329 ), .B1(n3811), .A0N(
        \D_cache/cache[6][90] ), .A1N(n3822), .Y(\D_cache/n1070 ) );
  OAI2BB2XL U8564 ( .B0(\D_cache/n329 ), .B1(n3829), .A0N(
        \D_cache/cache[5][90] ), .A1N(n3839), .Y(\D_cache/n1071 ) );
  OAI2BB2XL U8565 ( .B0(\D_cache/n329 ), .B1(n3849), .A0N(
        \D_cache/cache[4][90] ), .A1N(n3862), .Y(\D_cache/n1072 ) );
  OAI2BB2XL U8566 ( .B0(\D_cache/n329 ), .B1(n3868), .A0N(
        \D_cache/cache[3][90] ), .A1N(n3881), .Y(\D_cache/n1073 ) );
  OAI2BB2XL U8567 ( .B0(\D_cache/n329 ), .B1(n3891), .A0N(
        \D_cache/cache[2][90] ), .A1N(n3902), .Y(\D_cache/n1074 ) );
  OAI2BB2XL U8568 ( .B0(\D_cache/n329 ), .B1(n3911), .A0N(
        \D_cache/cache[1][90] ), .A1N(n3923), .Y(\D_cache/n1075 ) );
  OAI2BB2XL U8569 ( .B0(\D_cache/n329 ), .B1(n3931), .A0N(
        \D_cache/cache[0][90] ), .A1N(n3944), .Y(\D_cache/n1076 ) );
  OAI2BB2XL U8570 ( .B0(\D_cache/n331 ), .B1(n3785), .A0N(
        \D_cache/cache[7][89] ), .A1N(n3802), .Y(\D_cache/n1077 ) );
  OAI2BB2XL U8571 ( .B0(\D_cache/n331 ), .B1(n3805), .A0N(
        \D_cache/cache[6][89] ), .A1N(n3822), .Y(\D_cache/n1078 ) );
  OAI2BB2XL U8572 ( .B0(\D_cache/n331 ), .B1(n3824), .A0N(
        \D_cache/cache[5][89] ), .A1N(n3839), .Y(\D_cache/n1079 ) );
  OAI2BB2XL U8573 ( .B0(\D_cache/n331 ), .B1(n3846), .A0N(
        \D_cache/cache[4][89] ), .A1N(n3862), .Y(\D_cache/n1080 ) );
  OAI2BB2XL U8574 ( .B0(\D_cache/n331 ), .B1(n3864), .A0N(
        \D_cache/cache[3][89] ), .A1N(n3881), .Y(\D_cache/n1081 ) );
  OAI2BB2XL U8575 ( .B0(\D_cache/n331 ), .B1(n3885), .A0N(
        \D_cache/cache[2][89] ), .A1N(n3902), .Y(\D_cache/n1082 ) );
  OAI2BB2XL U8576 ( .B0(\D_cache/n331 ), .B1(n3905), .A0N(
        \D_cache/cache[1][89] ), .A1N(n3923), .Y(\D_cache/n1083 ) );
  OAI2BB2XL U8577 ( .B0(\D_cache/n331 ), .B1(n3925), .A0N(
        \D_cache/cache[0][89] ), .A1N(n3944), .Y(\D_cache/n1084 ) );
  OAI2BB2XL U8578 ( .B0(\D_cache/n333 ), .B1(n3785), .A0N(
        \D_cache/cache[7][88] ), .A1N(n3802), .Y(\D_cache/n1085 ) );
  OAI2BB2XL U8579 ( .B0(\D_cache/n333 ), .B1(n3805), .A0N(
        \D_cache/cache[6][88] ), .A1N(n3822), .Y(\D_cache/n1086 ) );
  OAI2BB2XL U8580 ( .B0(\D_cache/n333 ), .B1(n3824), .A0N(
        \D_cache/cache[5][88] ), .A1N(n3839), .Y(\D_cache/n1087 ) );
  OAI2BB2XL U8581 ( .B0(\D_cache/n333 ), .B1(n3851), .A0N(
        \D_cache/cache[4][88] ), .A1N(n3862), .Y(\D_cache/n1088 ) );
  OAI2BB2XL U8582 ( .B0(\D_cache/n333 ), .B1(n3864), .A0N(
        \D_cache/cache[3][88] ), .A1N(n3881), .Y(\D_cache/n1089 ) );
  OAI2BB2XL U8583 ( .B0(\D_cache/n333 ), .B1(n3885), .A0N(
        \D_cache/cache[2][88] ), .A1N(n3902), .Y(\D_cache/n1090 ) );
  OAI2BB2XL U8584 ( .B0(\D_cache/n333 ), .B1(n3905), .A0N(
        \D_cache/cache[1][88] ), .A1N(n3923), .Y(\D_cache/n1091 ) );
  OAI2BB2XL U8585 ( .B0(\D_cache/n333 ), .B1(n3925), .A0N(
        \D_cache/cache[0][88] ), .A1N(n3944), .Y(\D_cache/n1092 ) );
  OAI2BB2XL U8586 ( .B0(\D_cache/n335 ), .B1(n3785), .A0N(
        \D_cache/cache[7][87] ), .A1N(n3802), .Y(\D_cache/n1093 ) );
  OAI2BB2XL U8587 ( .B0(\D_cache/n335 ), .B1(n3805), .A0N(
        \D_cache/cache[6][87] ), .A1N(n3822), .Y(\D_cache/n1094 ) );
  OAI2BB2XL U8588 ( .B0(\D_cache/n335 ), .B1(n3824), .A0N(
        \D_cache/cache[5][87] ), .A1N(n3839), .Y(\D_cache/n1095 ) );
  OAI2BB2XL U8589 ( .B0(\D_cache/n335 ), .B1(n3850), .A0N(
        \D_cache/cache[4][87] ), .A1N(n3862), .Y(\D_cache/n1096 ) );
  OAI2BB2XL U8590 ( .B0(\D_cache/n335 ), .B1(n3864), .A0N(
        \D_cache/cache[3][87] ), .A1N(n3881), .Y(\D_cache/n1097 ) );
  OAI2BB2XL U8591 ( .B0(\D_cache/n335 ), .B1(n3885), .A0N(
        \D_cache/cache[2][87] ), .A1N(n3902), .Y(\D_cache/n1098 ) );
  OAI2BB2XL U8592 ( .B0(\D_cache/n335 ), .B1(n3905), .A0N(
        \D_cache/cache[1][87] ), .A1N(n3923), .Y(\D_cache/n1099 ) );
  OAI2BB2XL U8593 ( .B0(\D_cache/n335 ), .B1(n3925), .A0N(
        \D_cache/cache[0][87] ), .A1N(n3944), .Y(\D_cache/n1100 ) );
  OAI2BB2XL U8594 ( .B0(\D_cache/n337 ), .B1(n3786), .A0N(
        \D_cache/cache[7][86] ), .A1N(n3802), .Y(\D_cache/n1101 ) );
  OAI2BB2XL U8595 ( .B0(\D_cache/n337 ), .B1(n3806), .A0N(
        \D_cache/cache[6][86] ), .A1N(n3822), .Y(\D_cache/n1102 ) );
  OAI2BB2XL U8596 ( .B0(\D_cache/n337 ), .B1(n3825), .A0N(
        \D_cache/cache[5][86] ), .A1N(n3839), .Y(\D_cache/n1103 ) );
  OAI2BB2XL U8597 ( .B0(\D_cache/n337 ), .B1(n3844), .A0N(
        \D_cache/cache[4][86] ), .A1N(n3862), .Y(\D_cache/n1104 ) );
  OAI2BB2XL U8598 ( .B0(\D_cache/n337 ), .B1(n3865), .A0N(
        \D_cache/cache[3][86] ), .A1N(n3881), .Y(\D_cache/n1105 ) );
  OAI2BB2XL U8599 ( .B0(\D_cache/n337 ), .B1(n3886), .A0N(
        \D_cache/cache[2][86] ), .A1N(n3902), .Y(\D_cache/n1106 ) );
  OAI2BB2XL U8600 ( .B0(\D_cache/n337 ), .B1(n3906), .A0N(
        \D_cache/cache[1][86] ), .A1N(n3923), .Y(\D_cache/n1107 ) );
  OAI2BB2XL U8601 ( .B0(\D_cache/n337 ), .B1(n3926), .A0N(
        \D_cache/cache[0][86] ), .A1N(n3944), .Y(\D_cache/n1108 ) );
  OAI2BB2XL U8602 ( .B0(\D_cache/n339 ), .B1(n3786), .A0N(
        \D_cache/cache[7][85] ), .A1N(n3802), .Y(\D_cache/n1109 ) );
  OAI2BB2XL U8603 ( .B0(\D_cache/n339 ), .B1(n3806), .A0N(
        \D_cache/cache[6][85] ), .A1N(n3822), .Y(\D_cache/n1110 ) );
  OAI2BB2XL U8604 ( .B0(\D_cache/n339 ), .B1(n3825), .A0N(
        \D_cache/cache[5][85] ), .A1N(n3839), .Y(\D_cache/n1111 ) );
  OAI2BB2XL U8605 ( .B0(\D_cache/n339 ), .B1(n3844), .A0N(
        \D_cache/cache[4][85] ), .A1N(n3862), .Y(\D_cache/n1112 ) );
  OAI2BB2XL U8606 ( .B0(\D_cache/n339 ), .B1(n3865), .A0N(
        \D_cache/cache[3][85] ), .A1N(n3881), .Y(\D_cache/n1113 ) );
  OAI2BB2XL U8607 ( .B0(\D_cache/n339 ), .B1(n3886), .A0N(
        \D_cache/cache[2][85] ), .A1N(n3902), .Y(\D_cache/n1114 ) );
  OAI2BB2XL U8608 ( .B0(\D_cache/n339 ), .B1(n3906), .A0N(
        \D_cache/cache[1][85] ), .A1N(n3923), .Y(\D_cache/n1115 ) );
  OAI2BB2XL U8609 ( .B0(\D_cache/n339 ), .B1(n3926), .A0N(
        \D_cache/cache[0][85] ), .A1N(n3944), .Y(\D_cache/n1116 ) );
  OAI2BB2XL U8610 ( .B0(\D_cache/n341 ), .B1(n3786), .A0N(
        \D_cache/cache[7][84] ), .A1N(n3802), .Y(\D_cache/n1117 ) );
  OAI2BB2XL U8611 ( .B0(\D_cache/n341 ), .B1(n3806), .A0N(
        \D_cache/cache[6][84] ), .A1N(n3822), .Y(\D_cache/n1118 ) );
  OAI2BB2XL U8612 ( .B0(\D_cache/n341 ), .B1(n3825), .A0N(
        \D_cache/cache[5][84] ), .A1N(n3839), .Y(\D_cache/n1119 ) );
  OAI2BB2XL U8613 ( .B0(\D_cache/n341 ), .B1(n3844), .A0N(
        \D_cache/cache[4][84] ), .A1N(n3862), .Y(\D_cache/n1120 ) );
  OAI2BB2XL U8614 ( .B0(\D_cache/n341 ), .B1(n3865), .A0N(
        \D_cache/cache[3][84] ), .A1N(n3881), .Y(\D_cache/n1121 ) );
  OAI2BB2XL U8615 ( .B0(\D_cache/n341 ), .B1(n3886), .A0N(
        \D_cache/cache[2][84] ), .A1N(n3902), .Y(\D_cache/n1122 ) );
  OAI2BB2XL U8616 ( .B0(\D_cache/n341 ), .B1(n3906), .A0N(
        \D_cache/cache[1][84] ), .A1N(n3923), .Y(\D_cache/n1123 ) );
  OAI2BB2XL U8617 ( .B0(\D_cache/n341 ), .B1(n3926), .A0N(
        \D_cache/cache[0][84] ), .A1N(n3944), .Y(\D_cache/n1124 ) );
  OAI2BB2XL U8618 ( .B0(\D_cache/n343 ), .B1(n3786), .A0N(
        \D_cache/cache[7][83] ), .A1N(n3801), .Y(\D_cache/n1125 ) );
  OAI2BB2XL U8619 ( .B0(\D_cache/n343 ), .B1(n3806), .A0N(
        \D_cache/cache[6][83] ), .A1N(n3821), .Y(\D_cache/n1126 ) );
  OAI2BB2XL U8620 ( .B0(\D_cache/n343 ), .B1(n3825), .A0N(
        \D_cache/cache[5][83] ), .A1N(n3838), .Y(\D_cache/n1127 ) );
  OAI2BB2XL U8621 ( .B0(\D_cache/n343 ), .B1(n3844), .A0N(
        \D_cache/cache[4][83] ), .A1N(n3861), .Y(\D_cache/n1128 ) );
  OAI2BB2XL U8622 ( .B0(\D_cache/n343 ), .B1(n3865), .A0N(
        \D_cache/cache[3][83] ), .A1N(n3880), .Y(\D_cache/n1129 ) );
  OAI2BB2XL U8623 ( .B0(\D_cache/n343 ), .B1(n3886), .A0N(
        \D_cache/cache[2][83] ), .A1N(n3901), .Y(\D_cache/n1130 ) );
  OAI2BB2XL U8624 ( .B0(\D_cache/n343 ), .B1(n3906), .A0N(
        \D_cache/cache[1][83] ), .A1N(n3922), .Y(\D_cache/n1131 ) );
  OAI2BB2XL U8625 ( .B0(\D_cache/n343 ), .B1(n3926), .A0N(
        \D_cache/cache[0][83] ), .A1N(n3943), .Y(\D_cache/n1132 ) );
  OAI2BB2XL U8626 ( .B0(\D_cache/n345 ), .B1(n3786), .A0N(
        \D_cache/cache[7][82] ), .A1N(n3801), .Y(\D_cache/n1133 ) );
  OAI2BB2XL U8627 ( .B0(\D_cache/n345 ), .B1(n3806), .A0N(
        \D_cache/cache[6][82] ), .A1N(n3821), .Y(\D_cache/n1134 ) );
  OAI2BB2XL U8628 ( .B0(\D_cache/n345 ), .B1(n3825), .A0N(
        \D_cache/cache[5][82] ), .A1N(n3838), .Y(\D_cache/n1135 ) );
  OAI2BB2XL U8629 ( .B0(\D_cache/n345 ), .B1(n3844), .A0N(
        \D_cache/cache[4][82] ), .A1N(n3861), .Y(\D_cache/n1136 ) );
  OAI2BB2XL U8630 ( .B0(\D_cache/n345 ), .B1(n3865), .A0N(
        \D_cache/cache[3][82] ), .A1N(n3880), .Y(\D_cache/n1137 ) );
  OAI2BB2XL U8631 ( .B0(\D_cache/n345 ), .B1(n3886), .A0N(
        \D_cache/cache[2][82] ), .A1N(n3901), .Y(\D_cache/n1138 ) );
  OAI2BB2XL U8632 ( .B0(\D_cache/n345 ), .B1(n3906), .A0N(
        \D_cache/cache[1][82] ), .A1N(n3922), .Y(\D_cache/n1139 ) );
  OAI2BB2XL U8633 ( .B0(\D_cache/n345 ), .B1(n3926), .A0N(
        \D_cache/cache[0][82] ), .A1N(n3943), .Y(\D_cache/n1140 ) );
  OAI2BB2XL U8634 ( .B0(\D_cache/n347 ), .B1(n3786), .A0N(
        \D_cache/cache[7][81] ), .A1N(n3801), .Y(\D_cache/n1141 ) );
  OAI2BB2XL U8635 ( .B0(\D_cache/n347 ), .B1(n3806), .A0N(
        \D_cache/cache[6][81] ), .A1N(n3821), .Y(\D_cache/n1142 ) );
  OAI2BB2XL U8636 ( .B0(\D_cache/n347 ), .B1(n3825), .A0N(
        \D_cache/cache[5][81] ), .A1N(n3838), .Y(\D_cache/n1143 ) );
  OAI2BB2XL U8637 ( .B0(\D_cache/n347 ), .B1(n3844), .A0N(
        \D_cache/cache[4][81] ), .A1N(n3861), .Y(\D_cache/n1144 ) );
  OAI2BB2XL U8638 ( .B0(\D_cache/n347 ), .B1(n3865), .A0N(
        \D_cache/cache[3][81] ), .A1N(n3880), .Y(\D_cache/n1145 ) );
  OAI2BB2XL U8639 ( .B0(\D_cache/n347 ), .B1(n3886), .A0N(
        \D_cache/cache[2][81] ), .A1N(n3901), .Y(\D_cache/n1146 ) );
  OAI2BB2XL U8640 ( .B0(\D_cache/n347 ), .B1(n3906), .A0N(
        \D_cache/cache[1][81] ), .A1N(n3922), .Y(\D_cache/n1147 ) );
  OAI2BB2XL U8641 ( .B0(\D_cache/n347 ), .B1(n3926), .A0N(
        \D_cache/cache[0][81] ), .A1N(n3943), .Y(\D_cache/n1148 ) );
  OAI2BB2XL U8642 ( .B0(\D_cache/n349 ), .B1(n3786), .A0N(
        \D_cache/cache[7][80] ), .A1N(n3801), .Y(\D_cache/n1149 ) );
  OAI2BB2XL U8643 ( .B0(\D_cache/n349 ), .B1(n3806), .A0N(
        \D_cache/cache[6][80] ), .A1N(n3821), .Y(\D_cache/n1150 ) );
  OAI2BB2XL U8644 ( .B0(\D_cache/n349 ), .B1(n3825), .A0N(
        \D_cache/cache[5][80] ), .A1N(n3838), .Y(\D_cache/n1151 ) );
  OAI2BB2XL U8645 ( .B0(\D_cache/n349 ), .B1(n3844), .A0N(
        \D_cache/cache[4][80] ), .A1N(n3861), .Y(\D_cache/n1152 ) );
  OAI2BB2XL U8646 ( .B0(\D_cache/n349 ), .B1(n3865), .A0N(
        \D_cache/cache[3][80] ), .A1N(n3880), .Y(\D_cache/n1153 ) );
  OAI2BB2XL U8647 ( .B0(\D_cache/n349 ), .B1(n3886), .A0N(
        \D_cache/cache[2][80] ), .A1N(n3901), .Y(\D_cache/n1154 ) );
  OAI2BB2XL U8648 ( .B0(\D_cache/n349 ), .B1(n3906), .A0N(
        \D_cache/cache[1][80] ), .A1N(n3922), .Y(\D_cache/n1155 ) );
  OAI2BB2XL U8649 ( .B0(\D_cache/n349 ), .B1(n3926), .A0N(
        \D_cache/cache[0][80] ), .A1N(n3943), .Y(\D_cache/n1156 ) );
  OAI2BB2XL U8650 ( .B0(\D_cache/n351 ), .B1(n3786), .A0N(
        \D_cache/cache[7][79] ), .A1N(n3801), .Y(\D_cache/n1157 ) );
  OAI2BB2XL U8651 ( .B0(\D_cache/n351 ), .B1(n3806), .A0N(
        \D_cache/cache[6][79] ), .A1N(n3821), .Y(\D_cache/n1158 ) );
  OAI2BB2XL U8652 ( .B0(\D_cache/n351 ), .B1(n3825), .A0N(
        \D_cache/cache[5][79] ), .A1N(n3838), .Y(\D_cache/n1159 ) );
  OAI2BB2XL U8653 ( .B0(\D_cache/n351 ), .B1(n3844), .A0N(
        \D_cache/cache[4][79] ), .A1N(n3861), .Y(\D_cache/n1160 ) );
  OAI2BB2XL U8654 ( .B0(\D_cache/n351 ), .B1(n3865), .A0N(
        \D_cache/cache[3][79] ), .A1N(n3880), .Y(\D_cache/n1161 ) );
  OAI2BB2XL U8655 ( .B0(\D_cache/n351 ), .B1(n3886), .A0N(
        \D_cache/cache[2][79] ), .A1N(n3901), .Y(\D_cache/n1162 ) );
  OAI2BB2XL U8656 ( .B0(\D_cache/n351 ), .B1(n3906), .A0N(
        \D_cache/cache[1][79] ), .A1N(n3922), .Y(\D_cache/n1163 ) );
  OAI2BB2XL U8657 ( .B0(\D_cache/n351 ), .B1(n3926), .A0N(
        \D_cache/cache[0][79] ), .A1N(n3943), .Y(\D_cache/n1164 ) );
  OAI2BB2XL U8658 ( .B0(\D_cache/n353 ), .B1(n3787), .A0N(
        \D_cache/cache[7][78] ), .A1N(n3801), .Y(\D_cache/n1165 ) );
  OAI2BB2XL U8659 ( .B0(\D_cache/n353 ), .B1(n3807), .A0N(
        \D_cache/cache[6][78] ), .A1N(n3821), .Y(\D_cache/n1166 ) );
  OAI2BB2XL U8660 ( .B0(\D_cache/n353 ), .B1(n3826), .A0N(
        \D_cache/cache[5][78] ), .A1N(n3838), .Y(\D_cache/n1167 ) );
  OAI2BB2XL U8661 ( .B0(\D_cache/n353 ), .B1(n3845), .A0N(
        \D_cache/cache[4][78] ), .A1N(n3861), .Y(\D_cache/n1168 ) );
  OAI2BB2XL U8662 ( .B0(\D_cache/n353 ), .B1(n3867), .A0N(
        \D_cache/cache[3][78] ), .A1N(n3880), .Y(\D_cache/n1169 ) );
  OAI2BB2XL U8663 ( .B0(\D_cache/n353 ), .B1(n3887), .A0N(
        \D_cache/cache[2][78] ), .A1N(n3901), .Y(\D_cache/n1170 ) );
  OAI2BB2XL U8664 ( .B0(\D_cache/n353 ), .B1(n3907), .A0N(
        \D_cache/cache[1][78] ), .A1N(n3922), .Y(\D_cache/n1171 ) );
  OAI2BB2XL U8665 ( .B0(\D_cache/n353 ), .B1(n3927), .A0N(
        \D_cache/cache[0][78] ), .A1N(n3943), .Y(\D_cache/n1172 ) );
  OAI2BB2XL U8666 ( .B0(\D_cache/n355 ), .B1(n3787), .A0N(
        \D_cache/cache[7][77] ), .A1N(n3801), .Y(\D_cache/n1173 ) );
  OAI2BB2XL U8667 ( .B0(\D_cache/n355 ), .B1(n3807), .A0N(
        \D_cache/cache[6][77] ), .A1N(n3821), .Y(\D_cache/n1174 ) );
  OAI2BB2XL U8668 ( .B0(\D_cache/n355 ), .B1(n3826), .A0N(
        \D_cache/cache[5][77] ), .A1N(n3838), .Y(\D_cache/n1175 ) );
  OAI2BB2XL U8669 ( .B0(\D_cache/n355 ), .B1(n3845), .A0N(
        \D_cache/cache[4][77] ), .A1N(n3861), .Y(\D_cache/n1176 ) );
  OAI2BB2XL U8670 ( .B0(\D_cache/n355 ), .B1(n3872), .A0N(
        \D_cache/cache[3][77] ), .A1N(n3880), .Y(\D_cache/n1177 ) );
  OAI2BB2XL U8671 ( .B0(\D_cache/n355 ), .B1(n3887), .A0N(
        \D_cache/cache[2][77] ), .A1N(n3901), .Y(\D_cache/n1178 ) );
  OAI2BB2XL U8672 ( .B0(\D_cache/n355 ), .B1(n3907), .A0N(
        \D_cache/cache[1][77] ), .A1N(n3922), .Y(\D_cache/n1179 ) );
  OAI2BB2XL U8673 ( .B0(\D_cache/n355 ), .B1(n3927), .A0N(
        \D_cache/cache[0][77] ), .A1N(n3943), .Y(\D_cache/n1180 ) );
  OAI2BB2XL U8674 ( .B0(\D_cache/n357 ), .B1(n3787), .A0N(
        \D_cache/cache[7][76] ), .A1N(n3801), .Y(\D_cache/n1181 ) );
  OAI2BB2XL U8675 ( .B0(\D_cache/n357 ), .B1(n3807), .A0N(
        \D_cache/cache[6][76] ), .A1N(n3821), .Y(\D_cache/n1182 ) );
  OAI2BB2XL U8676 ( .B0(\D_cache/n357 ), .B1(n3826), .A0N(
        \D_cache/cache[5][76] ), .A1N(n3838), .Y(\D_cache/n1183 ) );
  OAI2BB2XL U8677 ( .B0(\D_cache/n357 ), .B1(n3845), .A0N(
        \D_cache/cache[4][76] ), .A1N(n3861), .Y(\D_cache/n1184 ) );
  OAI2BB2XL U8678 ( .B0(\D_cache/n357 ), .B1(n3870), .A0N(
        \D_cache/cache[3][76] ), .A1N(n3880), .Y(\D_cache/n1185 ) );
  OAI2BB2XL U8679 ( .B0(\D_cache/n357 ), .B1(n3887), .A0N(
        \D_cache/cache[2][76] ), .A1N(n3901), .Y(\D_cache/n1186 ) );
  OAI2BB2XL U8680 ( .B0(\D_cache/n357 ), .B1(n3907), .A0N(
        \D_cache/cache[1][76] ), .A1N(n3922), .Y(\D_cache/n1187 ) );
  OAI2BB2XL U8681 ( .B0(\D_cache/n357 ), .B1(n3927), .A0N(
        \D_cache/cache[0][76] ), .A1N(n3943), .Y(\D_cache/n1188 ) );
  OAI2BB2XL U8682 ( .B0(\D_cache/n359 ), .B1(n3787), .A0N(
        \D_cache/cache[7][75] ), .A1N(n3801), .Y(\D_cache/n1189 ) );
  OAI2BB2XL U8683 ( .B0(\D_cache/n359 ), .B1(n3807), .A0N(
        \D_cache/cache[6][75] ), .A1N(n3821), .Y(\D_cache/n1190 ) );
  OAI2BB2XL U8684 ( .B0(\D_cache/n359 ), .B1(n3826), .A0N(
        \D_cache/cache[5][75] ), .A1N(n3838), .Y(\D_cache/n1191 ) );
  OAI2BB2XL U8685 ( .B0(\D_cache/n359 ), .B1(n3845), .A0N(
        \D_cache/cache[4][75] ), .A1N(n3861), .Y(\D_cache/n1192 ) );
  OAI2BB2XL U8686 ( .B0(\D_cache/n359 ), .B1(n3869), .A0N(
        \D_cache/cache[3][75] ), .A1N(n3880), .Y(\D_cache/n1193 ) );
  OAI2BB2XL U8687 ( .B0(\D_cache/n359 ), .B1(n3887), .A0N(
        \D_cache/cache[2][75] ), .A1N(n3901), .Y(\D_cache/n1194 ) );
  OAI2BB2XL U8688 ( .B0(\D_cache/n359 ), .B1(n3907), .A0N(
        \D_cache/cache[1][75] ), .A1N(n3922), .Y(\D_cache/n1195 ) );
  OAI2BB2XL U8689 ( .B0(\D_cache/n359 ), .B1(n3927), .A0N(
        \D_cache/cache[0][75] ), .A1N(n3943), .Y(\D_cache/n1196 ) );
  OAI2BB2XL U8690 ( .B0(\D_cache/n361 ), .B1(n3787), .A0N(
        \D_cache/cache[7][74] ), .A1N(n3801), .Y(\D_cache/n1197 ) );
  OAI2BB2XL U8691 ( .B0(\D_cache/n361 ), .B1(n3807), .A0N(
        \D_cache/cache[6][74] ), .A1N(n3821), .Y(\D_cache/n1198 ) );
  OAI2BB2XL U8692 ( .B0(\D_cache/n361 ), .B1(n3826), .A0N(
        \D_cache/cache[5][74] ), .A1N(n3838), .Y(\D_cache/n1199 ) );
  OAI2BB2XL U8693 ( .B0(\D_cache/n361 ), .B1(n3845), .A0N(
        \D_cache/cache[4][74] ), .A1N(n3861), .Y(\D_cache/n1200 ) );
  OAI2BB2XL U8694 ( .B0(\D_cache/n361 ), .B1(n3871), .A0N(
        \D_cache/cache[3][74] ), .A1N(n3880), .Y(\D_cache/n1201 ) );
  OAI2BB2XL U8695 ( .B0(\D_cache/n361 ), .B1(n3887), .A0N(
        \D_cache/cache[2][74] ), .A1N(n3901), .Y(\D_cache/n1202 ) );
  OAI2BB2XL U8696 ( .B0(\D_cache/n361 ), .B1(n3907), .A0N(
        \D_cache/cache[1][74] ), .A1N(n3922), .Y(\D_cache/n1203 ) );
  OAI2BB2XL U8697 ( .B0(\D_cache/n361 ), .B1(n3927), .A0N(
        \D_cache/cache[0][74] ), .A1N(n3943), .Y(\D_cache/n1204 ) );
  OAI2BB2XL U8698 ( .B0(\D_cache/n363 ), .B1(n3787), .A0N(
        \D_cache/cache[7][73] ), .A1N(n3801), .Y(\D_cache/n1205 ) );
  OAI2BB2XL U8699 ( .B0(\D_cache/n363 ), .B1(n3807), .A0N(
        \D_cache/cache[6][73] ), .A1N(n3821), .Y(\D_cache/n1206 ) );
  OAI2BB2XL U8700 ( .B0(\D_cache/n363 ), .B1(n3826), .A0N(
        \D_cache/cache[5][73] ), .A1N(n3838), .Y(\D_cache/n1207 ) );
  OAI2BB2XL U8701 ( .B0(\D_cache/n363 ), .B1(n3845), .A0N(
        \D_cache/cache[4][73] ), .A1N(n3861), .Y(\D_cache/n1208 ) );
  OAI2BB2XL U8702 ( .B0(\D_cache/n363 ), .B1(n3866), .A0N(
        \D_cache/cache[3][73] ), .A1N(n3880), .Y(\D_cache/n1209 ) );
  OAI2BB2XL U8703 ( .B0(\D_cache/n363 ), .B1(n3887), .A0N(
        \D_cache/cache[2][73] ), .A1N(n3901), .Y(\D_cache/n1210 ) );
  OAI2BB2XL U8704 ( .B0(\D_cache/n363 ), .B1(n3907), .A0N(
        \D_cache/cache[1][73] ), .A1N(n3922), .Y(\D_cache/n1211 ) );
  OAI2BB2XL U8705 ( .B0(\D_cache/n363 ), .B1(n3927), .A0N(
        \D_cache/cache[0][73] ), .A1N(n3943), .Y(\D_cache/n1212 ) );
  OAI2BB2XL U8706 ( .B0(\D_cache/n365 ), .B1(n3787), .A0N(
        \D_cache/cache[7][72] ), .A1N(n3801), .Y(\D_cache/n1213 ) );
  OAI2BB2XL U8707 ( .B0(\D_cache/n365 ), .B1(n3807), .A0N(
        \D_cache/cache[6][72] ), .A1N(n3821), .Y(\D_cache/n1214 ) );
  OAI2BB2XL U8708 ( .B0(\D_cache/n365 ), .B1(n3826), .A0N(
        \D_cache/cache[5][72] ), .A1N(n3838), .Y(\D_cache/n1215 ) );
  OAI2BB2XL U8709 ( .B0(\D_cache/n365 ), .B1(n3845), .A0N(
        \D_cache/cache[4][72] ), .A1N(n3861), .Y(\D_cache/n1216 ) );
  OAI2BB2XL U8710 ( .B0(\D_cache/n365 ), .B1(n3864), .A0N(
        \D_cache/cache[3][72] ), .A1N(n3880), .Y(\D_cache/n1217 ) );
  OAI2BB2XL U8711 ( .B0(\D_cache/n365 ), .B1(n3887), .A0N(
        \D_cache/cache[2][72] ), .A1N(n3901), .Y(\D_cache/n1218 ) );
  OAI2BB2XL U8712 ( .B0(\D_cache/n365 ), .B1(n3907), .A0N(
        \D_cache/cache[1][72] ), .A1N(n3922), .Y(\D_cache/n1219 ) );
  OAI2BB2XL U8713 ( .B0(\D_cache/n365 ), .B1(n3927), .A0N(
        \D_cache/cache[0][72] ), .A1N(n3943), .Y(\D_cache/n1220 ) );
  OAI2BB2XL U8714 ( .B0(\D_cache/n367 ), .B1(n3787), .A0N(
        \D_cache/cache[7][71] ), .A1N(n3801), .Y(\D_cache/n1221 ) );
  OAI2BB2XL U8715 ( .B0(\D_cache/n367 ), .B1(n3807), .A0N(
        \D_cache/cache[6][71] ), .A1N(n3821), .Y(\D_cache/n1222 ) );
  OAI2BB2XL U8716 ( .B0(\D_cache/n367 ), .B1(n3826), .A0N(
        \D_cache/cache[5][71] ), .A1N(n3838), .Y(\D_cache/n1223 ) );
  OAI2BB2XL U8717 ( .B0(\D_cache/n367 ), .B1(n3845), .A0N(
        \D_cache/cache[4][71] ), .A1N(n3861), .Y(\D_cache/n1224 ) );
  OAI2BB2XL U8718 ( .B0(\D_cache/n367 ), .B1(n3865), .A0N(
        \D_cache/cache[3][71] ), .A1N(n3880), .Y(\D_cache/n1225 ) );
  OAI2BB2XL U8719 ( .B0(\D_cache/n367 ), .B1(n3887), .A0N(
        \D_cache/cache[2][71] ), .A1N(n3901), .Y(\D_cache/n1226 ) );
  OAI2BB2XL U8720 ( .B0(\D_cache/n367 ), .B1(n3907), .A0N(
        \D_cache/cache[1][71] ), .A1N(n3922), .Y(\D_cache/n1227 ) );
  OAI2BB2XL U8721 ( .B0(\D_cache/n367 ), .B1(n3927), .A0N(
        \D_cache/cache[0][71] ), .A1N(n3943), .Y(\D_cache/n1228 ) );
  OAI2BB2XL U8722 ( .B0(\D_cache/n369 ), .B1(n3788), .A0N(
        \D_cache/cache[7][70] ), .A1N(n3801), .Y(\D_cache/n1229 ) );
  OAI2BB2XL U8723 ( .B0(\D_cache/n369 ), .B1(n3808), .A0N(
        \D_cache/cache[6][70] ), .A1N(n3821), .Y(\D_cache/n1230 ) );
  OAI2BB2XL U8724 ( .B0(\D_cache/n369 ), .B1(n3827), .A0N(
        \D_cache/cache[5][70] ), .A1N(n3838), .Y(\D_cache/n1231 ) );
  OAI2BB2XL U8725 ( .B0(\D_cache/n369 ), .B1(n3846), .A0N(
        \D_cache/cache[4][70] ), .A1N(n3861), .Y(\D_cache/n1232 ) );
  OAI2BB2XL U8726 ( .B0(\D_cache/n369 ), .B1(n3867), .A0N(
        \D_cache/cache[3][70] ), .A1N(n3880), .Y(\D_cache/n1233 ) );
  OAI2BB2XL U8727 ( .B0(\D_cache/n369 ), .B1(n3888), .A0N(
        \D_cache/cache[2][70] ), .A1N(n3901), .Y(\D_cache/n1234 ) );
  OAI2BB2XL U8728 ( .B0(\D_cache/n369 ), .B1(n3908), .A0N(
        \D_cache/cache[1][70] ), .A1N(n3922), .Y(\D_cache/n1235 ) );
  OAI2BB2XL U8729 ( .B0(\D_cache/n369 ), .B1(n3928), .A0N(
        \D_cache/cache[0][70] ), .A1N(n3943), .Y(\D_cache/n1236 ) );
  OAI2BB2XL U8730 ( .B0(\D_cache/n371 ), .B1(n3788), .A0N(
        \D_cache/cache[7][69] ), .A1N(n3801), .Y(\D_cache/n1237 ) );
  OAI2BB2XL U8731 ( .B0(\D_cache/n371 ), .B1(n3808), .A0N(
        \D_cache/cache[6][69] ), .A1N(n3821), .Y(\D_cache/n1238 ) );
  OAI2BB2XL U8732 ( .B0(\D_cache/n371 ), .B1(n3827), .A0N(
        \D_cache/cache[5][69] ), .A1N(n3838), .Y(\D_cache/n1239 ) );
  OAI2BB2XL U8733 ( .B0(\D_cache/n371 ), .B1(n3846), .A0N(
        \D_cache/cache[4][69] ), .A1N(n3861), .Y(\D_cache/n1240 ) );
  OAI2BB2XL U8734 ( .B0(\D_cache/n371 ), .B1(n3872), .A0N(
        \D_cache/cache[3][69] ), .A1N(n3880), .Y(\D_cache/n1241 ) );
  OAI2BB2XL U8735 ( .B0(\D_cache/n371 ), .B1(n3888), .A0N(
        \D_cache/cache[2][69] ), .A1N(n3901), .Y(\D_cache/n1242 ) );
  OAI2BB2XL U8736 ( .B0(\D_cache/n371 ), .B1(n3908), .A0N(
        \D_cache/cache[1][69] ), .A1N(n3922), .Y(\D_cache/n1243 ) );
  OAI2BB2XL U8737 ( .B0(\D_cache/n371 ), .B1(n3928), .A0N(
        \D_cache/cache[0][69] ), .A1N(n3943), .Y(\D_cache/n1244 ) );
  OAI2BB2XL U8738 ( .B0(\D_cache/n373 ), .B1(n3788), .A0N(
        \D_cache/cache[7][68] ), .A1N(n3801), .Y(\D_cache/n1245 ) );
  OAI2BB2XL U8739 ( .B0(\D_cache/n373 ), .B1(n3808), .A0N(
        \D_cache/cache[6][68] ), .A1N(n3821), .Y(\D_cache/n1246 ) );
  OAI2BB2XL U8740 ( .B0(\D_cache/n373 ), .B1(n3827), .A0N(
        \D_cache/cache[5][68] ), .A1N(n3838), .Y(\D_cache/n1247 ) );
  OAI2BB2XL U8741 ( .B0(\D_cache/n373 ), .B1(n3846), .A0N(
        \D_cache/cache[4][68] ), .A1N(n3861), .Y(\D_cache/n1248 ) );
  OAI2BB2XL U8742 ( .B0(\D_cache/n373 ), .B1(n3868), .A0N(
        \D_cache/cache[3][68] ), .A1N(n3880), .Y(\D_cache/n1249 ) );
  OAI2BB2XL U8743 ( .B0(\D_cache/n373 ), .B1(n3888), .A0N(
        \D_cache/cache[2][68] ), .A1N(n3901), .Y(\D_cache/n1250 ) );
  OAI2BB2XL U8744 ( .B0(\D_cache/n373 ), .B1(n3908), .A0N(
        \D_cache/cache[1][68] ), .A1N(n3922), .Y(\D_cache/n1251 ) );
  OAI2BB2XL U8745 ( .B0(\D_cache/n373 ), .B1(n3928), .A0N(
        \D_cache/cache[0][68] ), .A1N(n3943), .Y(\D_cache/n1252 ) );
  OAI2BB2XL U8746 ( .B0(\D_cache/n375 ), .B1(n3788), .A0N(
        \D_cache/cache[7][67] ), .A1N(n3801), .Y(\D_cache/n1253 ) );
  OAI2BB2XL U8747 ( .B0(\D_cache/n375 ), .B1(n3808), .A0N(
        \D_cache/cache[6][67] ), .A1N(n3821), .Y(\D_cache/n1254 ) );
  OAI2BB2XL U8748 ( .B0(\D_cache/n375 ), .B1(n3827), .A0N(
        \D_cache/cache[5][67] ), .A1N(n3838), .Y(\D_cache/n1255 ) );
  OAI2BB2XL U8749 ( .B0(\D_cache/n375 ), .B1(n3846), .A0N(
        \D_cache/cache[4][67] ), .A1N(n3861), .Y(\D_cache/n1256 ) );
  OAI2BB2XL U8750 ( .B0(\D_cache/n375 ), .B1(n3864), .A0N(
        \D_cache/cache[3][67] ), .A1N(n3880), .Y(\D_cache/n1257 ) );
  OAI2BB2XL U8751 ( .B0(\D_cache/n375 ), .B1(n3888), .A0N(
        \D_cache/cache[2][67] ), .A1N(n3901), .Y(\D_cache/n1258 ) );
  OAI2BB2XL U8752 ( .B0(\D_cache/n375 ), .B1(n3908), .A0N(
        \D_cache/cache[1][67] ), .A1N(n3922), .Y(\D_cache/n1259 ) );
  OAI2BB2XL U8753 ( .B0(\D_cache/n375 ), .B1(n3928), .A0N(
        \D_cache/cache[0][67] ), .A1N(n3943), .Y(\D_cache/n1260 ) );
  OAI2BB2XL U8754 ( .B0(\D_cache/n377 ), .B1(n3788), .A0N(
        \D_cache/cache[7][66] ), .A1N(n3801), .Y(\D_cache/n1261 ) );
  OAI2BB2XL U8755 ( .B0(\D_cache/n377 ), .B1(n3808), .A0N(
        \D_cache/cache[6][66] ), .A1N(n3821), .Y(\D_cache/n1262 ) );
  OAI2BB2XL U8756 ( .B0(\D_cache/n377 ), .B1(n3827), .A0N(
        \D_cache/cache[5][66] ), .A1N(n3838), .Y(\D_cache/n1263 ) );
  OAI2BB2XL U8757 ( .B0(\D_cache/n377 ), .B1(n3846), .A0N(
        \D_cache/cache[4][66] ), .A1N(n3861), .Y(\D_cache/n1264 ) );
  OAI2BB2XL U8758 ( .B0(\D_cache/n377 ), .B1(n3870), .A0N(
        \D_cache/cache[3][66] ), .A1N(n3880), .Y(\D_cache/n1265 ) );
  OAI2BB2XL U8759 ( .B0(\D_cache/n377 ), .B1(n3888), .A0N(
        \D_cache/cache[2][66] ), .A1N(n3901), .Y(\D_cache/n1266 ) );
  OAI2BB2XL U8760 ( .B0(\D_cache/n377 ), .B1(n3908), .A0N(
        \D_cache/cache[1][66] ), .A1N(n3922), .Y(\D_cache/n1267 ) );
  OAI2BB2XL U8761 ( .B0(\D_cache/n377 ), .B1(n3928), .A0N(
        \D_cache/cache[0][66] ), .A1N(n3943), .Y(\D_cache/n1268 ) );
  OAI2BB2XL U8762 ( .B0(\D_cache/n379 ), .B1(n3788), .A0N(
        \D_cache/cache[7][65] ), .A1N(n3801), .Y(\D_cache/n1269 ) );
  OAI2BB2XL U8763 ( .B0(\D_cache/n379 ), .B1(n3808), .A0N(
        \D_cache/cache[6][65] ), .A1N(n3821), .Y(\D_cache/n1270 ) );
  OAI2BB2XL U8764 ( .B0(\D_cache/n379 ), .B1(n3827), .A0N(
        \D_cache/cache[5][65] ), .A1N(n3838), .Y(\D_cache/n1271 ) );
  OAI2BB2XL U8765 ( .B0(\D_cache/n379 ), .B1(n3846), .A0N(
        \D_cache/cache[4][65] ), .A1N(n3861), .Y(\D_cache/n1272 ) );
  OAI2BB2XL U8766 ( .B0(\D_cache/n379 ), .B1(n3869), .A0N(
        \D_cache/cache[3][65] ), .A1N(n3880), .Y(\D_cache/n1273 ) );
  OAI2BB2XL U8767 ( .B0(\D_cache/n379 ), .B1(n3888), .A0N(
        \D_cache/cache[2][65] ), .A1N(n3901), .Y(\D_cache/n1274 ) );
  OAI2BB2XL U8768 ( .B0(\D_cache/n379 ), .B1(n3908), .A0N(
        \D_cache/cache[1][65] ), .A1N(n3922), .Y(\D_cache/n1275 ) );
  OAI2BB2XL U8769 ( .B0(\D_cache/n379 ), .B1(n3928), .A0N(
        \D_cache/cache[0][65] ), .A1N(n3943), .Y(\D_cache/n1276 ) );
  OAI2BB2XL U8770 ( .B0(\D_cache/n381 ), .B1(n3788), .A0N(
        \D_cache/cache[7][64] ), .A1N(n3800), .Y(\D_cache/n1277 ) );
  OAI2BB2XL U8771 ( .B0(\D_cache/n381 ), .B1(n3808), .A0N(
        \D_cache/cache[6][64] ), .A1N(n3820), .Y(\D_cache/n1278 ) );
  OAI2BB2XL U8772 ( .B0(\D_cache/n381 ), .B1(n3827), .A0N(
        \D_cache/cache[5][64] ), .A1N(n3827), .Y(\D_cache/n1279 ) );
  OAI2BB2XL U8773 ( .B0(\D_cache/n381 ), .B1(n3846), .A0N(
        \D_cache/cache[4][64] ), .A1N(n3860), .Y(\D_cache/n1280 ) );
  OAI2BB2XL U8774 ( .B0(\D_cache/n381 ), .B1(n3871), .A0N(
        \D_cache/cache[3][64] ), .A1N(n3879), .Y(\D_cache/n1281 ) );
  OAI2BB2XL U8775 ( .B0(\D_cache/n381 ), .B1(n3888), .A0N(
        \D_cache/cache[2][64] ), .A1N(n3900), .Y(\D_cache/n1282 ) );
  OAI2BB2XL U8776 ( .B0(\D_cache/n381 ), .B1(n3908), .A0N(
        \D_cache/cache[1][64] ), .A1N(n3921), .Y(\D_cache/n1283 ) );
  OAI2BB2XL U8777 ( .B0(\D_cache/n381 ), .B1(n3928), .A0N(
        \D_cache/cache[0][64] ), .A1N(n3942), .Y(\D_cache/n1284 ) );
  OAI2BB2XL U8778 ( .B0(\D_cache/n452 ), .B1(n3793), .A0N(
        \D_cache/cache[7][31] ), .A1N(n3799), .Y(\D_cache/n1541 ) );
  OAI2BB2XL U8779 ( .B0(\D_cache/n452 ), .B1(n3813), .A0N(
        \D_cache/cache[6][31] ), .A1N(n3819), .Y(\D_cache/n1542 ) );
  OAI2BB2XL U8780 ( .B0(\D_cache/n452 ), .B1(n3831), .A0N(
        \D_cache/cache[5][31] ), .A1N(n3837), .Y(\D_cache/n1543 ) );
  OAI2BB2XL U8781 ( .B0(\D_cache/n452 ), .B1(n3853), .A0N(
        \D_cache/cache[4][31] ), .A1N(n3859), .Y(\D_cache/n1544 ) );
  OAI2BB2XL U8782 ( .B0(\D_cache/n452 ), .B1(n3872), .A0N(
        \D_cache/cache[3][31] ), .A1N(n3878), .Y(\D_cache/n1545 ) );
  OAI2BB2XL U8783 ( .B0(\D_cache/n452 ), .B1(n3893), .A0N(
        \D_cache/cache[2][31] ), .A1N(n3899), .Y(\D_cache/n1546 ) );
  OAI2BB2XL U8784 ( .B0(\D_cache/n452 ), .B1(n3914), .A0N(
        \D_cache/cache[1][31] ), .A1N(n3920), .Y(\D_cache/n1547 ) );
  OAI2BB2XL U8785 ( .B0(\D_cache/n452 ), .B1(n3935), .A0N(
        \D_cache/cache[0][31] ), .A1N(n3941), .Y(\D_cache/n1548 ) );
  OAI2BB2XL U8786 ( .B0(\D_cache/n456 ), .B1(n3793), .A0N(
        \D_cache/cache[7][30] ), .A1N(n3799), .Y(\D_cache/n1549 ) );
  OAI2BB2XL U8787 ( .B0(\D_cache/n456 ), .B1(n3813), .A0N(
        \D_cache/cache[6][30] ), .A1N(n3819), .Y(\D_cache/n1550 ) );
  OAI2BB2XL U8788 ( .B0(\D_cache/n456 ), .B1(n3831), .A0N(
        \D_cache/cache[5][30] ), .A1N(n3837), .Y(\D_cache/n1551 ) );
  OAI2BB2XL U8789 ( .B0(\D_cache/n456 ), .B1(n3853), .A0N(
        \D_cache/cache[4][30] ), .A1N(n3859), .Y(\D_cache/n1552 ) );
  OAI2BB2XL U8790 ( .B0(\D_cache/n456 ), .B1(n3872), .A0N(
        \D_cache/cache[3][30] ), .A1N(n3878), .Y(\D_cache/n1553 ) );
  OAI2BB2XL U8791 ( .B0(\D_cache/n456 ), .B1(n3893), .A0N(
        \D_cache/cache[2][30] ), .A1N(n3899), .Y(\D_cache/n1554 ) );
  OAI2BB2XL U8792 ( .B0(\D_cache/n456 ), .B1(n3914), .A0N(
        \D_cache/cache[1][30] ), .A1N(n3920), .Y(\D_cache/n1555 ) );
  OAI2BB2XL U8793 ( .B0(\D_cache/n456 ), .B1(n3935), .A0N(
        \D_cache/cache[0][30] ), .A1N(n3941), .Y(\D_cache/n1556 ) );
  OAI2BB2XL U8794 ( .B0(\D_cache/n458 ), .B1(n3793), .A0N(
        \D_cache/cache[7][29] ), .A1N(n3799), .Y(\D_cache/n1557 ) );
  OAI2BB2XL U8795 ( .B0(\D_cache/n458 ), .B1(n3813), .A0N(
        \D_cache/cache[6][29] ), .A1N(n3819), .Y(\D_cache/n1558 ) );
  OAI2BB2XL U8796 ( .B0(\D_cache/n458 ), .B1(n3831), .A0N(
        \D_cache/cache[5][29] ), .A1N(n3837), .Y(\D_cache/n1559 ) );
  OAI2BB2XL U8797 ( .B0(\D_cache/n458 ), .B1(n3853), .A0N(
        \D_cache/cache[4][29] ), .A1N(n3859), .Y(\D_cache/n1560 ) );
  OAI2BB2XL U8798 ( .B0(\D_cache/n458 ), .B1(n3872), .A0N(
        \D_cache/cache[3][29] ), .A1N(n3878), .Y(\D_cache/n1561 ) );
  OAI2BB2XL U8799 ( .B0(\D_cache/n458 ), .B1(n3893), .A0N(
        \D_cache/cache[2][29] ), .A1N(n3899), .Y(\D_cache/n1562 ) );
  OAI2BB2XL U8800 ( .B0(\D_cache/n458 ), .B1(n3914), .A0N(
        \D_cache/cache[1][29] ), .A1N(n3920), .Y(\D_cache/n1563 ) );
  OAI2BB2XL U8801 ( .B0(\D_cache/n458 ), .B1(n3935), .A0N(
        \D_cache/cache[0][29] ), .A1N(n3941), .Y(\D_cache/n1564 ) );
  OAI2BB2XL U8802 ( .B0(\D_cache/n460 ), .B1(n3792), .A0N(
        \D_cache/cache[7][28] ), .A1N(n3799), .Y(\D_cache/n1565 ) );
  OAI2BB2XL U8803 ( .B0(\D_cache/n460 ), .B1(n3812), .A0N(
        \D_cache/cache[6][28] ), .A1N(n3819), .Y(\D_cache/n1566 ) );
  OAI2BB2XL U8804 ( .B0(\D_cache/n460 ), .B1(n3831), .A0N(
        \D_cache/cache[5][28] ), .A1N(n3837), .Y(\D_cache/n1567 ) );
  OAI2BB2XL U8805 ( .B0(\D_cache/n460 ), .B1(n3852), .A0N(
        \D_cache/cache[4][28] ), .A1N(n3859), .Y(\D_cache/n1568 ) );
  OAI2BB2XL U8806 ( .B0(\D_cache/n460 ), .B1(n3871), .A0N(
        \D_cache/cache[3][28] ), .A1N(n3878), .Y(\D_cache/n1569 ) );
  OAI2BB2XL U8807 ( .B0(\D_cache/n460 ), .B1(n3892), .A0N(
        \D_cache/cache[2][28] ), .A1N(n3899), .Y(\D_cache/n1570 ) );
  OAI2BB2XL U8808 ( .B0(\D_cache/n460 ), .B1(n3913), .A0N(
        \D_cache/cache[1][28] ), .A1N(n3920), .Y(\D_cache/n1571 ) );
  OAI2BB2XL U8809 ( .B0(\D_cache/n460 ), .B1(n3934), .A0N(
        \D_cache/cache[0][28] ), .A1N(n3941), .Y(\D_cache/n1572 ) );
  OAI2BB2XL U8810 ( .B0(\D_cache/n462 ), .B1(n3792), .A0N(
        \D_cache/cache[7][27] ), .A1N(n3798), .Y(\D_cache/n1573 ) );
  OAI2BB2XL U8811 ( .B0(\D_cache/n462 ), .B1(n3812), .A0N(
        \D_cache/cache[6][27] ), .A1N(n3818), .Y(\D_cache/n1574 ) );
  OAI2BB2XL U8812 ( .B0(\D_cache/n462 ), .B1(n3825), .A0N(
        \D_cache/cache[5][27] ), .A1N(n3836), .Y(\D_cache/n1575 ) );
  OAI2BB2XL U8813 ( .B0(\D_cache/n462 ), .B1(n3852), .A0N(
        \D_cache/cache[4][27] ), .A1N(n3858), .Y(\D_cache/n1576 ) );
  OAI2BB2XL U8814 ( .B0(\D_cache/n462 ), .B1(n3871), .A0N(
        \D_cache/cache[3][27] ), .A1N(n3877), .Y(\D_cache/n1577 ) );
  OAI2BB2XL U8815 ( .B0(\D_cache/n462 ), .B1(n3892), .A0N(
        \D_cache/cache[2][27] ), .A1N(n3898), .Y(\D_cache/n1578 ) );
  OAI2BB2XL U8816 ( .B0(\D_cache/n462 ), .B1(n3913), .A0N(
        \D_cache/cache[1][27] ), .A1N(n3919), .Y(\D_cache/n1579 ) );
  OAI2BB2XL U8817 ( .B0(\D_cache/n462 ), .B1(n3934), .A0N(
        \D_cache/cache[0][27] ), .A1N(n3940), .Y(\D_cache/n1580 ) );
  OAI2BB2XL U8818 ( .B0(\D_cache/n464 ), .B1(n3792), .A0N(
        \D_cache/cache[7][26] ), .A1N(n3798), .Y(\D_cache/n1581 ) );
  OAI2BB2XL U8819 ( .B0(\D_cache/n464 ), .B1(n3812), .A0N(
        \D_cache/cache[6][26] ), .A1N(n3818), .Y(\D_cache/n1582 ) );
  OAI2BB2XL U8820 ( .B0(\D_cache/n464 ), .B1(n3826), .A0N(
        \D_cache/cache[5][26] ), .A1N(n3836), .Y(\D_cache/n1583 ) );
  OAI2BB2XL U8821 ( .B0(\D_cache/n464 ), .B1(n3852), .A0N(
        \D_cache/cache[4][26] ), .A1N(n3858), .Y(\D_cache/n1584 ) );
  OAI2BB2XL U8822 ( .B0(\D_cache/n464 ), .B1(n3871), .A0N(
        \D_cache/cache[3][26] ), .A1N(n3877), .Y(\D_cache/n1585 ) );
  OAI2BB2XL U8823 ( .B0(\D_cache/n464 ), .B1(n3892), .A0N(
        \D_cache/cache[2][26] ), .A1N(n3898), .Y(\D_cache/n1586 ) );
  OAI2BB2XL U8824 ( .B0(\D_cache/n464 ), .B1(n3913), .A0N(
        \D_cache/cache[1][26] ), .A1N(n3919), .Y(\D_cache/n1587 ) );
  OAI2BB2XL U8825 ( .B0(\D_cache/n464 ), .B1(n3934), .A0N(
        \D_cache/cache[0][26] ), .A1N(n3940), .Y(\D_cache/n1588 ) );
  OAI2BB2XL U8826 ( .B0(\D_cache/n466 ), .B1(n3792), .A0N(
        \D_cache/cache[7][25] ), .A1N(n3798), .Y(\D_cache/n1589 ) );
  OAI2BB2XL U8827 ( .B0(\D_cache/n466 ), .B1(n3812), .A0N(
        \D_cache/cache[6][25] ), .A1N(n3818), .Y(\D_cache/n1590 ) );
  OAI2BB2XL U8828 ( .B0(\D_cache/n466 ), .B1(n3829), .A0N(
        \D_cache/cache[5][25] ), .A1N(n3836), .Y(\D_cache/n1591 ) );
  OAI2BB2XL U8829 ( .B0(\D_cache/n466 ), .B1(n3852), .A0N(
        \D_cache/cache[4][25] ), .A1N(n3858), .Y(\D_cache/n1592 ) );
  OAI2BB2XL U8830 ( .B0(\D_cache/n466 ), .B1(n3871), .A0N(
        \D_cache/cache[3][25] ), .A1N(n3877), .Y(\D_cache/n1593 ) );
  OAI2BB2XL U8831 ( .B0(\D_cache/n466 ), .B1(n3892), .A0N(
        \D_cache/cache[2][25] ), .A1N(n3898), .Y(\D_cache/n1594 ) );
  OAI2BB2XL U8832 ( .B0(\D_cache/n466 ), .B1(n3913), .A0N(
        \D_cache/cache[1][25] ), .A1N(n3919), .Y(\D_cache/n1595 ) );
  OAI2BB2XL U8833 ( .B0(\D_cache/n466 ), .B1(n3934), .A0N(
        \D_cache/cache[0][25] ), .A1N(n3940), .Y(\D_cache/n1596 ) );
  OAI2BB2XL U8834 ( .B0(\D_cache/n468 ), .B1(n3792), .A0N(
        \D_cache/cache[7][24] ), .A1N(n3798), .Y(\D_cache/n1597 ) );
  OAI2BB2XL U8835 ( .B0(\D_cache/n468 ), .B1(n3812), .A0N(
        \D_cache/cache[6][24] ), .A1N(n3818), .Y(\D_cache/n1598 ) );
  OAI2BB2XL U8836 ( .B0(\D_cache/n468 ), .B1(n3828), .A0N(
        \D_cache/cache[5][24] ), .A1N(n3836), .Y(\D_cache/n1599 ) );
  OAI2BB2XL U8837 ( .B0(\D_cache/n468 ), .B1(n3852), .A0N(
        \D_cache/cache[4][24] ), .A1N(n3858), .Y(\D_cache/n1600 ) );
  OAI2BB2XL U8838 ( .B0(\D_cache/n468 ), .B1(n3871), .A0N(
        \D_cache/cache[3][24] ), .A1N(n3877), .Y(\D_cache/n1601 ) );
  OAI2BB2XL U8839 ( .B0(\D_cache/n468 ), .B1(n3892), .A0N(
        \D_cache/cache[2][24] ), .A1N(n3898), .Y(\D_cache/n1602 ) );
  OAI2BB2XL U8840 ( .B0(\D_cache/n468 ), .B1(n3913), .A0N(
        \D_cache/cache[1][24] ), .A1N(n3919), .Y(\D_cache/n1603 ) );
  OAI2BB2XL U8841 ( .B0(\D_cache/n468 ), .B1(n3934), .A0N(
        \D_cache/cache[0][24] ), .A1N(n3940), .Y(\D_cache/n1604 ) );
  OAI2BB2XL U8842 ( .B0(\D_cache/n470 ), .B1(n3792), .A0N(
        \D_cache/cache[7][23] ), .A1N(n3798), .Y(\D_cache/n1605 ) );
  OAI2BB2XL U8843 ( .B0(\D_cache/n470 ), .B1(n3812), .A0N(
        \D_cache/cache[6][23] ), .A1N(n3818), .Y(\D_cache/n1606 ) );
  OAI2BB2XL U8844 ( .B0(\D_cache/n470 ), .B1(n3827), .A0N(
        \D_cache/cache[5][23] ), .A1N(n3836), .Y(\D_cache/n1607 ) );
  OAI2BB2XL U8845 ( .B0(\D_cache/n470 ), .B1(n3852), .A0N(
        \D_cache/cache[4][23] ), .A1N(n3858), .Y(\D_cache/n1608 ) );
  OAI2BB2XL U8846 ( .B0(\D_cache/n470 ), .B1(n3871), .A0N(
        \D_cache/cache[3][23] ), .A1N(n3877), .Y(\D_cache/n1609 ) );
  OAI2BB2XL U8847 ( .B0(\D_cache/n470 ), .B1(n3892), .A0N(
        \D_cache/cache[2][23] ), .A1N(n3898), .Y(\D_cache/n1610 ) );
  OAI2BB2XL U8848 ( .B0(\D_cache/n470 ), .B1(n3913), .A0N(
        \D_cache/cache[1][23] ), .A1N(n3919), .Y(\D_cache/n1611 ) );
  OAI2BB2XL U8849 ( .B0(\D_cache/n470 ), .B1(n3934), .A0N(
        \D_cache/cache[0][23] ), .A1N(n3940), .Y(\D_cache/n1612 ) );
  OAI2BB2XL U8850 ( .B0(\D_cache/n472 ), .B1(n3792), .A0N(
        \D_cache/cache[7][22] ), .A1N(n3798), .Y(\D_cache/n1613 ) );
  OAI2BB2XL U8851 ( .B0(\D_cache/n472 ), .B1(n3812), .A0N(
        \D_cache/cache[6][22] ), .A1N(n3818), .Y(\D_cache/n1614 ) );
  OAI2BB2XL U8852 ( .B0(\D_cache/n472 ), .B1(n3831), .A0N(
        \D_cache/cache[5][22] ), .A1N(n3836), .Y(\D_cache/n1615 ) );
  OAI2BB2XL U8853 ( .B0(\D_cache/n472 ), .B1(n3852), .A0N(
        \D_cache/cache[4][22] ), .A1N(n3858), .Y(\D_cache/n1616 ) );
  OAI2BB2XL U8854 ( .B0(\D_cache/n472 ), .B1(n3871), .A0N(
        \D_cache/cache[3][22] ), .A1N(n3877), .Y(\D_cache/n1617 ) );
  OAI2BB2XL U8855 ( .B0(\D_cache/n472 ), .B1(n3892), .A0N(
        \D_cache/cache[2][22] ), .A1N(n3898), .Y(\D_cache/n1618 ) );
  OAI2BB2XL U8856 ( .B0(\D_cache/n472 ), .B1(n3913), .A0N(
        \D_cache/cache[1][22] ), .A1N(n3919), .Y(\D_cache/n1619 ) );
  OAI2BB2XL U8857 ( .B0(\D_cache/n472 ), .B1(n3934), .A0N(
        \D_cache/cache[0][22] ), .A1N(n3940), .Y(\D_cache/n1620 ) );
  OAI2BB2XL U8858 ( .B0(\D_cache/n474 ), .B1(n3792), .A0N(
        \D_cache/cache[7][21] ), .A1N(n3798), .Y(\D_cache/n1621 ) );
  OAI2BB2XL U8859 ( .B0(\D_cache/n474 ), .B1(n3812), .A0N(
        \D_cache/cache[6][21] ), .A1N(n3818), .Y(\D_cache/n1622 ) );
  OAI2BB2XL U8860 ( .B0(\D_cache/n474 ), .B1(n3825), .A0N(
        \D_cache/cache[5][21] ), .A1N(n3836), .Y(\D_cache/n1623 ) );
  OAI2BB2XL U8861 ( .B0(\D_cache/n474 ), .B1(n3852), .A0N(
        \D_cache/cache[4][21] ), .A1N(n3858), .Y(\D_cache/n1624 ) );
  OAI2BB2XL U8862 ( .B0(\D_cache/n474 ), .B1(n3871), .A0N(
        \D_cache/cache[3][21] ), .A1N(n3877), .Y(\D_cache/n1625 ) );
  OAI2BB2XL U8863 ( .B0(\D_cache/n474 ), .B1(n3892), .A0N(
        \D_cache/cache[2][21] ), .A1N(n3898), .Y(\D_cache/n1626 ) );
  OAI2BB2XL U8864 ( .B0(\D_cache/n474 ), .B1(n3913), .A0N(
        \D_cache/cache[1][21] ), .A1N(n3919), .Y(\D_cache/n1627 ) );
  OAI2BB2XL U8865 ( .B0(\D_cache/n474 ), .B1(n3934), .A0N(
        \D_cache/cache[0][21] ), .A1N(n3940), .Y(\D_cache/n1628 ) );
  OAI2BB2XL U8866 ( .B0(\D_cache/n476 ), .B1(n3791), .A0N(
        \D_cache/cache[7][20] ), .A1N(n3798), .Y(\D_cache/n1629 ) );
  OAI2BB2XL U8867 ( .B0(\D_cache/n476 ), .B1(n3811), .A0N(
        \D_cache/cache[6][20] ), .A1N(n3818), .Y(\D_cache/n1630 ) );
  OAI2BB2XL U8868 ( .B0(\D_cache/n476 ), .B1(n3830), .A0N(
        \D_cache/cache[5][20] ), .A1N(n3836), .Y(\D_cache/n1631 ) );
  OAI2BB2XL U8869 ( .B0(\D_cache/n476 ), .B1(n3851), .A0N(
        \D_cache/cache[4][20] ), .A1N(n3858), .Y(\D_cache/n1632 ) );
  OAI2BB2XL U8870 ( .B0(\D_cache/n476 ), .B1(n3870), .A0N(
        \D_cache/cache[3][20] ), .A1N(n3877), .Y(\D_cache/n1633 ) );
  OAI2BB2XL U8871 ( .B0(\D_cache/n476 ), .B1(n3891), .A0N(
        \D_cache/cache[2][20] ), .A1N(n3898), .Y(\D_cache/n1634 ) );
  OAI2BB2XL U8872 ( .B0(\D_cache/n476 ), .B1(n3911), .A0N(
        \D_cache/cache[1][20] ), .A1N(n3919), .Y(\D_cache/n1635 ) );
  OAI2BB2XL U8873 ( .B0(\D_cache/n476 ), .B1(n3933), .A0N(
        \D_cache/cache[0][20] ), .A1N(n3940), .Y(\D_cache/n1636 ) );
  OAI2BB2XL U8874 ( .B0(\D_cache/n478 ), .B1(n3786), .A0N(
        \D_cache/cache[7][19] ), .A1N(n3798), .Y(\D_cache/n1637 ) );
  OAI2BB2XL U8875 ( .B0(\D_cache/n478 ), .B1(n3806), .A0N(
        \D_cache/cache[6][19] ), .A1N(n3818), .Y(\D_cache/n1638 ) );
  OAI2BB2XL U8876 ( .B0(\D_cache/n478 ), .B1(n3830), .A0N(
        \D_cache/cache[5][19] ), .A1N(n3836), .Y(\D_cache/n1639 ) );
  OAI2BB2XL U8877 ( .B0(\D_cache/n478 ), .B1(n3851), .A0N(
        \D_cache/cache[4][19] ), .A1N(n3858), .Y(\D_cache/n1640 ) );
  OAI2BB2XL U8878 ( .B0(\D_cache/n478 ), .B1(n3870), .A0N(
        \D_cache/cache[3][19] ), .A1N(n3877), .Y(\D_cache/n1641 ) );
  OAI2BB2XL U8879 ( .B0(\D_cache/n478 ), .B1(n3886), .A0N(
        \D_cache/cache[2][19] ), .A1N(n3898), .Y(\D_cache/n1642 ) );
  OAI2BB2XL U8880 ( .B0(\D_cache/n478 ), .B1(n3906), .A0N(
        \D_cache/cache[1][19] ), .A1N(n3919), .Y(\D_cache/n1643 ) );
  OAI2BB2XL U8881 ( .B0(\D_cache/n478 ), .B1(n3933), .A0N(
        \D_cache/cache[0][19] ), .A1N(n3940), .Y(\D_cache/n1644 ) );
  OAI2BB2XL U8882 ( .B0(\D_cache/n480 ), .B1(n3785), .A0N(
        \D_cache/cache[7][18] ), .A1N(n3798), .Y(\D_cache/n1645 ) );
  OAI2BB2XL U8883 ( .B0(\D_cache/n480 ), .B1(n3805), .A0N(
        \D_cache/cache[6][18] ), .A1N(n3818), .Y(\D_cache/n1646 ) );
  OAI2BB2XL U8884 ( .B0(\D_cache/n480 ), .B1(n3830), .A0N(
        \D_cache/cache[5][18] ), .A1N(n3836), .Y(\D_cache/n1647 ) );
  OAI2BB2XL U8885 ( .B0(\D_cache/n480 ), .B1(n3851), .A0N(
        \D_cache/cache[4][18] ), .A1N(n3858), .Y(\D_cache/n1648 ) );
  OAI2BB2XL U8886 ( .B0(\D_cache/n480 ), .B1(n3870), .A0N(
        \D_cache/cache[3][18] ), .A1N(n3877), .Y(\D_cache/n1649 ) );
  OAI2BB2XL U8887 ( .B0(\D_cache/n480 ), .B1(n3885), .A0N(
        \D_cache/cache[2][18] ), .A1N(n3898), .Y(\D_cache/n1650 ) );
  OAI2BB2XL U8888 ( .B0(\D_cache/n480 ), .B1(n3905), .A0N(
        \D_cache/cache[1][18] ), .A1N(n3919), .Y(\D_cache/n1651 ) );
  OAI2BB2XL U8889 ( .B0(\D_cache/n480 ), .B1(n3933), .A0N(
        \D_cache/cache[0][18] ), .A1N(n3940), .Y(\D_cache/n1652 ) );
  OAI2BB2XL U8890 ( .B0(\D_cache/n482 ), .B1(n3791), .A0N(
        \D_cache/cache[7][17] ), .A1N(n3798), .Y(\D_cache/n1653 ) );
  OAI2BB2XL U8891 ( .B0(\D_cache/n482 ), .B1(n3811), .A0N(
        \D_cache/cache[6][17] ), .A1N(n3818), .Y(\D_cache/n1654 ) );
  OAI2BB2XL U8892 ( .B0(\D_cache/n482 ), .B1(n3830), .A0N(
        \D_cache/cache[5][17] ), .A1N(n3836), .Y(\D_cache/n1655 ) );
  OAI2BB2XL U8893 ( .B0(\D_cache/n482 ), .B1(n3851), .A0N(
        \D_cache/cache[4][17] ), .A1N(n3858), .Y(\D_cache/n1656 ) );
  OAI2BB2XL U8894 ( .B0(\D_cache/n482 ), .B1(n3870), .A0N(
        \D_cache/cache[3][17] ), .A1N(n3877), .Y(\D_cache/n1657 ) );
  OAI2BB2XL U8895 ( .B0(\D_cache/n482 ), .B1(n3891), .A0N(
        \D_cache/cache[2][17] ), .A1N(n3898), .Y(\D_cache/n1658 ) );
  OAI2BB2XL U8896 ( .B0(\D_cache/n482 ), .B1(n3911), .A0N(
        \D_cache/cache[1][17] ), .A1N(n3919), .Y(\D_cache/n1659 ) );
  OAI2BB2XL U8897 ( .B0(\D_cache/n482 ), .B1(n3933), .A0N(
        \D_cache/cache[0][17] ), .A1N(n3940), .Y(\D_cache/n1660 ) );
  OAI2BB2XL U8898 ( .B0(\D_cache/n484 ), .B1(n3786), .A0N(
        \D_cache/cache[7][16] ), .A1N(n3798), .Y(\D_cache/n1661 ) );
  OAI2BB2XL U8899 ( .B0(\D_cache/n484 ), .B1(n3806), .A0N(
        \D_cache/cache[6][16] ), .A1N(n3818), .Y(\D_cache/n1662 ) );
  OAI2BB2XL U8900 ( .B0(\D_cache/n484 ), .B1(n3830), .A0N(
        \D_cache/cache[5][16] ), .A1N(n3836), .Y(\D_cache/n1663 ) );
  OAI2BB2XL U8901 ( .B0(\D_cache/n484 ), .B1(n3851), .A0N(
        \D_cache/cache[4][16] ), .A1N(n3858), .Y(\D_cache/n1664 ) );
  OAI2BB2XL U8902 ( .B0(\D_cache/n484 ), .B1(n3870), .A0N(
        \D_cache/cache[3][16] ), .A1N(n3877), .Y(\D_cache/n1665 ) );
  OAI2BB2XL U8903 ( .B0(\D_cache/n484 ), .B1(n3886), .A0N(
        \D_cache/cache[2][16] ), .A1N(n3898), .Y(\D_cache/n1666 ) );
  OAI2BB2XL U8904 ( .B0(\D_cache/n484 ), .B1(n3906), .A0N(
        \D_cache/cache[1][16] ), .A1N(n3919), .Y(\D_cache/n1667 ) );
  OAI2BB2XL U8905 ( .B0(\D_cache/n484 ), .B1(n3933), .A0N(
        \D_cache/cache[0][16] ), .A1N(n3940), .Y(\D_cache/n1668 ) );
  OAI2BB2XL U8906 ( .B0(\D_cache/n486 ), .B1(n3785), .A0N(
        \D_cache/cache[7][15] ), .A1N(n3798), .Y(\D_cache/n1669 ) );
  OAI2BB2XL U8907 ( .B0(\D_cache/n486 ), .B1(n3805), .A0N(
        \D_cache/cache[6][15] ), .A1N(n3818), .Y(\D_cache/n1670 ) );
  OAI2BB2XL U8908 ( .B0(\D_cache/n486 ), .B1(n3830), .A0N(
        \D_cache/cache[5][15] ), .A1N(n3836), .Y(\D_cache/n1671 ) );
  OAI2BB2XL U8909 ( .B0(\D_cache/n486 ), .B1(n3851), .A0N(
        \D_cache/cache[4][15] ), .A1N(n3858), .Y(\D_cache/n1672 ) );
  OAI2BB2XL U8910 ( .B0(\D_cache/n486 ), .B1(n3870), .A0N(
        \D_cache/cache[3][15] ), .A1N(n3877), .Y(\D_cache/n1673 ) );
  OAI2BB2XL U8911 ( .B0(\D_cache/n486 ), .B1(n3885), .A0N(
        \D_cache/cache[2][15] ), .A1N(n3898), .Y(\D_cache/n1674 ) );
  OAI2BB2XL U8912 ( .B0(\D_cache/n486 ), .B1(n3905), .A0N(
        \D_cache/cache[1][15] ), .A1N(n3919), .Y(\D_cache/n1675 ) );
  OAI2BB2XL U8913 ( .B0(\D_cache/n486 ), .B1(n3933), .A0N(
        \D_cache/cache[0][15] ), .A1N(n3940), .Y(\D_cache/n1676 ) );
  OAI2BB2XL U8914 ( .B0(\D_cache/n488 ), .B1(n3791), .A0N(
        \D_cache/cache[7][14] ), .A1N(n3798), .Y(\D_cache/n1677 ) );
  OAI2BB2XL U8915 ( .B0(\D_cache/n488 ), .B1(n3811), .A0N(
        \D_cache/cache[6][14] ), .A1N(n3818), .Y(\D_cache/n1678 ) );
  OAI2BB2XL U8916 ( .B0(\D_cache/n488 ), .B1(n3830), .A0N(
        \D_cache/cache[5][14] ), .A1N(n3836), .Y(\D_cache/n1679 ) );
  OAI2BB2XL U8917 ( .B0(\D_cache/n488 ), .B1(n3851), .A0N(
        \D_cache/cache[4][14] ), .A1N(n3858), .Y(\D_cache/n1680 ) );
  OAI2BB2XL U8918 ( .B0(\D_cache/n488 ), .B1(n3870), .A0N(
        \D_cache/cache[3][14] ), .A1N(n3877), .Y(\D_cache/n1681 ) );
  OAI2BB2XL U8919 ( .B0(\D_cache/n488 ), .B1(n3891), .A0N(
        \D_cache/cache[2][14] ), .A1N(n3898), .Y(\D_cache/n1682 ) );
  OAI2BB2XL U8920 ( .B0(\D_cache/n488 ), .B1(n3911), .A0N(
        \D_cache/cache[1][14] ), .A1N(n3919), .Y(\D_cache/n1683 ) );
  OAI2BB2XL U8921 ( .B0(\D_cache/n488 ), .B1(n3933), .A0N(
        \D_cache/cache[0][14] ), .A1N(n3940), .Y(\D_cache/n1684 ) );
  OAI2BB2XL U8922 ( .B0(\D_cache/n490 ), .B1(n3786), .A0N(
        \D_cache/cache[7][13] ), .A1N(n3798), .Y(\D_cache/n1685 ) );
  OAI2BB2XL U8923 ( .B0(\D_cache/n490 ), .B1(n3806), .A0N(
        \D_cache/cache[6][13] ), .A1N(n3818), .Y(\D_cache/n1686 ) );
  OAI2BB2XL U8924 ( .B0(\D_cache/n490 ), .B1(n3830), .A0N(
        \D_cache/cache[5][13] ), .A1N(n3836), .Y(\D_cache/n1687 ) );
  OAI2BB2XL U8925 ( .B0(\D_cache/n490 ), .B1(n3851), .A0N(
        \D_cache/cache[4][13] ), .A1N(n3858), .Y(\D_cache/n1688 ) );
  OAI2BB2XL U8926 ( .B0(\D_cache/n490 ), .B1(n3870), .A0N(
        \D_cache/cache[3][13] ), .A1N(n3877), .Y(\D_cache/n1689 ) );
  OAI2BB2XL U8927 ( .B0(\D_cache/n490 ), .B1(n3886), .A0N(
        \D_cache/cache[2][13] ), .A1N(n3898), .Y(\D_cache/n1690 ) );
  OAI2BB2XL U8928 ( .B0(\D_cache/n490 ), .B1(n3906), .A0N(
        \D_cache/cache[1][13] ), .A1N(n3919), .Y(\D_cache/n1691 ) );
  OAI2BB2XL U8929 ( .B0(\D_cache/n490 ), .B1(n3933), .A0N(
        \D_cache/cache[0][13] ), .A1N(n3940), .Y(\D_cache/n1692 ) );
  OAI2BB2XL U8930 ( .B0(\D_cache/n492 ), .B1(n3791), .A0N(
        \D_cache/cache[7][12] ), .A1N(n3798), .Y(\D_cache/n1693 ) );
  OAI2BB2XL U8931 ( .B0(\D_cache/n492 ), .B1(n3811), .A0N(
        \D_cache/cache[6][12] ), .A1N(n3818), .Y(\D_cache/n1694 ) );
  OAI2BB2XL U8932 ( .B0(\D_cache/n492 ), .B1(n3827), .A0N(
        \D_cache/cache[5][12] ), .A1N(n3836), .Y(\D_cache/n1695 ) );
  OAI2BB2XL U8933 ( .B0(\D_cache/n492 ), .B1(n3850), .A0N(
        \D_cache/cache[4][12] ), .A1N(n3858), .Y(\D_cache/n1696 ) );
  OAI2BB2XL U8934 ( .B0(\D_cache/n492 ), .B1(n3869), .A0N(
        \D_cache/cache[3][12] ), .A1N(n3877), .Y(\D_cache/n1697 ) );
  OAI2BB2XL U8935 ( .B0(\D_cache/n492 ), .B1(n3891), .A0N(
        \D_cache/cache[2][12] ), .A1N(n3898), .Y(\D_cache/n1698 ) );
  OAI2BB2XL U8936 ( .B0(\D_cache/n492 ), .B1(n3912), .A0N(
        \D_cache/cache[1][12] ), .A1N(n3919), .Y(\D_cache/n1699 ) );
  OAI2BB2XL U8937 ( .B0(\D_cache/n492 ), .B1(n3932), .A0N(
        \D_cache/cache[0][12] ), .A1N(n3940), .Y(\D_cache/n1700 ) );
  OAI2BB2XL U8938 ( .B0(\D_cache/n494 ), .B1(n3786), .A0N(
        \D_cache/cache[7][11] ), .A1N(n3798), .Y(\D_cache/n1701 ) );
  OAI2BB2XL U8939 ( .B0(\D_cache/n494 ), .B1(n3806), .A0N(
        \D_cache/cache[6][11] ), .A1N(n3818), .Y(\D_cache/n1702 ) );
  OAI2BB2XL U8940 ( .B0(\D_cache/n494 ), .B1(n3831), .A0N(
        \D_cache/cache[5][11] ), .A1N(n3836), .Y(\D_cache/n1703 ) );
  OAI2BB2XL U8941 ( .B0(\D_cache/n494 ), .B1(n3850), .A0N(
        \D_cache/cache[4][11] ), .A1N(n3858), .Y(\D_cache/n1704 ) );
  OAI2BB2XL U8942 ( .B0(\D_cache/n494 ), .B1(n3869), .A0N(
        \D_cache/cache[3][11] ), .A1N(n3877), .Y(\D_cache/n1705 ) );
  OAI2BB2XL U8943 ( .B0(\D_cache/n494 ), .B1(n3886), .A0N(
        \D_cache/cache[2][11] ), .A1N(n3898), .Y(\D_cache/n1706 ) );
  OAI2BB2XL U8944 ( .B0(\D_cache/n494 ), .B1(n3912), .A0N(
        \D_cache/cache[1][11] ), .A1N(n3919), .Y(\D_cache/n1707 ) );
  OAI2BB2XL U8945 ( .B0(\D_cache/n494 ), .B1(n3932), .A0N(
        \D_cache/cache[0][11] ), .A1N(n3940), .Y(\D_cache/n1708 ) );
  OAI2BB2XL U8946 ( .B0(\D_cache/n496 ), .B1(n3785), .A0N(
        \D_cache/cache[7][10] ), .A1N(n3798), .Y(\D_cache/n1709 ) );
  OAI2BB2XL U8947 ( .B0(\D_cache/n496 ), .B1(n3805), .A0N(
        \D_cache/cache[6][10] ), .A1N(n3818), .Y(\D_cache/n1710 ) );
  OAI2BB2XL U8948 ( .B0(\D_cache/n496 ), .B1(n3826), .A0N(
        \D_cache/cache[5][10] ), .A1N(n3836), .Y(\D_cache/n1711 ) );
  OAI2BB2XL U8949 ( .B0(\D_cache/n496 ), .B1(n3850), .A0N(
        \D_cache/cache[4][10] ), .A1N(n3858), .Y(\D_cache/n1712 ) );
  OAI2BB2XL U8950 ( .B0(\D_cache/n496 ), .B1(n3869), .A0N(
        \D_cache/cache[3][10] ), .A1N(n3877), .Y(\D_cache/n1713 ) );
  OAI2BB2XL U8951 ( .B0(\D_cache/n496 ), .B1(n3885), .A0N(
        \D_cache/cache[2][10] ), .A1N(n3898), .Y(\D_cache/n1714 ) );
  OAI2BB2XL U8952 ( .B0(\D_cache/n496 ), .B1(n3912), .A0N(
        \D_cache/cache[1][10] ), .A1N(n3919), .Y(\D_cache/n1715 ) );
  OAI2BB2XL U8953 ( .B0(\D_cache/n496 ), .B1(n3932), .A0N(
        \D_cache/cache[0][10] ), .A1N(n3940), .Y(\D_cache/n1716 ) );
  OAI2BB2XL U8954 ( .B0(\D_cache/n498 ), .B1(n3791), .A0N(
        \D_cache/cache[7][9] ), .A1N(n3798), .Y(\D_cache/n1717 ) );
  OAI2BB2XL U8955 ( .B0(\D_cache/n498 ), .B1(n3811), .A0N(
        \D_cache/cache[6][9] ), .A1N(n3818), .Y(\D_cache/n1718 ) );
  OAI2BB2XL U8956 ( .B0(\D_cache/n498 ), .B1(n3830), .A0N(
        \D_cache/cache[5][9] ), .A1N(n3836), .Y(\D_cache/n1719 ) );
  OAI2BB2XL U8957 ( .B0(\D_cache/n498 ), .B1(n3850), .A0N(
        \D_cache/cache[4][9] ), .A1N(n3858), .Y(\D_cache/n1720 ) );
  OAI2BB2XL U8958 ( .B0(\D_cache/n498 ), .B1(n3869), .A0N(
        \D_cache/cache[3][9] ), .A1N(n3877), .Y(\D_cache/n1721 ) );
  OAI2BB2XL U8959 ( .B0(\D_cache/n498 ), .B1(n3891), .A0N(
        \D_cache/cache[2][9] ), .A1N(n3898), .Y(\D_cache/n1722 ) );
  OAI2BB2XL U8960 ( .B0(\D_cache/n498 ), .B1(n3912), .A0N(
        \D_cache/cache[1][9] ), .A1N(n3919), .Y(\D_cache/n1723 ) );
  OAI2BB2XL U8961 ( .B0(\D_cache/n498 ), .B1(n3932), .A0N(
        \D_cache/cache[0][9] ), .A1N(n3940), .Y(\D_cache/n1724 ) );
  OAI2BB2XL U8962 ( .B0(\D_cache/n500 ), .B1(n3786), .A0N(
        \D_cache/cache[7][8] ), .A1N(n3797), .Y(\D_cache/n1725 ) );
  OAI2BB2XL U8963 ( .B0(\D_cache/n500 ), .B1(n3806), .A0N(
        \D_cache/cache[6][8] ), .A1N(n3817), .Y(\D_cache/n1726 ) );
  OAI2BB2XL U8964 ( .B0(\D_cache/n500 ), .B1(n3829), .A0N(
        \D_cache/cache[5][8] ), .A1N(n3835), .Y(\D_cache/n1727 ) );
  OAI2BB2XL U8965 ( .B0(\D_cache/n500 ), .B1(n3850), .A0N(
        \D_cache/cache[4][8] ), .A1N(n3857), .Y(\D_cache/n1728 ) );
  OAI2BB2XL U8966 ( .B0(\D_cache/n500 ), .B1(n3869), .A0N(
        \D_cache/cache[3][8] ), .A1N(n3876), .Y(\D_cache/n1729 ) );
  OAI2BB2XL U8967 ( .B0(\D_cache/n500 ), .B1(n3886), .A0N(
        \D_cache/cache[2][8] ), .A1N(n3897), .Y(\D_cache/n1730 ) );
  OAI2BB2XL U8968 ( .B0(\D_cache/n500 ), .B1(n3912), .A0N(
        \D_cache/cache[1][8] ), .A1N(n3918), .Y(\D_cache/n1731 ) );
  OAI2BB2XL U8969 ( .B0(\D_cache/n500 ), .B1(n3932), .A0N(
        \D_cache/cache[0][8] ), .A1N(n3939), .Y(\D_cache/n1732 ) );
  OAI2BB2XL U8970 ( .B0(\D_cache/n502 ), .B1(n3785), .A0N(
        \D_cache/cache[7][7] ), .A1N(n3797), .Y(\D_cache/n1733 ) );
  OAI2BB2XL U8971 ( .B0(\D_cache/n502 ), .B1(n3805), .A0N(
        \D_cache/cache[6][7] ), .A1N(n3817), .Y(\D_cache/n1734 ) );
  OAI2BB2XL U8972 ( .B0(\D_cache/n502 ), .B1(n3828), .A0N(
        \D_cache/cache[5][7] ), .A1N(n3835), .Y(\D_cache/n1735 ) );
  OAI2BB2XL U8973 ( .B0(\D_cache/n502 ), .B1(n3850), .A0N(
        \D_cache/cache[4][7] ), .A1N(n3857), .Y(\D_cache/n1736 ) );
  OAI2BB2XL U8974 ( .B0(\D_cache/n502 ), .B1(n3869), .A0N(
        \D_cache/cache[3][7] ), .A1N(n3876), .Y(\D_cache/n1737 ) );
  OAI2BB2XL U8975 ( .B0(\D_cache/n502 ), .B1(n3885), .A0N(
        \D_cache/cache[2][7] ), .A1N(n3897), .Y(\D_cache/n1738 ) );
  OAI2BB2XL U8976 ( .B0(\D_cache/n502 ), .B1(n3912), .A0N(
        \D_cache/cache[1][7] ), .A1N(n3918), .Y(\D_cache/n1739 ) );
  OAI2BB2XL U8977 ( .B0(\D_cache/n502 ), .B1(n3932), .A0N(
        \D_cache/cache[0][7] ), .A1N(n3939), .Y(\D_cache/n1740 ) );
  OAI2BB2XL U8978 ( .B0(\D_cache/n504 ), .B1(n3791), .A0N(
        \D_cache/cache[7][6] ), .A1N(n3797), .Y(\D_cache/n1741 ) );
  OAI2BB2XL U8979 ( .B0(\D_cache/n504 ), .B1(n3811), .A0N(
        \D_cache/cache[6][6] ), .A1N(n3817), .Y(\D_cache/n1742 ) );
  OAI2BB2XL U8980 ( .B0(\D_cache/n504 ), .B1(n3825), .A0N(
        \D_cache/cache[5][6] ), .A1N(n3835), .Y(\D_cache/n1743 ) );
  OAI2BB2XL U8981 ( .B0(\D_cache/n504 ), .B1(n3850), .A0N(
        \D_cache/cache[4][6] ), .A1N(n3857), .Y(\D_cache/n1744 ) );
  OAI2BB2XL U8982 ( .B0(\D_cache/n504 ), .B1(n3869), .A0N(
        \D_cache/cache[3][6] ), .A1N(n3876), .Y(\D_cache/n1745 ) );
  OAI2BB2XL U8983 ( .B0(\D_cache/n504 ), .B1(n3891), .A0N(
        \D_cache/cache[2][6] ), .A1N(n3897), .Y(\D_cache/n1746 ) );
  OAI2BB2XL U8984 ( .B0(\D_cache/n504 ), .B1(n3912), .A0N(
        \D_cache/cache[1][6] ), .A1N(n3918), .Y(\D_cache/n1747 ) );
  OAI2BB2XL U8985 ( .B0(\D_cache/n504 ), .B1(n3932), .A0N(
        \D_cache/cache[0][6] ), .A1N(n3939), .Y(\D_cache/n1748 ) );
  OAI2BB2XL U8986 ( .B0(\D_cache/n506 ), .B1(n3786), .A0N(
        \D_cache/cache[7][5] ), .A1N(n3797), .Y(\D_cache/n1749 ) );
  OAI2BB2XL U8987 ( .B0(\D_cache/n506 ), .B1(n3806), .A0N(
        \D_cache/cache[6][5] ), .A1N(n3817), .Y(\D_cache/n1750 ) );
  OAI2BB2XL U8988 ( .B0(\D_cache/n506 ), .B1(n3827), .A0N(
        \D_cache/cache[5][5] ), .A1N(n3835), .Y(\D_cache/n1751 ) );
  OAI2BB2XL U8989 ( .B0(\D_cache/n506 ), .B1(n3850), .A0N(
        \D_cache/cache[4][5] ), .A1N(n3857), .Y(\D_cache/n1752 ) );
  OAI2BB2XL U8990 ( .B0(\D_cache/n506 ), .B1(n3869), .A0N(
        \D_cache/cache[3][5] ), .A1N(n3876), .Y(\D_cache/n1753 ) );
  OAI2BB2XL U8991 ( .B0(\D_cache/n506 ), .B1(n3886), .A0N(
        \D_cache/cache[2][5] ), .A1N(n3897), .Y(\D_cache/n1754 ) );
  OAI2BB2XL U8992 ( .B0(\D_cache/n506 ), .B1(n3912), .A0N(
        \D_cache/cache[1][5] ), .A1N(n3918), .Y(\D_cache/n1755 ) );
  OAI2BB2XL U8993 ( .B0(\D_cache/n506 ), .B1(n3932), .A0N(
        \D_cache/cache[0][5] ), .A1N(n3939), .Y(\D_cache/n1756 ) );
  OAI2BB2XL U8994 ( .B0(\D_cache/n508 ), .B1(n3791), .A0N(
        \D_cache/cache[7][4] ), .A1N(n3797), .Y(\D_cache/n1757 ) );
  OAI2BB2XL U8995 ( .B0(\D_cache/n508 ), .B1(n3811), .A0N(
        \D_cache/cache[6][4] ), .A1N(n3817), .Y(\D_cache/n1758 ) );
  OAI2BB2XL U8996 ( .B0(\D_cache/n508 ), .B1(n3829), .A0N(
        \D_cache/cache[5][4] ), .A1N(n3835), .Y(\D_cache/n1759 ) );
  OAI2BB2XL U8997 ( .B0(\D_cache/n508 ), .B1(n3849), .A0N(
        \D_cache/cache[4][4] ), .A1N(n3857), .Y(\D_cache/n1760 ) );
  OAI2BB2XL U8998 ( .B0(\D_cache/n508 ), .B1(n3868), .A0N(
        \D_cache/cache[3][4] ), .A1N(n3876), .Y(\D_cache/n1761 ) );
  OAI2BB2XL U8999 ( .B0(\D_cache/n508 ), .B1(n3891), .A0N(
        \D_cache/cache[2][4] ), .A1N(n3897), .Y(\D_cache/n1762 ) );
  OAI2BB2XL U9000 ( .B0(\D_cache/n508 ), .B1(n3911), .A0N(
        \D_cache/cache[1][4] ), .A1N(n3918), .Y(\D_cache/n1763 ) );
  OAI2BB2XL U9001 ( .B0(\D_cache/n508 ), .B1(n3931), .A0N(
        \D_cache/cache[0][4] ), .A1N(n3939), .Y(\D_cache/n1764 ) );
  OAI2BB2XL U9002 ( .B0(\D_cache/n510 ), .B1(n3791), .A0N(
        \D_cache/cache[7][3] ), .A1N(n3797), .Y(\D_cache/n1765 ) );
  OAI2BB2XL U9003 ( .B0(\D_cache/n510 ), .B1(n3811), .A0N(
        \D_cache/cache[6][3] ), .A1N(n3817), .Y(\D_cache/n1766 ) );
  OAI2BB2XL U9004 ( .B0(\D_cache/n510 ), .B1(n3829), .A0N(
        \D_cache/cache[5][3] ), .A1N(n3835), .Y(\D_cache/n1767 ) );
  OAI2BB2XL U9005 ( .B0(\D_cache/n510 ), .B1(n3849), .A0N(
        \D_cache/cache[4][3] ), .A1N(n3857), .Y(\D_cache/n1768 ) );
  OAI2BB2XL U9006 ( .B0(\D_cache/n510 ), .B1(n3868), .A0N(
        \D_cache/cache[3][3] ), .A1N(n3876), .Y(\D_cache/n1769 ) );
  OAI2BB2XL U9007 ( .B0(\D_cache/n510 ), .B1(n3891), .A0N(
        \D_cache/cache[2][3] ), .A1N(n3897), .Y(\D_cache/n1770 ) );
  OAI2BB2XL U9008 ( .B0(\D_cache/n510 ), .B1(n3911), .A0N(
        \D_cache/cache[1][3] ), .A1N(n3918), .Y(\D_cache/n1771 ) );
  OAI2BB2XL U9009 ( .B0(\D_cache/n510 ), .B1(n3931), .A0N(
        \D_cache/cache[0][3] ), .A1N(n3939), .Y(\D_cache/n1772 ) );
  OAI2BB2XL U9010 ( .B0(\D_cache/n512 ), .B1(n3791), .A0N(
        \D_cache/cache[7][2] ), .A1N(n3800), .Y(\D_cache/n1773 ) );
  OAI2BB2XL U9011 ( .B0(\D_cache/n512 ), .B1(n3811), .A0N(
        \D_cache/cache[6][2] ), .A1N(n3820), .Y(\D_cache/n1774 ) );
  OAI2BB2XL U9012 ( .B0(\D_cache/n512 ), .B1(n3829), .A0N(
        \D_cache/cache[5][2] ), .A1N(n3831), .Y(\D_cache/n1775 ) );
  OAI2BB2XL U9013 ( .B0(\D_cache/n512 ), .B1(n3849), .A0N(
        \D_cache/cache[4][2] ), .A1N(n3860), .Y(\D_cache/n1776 ) );
  OAI2BB2XL U9014 ( .B0(\D_cache/n512 ), .B1(n3868), .A0N(
        \D_cache/cache[3][2] ), .A1N(n3879), .Y(\D_cache/n1777 ) );
  OAI2BB2XL U9015 ( .B0(\D_cache/n512 ), .B1(n3891), .A0N(
        \D_cache/cache[2][2] ), .A1N(n3900), .Y(\D_cache/n1778 ) );
  OAI2BB2XL U9016 ( .B0(\D_cache/n512 ), .B1(n3911), .A0N(
        \D_cache/cache[1][2] ), .A1N(n3921), .Y(\D_cache/n1779 ) );
  OAI2BB2XL U9017 ( .B0(\D_cache/n512 ), .B1(n3931), .A0N(
        \D_cache/cache[0][2] ), .A1N(n3942), .Y(\D_cache/n1780 ) );
  OAI2BB2XL U9018 ( .B0(\D_cache/n514 ), .B1(n3791), .A0N(
        \D_cache/cache[7][1] ), .A1N(n3797), .Y(\D_cache/n1781 ) );
  OAI2BB2XL U9019 ( .B0(\D_cache/n514 ), .B1(n3811), .A0N(
        \D_cache/cache[6][1] ), .A1N(n3817), .Y(\D_cache/n1782 ) );
  OAI2BB2XL U9020 ( .B0(\D_cache/n514 ), .B1(n3829), .A0N(
        \D_cache/cache[5][1] ), .A1N(n3835), .Y(\D_cache/n1783 ) );
  OAI2BB2XL U9021 ( .B0(\D_cache/n514 ), .B1(n3849), .A0N(
        \D_cache/cache[4][1] ), .A1N(n3857), .Y(\D_cache/n1784 ) );
  OAI2BB2XL U9022 ( .B0(\D_cache/n514 ), .B1(n3868), .A0N(
        \D_cache/cache[3][1] ), .A1N(n3876), .Y(\D_cache/n1785 ) );
  OAI2BB2XL U9023 ( .B0(\D_cache/n514 ), .B1(n3891), .A0N(
        \D_cache/cache[2][1] ), .A1N(n3897), .Y(\D_cache/n1786 ) );
  OAI2BB2XL U9024 ( .B0(\D_cache/n514 ), .B1(n3911), .A0N(
        \D_cache/cache[1][1] ), .A1N(n3918), .Y(\D_cache/n1787 ) );
  OAI2BB2XL U9025 ( .B0(\D_cache/n514 ), .B1(n3931), .A0N(
        \D_cache/cache[0][1] ), .A1N(n3939), .Y(\D_cache/n1788 ) );
  OAI2BB2XL U9026 ( .B0(\D_cache/n516 ), .B1(n3792), .A0N(
        \D_cache/cache[7][0] ), .A1N(n3797), .Y(\D_cache/n1796 ) );
  OAI2BB2XL U9027 ( .B0(\D_cache/n516 ), .B1(n3812), .A0N(
        \D_cache/cache[6][0] ), .A1N(n3817), .Y(\D_cache/n1789 ) );
  OAI2BB2XL U9028 ( .B0(\D_cache/n516 ), .B1(n3826), .A0N(
        \D_cache/cache[5][0] ), .A1N(n3835), .Y(\D_cache/n1790 ) );
  OAI2BB2XL U9029 ( .B0(\D_cache/n516 ), .B1(n3852), .A0N(
        \D_cache/cache[4][0] ), .A1N(n3857), .Y(\D_cache/n1791 ) );
  OAI2BB2XL U9030 ( .B0(\D_cache/n516 ), .B1(n3871), .A0N(
        \D_cache/cache[3][0] ), .A1N(n3876), .Y(\D_cache/n1792 ) );
  OAI2BB2XL U9031 ( .B0(\D_cache/n516 ), .B1(n3892), .A0N(
        \D_cache/cache[2][0] ), .A1N(n3897), .Y(\D_cache/n1793 ) );
  OAI2BB2XL U9032 ( .B0(\D_cache/n516 ), .B1(n3913), .A0N(
        \D_cache/cache[1][0] ), .A1N(n3918), .Y(\D_cache/n1794 ) );
  OAI2BB2XL U9033 ( .B0(\D_cache/n516 ), .B1(n3934), .A0N(
        \D_cache/cache[0][0] ), .A1N(n3939), .Y(\D_cache/n1795 ) );
  AOI2BB2X1 U9034 ( .B0(\i_MIPS/IF_ID[92] ), .B1(n2157), .A0N(n3595), .A1N(
        \i_MIPS/n207 ), .Y(n8204) );
  OA22X1 U9035 ( .A0(n8202), .A1(n3599), .B0(n2158), .B1(n8267), .Y(n8203) );
  AOI2BB2X1 U9036 ( .B0(\i_MIPS/IF_ID[88] ), .B1(n2157), .A0N(n3595), .A1N(
        \i_MIPS/n203 ), .Y(n8097) );
  AOI2BB2X1 U9037 ( .B0(\i_MIPS/IF_ID[84] ), .B1(n2157), .A0N(n3594), .A1N(
        \i_MIPS/n199 ), .Y(n8034) );
  AOI2BB2X1 U9038 ( .B0(\i_MIPS/IF_ID[83] ), .B1(n2157), .A0N(n3594), .A1N(
        \i_MIPS/n198 ), .Y(n8007) );
  OA22X1 U9039 ( .A0(n8005), .A1(n3598), .B0(n2158), .B1(n8025), .Y(n8006) );
  AOI2BB2X1 U9040 ( .B0(\i_MIPS/IF_ID[82] ), .B1(n2157), .A0N(n3594), .A1N(
        \i_MIPS/n197 ), .Y(n7992) );
  OA22X1 U9041 ( .A0(n3580), .A1(n3598), .B0(n2158), .B1(n7996), .Y(n7991) );
  AOI2BB2X1 U9042 ( .B0(\i_MIPS/IF_ID[80] ), .B1(n2157), .A0N(n3594), .A1N(
        \i_MIPS/n195 ), .Y(n7961) );
  OA22X1 U9043 ( .A0(n7966), .A1(n3598), .B0(n2158), .B1(n7965), .Y(n7960) );
  AOI2BB2X1 U9044 ( .B0(\i_MIPS/IF_ID[79] ), .B1(n2157), .A0N(n3594), .A1N(
        \i_MIPS/n194 ), .Y(n7941) );
  OA22X1 U9045 ( .A0(n7945), .A1(n3598), .B0(n2158), .B1(n7944), .Y(n7940) );
  AOI2BB2X1 U9046 ( .B0(\i_MIPS/IF_ID[78] ), .B1(n2157), .A0N(n3594), .A1N(
        \i_MIPS/n193 ), .Y(n7926) );
  OA22X1 U9047 ( .A0(n7931), .A1(n3598), .B0(n2158), .B1(n7930), .Y(n7925) );
  AOI2BB2X1 U9048 ( .B0(\i_MIPS/IF_ID[76] ), .B1(n2157), .A0N(n3594), .A1N(
        \i_MIPS/n191 ), .Y(n7906) );
  OA22X1 U9049 ( .A0(n7915), .A1(n3598), .B0(n2158), .B1(n7914), .Y(n7905) );
  AOI2BB2X1 U9050 ( .B0(\i_MIPS/IF_ID[75] ), .B1(n2157), .A0N(n3594), .A1N(
        \i_MIPS/n190 ), .Y(n7890) );
  OA22X1 U9051 ( .A0(n7896), .A1(n3598), .B0(n2158), .B1(n7895), .Y(n7889) );
  AOI2BB2X1 U9052 ( .B0(\i_MIPS/IF_ID[74] ), .B1(n2157), .A0N(n3594), .A1N(
        \i_MIPS/n189 ), .Y(n7878) );
  OA22X1 U9053 ( .A0(n7849), .A1(n3598), .B0(n2158), .B1(n7848), .Y(n7843) );
  AOI33X1 U9054 ( .A0(\i_MIPS/Hazard_detection/n7 ), .A1(n7085), .A2(n7084), 
        .B0(\i_MIPS/Hazard_detection/n4 ), .B1(n7083), .B2(n7082), .Y(n7086)
         );
  OAI2BB2XL U9055 ( .B0(n3030), .B1(n3759), .A0N(
        \i_MIPS/Register/register[7][5] ), .A1N(n3761), .Y(
        \i_MIPS/Register/n889 ) );
  OAI2BB2XL U9056 ( .B0(n3030), .B1(n3756), .A0N(
        \i_MIPS/Register/register[8][5] ), .A1N(n3758), .Y(
        \i_MIPS/Register/n857 ) );
  OAI2BB2XL U9057 ( .B0(n3030), .B1(n3753), .A0N(
        \i_MIPS/Register/register[9][5] ), .A1N(n3755), .Y(
        \i_MIPS/Register/n825 ) );
  OAI2BB2XL U9058 ( .B0(n3030), .B1(n3750), .A0N(
        \i_MIPS/Register/register[10][5] ), .A1N(n3752), .Y(
        \i_MIPS/Register/n793 ) );
  OAI2BB2XL U9059 ( .B0(n3030), .B1(n3747), .A0N(
        \i_MIPS/Register/register[11][5] ), .A1N(n3749), .Y(
        \i_MIPS/Register/n761 ) );
  OAI2BB2XL U9060 ( .B0(n3030), .B1(n3744), .A0N(
        \i_MIPS/Register/register[12][5] ), .A1N(n3746), .Y(
        \i_MIPS/Register/n729 ) );
  OAI2BB2XL U9061 ( .B0(n3030), .B1(n3741), .A0N(
        \i_MIPS/Register/register[13][5] ), .A1N(n3743), .Y(
        \i_MIPS/Register/n697 ) );
  OAI2BB2XL U9062 ( .B0(n3030), .B1(n3738), .A0N(
        \i_MIPS/Register/register[14][5] ), .A1N(n3740), .Y(
        \i_MIPS/Register/n665 ) );
  OAI2BB2XL U9063 ( .B0(n3030), .B1(n3735), .A0N(
        \i_MIPS/Register/register[15][5] ), .A1N(n3737), .Y(
        \i_MIPS/Register/n633 ) );
  OAI2BB2XL U9064 ( .B0(n3030), .B1(n3732), .A0N(
        \i_MIPS/Register/register[16][5] ), .A1N(n3734), .Y(
        \i_MIPS/Register/n601 ) );
  OAI2BB2XL U9065 ( .B0(n3030), .B1(n3729), .A0N(
        \i_MIPS/Register/register[17][5] ), .A1N(n3731), .Y(
        \i_MIPS/Register/n569 ) );
  OAI2BB2XL U9066 ( .B0(n3679), .B1(n3726), .A0N(
        \i_MIPS/Register/register[18][5] ), .A1N(n3728), .Y(
        \i_MIPS/Register/n537 ) );
  OAI2BB2XL U9067 ( .B0(n3679), .B1(n3723), .A0N(
        \i_MIPS/Register/register[19][5] ), .A1N(n3725), .Y(
        \i_MIPS/Register/n505 ) );
  OAI2BB2XL U9068 ( .B0(n3679), .B1(n3720), .A0N(
        \i_MIPS/Register/register[20][5] ), .A1N(n3722), .Y(
        \i_MIPS/Register/n473 ) );
  OAI2BB2XL U9069 ( .B0(n3679), .B1(n3717), .A0N(
        \i_MIPS/Register/register[21][5] ), .A1N(n3719), .Y(
        \i_MIPS/Register/n441 ) );
  OAI2BB2XL U9070 ( .B0(n3679), .B1(n3714), .A0N(
        \i_MIPS/Register/register[22][5] ), .A1N(n3716), .Y(
        \i_MIPS/Register/n409 ) );
  OAI2BB2XL U9071 ( .B0(n3679), .B1(n3711), .A0N(
        \i_MIPS/Register/register[23][5] ), .A1N(n3713), .Y(
        \i_MIPS/Register/n377 ) );
  OAI2BB2XL U9072 ( .B0(n3679), .B1(n3708), .A0N(
        \i_MIPS/Register/register[24][5] ), .A1N(n3710), .Y(
        \i_MIPS/Register/n345 ) );
  OAI2BB2XL U9073 ( .B0(n3679), .B1(n3705), .A0N(
        \i_MIPS/Register/register[25][5] ), .A1N(n3707), .Y(
        \i_MIPS/Register/n313 ) );
  OAI2BB2XL U9074 ( .B0(n3679), .B1(n3702), .A0N(
        \i_MIPS/Register/register[26][5] ), .A1N(n3704), .Y(
        \i_MIPS/Register/n281 ) );
  OAI2BB2XL U9075 ( .B0(n3679), .B1(n3699), .A0N(
        \i_MIPS/Register/register[27][5] ), .A1N(n3701), .Y(
        \i_MIPS/Register/n249 ) );
  OAI2BB2XL U9076 ( .B0(n3679), .B1(n3696), .A0N(
        \i_MIPS/Register/register[28][5] ), .A1N(n3698), .Y(
        \i_MIPS/Register/n217 ) );
  OAI2BB2XL U9077 ( .B0(n3679), .B1(n3693), .A0N(
        \i_MIPS/Register/register[29][5] ), .A1N(n3695), .Y(
        \i_MIPS/Register/n185 ) );
  OAI2BB2XL U9078 ( .B0(n3030), .B1(n3690), .A0N(
        \i_MIPS/Register/register[30][5] ), .A1N(n3692), .Y(
        \i_MIPS/Register/n153 ) );
  OAI21XL U9079 ( .A0(\i_MIPS/n180 ), .A1(n3613), .B0(n8261), .Y(\i_MIPS/N23 )
         );
  OAI21XL U9080 ( .A0(\i_MIPS/n181 ), .A1(n3611), .B0(n8238), .Y(\i_MIPS/N24 )
         );
  OAI21XL U9081 ( .A0(\i_MIPS/n234 ), .A1(n3610), .B0(n8261), .Y(\i_MIPS/N88 )
         );
  XOR2X1 U9082 ( .A(n7964), .B(ICACHE_addr[14]), .Y(n7982) );
  XOR2X1 U9083 ( .A(n7917), .B(ICACHE_addr[10]), .Y(n8216) );
  CLKXOR2X2 U9084 ( .A(n8041), .B(ICACHE_addr[18]), .Y(n8051) );
  AOI2BB2X1 U9085 ( .B0(\i_MIPS/IF_ID[85] ), .B1(n2157), .A0N(n3595), .A1N(
        \i_MIPS/n200 ), .Y(n8054) );
  OA22X1 U9086 ( .A0(n8052), .A1(n3598), .B0(n2158), .B1(n8051), .Y(n8053) );
  AOI2BB2X1 U9087 ( .B0(\i_MIPS/IF_ID[81] ), .B1(n2157), .A0N(n3594), .A1N(
        \i_MIPS/n196 ), .Y(n7974) );
  OA22X1 U9088 ( .A0(n7983), .A1(n3598), .B0(n2158), .B1(n7982), .Y(n7973) );
  OA22X2 U9089 ( .A0(n3462), .A1(n170), .B0(n3415), .B1(n1067), .Y(n4517) );
  NAND3X4 U9090 ( .A(n4419), .B(n4418), .C(n4417), .Y(n4431) );
  NOR2X4 U9091 ( .A(n4402), .B(n4401), .Y(n4419) );
  AOI2BB2X1 U9092 ( .B0(\i_MIPS/IF_ID[73] ), .B1(n2157), .A0N(n3594), .A1N(
        \i_MIPS/n188 ), .Y(n7859) );
  OA22X1 U9093 ( .A0(n7867), .A1(n3598), .B0(n2158), .B1(n7866), .Y(n7858) );
  AOI2BB2X1 U9094 ( .B0(\i_MIPS/IF_ID[91] ), .B1(n2157), .A0N(n3595), .A1N(
        \i_MIPS/n206 ), .Y(n8183) );
  AOI2BB2X1 U9095 ( .B0(\i_MIPS/IF_ID[87] ), .B1(n2157), .A0N(n3595), .A1N(
        \i_MIPS/n202 ), .Y(n8078) );
  AOI2BB2X1 U9096 ( .B0(\i_MIPS/IF_ID[89] ), .B1(n2157), .A0N(n3595), .A1N(
        \i_MIPS/n204 ), .Y(n8140) );
  AND2X2 U9097 ( .A(\i_MIPS/ID_EX[80] ), .B(n54), .Y(n2907) );
  OA22X2 U9098 ( .A0(n3462), .A1(n171), .B0(n3415), .B1(n1068), .Y(n4521) );
  AOI2BB2X1 U9099 ( .B0(\i_MIPS/IF_ID[86] ), .B1(n2157), .A0N(n3595), .A1N(
        \i_MIPS/n201 ), .Y(n8424) );
  AND3X2 U9100 ( .A(n2888), .B(n964), .C(n4608), .Y(n4609) );
  OA22X1 U9101 ( .A0(n3550), .A1(n521), .B0(n3509), .B1(n1439), .Y(n4564) );
  OA22X1 U9102 ( .A0(n3550), .A1(n522), .B0(n3509), .B1(n1440), .Y(n4554) );
  OA22X1 U9103 ( .A0(n3554), .A1(n691), .B0(n3512), .B1(n1612), .Y(n7367) );
  OA22X1 U9104 ( .A0(n3555), .A1(n692), .B0(n3513), .B1(n1613), .Y(n7375) );
  OA22X1 U9105 ( .A0(n3555), .A1(n693), .B0(n3513), .B1(n1614), .Y(n7379) );
  OA22X1 U9106 ( .A0(n3555), .A1(n694), .B0(n3513), .B1(n1615), .Y(n7371) );
  OA22X1 U9107 ( .A0(n3473), .A1(n523), .B0(n3426), .B1(n1441), .Y(n7551) );
  OA22X1 U9108 ( .A0(n3472), .A1(n524), .B0(n3425), .B1(n1442), .Y(n7546) );
  OA22X1 U9109 ( .A0(n3467), .A1(n525), .B0(n3420), .B1(n1443), .Y(n7324) );
  AOI2BB2X1 U9110 ( .B0(\i_MIPS/IF_ID[90] ), .B1(n2157), .A0N(n3595), .A1N(
        \i_MIPS/n205 ), .Y(n8156) );
  OAI221X1 U9111 ( .A0(\D_cache/n164 ), .A1(n8859), .B0(n3074), .B1(n8840), 
        .C0(\D_cache/n197 ), .Y(DCACHE_rdata[11]) );
  CLKINVX1 U9112 ( .A(\i_MIPS/n316 ), .Y(n7164) );
  CLKINVX1 U9113 ( .A(\i_MIPS/n314 ), .Y(n7091) );
  XOR2X1 U9114 ( .A(\i_MIPS/PC/n4 ), .B(ICACHE_addr[1]), .Y(n8340) );
  XOR2X1 U9115 ( .A(n7847), .B(ICACHE_addr[6]), .Y(n7866) );
  XOR2X1 U9116 ( .A(n7892), .B(ICACHE_addr[9]), .Y(n7914) );
  XOR2X1 U9117 ( .A(n7818), .B(ICACHE_addr[5]), .Y(n7848) );
  XOR2X1 U9118 ( .A(n7861), .B(ICACHE_addr[7]), .Y(n7880) );
  XOR2X1 U9119 ( .A(n7823), .B(ICACHE_addr[4]), .Y(n8358) );
  XOR2X1 U9120 ( .A(n7817), .B(ICACHE_addr[8]), .Y(n7895) );
  OAI221X1 U9121 ( .A0(\i_MIPS/ALUin1[12] ), .A1(n14), .B0(\i_MIPS/ALUin1[11] ), .B1(n3077), .C0(n4984), .Y(n5269) );
  OAI221XL U9122 ( .A0(\i_MIPS/ALUin1[20] ), .A1(n3082), .B0(
        \i_MIPS/ALUin1[21] ), .B1(n3077), .C0(n5466), .Y(n5823) );
  OAI221XL U9123 ( .A0(\i_MIPS/ALUin1[19] ), .A1(n3091), .B0(
        \i_MIPS/ALUin1[20] ), .B1(n3086), .C0(n6049), .Y(n6675) );
  OAI221XL U9124 ( .A0(\i_MIPS/ALUin1[19] ), .A1(n3082), .B0(
        \i_MIPS/ALUin1[20] ), .B1(n3077), .C0(n4814), .Y(n5963) );
  OAI221XL U9125 ( .A0(\i_MIPS/ALUin1[20] ), .A1(n3091), .B0(
        \i_MIPS/ALUin1[21] ), .B1(n3086), .C0(n4711), .Y(n6757) );
  OAI221XL U9126 ( .A0(\i_MIPS/ALUin1[18] ), .A1(n3082), .B0(
        \i_MIPS/ALUin1[19] ), .B1(n3077), .C0(n4712), .Y(n5620) );
  CLKMX2X2 U9127 ( .A(n2928), .B(n2929), .S0(n3067), .Y(\D_cache/N152 ) );
  OAI221XL U9128 ( .A0(\i_MIPS/ALUin1[9] ), .A1(n3091), .B0(\i_MIPS/ALUin1[8] ), .B1(n3086), .C0(n4910), .Y(n6613) );
  OAI211X1 U9129 ( .A0(\i_MIPS/ID_EX[80] ), .A1(n6528), .B0(n5463), .C0(n5118), 
        .Y(n5401) );
  OAI221XL U9130 ( .A0(\i_MIPS/ALUin1[7] ), .A1(n3091), .B0(\i_MIPS/ALUin1[6] ), .B1(n3086), .C0(n5038), .Y(n5330) );
  OAI222XL U9131 ( .A0(n8334), .A1(n66), .B0(n3638), .B1(n8333), .C0(n3688), 
        .C1(\i_MIPS/n211 ), .Y(n8773) );
  OAI222XL U9132 ( .A0(n3585), .A1(n67), .B0(n3643), .B1(n8333), .C0(n3688), 
        .C1(\i_MIPS/n208 ), .Y(n8776) );
  AO22X2 U9133 ( .A0(mem_rdata_I[31]), .A1(n3605), .B0(n3591), .B1(n8585), .Y(
        n8409) );
  AO22X2 U9134 ( .A0(mem_rdata_I[30]), .A1(n3605), .B0(n3589), .B1(n8584), .Y(
        n7275) );
  AO22X2 U9135 ( .A0(mem_rdata_I[29]), .A1(n3604), .B0(n3589), .B1(n8583), .Y(
        n7251) );
  AO22X2 U9136 ( .A0(mem_rdata_I[28]), .A1(n3604), .B0(n3588), .B1(n8582), .Y(
        n7227) );
  AO22X2 U9137 ( .A0(mem_rdata_I[27]), .A1(n3604), .B0(n3588), .B1(n8581), .Y(
        n7203) );
  AO22X2 U9138 ( .A0(mem_rdata_I[26]), .A1(n3604), .B0(n3588), .B1(n8580), .Y(
        n7179) );
  AO22X2 U9139 ( .A0(mem_rdata_I[25]), .A1(n3607), .B0(n3591), .B1(n8579), .Y(
        n7651) );
  AO22X2 U9140 ( .A0(mem_rdata_I[24]), .A1(n3605), .B0(n3590), .B1(n8578), .Y(
        n7429) );
  AO22X2 U9141 ( .A0(mem_rdata_I[23]), .A1(n3605), .B0(n3590), .B1(n8577), .Y(
        n7453) );
  AO22X2 U9142 ( .A0(mem_rdata_I[22]), .A1(n3606), .B0(n3592), .B1(n8576), .Y(
        n8113) );
  AO22X2 U9143 ( .A0(mem_rdata_I[21]), .A1(n3605), .B0(n3590), .B1(n8575), .Y(
        n7477) );
  AO22X2 U9144 ( .A0(mem_rdata_I[20]), .A1(n8453), .B0(n3588), .B1(n8574), .Y(
        n7501) );
  AO22X2 U9145 ( .A0(mem_rdata_I[19]), .A1(n3603), .B0(n3587), .B1(n8573), .Y(
        n7130) );
  AO22X2 U9146 ( .A0(mem_rdata_I[18]), .A1(n3603), .B0(n3587), .B1(n8572), .Y(
        n7154) );
  AO22X2 U9147 ( .A0(mem_rdata_I[17]), .A1(n3602), .B0(n3586), .B1(n8571), .Y(
        n4583) );
  AO22X2 U9148 ( .A0(mem_rdata_I[16]), .A1(n3603), .B0(n3587), .B1(n8570), .Y(
        n7106) );
  AO22X2 U9149 ( .A0(mem_rdata_I[14]), .A1(n3608), .B0(n3592), .B1(n8568), .Y(
        n7525) );
  AO22X2 U9150 ( .A0(mem_rdata_I[13]), .A1(n3606), .B0(n3591), .B1(n8567), .Y(
        n7574) );
  AO22X2 U9151 ( .A0(mem_rdata_I[12]), .A1(n3606), .B0(n3591), .B1(n8566), .Y(
        n7622) );
  AO22X2 U9152 ( .A0(mem_rdata_I[11]), .A1(n3606), .B0(n3591), .B1(n8565), .Y(
        n7598) );
  AO22X2 U9153 ( .A0(mem_rdata_I[10]), .A1(n3607), .B0(n3591), .B1(n8564), .Y(
        n7676) );
  AO22X2 U9154 ( .A0(mem_rdata_I[9]), .A1(n3607), .B0(n3591), .B1(n8563), .Y(
        n7699) );
  AO22X2 U9155 ( .A0(mem_rdata_I[8]), .A1(n3608), .B0(n3589), .B1(n8562), .Y(
        n7723) );
  AO22X2 U9156 ( .A0(mem_rdata_I[7]), .A1(n3608), .B0(n3589), .B1(n8561), .Y(
        n7749) );
  AO22X2 U9157 ( .A0(mem_rdata_I[6]), .A1(n3608), .B0(n3589), .B1(n8560), .Y(
        n7772) );
  AO22X2 U9158 ( .A0(mem_rdata_I[5]), .A1(n3604), .B0(n3589), .B1(n8559), .Y(
        n7401) );
  AO22X2 U9159 ( .A0(mem_rdata_I[4]), .A1(n3609), .B0(n3592), .B1(n8558), .Y(
        n8346) );
  AO22X2 U9160 ( .A0(mem_rdata_I[3]), .A1(n3605), .B0(n3592), .B1(n8557), .Y(
        n8365) );
  AO22X2 U9161 ( .A0(mem_rdata_I[2]), .A1(n3607), .B0(n3592), .B1(n8556), .Y(
        n8379) );
  AO22X2 U9162 ( .A0(mem_rdata_I[1]), .A1(n3602), .B0(n3590), .B1(n8555), .Y(
        n4563) );
  AO22X2 U9163 ( .A0(mem_rdata_I[0]), .A1(n8453), .B0(n3587), .B1(n8554), .Y(
        n8397) );
  AO22X2 U9164 ( .A0(mem_rdata_I[63]), .A1(n3604), .B0(n3591), .B1(n8617), .Y(
        n8411) );
  AO22X2 U9165 ( .A0(mem_rdata_I[62]), .A1(n3605), .B0(n3589), .B1(n8616), .Y(
        n7280) );
  AO22X2 U9166 ( .A0(mem_rdata_I[61]), .A1(n3604), .B0(n3589), .B1(n8615), .Y(
        n7256) );
  AO22X2 U9167 ( .A0(mem_rdata_I[60]), .A1(n3604), .B0(n3588), .B1(n8614), .Y(
        n7232) );
  AO22X2 U9168 ( .A0(mem_rdata_I[59]), .A1(n3604), .B0(n3588), .B1(n8613), .Y(
        n7208) );
  AO22X2 U9169 ( .A0(mem_rdata_I[58]), .A1(n3604), .B0(n3588), .B1(n8612), .Y(
        n7184) );
  AO22X2 U9170 ( .A0(mem_rdata_I[57]), .A1(n3607), .B0(n3587), .B1(n8611), .Y(
        n7656) );
  AO22X2 U9171 ( .A0(mem_rdata_I[56]), .A1(n3605), .B0(n3590), .B1(n8610), .Y(
        n7434) );
  AO22X2 U9172 ( .A0(mem_rdata_I[55]), .A1(n3605), .B0(n3590), .B1(n8609), .Y(
        n7458) );
  AO22X2 U9173 ( .A0(mem_rdata_I[54]), .A1(n3606), .B0(n3592), .B1(n8608), .Y(
        n8119) );
  AO22X2 U9174 ( .A0(mem_rdata_I[53]), .A1(n3605), .B0(n3590), .B1(n8607), .Y(
        n7482) );
  AO22X2 U9175 ( .A0(mem_rdata_I[52]), .A1(n3605), .B0(n3590), .B1(n8606), .Y(
        n7506) );
  AO22X2 U9176 ( .A0(mem_rdata_I[51]), .A1(n3603), .B0(n3587), .B1(n8605), .Y(
        n7135) );
  AO22X2 U9177 ( .A0(mem_rdata_I[50]), .A1(n3603), .B0(n3587), .B1(n8604), .Y(
        n7159) );
  AO22X2 U9178 ( .A0(mem_rdata_I[49]), .A1(n3602), .B0(n3590), .B1(n8603), .Y(
        n4588) );
  AO22X2 U9179 ( .A0(mem_rdata_I[48]), .A1(n3603), .B0(n3587), .B1(n8602), .Y(
        n7111) );
  AO22X2 U9180 ( .A0(mem_rdata_I[46]), .A1(n3606), .B0(n3592), .B1(n8600), .Y(
        n7530) );
  AO22X2 U9181 ( .A0(mem_rdata_I[45]), .A1(n3606), .B0(n3591), .B1(n8599), .Y(
        n7579) );
  AO22X2 U9182 ( .A0(mem_rdata_I[44]), .A1(n3606), .B0(n3591), .B1(n8598), .Y(
        n7627) );
  AO22X2 U9183 ( .A0(mem_rdata_I[43]), .A1(n3606), .B0(n3591), .B1(n8597), .Y(
        n7603) );
  AO22X2 U9184 ( .A0(mem_rdata_I[42]), .A1(n3607), .B0(n3591), .B1(n8596), .Y(
        n7681) );
  AO22X2 U9185 ( .A0(mem_rdata_I[41]), .A1(n3607), .B0(n3587), .B1(n8595), .Y(
        n7704) );
  AO22X2 U9186 ( .A0(mem_rdata_I[40]), .A1(n3608), .B0(n3589), .B1(n8594), .Y(
        n7727) );
  AO22X2 U9187 ( .A0(mem_rdata_I[39]), .A1(n3608), .B0(n3587), .B1(n8593), .Y(
        n7754) );
  AO22X2 U9188 ( .A0(mem_rdata_I[38]), .A1(n3608), .B0(n3589), .B1(n8592), .Y(
        n7777) );
  AO22X2 U9189 ( .A0(mem_rdata_I[37]), .A1(n3605), .B0(n3589), .B1(n8591), .Y(
        n7406) );
  AO22X2 U9190 ( .A0(mem_rdata_I[36]), .A1(n3607), .B0(n3592), .B1(n8590), .Y(
        n8347) );
  AO22X2 U9191 ( .A0(mem_rdata_I[35]), .A1(n3604), .B0(n3592), .B1(n8589), .Y(
        n8366) );
  AO22X2 U9192 ( .A0(mem_rdata_I[34]), .A1(n3609), .B0(n3592), .B1(n8588), .Y(
        n8380) );
  AO22X2 U9193 ( .A0(mem_rdata_I[33]), .A1(n3602), .B0(n3588), .B1(n8587), .Y(
        n4568) );
  AO22X2 U9194 ( .A0(mem_rdata_I[32]), .A1(n8453), .B0(n3589), .B1(n8586), .Y(
        n8398) );
  AO22X2 U9195 ( .A0(mem_rdata_I[95]), .A1(n3605), .B0(n3586), .B1(n8649), .Y(
        n8408) );
  AO22X2 U9196 ( .A0(mem_rdata_I[94]), .A1(n3605), .B0(n3589), .B1(n8648), .Y(
        n7270) );
  AO22X2 U9197 ( .A0(mem_rdata_I[93]), .A1(n3604), .B0(n3588), .B1(n8647), .Y(
        n7246) );
  AO22X2 U9198 ( .A0(mem_rdata_I[92]), .A1(n3604), .B0(n3588), .B1(n8646), .Y(
        n7222) );
  AO22X2 U9199 ( .A0(mem_rdata_I[91]), .A1(n3604), .B0(n3588), .B1(n8645), .Y(
        n7198) );
  AO22X2 U9200 ( .A0(mem_rdata_I[90]), .A1(n3603), .B0(n3587), .B1(n8644), .Y(
        n7174) );
  AO22X2 U9201 ( .A0(mem_rdata_I[89]), .A1(n3606), .B0(n3591), .B1(n8643), .Y(
        n7646) );
  AO22X2 U9202 ( .A0(mem_rdata_I[88]), .A1(n3604), .B0(n3589), .B1(n8642), .Y(
        n7424) );
  AO22X2 U9203 ( .A0(mem_rdata_I[87]), .A1(n3605), .B0(n3590), .B1(n8641), .Y(
        n7448) );
  AO22X2 U9204 ( .A0(mem_rdata_I[86]), .A1(n3608), .B0(n3592), .B1(n8640), .Y(
        n8108) );
  AO22X2 U9205 ( .A0(mem_rdata_I[85]), .A1(n3605), .B0(n3590), .B1(n8639), .Y(
        n7472) );
  AO22X2 U9206 ( .A0(mem_rdata_I[84]), .A1(n3605), .B0(n3590), .B1(n8638), .Y(
        n7496) );
  AO22X2 U9207 ( .A0(mem_rdata_I[83]), .A1(n3603), .B0(n3587), .B1(n8637), .Y(
        n7125) );
  AO22X2 U9208 ( .A0(mem_rdata_I[82]), .A1(n3603), .B0(n3587), .B1(n8636), .Y(
        n7149) );
  AO22X2 U9209 ( .A0(mem_rdata_I[81]), .A1(n3602), .B0(n3592), .B1(n8635), .Y(
        n4578) );
  AO22X2 U9210 ( .A0(mem_rdata_I[80]), .A1(n3602), .B0(n3586), .B1(n8634), .Y(
        n7101) );
  AO22X2 U9211 ( .A0(mem_rdata_I[78]), .A1(n3609), .B0(n3588), .B1(n8632), .Y(
        n7520) );
  AO22X2 U9212 ( .A0(mem_rdata_I[77]), .A1(n3604), .B0(n3590), .B1(n8631), .Y(
        n7569) );
  AO22X2 U9213 ( .A0(mem_rdata_I[76]), .A1(n3606), .B0(n3591), .B1(n8630), .Y(
        n7618) );
  AO22X2 U9214 ( .A0(mem_rdata_I[75]), .A1(n3606), .B0(n3591), .B1(n8629), .Y(
        n7593) );
  AO22X2 U9215 ( .A0(mem_rdata_I[74]), .A1(n3607), .B0(n3587), .B1(n8628), .Y(
        n7671) );
  AO22X2 U9216 ( .A0(mem_rdata_I[73]), .A1(n3607), .B0(n3591), .B1(n8627), .Y(
        n7695) );
  AO22X2 U9217 ( .A0(mem_rdata_I[72]), .A1(n3607), .B0(n3587), .B1(n8626), .Y(
        n7718) );
  AO22X2 U9218 ( .A0(mem_rdata_I[71]), .A1(n3608), .B0(n3586), .B1(n8625), .Y(
        n7744) );
  AO22X2 U9219 ( .A0(mem_rdata_I[70]), .A1(n3608), .B0(n3588), .B1(n8624), .Y(
        n7768) );
  AO22X2 U9220 ( .A0(mem_rdata_I[69]), .A1(n3602), .B0(n3589), .B1(n8623), .Y(
        n7396) );
  AO22X2 U9221 ( .A0(mem_rdata_I[68]), .A1(n3602), .B0(n3592), .B1(n8622), .Y(
        n8345) );
  AO22X2 U9222 ( .A0(mem_rdata_I[67]), .A1(n3603), .B0(n3592), .B1(n8621), .Y(
        n8364) );
  AO22X2 U9223 ( .A0(mem_rdata_I[66]), .A1(n3603), .B0(n3592), .B1(n8620), .Y(
        n8378) );
  AO22X2 U9224 ( .A0(mem_rdata_I[65]), .A1(n3602), .B0(n3590), .B1(n8619), .Y(
        n4558) );
  AO22X2 U9225 ( .A0(mem_rdata_I[64]), .A1(n8453), .B0(n3586), .B1(n8618), .Y(
        n8396) );
  AO22X2 U9226 ( .A0(mem_rdata_I[127]), .A1(n3609), .B0(n3586), .B1(n8681), 
        .Y(n8407) );
  AO22X2 U9227 ( .A0(mem_rdata_I[126]), .A1(n3603), .B0(n3589), .B1(n8680), 
        .Y(n7265) );
  AO22X2 U9228 ( .A0(mem_rdata_I[125]), .A1(n3604), .B0(n3588), .B1(n8679), 
        .Y(n7241) );
  AO22X2 U9229 ( .A0(mem_rdata_I[124]), .A1(n3604), .B0(n3588), .B1(n8678), 
        .Y(n7217) );
  AO22X2 U9230 ( .A0(mem_rdata_I[123]), .A1(n3604), .B0(n3588), .B1(n8677), 
        .Y(n7193) );
  AO22X2 U9231 ( .A0(mem_rdata_I[122]), .A1(n3603), .B0(n3587), .B1(n8676), 
        .Y(n7169) );
  AO22X2 U9232 ( .A0(mem_rdata_I[121]), .A1(n3606), .B0(n3591), .B1(n8675), 
        .Y(n7641) );
  AO22X2 U9233 ( .A0(mem_rdata_I[120]), .A1(n3604), .B0(n3589), .B1(n8674), 
        .Y(n7419) );
  AO22X2 U9234 ( .A0(mem_rdata_I[119]), .A1(n3605), .B0(n3590), .B1(n8673), 
        .Y(n7443) );
  AO22X2 U9235 ( .A0(mem_rdata_I[118]), .A1(n3608), .B0(n3590), .B1(n8672), 
        .Y(n8103) );
  AO22X2 U9236 ( .A0(mem_rdata_I[117]), .A1(n3605), .B0(n3590), .B1(n8671), 
        .Y(n7467) );
  AO22X2 U9237 ( .A0(mem_rdata_I[116]), .A1(n3605), .B0(n3590), .B1(n8670), 
        .Y(n7491) );
  AO22X2 U9238 ( .A0(mem_rdata_I[115]), .A1(n3603), .B0(n3587), .B1(n8669), 
        .Y(n7120) );
  AO22X2 U9239 ( .A0(mem_rdata_I[114]), .A1(n3603), .B0(n3587), .B1(n8668), 
        .Y(n7144) );
  AO22X2 U9240 ( .A0(mem_rdata_I[113]), .A1(n3602), .B0(n3588), .B1(n8667), 
        .Y(n4573) );
  AO22X2 U9241 ( .A0(mem_rdata_I[112]), .A1(n3602), .B0(n3592), .B1(n8666), 
        .Y(n7096) );
  AO22X2 U9242 ( .A0(mem_rdata_I[110]), .A1(n3609), .B0(n3590), .B1(n8664), 
        .Y(n7515) );
  AO22X2 U9243 ( .A0(mem_rdata_I[109]), .A1(n3607), .B0(n3592), .B1(n8663), 
        .Y(n7564) );
  AO22X2 U9244 ( .A0(mem_rdata_I[108]), .A1(n3606), .B0(n3591), .B1(n8662), 
        .Y(n7613) );
  AO22X2 U9245 ( .A0(mem_rdata_I[107]), .A1(n3606), .B0(n3591), .B1(n8661), 
        .Y(n7588) );
  AO22X2 U9246 ( .A0(mem_rdata_I[106]), .A1(n3607), .B0(n3591), .B1(n8660), 
        .Y(n7666) );
  AO22X2 U9247 ( .A0(mem_rdata_I[105]), .A1(n3607), .B0(n3587), .B1(n8659), 
        .Y(n7690) );
  AO22X2 U9248 ( .A0(mem_rdata_I[104]), .A1(n3607), .B0(n3586), .B1(n8658), 
        .Y(n7713) );
  AO22X2 U9249 ( .A0(mem_rdata_I[103]), .A1(n3608), .B0(n3586), .B1(n8657), 
        .Y(n7739) );
  AO22X2 U9250 ( .A0(mem_rdata_I[102]), .A1(n3608), .B0(n3589), .B1(n8656), 
        .Y(n7763) );
  AO22X2 U9251 ( .A0(mem_rdata_I[101]), .A1(n3608), .B0(n3589), .B1(n8655), 
        .Y(n7391) );
  AO22X2 U9252 ( .A0(mem_rdata_I[100]), .A1(n3602), .B0(n3588), .B1(n8654), 
        .Y(n4548) );
  AO22X2 U9253 ( .A0(mem_rdata_I[99]), .A1(n3602), .B0(n3592), .B1(n8653), .Y(
        n8363) );
  AO22X2 U9254 ( .A0(mem_rdata_I[98]), .A1(n3608), .B0(n3592), .B1(n8652), .Y(
        n8377) );
  AO22X2 U9255 ( .A0(mem_rdata_I[97]), .A1(n3602), .B0(n8410), .B1(n8651), .Y(
        n4553) );
  AO22X2 U9256 ( .A0(mem_rdata_I[96]), .A1(n8453), .B0(n3589), .B1(n8650), .Y(
        n8395) );
  AO22X2 U9257 ( .A0(mem_rdata_I[15]), .A1(n3603), .B0(n3588), .B1(n8569), .Y(
        n7549) );
  AO22X2 U9258 ( .A0(mem_rdata_I[47]), .A1(n3608), .B0(n3588), .B1(n8601), .Y(
        n7554) );
  AO22X2 U9259 ( .A0(mem_rdata_I[79]), .A1(n3606), .B0(n3590), .B1(n8633), .Y(
        n7544) );
  AO22X2 U9260 ( .A0(mem_rdata_I[111]), .A1(n3602), .B0(n3592), .B1(n8665), 
        .Y(n7539) );
  NAND2X1 U9261 ( .A(\i_MIPS/ALUin1[26] ), .B(n4630), .Y(n6064) );
  OAI221XL U9262 ( .A0(\i_MIPS/Register/register[2][12] ), .A1(n3175), .B0(
        \i_MIPS/Register/register[10][12] ), .B1(n16), .C0(n6298), .Y(n6306)
         );
  OAI221XL U9263 ( .A0(\i_MIPS/Register/register[2][13] ), .A1(n3175), .B0(
        \i_MIPS/Register/register[10][13] ), .B1(n16), .C0(n6433), .Y(n6441)
         );
  OAI221XL U9264 ( .A0(\i_MIPS/Register/register[2][4] ), .A1(n3123), .B0(
        \i_MIPS/Register/register[10][4] ), .B1(n2790), .C0(n5337), .Y(n5345)
         );
  OAI221XL U9265 ( .A0(\i_MIPS/Register/register[2][0] ), .A1(n3122), .B0(
        \i_MIPS/Register/register[10][0] ), .B1(n3119), .C0(n5063), .Y(n5071)
         );
  OAI221XL U9266 ( .A0(\i_MIPS/Register/register[18][8] ), .A1(n3124), .B0(
        \i_MIPS/Register/register[26][8] ), .B1(n3121), .C0(n6154), .Y(n6162)
         );
  OA22X1 U9267 ( .A0(\i_MIPS/Register/register[22][8] ), .A1(n3117), .B0(
        \i_MIPS/Register/register[30][8] ), .B1(n3115), .Y(n6154) );
  OAI221XL U9268 ( .A0(\i_MIPS/Register/register[2][8] ), .A1(n3124), .B0(
        \i_MIPS/Register/register[10][8] ), .B1(n3121), .C0(n6145), .Y(n6153)
         );
  OA22X1 U9269 ( .A0(\i_MIPS/Register/register[6][8] ), .A1(n3116), .B0(
        \i_MIPS/Register/register[14][8] ), .B1(n3115), .Y(n6145) );
  OAI221XL U9270 ( .A0(\i_MIPS/Register/register[18][9] ), .A1(n3124), .B0(
        \i_MIPS/Register/register[26][9] ), .B1(n3121), .C0(n6223), .Y(n6231)
         );
  OA22X1 U9271 ( .A0(\i_MIPS/Register/register[22][9] ), .A1(n3117), .B0(
        \i_MIPS/Register/register[30][9] ), .B1(n3113), .Y(n6223) );
  OAI221XL U9272 ( .A0(\i_MIPS/Register/register[2][9] ), .A1(n3123), .B0(
        \i_MIPS/Register/register[10][9] ), .B1(n3121), .C0(n6214), .Y(n6222)
         );
  OA22X1 U9273 ( .A0(\i_MIPS/Register/register[6][9] ), .A1(n3117), .B0(
        \i_MIPS/Register/register[14][9] ), .B1(n3114), .Y(n6214) );
  OAI221XL U9274 ( .A0(\i_MIPS/Register/register[2][9] ), .A1(n3175), .B0(
        \i_MIPS/Register/register[10][9] ), .B1(n16), .C0(n6235), .Y(n6243) );
  OA22X1 U9275 ( .A0(\i_MIPS/Register/register[6][9] ), .A1(n3172), .B0(
        \i_MIPS/Register/register[14][9] ), .B1(n3169), .Y(n6235) );
  OAI221XL U9276 ( .A0(\i_MIPS/Register/register[18][13] ), .A1(n3122), .B0(
        \i_MIPS/Register/register[26][13] ), .B1(n3121), .C0(n6421), .Y(n6429)
         );
  OA22X1 U9277 ( .A0(\i_MIPS/Register/register[22][13] ), .A1(n3117), .B0(
        \i_MIPS/Register/register[30][13] ), .B1(n3115), .Y(n6421) );
  OAI221XL U9278 ( .A0(\i_MIPS/Register/register[2][13] ), .A1(n2791), .B0(
        \i_MIPS/Register/register[10][13] ), .B1(n3121), .C0(n6412), .Y(n6420)
         );
  OA22X1 U9279 ( .A0(\i_MIPS/Register/register[6][13] ), .A1(n3117), .B0(
        \i_MIPS/Register/register[14][13] ), .B1(n3114), .Y(n6412) );
  OAI221XL U9280 ( .A0(\i_MIPS/Register/register[18][14] ), .A1(n3175), .B0(
        \i_MIPS/Register/register[26][14] ), .B1(n16), .C0(n6376), .Y(n6384)
         );
  OA22X1 U9281 ( .A0(\i_MIPS/Register/register[22][14] ), .A1(n3172), .B0(
        \i_MIPS/Register/register[30][14] ), .B1(n3169), .Y(n6376) );
  OAI221XL U9282 ( .A0(\i_MIPS/Register/register[2][14] ), .A1(n3175), .B0(
        \i_MIPS/Register/register[10][14] ), .B1(n16), .C0(n6367), .Y(n6375)
         );
  OA22X1 U9283 ( .A0(\i_MIPS/Register/register[6][14] ), .A1(n3172), .B0(
        \i_MIPS/Register/register[14][14] ), .B1(n3169), .Y(n6367) );
  OAI221XL U9284 ( .A0(\i_MIPS/Register/register[18][14] ), .A1(n3122), .B0(
        \i_MIPS/Register/register[26][14] ), .B1(n3121), .C0(n6355), .Y(n6363)
         );
  OA22X1 U9285 ( .A0(\i_MIPS/Register/register[22][14] ), .A1(n3117), .B0(
        \i_MIPS/Register/register[30][14] ), .B1(n2782), .Y(n6355) );
  OAI221XL U9286 ( .A0(\i_MIPS/Register/register[2][14] ), .A1(n3124), .B0(
        \i_MIPS/Register/register[10][14] ), .B1(n3121), .C0(n6346), .Y(n6354)
         );
  OA22X1 U9287 ( .A0(\i_MIPS/Register/register[6][14] ), .A1(n3117), .B0(
        \i_MIPS/Register/register[14][14] ), .B1(n3113), .Y(n6346) );
  OAI221XL U9288 ( .A0(\i_MIPS/Register/register[18][4] ), .A1(n3173), .B0(
        \i_MIPS/Register/register[26][4] ), .B1(n16), .C0(n5367), .Y(n5375) );
  OAI221XL U9289 ( .A0(\i_MIPS/Register/register[2][4] ), .A1(n3173), .B0(
        \i_MIPS/Register/register[10][4] ), .B1(n16), .C0(n5358), .Y(n5366) );
  OAI221XL U9290 ( .A0(\i_MIPS/Register/register[18][11] ), .A1(n3123), .B0(
        \i_MIPS/Register/register[26][11] ), .B1(n3119), .C0(n5285), .Y(n5293)
         );
  OA22X1 U9291 ( .A0(\i_MIPS/Register/register[22][11] ), .A1(n2776), .B0(
        \i_MIPS/Register/register[30][11] ), .B1(n3114), .Y(n5285) );
  OAI221XL U9292 ( .A0(\i_MIPS/Register/register[2][11] ), .A1(n3123), .B0(
        \i_MIPS/Register/register[10][11] ), .B1(n3121), .C0(n5276), .Y(n5284)
         );
  OA22X1 U9293 ( .A0(\i_MIPS/Register/register[6][11] ), .A1(n2776), .B0(
        \i_MIPS/Register/register[14][11] ), .B1(n3114), .Y(n5276) );
  OAI221XL U9294 ( .A0(\i_MIPS/Register/register[18][10] ), .A1(n3173), .B0(
        \i_MIPS/Register/register[26][10] ), .B1(n16), .C0(n5241), .Y(n5249)
         );
  OA22X1 U9295 ( .A0(\i_MIPS/Register/register[22][10] ), .A1(n3171), .B0(
        \i_MIPS/Register/register[30][10] ), .B1(n3167), .Y(n5241) );
  OAI221XL U9296 ( .A0(\i_MIPS/Register/register[2][10] ), .A1(n3173), .B0(
        \i_MIPS/Register/register[10][10] ), .B1(n16), .C0(n5232), .Y(n5240)
         );
  OA22X1 U9297 ( .A0(\i_MIPS/Register/register[6][10] ), .A1(n3170), .B0(
        \i_MIPS/Register/register[14][10] ), .B1(n3169), .Y(n5232) );
  OAI221XL U9298 ( .A0(\i_MIPS/Register/register[18][10] ), .A1(n3123), .B0(
        \i_MIPS/Register/register[26][10] ), .B1(n3119), .C0(n5220), .Y(n5228)
         );
  OA22X1 U9299 ( .A0(\i_MIPS/Register/register[22][10] ), .A1(n3116), .B0(
        \i_MIPS/Register/register[30][10] ), .B1(n3114), .Y(n5220) );
  OAI221XL U9300 ( .A0(\i_MIPS/Register/register[2][10] ), .A1(n3122), .B0(
        \i_MIPS/Register/register[10][10] ), .B1(n2790), .C0(n5211), .Y(n5219)
         );
  OA22X1 U9301 ( .A0(\i_MIPS/Register/register[6][10] ), .A1(n3116), .B0(
        \i_MIPS/Register/register[14][10] ), .B1(n3113), .Y(n5211) );
  OAI221XL U9302 ( .A0(\i_MIPS/Register/register[18][5] ), .A1(n3173), .B0(
        \i_MIPS/Register/register[26][5] ), .B1(n16), .C0(n5436), .Y(n5444) );
  OA22X1 U9303 ( .A0(\i_MIPS/Register/register[22][5] ), .A1(n3171), .B0(
        \i_MIPS/Register/register[30][5] ), .B1(n3167), .Y(n5436) );
  OAI221XL U9304 ( .A0(\i_MIPS/Register/register[2][5] ), .A1(n3173), .B0(
        \i_MIPS/Register/register[10][5] ), .B1(n16), .C0(n5427), .Y(n5435) );
  OA22X1 U9305 ( .A0(\i_MIPS/Register/register[6][5] ), .A1(n3171), .B0(
        \i_MIPS/Register/register[14][5] ), .B1(n3167), .Y(n5427) );
  OAI221XL U9306 ( .A0(\i_MIPS/Register/register[18][5] ), .A1(n3123), .B0(
        \i_MIPS/Register/register[26][5] ), .B1(n3120), .C0(n5415), .Y(n5423)
         );
  OA22X1 U9307 ( .A0(\i_MIPS/Register/register[22][5] ), .A1(n3117), .B0(
        \i_MIPS/Register/register[30][5] ), .B1(n3114), .Y(n5415) );
  OAI221XL U9308 ( .A0(\i_MIPS/Register/register[2][5] ), .A1(n3123), .B0(
        \i_MIPS/Register/register[10][5] ), .B1(n3120), .C0(n5406), .Y(n5414)
         );
  OA22X1 U9309 ( .A0(\i_MIPS/Register/register[6][5] ), .A1(n3118), .B0(
        \i_MIPS/Register/register[14][5] ), .B1(n3114), .Y(n5406) );
  OAI221XL U9310 ( .A0(\i_MIPS/Register/register[18][7] ), .A1(n2792), .B0(
        \i_MIPS/Register/register[26][7] ), .B1(n16), .C0(n5023), .Y(n5031) );
  OA22X1 U9311 ( .A0(\i_MIPS/Register/register[22][7] ), .A1(n3170), .B0(
        \i_MIPS/Register/register[30][7] ), .B1(n2773), .Y(n5023) );
  OAI221XL U9312 ( .A0(\i_MIPS/Register/register[2][7] ), .A1(n2792), .B0(
        \i_MIPS/Register/register[10][7] ), .B1(n16), .C0(n5014), .Y(n5022) );
  OA22X1 U9313 ( .A0(\i_MIPS/Register/register[6][7] ), .A1(n3170), .B0(
        \i_MIPS/Register/register[14][7] ), .B1(n2773), .Y(n5014) );
  OAI221XL U9314 ( .A0(\i_MIPS/Register/register[18][7] ), .A1(n3122), .B0(
        \i_MIPS/Register/register[26][7] ), .B1(n3119), .C0(n5002), .Y(n5010)
         );
  OA22X1 U9315 ( .A0(\i_MIPS/Register/register[22][7] ), .A1(n3116), .B0(
        \i_MIPS/Register/register[30][7] ), .B1(n3113), .Y(n5002) );
  OAI221XL U9316 ( .A0(\i_MIPS/Register/register[2][7] ), .A1(n3122), .B0(
        \i_MIPS/Register/register[10][7] ), .B1(n3119), .C0(n4993), .Y(n5001)
         );
  OA22X1 U9317 ( .A0(\i_MIPS/Register/register[6][7] ), .A1(n3116), .B0(
        \i_MIPS/Register/register[14][7] ), .B1(n3113), .Y(n4993) );
  OAI221XL U9318 ( .A0(\i_MIPS/Register/register[18][6] ), .A1(n3174), .B0(
        \i_MIPS/Register/register[26][6] ), .B1(n16), .C0(n4953), .Y(n4961) );
  OA22X1 U9319 ( .A0(\i_MIPS/Register/register[22][6] ), .A1(n3170), .B0(
        \i_MIPS/Register/register[30][6] ), .B1(n3168), .Y(n4953) );
  OAI221XL U9320 ( .A0(\i_MIPS/Register/register[2][6] ), .A1(n3173), .B0(
        \i_MIPS/Register/register[10][6] ), .B1(n16), .C0(n4944), .Y(n4952) );
  OA22X1 U9321 ( .A0(\i_MIPS/Register/register[6][6] ), .A1(n3170), .B0(
        \i_MIPS/Register/register[14][6] ), .B1(n3167), .Y(n4944) );
  OAI221XL U9322 ( .A0(\i_MIPS/Register/register[18][6] ), .A1(n3122), .B0(
        \i_MIPS/Register/register[26][6] ), .B1(n3119), .C0(n4932), .Y(n4940)
         );
  OA22X1 U9323 ( .A0(\i_MIPS/Register/register[22][6] ), .A1(n3116), .B0(
        \i_MIPS/Register/register[30][6] ), .B1(n3113), .Y(n4932) );
  OAI221XL U9324 ( .A0(\i_MIPS/Register/register[2][6] ), .A1(n3122), .B0(
        \i_MIPS/Register/register[10][6] ), .B1(n3119), .C0(n4923), .Y(n4931)
         );
  OA22X1 U9325 ( .A0(\i_MIPS/Register/register[6][6] ), .A1(n3116), .B0(
        \i_MIPS/Register/register[14][6] ), .B1(n3113), .Y(n4923) );
  OAI221XL U9326 ( .A0(\i_MIPS/Register/register[18][1] ), .A1(n3174), .B0(
        \i_MIPS/Register/register[26][1] ), .B1(n16), .C0(n5165), .Y(n5173) );
  OA22X1 U9327 ( .A0(\i_MIPS/Register/register[22][1] ), .A1(n3170), .B0(
        \i_MIPS/Register/register[30][1] ), .B1(n3169), .Y(n5165) );
  OAI221XL U9328 ( .A0(\i_MIPS/Register/register[2][1] ), .A1(n2792), .B0(
        \i_MIPS/Register/register[10][1] ), .B1(n16), .C0(n5156), .Y(n5164) );
  OA22X1 U9329 ( .A0(\i_MIPS/Register/register[6][1] ), .A1(n3170), .B0(
        \i_MIPS/Register/register[14][1] ), .B1(n2773), .Y(n5156) );
  OAI221XL U9330 ( .A0(\i_MIPS/Register/register[18][1] ), .A1(n3122), .B0(
        \i_MIPS/Register/register[26][1] ), .B1(n3119), .C0(n5144), .Y(n5152)
         );
  OA22X1 U9331 ( .A0(\i_MIPS/Register/register[22][1] ), .A1(n3116), .B0(
        \i_MIPS/Register/register[30][1] ), .B1(n3113), .Y(n5144) );
  OAI221XL U9332 ( .A0(\i_MIPS/Register/register[2][1] ), .A1(n3122), .B0(
        \i_MIPS/Register/register[10][1] ), .B1(n3119), .C0(n5135), .Y(n5143)
         );
  OA22X1 U9333 ( .A0(\i_MIPS/Register/register[6][1] ), .A1(n3116), .B0(
        \i_MIPS/Register/register[14][1] ), .B1(n3113), .Y(n5135) );
  OAI221XL U9334 ( .A0(\i_MIPS/Register/register[18][0] ), .A1(n3175), .B0(
        \i_MIPS/Register/register[26][0] ), .B1(n16), .C0(n5093), .Y(n5101) );
  OAI221XL U9335 ( .A0(\i_MIPS/Register/register[2][0] ), .A1(n3174), .B0(
        \i_MIPS/Register/register[10][0] ), .B1(n16), .C0(n5084), .Y(n5092) );
  OAI221XL U9336 ( .A0(\i_MIPS/Register/register[18][2] ), .A1(n3173), .B0(
        \i_MIPS/Register/register[26][2] ), .B1(n16), .C0(n6657), .Y(n6665) );
  OA22X1 U9337 ( .A0(\i_MIPS/Register/register[22][2] ), .A1(n3172), .B0(
        \i_MIPS/Register/register[30][2] ), .B1(n3169), .Y(n6657) );
  OAI221XL U9338 ( .A0(\i_MIPS/Register/register[2][2] ), .A1(n3175), .B0(
        \i_MIPS/Register/register[10][2] ), .B1(n16), .C0(n6648), .Y(n6656) );
  OA22X1 U9339 ( .A0(\i_MIPS/Register/register[6][2] ), .A1(n3172), .B0(
        \i_MIPS/Register/register[14][2] ), .B1(n3167), .Y(n6648) );
  OAI221XL U9340 ( .A0(\i_MIPS/Register/register[18][2] ), .A1(n3122), .B0(
        \i_MIPS/Register/register[26][2] ), .B1(n3120), .C0(n6636), .Y(n6644)
         );
  OAI221XL U9341 ( .A0(\i_MIPS/Register/register[2][2] ), .A1(n3124), .B0(
        \i_MIPS/Register/register[10][2] ), .B1(n3121), .C0(n6627), .Y(n6635)
         );
  OAI221XL U9342 ( .A0(\i_MIPS/Register/register[18][3] ), .A1(n3175), .B0(
        \i_MIPS/Register/register[26][3] ), .B1(n16), .C0(n6585), .Y(n6593) );
  OAI221XL U9343 ( .A0(\i_MIPS/Register/register[2][3] ), .A1(n3175), .B0(
        \i_MIPS/Register/register[10][3] ), .B1(n16), .C0(n6576), .Y(n6584) );
  OAI221XL U9344 ( .A0(\i_MIPS/Register/register[18][3] ), .A1(n3122), .B0(
        \i_MIPS/Register/register[26][3] ), .B1(n3120), .C0(n6564), .Y(n6572)
         );
  OAI221XL U9345 ( .A0(\i_MIPS/Register/register[2][3] ), .A1(n3124), .B0(
        \i_MIPS/Register/register[10][3] ), .B1(n3121), .C0(n6555), .Y(n6563)
         );
  OAI221XL U9346 ( .A0(\i_MIPS/Register/register[2][16] ), .A1(n2791), .B0(
        \i_MIPS/Register/register[10][16] ), .B1(n3119), .C0(n6950), .Y(n6958)
         );
  OA22X1 U9347 ( .A0(\i_MIPS/Register/register[6][16] ), .A1(n3118), .B0(
        \i_MIPS/Register/register[14][16] ), .B1(n2782), .Y(n6950) );
  OAI221XL U9348 ( .A0(\i_MIPS/Register/register[18][18] ), .A1(n3174), .B0(
        \i_MIPS/Register/register[26][18] ), .B1(n16), .C0(n5791), .Y(n5799)
         );
  OAI221XL U9349 ( .A0(\i_MIPS/Register/register[2][18] ), .A1(n3174), .B0(
        \i_MIPS/Register/register[10][18] ), .B1(n16), .C0(n5782), .Y(n5790)
         );
  OAI221XL U9350 ( .A0(\i_MIPS/Register/register[18][17] ), .A1(n3174), .B0(
        \i_MIPS/Register/register[26][17] ), .B1(n16), .C0(n5719), .Y(n5727)
         );
  OAI221XL U9351 ( .A0(\i_MIPS/Register/register[2][17] ), .A1(n3174), .B0(
        \i_MIPS/Register/register[10][17] ), .B1(n16), .C0(n5710), .Y(n5718)
         );
  OAI221XL U9352 ( .A0(\i_MIPS/Register/register[18][25] ), .A1(n3173), .B0(
        \i_MIPS/Register/register[26][25] ), .B1(n16), .C0(n5521), .Y(n5529)
         );
  OAI221XL U9353 ( .A0(\i_MIPS/Register/register[2][25] ), .A1(n3173), .B0(
        \i_MIPS/Register/register[10][25] ), .B1(n16), .C0(n5512), .Y(n5520)
         );
  OAI221XL U9354 ( .A0(\i_MIPS/Register/register[18][25] ), .A1(n3123), .B0(
        \i_MIPS/Register/register[26][25] ), .B1(n3119), .C0(n5498), .Y(n5506)
         );
  OAI221XL U9355 ( .A0(\i_MIPS/Register/register[2][25] ), .A1(n3123), .B0(
        \i_MIPS/Register/register[10][25] ), .B1(n3121), .C0(n5489), .Y(n5497)
         );
  OAI221XL U9356 ( .A0(\i_MIPS/Register/register[18][15] ), .A1(n3173), .B0(
        \i_MIPS/Register/register[26][15] ), .B1(n16), .C0(n5586), .Y(n5594)
         );
  OA22X1 U9357 ( .A0(\i_MIPS/Register/register[22][15] ), .A1(n3171), .B0(
        \i_MIPS/Register/register[30][15] ), .B1(n3167), .Y(n5586) );
  OAI221XL U9358 ( .A0(\i_MIPS/Register/register[2][15] ), .A1(n3173), .B0(
        \i_MIPS/Register/register[10][15] ), .B1(n16), .C0(n5577), .Y(n5585)
         );
  OA22X1 U9359 ( .A0(\i_MIPS/Register/register[6][15] ), .A1(n3171), .B0(
        \i_MIPS/Register/register[14][15] ), .B1(n3167), .Y(n5577) );
  OAI221XL U9360 ( .A0(\i_MIPS/Register/register[18][15] ), .A1(n3123), .B0(
        \i_MIPS/Register/register[26][15] ), .B1(n3121), .C0(n5565), .Y(n5573)
         );
  OA22X1 U9361 ( .A0(\i_MIPS/Register/register[22][15] ), .A1(n2776), .B0(
        \i_MIPS/Register/register[30][15] ), .B1(n3114), .Y(n5565) );
  OAI221XL U9362 ( .A0(\i_MIPS/Register/register[2][15] ), .A1(n3123), .B0(
        \i_MIPS/Register/register[10][15] ), .B1(n3120), .C0(n5556), .Y(n5564)
         );
  OA22X1 U9363 ( .A0(\i_MIPS/Register/register[6][15] ), .A1(n2776), .B0(
        \i_MIPS/Register/register[14][15] ), .B1(n3114), .Y(n5556) );
  OAI221XL U9364 ( .A0(\i_MIPS/Register/register[18][21] ), .A1(n3122), .B0(
        \i_MIPS/Register/register[26][21] ), .B1(n3121), .C0(n6491), .Y(n6499)
         );
  OAI221XL U9365 ( .A0(\i_MIPS/Register/register[2][21] ), .A1(n3123), .B0(
        \i_MIPS/Register/register[10][21] ), .B1(n3120), .C0(n6482), .Y(n6490)
         );
  OAI221XL U9366 ( .A0(\i_MIPS/Register/register[18][22] ), .A1(n3173), .B0(
        \i_MIPS/Register/register[26][22] ), .B1(n16), .C0(n6714), .Y(n6722)
         );
  OAI221XL U9367 ( .A0(\i_MIPS/Register/register[2][22] ), .A1(n3174), .B0(
        \i_MIPS/Register/register[10][22] ), .B1(n16), .C0(n6705), .Y(n6713)
         );
  OAI221XL U9368 ( .A0(\i_MIPS/Register/register[18][24] ), .A1(n3174), .B0(
        \i_MIPS/Register/register[26][24] ), .B1(n16), .C0(n6033), .Y(n6041)
         );
  OAI221XL U9369 ( .A0(\i_MIPS/Register/register[2][24] ), .A1(n3174), .B0(
        \i_MIPS/Register/register[10][24] ), .B1(n16), .C0(n6024), .Y(n6032)
         );
  OAI221XL U9370 ( .A0(\i_MIPS/Register/register[18][24] ), .A1(n3124), .B0(
        \i_MIPS/Register/register[26][24] ), .B1(n3120), .C0(n6010), .Y(n6018)
         );
  OAI221XL U9371 ( .A0(\i_MIPS/Register/register[2][24] ), .A1(n3124), .B0(
        \i_MIPS/Register/register[10][24] ), .B1(n3120), .C0(n6001), .Y(n6009)
         );
  OAI221XL U9372 ( .A0(\i_MIPS/Register/register[18][26] ), .A1(n3174), .B0(
        \i_MIPS/Register/register[26][26] ), .B1(n16), .C0(n6108), .Y(n6116)
         );
  OAI221XL U9373 ( .A0(\i_MIPS/Register/register[2][26] ), .A1(n3174), .B0(
        \i_MIPS/Register/register[10][26] ), .B1(n16), .C0(n6099), .Y(n6107)
         );
  OAI221XL U9374 ( .A0(\i_MIPS/Register/register[18][26] ), .A1(n3124), .B0(
        \i_MIPS/Register/register[26][26] ), .B1(n3121), .C0(n6085), .Y(n6093)
         );
  OAI221XL U9375 ( .A0(\i_MIPS/Register/register[2][26] ), .A1(n3124), .B0(
        \i_MIPS/Register/register[10][26] ), .B1(n3121), .C0(n6076), .Y(n6084)
         );
  OAI221XL U9376 ( .A0(\i_MIPS/Register/register[18][23] ), .A1(n3175), .B0(
        \i_MIPS/Register/register[26][23] ), .B1(n16), .C0(n6867), .Y(n6875)
         );
  OAI221XL U9377 ( .A0(\i_MIPS/Register/register[2][23] ), .A1(n3173), .B0(
        \i_MIPS/Register/register[10][23] ), .B1(n16), .C0(n6858), .Y(n6866)
         );
  OAI221XL U9378 ( .A0(\i_MIPS/Register/register[18][16] ), .A1(n3173), .B0(
        \i_MIPS/Register/register[26][16] ), .B1(n16), .C0(n6938), .Y(n6946)
         );
  OA22X1 U9379 ( .A0(\i_MIPS/Register/register[22][16] ), .A1(n2777), .B0(
        \i_MIPS/Register/register[30][16] ), .B1(n3167), .Y(n6938) );
  OAI221XL U9380 ( .A0(\i_MIPS/Register/register[2][16] ), .A1(n3175), .B0(
        \i_MIPS/Register/register[10][16] ), .B1(n16), .C0(n6929), .Y(n6937)
         );
  OA22X1 U9381 ( .A0(\i_MIPS/Register/register[6][16] ), .A1(n2777), .B0(
        \i_MIPS/Register/register[14][16] ), .B1(n3169), .Y(n6929) );
  OAI221XL U9382 ( .A0(\i_MIPS/Register/register[18][19] ), .A1(n3173), .B0(
        \i_MIPS/Register/register[26][19] ), .B1(n16), .C0(n5659), .Y(n5667)
         );
  OAI221XL U9383 ( .A0(\i_MIPS/Register/register[2][19] ), .A1(n3173), .B0(
        \i_MIPS/Register/register[10][19] ), .B1(n16), .C0(n5650), .Y(n5658)
         );
  OAI221XL U9384 ( .A0(\i_MIPS/Register/register[18][19] ), .A1(n3123), .B0(
        \i_MIPS/Register/register[26][19] ), .B1(n3120), .C0(n5636), .Y(n5644)
         );
  OAI221XL U9385 ( .A0(\i_MIPS/Register/register[2][19] ), .A1(n3123), .B0(
        \i_MIPS/Register/register[10][19] ), .B1(n3120), .C0(n5627), .Y(n5635)
         );
  OAI221XL U9386 ( .A0(\i_MIPS/Register/register[18][27] ), .A1(n3175), .B0(
        \i_MIPS/Register/register[26][27] ), .B1(n16), .C0(n6811), .Y(n6819)
         );
  OAI221XL U9387 ( .A0(\i_MIPS/Register/register[2][27] ), .A1(n3173), .B0(
        \i_MIPS/Register/register[10][27] ), .B1(n16), .C0(n6802), .Y(n6810)
         );
  OAI221XL U9388 ( .A0(\i_MIPS/Register/register[18][27] ), .A1(n3123), .B0(
        \i_MIPS/Register/register[26][27] ), .B1(n3121), .C0(n6788), .Y(n6796)
         );
  OAI221XL U9389 ( .A0(\i_MIPS/Register/register[2][27] ), .A1(n3124), .B0(
        \i_MIPS/Register/register[10][27] ), .B1(n3121), .C0(n6779), .Y(n6787)
         );
  OAI221XL U9390 ( .A0(\i_MIPS/Register/register[18][29] ), .A1(n3174), .B0(
        \i_MIPS/Register/register[26][29] ), .B1(n16), .C0(n5871), .Y(n5879)
         );
  OAI221XL U9391 ( .A0(\i_MIPS/Register/register[2][29] ), .A1(n3174), .B0(
        \i_MIPS/Register/register[10][29] ), .B1(n16), .C0(n5862), .Y(n5870)
         );
  OAI221XL U9392 ( .A0(\i_MIPS/Register/register[18][29] ), .A1(n3124), .B0(
        \i_MIPS/Register/register[26][29] ), .B1(n3120), .C0(n5848), .Y(n5856)
         );
  OAI221XL U9393 ( .A0(\i_MIPS/Register/register[2][29] ), .A1(n3124), .B0(
        \i_MIPS/Register/register[10][29] ), .B1(n3120), .C0(n5839), .Y(n5847)
         );
  OAI221XL U9394 ( .A0(\i_MIPS/Register/register[18][20] ), .A1(n3175), .B0(
        \i_MIPS/Register/register[26][20] ), .B1(n16), .C0(n4855), .Y(n4863)
         );
  OAI221XL U9395 ( .A0(\i_MIPS/Register/register[2][20] ), .A1(n3174), .B0(
        \i_MIPS/Register/register[10][20] ), .B1(n16), .C0(n4846), .Y(n4854)
         );
  OAI221XL U9396 ( .A0(\i_MIPS/Register/register[18][28] ), .A1(n3174), .B0(
        \i_MIPS/Register/register[26][28] ), .B1(n16), .C0(n5944), .Y(n5952)
         );
  OAI221XL U9397 ( .A0(\i_MIPS/Register/register[2][28] ), .A1(n3174), .B0(
        \i_MIPS/Register/register[10][28] ), .B1(n16), .C0(n5935), .Y(n5943)
         );
  OAI221XL U9398 ( .A0(\i_MIPS/Register/register[18][28] ), .A1(n3124), .B0(
        \i_MIPS/Register/register[26][28] ), .B1(n3120), .C0(n5921), .Y(n5929)
         );
  OAI221XL U9399 ( .A0(\i_MIPS/Register/register[2][28] ), .A1(n3124), .B0(
        \i_MIPS/Register/register[10][28] ), .B1(n3120), .C0(n5912), .Y(n5920)
         );
  OAI221XL U9400 ( .A0(\i_MIPS/Register/register[18][31] ), .A1(n3173), .B0(
        \i_MIPS/Register/register[26][31] ), .B1(n16), .C0(n4791), .Y(n4799)
         );
  OAI221XL U9401 ( .A0(\i_MIPS/Register/register[2][31] ), .A1(n3175), .B0(
        \i_MIPS/Register/register[10][31] ), .B1(n16), .C0(n4782), .Y(n4790)
         );
  OAI221XL U9402 ( .A0(\i_MIPS/Register/register[18][30] ), .A1(n3175), .B0(
        \i_MIPS/Register/register[26][30] ), .B1(n16), .C0(n7058), .Y(n7066)
         );
  OAI221XL U9403 ( .A0(\i_MIPS/Register/register[2][30] ), .A1(n3174), .B0(
        \i_MIPS/Register/register[10][30] ), .B1(n16), .C0(n7049), .Y(n7057)
         );
  OAI221XL U9404 ( .A0(\i_MIPS/Register/register[18][31] ), .A1(n3122), .B0(
        \i_MIPS/Register/register[26][31] ), .B1(n3119), .C0(n4753), .Y(n4761)
         );
  OAI221XL U9405 ( .A0(\i_MIPS/Register/register[2][31] ), .A1(n3122), .B0(
        \i_MIPS/Register/register[10][31] ), .B1(n3119), .C0(n4744), .Y(n4752)
         );
  OAI221XL U9406 ( .A0(\i_MIPS/Register/register[18][30] ), .A1(n3122), .B0(
        \i_MIPS/Register/register[26][30] ), .B1(n3120), .C0(n7031), .Y(n7039)
         );
  OAI221XL U9407 ( .A0(\i_MIPS/Register/register[2][30] ), .A1(n3123), .B0(
        \i_MIPS/Register/register[10][30] ), .B1(n3119), .C0(n7022), .Y(n7030)
         );
  OAI221XL U9408 ( .A0(\i_MIPS/Register/register[2][22] ), .A1(n3122), .B0(
        \i_MIPS/Register/register[10][22] ), .B1(n3120), .C0(n6726), .Y(n6734)
         );
  OAI221XL U9409 ( .A0(\i_MIPS/Register/register[2][23] ), .A1(n3123), .B0(
        \i_MIPS/Register/register[10][23] ), .B1(n3120), .C0(n6881), .Y(n6889)
         );
  OA22X1 U9410 ( .A0(\i_MIPS/Register/register[6][23] ), .A1(n3118), .B0(
        \i_MIPS/Register/register[14][23] ), .B1(n3113), .Y(n6881) );
  OAI221XL U9411 ( .A0(\i_MIPS/Register/register[2][20] ), .A1(n3122), .B0(
        \i_MIPS/Register/register[10][20] ), .B1(n3119), .C0(n4869), .Y(n4877)
         );
  OAI221XL U9412 ( .A0(\i_MIPS/Register/register[2][18] ), .A1(n3124), .B0(
        \i_MIPS/Register/register[10][18] ), .B1(n3120), .C0(n5761), .Y(n5769)
         );
  OAI221XL U9413 ( .A0(\i_MIPS/Register/register[2][17] ), .A1(n3124), .B0(
        \i_MIPS/Register/register[10][17] ), .B1(n3120), .C0(n5689), .Y(n5697)
         );
  OA22X1 U9414 ( .A0(\i_MIPS/Register/register[6][17] ), .A1(n3117), .B0(
        \i_MIPS/Register/register[14][17] ), .B1(n3115), .Y(n5689) );
  OAI2BB1X1 U9415 ( .A0N(n3084), .A1N(\i_MIPS/ALU/N303 ), .B0(n6995), .Y(n6686) );
  NAND3BX1 U9416 ( .AN(n2880), .B(n5465), .C(n4985), .Y(n5268) );
  NAND3BX1 U9417 ( .AN(n2879), .B(n5040), .C(n4815), .Y(n5962) );
  OAI2BB2XL U9418 ( .B0(n3677), .B1(n3780), .A0N(
        \i_MIPS/Register/register[0][7] ), .A1N(n3782), .Y(
        \i_MIPS/Register/n1115 ) );
  OAI2BB2XL U9419 ( .B0(n3677), .B1(n3777), .A0N(
        \i_MIPS/Register/register[1][7] ), .A1N(n3779), .Y(
        \i_MIPS/Register/n1083 ) );
  OAI2BB2XL U9420 ( .B0(n3677), .B1(n3774), .A0N(
        \i_MIPS/Register/register[2][7] ), .A1N(n3776), .Y(
        \i_MIPS/Register/n1051 ) );
  OAI2BB2XL U9421 ( .B0(n3677), .B1(n3771), .A0N(
        \i_MIPS/Register/register[3][7] ), .A1N(n3773), .Y(
        \i_MIPS/Register/n1019 ) );
  OAI2BB2XL U9422 ( .B0(n3677), .B1(n3768), .A0N(
        \i_MIPS/Register/register[4][7] ), .A1N(n3770), .Y(
        \i_MIPS/Register/n987 ) );
  OAI2BB2XL U9423 ( .B0(n3677), .B1(n3765), .A0N(
        \i_MIPS/Register/register[5][7] ), .A1N(n3767), .Y(
        \i_MIPS/Register/n955 ) );
  OAI2BB2XL U9424 ( .B0(n3677), .B1(n3762), .A0N(
        \i_MIPS/Register/register[6][7] ), .A1N(n3764), .Y(
        \i_MIPS/Register/n923 ) );
  OAI2BB2XL U9425 ( .B0(n3680), .B1(n3780), .A0N(
        \i_MIPS/Register/register[0][11] ), .A1N(n3782), .Y(
        \i_MIPS/Register/n1119 ) );
  OAI2BB2XL U9426 ( .B0(n3680), .B1(n3777), .A0N(
        \i_MIPS/Register/register[1][11] ), .A1N(n3779), .Y(
        \i_MIPS/Register/n1087 ) );
  OAI2BB2XL U9427 ( .B0(n3680), .B1(n3774), .A0N(
        \i_MIPS/Register/register[2][11] ), .A1N(n3776), .Y(
        \i_MIPS/Register/n1055 ) );
  OAI2BB2XL U9428 ( .B0(n3680), .B1(n3768), .A0N(
        \i_MIPS/Register/register[4][11] ), .A1N(n3770), .Y(
        \i_MIPS/Register/n991 ) );
  OAI2BB2XL U9429 ( .B0(n3680), .B1(n3762), .A0N(
        \i_MIPS/Register/register[6][11] ), .A1N(n3764), .Y(
        \i_MIPS/Register/n927 ) );
  OAI2BB2XL U9430 ( .B0(n3658), .B1(n3781), .A0N(
        \i_MIPS/Register/register[0][16] ), .A1N(n3782), .Y(
        \i_MIPS/Register/n1124 ) );
  OAI2BB2XL U9431 ( .B0(n3657), .B1(n3778), .A0N(
        \i_MIPS/Register/register[1][16] ), .A1N(n3779), .Y(
        \i_MIPS/Register/n1092 ) );
  OAI2BB2XL U9432 ( .B0(n3657), .B1(n3775), .A0N(
        \i_MIPS/Register/register[2][16] ), .A1N(n3776), .Y(
        \i_MIPS/Register/n1060 ) );
  OAI2BB2XL U9433 ( .B0(n3657), .B1(n3772), .A0N(
        \i_MIPS/Register/register[3][16] ), .A1N(n3773), .Y(
        \i_MIPS/Register/n1028 ) );
  OAI2BB2XL U9434 ( .B0(n3657), .B1(n3769), .A0N(
        \i_MIPS/Register/register[4][16] ), .A1N(n3770), .Y(
        \i_MIPS/Register/n996 ) );
  OAI2BB2XL U9435 ( .B0(n3657), .B1(n3766), .A0N(
        \i_MIPS/Register/register[5][16] ), .A1N(n3767), .Y(
        \i_MIPS/Register/n964 ) );
  OAI2BB2XL U9436 ( .B0(n3657), .B1(n3763), .A0N(
        \i_MIPS/Register/register[6][16] ), .A1N(n3764), .Y(
        \i_MIPS/Register/n932 ) );
  OAI2BB2XL U9437 ( .B0(n3657), .B1(n3727), .A0N(
        \i_MIPS/Register/register[18][16] ), .A1N(n3728), .Y(
        \i_MIPS/Register/n548 ) );
  OAI2BB2XL U9438 ( .B0(n3657), .B1(n3724), .A0N(
        \i_MIPS/Register/register[19][16] ), .A1N(n3725), .Y(
        \i_MIPS/Register/n516 ) );
  OAI2BB2XL U9439 ( .B0(n3657), .B1(n3721), .A0N(
        \i_MIPS/Register/register[20][16] ), .A1N(n3722), .Y(
        \i_MIPS/Register/n484 ) );
  OAI2BB2XL U9440 ( .B0(n3657), .B1(n3718), .A0N(
        \i_MIPS/Register/register[21][16] ), .A1N(n3719), .Y(
        \i_MIPS/Register/n452 ) );
  OAI2BB2XL U9441 ( .B0(n3657), .B1(n3715), .A0N(
        \i_MIPS/Register/register[22][16] ), .A1N(n3716), .Y(
        \i_MIPS/Register/n420 ) );
  OAI2BB2XL U9442 ( .B0(n3657), .B1(n3712), .A0N(
        \i_MIPS/Register/register[23][16] ), .A1N(n3713), .Y(
        \i_MIPS/Register/n388 ) );
  OAI2BB2XL U9443 ( .B0(n3658), .B1(n3709), .A0N(
        \i_MIPS/Register/register[24][16] ), .A1N(n3710), .Y(
        \i_MIPS/Register/n356 ) );
  OAI2BB2XL U9444 ( .B0(n3658), .B1(n3706), .A0N(
        \i_MIPS/Register/register[25][16] ), .A1N(n3707), .Y(
        \i_MIPS/Register/n324 ) );
  OAI2BB2XL U9445 ( .B0(n3658), .B1(n3703), .A0N(
        \i_MIPS/Register/register[26][16] ), .A1N(n3704), .Y(
        \i_MIPS/Register/n292 ) );
  OAI2BB2XL U9446 ( .B0(n3658), .B1(n3700), .A0N(
        \i_MIPS/Register/register[27][16] ), .A1N(n3701), .Y(
        \i_MIPS/Register/n260 ) );
  OAI2BB2XL U9447 ( .B0(n3658), .B1(n3697), .A0N(
        \i_MIPS/Register/register[28][16] ), .A1N(n3698), .Y(
        \i_MIPS/Register/n228 ) );
  OAI2BB2XL U9448 ( .B0(n3658), .B1(n3694), .A0N(
        \i_MIPS/Register/register[29][16] ), .A1N(n3695), .Y(
        \i_MIPS/Register/n196 ) );
  OAI2BB2XL U9449 ( .B0(n965), .B1(n3791), .A0N(\D_cache/cache[7][152] ), 
        .A1N(n3796), .Y(\D_cache/n573 ) );
  OAI2BB2XL U9450 ( .B0(n965), .B1(n3811), .A0N(\D_cache/cache[6][152] ), 
        .A1N(n3816), .Y(\D_cache/n574 ) );
  OAI2BB2XL U9451 ( .B0(n965), .B1(n3829), .A0N(\D_cache/cache[5][152] ), 
        .A1N(n3834), .Y(\D_cache/n575 ) );
  OAI2BB2XL U9452 ( .B0(n965), .B1(n3849), .A0N(\D_cache/cache[4][152] ), 
        .A1N(n3856), .Y(\D_cache/n576 ) );
  OAI2BB2XL U9453 ( .B0(n965), .B1(n3868), .A0N(\D_cache/cache[3][152] ), 
        .A1N(n3875), .Y(\D_cache/n577 ) );
  OAI2BB2XL U9454 ( .B0(n965), .B1(n3891), .A0N(\D_cache/cache[2][152] ), 
        .A1N(n3896), .Y(\D_cache/n578 ) );
  OAI2BB2XL U9455 ( .B0(n965), .B1(n3911), .A0N(\D_cache/cache[1][152] ), 
        .A1N(n3917), .Y(\D_cache/n579 ) );
  OAI2BB2XL U9456 ( .B0(n965), .B1(n3931), .A0N(\D_cache/cache[0][152] ), 
        .A1N(n3938), .Y(\D_cache/n580 ) );
  AO22X1 U9457 ( .A0(n3080), .A1(\i_MIPS/ALUin1[1] ), .B0(n3084), .B1(
        \i_MIPS/ALUin1[0] ), .Y(n5815) );
  OAI2BB2XL U9458 ( .B0(n3656), .B1(n3781), .A0N(
        \i_MIPS/Register/register[0][17] ), .A1N(n3780), .Y(
        \i_MIPS/Register/n1125 ) );
  OAI2BB2XL U9459 ( .B0(n3649), .B1(n3781), .A0N(
        \i_MIPS/Register/register[0][14] ), .A1N(n3782), .Y(
        \i_MIPS/Register/n1122 ) );
  OAI2BB2XL U9460 ( .B0(n3670), .B1(n3780), .A0N(
        \i_MIPS/Register/register[0][3] ), .A1N(n3782), .Y(
        \i_MIPS/Register/n1111 ) );
  OAI2BB2XL U9461 ( .B0(n3656), .B1(n3775), .A0N(
        \i_MIPS/Register/register[2][17] ), .A1N(n3774), .Y(
        \i_MIPS/Register/n1061 ) );
  OAI2BB2XL U9462 ( .B0(n3648), .B1(n3775), .A0N(
        \i_MIPS/Register/register[2][14] ), .A1N(n3776), .Y(
        \i_MIPS/Register/n1058 ) );
  OAI2BB2XL U9463 ( .B0(n3669), .B1(n3774), .A0N(
        \i_MIPS/Register/register[2][3] ), .A1N(n3776), .Y(
        \i_MIPS/Register/n1047 ) );
  OAI2BB2XL U9464 ( .B0(n3656), .B1(n3769), .A0N(
        \i_MIPS/Register/register[4][17] ), .A1N(n3768), .Y(
        \i_MIPS/Register/n997 ) );
  OAI2BB2XL U9465 ( .B0(n3648), .B1(n3769), .A0N(
        \i_MIPS/Register/register[4][14] ), .A1N(n3770), .Y(
        \i_MIPS/Register/n994 ) );
  OAI2BB2XL U9466 ( .B0(n3669), .B1(n3768), .A0N(
        \i_MIPS/Register/register[4][3] ), .A1N(n3770), .Y(
        \i_MIPS/Register/n983 ) );
  OAI2BB2XL U9467 ( .B0(n3656), .B1(n3763), .A0N(
        \i_MIPS/Register/register[6][17] ), .A1N(n3762), .Y(
        \i_MIPS/Register/n933 ) );
  OAI2BB2XL U9468 ( .B0(n3648), .B1(n3763), .A0N(
        \i_MIPS/Register/register[6][14] ), .A1N(n3764), .Y(
        \i_MIPS/Register/n930 ) );
  OAI2BB2XL U9469 ( .B0(n3669), .B1(n3762), .A0N(
        \i_MIPS/Register/register[6][3] ), .A1N(n3764), .Y(
        \i_MIPS/Register/n919 ) );
  OAI2BB2XL U9470 ( .B0(n3656), .B1(n3760), .A0N(
        \i_MIPS/Register/register[7][17] ), .A1N(n3760), .Y(
        \i_MIPS/Register/n901 ) );
  OAI2BB2XL U9471 ( .B0(n3648), .B1(n3760), .A0N(
        \i_MIPS/Register/register[7][14] ), .A1N(n3761), .Y(
        \i_MIPS/Register/n898 ) );
  OAI2BB2XL U9472 ( .B0(n3669), .B1(n3759), .A0N(
        \i_MIPS/Register/register[7][3] ), .A1N(n3761), .Y(
        \i_MIPS/Register/n887 ) );
  OAI2BB2XL U9473 ( .B0(n3656), .B1(n3757), .A0N(
        \i_MIPS/Register/register[8][17] ), .A1N(n3756), .Y(
        \i_MIPS/Register/n869 ) );
  OAI2BB2XL U9474 ( .B0(n3648), .B1(n3757), .A0N(
        \i_MIPS/Register/register[8][14] ), .A1N(n3758), .Y(
        \i_MIPS/Register/n866 ) );
  OAI2BB2XL U9475 ( .B0(n3669), .B1(n3756), .A0N(
        \i_MIPS/Register/register[8][3] ), .A1N(n3758), .Y(
        \i_MIPS/Register/n855 ) );
  OAI2BB2XL U9476 ( .B0(n3656), .B1(n3754), .A0N(
        \i_MIPS/Register/register[9][17] ), .A1N(n3754), .Y(
        \i_MIPS/Register/n837 ) );
  OAI2BB2XL U9477 ( .B0(n3648), .B1(n3754), .A0N(
        \i_MIPS/Register/register[9][14] ), .A1N(n3755), .Y(
        \i_MIPS/Register/n834 ) );
  OAI2BB2XL U9478 ( .B0(n3669), .B1(n3753), .A0N(
        \i_MIPS/Register/register[9][3] ), .A1N(n3755), .Y(
        \i_MIPS/Register/n823 ) );
  OAI2BB2XL U9479 ( .B0(n3656), .B1(n3751), .A0N(
        \i_MIPS/Register/register[10][17] ), .A1N(n3751), .Y(
        \i_MIPS/Register/n805 ) );
  OAI2BB2XL U9480 ( .B0(n3648), .B1(n3751), .A0N(
        \i_MIPS/Register/register[10][14] ), .A1N(n3752), .Y(
        \i_MIPS/Register/n802 ) );
  OAI2BB2XL U9481 ( .B0(n3669), .B1(n3750), .A0N(
        \i_MIPS/Register/register[10][3] ), .A1N(n3752), .Y(
        \i_MIPS/Register/n791 ) );
  OAI2BB2XL U9482 ( .B0(n3656), .B1(n3748), .A0N(
        \i_MIPS/Register/register[11][17] ), .A1N(n3748), .Y(
        \i_MIPS/Register/n773 ) );
  OAI2BB2XL U9483 ( .B0(n3648), .B1(n3748), .A0N(
        \i_MIPS/Register/register[11][14] ), .A1N(n3749), .Y(
        \i_MIPS/Register/n770 ) );
  OAI2BB2XL U9484 ( .B0(n3669), .B1(n3747), .A0N(
        \i_MIPS/Register/register[11][3] ), .A1N(n3749), .Y(
        \i_MIPS/Register/n759 ) );
  OAI2BB2XL U9485 ( .B0(n3656), .B1(n3745), .A0N(
        \i_MIPS/Register/register[12][17] ), .A1N(n3745), .Y(
        \i_MIPS/Register/n741 ) );
  OAI2BB2XL U9486 ( .B0(n3648), .B1(n3745), .A0N(
        \i_MIPS/Register/register[12][14] ), .A1N(n3746), .Y(
        \i_MIPS/Register/n738 ) );
  OAI2BB2XL U9487 ( .B0(n3669), .B1(n3744), .A0N(
        \i_MIPS/Register/register[12][3] ), .A1N(n3746), .Y(
        \i_MIPS/Register/n727 ) );
  OAI2BB2XL U9488 ( .B0(n3656), .B1(n3742), .A0N(
        \i_MIPS/Register/register[13][17] ), .A1N(n3742), .Y(
        \i_MIPS/Register/n709 ) );
  OAI2BB2XL U9489 ( .B0(n3648), .B1(n3742), .A0N(
        \i_MIPS/Register/register[13][14] ), .A1N(n3743), .Y(
        \i_MIPS/Register/n706 ) );
  OAI2BB2XL U9490 ( .B0(n3669), .B1(n3741), .A0N(
        \i_MIPS/Register/register[13][3] ), .A1N(n3743), .Y(
        \i_MIPS/Register/n695 ) );
  OAI2BB2XL U9491 ( .B0(n3656), .B1(n3739), .A0N(
        \i_MIPS/Register/register[14][17] ), .A1N(n3739), .Y(
        \i_MIPS/Register/n677 ) );
  OAI2BB2XL U9492 ( .B0(n3648), .B1(n3739), .A0N(
        \i_MIPS/Register/register[14][14] ), .A1N(n3740), .Y(
        \i_MIPS/Register/n674 ) );
  OAI2BB2XL U9493 ( .B0(n3669), .B1(n3738), .A0N(
        \i_MIPS/Register/register[14][3] ), .A1N(n3740), .Y(
        \i_MIPS/Register/n663 ) );
  OAI2BB2XL U9494 ( .B0(n3656), .B1(n3736), .A0N(
        \i_MIPS/Register/register[15][17] ), .A1N(n3736), .Y(
        \i_MIPS/Register/n645 ) );
  OAI2BB2XL U9495 ( .B0(n3648), .B1(n3736), .A0N(
        \i_MIPS/Register/register[15][14] ), .A1N(n3737), .Y(
        \i_MIPS/Register/n642 ) );
  OAI2BB2XL U9496 ( .B0(n3669), .B1(n3735), .A0N(
        \i_MIPS/Register/register[15][3] ), .A1N(n3737), .Y(
        \i_MIPS/Register/n631 ) );
  OAI2BB2XL U9497 ( .B0(n3656), .B1(n3733), .A0N(
        \i_MIPS/Register/register[16][17] ), .A1N(n3732), .Y(
        \i_MIPS/Register/n613 ) );
  OAI2BB2XL U9498 ( .B0(n3649), .B1(n3733), .A0N(
        \i_MIPS/Register/register[16][14] ), .A1N(n3734), .Y(
        \i_MIPS/Register/n610 ) );
  OAI2BB2XL U9499 ( .B0(n3670), .B1(n3732), .A0N(
        \i_MIPS/Register/register[16][3] ), .A1N(n3734), .Y(
        \i_MIPS/Register/n599 ) );
  OAI2BB2XL U9500 ( .B0(n3656), .B1(n3730), .A0N(
        \i_MIPS/Register/register[17][17] ), .A1N(n3729), .Y(
        \i_MIPS/Register/n581 ) );
  OAI2BB2XL U9501 ( .B0(n3649), .B1(n3730), .A0N(
        \i_MIPS/Register/register[17][14] ), .A1N(n3731), .Y(
        \i_MIPS/Register/n578 ) );
  OAI2BB2XL U9502 ( .B0(n3670), .B1(n3729), .A0N(
        \i_MIPS/Register/register[17][3] ), .A1N(n3731), .Y(
        \i_MIPS/Register/n567 ) );
  OAI2BB2XL U9503 ( .B0(n3656), .B1(n3691), .A0N(
        \i_MIPS/Register/register[30][17] ), .A1N(n3691), .Y(
        \i_MIPS/Register/n165 ) );
  OAI2BB2XL U9504 ( .B0(n3649), .B1(n3691), .A0N(
        \i_MIPS/Register/register[30][14] ), .A1N(n3692), .Y(
        \i_MIPS/Register/n162 ) );
  OAI2BB2XL U9505 ( .B0(n3670), .B1(n3690), .A0N(
        \i_MIPS/Register/register[30][3] ), .A1N(n3692), .Y(
        \i_MIPS/Register/n151 ) );
  OAI2BB2XL U9506 ( .B0(n3655), .B1(n3778), .A0N(
        \i_MIPS/Register/register[1][17] ), .A1N(n3777), .Y(
        \i_MIPS/Register/n1093 ) );
  OAI2BB2XL U9507 ( .B0(n3649), .B1(n3778), .A0N(
        \i_MIPS/Register/register[1][14] ), .A1N(n3779), .Y(
        \i_MIPS/Register/n1090 ) );
  OAI2BB2XL U9508 ( .B0(n3670), .B1(n3777), .A0N(
        \i_MIPS/Register/register[1][3] ), .A1N(n3779), .Y(
        \i_MIPS/Register/n1079 ) );
  OAI2BB2XL U9509 ( .B0(n3655), .B1(n3772), .A0N(
        \i_MIPS/Register/register[3][17] ), .A1N(n3771), .Y(
        \i_MIPS/Register/n1029 ) );
  OAI2BB2XL U9510 ( .B0(n3649), .B1(n3772), .A0N(
        \i_MIPS/Register/register[3][14] ), .A1N(n3773), .Y(
        \i_MIPS/Register/n1026 ) );
  OAI2BB2XL U9511 ( .B0(n3670), .B1(n3771), .A0N(
        \i_MIPS/Register/register[3][3] ), .A1N(n3773), .Y(
        \i_MIPS/Register/n1015 ) );
  OAI2BB2XL U9512 ( .B0(n3655), .B1(n3766), .A0N(
        \i_MIPS/Register/register[5][17] ), .A1N(n3765), .Y(
        \i_MIPS/Register/n965 ) );
  OAI2BB2XL U9513 ( .B0(n3649), .B1(n3766), .A0N(
        \i_MIPS/Register/register[5][14] ), .A1N(n3767), .Y(
        \i_MIPS/Register/n962 ) );
  OAI2BB2XL U9514 ( .B0(n3670), .B1(n3765), .A0N(
        \i_MIPS/Register/register[5][3] ), .A1N(n3767), .Y(
        \i_MIPS/Register/n951 ) );
  OAI2BB2XL U9515 ( .B0(n3655), .B1(n3727), .A0N(
        \i_MIPS/Register/register[18][17] ), .A1N(n3727), .Y(
        \i_MIPS/Register/n549 ) );
  OAI2BB2XL U9516 ( .B0(n3649), .B1(n3727), .A0N(
        \i_MIPS/Register/register[18][14] ), .A1N(n3728), .Y(
        \i_MIPS/Register/n546 ) );
  OAI2BB2XL U9517 ( .B0(n3670), .B1(n3726), .A0N(
        \i_MIPS/Register/register[18][3] ), .A1N(n3728), .Y(
        \i_MIPS/Register/n535 ) );
  OAI2BB2XL U9518 ( .B0(n3655), .B1(n3724), .A0N(
        \i_MIPS/Register/register[19][17] ), .A1N(n3724), .Y(
        \i_MIPS/Register/n517 ) );
  OAI2BB2XL U9519 ( .B0(n3649), .B1(n3724), .A0N(
        \i_MIPS/Register/register[19][14] ), .A1N(n3725), .Y(
        \i_MIPS/Register/n514 ) );
  OAI2BB2XL U9520 ( .B0(n3670), .B1(n3723), .A0N(
        \i_MIPS/Register/register[19][3] ), .A1N(n3725), .Y(
        \i_MIPS/Register/n503 ) );
  OAI2BB2XL U9521 ( .B0(n3655), .B1(n3721), .A0N(
        \i_MIPS/Register/register[20][17] ), .A1N(n3721), .Y(
        \i_MIPS/Register/n485 ) );
  OAI2BB2XL U9522 ( .B0(n3649), .B1(n3721), .A0N(
        \i_MIPS/Register/register[20][14] ), .A1N(n3722), .Y(
        \i_MIPS/Register/n482 ) );
  OAI2BB2XL U9523 ( .B0(n3670), .B1(n3720), .A0N(
        \i_MIPS/Register/register[20][3] ), .A1N(n3722), .Y(
        \i_MIPS/Register/n471 ) );
  OAI2BB2XL U9524 ( .B0(n3655), .B1(n3718), .A0N(
        \i_MIPS/Register/register[21][17] ), .A1N(n3718), .Y(
        \i_MIPS/Register/n453 ) );
  OAI2BB2XL U9525 ( .B0(n3649), .B1(n3718), .A0N(
        \i_MIPS/Register/register[21][14] ), .A1N(n3719), .Y(
        \i_MIPS/Register/n450 ) );
  OAI2BB2XL U9526 ( .B0(n3670), .B1(n3717), .A0N(
        \i_MIPS/Register/register[21][3] ), .A1N(n3719), .Y(
        \i_MIPS/Register/n439 ) );
  OAI2BB2XL U9527 ( .B0(n3655), .B1(n3715), .A0N(
        \i_MIPS/Register/register[22][17] ), .A1N(n3715), .Y(
        \i_MIPS/Register/n421 ) );
  OAI2BB2XL U9528 ( .B0(n3649), .B1(n3715), .A0N(
        \i_MIPS/Register/register[22][14] ), .A1N(n3716), .Y(
        \i_MIPS/Register/n418 ) );
  OAI2BB2XL U9529 ( .B0(n3670), .B1(n3714), .A0N(
        \i_MIPS/Register/register[22][3] ), .A1N(n3716), .Y(
        \i_MIPS/Register/n407 ) );
  OAI2BB2XL U9530 ( .B0(n3655), .B1(n3712), .A0N(
        \i_MIPS/Register/register[23][17] ), .A1N(n3712), .Y(
        \i_MIPS/Register/n389 ) );
  OAI2BB2XL U9531 ( .B0(n3649), .B1(n3712), .A0N(
        \i_MIPS/Register/register[23][14] ), .A1N(n3713), .Y(
        \i_MIPS/Register/n386 ) );
  OAI2BB2XL U9532 ( .B0(n3670), .B1(n3711), .A0N(
        \i_MIPS/Register/register[23][3] ), .A1N(n3713), .Y(
        \i_MIPS/Register/n375 ) );
  OAI2BB2XL U9533 ( .B0(n3655), .B1(n3709), .A0N(
        \i_MIPS/Register/register[24][17] ), .A1N(n3709), .Y(
        \i_MIPS/Register/n357 ) );
  OAI2BB2XL U9534 ( .B0(n3649), .B1(n3709), .A0N(
        \i_MIPS/Register/register[24][14] ), .A1N(n3710), .Y(
        \i_MIPS/Register/n354 ) );
  OAI2BB2XL U9535 ( .B0(n3670), .B1(n3708), .A0N(
        \i_MIPS/Register/register[24][3] ), .A1N(n3710), .Y(
        \i_MIPS/Register/n343 ) );
  OAI2BB2XL U9536 ( .B0(n3655), .B1(n3706), .A0N(
        \i_MIPS/Register/register[25][17] ), .A1N(n3706), .Y(
        \i_MIPS/Register/n325 ) );
  OAI2BB2XL U9537 ( .B0(n3649), .B1(n3706), .A0N(
        \i_MIPS/Register/register[25][14] ), .A1N(n3707), .Y(
        \i_MIPS/Register/n322 ) );
  OAI2BB2XL U9538 ( .B0(n3670), .B1(n3705), .A0N(
        \i_MIPS/Register/register[25][3] ), .A1N(n3707), .Y(
        \i_MIPS/Register/n311 ) );
  OAI2BB2XL U9539 ( .B0(n3655), .B1(n3703), .A0N(
        \i_MIPS/Register/register[26][17] ), .A1N(n3703), .Y(
        \i_MIPS/Register/n293 ) );
  OAI2BB2XL U9540 ( .B0(n3649), .B1(n3703), .A0N(
        \i_MIPS/Register/register[26][14] ), .A1N(n3704), .Y(
        \i_MIPS/Register/n290 ) );
  OAI2BB2XL U9541 ( .B0(n3670), .B1(n3702), .A0N(
        \i_MIPS/Register/register[26][3] ), .A1N(n3704), .Y(
        \i_MIPS/Register/n279 ) );
  OAI2BB2XL U9542 ( .B0(n3655), .B1(n3700), .A0N(
        \i_MIPS/Register/register[27][17] ), .A1N(n3700), .Y(
        \i_MIPS/Register/n261 ) );
  OAI2BB2XL U9543 ( .B0(n3649), .B1(n3700), .A0N(
        \i_MIPS/Register/register[27][14] ), .A1N(n3701), .Y(
        \i_MIPS/Register/n258 ) );
  OAI2BB2XL U9544 ( .B0(n3670), .B1(n3699), .A0N(
        \i_MIPS/Register/register[27][3] ), .A1N(n3701), .Y(
        \i_MIPS/Register/n247 ) );
  OAI2BB2XL U9545 ( .B0(n3655), .B1(n3697), .A0N(
        \i_MIPS/Register/register[28][17] ), .A1N(n3697), .Y(
        \i_MIPS/Register/n229 ) );
  OAI2BB2XL U9546 ( .B0(n3649), .B1(n3697), .A0N(
        \i_MIPS/Register/register[28][14] ), .A1N(n3698), .Y(
        \i_MIPS/Register/n226 ) );
  OAI2BB2XL U9547 ( .B0(n3670), .B1(n3696), .A0N(
        \i_MIPS/Register/register[28][3] ), .A1N(n3698), .Y(
        \i_MIPS/Register/n215 ) );
  OAI2BB2XL U9548 ( .B0(n3655), .B1(n3694), .A0N(
        \i_MIPS/Register/register[29][17] ), .A1N(n3694), .Y(
        \i_MIPS/Register/n197 ) );
  OAI2BB2XL U9549 ( .B0(n3649), .B1(n3694), .A0N(
        \i_MIPS/Register/register[29][14] ), .A1N(n3695), .Y(
        \i_MIPS/Register/n194 ) );
  OAI2BB2XL U9550 ( .B0(n3670), .B1(n3693), .A0N(
        \i_MIPS/Register/register[29][3] ), .A1N(n3695), .Y(
        \i_MIPS/Register/n183 ) );
  OAI2BB2XL U9551 ( .B0(n3661), .B1(n3769), .A0N(
        \i_MIPS/Register/register[4][18] ), .A1N(n3770), .Y(
        \i_MIPS/Register/n998 ) );
  OAI2BB2XL U9552 ( .B0(n3663), .B1(n3768), .A0N(
        \i_MIPS/Register/register[4][2] ), .A1N(n3769), .Y(
        \i_MIPS/Register/n982 ) );
  OAI2BB2XL U9553 ( .B0(n3661), .B1(n3766), .A0N(
        \i_MIPS/Register/register[5][18] ), .A1N(n3767), .Y(
        \i_MIPS/Register/n966 ) );
  OAI2BB2XL U9554 ( .B0(n3663), .B1(n3765), .A0N(
        \i_MIPS/Register/register[5][2] ), .A1N(n3766), .Y(
        \i_MIPS/Register/n950 ) );
  OAI2BB2XL U9555 ( .B0(n3661), .B1(n3763), .A0N(
        \i_MIPS/Register/register[6][18] ), .A1N(n3764), .Y(
        \i_MIPS/Register/n934 ) );
  OAI2BB2XL U9556 ( .B0(n3663), .B1(n3762), .A0N(
        \i_MIPS/Register/register[6][2] ), .A1N(n3763), .Y(
        \i_MIPS/Register/n918 ) );
  OAI2BB2XL U9557 ( .B0(n3687), .B1(n3768), .A0N(
        \i_MIPS/Register/register[4][8] ), .A1N(n3770), .Y(
        \i_MIPS/Register/n988 ) );
  OAI2BB2XL U9558 ( .B0(n3687), .B1(n3765), .A0N(
        \i_MIPS/Register/register[5][8] ), .A1N(n3767), .Y(
        \i_MIPS/Register/n956 ) );
  OAI2BB2XL U9559 ( .B0(n3687), .B1(n3762), .A0N(
        \i_MIPS/Register/register[6][8] ), .A1N(n3764), .Y(
        \i_MIPS/Register/n924 ) );
  OAI21XL U9560 ( .A0(n8808), .A1(n8809), .B0(mem_ready_D), .Y(\D_cache/n247 )
         );
  MXI2X1 U9561 ( .A(\i_MIPS/n359 ), .B(n8248), .S0(n3618), .Y(\i_MIPS/n550 )
         );
  OAI2BB2XL U9562 ( .B0(n3660), .B1(n3780), .A0N(
        \i_MIPS/Register/register[0][23] ), .A1N(n3780), .Y(
        \i_MIPS/Register/n1131 ) );
  OAI2BB2XL U9563 ( .B0(n3017), .B1(n3781), .A0N(
        \i_MIPS/Register/register[0][22] ), .A1N(n3782), .Y(
        \i_MIPS/Register/n1130 ) );
  OAI2BB2XL U9564 ( .B0(n3660), .B1(n3777), .A0N(
        \i_MIPS/Register/register[1][23] ), .A1N(n3779), .Y(
        \i_MIPS/Register/n1099 ) );
  OAI2BB2XL U9565 ( .B0(n3017), .B1(n3778), .A0N(
        \i_MIPS/Register/register[1][22] ), .A1N(n3779), .Y(
        \i_MIPS/Register/n1098 ) );
  OAI2BB2XL U9566 ( .B0(n3660), .B1(n3774), .A0N(
        \i_MIPS/Register/register[2][23] ), .A1N(n3776), .Y(
        \i_MIPS/Register/n1067 ) );
  OAI2BB2XL U9567 ( .B0(n3017), .B1(n3775), .A0N(
        \i_MIPS/Register/register[2][22] ), .A1N(n3776), .Y(
        \i_MIPS/Register/n1066 ) );
  OAI2BB2XL U9568 ( .B0(n3660), .B1(n3768), .A0N(
        \i_MIPS/Register/register[4][23] ), .A1N(n3770), .Y(
        \i_MIPS/Register/n1003 ) );
  OAI2BB2XL U9569 ( .B0(n3017), .B1(n3769), .A0N(
        \i_MIPS/Register/register[4][22] ), .A1N(n3770), .Y(
        \i_MIPS/Register/n1002 ) );
  MXI2X1 U9570 ( .A(\i_MIPS/n363 ), .B(n8232), .S0(n3619), .Y(\i_MIPS/n554 )
         );
  NAND4BX1 U9571 ( .AN(n6174), .B(n6173), .C(n6172), .D(n6171), .Y(n6185) );
  OA22X1 U9572 ( .A0(\i_MIPS/Register/register[4][8] ), .A1(n3180), .B0(
        \i_MIPS/Register/register[12][8] ), .B1(n3177), .Y(n6173) );
  OA22X1 U9573 ( .A0(\i_MIPS/Register/register[0][8] ), .A1(n3186), .B0(
        \i_MIPS/Register/register[8][8] ), .B1(n3183), .Y(n6172) );
  OAI221XL U9574 ( .A0(\i_MIPS/Register/register[2][8] ), .A1(n3174), .B0(
        \i_MIPS/Register/register[10][8] ), .B1(n16), .C0(n6166), .Y(n6174) );
  NAND4BX1 U9575 ( .AN(n5305), .B(n5304), .C(n5303), .D(n5302), .Y(n5316) );
  OA22X1 U9576 ( .A0(\i_MIPS/Register/register[4][11] ), .A1(n3180), .B0(
        \i_MIPS/Register/register[12][11] ), .B1(n3176), .Y(n5304) );
  OA22X1 U9577 ( .A0(\i_MIPS/Register/register[0][11] ), .A1(n3185), .B0(
        \i_MIPS/Register/register[8][11] ), .B1(n3182), .Y(n5303) );
  OAI221XL U9578 ( .A0(\i_MIPS/Register/register[2][11] ), .A1(n3173), .B0(
        \i_MIPS/Register/register[10][11] ), .B1(n16), .C0(n5297), .Y(n5305)
         );
  NAND4BX1 U9579 ( .AN(n6513), .B(n6512), .C(n6511), .D(n6510), .Y(n6524) );
  OAI221XL U9580 ( .A0(\i_MIPS/Register/register[2][21] ), .A1(n3175), .B0(
        \i_MIPS/Register/register[10][21] ), .B1(n16), .C0(n6505), .Y(n6513)
         );
  NAND4BX1 U9581 ( .AN(n6183), .B(n6182), .C(n6181), .D(n6180), .Y(n6184) );
  OA22X1 U9582 ( .A0(\i_MIPS/Register/register[20][8] ), .A1(n3181), .B0(
        \i_MIPS/Register/register[28][8] ), .B1(n3178), .Y(n6182) );
  OA22X1 U9583 ( .A0(\i_MIPS/Register/register[16][8] ), .A1(n3187), .B0(
        \i_MIPS/Register/register[24][8] ), .B1(n3184), .Y(n6181) );
  OAI221XL U9584 ( .A0(\i_MIPS/Register/register[18][8] ), .A1(n3175), .B0(
        \i_MIPS/Register/register[26][8] ), .B1(n16), .C0(n6175), .Y(n6183) );
  NAND4BX1 U9585 ( .AN(n5314), .B(n5313), .C(n5312), .D(n5311), .Y(n5315) );
  OA22X1 U9586 ( .A0(\i_MIPS/Register/register[20][11] ), .A1(n3180), .B0(
        \i_MIPS/Register/register[28][11] ), .B1(n3176), .Y(n5313) );
  OA22X1 U9587 ( .A0(\i_MIPS/Register/register[16][11] ), .A1(n3185), .B0(
        \i_MIPS/Register/register[24][11] ), .B1(n3182), .Y(n5312) );
  OAI221XL U9588 ( .A0(\i_MIPS/Register/register[18][11] ), .A1(n3173), .B0(
        \i_MIPS/Register/register[26][11] ), .B1(n16), .C0(n5306), .Y(n5314)
         );
  NAND4BX1 U9589 ( .AN(n6315), .B(n6314), .C(n6313), .D(n6312), .Y(n6316) );
  OAI221XL U9590 ( .A0(\i_MIPS/Register/register[18][12] ), .A1(n3175), .B0(
        \i_MIPS/Register/register[26][12] ), .B1(n16), .C0(n6307), .Y(n6315)
         );
  NAND4BX1 U9591 ( .AN(n6294), .B(n6293), .C(n6292), .D(n6291), .Y(n6295) );
  OAI221XL U9592 ( .A0(\i_MIPS/Register/register[18][12] ), .A1(n3123), .B0(
        \i_MIPS/Register/register[26][12] ), .B1(n3121), .C0(n6286), .Y(n6294)
         );
  NAND4BX1 U9593 ( .AN(n6450), .B(n6449), .C(n6448), .D(n6447), .Y(n6451) );
  OAI221XL U9594 ( .A0(\i_MIPS/Register/register[18][13] ), .A1(n3175), .B0(
        \i_MIPS/Register/register[26][13] ), .B1(n16), .C0(n6442), .Y(n6450)
         );
  NAND4BX1 U9595 ( .AN(n5354), .B(n5353), .C(n5352), .D(n5351), .Y(n5355) );
  OAI221XL U9596 ( .A0(\i_MIPS/Register/register[18][4] ), .A1(n3123), .B0(
        \i_MIPS/Register/register[26][4] ), .B1(n2790), .C0(n5346), .Y(n5354)
         );
  NAND4BX1 U9597 ( .AN(n5080), .B(n5079), .C(n5078), .D(n5077), .Y(n5081) );
  OAI221XL U9598 ( .A0(\i_MIPS/Register/register[18][0] ), .A1(n3122), .B0(
        \i_MIPS/Register/register[26][0] ), .B1(n3119), .C0(n5072), .Y(n5080)
         );
  NAND4BX1 U9599 ( .AN(n6252), .B(n6251), .C(n6250), .D(n6249), .Y(n6253) );
  OA22X1 U9600 ( .A0(\i_MIPS/Register/register[20][9] ), .A1(n2786), .B0(
        \i_MIPS/Register/register[28][9] ), .B1(n3178), .Y(n6251) );
  OA22X1 U9601 ( .A0(\i_MIPS/Register/register[16][9] ), .A1(n3187), .B0(
        \i_MIPS/Register/register[24][9] ), .B1(n3184), .Y(n6250) );
  OAI221XL U9602 ( .A0(\i_MIPS/Register/register[18][9] ), .A1(n3175), .B0(
        \i_MIPS/Register/register[26][9] ), .B1(n16), .C0(n6244), .Y(n6252) );
  NAND4BX1 U9603 ( .AN(n6522), .B(n6521), .C(n6520), .D(n6519), .Y(n6523) );
  OAI221XL U9604 ( .A0(\i_MIPS/Register/register[18][21] ), .A1(n3175), .B0(
        \i_MIPS/Register/register[26][21] ), .B1(n16), .C0(n6514), .Y(n6522)
         );
  NAND4BX1 U9605 ( .AN(n6967), .B(n6966), .C(n6965), .D(n6964), .Y(n6968) );
  OA22X1 U9606 ( .A0(\i_MIPS/Register/register[20][16] ), .A1(n2789), .B0(
        \i_MIPS/Register/register[28][16] ), .B1(n2787), .Y(n6966) );
  OA22X1 U9607 ( .A0(\i_MIPS/Register/register[16][16] ), .A1(n3136), .B0(
        \i_MIPS/Register/register[24][16] ), .B1(n2788), .Y(n6965) );
  OAI221XL U9608 ( .A0(\i_MIPS/Register/register[18][16] ), .A1(n2791), .B0(
        \i_MIPS/Register/register[26][16] ), .B1(n3119), .C0(n6959), .Y(n6967)
         );
  NAND4BX1 U9609 ( .AN(n6743), .B(n6742), .C(n6741), .D(n6740), .Y(n6744) );
  OAI221XL U9610 ( .A0(\i_MIPS/Register/register[18][22] ), .A1(n3123), .B0(
        \i_MIPS/Register/register[26][22] ), .B1(n3119), .C0(n6735), .Y(n6743)
         );
  NAND4BX1 U9611 ( .AN(n6898), .B(n6897), .C(n6896), .D(n6895), .Y(n6899) );
  OA22X1 U9612 ( .A0(\i_MIPS/Register/register[20][23] ), .A1(n2789), .B0(
        \i_MIPS/Register/register[28][23] ), .B1(n3125), .Y(n6897) );
  OA22X1 U9613 ( .A0(\i_MIPS/Register/register[16][23] ), .A1(n3135), .B0(
        \i_MIPS/Register/register[24][23] ), .B1(n3131), .Y(n6896) );
  OAI221XL U9614 ( .A0(\i_MIPS/Register/register[18][23] ), .A1(n3124), .B0(
        \i_MIPS/Register/register[26][23] ), .B1(n3121), .C0(n6890), .Y(n6898)
         );
  NAND4BX1 U9615 ( .AN(n4886), .B(n4885), .C(n4884), .D(n4883), .Y(n4887) );
  OAI221XL U9616 ( .A0(\i_MIPS/Register/register[18][20] ), .A1(n3122), .B0(
        \i_MIPS/Register/register[26][20] ), .B1(n3119), .C0(n4878), .Y(n4886)
         );
  NAND4BX1 U9617 ( .AN(n5778), .B(n5777), .C(n5776), .D(n5775), .Y(n5779) );
  OAI221XL U9618 ( .A0(\i_MIPS/Register/register[18][18] ), .A1(n3124), .B0(
        \i_MIPS/Register/register[26][18] ), .B1(n3120), .C0(n5770), .Y(n5778)
         );
  NAND4BX1 U9619 ( .AN(n5706), .B(n5705), .C(n5704), .D(n5703), .Y(n5707) );
  OA22X1 U9620 ( .A0(\i_MIPS/Register/register[20][17] ), .A1(n3130), .B0(
        \i_MIPS/Register/register[28][17] ), .B1(n3127), .Y(n5705) );
  OA22X1 U9621 ( .A0(\i_MIPS/Register/register[16][17] ), .A1(n3136), .B0(
        \i_MIPS/Register/register[24][17] ), .B1(n3132), .Y(n5704) );
  OAI221XL U9622 ( .A0(\i_MIPS/Register/register[18][17] ), .A1(n3124), .B0(
        \i_MIPS/Register/register[26][17] ), .B1(n3120), .C0(n5698), .Y(n5706)
         );
  MXI2X1 U9623 ( .A(\i_MIPS/n336 ), .B(\i_MIPS/n337 ), .S0(n3618), .Y(
        \i_MIPS/n526 ) );
  OAI2BB2XL U9624 ( .B0(n3658), .B1(n3760), .A0N(
        \i_MIPS/Register/register[7][16] ), .A1N(n3761), .Y(
        \i_MIPS/Register/n900 ) );
  OAI2BB2XL U9625 ( .B0(n3658), .B1(n3757), .A0N(
        \i_MIPS/Register/register[8][16] ), .A1N(n3758), .Y(
        \i_MIPS/Register/n868 ) );
  OAI2BB2XL U9626 ( .B0(n3658), .B1(n3754), .A0N(
        \i_MIPS/Register/register[9][16] ), .A1N(n3755), .Y(
        \i_MIPS/Register/n836 ) );
  OAI2BB2XL U9627 ( .B0(n3658), .B1(n3751), .A0N(
        \i_MIPS/Register/register[10][16] ), .A1N(n3752), .Y(
        \i_MIPS/Register/n804 ) );
  OAI2BB2XL U9628 ( .B0(n3658), .B1(n3748), .A0N(
        \i_MIPS/Register/register[11][16] ), .A1N(n3749), .Y(
        \i_MIPS/Register/n772 ) );
  OAI2BB2XL U9629 ( .B0(n3658), .B1(n3745), .A0N(
        \i_MIPS/Register/register[12][16] ), .A1N(n3746), .Y(
        \i_MIPS/Register/n740 ) );
  OAI2BB2XL U9630 ( .B0(n3658), .B1(n3742), .A0N(
        \i_MIPS/Register/register[13][16] ), .A1N(n3743), .Y(
        \i_MIPS/Register/n708 ) );
  OAI2BB2XL U9631 ( .B0(n3658), .B1(n3739), .A0N(
        \i_MIPS/Register/register[14][16] ), .A1N(n3740), .Y(
        \i_MIPS/Register/n676 ) );
  OAI2BB2XL U9632 ( .B0(n3658), .B1(n3736), .A0N(
        \i_MIPS/Register/register[15][16] ), .A1N(n3737), .Y(
        \i_MIPS/Register/n644 ) );
  OAI2BB2XL U9633 ( .B0(n3658), .B1(n3733), .A0N(
        \i_MIPS/Register/register[16][16] ), .A1N(n3734), .Y(
        \i_MIPS/Register/n612 ) );
  OAI2BB2XL U9634 ( .B0(n3658), .B1(n3730), .A0N(
        \i_MIPS/Register/register[17][16] ), .A1N(n3731), .Y(
        \i_MIPS/Register/n580 ) );
  OAI2BB2XL U9635 ( .B0(n3658), .B1(n3691), .A0N(
        \i_MIPS/Register/register[30][16] ), .A1N(n3692), .Y(
        \i_MIPS/Register/n164 ) );
  OAI2BB2XL U9636 ( .B0(n3647), .B1(n3760), .A0N(
        \i_MIPS/Register/register[7][15] ), .A1N(n3759), .Y(
        \i_MIPS/Register/n899 ) );
  OAI2BB2XL U9637 ( .B0(n3646), .B1(n3757), .A0N(
        \i_MIPS/Register/register[8][15] ), .A1N(n3758), .Y(
        \i_MIPS/Register/n867 ) );
  OAI2BB2XL U9638 ( .B0(n3646), .B1(n3754), .A0N(
        \i_MIPS/Register/register[9][15] ), .A1N(n3755), .Y(
        \i_MIPS/Register/n835 ) );
  OAI2BB2XL U9639 ( .B0(n3646), .B1(n3751), .A0N(
        \i_MIPS/Register/register[10][15] ), .A1N(n3752), .Y(
        \i_MIPS/Register/n803 ) );
  OAI2BB2XL U9640 ( .B0(n3646), .B1(n3748), .A0N(
        \i_MIPS/Register/register[11][15] ), .A1N(n3749), .Y(
        \i_MIPS/Register/n771 ) );
  OAI2BB2XL U9641 ( .B0(n3646), .B1(n3745), .A0N(
        \i_MIPS/Register/register[12][15] ), .A1N(n3746), .Y(
        \i_MIPS/Register/n739 ) );
  OAI2BB2XL U9642 ( .B0(n3646), .B1(n3742), .A0N(
        \i_MIPS/Register/register[13][15] ), .A1N(n3743), .Y(
        \i_MIPS/Register/n707 ) );
  OAI2BB2XL U9643 ( .B0(n3646), .B1(n3739), .A0N(
        \i_MIPS/Register/register[14][15] ), .A1N(n3740), .Y(
        \i_MIPS/Register/n675 ) );
  OAI2BB2XL U9644 ( .B0(n3646), .B1(n3736), .A0N(
        \i_MIPS/Register/register[15][15] ), .A1N(n3737), .Y(
        \i_MIPS/Register/n643 ) );
  OAI2BB2XL U9645 ( .B0(n3646), .B1(n3733), .A0N(
        \i_MIPS/Register/register[16][15] ), .A1N(n3734), .Y(
        \i_MIPS/Register/n611 ) );
  OAI2BB2XL U9646 ( .B0(n3646), .B1(n3730), .A0N(
        \i_MIPS/Register/register[17][15] ), .A1N(n3731), .Y(
        \i_MIPS/Register/n579 ) );
  OAI2BB2XL U9647 ( .B0(n3646), .B1(n3691), .A0N(
        \i_MIPS/Register/register[30][15] ), .A1N(n3692), .Y(
        \i_MIPS/Register/n163 ) );
  OAI2BB2XL U9648 ( .B0(n3665), .B1(n3780), .A0N(
        \i_MIPS/Register/register[0][9] ), .A1N(n3782), .Y(
        \i_MIPS/Register/n1117 ) );
  OAI2BB2XL U9649 ( .B0(n3665), .B1(n3771), .A0N(
        \i_MIPS/Register/register[3][9] ), .A1N(n3773), .Y(
        \i_MIPS/Register/n1021 ) );
  OAI2BB2XL U9650 ( .B0(n3665), .B1(n3762), .A0N(
        \i_MIPS/Register/register[6][9] ), .A1N(n3764), .Y(
        \i_MIPS/Register/n925 ) );
  OAI2BB2XL U9651 ( .B0(n3665), .B1(n3744), .A0N(
        \i_MIPS/Register/register[12][9] ), .A1N(n3746), .Y(
        \i_MIPS/Register/n733 ) );
  OAI2BB2XL U9652 ( .B0(n3665), .B1(n3735), .A0N(
        \i_MIPS/Register/register[15][9] ), .A1N(n3737), .Y(
        \i_MIPS/Register/n637 ) );
  MXI2X1 U9653 ( .A(\i_MIPS/n290 ), .B(\i_MIPS/n291 ), .S0(n3619), .Y(
        \i_MIPS/n418 ) );
  MXI2X1 U9654 ( .A(\i_MIPS/n347 ), .B(n8128), .S0(n3618), .Y(\i_MIPS/n538 )
         );
  MXI2X1 U9655 ( .A(\i_MIPS/n346 ), .B(n8158), .S0(n3618), .Y(\i_MIPS/n537 )
         );
  MXI2X1 U9656 ( .A(\i_MIPS/n345 ), .B(n8264), .S0(n3618), .Y(\i_MIPS/n536 )
         );
  MXI2X1 U9657 ( .A(\i_MIPS/n364 ), .B(n8010), .S0(n3617), .Y(\i_MIPS/n555 )
         );
  MXI2X1 U9658 ( .A(\i_MIPS/n362 ), .B(n8245), .S0(n3619), .Y(\i_MIPS/n553 )
         );
  MXI2X1 U9659 ( .A(\i_MIPS/n361 ), .B(n8013), .S0(n3617), .Y(\i_MIPS/n552 )
         );
  MXI2X1 U9660 ( .A(\i_MIPS/n360 ), .B(n8247), .S0(n3618), .Y(\i_MIPS/n551 )
         );
  MXI2X1 U9661 ( .A(\i_MIPS/n352 ), .B(n8036), .S0(n3618), .Y(\i_MIPS/n543 )
         );
  MXI2X1 U9662 ( .A(\i_MIPS/n350 ), .B(n8416), .S0(n3617), .Y(\i_MIPS/n541 )
         );
  CLKINVX1 U9663 ( .A(n6048), .Y(n7007) );
  OAI221XL U9664 ( .A0(\i_MIPS/ALUin1[23] ), .A1(n3091), .B0(
        \i_MIPS/ALUin1[24] ), .B1(n3085), .C0(n6047), .Y(n6048) );
  OA22X1 U9665 ( .A0(\i_MIPS/ALUin1[25] ), .A1(n14), .B0(\i_MIPS/ALUin1[26] ), 
        .B1(n3078), .Y(n6047) );
  MXI2X1 U9666 ( .A(\i_MIPS/n340 ), .B(n8329), .S0(n3617), .Y(\i_MIPS/n531 )
         );
  OAI2BB2XL U9667 ( .B0(n3665), .B1(n3777), .A0N(
        \i_MIPS/Register/register[1][9] ), .A1N(n3779), .Y(
        \i_MIPS/Register/n1085 ) );
  OAI2BB2XL U9668 ( .B0(n3664), .B1(n3768), .A0N(
        \i_MIPS/Register/register[4][9] ), .A1N(n3770), .Y(
        \i_MIPS/Register/n989 ) );
  OAI2BB2XL U9669 ( .B0(n3664), .B1(n3741), .A0N(
        \i_MIPS/Register/register[13][9] ), .A1N(n3743), .Y(
        \i_MIPS/Register/n701 ) );
  OAI2BB2XL U9670 ( .B0(n3664), .B1(n3732), .A0N(
        \i_MIPS/Register/register[16][9] ), .A1N(n3734), .Y(
        \i_MIPS/Register/n605 ) );
  CLKINVX1 U9671 ( .A(n4982), .Y(n6529) );
  OAI221XL U9672 ( .A0(\i_MIPS/ALUin1[10] ), .A1(n3091), .B0(
        \i_MIPS/ALUin1[9] ), .B1(n3086), .C0(n4981), .Y(n4982) );
  OAI2BB2XL U9673 ( .B0(\D_cache/n240 ), .B1(n3794), .A0N(
        \D_cache/cache[7][133] ), .A1N(n3797), .Y(\D_cache/n725 ) );
  OAI2BB2XL U9674 ( .B0(\D_cache/n240 ), .B1(n3814), .A0N(
        \D_cache/cache[6][133] ), .A1N(n3817), .Y(\D_cache/n726 ) );
  OAI2BB2XL U9675 ( .B0(\D_cache/n240 ), .B1(n3832), .A0N(
        \D_cache/cache[5][133] ), .A1N(n3835), .Y(\D_cache/n727 ) );
  OAI2BB2XL U9676 ( .B0(\D_cache/n240 ), .B1(n3854), .A0N(
        \D_cache/cache[4][133] ), .A1N(n3857), .Y(\D_cache/n728 ) );
  OAI2BB2XL U9677 ( .B0(\D_cache/n240 ), .B1(n3873), .A0N(
        \D_cache/cache[3][133] ), .A1N(n3876), .Y(\D_cache/n729 ) );
  OAI2BB2XL U9678 ( .B0(\D_cache/n240 ), .B1(n3894), .A0N(
        \D_cache/cache[2][133] ), .A1N(n3897), .Y(\D_cache/n730 ) );
  OAI2BB2XL U9679 ( .B0(\D_cache/n240 ), .B1(n3915), .A0N(
        \D_cache/cache[1][133] ), .A1N(n3918), .Y(\D_cache/n731 ) );
  OAI2BB2XL U9680 ( .B0(\D_cache/n240 ), .B1(n3936), .A0N(
        \D_cache/cache[0][133] ), .A1N(n3939), .Y(\D_cache/n732 ) );
  OAI2BB2XL U9681 ( .B0(\D_cache/n239 ), .B1(n3793), .A0N(
        \D_cache/cache[7][134] ), .A1N(n3797), .Y(\D_cache/n717 ) );
  OAI2BB2XL U9682 ( .B0(\D_cache/n239 ), .B1(n3813), .A0N(
        \D_cache/cache[6][134] ), .A1N(n3817), .Y(\D_cache/n718 ) );
  OAI2BB2XL U9683 ( .B0(\D_cache/n239 ), .B1(n3831), .A0N(
        \D_cache/cache[5][134] ), .A1N(n3835), .Y(\D_cache/n719 ) );
  OAI2BB2XL U9684 ( .B0(\D_cache/n239 ), .B1(n3853), .A0N(
        \D_cache/cache[4][134] ), .A1N(n3857), .Y(\D_cache/n720 ) );
  OAI2BB2XL U9685 ( .B0(\D_cache/n239 ), .B1(n3872), .A0N(
        \D_cache/cache[3][134] ), .A1N(n3876), .Y(\D_cache/n721 ) );
  OAI2BB2XL U9686 ( .B0(\D_cache/n239 ), .B1(n3893), .A0N(
        \D_cache/cache[2][134] ), .A1N(n3897), .Y(\D_cache/n722 ) );
  OAI2BB2XL U9687 ( .B0(\D_cache/n239 ), .B1(n3914), .A0N(
        \D_cache/cache[1][134] ), .A1N(n3918), .Y(\D_cache/n723 ) );
  OAI2BB2XL U9688 ( .B0(\D_cache/n239 ), .B1(n3935), .A0N(
        \D_cache/cache[0][134] ), .A1N(n3939), .Y(\D_cache/n724 ) );
  OAI2BB2XL U9689 ( .B0(\D_cache/n235 ), .B1(n3794), .A0N(
        \D_cache/cache[7][138] ), .A1N(n3795), .Y(\D_cache/n685 ) );
  OAI2BB2XL U9690 ( .B0(\D_cache/n235 ), .B1(n3814), .A0N(
        \D_cache/cache[6][138] ), .A1N(n3815), .Y(\D_cache/n686 ) );
  OAI2BB2XL U9691 ( .B0(\D_cache/n235 ), .B1(n3832), .A0N(
        \D_cache/cache[5][138] ), .A1N(n3833), .Y(\D_cache/n687 ) );
  OAI2BB2XL U9692 ( .B0(\D_cache/n235 ), .B1(n3854), .A0N(
        \D_cache/cache[4][138] ), .A1N(n3855), .Y(\D_cache/n688 ) );
  OAI2BB2XL U9693 ( .B0(\D_cache/n235 ), .B1(n3873), .A0N(
        \D_cache/cache[3][138] ), .A1N(n3874), .Y(\D_cache/n689 ) );
  OAI2BB2XL U9694 ( .B0(\D_cache/n235 ), .B1(n3894), .A0N(
        \D_cache/cache[2][138] ), .A1N(n3895), .Y(\D_cache/n690 ) );
  OAI2BB2XL U9695 ( .B0(\D_cache/n235 ), .B1(n3915), .A0N(
        \D_cache/cache[1][138] ), .A1N(n3916), .Y(\D_cache/n691 ) );
  OAI2BB2XL U9696 ( .B0(\D_cache/n235 ), .B1(n3936), .A0N(
        \D_cache/cache[0][138] ), .A1N(n3937), .Y(\D_cache/n692 ) );
  OAI2BB2XL U9697 ( .B0(\D_cache/n241 ), .B1(n3791), .A0N(
        \D_cache/cache[7][132] ), .A1N(n3797), .Y(\D_cache/n733 ) );
  OAI2BB2XL U9698 ( .B0(\D_cache/n241 ), .B1(n3811), .A0N(
        \D_cache/cache[6][132] ), .A1N(n3817), .Y(\D_cache/n734 ) );
  OAI2BB2XL U9699 ( .B0(\D_cache/n241 ), .B1(n3829), .A0N(
        \D_cache/cache[5][132] ), .A1N(n3835), .Y(\D_cache/n735 ) );
  OAI2BB2XL U9700 ( .B0(\D_cache/n241 ), .B1(n3849), .A0N(
        \D_cache/cache[4][132] ), .A1N(n3857), .Y(\D_cache/n736 ) );
  OAI2BB2XL U9701 ( .B0(\D_cache/n241 ), .B1(n3868), .A0N(
        \D_cache/cache[3][132] ), .A1N(n3876), .Y(\D_cache/n737 ) );
  OAI2BB2XL U9702 ( .B0(\D_cache/n241 ), .B1(n3891), .A0N(
        \D_cache/cache[2][132] ), .A1N(n3897), .Y(\D_cache/n738 ) );
  OAI2BB2XL U9703 ( .B0(\D_cache/n241 ), .B1(n3911), .A0N(
        \D_cache/cache[1][132] ), .A1N(n3918), .Y(\D_cache/n739 ) );
  OAI2BB2XL U9704 ( .B0(\D_cache/n241 ), .B1(n3931), .A0N(
        \D_cache/cache[0][132] ), .A1N(n3939), .Y(\D_cache/n740 ) );
  OAI2BB2XL U9705 ( .B0(\D_cache/n243 ), .B1(n3790), .A0N(
        \D_cache/cache[7][130] ), .A1N(n3796), .Y(\D_cache/n749 ) );
  OAI2BB2XL U9706 ( .B0(\D_cache/n243 ), .B1(n3810), .A0N(
        \D_cache/cache[6][130] ), .A1N(n3816), .Y(\D_cache/n750 ) );
  OAI2BB2XL U9707 ( .B0(\D_cache/n243 ), .B1(n3831), .A0N(
        \D_cache/cache[5][130] ), .A1N(n3834), .Y(\D_cache/n751 ) );
  OAI2BB2XL U9708 ( .B0(\D_cache/n243 ), .B1(n3848), .A0N(
        \D_cache/cache[4][130] ), .A1N(n3856), .Y(\D_cache/n752 ) );
  OAI2BB2XL U9709 ( .B0(\D_cache/n243 ), .B1(n3867), .A0N(
        \D_cache/cache[3][130] ), .A1N(n3875), .Y(\D_cache/n753 ) );
  OAI2BB2XL U9710 ( .B0(\D_cache/n243 ), .B1(n3890), .A0N(
        \D_cache/cache[2][130] ), .A1N(n3896), .Y(\D_cache/n754 ) );
  OAI2BB2XL U9711 ( .B0(\D_cache/n243 ), .B1(n3910), .A0N(
        \D_cache/cache[1][130] ), .A1N(n3917), .Y(\D_cache/n755 ) );
  OAI2BB2XL U9712 ( .B0(\D_cache/n243 ), .B1(n3930), .A0N(
        \D_cache/cache[0][130] ), .A1N(n3938), .Y(\D_cache/n756 ) );
  OAI2BB2XL U9713 ( .B0(\D_cache/n244 ), .B1(n3790), .A0N(
        \D_cache/cache[7][129] ), .A1N(n3796), .Y(\D_cache/n757 ) );
  OAI2BB2XL U9714 ( .B0(\D_cache/n244 ), .B1(n3810), .A0N(
        \D_cache/cache[6][129] ), .A1N(n3816), .Y(\D_cache/n758 ) );
  OAI2BB2XL U9715 ( .B0(\D_cache/n244 ), .B1(n3825), .A0N(
        \D_cache/cache[5][129] ), .A1N(n3834), .Y(\D_cache/n759 ) );
  OAI2BB2XL U9716 ( .B0(\D_cache/n244 ), .B1(n3848), .A0N(
        \D_cache/cache[4][129] ), .A1N(n3856), .Y(\D_cache/n760 ) );
  OAI2BB2XL U9717 ( .B0(\D_cache/n244 ), .B1(n3867), .A0N(
        \D_cache/cache[3][129] ), .A1N(n3875), .Y(\D_cache/n761 ) );
  OAI2BB2XL U9718 ( .B0(\D_cache/n244 ), .B1(n3890), .A0N(
        \D_cache/cache[2][129] ), .A1N(n3896), .Y(\D_cache/n762 ) );
  OAI2BB2XL U9719 ( .B0(\D_cache/n244 ), .B1(n3910), .A0N(
        \D_cache/cache[1][129] ), .A1N(n3917), .Y(\D_cache/n763 ) );
  OAI2BB2XL U9720 ( .B0(\D_cache/n244 ), .B1(n3930), .A0N(
        \D_cache/cache[0][129] ), .A1N(n3938), .Y(\D_cache/n764 ) );
  OAI2BB2XL U9721 ( .B0(\D_cache/n237 ), .B1(n3794), .A0N(
        \D_cache/cache[7][136] ), .A1N(n3796), .Y(\D_cache/n701 ) );
  OAI2BB2XL U9722 ( .B0(\D_cache/n237 ), .B1(n3814), .A0N(
        \D_cache/cache[6][136] ), .A1N(n3816), .Y(\D_cache/n702 ) );
  OAI2BB2XL U9723 ( .B0(\D_cache/n237 ), .B1(n3832), .A0N(
        \D_cache/cache[5][136] ), .A1N(n3834), .Y(\D_cache/n703 ) );
  OAI2BB2XL U9724 ( .B0(\D_cache/n237 ), .B1(n3854), .A0N(
        \D_cache/cache[4][136] ), .A1N(n3856), .Y(\D_cache/n704 ) );
  OAI2BB2XL U9725 ( .B0(\D_cache/n237 ), .B1(n3873), .A0N(
        \D_cache/cache[3][136] ), .A1N(n3875), .Y(\D_cache/n705 ) );
  OAI2BB2XL U9726 ( .B0(\D_cache/n237 ), .B1(n3894), .A0N(
        \D_cache/cache[2][136] ), .A1N(n3896), .Y(\D_cache/n706 ) );
  OAI2BB2XL U9727 ( .B0(\D_cache/n237 ), .B1(n3915), .A0N(
        \D_cache/cache[1][136] ), .A1N(n3917), .Y(\D_cache/n707 ) );
  OAI2BB2XL U9728 ( .B0(\D_cache/n237 ), .B1(n3936), .A0N(
        \D_cache/cache[0][136] ), .A1N(n3938), .Y(\D_cache/n708 ) );
  OAI2BB2XL U9729 ( .B0(\D_cache/n245 ), .B1(n3790), .A0N(
        \D_cache/cache[7][128] ), .A1N(n3796), .Y(\D_cache/n765 ) );
  OAI2BB2XL U9730 ( .B0(\D_cache/n234 ), .B1(n3793), .A0N(
        \D_cache/cache[7][139] ), .A1N(n3795), .Y(\D_cache/n677 ) );
  OAI2BB2XL U9731 ( .B0(\D_cache/n234 ), .B1(n3813), .A0N(
        \D_cache/cache[6][139] ), .A1N(n3815), .Y(\D_cache/n678 ) );
  OAI2BB2XL U9732 ( .B0(\D_cache/n234 ), .B1(n3831), .A0N(
        \D_cache/cache[5][139] ), .A1N(n3833), .Y(\D_cache/n679 ) );
  OAI2BB2XL U9733 ( .B0(\D_cache/n234 ), .B1(n3853), .A0N(
        \D_cache/cache[4][139] ), .A1N(n3855), .Y(\D_cache/n680 ) );
  OAI2BB2XL U9734 ( .B0(\D_cache/n234 ), .B1(n3872), .A0N(
        \D_cache/cache[3][139] ), .A1N(n3874), .Y(\D_cache/n681 ) );
  OAI2BB2XL U9735 ( .B0(\D_cache/n234 ), .B1(n3893), .A0N(
        \D_cache/cache[2][139] ), .A1N(n3895), .Y(\D_cache/n682 ) );
  OAI2BB2XL U9736 ( .B0(\D_cache/n234 ), .B1(n3914), .A0N(
        \D_cache/cache[1][139] ), .A1N(n3916), .Y(\D_cache/n683 ) );
  OAI2BB2XL U9737 ( .B0(\D_cache/n234 ), .B1(n3935), .A0N(
        \D_cache/cache[0][139] ), .A1N(n3937), .Y(\D_cache/n684 ) );
  OAI2BB2XL U9738 ( .B0(\D_cache/n245 ), .B1(n3810), .A0N(
        \D_cache/cache[6][128] ), .A1N(n3816), .Y(\D_cache/n766 ) );
  OAI2BB2XL U9739 ( .B0(\D_cache/n245 ), .B1(n3826), .A0N(
        \D_cache/cache[5][128] ), .A1N(n3834), .Y(\D_cache/n767 ) );
  OAI2BB2XL U9740 ( .B0(\D_cache/n245 ), .B1(n3848), .A0N(
        \D_cache/cache[4][128] ), .A1N(n3856), .Y(\D_cache/n768 ) );
  OAI2BB2XL U9741 ( .B0(\D_cache/n245 ), .B1(n3867), .A0N(
        \D_cache/cache[3][128] ), .A1N(n3875), .Y(\D_cache/n769 ) );
  OAI2BB2XL U9742 ( .B0(\D_cache/n245 ), .B1(n3890), .A0N(
        \D_cache/cache[2][128] ), .A1N(n3896), .Y(\D_cache/n770 ) );
  OAI2BB2XL U9743 ( .B0(\D_cache/n245 ), .B1(n3910), .A0N(
        \D_cache/cache[1][128] ), .A1N(n3917), .Y(\D_cache/n771 ) );
  OAI2BB2XL U9744 ( .B0(\D_cache/n245 ), .B1(n3930), .A0N(
        \D_cache/cache[0][128] ), .A1N(n3938), .Y(\D_cache/n772 ) );
  OAI2BB2XL U9745 ( .B0(\D_cache/n222 ), .B1(n3785), .A0N(
        \D_cache/cache[7][151] ), .A1N(n3796), .Y(\D_cache/n581 ) );
  OAI2BB2XL U9746 ( .B0(\D_cache/n222 ), .B1(n3805), .A0N(
        \D_cache/cache[6][151] ), .A1N(n3816), .Y(\D_cache/n582 ) );
  OAI2BB2XL U9747 ( .B0(\D_cache/n222 ), .B1(n3831), .A0N(
        \D_cache/cache[5][151] ), .A1N(n3834), .Y(\D_cache/n583 ) );
  OAI2BB2XL U9748 ( .B0(\D_cache/n222 ), .B1(n3850), .A0N(
        \D_cache/cache[4][151] ), .A1N(n3856), .Y(\D_cache/n584 ) );
  OAI2BB2XL U9749 ( .B0(\D_cache/n222 ), .B1(n3869), .A0N(
        \D_cache/cache[3][151] ), .A1N(n3875), .Y(\D_cache/n585 ) );
  OAI2BB2XL U9750 ( .B0(\D_cache/n222 ), .B1(n3885), .A0N(
        \D_cache/cache[2][151] ), .A1N(n3896), .Y(\D_cache/n586 ) );
  OAI2BB2XL U9751 ( .B0(\D_cache/n222 ), .B1(n3912), .A0N(
        \D_cache/cache[1][151] ), .A1N(n3917), .Y(\D_cache/n587 ) );
  OAI2BB2XL U9752 ( .B0(\D_cache/n222 ), .B1(n3932), .A0N(
        \D_cache/cache[0][151] ), .A1N(n3938), .Y(\D_cache/n588 ) );
  OAI2BB2XL U9753 ( .B0(\D_cache/n223 ), .B1(n3791), .A0N(
        \D_cache/cache[7][150] ), .A1N(n3796), .Y(\D_cache/n589 ) );
  OAI2BB2XL U9754 ( .B0(\D_cache/n223 ), .B1(n3811), .A0N(
        \D_cache/cache[6][150] ), .A1N(n3816), .Y(\D_cache/n590 ) );
  OAI2BB2XL U9755 ( .B0(\D_cache/n223 ), .B1(n3826), .A0N(
        \D_cache/cache[5][150] ), .A1N(n3834), .Y(\D_cache/n591 ) );
  OAI2BB2XL U9756 ( .B0(\D_cache/n223 ), .B1(n3850), .A0N(
        \D_cache/cache[4][150] ), .A1N(n3856), .Y(\D_cache/n592 ) );
  OAI2BB2XL U9757 ( .B0(\D_cache/n223 ), .B1(n3869), .A0N(
        \D_cache/cache[3][150] ), .A1N(n3875), .Y(\D_cache/n593 ) );
  OAI2BB2XL U9758 ( .B0(\D_cache/n223 ), .B1(n3891), .A0N(
        \D_cache/cache[2][150] ), .A1N(n3896), .Y(\D_cache/n594 ) );
  OAI2BB2XL U9759 ( .B0(\D_cache/n223 ), .B1(n3912), .A0N(
        \D_cache/cache[1][150] ), .A1N(n3917), .Y(\D_cache/n595 ) );
  OAI2BB2XL U9760 ( .B0(\D_cache/n223 ), .B1(n3932), .A0N(
        \D_cache/cache[0][150] ), .A1N(n3938), .Y(\D_cache/n596 ) );
  OAI2BB2XL U9761 ( .B0(\D_cache/n224 ), .B1(n3786), .A0N(
        \D_cache/cache[7][149] ), .A1N(n3796), .Y(\D_cache/n597 ) );
  OAI2BB2XL U9762 ( .B0(\D_cache/n224 ), .B1(n3806), .A0N(
        \D_cache/cache[6][149] ), .A1N(n3816), .Y(\D_cache/n598 ) );
  OAI2BB2XL U9763 ( .B0(\D_cache/n224 ), .B1(n3830), .A0N(
        \D_cache/cache[5][149] ), .A1N(n3834), .Y(\D_cache/n599 ) );
  OAI2BB2XL U9764 ( .B0(\D_cache/n224 ), .B1(n3850), .A0N(
        \D_cache/cache[4][149] ), .A1N(n3856), .Y(\D_cache/n600 ) );
  OAI2BB2XL U9765 ( .B0(\D_cache/n224 ), .B1(n3869), .A0N(
        \D_cache/cache[3][149] ), .A1N(n3875), .Y(\D_cache/n601 ) );
  OAI2BB2XL U9766 ( .B0(\D_cache/n224 ), .B1(n3886), .A0N(
        \D_cache/cache[2][149] ), .A1N(n3896), .Y(\D_cache/n602 ) );
  OAI2BB2XL U9767 ( .B0(\D_cache/n224 ), .B1(n3912), .A0N(
        \D_cache/cache[1][149] ), .A1N(n3917), .Y(\D_cache/n603 ) );
  OAI2BB2XL U9768 ( .B0(\D_cache/n224 ), .B1(n3932), .A0N(
        \D_cache/cache[0][149] ), .A1N(n3938), .Y(\D_cache/n604 ) );
  OAI2BB2XL U9769 ( .B0(\D_cache/n225 ), .B1(n3785), .A0N(
        \D_cache/cache[7][148] ), .A1N(n3796), .Y(\D_cache/n605 ) );
  OAI2BB2XL U9770 ( .B0(\D_cache/n225 ), .B1(n3805), .A0N(
        \D_cache/cache[6][148] ), .A1N(n3816), .Y(\D_cache/n606 ) );
  OAI2BB2XL U9771 ( .B0(\D_cache/n225 ), .B1(n3824), .A0N(
        \D_cache/cache[5][148] ), .A1N(n3834), .Y(\D_cache/n607 ) );
  OAI2BB2XL U9772 ( .B0(\D_cache/n225 ), .B1(n3850), .A0N(
        \D_cache/cache[4][148] ), .A1N(n3856), .Y(\D_cache/n608 ) );
  OAI2BB2XL U9773 ( .B0(\D_cache/n225 ), .B1(n3869), .A0N(
        \D_cache/cache[3][148] ), .A1N(n3875), .Y(\D_cache/n609 ) );
  OAI2BB2XL U9774 ( .B0(\D_cache/n225 ), .B1(n3885), .A0N(
        \D_cache/cache[2][148] ), .A1N(n3896), .Y(\D_cache/n610 ) );
  OAI2BB2XL U9775 ( .B0(\D_cache/n225 ), .B1(n3912), .A0N(
        \D_cache/cache[1][148] ), .A1N(n3917), .Y(\D_cache/n611 ) );
  OAI2BB2XL U9776 ( .B0(\D_cache/n225 ), .B1(n3932), .A0N(
        \D_cache/cache[0][148] ), .A1N(n3938), .Y(\D_cache/n612 ) );
  OAI2BB2XL U9777 ( .B0(\D_cache/n226 ), .B1(n3785), .A0N(
        \D_cache/cache[7][147] ), .A1N(n3795), .Y(\D_cache/n613 ) );
  OAI2BB2XL U9778 ( .B0(\D_cache/n226 ), .B1(n3805), .A0N(
        \D_cache/cache[6][147] ), .A1N(n3815), .Y(\D_cache/n614 ) );
  OAI2BB2XL U9779 ( .B0(\D_cache/n226 ), .B1(n3830), .A0N(
        \D_cache/cache[5][147] ), .A1N(n3833), .Y(\D_cache/n615 ) );
  OAI2BB2XL U9780 ( .B0(\D_cache/n226 ), .B1(n3851), .A0N(
        \D_cache/cache[4][147] ), .A1N(n3855), .Y(\D_cache/n616 ) );
  OAI2BB2XL U9781 ( .B0(\D_cache/n226 ), .B1(n3870), .A0N(
        \D_cache/cache[3][147] ), .A1N(n3874), .Y(\D_cache/n617 ) );
  OAI2BB2XL U9782 ( .B0(\D_cache/n226 ), .B1(n3885), .A0N(
        \D_cache/cache[2][147] ), .A1N(n3895), .Y(\D_cache/n618 ) );
  OAI2BB2XL U9783 ( .B0(\D_cache/n226 ), .B1(n3905), .A0N(
        \D_cache/cache[1][147] ), .A1N(n3916), .Y(\D_cache/n619 ) );
  OAI2BB2XL U9784 ( .B0(\D_cache/n226 ), .B1(n3933), .A0N(
        \D_cache/cache[0][147] ), .A1N(n3937), .Y(\D_cache/n620 ) );
  OAI2BB2XL U9785 ( .B0(\D_cache/n227 ), .B1(n3791), .A0N(
        \D_cache/cache[7][146] ), .A1N(n3795), .Y(\D_cache/n621 ) );
  OAI2BB2XL U9786 ( .B0(\D_cache/n227 ), .B1(n3811), .A0N(
        \D_cache/cache[6][146] ), .A1N(n3815), .Y(\D_cache/n622 ) );
  OAI2BB2XL U9787 ( .B0(\D_cache/n227 ), .B1(n3830), .A0N(
        \D_cache/cache[5][146] ), .A1N(n3833), .Y(\D_cache/n623 ) );
  OAI2BB2XL U9788 ( .B0(\D_cache/n227 ), .B1(n3851), .A0N(
        \D_cache/cache[4][146] ), .A1N(n3855), .Y(\D_cache/n624 ) );
  OAI2BB2XL U9789 ( .B0(\D_cache/n227 ), .B1(n3870), .A0N(
        \D_cache/cache[3][146] ), .A1N(n3874), .Y(\D_cache/n625 ) );
  OAI2BB2XL U9790 ( .B0(\D_cache/n227 ), .B1(n3891), .A0N(
        \D_cache/cache[2][146] ), .A1N(n3895), .Y(\D_cache/n626 ) );
  OAI2BB2XL U9791 ( .B0(\D_cache/n227 ), .B1(n3911), .A0N(
        \D_cache/cache[1][146] ), .A1N(n3916), .Y(\D_cache/n627 ) );
  OAI2BB2XL U9792 ( .B0(\D_cache/n227 ), .B1(n3933), .A0N(
        \D_cache/cache[0][146] ), .A1N(n3937), .Y(\D_cache/n628 ) );
  OAI2BB2XL U9793 ( .B0(\D_cache/n228 ), .B1(n3786), .A0N(
        \D_cache/cache[7][145] ), .A1N(n3795), .Y(\D_cache/n629 ) );
  OAI2BB2XL U9794 ( .B0(\D_cache/n228 ), .B1(n3806), .A0N(
        \D_cache/cache[6][145] ), .A1N(n3815), .Y(\D_cache/n630 ) );
  OAI2BB2XL U9795 ( .B0(\D_cache/n228 ), .B1(n3830), .A0N(
        \D_cache/cache[5][145] ), .A1N(n3833), .Y(\D_cache/n631 ) );
  OAI2BB2XL U9796 ( .B0(\D_cache/n228 ), .B1(n3851), .A0N(
        \D_cache/cache[4][145] ), .A1N(n3855), .Y(\D_cache/n632 ) );
  OAI2BB2XL U9797 ( .B0(\D_cache/n228 ), .B1(n3870), .A0N(
        \D_cache/cache[3][145] ), .A1N(n3874), .Y(\D_cache/n633 ) );
  OAI2BB2XL U9798 ( .B0(\D_cache/n228 ), .B1(n3886), .A0N(
        \D_cache/cache[2][145] ), .A1N(n3895), .Y(\D_cache/n634 ) );
  OAI2BB2XL U9799 ( .B0(\D_cache/n228 ), .B1(n3906), .A0N(
        \D_cache/cache[1][145] ), .A1N(n3916), .Y(\D_cache/n635 ) );
  OAI2BB2XL U9800 ( .B0(\D_cache/n228 ), .B1(n3933), .A0N(
        \D_cache/cache[0][145] ), .A1N(n3937), .Y(\D_cache/n636 ) );
  OAI2BB2XL U9801 ( .B0(\D_cache/n229 ), .B1(n3785), .A0N(
        \D_cache/cache[7][144] ), .A1N(n3795), .Y(\D_cache/n637 ) );
  OAI2BB2XL U9802 ( .B0(\D_cache/n229 ), .B1(n3805), .A0N(
        \D_cache/cache[6][144] ), .A1N(n3815), .Y(\D_cache/n638 ) );
  OAI2BB2XL U9803 ( .B0(\D_cache/n229 ), .B1(n3830), .A0N(
        \D_cache/cache[5][144] ), .A1N(n3833), .Y(\D_cache/n639 ) );
  OAI2BB2XL U9804 ( .B0(\D_cache/n229 ), .B1(n3851), .A0N(
        \D_cache/cache[4][144] ), .A1N(n3855), .Y(\D_cache/n640 ) );
  OAI2BB2XL U9805 ( .B0(\D_cache/n229 ), .B1(n3870), .A0N(
        \D_cache/cache[3][144] ), .A1N(n3874), .Y(\D_cache/n641 ) );
  OAI2BB2XL U9806 ( .B0(\D_cache/n229 ), .B1(n3885), .A0N(
        \D_cache/cache[2][144] ), .A1N(n3895), .Y(\D_cache/n642 ) );
  OAI2BB2XL U9807 ( .B0(\D_cache/n229 ), .B1(n3905), .A0N(
        \D_cache/cache[1][144] ), .A1N(n3916), .Y(\D_cache/n643 ) );
  OAI2BB2XL U9808 ( .B0(\D_cache/n229 ), .B1(n3933), .A0N(
        \D_cache/cache[0][144] ), .A1N(n3937), .Y(\D_cache/n644 ) );
  OAI2BB2XL U9809 ( .B0(\D_cache/n230 ), .B1(n3792), .A0N(
        \D_cache/cache[7][143] ), .A1N(n3795), .Y(\D_cache/n645 ) );
  OAI2BB2XL U9810 ( .B0(\D_cache/n230 ), .B1(n3812), .A0N(
        \D_cache/cache[6][143] ), .A1N(n3815), .Y(\D_cache/n646 ) );
  OAI2BB2XL U9811 ( .B0(\D_cache/n230 ), .B1(n3829), .A0N(
        \D_cache/cache[5][143] ), .A1N(n3833), .Y(\D_cache/n647 ) );
  OAI2BB2XL U9812 ( .B0(\D_cache/n230 ), .B1(n3852), .A0N(
        \D_cache/cache[4][143] ), .A1N(n3855), .Y(\D_cache/n648 ) );
  OAI2BB2XL U9813 ( .B0(\D_cache/n230 ), .B1(n3871), .A0N(
        \D_cache/cache[3][143] ), .A1N(n3874), .Y(\D_cache/n649 ) );
  OAI2BB2XL U9814 ( .B0(\D_cache/n230 ), .B1(n3892), .A0N(
        \D_cache/cache[2][143] ), .A1N(n3895), .Y(\D_cache/n650 ) );
  OAI2BB2XL U9815 ( .B0(\D_cache/n230 ), .B1(n3913), .A0N(
        \D_cache/cache[1][143] ), .A1N(n3916), .Y(\D_cache/n651 ) );
  OAI2BB2XL U9816 ( .B0(\D_cache/n230 ), .B1(n3934), .A0N(
        \D_cache/cache[0][143] ), .A1N(n3937), .Y(\D_cache/n652 ) );
  OAI2BB2XL U9817 ( .B0(\D_cache/n231 ), .B1(n3792), .A0N(
        \D_cache/cache[7][142] ), .A1N(n3795), .Y(\D_cache/n653 ) );
  OAI2BB2XL U9818 ( .B0(\D_cache/n231 ), .B1(n3812), .A0N(
        \D_cache/cache[6][142] ), .A1N(n3815), .Y(\D_cache/n654 ) );
  OAI2BB2XL U9819 ( .B0(\D_cache/n231 ), .B1(n3828), .A0N(
        \D_cache/cache[5][142] ), .A1N(n3833), .Y(\D_cache/n655 ) );
  OAI2BB2XL U9820 ( .B0(\D_cache/n231 ), .B1(n3852), .A0N(
        \D_cache/cache[4][142] ), .A1N(n3855), .Y(\D_cache/n656 ) );
  OAI2BB2XL U9821 ( .B0(\D_cache/n231 ), .B1(n3871), .A0N(
        \D_cache/cache[3][142] ), .A1N(n3874), .Y(\D_cache/n657 ) );
  OAI2BB2XL U9822 ( .B0(\D_cache/n231 ), .B1(n3892), .A0N(
        \D_cache/cache[2][142] ), .A1N(n3895), .Y(\D_cache/n658 ) );
  OAI2BB2XL U9823 ( .B0(\D_cache/n231 ), .B1(n3913), .A0N(
        \D_cache/cache[1][142] ), .A1N(n3916), .Y(\D_cache/n659 ) );
  OAI2BB2XL U9824 ( .B0(\D_cache/n231 ), .B1(n3934), .A0N(
        \D_cache/cache[0][142] ), .A1N(n3937), .Y(\D_cache/n660 ) );
  OAI2BB2XL U9825 ( .B0(\D_cache/n232 ), .B1(n3792), .A0N(
        \D_cache/cache[7][141] ), .A1N(n3794), .Y(\D_cache/n661 ) );
  OAI2BB2XL U9826 ( .B0(\D_cache/n232 ), .B1(n3812), .A0N(
        \D_cache/cache[6][141] ), .A1N(n3814), .Y(\D_cache/n662 ) );
  OAI2BB2XL U9827 ( .B0(\D_cache/n232 ), .B1(n3827), .A0N(
        \D_cache/cache[5][141] ), .A1N(n3832), .Y(\D_cache/n663 ) );
  OAI2BB2XL U9828 ( .B0(\D_cache/n232 ), .B1(n3852), .A0N(
        \D_cache/cache[4][141] ), .A1N(n3854), .Y(\D_cache/n664 ) );
  OAI2BB2XL U9829 ( .B0(\D_cache/n232 ), .B1(n3871), .A0N(
        \D_cache/cache[3][141] ), .A1N(n3873), .Y(\D_cache/n665 ) );
  OAI2BB2XL U9830 ( .B0(\D_cache/n232 ), .B1(n3892), .A0N(
        \D_cache/cache[2][141] ), .A1N(n3894), .Y(\D_cache/n666 ) );
  OAI2BB2XL U9831 ( .B0(\D_cache/n232 ), .B1(n3913), .A0N(
        \D_cache/cache[1][141] ), .A1N(n3915), .Y(\D_cache/n667 ) );
  OAI2BB2XL U9832 ( .B0(\D_cache/n232 ), .B1(n3934), .A0N(
        \D_cache/cache[0][141] ), .A1N(n3936), .Y(\D_cache/n668 ) );
  OAI2BB2XL U9833 ( .B0(\D_cache/n233 ), .B1(n3793), .A0N(
        \D_cache/cache[7][140] ), .A1N(n3795), .Y(\D_cache/n669 ) );
  OAI2BB2XL U9834 ( .B0(\D_cache/n233 ), .B1(n3813), .A0N(
        \D_cache/cache[6][140] ), .A1N(n3815), .Y(\D_cache/n670 ) );
  OAI2BB2XL U9835 ( .B0(\D_cache/n233 ), .B1(n3831), .A0N(
        \D_cache/cache[5][140] ), .A1N(n3833), .Y(\D_cache/n671 ) );
  OAI2BB2XL U9836 ( .B0(\D_cache/n233 ), .B1(n3853), .A0N(
        \D_cache/cache[4][140] ), .A1N(n3855), .Y(\D_cache/n672 ) );
  OAI2BB2XL U9837 ( .B0(\D_cache/n233 ), .B1(n3872), .A0N(
        \D_cache/cache[3][140] ), .A1N(n3874), .Y(\D_cache/n673 ) );
  OAI2BB2XL U9838 ( .B0(\D_cache/n233 ), .B1(n3893), .A0N(
        \D_cache/cache[2][140] ), .A1N(n3895), .Y(\D_cache/n674 ) );
  OAI2BB2XL U9839 ( .B0(\D_cache/n233 ), .B1(n3914), .A0N(
        \D_cache/cache[1][140] ), .A1N(n3916), .Y(\D_cache/n675 ) );
  OAI2BB2XL U9840 ( .B0(\D_cache/n233 ), .B1(n3935), .A0N(
        \D_cache/cache[0][140] ), .A1N(n3937), .Y(\D_cache/n676 ) );
  OAI2BB2XL U9841 ( .B0(\D_cache/n236 ), .B1(n3793), .A0N(
        \D_cache/cache[7][137] ), .A1N(n3795), .Y(\D_cache/n693 ) );
  OAI2BB2XL U9842 ( .B0(\D_cache/n236 ), .B1(n3813), .A0N(
        \D_cache/cache[6][137] ), .A1N(n3815), .Y(\D_cache/n694 ) );
  OAI2BB2XL U9843 ( .B0(\D_cache/n236 ), .B1(n3831), .A0N(
        \D_cache/cache[5][137] ), .A1N(n3833), .Y(\D_cache/n695 ) );
  OAI2BB2XL U9844 ( .B0(\D_cache/n236 ), .B1(n3853), .A0N(
        \D_cache/cache[4][137] ), .A1N(n3855), .Y(\D_cache/n696 ) );
  OAI2BB2XL U9845 ( .B0(\D_cache/n236 ), .B1(n3872), .A0N(
        \D_cache/cache[3][137] ), .A1N(n3874), .Y(\D_cache/n697 ) );
  OAI2BB2XL U9846 ( .B0(\D_cache/n236 ), .B1(n3893), .A0N(
        \D_cache/cache[2][137] ), .A1N(n3895), .Y(\D_cache/n698 ) );
  OAI2BB2XL U9847 ( .B0(\D_cache/n236 ), .B1(n3914), .A0N(
        \D_cache/cache[1][137] ), .A1N(n3916), .Y(\D_cache/n699 ) );
  OAI2BB2XL U9848 ( .B0(\D_cache/n236 ), .B1(n3935), .A0N(
        \D_cache/cache[0][137] ), .A1N(n3937), .Y(\D_cache/n700 ) );
  OAI2BB2XL U9849 ( .B0(\D_cache/n238 ), .B1(n3793), .A0N(
        \D_cache/cache[7][135] ), .A1N(n3796), .Y(\D_cache/n709 ) );
  OAI2BB2XL U9850 ( .B0(\D_cache/n238 ), .B1(n3813), .A0N(
        \D_cache/cache[6][135] ), .A1N(n3816), .Y(\D_cache/n710 ) );
  OAI2BB2XL U9851 ( .B0(\D_cache/n238 ), .B1(n3831), .A0N(
        \D_cache/cache[5][135] ), .A1N(n3834), .Y(\D_cache/n711 ) );
  OAI2BB2XL U9852 ( .B0(\D_cache/n238 ), .B1(n3853), .A0N(
        \D_cache/cache[4][135] ), .A1N(n3856), .Y(\D_cache/n712 ) );
  OAI2BB2XL U9853 ( .B0(\D_cache/n238 ), .B1(n3872), .A0N(
        \D_cache/cache[3][135] ), .A1N(n3875), .Y(\D_cache/n713 ) );
  OAI2BB2XL U9854 ( .B0(\D_cache/n238 ), .B1(n3893), .A0N(
        \D_cache/cache[2][135] ), .A1N(n3896), .Y(\D_cache/n714 ) );
  OAI2BB2XL U9855 ( .B0(\D_cache/n238 ), .B1(n3914), .A0N(
        \D_cache/cache[1][135] ), .A1N(n3917), .Y(\D_cache/n715 ) );
  OAI2BB2XL U9856 ( .B0(\D_cache/n238 ), .B1(n3935), .A0N(
        \D_cache/cache[0][135] ), .A1N(n3938), .Y(\D_cache/n716 ) );
  OAI2BB2XL U9857 ( .B0(\D_cache/n242 ), .B1(n3791), .A0N(
        \D_cache/cache[7][131] ), .A1N(n3797), .Y(\D_cache/n741 ) );
  OAI2BB2XL U9858 ( .B0(\D_cache/n242 ), .B1(n3811), .A0N(
        \D_cache/cache[6][131] ), .A1N(n3817), .Y(\D_cache/n742 ) );
  OAI2BB2XL U9859 ( .B0(\D_cache/n242 ), .B1(n3829), .A0N(
        \D_cache/cache[5][131] ), .A1N(n3835), .Y(\D_cache/n743 ) );
  OAI2BB2XL U9860 ( .B0(\D_cache/n242 ), .B1(n3849), .A0N(
        \D_cache/cache[4][131] ), .A1N(n3857), .Y(\D_cache/n744 ) );
  OAI2BB2XL U9861 ( .B0(\D_cache/n242 ), .B1(n3868), .A0N(
        \D_cache/cache[3][131] ), .A1N(n3876), .Y(\D_cache/n745 ) );
  OAI2BB2XL U9862 ( .B0(\D_cache/n242 ), .B1(n3891), .A0N(
        \D_cache/cache[2][131] ), .A1N(n3897), .Y(\D_cache/n746 ) );
  OAI2BB2XL U9863 ( .B0(\D_cache/n242 ), .B1(n3911), .A0N(
        \D_cache/cache[1][131] ), .A1N(n3918), .Y(\D_cache/n747 ) );
  OAI2BB2XL U9864 ( .B0(\D_cache/n242 ), .B1(n3931), .A0N(
        \D_cache/cache[0][131] ), .A1N(n3939), .Y(\D_cache/n748 ) );
  NOR2X1 U9865 ( .A(n8809), .B(mem_ready_D), .Y(\D_cache/n218 ) );
  OAI2BB2XL U9866 ( .B0(\D_cache/n215 ), .B1(n3791), .A0N(
        \D_cache/cache[7][153] ), .A1N(n3797), .Y(\D_cache/n565 ) );
  OAI2BB2XL U9867 ( .B0(\D_cache/n215 ), .B1(n3811), .A0N(
        \D_cache/cache[6][153] ), .A1N(n3817), .Y(\D_cache/n566 ) );
  OAI2BB2XL U9868 ( .B0(\D_cache/n215 ), .B1(n3829), .A0N(
        \D_cache/cache[5][153] ), .A1N(n3835), .Y(\D_cache/n567 ) );
  OAI2BB2XL U9869 ( .B0(\D_cache/n215 ), .B1(n3849), .A0N(
        \D_cache/cache[4][153] ), .A1N(n3857), .Y(\D_cache/n568 ) );
  OAI2BB2XL U9870 ( .B0(\D_cache/n215 ), .B1(n3868), .A0N(
        \D_cache/cache[3][153] ), .A1N(n3876), .Y(\D_cache/n569 ) );
  OAI2BB2XL U9871 ( .B0(\D_cache/n215 ), .B1(n3891), .A0N(
        \D_cache/cache[2][153] ), .A1N(n3897), .Y(\D_cache/n570 ) );
  OAI2BB2XL U9872 ( .B0(\D_cache/n215 ), .B1(n3911), .A0N(
        \D_cache/cache[1][153] ), .A1N(n3918), .Y(\D_cache/n571 ) );
  OAI2BB2XL U9873 ( .B0(\D_cache/n215 ), .B1(n3931), .A0N(
        \D_cache/cache[0][153] ), .A1N(n3939), .Y(\D_cache/n572 ) );
  MXI2X1 U9874 ( .A(\i_MIPS/n373 ), .B(\i_MIPS/n372 ), .S0(n3617), .Y(
        \i_MIPS/n563 ) );
  MXI2X1 U9875 ( .A(\i_MIPS/n338 ), .B(\i_MIPS/n339 ), .S0(n3621), .Y(
        \i_MIPS/n529 ) );
  MXI2X1 U9876 ( .A(\i_MIPS/n334 ), .B(\i_MIPS/n335 ), .S0(n3621), .Y(
        \i_MIPS/n524 ) );
  MXI2X1 U9877 ( .A(\i_MIPS/n333 ), .B(\i_MIPS/n332 ), .S0(n3621), .Y(
        \i_MIPS/n523 ) );
  MXI2X1 U9878 ( .A(\i_MIPS/n331 ), .B(\i_MIPS/n330 ), .S0(n3621), .Y(
        \i_MIPS/n522 ) );
  MXI2X1 U9879 ( .A(\i_MIPS/n321 ), .B(\i_MIPS/n320 ), .S0(n3618), .Y(
        \i_MIPS/n517 ) );
  MXI2X1 U9880 ( .A(\i_MIPS/n319 ), .B(\i_MIPS/n318 ), .S0(n3618), .Y(
        \i_MIPS/n516 ) );
  MXI2X1 U9881 ( .A(\i_MIPS/n317 ), .B(\i_MIPS/n316 ), .S0(n3618), .Y(
        \i_MIPS/n515 ) );
  MXI2X1 U9882 ( .A(\i_MIPS/n315 ), .B(\i_MIPS/n314 ), .S0(n3620), .Y(
        \i_MIPS/n514 ) );
  MXI2X1 U9883 ( .A(\i_MIPS/n313 ), .B(\i_MIPS/n312 ), .S0(n3617), .Y(
        \i_MIPS/n513 ) );
  MXI2X1 U9884 ( .A(\i_MIPS/n310 ), .B(\i_MIPS/n311 ), .S0(n3617), .Y(
        \i_MIPS/n479 ) );
  MXI2X1 U9885 ( .A(\i_MIPS/n296 ), .B(\i_MIPS/n297 ), .S0(n3620), .Y(
        \i_MIPS/n424 ) );
  MXI2X1 U9886 ( .A(\i_MIPS/n292 ), .B(\i_MIPS/n293 ), .S0(n3619), .Y(
        \i_MIPS/n420 ) );
  MXI2X1 U9887 ( .A(\i_MIPS/n286 ), .B(\i_MIPS/n287 ), .S0(n3619), .Y(
        \i_MIPS/n414 ) );
  MXI2X1 U9888 ( .A(\i_MIPS/n276 ), .B(\i_MIPS/n277 ), .S0(n3621), .Y(
        \i_MIPS/n404 ) );
  MXI2X1 U9889 ( .A(\i_MIPS/n274 ), .B(\i_MIPS/n275 ), .S0(n3621), .Y(
        \i_MIPS/n402 ) );
  MXI2X1 U9890 ( .A(\i_MIPS/n272 ), .B(\i_MIPS/n273 ), .S0(n3621), .Y(
        \i_MIPS/n400 ) );
  MXI2X1 U9891 ( .A(\i_MIPS/n270 ), .B(\i_MIPS/n271 ), .S0(n3621), .Y(
        \i_MIPS/n398 ) );
  MXI2X1 U9892 ( .A(\i_MIPS/n268 ), .B(\i_MIPS/n269 ), .S0(n3621), .Y(
        \i_MIPS/n396 ) );
  MXI2X1 U9893 ( .A(\i_MIPS/n266 ), .B(\i_MIPS/n267 ), .S0(n3620), .Y(
        \i_MIPS/n394 ) );
  MXI2X1 U9894 ( .A(\i_MIPS/n264 ), .B(\i_MIPS/n265 ), .S0(n3620), .Y(
        \i_MIPS/n392 ) );
  MXI2X1 U9895 ( .A(\i_MIPS/n262 ), .B(\i_MIPS/n263 ), .S0(n3620), .Y(
        \i_MIPS/n390 ) );
  MXI2X1 U9896 ( .A(\i_MIPS/n260 ), .B(\i_MIPS/n261 ), .S0(n3619), .Y(
        \i_MIPS/n388 ) );
  MXI2X1 U9897 ( .A(\i_MIPS/n256 ), .B(\i_MIPS/n257 ), .S0(n3620), .Y(
        \i_MIPS/n384 ) );
  MXI2X1 U9898 ( .A(\i_MIPS/n252 ), .B(\i_MIPS/n253 ), .S0(n3621), .Y(
        \i_MIPS/n380 ) );
  MXI2X1 U9899 ( .A(\i_MIPS/n248 ), .B(\i_MIPS/n249 ), .S0(n3627), .Y(
        \i_MIPS/n376 ) );
  OAI2BB2XL U9900 ( .B0(n3017), .B1(n3772), .A0N(
        \i_MIPS/Register/register[3][22] ), .A1N(n3773), .Y(
        \i_MIPS/Register/n1034 ) );
  OAI2BB2XL U9901 ( .B0(n3660), .B1(n3771), .A0N(
        \i_MIPS/Register/register[3][23] ), .A1N(n3773), .Y(
        \i_MIPS/Register/n1035 ) );
  OAI2BB2XL U9902 ( .B0(n3683), .B1(n3780), .A0N(
        \i_MIPS/Register/register[0][10] ), .A1N(n3782), .Y(
        \i_MIPS/Register/n1118 ) );
  OAI2BB2XL U9903 ( .B0(n3682), .B1(n3777), .A0N(
        \i_MIPS/Register/register[1][10] ), .A1N(n3779), .Y(
        \i_MIPS/Register/n1086 ) );
  OAI2BB2XL U9904 ( .B0(n3682), .B1(n3768), .A0N(
        \i_MIPS/Register/register[4][10] ), .A1N(n3770), .Y(
        \i_MIPS/Register/n990 ) );
  OAI2BB2XL U9905 ( .B0(n3682), .B1(n3765), .A0N(
        \i_MIPS/Register/register[5][10] ), .A1N(n3767), .Y(
        \i_MIPS/Register/n958 ) );
  OAI2BB2XL U9906 ( .B0(n3682), .B1(n3759), .A0N(
        \i_MIPS/Register/register[7][10] ), .A1N(n3761), .Y(
        \i_MIPS/Register/n894 ) );
  OAI2BB2XL U9907 ( .B0(n3682), .B1(n3756), .A0N(
        \i_MIPS/Register/register[8][10] ), .A1N(n3758), .Y(
        \i_MIPS/Register/n862 ) );
  OAI2BB2XL U9908 ( .B0(n3682), .B1(n3753), .A0N(
        \i_MIPS/Register/register[9][10] ), .A1N(n3755), .Y(
        \i_MIPS/Register/n830 ) );
  OAI2BB2XL U9909 ( .B0(n3682), .B1(n3750), .A0N(
        \i_MIPS/Register/register[10][10] ), .A1N(n3752), .Y(
        \i_MIPS/Register/n798 ) );
  OAI2BB2XL U9910 ( .B0(n3682), .B1(n3747), .A0N(
        \i_MIPS/Register/register[11][10] ), .A1N(n3749), .Y(
        \i_MIPS/Register/n766 ) );
  OAI2BB2XL U9911 ( .B0(n3682), .B1(n3744), .A0N(
        \i_MIPS/Register/register[12][10] ), .A1N(n3746), .Y(
        \i_MIPS/Register/n734 ) );
  OAI2BB2XL U9912 ( .B0(n3682), .B1(n3741), .A0N(
        \i_MIPS/Register/register[13][10] ), .A1N(n3743), .Y(
        \i_MIPS/Register/n702 ) );
  OAI2BB2XL U9913 ( .B0(n3682), .B1(n3738), .A0N(
        \i_MIPS/Register/register[14][10] ), .A1N(n3740), .Y(
        \i_MIPS/Register/n670 ) );
  OAI2BB2XL U9914 ( .B0(n3682), .B1(n3735), .A0N(
        \i_MIPS/Register/register[15][10] ), .A1N(n3737), .Y(
        \i_MIPS/Register/n638 ) );
  OAI2BB2XL U9915 ( .B0(n3683), .B1(n3732), .A0N(
        \i_MIPS/Register/register[16][10] ), .A1N(n3734), .Y(
        \i_MIPS/Register/n606 ) );
  OAI2BB2XL U9916 ( .B0(n3683), .B1(n3729), .A0N(
        \i_MIPS/Register/register[17][10] ), .A1N(n3731), .Y(
        \i_MIPS/Register/n574 ) );
  OAI2BB2XL U9917 ( .B0(n3683), .B1(n3690), .A0N(
        \i_MIPS/Register/register[30][10] ), .A1N(n3692), .Y(
        \i_MIPS/Register/n158 ) );
  OAI2BB2XL U9918 ( .B0(n3683), .B1(n3774), .A0N(
        \i_MIPS/Register/register[2][10] ), .A1N(n3776), .Y(
        \i_MIPS/Register/n1054 ) );
  OAI2BB2XL U9919 ( .B0(n3683), .B1(n3771), .A0N(
        \i_MIPS/Register/register[3][10] ), .A1N(n3773), .Y(
        \i_MIPS/Register/n1022 ) );
  OAI2BB2XL U9920 ( .B0(n3683), .B1(n3762), .A0N(
        \i_MIPS/Register/register[6][10] ), .A1N(n3764), .Y(
        \i_MIPS/Register/n926 ) );
  OAI2BB2XL U9921 ( .B0(n3683), .B1(n3726), .A0N(
        \i_MIPS/Register/register[18][10] ), .A1N(n3728), .Y(
        \i_MIPS/Register/n542 ) );
  OAI2BB2XL U9922 ( .B0(n3683), .B1(n3723), .A0N(
        \i_MIPS/Register/register[19][10] ), .A1N(n3725), .Y(
        \i_MIPS/Register/n510 ) );
  OAI2BB2XL U9923 ( .B0(n3683), .B1(n3720), .A0N(
        \i_MIPS/Register/register[20][10] ), .A1N(n3722), .Y(
        \i_MIPS/Register/n478 ) );
  OAI2BB2XL U9924 ( .B0(n3683), .B1(n3717), .A0N(
        \i_MIPS/Register/register[21][10] ), .A1N(n3719), .Y(
        \i_MIPS/Register/n446 ) );
  OAI2BB2XL U9925 ( .B0(n3683), .B1(n3714), .A0N(
        \i_MIPS/Register/register[22][10] ), .A1N(n3716), .Y(
        \i_MIPS/Register/n414 ) );
  OAI2BB2XL U9926 ( .B0(n3683), .B1(n3711), .A0N(
        \i_MIPS/Register/register[23][10] ), .A1N(n3713), .Y(
        \i_MIPS/Register/n382 ) );
  OAI2BB2XL U9927 ( .B0(n3683), .B1(n3708), .A0N(
        \i_MIPS/Register/register[24][10] ), .A1N(n3710), .Y(
        \i_MIPS/Register/n350 ) );
  OAI2BB2XL U9928 ( .B0(n3683), .B1(n3705), .A0N(
        \i_MIPS/Register/register[25][10] ), .A1N(n3707), .Y(
        \i_MIPS/Register/n318 ) );
  OAI2BB2XL U9929 ( .B0(n3683), .B1(n3702), .A0N(
        \i_MIPS/Register/register[26][10] ), .A1N(n3704), .Y(
        \i_MIPS/Register/n286 ) );
  OAI2BB2XL U9930 ( .B0(n3683), .B1(n3699), .A0N(
        \i_MIPS/Register/register[27][10] ), .A1N(n3701), .Y(
        \i_MIPS/Register/n254 ) );
  OAI2BB2XL U9931 ( .B0(n3683), .B1(n3696), .A0N(
        \i_MIPS/Register/register[28][10] ), .A1N(n3698), .Y(
        \i_MIPS/Register/n222 ) );
  OAI2BB2XL U9932 ( .B0(n3683), .B1(n3693), .A0N(
        \i_MIPS/Register/register[29][10] ), .A1N(n3695), .Y(
        \i_MIPS/Register/n190 ) );
  OAI2BB2XL U9933 ( .B0(n3659), .B1(n3759), .A0N(
        \i_MIPS/Register/register[7][12] ), .A1N(n3761), .Y(
        \i_MIPS/Register/n896 ) );
  OAI2BB2XL U9934 ( .B0(n8729), .B1(n3756), .A0N(
        \i_MIPS/Register/register[8][12] ), .A1N(n3758), .Y(
        \i_MIPS/Register/n864 ) );
  OAI2BB2XL U9935 ( .B0(n8729), .B1(n3753), .A0N(
        \i_MIPS/Register/register[9][12] ), .A1N(n3755), .Y(
        \i_MIPS/Register/n832 ) );
  OAI2BB2XL U9936 ( .B0(n8729), .B1(n3750), .A0N(
        \i_MIPS/Register/register[10][12] ), .A1N(n3752), .Y(
        \i_MIPS/Register/n800 ) );
  OAI2BB2XL U9937 ( .B0(n8729), .B1(n3747), .A0N(
        \i_MIPS/Register/register[11][12] ), .A1N(n3749), .Y(
        \i_MIPS/Register/n768 ) );
  OAI2BB2XL U9938 ( .B0(n8729), .B1(n3744), .A0N(
        \i_MIPS/Register/register[12][12] ), .A1N(n3746), .Y(
        \i_MIPS/Register/n736 ) );
  OAI2BB2XL U9939 ( .B0(n3659), .B1(n3741), .A0N(
        \i_MIPS/Register/register[13][12] ), .A1N(n3743), .Y(
        \i_MIPS/Register/n704 ) );
  OAI2BB2XL U9940 ( .B0(n3659), .B1(n3738), .A0N(
        \i_MIPS/Register/register[14][12] ), .A1N(n3740), .Y(
        \i_MIPS/Register/n672 ) );
  OAI2BB2XL U9941 ( .B0(n3659), .B1(n3735), .A0N(
        \i_MIPS/Register/register[15][12] ), .A1N(n3737), .Y(
        \i_MIPS/Register/n640 ) );
  OAI2BB2XL U9942 ( .B0(n3659), .B1(n3732), .A0N(
        \i_MIPS/Register/register[16][12] ), .A1N(n3734), .Y(
        \i_MIPS/Register/n608 ) );
  OAI2BB2XL U9943 ( .B0(n3659), .B1(n3729), .A0N(
        \i_MIPS/Register/register[17][12] ), .A1N(n3731), .Y(
        \i_MIPS/Register/n576 ) );
  OAI2BB2XL U9944 ( .B0(n3659), .B1(n3726), .A0N(
        \i_MIPS/Register/register[18][12] ), .A1N(n3728), .Y(
        \i_MIPS/Register/n544 ) );
  OAI2BB2XL U9945 ( .B0(n3659), .B1(n3723), .A0N(
        \i_MIPS/Register/register[19][12] ), .A1N(n3725), .Y(
        \i_MIPS/Register/n512 ) );
  OAI2BB2XL U9946 ( .B0(n3659), .B1(n3720), .A0N(
        \i_MIPS/Register/register[20][12] ), .A1N(n3722), .Y(
        \i_MIPS/Register/n480 ) );
  OAI2BB2XL U9947 ( .B0(n3659), .B1(n3717), .A0N(
        \i_MIPS/Register/register[21][12] ), .A1N(n3719), .Y(
        \i_MIPS/Register/n448 ) );
  OAI2BB2XL U9948 ( .B0(n3659), .B1(n3714), .A0N(
        \i_MIPS/Register/register[22][12] ), .A1N(n3716), .Y(
        \i_MIPS/Register/n416 ) );
  OAI2BB2XL U9949 ( .B0(n3659), .B1(n3711), .A0N(
        \i_MIPS/Register/register[23][12] ), .A1N(n3713), .Y(
        \i_MIPS/Register/n384 ) );
  OAI2BB2XL U9950 ( .B0(n3659), .B1(n3708), .A0N(
        \i_MIPS/Register/register[24][12] ), .A1N(n3710), .Y(
        \i_MIPS/Register/n352 ) );
  OAI2BB2XL U9951 ( .B0(n3659), .B1(n3705), .A0N(
        \i_MIPS/Register/register[25][12] ), .A1N(n3707), .Y(
        \i_MIPS/Register/n320 ) );
  OAI2BB2XL U9952 ( .B0(n3659), .B1(n3702), .A0N(
        \i_MIPS/Register/register[26][12] ), .A1N(n3704), .Y(
        \i_MIPS/Register/n288 ) );
  OAI2BB2XL U9953 ( .B0(n3659), .B1(n3699), .A0N(
        \i_MIPS/Register/register[27][12] ), .A1N(n3701), .Y(
        \i_MIPS/Register/n256 ) );
  OAI2BB2XL U9954 ( .B0(n3659), .B1(n3696), .A0N(
        \i_MIPS/Register/register[28][12] ), .A1N(n3698), .Y(
        \i_MIPS/Register/n224 ) );
  OAI2BB2XL U9955 ( .B0(n3659), .B1(n3693), .A0N(
        \i_MIPS/Register/register[29][12] ), .A1N(n3695), .Y(
        \i_MIPS/Register/n192 ) );
  OAI2BB2XL U9956 ( .B0(n3659), .B1(n3690), .A0N(
        \i_MIPS/Register/register[30][12] ), .A1N(n3692), .Y(
        \i_MIPS/Register/n160 ) );
  OAI2BB2XL U9957 ( .B0(n3638), .B1(n3760), .A0N(
        \i_MIPS/Register/register[7][31] ), .A1N(n3760), .Y(
        \i_MIPS/Register/n915 ) );
  OAI2BB2XL U9958 ( .B0(n3643), .B1(n3759), .A0N(
        \i_MIPS/Register/register[7][28] ), .A1N(n3761), .Y(
        \i_MIPS/Register/n912 ) );
  OAI2BB2XL U9959 ( .B0(n3660), .B1(n3759), .A0N(
        \i_MIPS/Register/register[7][23] ), .A1N(n3761), .Y(
        \i_MIPS/Register/n907 ) );
  OAI2BB2XL U9960 ( .B0(n3017), .B1(n3760), .A0N(
        \i_MIPS/Register/register[7][22] ), .A1N(n3761), .Y(
        \i_MIPS/Register/n906 ) );
  OAI2BB2XL U9961 ( .B0(n3638), .B1(n3756), .A0N(
        \i_MIPS/Register/register[8][31] ), .A1N(n3757), .Y(
        \i_MIPS/Register/n883 ) );
  OAI2BB2XL U9962 ( .B0(n3643), .B1(n3757), .A0N(
        \i_MIPS/Register/register[8][28] ), .A1N(n3758), .Y(
        \i_MIPS/Register/n880 ) );
  OAI2BB2XL U9963 ( .B0(n3660), .B1(n3757), .A0N(
        \i_MIPS/Register/register[8][23] ), .A1N(n3758), .Y(
        \i_MIPS/Register/n875 ) );
  OAI2BB2XL U9964 ( .B0(n3017), .B1(n3757), .A0N(
        \i_MIPS/Register/register[8][22] ), .A1N(n3758), .Y(
        \i_MIPS/Register/n874 ) );
  OAI2BB2XL U9965 ( .B0(n3638), .B1(n42), .A0N(
        \i_MIPS/Register/register[9][31] ), .A1N(n3754), .Y(
        \i_MIPS/Register/n851 ) );
  OAI2BB2XL U9966 ( .B0(n3643), .B1(n42), .A0N(
        \i_MIPS/Register/register[9][28] ), .A1N(n3755), .Y(
        \i_MIPS/Register/n848 ) );
  OAI2BB2XL U9967 ( .B0(n3660), .B1(n3754), .A0N(
        \i_MIPS/Register/register[9][23] ), .A1N(n3755), .Y(
        \i_MIPS/Register/n843 ) );
  OAI2BB2XL U9968 ( .B0(n3017), .B1(n3754), .A0N(
        \i_MIPS/Register/register[9][22] ), .A1N(n3755), .Y(
        \i_MIPS/Register/n842 ) );
  OAI2BB2XL U9969 ( .B0(n3638), .B1(n41), .A0N(
        \i_MIPS/Register/register[10][31] ), .A1N(n3750), .Y(
        \i_MIPS/Register/n819 ) );
  OAI2BB2XL U9970 ( .B0(n3643), .B1(n41), .A0N(
        \i_MIPS/Register/register[10][28] ), .A1N(n3752), .Y(
        \i_MIPS/Register/n816 ) );
  OAI2BB2XL U9971 ( .B0(n3660), .B1(n3751), .A0N(
        \i_MIPS/Register/register[10][23] ), .A1N(n3752), .Y(
        \i_MIPS/Register/n811 ) );
  OAI2BB2XL U9972 ( .B0(n3017), .B1(n3751), .A0N(
        \i_MIPS/Register/register[10][22] ), .A1N(n3752), .Y(
        \i_MIPS/Register/n810 ) );
  OAI2BB2XL U9973 ( .B0(n3637), .B1(n40), .A0N(
        \i_MIPS/Register/register[11][31] ), .A1N(n3748), .Y(
        \i_MIPS/Register/n787 ) );
  OAI2BB2XL U9974 ( .B0(n3643), .B1(n40), .A0N(
        \i_MIPS/Register/register[11][28] ), .A1N(n3749), .Y(
        \i_MIPS/Register/n784 ) );
  OAI2BB2XL U9975 ( .B0(n3660), .B1(n3748), .A0N(
        \i_MIPS/Register/register[11][23] ), .A1N(n3749), .Y(
        \i_MIPS/Register/n779 ) );
  OAI2BB2XL U9976 ( .B0(n3017), .B1(n3748), .A0N(
        \i_MIPS/Register/register[11][22] ), .A1N(n3749), .Y(
        \i_MIPS/Register/n778 ) );
  OAI2BB2XL U9977 ( .B0(n3638), .B1(n39), .A0N(
        \i_MIPS/Register/register[12][31] ), .A1N(n3744), .Y(
        \i_MIPS/Register/n755 ) );
  OAI2BB2XL U9978 ( .B0(n3643), .B1(n39), .A0N(
        \i_MIPS/Register/register[12][28] ), .A1N(n3746), .Y(
        \i_MIPS/Register/n752 ) );
  OAI2BB2XL U9979 ( .B0(n3660), .B1(n3745), .A0N(
        \i_MIPS/Register/register[12][23] ), .A1N(n3746), .Y(
        \i_MIPS/Register/n747 ) );
  OAI2BB2XL U9980 ( .B0(n3017), .B1(n3745), .A0N(
        \i_MIPS/Register/register[12][22] ), .A1N(n3746), .Y(
        \i_MIPS/Register/n746 ) );
  OAI2BB2XL U9981 ( .B0(n3638), .B1(n38), .A0N(
        \i_MIPS/Register/register[13][31] ), .A1N(n3742), .Y(
        \i_MIPS/Register/n723 ) );
  OAI2BB2XL U9982 ( .B0(n3643), .B1(n38), .A0N(
        \i_MIPS/Register/register[13][28] ), .A1N(n3743), .Y(
        \i_MIPS/Register/n720 ) );
  OAI2BB2XL U9983 ( .B0(n3660), .B1(n3742), .A0N(
        \i_MIPS/Register/register[13][23] ), .A1N(n3743), .Y(
        \i_MIPS/Register/n715 ) );
  OAI2BB2XL U9984 ( .B0(n3017), .B1(n3742), .A0N(
        \i_MIPS/Register/register[13][22] ), .A1N(n3743), .Y(
        \i_MIPS/Register/n714 ) );
  OAI2BB2XL U9985 ( .B0(n3638), .B1(n37), .A0N(
        \i_MIPS/Register/register[14][31] ), .A1N(n3738), .Y(
        \i_MIPS/Register/n691 ) );
  OAI2BB2XL U9986 ( .B0(n3643), .B1(n37), .A0N(
        \i_MIPS/Register/register[14][28] ), .A1N(n3740), .Y(
        \i_MIPS/Register/n688 ) );
  OAI2BB2XL U9987 ( .B0(n3660), .B1(n3739), .A0N(
        \i_MIPS/Register/register[14][23] ), .A1N(n3739), .Y(
        \i_MIPS/Register/n683 ) );
  OAI2BB2XL U9988 ( .B0(n3017), .B1(n3739), .A0N(
        \i_MIPS/Register/register[14][22] ), .A1N(n3740), .Y(
        \i_MIPS/Register/n682 ) );
  OAI2BB2XL U9989 ( .B0(n3637), .B1(n36), .A0N(
        \i_MIPS/Register/register[15][31] ), .A1N(n3735), .Y(
        \i_MIPS/Register/n659 ) );
  OAI2BB2XL U9990 ( .B0(n3643), .B1(n36), .A0N(
        \i_MIPS/Register/register[15][28] ), .A1N(n3737), .Y(
        \i_MIPS/Register/n656 ) );
  OAI2BB2XL U9991 ( .B0(n3660), .B1(n3736), .A0N(
        \i_MIPS/Register/register[15][23] ), .A1N(n3737), .Y(
        \i_MIPS/Register/n651 ) );
  OAI2BB2XL U9992 ( .B0(n3017), .B1(n3736), .A0N(
        \i_MIPS/Register/register[15][22] ), .A1N(n3737), .Y(
        \i_MIPS/Register/n650 ) );
  OAI2BB2XL U9993 ( .B0(n3638), .B1(n35), .A0N(
        \i_MIPS/Register/register[16][31] ), .A1N(n3732), .Y(
        \i_MIPS/Register/n627 ) );
  OAI2BB2XL U9994 ( .B0(n8721), .B1(n35), .A0N(
        \i_MIPS/Register/register[16][28] ), .A1N(n3734), .Y(
        \i_MIPS/Register/n624 ) );
  OAI2BB2XL U9995 ( .B0(n3660), .B1(n3732), .A0N(
        \i_MIPS/Register/register[16][23] ), .A1N(n3732), .Y(
        \i_MIPS/Register/n619 ) );
  OAI2BB2XL U9996 ( .B0(n3017), .B1(n3733), .A0N(
        \i_MIPS/Register/register[16][22] ), .A1N(n3734), .Y(
        \i_MIPS/Register/n618 ) );
  OAI2BB2XL U9997 ( .B0(n3638), .B1(n34), .A0N(
        \i_MIPS/Register/register[17][31] ), .A1N(n3729), .Y(
        \i_MIPS/Register/n595 ) );
  OAI2BB2XL U9998 ( .B0(n8721), .B1(n34), .A0N(
        \i_MIPS/Register/register[17][28] ), .A1N(n3731), .Y(
        \i_MIPS/Register/n592 ) );
  OAI2BB2XL U9999 ( .B0(n3660), .B1(n3729), .A0N(
        \i_MIPS/Register/register[17][23] ), .A1N(n3731), .Y(
        \i_MIPS/Register/n587 ) );
  OAI2BB2XL U10000 ( .B0(n3017), .B1(n3730), .A0N(
        \i_MIPS/Register/register[17][22] ), .A1N(n3731), .Y(
        \i_MIPS/Register/n586 ) );
  OAI2BB2XL U10001 ( .B0(n3638), .B1(n3726), .A0N(
        \i_MIPS/Register/register[18][31] ), .A1N(n3727), .Y(
        \i_MIPS/Register/n563 ) );
  OAI2BB2XL U10002 ( .B0(n3643), .B1(n3727), .A0N(
        \i_MIPS/Register/register[18][28] ), .A1N(n3728), .Y(
        \i_MIPS/Register/n560 ) );
  OAI2BB2XL U10003 ( .B0(n3660), .B1(n3726), .A0N(
        \i_MIPS/Register/register[18][23] ), .A1N(n3727), .Y(
        \i_MIPS/Register/n555 ) );
  OAI2BB2XL U10004 ( .B0(n3017), .B1(n3727), .A0N(
        \i_MIPS/Register/register[18][22] ), .A1N(n3728), .Y(
        \i_MIPS/Register/n554 ) );
  OAI2BB2XL U10005 ( .B0(n3638), .B1(n3723), .A0N(
        \i_MIPS/Register/register[19][31] ), .A1N(n3723), .Y(
        \i_MIPS/Register/n531 ) );
  OAI2BB2XL U10006 ( .B0(n3643), .B1(n3724), .A0N(
        \i_MIPS/Register/register[19][28] ), .A1N(n3725), .Y(
        \i_MIPS/Register/n528 ) );
  OAI2BB2XL U10007 ( .B0(n3660), .B1(n3723), .A0N(
        \i_MIPS/Register/register[19][23] ), .A1N(n3723), .Y(
        \i_MIPS/Register/n523 ) );
  OAI2BB2XL U10008 ( .B0(n3017), .B1(n3724), .A0N(
        \i_MIPS/Register/register[19][22] ), .A1N(n3725), .Y(
        \i_MIPS/Register/n522 ) );
  OAI2BB2XL U10009 ( .B0(n3638), .B1(n3720), .A0N(
        \i_MIPS/Register/register[20][31] ), .A1N(n3721), .Y(
        \i_MIPS/Register/n499 ) );
  OAI2BB2XL U10010 ( .B0(n3643), .B1(n3721), .A0N(
        \i_MIPS/Register/register[20][28] ), .A1N(n3722), .Y(
        \i_MIPS/Register/n496 ) );
  OAI2BB2XL U10011 ( .B0(n3660), .B1(n3720), .A0N(
        \i_MIPS/Register/register[20][23] ), .A1N(n3721), .Y(
        \i_MIPS/Register/n491 ) );
  OAI2BB2XL U10012 ( .B0(n3017), .B1(n3721), .A0N(
        \i_MIPS/Register/register[20][22] ), .A1N(n3722), .Y(
        \i_MIPS/Register/n490 ) );
  OAI2BB2XL U10013 ( .B0(n3638), .B1(n3717), .A0N(
        \i_MIPS/Register/register[21][31] ), .A1N(n3717), .Y(
        \i_MIPS/Register/n467 ) );
  OAI2BB2XL U10014 ( .B0(n3643), .B1(n3718), .A0N(
        \i_MIPS/Register/register[21][28] ), .A1N(n3719), .Y(
        \i_MIPS/Register/n464 ) );
  OAI2BB2XL U10015 ( .B0(n3660), .B1(n3717), .A0N(
        \i_MIPS/Register/register[21][23] ), .A1N(n3717), .Y(
        \i_MIPS/Register/n459 ) );
  OAI2BB2XL U10016 ( .B0(n3017), .B1(n3718), .A0N(
        \i_MIPS/Register/register[21][22] ), .A1N(n3719), .Y(
        \i_MIPS/Register/n458 ) );
  OAI2BB2XL U10017 ( .B0(n3637), .B1(n3714), .A0N(
        \i_MIPS/Register/register[22][31] ), .A1N(n3715), .Y(
        \i_MIPS/Register/n435 ) );
  OAI2BB2XL U10018 ( .B0(n3643), .B1(n3715), .A0N(
        \i_MIPS/Register/register[22][28] ), .A1N(n3716), .Y(
        \i_MIPS/Register/n432 ) );
  OAI2BB2XL U10019 ( .B0(n3660), .B1(n3714), .A0N(
        \i_MIPS/Register/register[22][23] ), .A1N(n3715), .Y(
        \i_MIPS/Register/n427 ) );
  OAI2BB2XL U10020 ( .B0(n3017), .B1(n3715), .A0N(
        \i_MIPS/Register/register[22][22] ), .A1N(n3716), .Y(
        \i_MIPS/Register/n426 ) );
  OAI2BB2XL U10021 ( .B0(n3638), .B1(n3711), .A0N(
        \i_MIPS/Register/register[23][31] ), .A1N(n3712), .Y(
        \i_MIPS/Register/n403 ) );
  OAI2BB2XL U10022 ( .B0(n3643), .B1(n3712), .A0N(
        \i_MIPS/Register/register[23][28] ), .A1N(n3713), .Y(
        \i_MIPS/Register/n400 ) );
  OAI2BB2XL U10023 ( .B0(n3660), .B1(n3711), .A0N(
        \i_MIPS/Register/register[23][23] ), .A1N(n3711), .Y(
        \i_MIPS/Register/n395 ) );
  OAI2BB2XL U10024 ( .B0(n3017), .B1(n3712), .A0N(
        \i_MIPS/Register/register[23][22] ), .A1N(n3713), .Y(
        \i_MIPS/Register/n394 ) );
  OAI2BB2XL U10025 ( .B0(n3638), .B1(n3708), .A0N(
        \i_MIPS/Register/register[24][31] ), .A1N(n3708), .Y(
        \i_MIPS/Register/n371 ) );
  OAI2BB2XL U10026 ( .B0(n3643), .B1(n3709), .A0N(
        \i_MIPS/Register/register[24][28] ), .A1N(n3710), .Y(
        \i_MIPS/Register/n368 ) );
  OAI2BB2XL U10027 ( .B0(n3660), .B1(n3708), .A0N(
        \i_MIPS/Register/register[24][23] ), .A1N(n3709), .Y(
        \i_MIPS/Register/n363 ) );
  OAI2BB2XL U10028 ( .B0(n3017), .B1(n3709), .A0N(
        \i_MIPS/Register/register[24][22] ), .A1N(n3710), .Y(
        \i_MIPS/Register/n362 ) );
  OAI2BB2XL U10029 ( .B0(n3638), .B1(n3705), .A0N(
        \i_MIPS/Register/register[25][31] ), .A1N(n3705), .Y(
        \i_MIPS/Register/n339 ) );
  OAI2BB2XL U10030 ( .B0(n3643), .B1(n3706), .A0N(
        \i_MIPS/Register/register[25][28] ), .A1N(n3707), .Y(
        \i_MIPS/Register/n336 ) );
  OAI2BB2XL U10031 ( .B0(n3660), .B1(n3705), .A0N(
        \i_MIPS/Register/register[25][23] ), .A1N(n3706), .Y(
        \i_MIPS/Register/n331 ) );
  OAI2BB2XL U10032 ( .B0(n3017), .B1(n3706), .A0N(
        \i_MIPS/Register/register[25][22] ), .A1N(n3707), .Y(
        \i_MIPS/Register/n330 ) );
  OAI2BB2XL U10033 ( .B0(n3638), .B1(n3702), .A0N(
        \i_MIPS/Register/register[26][31] ), .A1N(n3703), .Y(
        \i_MIPS/Register/n307 ) );
  OAI2BB2XL U10034 ( .B0(n3643), .B1(n3703), .A0N(
        \i_MIPS/Register/register[26][28] ), .A1N(n3704), .Y(
        \i_MIPS/Register/n304 ) );
  OAI2BB2XL U10035 ( .B0(n3660), .B1(n3702), .A0N(
        \i_MIPS/Register/register[26][23] ), .A1N(n3703), .Y(
        \i_MIPS/Register/n299 ) );
  OAI2BB2XL U10036 ( .B0(n3017), .B1(n3703), .A0N(
        \i_MIPS/Register/register[26][22] ), .A1N(n3704), .Y(
        \i_MIPS/Register/n298 ) );
  OAI2BB2XL U10037 ( .B0(n3637), .B1(n3699), .A0N(
        \i_MIPS/Register/register[27][31] ), .A1N(n3699), .Y(
        \i_MIPS/Register/n275 ) );
  OAI2BB2XL U10038 ( .B0(n3643), .B1(n3700), .A0N(
        \i_MIPS/Register/register[27][28] ), .A1N(n3701), .Y(
        \i_MIPS/Register/n272 ) );
  OAI2BB2XL U10039 ( .B0(n3660), .B1(n3699), .A0N(
        \i_MIPS/Register/register[27][23] ), .A1N(n3700), .Y(
        \i_MIPS/Register/n267 ) );
  OAI2BB2XL U10040 ( .B0(n3017), .B1(n3700), .A0N(
        \i_MIPS/Register/register[27][22] ), .A1N(n3701), .Y(
        \i_MIPS/Register/n266 ) );
  OAI2BB2XL U10041 ( .B0(n3638), .B1(n3696), .A0N(
        \i_MIPS/Register/register[28][31] ), .A1N(n3696), .Y(
        \i_MIPS/Register/n243 ) );
  OAI2BB2XL U10042 ( .B0(n3643), .B1(n3697), .A0N(
        \i_MIPS/Register/register[28][28] ), .A1N(n3698), .Y(
        \i_MIPS/Register/n240 ) );
  OAI2BB2XL U10043 ( .B0(n3660), .B1(n3696), .A0N(
        \i_MIPS/Register/register[28][23] ), .A1N(n3697), .Y(
        \i_MIPS/Register/n235 ) );
  OAI2BB2XL U10044 ( .B0(n3017), .B1(n3697), .A0N(
        \i_MIPS/Register/register[28][22] ), .A1N(n3698), .Y(
        \i_MIPS/Register/n234 ) );
  OAI2BB2XL U10045 ( .B0(n3638), .B1(n3693), .A0N(
        \i_MIPS/Register/register[29][31] ), .A1N(n3693), .Y(
        \i_MIPS/Register/n211 ) );
  OAI2BB2XL U10046 ( .B0(n3643), .B1(n3694), .A0N(
        \i_MIPS/Register/register[29][28] ), .A1N(n3695), .Y(
        \i_MIPS/Register/n208 ) );
  OAI2BB2XL U10047 ( .B0(n3660), .B1(n3693), .A0N(
        \i_MIPS/Register/register[29][23] ), .A1N(n3693), .Y(
        \i_MIPS/Register/n203 ) );
  OAI2BB2XL U10048 ( .B0(n3017), .B1(n3694), .A0N(
        \i_MIPS/Register/register[29][22] ), .A1N(n3695), .Y(
        \i_MIPS/Register/n202 ) );
  OAI2BB2XL U10049 ( .B0(n3637), .B1(\i_MIPS/Register/n106 ), .A0N(
        \i_MIPS/Register/register[30][31] ), .A1N(n3691), .Y(
        \i_MIPS/Register/n179 ) );
  OAI2BB2XL U10050 ( .B0(n8721), .B1(\i_MIPS/Register/n106 ), .A0N(
        \i_MIPS/Register/register[30][28] ), .A1N(n3692), .Y(
        \i_MIPS/Register/n176 ) );
  OAI2BB2XL U10051 ( .B0(n3660), .B1(n3691), .A0N(
        \i_MIPS/Register/register[30][23] ), .A1N(n3691), .Y(
        \i_MIPS/Register/n171 ) );
  OAI2BB2XL U10052 ( .B0(n3017), .B1(n3691), .A0N(
        \i_MIPS/Register/register[30][22] ), .A1N(n3692), .Y(
        \i_MIPS/Register/n170 ) );
  OAI2BB2XL U10053 ( .B0(n3678), .B1(n3759), .A0N(
        \i_MIPS/Register/register[7][7] ), .A1N(n3761), .Y(
        \i_MIPS/Register/n891 ) );
  OAI2BB2XL U10054 ( .B0(n3677), .B1(n3756), .A0N(
        \i_MIPS/Register/register[8][7] ), .A1N(n3758), .Y(
        \i_MIPS/Register/n859 ) );
  OAI2BB2XL U10055 ( .B0(n3677), .B1(n3753), .A0N(
        \i_MIPS/Register/register[9][7] ), .A1N(n3755), .Y(
        \i_MIPS/Register/n827 ) );
  OAI2BB2XL U10056 ( .B0(n3677), .B1(n3750), .A0N(
        \i_MIPS/Register/register[10][7] ), .A1N(n3752), .Y(
        \i_MIPS/Register/n795 ) );
  OAI2BB2XL U10057 ( .B0(n3677), .B1(n3747), .A0N(
        \i_MIPS/Register/register[11][7] ), .A1N(n3749), .Y(
        \i_MIPS/Register/n763 ) );
  OAI2BB2XL U10058 ( .B0(n3677), .B1(n3744), .A0N(
        \i_MIPS/Register/register[12][7] ), .A1N(n3746), .Y(
        \i_MIPS/Register/n731 ) );
  OAI2BB2XL U10059 ( .B0(n3678), .B1(n3741), .A0N(
        \i_MIPS/Register/register[13][7] ), .A1N(n3743), .Y(
        \i_MIPS/Register/n699 ) );
  OAI2BB2XL U10060 ( .B0(n3678), .B1(n3738), .A0N(
        \i_MIPS/Register/register[14][7] ), .A1N(n3740), .Y(
        \i_MIPS/Register/n667 ) );
  OAI2BB2XL U10061 ( .B0(n3678), .B1(n3735), .A0N(
        \i_MIPS/Register/register[15][7] ), .A1N(n3737), .Y(
        \i_MIPS/Register/n635 ) );
  OAI2BB2XL U10062 ( .B0(n3678), .B1(n3732), .A0N(
        \i_MIPS/Register/register[16][7] ), .A1N(n3734), .Y(
        \i_MIPS/Register/n603 ) );
  OAI2BB2XL U10063 ( .B0(n3678), .B1(n3729), .A0N(
        \i_MIPS/Register/register[17][7] ), .A1N(n3731), .Y(
        \i_MIPS/Register/n571 ) );
  OAI2BB2XL U10064 ( .B0(n3678), .B1(n3726), .A0N(
        \i_MIPS/Register/register[18][7] ), .A1N(n3728), .Y(
        \i_MIPS/Register/n539 ) );
  OAI2BB2XL U10065 ( .B0(n3678), .B1(n3723), .A0N(
        \i_MIPS/Register/register[19][7] ), .A1N(n3725), .Y(
        \i_MIPS/Register/n507 ) );
  OAI2BB2XL U10066 ( .B0(n3678), .B1(n3720), .A0N(
        \i_MIPS/Register/register[20][7] ), .A1N(n3722), .Y(
        \i_MIPS/Register/n475 ) );
  OAI2BB2XL U10067 ( .B0(n3678), .B1(n3717), .A0N(
        \i_MIPS/Register/register[21][7] ), .A1N(n3719), .Y(
        \i_MIPS/Register/n443 ) );
  OAI2BB2XL U10068 ( .B0(n3678), .B1(n3714), .A0N(
        \i_MIPS/Register/register[22][7] ), .A1N(n3716), .Y(
        \i_MIPS/Register/n411 ) );
  OAI2BB2XL U10069 ( .B0(n3678), .B1(n3711), .A0N(
        \i_MIPS/Register/register[23][7] ), .A1N(n3713), .Y(
        \i_MIPS/Register/n379 ) );
  OAI2BB2XL U10070 ( .B0(n3678), .B1(n3708), .A0N(
        \i_MIPS/Register/register[24][7] ), .A1N(n3710), .Y(
        \i_MIPS/Register/n347 ) );
  OAI2BB2XL U10071 ( .B0(n3678), .B1(n3705), .A0N(
        \i_MIPS/Register/register[25][7] ), .A1N(n3707), .Y(
        \i_MIPS/Register/n315 ) );
  OAI2BB2XL U10072 ( .B0(n3678), .B1(n3702), .A0N(
        \i_MIPS/Register/register[26][7] ), .A1N(n3704), .Y(
        \i_MIPS/Register/n283 ) );
  OAI2BB2XL U10073 ( .B0(n3678), .B1(n3699), .A0N(
        \i_MIPS/Register/register[27][7] ), .A1N(n3701), .Y(
        \i_MIPS/Register/n251 ) );
  OAI2BB2XL U10074 ( .B0(n3678), .B1(n3696), .A0N(
        \i_MIPS/Register/register[28][7] ), .A1N(n3698), .Y(
        \i_MIPS/Register/n219 ) );
  OAI2BB2XL U10075 ( .B0(n3678), .B1(n3693), .A0N(
        \i_MIPS/Register/register[29][7] ), .A1N(n3695), .Y(
        \i_MIPS/Register/n187 ) );
  OAI2BB2XL U10076 ( .B0(n3678), .B1(n3690), .A0N(
        \i_MIPS/Register/register[30][7] ), .A1N(n3692), .Y(
        \i_MIPS/Register/n155 ) );
  OAI2BB2XL U10077 ( .B0(n3016), .B1(n3780), .A0N(
        \i_MIPS/Register/register[0][4] ), .A1N(n3780), .Y(
        \i_MIPS/Register/n1112 ) );
  OAI2BB2XL U10078 ( .B0(n3016), .B1(n3777), .A0N(
        \i_MIPS/Register/register[1][4] ), .A1N(n3777), .Y(
        \i_MIPS/Register/n1080 ) );
  OAI2BB2XL U10079 ( .B0(n3016), .B1(n3774), .A0N(
        \i_MIPS/Register/register[2][4] ), .A1N(n3774), .Y(
        \i_MIPS/Register/n1048 ) );
  OAI2BB2XL U10080 ( .B0(n3016), .B1(n3771), .A0N(
        \i_MIPS/Register/register[3][4] ), .A1N(n3771), .Y(
        \i_MIPS/Register/n1016 ) );
  OAI2BB2XL U10081 ( .B0(n3016), .B1(n3768), .A0N(
        \i_MIPS/Register/register[4][4] ), .A1N(n3768), .Y(
        \i_MIPS/Register/n984 ) );
  OAI2BB2XL U10082 ( .B0(n3016), .B1(n3765), .A0N(
        \i_MIPS/Register/register[5][4] ), .A1N(n3765), .Y(
        \i_MIPS/Register/n952 ) );
  OAI2BB2XL U10083 ( .B0(n3016), .B1(n3762), .A0N(
        \i_MIPS/Register/register[6][4] ), .A1N(n3762), .Y(
        \i_MIPS/Register/n920 ) );
  OAI2BB2XL U10084 ( .B0(n3016), .B1(n3759), .A0N(
        \i_MIPS/Register/register[7][4] ), .A1N(n3759), .Y(
        \i_MIPS/Register/n888 ) );
  OAI2BB2XL U10085 ( .B0(n3016), .B1(n3756), .A0N(
        \i_MIPS/Register/register[8][4] ), .A1N(n3757), .Y(
        \i_MIPS/Register/n856 ) );
  OAI2BB2XL U10086 ( .B0(n3016), .B1(n3753), .A0N(
        \i_MIPS/Register/register[9][4] ), .A1N(n3754), .Y(
        \i_MIPS/Register/n824 ) );
  OAI2BB2XL U10087 ( .B0(n3016), .B1(n3750), .A0N(
        \i_MIPS/Register/register[10][4] ), .A1N(n3751), .Y(
        \i_MIPS/Register/n792 ) );
  OAI2BB2XL U10088 ( .B0(n3016), .B1(n3747), .A0N(
        \i_MIPS/Register/register[11][4] ), .A1N(n3748), .Y(
        \i_MIPS/Register/n760 ) );
  OAI2BB2XL U10089 ( .B0(n3016), .B1(n3744), .A0N(
        \i_MIPS/Register/register[12][4] ), .A1N(n3745), .Y(
        \i_MIPS/Register/n728 ) );
  OAI2BB2XL U10090 ( .B0(n3016), .B1(n3741), .A0N(
        \i_MIPS/Register/register[13][4] ), .A1N(n3742), .Y(
        \i_MIPS/Register/n696 ) );
  OAI2BB2XL U10091 ( .B0(n3668), .B1(n3738), .A0N(
        \i_MIPS/Register/register[14][4] ), .A1N(n3739), .Y(
        \i_MIPS/Register/n664 ) );
  OAI2BB2XL U10092 ( .B0(n3016), .B1(n3735), .A0N(
        \i_MIPS/Register/register[15][4] ), .A1N(n3736), .Y(
        \i_MIPS/Register/n632 ) );
  OAI2BB2XL U10093 ( .B0(n8735), .B1(n3732), .A0N(
        \i_MIPS/Register/register[16][4] ), .A1N(n3732), .Y(
        \i_MIPS/Register/n600 ) );
  OAI2BB2XL U10094 ( .B0(n3668), .B1(n3729), .A0N(
        \i_MIPS/Register/register[17][4] ), .A1N(n3730), .Y(
        \i_MIPS/Register/n568 ) );
  OAI2BB2XL U10095 ( .B0(n3016), .B1(n3726), .A0N(
        \i_MIPS/Register/register[18][4] ), .A1N(n3726), .Y(
        \i_MIPS/Register/n536 ) );
  OAI2BB2XL U10096 ( .B0(n3016), .B1(n3723), .A0N(
        \i_MIPS/Register/register[19][4] ), .A1N(n3723), .Y(
        \i_MIPS/Register/n504 ) );
  OAI2BB2XL U10097 ( .B0(n3016), .B1(n3720), .A0N(
        \i_MIPS/Register/register[20][4] ), .A1N(n3720), .Y(
        \i_MIPS/Register/n472 ) );
  OAI2BB2XL U10098 ( .B0(n3016), .B1(n3717), .A0N(
        \i_MIPS/Register/register[21][4] ), .A1N(n3717), .Y(
        \i_MIPS/Register/n440 ) );
  OAI2BB2XL U10099 ( .B0(n3016), .B1(n3714), .A0N(
        \i_MIPS/Register/register[22][4] ), .A1N(n3714), .Y(
        \i_MIPS/Register/n408 ) );
  OAI2BB2XL U10100 ( .B0(n3016), .B1(n3690), .A0N(
        \i_MIPS/Register/register[30][4] ), .A1N(n3691), .Y(
        \i_MIPS/Register/n152 ) );
  OAI2BB2XL U10101 ( .B0(n3686), .B1(n3760), .A0N(
        \i_MIPS/Register/register[7][20] ), .A1N(n3761), .Y(
        \i_MIPS/Register/n904 ) );
  OAI2BB2XL U10102 ( .B0(n3686), .B1(n3757), .A0N(
        \i_MIPS/Register/register[8][20] ), .A1N(n3756), .Y(
        \i_MIPS/Register/n872 ) );
  OAI2BB2XL U10103 ( .B0(n8744), .B1(n3754), .A0N(
        \i_MIPS/Register/register[9][20] ), .A1N(n3753), .Y(
        \i_MIPS/Register/n840 ) );
  OAI2BB2XL U10104 ( .B0(n8744), .B1(n3751), .A0N(
        \i_MIPS/Register/register[10][20] ), .A1N(n3750), .Y(
        \i_MIPS/Register/n808 ) );
  OAI2BB2XL U10105 ( .B0(n8744), .B1(n3748), .A0N(
        \i_MIPS/Register/register[11][20] ), .A1N(n3747), .Y(
        \i_MIPS/Register/n776 ) );
  OAI2BB2XL U10106 ( .B0(n8744), .B1(n3745), .A0N(
        \i_MIPS/Register/register[12][20] ), .A1N(n3744), .Y(
        \i_MIPS/Register/n744 ) );
  OAI2BB2XL U10107 ( .B0(n8744), .B1(n3742), .A0N(
        \i_MIPS/Register/register[13][20] ), .A1N(n3741), .Y(
        \i_MIPS/Register/n712 ) );
  OAI2BB2XL U10108 ( .B0(n8744), .B1(n3739), .A0N(
        \i_MIPS/Register/register[14][20] ), .A1N(n3738), .Y(
        \i_MIPS/Register/n680 ) );
  OAI2BB2XL U10109 ( .B0(n8744), .B1(n3736), .A0N(
        \i_MIPS/Register/register[15][20] ), .A1N(n3735), .Y(
        \i_MIPS/Register/n648 ) );
  OAI2BB2XL U10110 ( .B0(n8744), .B1(n3733), .A0N(
        \i_MIPS/Register/register[16][20] ), .A1N(n3733), .Y(
        \i_MIPS/Register/n616 ) );
  OAI2BB2XL U10111 ( .B0(n8744), .B1(n3730), .A0N(
        \i_MIPS/Register/register[17][20] ), .A1N(n3730), .Y(
        \i_MIPS/Register/n584 ) );
  OAI2BB2XL U10112 ( .B0(n3686), .B1(n3727), .A0N(
        \i_MIPS/Register/register[18][20] ), .A1N(n3728), .Y(
        \i_MIPS/Register/n552 ) );
  OAI2BB2XL U10113 ( .B0(n3686), .B1(n3724), .A0N(
        \i_MIPS/Register/register[19][20] ), .A1N(n3725), .Y(
        \i_MIPS/Register/n520 ) );
  OAI2BB2XL U10114 ( .B0(n3686), .B1(n3721), .A0N(
        \i_MIPS/Register/register[20][20] ), .A1N(n3722), .Y(
        \i_MIPS/Register/n488 ) );
  OAI2BB2XL U10115 ( .B0(n3686), .B1(n3718), .A0N(
        \i_MIPS/Register/register[21][20] ), .A1N(n3719), .Y(
        \i_MIPS/Register/n456 ) );
  OAI2BB2XL U10116 ( .B0(n3686), .B1(n3715), .A0N(
        \i_MIPS/Register/register[22][20] ), .A1N(n3716), .Y(
        \i_MIPS/Register/n424 ) );
  OAI2BB2XL U10117 ( .B0(n3686), .B1(n3712), .A0N(
        \i_MIPS/Register/register[23][20] ), .A1N(n3713), .Y(
        \i_MIPS/Register/n392 ) );
  OAI2BB2XL U10118 ( .B0(n3686), .B1(n3709), .A0N(
        \i_MIPS/Register/register[24][20] ), .A1N(n3710), .Y(
        \i_MIPS/Register/n360 ) );
  OAI2BB2XL U10119 ( .B0(n3686), .B1(n3706), .A0N(
        \i_MIPS/Register/register[25][20] ), .A1N(n3707), .Y(
        \i_MIPS/Register/n328 ) );
  OAI2BB2XL U10120 ( .B0(n3686), .B1(n3703), .A0N(
        \i_MIPS/Register/register[26][20] ), .A1N(n3704), .Y(
        \i_MIPS/Register/n296 ) );
  OAI2BB2XL U10121 ( .B0(n3686), .B1(n3700), .A0N(
        \i_MIPS/Register/register[27][20] ), .A1N(n3701), .Y(
        \i_MIPS/Register/n264 ) );
  OAI2BB2XL U10122 ( .B0(n3686), .B1(n3697), .A0N(
        \i_MIPS/Register/register[28][20] ), .A1N(n3698), .Y(
        \i_MIPS/Register/n232 ) );
  OAI2BB2XL U10123 ( .B0(n3686), .B1(n3694), .A0N(
        \i_MIPS/Register/register[29][20] ), .A1N(n3695), .Y(
        \i_MIPS/Register/n200 ) );
  OAI2BB2XL U10124 ( .B0(n8744), .B1(n3691), .A0N(
        \i_MIPS/Register/register[30][20] ), .A1N(n3690), .Y(
        \i_MIPS/Register/n168 ) );
  OAI2BB2XL U10125 ( .B0(n3660), .B1(n3765), .A0N(
        \i_MIPS/Register/register[5][23] ), .A1N(n3767), .Y(
        \i_MIPS/Register/n971 ) );
  OAI2BB2XL U10126 ( .B0(n3017), .B1(n3766), .A0N(
        \i_MIPS/Register/register[5][22] ), .A1N(n3767), .Y(
        \i_MIPS/Register/n970 ) );
  OAI2BB2XL U10127 ( .B0(n3660), .B1(n3762), .A0N(
        \i_MIPS/Register/register[6][23] ), .A1N(n3764), .Y(
        \i_MIPS/Register/n939 ) );
  OAI2BB2XL U10128 ( .B0(n3017), .B1(n3763), .A0N(
        \i_MIPS/Register/register[6][22] ), .A1N(n3764), .Y(
        \i_MIPS/Register/n938 ) );
  OAI2BB2XL U10129 ( .B0(n3638), .B1(n51), .A0N(
        \i_MIPS/Register/register[0][31] ), .A1N(n3781), .Y(
        \i_MIPS/Register/n1139 ) );
  OAI2BB2XL U10130 ( .B0(n3643), .B1(n51), .A0N(
        \i_MIPS/Register/register[0][28] ), .A1N(n3782), .Y(
        \i_MIPS/Register/n1136 ) );
  OAI2BB2XL U10131 ( .B0(n3638), .B1(n50), .A0N(
        \i_MIPS/Register/register[1][31] ), .A1N(n3777), .Y(
        \i_MIPS/Register/n1107 ) );
  OAI2BB2XL U10132 ( .B0(n3643), .B1(n50), .A0N(
        \i_MIPS/Register/register[1][28] ), .A1N(n3779), .Y(
        \i_MIPS/Register/n1104 ) );
  OAI2BB2XL U10133 ( .B0(n3638), .B1(n49), .A0N(
        \i_MIPS/Register/register[2][31] ), .A1N(n3775), .Y(
        \i_MIPS/Register/n1075 ) );
  OAI2BB2XL U10134 ( .B0(n3643), .B1(n49), .A0N(
        \i_MIPS/Register/register[2][28] ), .A1N(n3776), .Y(
        \i_MIPS/Register/n1072 ) );
  OAI2BB2XL U10135 ( .B0(n3638), .B1(n48), .A0N(
        \i_MIPS/Register/register[3][31] ), .A1N(n3771), .Y(
        \i_MIPS/Register/n1043 ) );
  OAI2BB2XL U10136 ( .B0(n3643), .B1(n48), .A0N(
        \i_MIPS/Register/register[3][28] ), .A1N(n3773), .Y(
        \i_MIPS/Register/n1040 ) );
  OAI2BB2XL U10137 ( .B0(n3637), .B1(n47), .A0N(
        \i_MIPS/Register/register[4][31] ), .A1N(n3768), .Y(
        \i_MIPS/Register/n1011 ) );
  OAI2BB2XL U10138 ( .B0(n3643), .B1(n47), .A0N(
        \i_MIPS/Register/register[4][28] ), .A1N(n3770), .Y(
        \i_MIPS/Register/n1008 ) );
  OAI2BB2XL U10139 ( .B0(n3638), .B1(n46), .A0N(
        \i_MIPS/Register/register[5][31] ), .A1N(n3765), .Y(
        \i_MIPS/Register/n979 ) );
  OAI2BB2XL U10140 ( .B0(n3643), .B1(n46), .A0N(
        \i_MIPS/Register/register[5][28] ), .A1N(n3767), .Y(
        \i_MIPS/Register/n976 ) );
  OAI2BB2XL U10141 ( .B0(n3638), .B1(n45), .A0N(
        \i_MIPS/Register/register[6][31] ), .A1N(n3762), .Y(
        \i_MIPS/Register/n947 ) );
  OAI2BB2XL U10142 ( .B0(n3643), .B1(n45), .A0N(
        \i_MIPS/Register/register[6][28] ), .A1N(n3764), .Y(
        \i_MIPS/Register/n944 ) );
  OAI2BB2XL U10143 ( .B0(n3668), .B1(n3711), .A0N(
        \i_MIPS/Register/register[23][4] ), .A1N(n3712), .Y(
        \i_MIPS/Register/n376 ) );
  OAI2BB2XL U10144 ( .B0(n3668), .B1(n3708), .A0N(
        \i_MIPS/Register/register[24][4] ), .A1N(n3708), .Y(
        \i_MIPS/Register/n344 ) );
  OAI2BB2XL U10145 ( .B0(n3668), .B1(n3705), .A0N(
        \i_MIPS/Register/register[25][4] ), .A1N(n3705), .Y(
        \i_MIPS/Register/n312 ) );
  OAI2BB2XL U10146 ( .B0(n3668), .B1(n3702), .A0N(
        \i_MIPS/Register/register[26][4] ), .A1N(n3702), .Y(
        \i_MIPS/Register/n280 ) );
  OAI2BB2XL U10147 ( .B0(n3668), .B1(n3699), .A0N(
        \i_MIPS/Register/register[27][4] ), .A1N(n3699), .Y(
        \i_MIPS/Register/n248 ) );
  OAI2BB2XL U10148 ( .B0(n3668), .B1(n3696), .A0N(
        \i_MIPS/Register/register[28][4] ), .A1N(n3696), .Y(
        \i_MIPS/Register/n216 ) );
  OAI2BB2XL U10149 ( .B0(n3668), .B1(n3693), .A0N(
        \i_MIPS/Register/register[29][4] ), .A1N(n3693), .Y(
        \i_MIPS/Register/n184 ) );
  OAI2BB2XL U10150 ( .B0(n8744), .B1(n3781), .A0N(
        \i_MIPS/Register/register[0][20] ), .A1N(n3781), .Y(
        \i_MIPS/Register/n1128 ) );
  OAI2BB2XL U10151 ( .B0(n8744), .B1(n3778), .A0N(
        \i_MIPS/Register/register[1][20] ), .A1N(n3778), .Y(
        \i_MIPS/Register/n1096 ) );
  OAI2BB2XL U10152 ( .B0(n8744), .B1(n3775), .A0N(
        \i_MIPS/Register/register[2][20] ), .A1N(n3775), .Y(
        \i_MIPS/Register/n1064 ) );
  OAI2BB2XL U10153 ( .B0(n8744), .B1(n3772), .A0N(
        \i_MIPS/Register/register[3][20] ), .A1N(n3772), .Y(
        \i_MIPS/Register/n1032 ) );
  OAI2BB2XL U10154 ( .B0(n8744), .B1(n3769), .A0N(
        \i_MIPS/Register/register[4][20] ), .A1N(n3769), .Y(
        \i_MIPS/Register/n1000 ) );
  OAI2BB2XL U10155 ( .B0(n8744), .B1(n3766), .A0N(
        \i_MIPS/Register/register[5][20] ), .A1N(n3766), .Y(
        \i_MIPS/Register/n968 ) );
  OAI2BB2XL U10156 ( .B0(n8744), .B1(n3763), .A0N(
        \i_MIPS/Register/register[6][20] ), .A1N(n3763), .Y(
        \i_MIPS/Register/n936 ) );
  NAND4BX1 U10157 ( .AN(n5092), .B(n5091), .C(n5090), .D(n5089), .Y(n5103) );
  NAND4BX1 U10158 ( .AN(n5101), .B(n5100), .C(n5099), .D(n5098), .Y(n5102) );
  CLKMX2X2 U10159 ( .A(n5377), .B(n5376), .S0(n4014), .Y(n5378) );
  NAND4BX1 U10160 ( .AN(n5366), .B(n5365), .C(n5364), .D(n5363), .Y(n5377) );
  NAND4BX1 U10161 ( .AN(n5375), .B(n5374), .C(n5373), .D(n5372), .Y(n5376) );
  CLKMX2X2 U10162 ( .A(n5596), .B(n5595), .S0(n4014), .Y(n5597) );
  NAND4BX1 U10163 ( .AN(n5585), .B(n5584), .C(n5583), .D(n5582), .Y(n5596) );
  NAND4BX1 U10164 ( .AN(n5594), .B(n5593), .C(n5592), .D(n5591), .Y(n5595) );
  OA22X1 U10165 ( .A0(\i_MIPS/Register/register[4][15] ), .A1(n3180), .B0(
        \i_MIPS/Register/register[12][15] ), .B1(n3176), .Y(n5584) );
  CLKMX2X2 U10166 ( .A(n6948), .B(n6947), .S0(n4015), .Y(n6949) );
  NAND4BX1 U10167 ( .AN(n6937), .B(n6936), .C(n6935), .D(n6934), .Y(n6948) );
  NAND4BX1 U10168 ( .AN(n6946), .B(n6945), .C(n6944), .D(n6943), .Y(n6947) );
  OA22X1 U10169 ( .A0(\i_MIPS/Register/register[4][16] ), .A1(n3181), .B0(
        \i_MIPS/Register/register[12][16] ), .B1(n3176), .Y(n6936) );
  CLKMX2X2 U10170 ( .A(n5575), .B(n5574), .S0(n4012), .Y(n5576) );
  NAND4BX1 U10171 ( .AN(n5564), .B(n5563), .C(n5562), .D(n5561), .Y(n5575) );
  NAND4BX1 U10172 ( .AN(n5573), .B(n5572), .C(n5571), .D(n5570), .Y(n5574) );
  OA22X1 U10173 ( .A0(\i_MIPS/Register/register[4][15] ), .A1(n3129), .B0(
        \i_MIPS/Register/register[12][15] ), .B1(n3126), .Y(n5563) );
  AND3X2 U10174 ( .A(n3611), .B(\i_MIPS/n326 ), .C(\i_MIPS/n330 ), .Y(n7634)
         );
  MX2XL U10175 ( .A(n10298), .B(n8300), .S0(n3627), .Y(\i_MIPS/n439 ) );
  OAI222XL U10176 ( .A0(n3584), .A1(n68), .B0(n3640), .B1(n3582), .C0(n3688), 
        .C1(\i_MIPS/n210 ), .Y(n8774) );
  OAI222XL U10177 ( .A0(n3584), .A1(n69), .B0(n3642), .B1(n3583), .C0(n3688), 
        .C1(\i_MIPS/n209 ), .Y(n8775) );
  MX2XL U10178 ( .A(DCACHE_addr[1]), .B(n8240), .S0(n3624), .Y(\i_MIPS/n466 )
         );
  MX2XL U10179 ( .A(n10323), .B(n8233), .S0(n3624), .Y(\i_MIPS/n467 ) );
  MX2XL U10180 ( .A(n10309), .B(n8015), .S0(n3624), .Y(\i_MIPS/n450 ) );
  MX2XL U10181 ( .A(n10305), .B(n8227), .S0(n3625), .Y(\i_MIPS/n446 ) );
  MX2XL U10182 ( .A(n10302), .B(n8263), .S0(n3625), .Y(\i_MIPS/n443 ) );
  MX2XL U10183 ( .A(n10301), .B(n8167), .S0(n3625), .Y(\i_MIPS/n442 ) );
  MX2XL U10184 ( .A(n10300), .B(n8266), .S0(n3625), .Y(\i_MIPS/n441 ) );
  CLKBUFX3 U10185 ( .A(\i_MIPS/EX_MEM_1 ), .Y(n4023) );
  OA22X1 U10186 ( .A0(n3568), .A1(n175), .B0(n3526), .B1(n1444), .Y(n4389) );
  OA22X1 U10187 ( .A0(n3570), .A1(n811), .B0(n3510), .B1(n1744), .Y(n7165) );
  OA22X1 U10188 ( .A0(n3570), .A1(n812), .B0(n3510), .B1(n1745), .Y(n7180) );
  OA22X1 U10189 ( .A0(n3570), .A1(n813), .B0(n3510), .B1(n1746), .Y(n7170) );
  OA22X1 U10190 ( .A0(n3570), .A1(n814), .B0(n3510), .B1(n1747), .Y(n7175) );
  OA22X1 U10191 ( .A0(n3552), .A1(n815), .B0(n3510), .B1(n1748), .Y(n7237) );
  OA22X1 U10192 ( .A0(n3552), .A1(n816), .B0(n3510), .B1(n1749), .Y(n7247) );
  OA22X1 U10193 ( .A0(n3552), .A1(n817), .B0(n3510), .B1(n1750), .Y(n7252) );
  OA22X1 U10194 ( .A0(n3552), .A1(n818), .B0(n3510), .B1(n1751), .Y(n7242) );
  OA22X1 U10195 ( .A0(n3552), .A1(n819), .B0(n3510), .B1(n1752), .Y(n7285) );
  OA22X1 U10196 ( .A0(n3552), .A1(n820), .B0(n3510), .B1(n1753), .Y(n7293) );
  OA22X1 U10197 ( .A0(n3552), .A1(n821), .B0(n3510), .B1(n1754), .Y(n7289) );
  OA22X1 U10198 ( .A0(n3552), .A1(n822), .B0(n3513), .B1(n1755), .Y(n7261) );
  OA22X1 U10199 ( .A0(n3552), .A1(n823), .B0(n3510), .B1(n1756), .Y(n7271) );
  OA22X1 U10200 ( .A0(n3552), .A1(n824), .B0(n3510), .B1(n1757), .Y(n7276) );
  OA22X1 U10201 ( .A0(n3552), .A1(n825), .B0(n3510), .B1(n1758), .Y(n7266) );
  OA22X1 U10202 ( .A0(n3552), .A1(n826), .B0(n3510), .B1(n1759), .Y(n7213) );
  OA22X1 U10203 ( .A0(n3570), .A1(n827), .B0(n3513), .B1(n1760), .Y(n7228) );
  OA22X1 U10204 ( .A0(n3551), .A1(n828), .B0(n3510), .B1(n1761), .Y(n7218) );
  OA22X1 U10205 ( .A0(n3570), .A1(n829), .B0(n3510), .B1(n1762), .Y(n7223) );
  OA22X1 U10206 ( .A0(n3552), .A1(n830), .B0(n3509), .B1(n1763), .Y(n7189) );
  OA22X1 U10207 ( .A0(n3552), .A1(n831), .B0(n3510), .B1(n1764), .Y(n7204) );
  OA22X1 U10208 ( .A0(n3570), .A1(n832), .B0(n3510), .B1(n1765), .Y(n7194) );
  OA22X1 U10209 ( .A0(n3570), .A1(n833), .B0(n3510), .B1(n1766), .Y(n7199) );
  OA22X1 U10210 ( .A0(n3552), .A1(n834), .B0(n3520), .B1(n1767), .Y(n7131) );
  OA22X1 U10211 ( .A0(n3552), .A1(n835), .B0(n3515), .B1(n1768), .Y(n7121) );
  OA22X1 U10212 ( .A0(n3570), .A1(n836), .B0(n3509), .B1(n1769), .Y(n7126) );
  OA22X1 U10213 ( .A0(n3551), .A1(n837), .B0(n3522), .B1(n1770), .Y(n7116) );
  OA22X1 U10214 ( .A0(n3551), .A1(n838), .B0(n3509), .B1(n1771), .Y(n7449) );
  OA22X1 U10215 ( .A0(n3552), .A1(n839), .B0(n3510), .B1(n1772), .Y(n7454) );
  OA22X1 U10216 ( .A0(n3551), .A1(n840), .B0(n3509), .B1(n1773), .Y(n7444) );
  OA22X1 U10217 ( .A0(n3551), .A1(n841), .B0(n3509), .B1(n1774), .Y(n7473) );
  OA22X1 U10218 ( .A0(n3552), .A1(n842), .B0(n3511), .B1(n1775), .Y(n7463) );
  OA22X1 U10219 ( .A0(n3570), .A1(n843), .B0(n3515), .B1(n1776), .Y(n7468) );
  OA22X1 U10220 ( .A0(n3551), .A1(n844), .B0(n3511), .B1(n1777), .Y(n7155) );
  OA22X1 U10221 ( .A0(n3570), .A1(n845), .B0(n3509), .B1(n1778), .Y(n7145) );
  OA22X1 U10222 ( .A0(n3552), .A1(n846), .B0(n3509), .B1(n1779), .Y(n7150) );
  OA22X1 U10223 ( .A0(n3552), .A1(n847), .B0(n3520), .B1(n1780), .Y(n7140) );
  OA22X1 U10224 ( .A0(n3551), .A1(n848), .B0(n3522), .B1(n1781), .Y(n4584) );
  OA22X1 U10225 ( .A0(n3551), .A1(n849), .B0(n3523), .B1(n1782), .Y(n7107) );
  OA22X1 U10226 ( .A0(n3551), .A1(n850), .B0(n3523), .B1(n1783), .Y(n7097) );
  OA22X1 U10227 ( .A0(n3551), .A1(n851), .B0(n3509), .B1(n1784), .Y(n7102) );
  OA22X1 U10228 ( .A0(n3551), .A1(n852), .B0(n3512), .B1(n1785), .Y(n7092) );
  OA22X1 U10229 ( .A0(\i_MIPS/Register/register[16][8] ), .A1(n3136), .B0(
        \i_MIPS/Register/register[24][8] ), .B1(n3133), .Y(n6160) );
  OA22X1 U10230 ( .A0(\i_MIPS/Register/register[0][8] ), .A1(n3134), .B0(
        \i_MIPS/Register/register[8][8] ), .B1(n3132), .Y(n6151) );
  OA22X1 U10231 ( .A0(\i_MIPS/Register/register[16][9] ), .A1(n3136), .B0(
        \i_MIPS/Register/register[24][9] ), .B1(n3133), .Y(n6229) );
  OA22X1 U10232 ( .A0(\i_MIPS/Register/register[0][9] ), .A1(n3136), .B0(
        \i_MIPS/Register/register[8][9] ), .B1(n3133), .Y(n6220) );
  OA22X1 U10233 ( .A0(\i_MIPS/Register/register[0][9] ), .A1(n3187), .B0(
        \i_MIPS/Register/register[8][9] ), .B1(n3184), .Y(n6241) );
  OA22X1 U10234 ( .A0(\i_MIPS/Register/register[16][13] ), .A1(n3136), .B0(
        \i_MIPS/Register/register[24][13] ), .B1(n3133), .Y(n6427) );
  OA22X1 U10235 ( .A0(\i_MIPS/Register/register[0][13] ), .A1(n3136), .B0(
        \i_MIPS/Register/register[8][13] ), .B1(n3133), .Y(n6418) );
  OA22X1 U10236 ( .A0(\i_MIPS/Register/register[16][14] ), .A1(n3136), .B0(
        \i_MIPS/Register/register[24][14] ), .B1(n3133), .Y(n6361) );
  OA22X1 U10237 ( .A0(\i_MIPS/Register/register[0][14] ), .A1(n3136), .B0(
        \i_MIPS/Register/register[8][14] ), .B1(n3133), .Y(n6352) );
  OA22X1 U10238 ( .A0(\i_MIPS/Register/register[16][11] ), .A1(n3135), .B0(
        \i_MIPS/Register/register[24][11] ), .B1(n2788), .Y(n5291) );
  OA22X1 U10239 ( .A0(\i_MIPS/Register/register[0][11] ), .A1(n3135), .B0(
        \i_MIPS/Register/register[8][11] ), .B1(n3131), .Y(n5282) );
  OA22X1 U10240 ( .A0(\i_MIPS/Register/register[16][10] ), .A1(n3185), .B0(
        \i_MIPS/Register/register[24][10] ), .B1(n3182), .Y(n5247) );
  OA22X1 U10241 ( .A0(\i_MIPS/Register/register[0][10] ), .A1(n3187), .B0(
        \i_MIPS/Register/register[8][10] ), .B1(n3184), .Y(n5238) );
  OA22X1 U10242 ( .A0(\i_MIPS/Register/register[16][10] ), .A1(n3135), .B0(
        \i_MIPS/Register/register[24][10] ), .B1(n3132), .Y(n5226) );
  OA22X1 U10243 ( .A0(\i_MIPS/Register/register[0][10] ), .A1(n3134), .B0(
        \i_MIPS/Register/register[8][10] ), .B1(n3131), .Y(n5217) );
  OA22X1 U10244 ( .A0(\i_MIPS/Register/register[16][5] ), .A1(n3185), .B0(
        \i_MIPS/Register/register[24][5] ), .B1(n3182), .Y(n5442) );
  OA22X1 U10245 ( .A0(\i_MIPS/Register/register[0][5] ), .A1(n3185), .B0(
        \i_MIPS/Register/register[8][5] ), .B1(n3182), .Y(n5433) );
  OA22X1 U10246 ( .A0(\i_MIPS/Register/register[16][5] ), .A1(n3135), .B0(
        \i_MIPS/Register/register[24][5] ), .B1(n3133), .Y(n5421) );
  OA22X1 U10247 ( .A0(\i_MIPS/Register/register[0][5] ), .A1(n3135), .B0(
        \i_MIPS/Register/register[8][5] ), .B1(n3133), .Y(n5412) );
  OA22X1 U10248 ( .A0(\i_MIPS/Register/register[16][7] ), .A1(n2764), .B0(
        \i_MIPS/Register/register[24][7] ), .B1(n2784), .Y(n5029) );
  OA22X1 U10249 ( .A0(\i_MIPS/Register/register[0][7] ), .A1(n2764), .B0(
        \i_MIPS/Register/register[8][7] ), .B1(n3184), .Y(n5020) );
  OA22X1 U10250 ( .A0(\i_MIPS/Register/register[16][7] ), .A1(n3134), .B0(
        \i_MIPS/Register/register[24][7] ), .B1(n3131), .Y(n5008) );
  OA22X1 U10251 ( .A0(\i_MIPS/Register/register[0][7] ), .A1(n3134), .B0(
        \i_MIPS/Register/register[8][7] ), .B1(n3131), .Y(n4999) );
  OA22X1 U10252 ( .A0(\i_MIPS/Register/register[16][6] ), .A1(n3185), .B0(
        \i_MIPS/Register/register[24][6] ), .B1(n3183), .Y(n4959) );
  OA22X1 U10253 ( .A0(\i_MIPS/Register/register[0][6] ), .A1(n3186), .B0(
        \i_MIPS/Register/register[8][6] ), .B1(n3182), .Y(n4950) );
  OA22X1 U10254 ( .A0(\i_MIPS/Register/register[16][6] ), .A1(n3134), .B0(
        \i_MIPS/Register/register[24][6] ), .B1(n3131), .Y(n4938) );
  OA22X1 U10255 ( .A0(\i_MIPS/Register/register[0][6] ), .A1(n3134), .B0(
        \i_MIPS/Register/register[8][6] ), .B1(n3131), .Y(n4929) );
  OA22X1 U10256 ( .A0(\i_MIPS/Register/register[16][2] ), .A1(n3187), .B0(
        \i_MIPS/Register/register[24][2] ), .B1(n3182), .Y(n6663) );
  OA22X1 U10257 ( .A0(\i_MIPS/Register/register[0][2] ), .A1(n3185), .B0(
        \i_MIPS/Register/register[8][2] ), .B1(n3183), .Y(n6654) );
  OA22X1 U10258 ( .A0(\i_MIPS/Register/register[0][16] ), .A1(n3136), .B0(
        \i_MIPS/Register/register[8][16] ), .B1(n2788), .Y(n6956) );
  OA22X1 U10259 ( .A0(\i_MIPS/Register/register[16][15] ), .A1(n3185), .B0(
        \i_MIPS/Register/register[24][15] ), .B1(n3182), .Y(n5592) );
  OA22X1 U10260 ( .A0(\i_MIPS/Register/register[0][15] ), .A1(n3185), .B0(
        \i_MIPS/Register/register[8][15] ), .B1(n3182), .Y(n5583) );
  OA22X1 U10261 ( .A0(\i_MIPS/Register/register[16][15] ), .A1(n3135), .B0(
        \i_MIPS/Register/register[24][15] ), .B1(n2788), .Y(n5571) );
  OA22X1 U10262 ( .A0(\i_MIPS/Register/register[16][16] ), .A1(n3185), .B0(
        \i_MIPS/Register/register[24][16] ), .B1(n2784), .Y(n6944) );
  OA22X1 U10263 ( .A0(\i_MIPS/Register/register[0][16] ), .A1(n3187), .B0(
        \i_MIPS/Register/register[8][16] ), .B1(n3184), .Y(n6935) );
  OA22X1 U10264 ( .A0(\i_MIPS/Register/register[0][23] ), .A1(n3134), .B0(
        \i_MIPS/Register/register[8][23] ), .B1(n3132), .Y(n6887) );
  OA22X1 U10265 ( .A0(\i_MIPS/Register/register[0][17] ), .A1(n2763), .B0(
        \i_MIPS/Register/register[8][17] ), .B1(n3132), .Y(n5695) );
  OA22X1 U10266 ( .A0(\i_MIPS/Register/register[16][1] ), .A1(n2764), .B0(
        \i_MIPS/Register/register[24][1] ), .B1(n3183), .Y(n5171) );
  OA22X1 U10267 ( .A0(\i_MIPS/Register/register[0][1] ), .A1(n3187), .B0(
        \i_MIPS/Register/register[8][1] ), .B1(n3182), .Y(n5162) );
  OA22X1 U10268 ( .A0(\i_MIPS/Register/register[16][1] ), .A1(n3134), .B0(
        \i_MIPS/Register/register[24][1] ), .B1(n3131), .Y(n5150) );
  OA22X1 U10269 ( .A0(\i_MIPS/Register/register[0][1] ), .A1(n3134), .B0(
        \i_MIPS/Register/register[8][1] ), .B1(n3131), .Y(n5141) );
  OA22X1 U10270 ( .A0(n3470), .A1(n526), .B0(n3423), .B1(n1445), .Y(n7403) );
  OA22X1 U10271 ( .A0(n3478), .A1(n527), .B0(n3431), .B1(n1446), .Y(n7770) );
  OA22X1 U10272 ( .A0(n3479), .A1(n528), .B0(n3432), .B1(n1447), .Y(n7774) );
  OA22X1 U10273 ( .A0(n3477), .A1(n529), .B0(n3430), .B1(n1448), .Y(n7725) );
  OA22X1 U10274 ( .A0(n3476), .A1(n530), .B0(n3429), .B1(n1449), .Y(n7697) );
  OA22X1 U10275 ( .A0(n3474), .A1(n531), .B0(n3427), .B1(n1450), .Y(n7620) );
  OA22X1 U10276 ( .A0(n3475), .A1(n532), .B0(n3428), .B1(n1451), .Y(n7624) );
  OA22X1 U10277 ( .A0(n3471), .A1(n533), .B0(n3424), .B1(n1452), .Y(n7512) );
  OA22X1 U10278 ( .A0(\i_MIPS/Register/register[22][8] ), .A1(n3172), .B0(
        \i_MIPS/Register/register[30][8] ), .B1(n3169), .Y(n6175) );
  OA22X1 U10279 ( .A0(\i_MIPS/Register/register[6][8] ), .A1(n3171), .B0(
        \i_MIPS/Register/register[14][8] ), .B1(n3168), .Y(n6166) );
  OA22X1 U10280 ( .A0(\i_MIPS/Register/register[22][11] ), .A1(n3171), .B0(
        \i_MIPS/Register/register[30][11] ), .B1(n3167), .Y(n5306) );
  OA22X1 U10281 ( .A0(\i_MIPS/Register/register[6][11] ), .A1(n3171), .B0(
        \i_MIPS/Register/register[14][11] ), .B1(n3167), .Y(n5297) );
  OA22X1 U10282 ( .A0(\i_MIPS/Register/register[22][9] ), .A1(n3172), .B0(
        \i_MIPS/Register/register[30][9] ), .B1(n3169), .Y(n6244) );
  OA22X1 U10283 ( .A0(\i_MIPS/Register/register[22][23] ), .A1(n3118), .B0(
        \i_MIPS/Register/register[30][23] ), .B1(n3115), .Y(n6890) );
  OA22X1 U10284 ( .A0(\i_MIPS/Register/register[22][17] ), .A1(n3118), .B0(
        \i_MIPS/Register/register[30][17] ), .B1(n3115), .Y(n5698) );
  OA22X1 U10285 ( .A0(\i_MIPS/Register/register[20][8] ), .A1(n3130), .B0(
        \i_MIPS/Register/register[28][8] ), .B1(n3125), .Y(n6161) );
  OA22X1 U10286 ( .A0(\i_MIPS/Register/register[4][8] ), .A1(n3128), .B0(
        \i_MIPS/Register/register[12][8] ), .B1(n3127), .Y(n6152) );
  OA22X1 U10287 ( .A0(\i_MIPS/Register/register[20][9] ), .A1(n3130), .B0(
        \i_MIPS/Register/register[28][9] ), .B1(n3125), .Y(n6230) );
  OA22X1 U10288 ( .A0(\i_MIPS/Register/register[4][9] ), .A1(n3130), .B0(
        \i_MIPS/Register/register[12][9] ), .B1(n3127), .Y(n6221) );
  OA22X1 U10289 ( .A0(\i_MIPS/Register/register[4][9] ), .A1(n2786), .B0(
        \i_MIPS/Register/register[12][9] ), .B1(n3178), .Y(n6242) );
  OA22X1 U10290 ( .A0(\i_MIPS/Register/register[20][13] ), .A1(n3130), .B0(
        \i_MIPS/Register/register[28][13] ), .B1(n3126), .Y(n6428) );
  OA22X1 U10291 ( .A0(\i_MIPS/Register/register[4][13] ), .A1(n3130), .B0(
        \i_MIPS/Register/register[12][13] ), .B1(n3125), .Y(n6419) );
  OA22X1 U10292 ( .A0(\i_MIPS/Register/register[20][14] ), .A1(n3130), .B0(
        \i_MIPS/Register/register[28][14] ), .B1(n3127), .Y(n6362) );
  OA22X1 U10293 ( .A0(\i_MIPS/Register/register[4][14] ), .A1(n3130), .B0(
        \i_MIPS/Register/register[12][14] ), .B1(n3126), .Y(n6353) );
  OA22X1 U10294 ( .A0(\i_MIPS/Register/register[20][11] ), .A1(n3129), .B0(
        \i_MIPS/Register/register[28][11] ), .B1(n3126), .Y(n5292) );
  OA22X1 U10295 ( .A0(\i_MIPS/Register/register[4][11] ), .A1(n3129), .B0(
        \i_MIPS/Register/register[12][11] ), .B1(n3126), .Y(n5283) );
  OA22X1 U10296 ( .A0(\i_MIPS/Register/register[20][10] ), .A1(n3180), .B0(
        \i_MIPS/Register/register[28][10] ), .B1(n3176), .Y(n5248) );
  OA22X1 U10297 ( .A0(\i_MIPS/Register/register[4][10] ), .A1(n3179), .B0(
        \i_MIPS/Register/register[12][10] ), .B1(n3177), .Y(n5239) );
  OA22X1 U10298 ( .A0(\i_MIPS/Register/register[20][10] ), .A1(n3129), .B0(
        \i_MIPS/Register/register[28][10] ), .B1(n3126), .Y(n5227) );
  OA22X1 U10299 ( .A0(\i_MIPS/Register/register[4][10] ), .A1(n3128), .B0(
        \i_MIPS/Register/register[12][10] ), .B1(n3125), .Y(n5218) );
  OA22X1 U10300 ( .A0(\i_MIPS/Register/register[20][5] ), .A1(n3180), .B0(
        \i_MIPS/Register/register[28][5] ), .B1(n3176), .Y(n5443) );
  OA22X1 U10301 ( .A0(\i_MIPS/Register/register[4][5] ), .A1(n3180), .B0(
        \i_MIPS/Register/register[12][5] ), .B1(n3176), .Y(n5434) );
  OA22X1 U10302 ( .A0(\i_MIPS/Register/register[20][5] ), .A1(n3129), .B0(
        \i_MIPS/Register/register[28][5] ), .B1(n3126), .Y(n5422) );
  OA22X1 U10303 ( .A0(\i_MIPS/Register/register[4][5] ), .A1(n3129), .B0(
        \i_MIPS/Register/register[12][5] ), .B1(n3126), .Y(n5413) );
  OA22X1 U10304 ( .A0(\i_MIPS/Register/register[20][7] ), .A1(n3179), .B0(
        \i_MIPS/Register/register[28][7] ), .B1(n2785), .Y(n5030) );
  OA22X1 U10305 ( .A0(\i_MIPS/Register/register[4][7] ), .A1(n3179), .B0(
        \i_MIPS/Register/register[12][7] ), .B1(n2785), .Y(n5021) );
  OA22X1 U10306 ( .A0(\i_MIPS/Register/register[20][7] ), .A1(n3128), .B0(
        \i_MIPS/Register/register[28][7] ), .B1(n3125), .Y(n5009) );
  OA22X1 U10307 ( .A0(\i_MIPS/Register/register[4][7] ), .A1(n3128), .B0(
        \i_MIPS/Register/register[12][7] ), .B1(n3125), .Y(n5000) );
  OA22X1 U10308 ( .A0(\i_MIPS/Register/register[20][6] ), .A1(n3179), .B0(
        \i_MIPS/Register/register[28][6] ), .B1(n3178), .Y(n4960) );
  OA22X1 U10309 ( .A0(\i_MIPS/Register/register[4][6] ), .A1(n3179), .B0(
        \i_MIPS/Register/register[12][6] ), .B1(n3176), .Y(n4951) );
  OA22X1 U10310 ( .A0(\i_MIPS/Register/register[20][6] ), .A1(n3128), .B0(
        \i_MIPS/Register/register[28][6] ), .B1(n3125), .Y(n4939) );
  OA22X1 U10311 ( .A0(\i_MIPS/Register/register[4][6] ), .A1(n3128), .B0(
        \i_MIPS/Register/register[12][6] ), .B1(n3125), .Y(n4930) );
  OA22X1 U10312 ( .A0(\i_MIPS/Register/register[20][2] ), .A1(n3181), .B0(
        \i_MIPS/Register/register[28][2] ), .B1(n3178), .Y(n6664) );
  OA22X1 U10313 ( .A0(\i_MIPS/Register/register[4][2] ), .A1(n3181), .B0(
        \i_MIPS/Register/register[12][2] ), .B1(n3176), .Y(n6655) );
  OA22X1 U10314 ( .A0(\i_MIPS/Register/register[4][16] ), .A1(n3130), .B0(
        \i_MIPS/Register/register[12][16] ), .B1(n2787), .Y(n6957) );
  OA22X1 U10315 ( .A0(\i_MIPS/Register/register[20][15] ), .A1(n3180), .B0(
        \i_MIPS/Register/register[28][15] ), .B1(n3176), .Y(n5593) );
  OA22X1 U10316 ( .A0(\i_MIPS/Register/register[20][15] ), .A1(n3129), .B0(
        \i_MIPS/Register/register[28][15] ), .B1(n3126), .Y(n5572) );
  OA22X1 U10317 ( .A0(\i_MIPS/Register/register[20][16] ), .A1(n3181), .B0(
        \i_MIPS/Register/register[28][16] ), .B1(n3178), .Y(n6945) );
  OA22X1 U10318 ( .A0(\i_MIPS/Register/register[4][23] ), .A1(n3129), .B0(
        \i_MIPS/Register/register[12][23] ), .B1(n3127), .Y(n6888) );
  OA22X1 U10319 ( .A0(\i_MIPS/Register/register[4][17] ), .A1(n3129), .B0(
        \i_MIPS/Register/register[12][17] ), .B1(n3127), .Y(n5696) );
  OA22X1 U10320 ( .A0(\i_MIPS/Register/register[20][1] ), .A1(n3179), .B0(
        \i_MIPS/Register/register[28][1] ), .B1(n2785), .Y(n5172) );
  OA22X1 U10321 ( .A0(\i_MIPS/Register/register[4][1] ), .A1(n3179), .B0(
        \i_MIPS/Register/register[12][1] ), .B1(n3177), .Y(n5163) );
  OA22X1 U10322 ( .A0(\i_MIPS/Register/register[20][1] ), .A1(n3128), .B0(
        \i_MIPS/Register/register[28][1] ), .B1(n3125), .Y(n5151) );
  OA22X1 U10323 ( .A0(\i_MIPS/Register/register[4][1] ), .A1(n3128), .B0(
        \i_MIPS/Register/register[12][1] ), .B1(n3125), .Y(n5142) );
  CLKMX2X2 U10324 ( .A(\I_cache/cache[7][127] ), .B(n8409), .S0(n3497), .Y(
        n9141) );
  CLKMX2X2 U10325 ( .A(\I_cache/cache[6][127] ), .B(n8409), .S0(n3541), .Y(
        n9142) );
  CLKMX2X2 U10326 ( .A(\I_cache/cache[5][127] ), .B(n8409), .S0(n3406), .Y(
        n9143) );
  CLKMX2X2 U10327 ( .A(\I_cache/cache[4][127] ), .B(n8409), .S0(n3452), .Y(
        n9144) );
  CLKMX2X2 U10328 ( .A(\I_cache/cache[3][127] ), .B(n8409), .S0(n3319), .Y(
        n9145) );
  CLKMX2X2 U10329 ( .A(\I_cache/cache[2][127] ), .B(n8409), .S0(n3362), .Y(
        n9146) );
  CLKMX2X2 U10330 ( .A(\I_cache/cache[1][127] ), .B(n8409), .S0(n3229), .Y(
        n9147) );
  CLKMX2X2 U10331 ( .A(\I_cache/cache[0][127] ), .B(n8409), .S0(n3274), .Y(
        n9148) );
  CLKMX2X2 U10332 ( .A(\I_cache/cache[7][126] ), .B(n7275), .S0(n3489), .Y(
        n9149) );
  CLKMX2X2 U10333 ( .A(\I_cache/cache[6][126] ), .B(n7275), .S0(n3533), .Y(
        n9150) );
  CLKMX2X2 U10334 ( .A(\I_cache/cache[5][126] ), .B(n7275), .S0(n3399), .Y(
        n9151) );
  CLKMX2X2 U10335 ( .A(\I_cache/cache[4][126] ), .B(n7275), .S0(n3443), .Y(
        n9152) );
  CLKMX2X2 U10336 ( .A(\I_cache/cache[3][126] ), .B(n7275), .S0(n3311), .Y(
        n9153) );
  CLKMX2X2 U10337 ( .A(\I_cache/cache[2][126] ), .B(n7275), .S0(n3354), .Y(
        n9154) );
  CLKMX2X2 U10338 ( .A(\I_cache/cache[1][126] ), .B(n7275), .S0(n3221), .Y(
        n9155) );
  CLKMX2X2 U10339 ( .A(\I_cache/cache[0][126] ), .B(n7275), .S0(n3266), .Y(
        n9156) );
  CLKMX2X2 U10340 ( .A(\I_cache/cache[7][125] ), .B(n7251), .S0(n3488), .Y(
        n9157) );
  CLKMX2X2 U10341 ( .A(\I_cache/cache[6][125] ), .B(n7251), .S0(n3532), .Y(
        n9158) );
  CLKMX2X2 U10342 ( .A(\I_cache/cache[5][125] ), .B(n7251), .S0(n3398), .Y(
        n9159) );
  CLKMX2X2 U10343 ( .A(\I_cache/cache[4][125] ), .B(n7251), .S0(n3443), .Y(
        n9160) );
  CLKMX2X2 U10344 ( .A(\I_cache/cache[3][125] ), .B(n7251), .S0(n3310), .Y(
        n9161) );
  CLKMX2X2 U10345 ( .A(\I_cache/cache[2][125] ), .B(n7251), .S0(n3353), .Y(
        n9162) );
  CLKMX2X2 U10346 ( .A(\I_cache/cache[1][125] ), .B(n7251), .S0(n3220), .Y(
        n9163) );
  CLKMX2X2 U10347 ( .A(\I_cache/cache[0][125] ), .B(n7251), .S0(n3270), .Y(
        n9164) );
  CLKMX2X2 U10348 ( .A(\I_cache/cache[7][124] ), .B(n7227), .S0(n3488), .Y(
        n9165) );
  CLKMX2X2 U10349 ( .A(\I_cache/cache[6][124] ), .B(n7227), .S0(n3532), .Y(
        n9166) );
  CLKMX2X2 U10350 ( .A(\I_cache/cache[5][124] ), .B(n7227), .S0(n3398), .Y(
        n9167) );
  CLKMX2X2 U10351 ( .A(\I_cache/cache[4][124] ), .B(n7227), .S0(n3443), .Y(
        n9168) );
  CLKMX2X2 U10352 ( .A(\I_cache/cache[3][124] ), .B(n7227), .S0(n3310), .Y(
        n9169) );
  CLKMX2X2 U10353 ( .A(\I_cache/cache[2][124] ), .B(n7227), .S0(n3353), .Y(
        n9170) );
  CLKMX2X2 U10354 ( .A(\I_cache/cache[1][124] ), .B(n7227), .S0(n3220), .Y(
        n9171) );
  CLKMX2X2 U10355 ( .A(\I_cache/cache[0][124] ), .B(n7227), .S0(n3265), .Y(
        n9172) );
  CLKMX2X2 U10356 ( .A(\I_cache/cache[7][123] ), .B(n7203), .S0(n3488), .Y(
        n9173) );
  CLKMX2X2 U10357 ( .A(\I_cache/cache[6][123] ), .B(n7203), .S0(n3532), .Y(
        n9174) );
  CLKMX2X2 U10358 ( .A(\I_cache/cache[5][123] ), .B(n7203), .S0(n3398), .Y(
        n9175) );
  CLKMX2X2 U10359 ( .A(\I_cache/cache[4][123] ), .B(n7203), .S0(n3443), .Y(
        n9176) );
  CLKMX2X2 U10360 ( .A(\I_cache/cache[3][123] ), .B(n7203), .S0(n3310), .Y(
        n9177) );
  CLKMX2X2 U10361 ( .A(\I_cache/cache[2][123] ), .B(n7203), .S0(n3353), .Y(
        n9178) );
  CLKMX2X2 U10362 ( .A(\I_cache/cache[1][123] ), .B(n7203), .S0(n3220), .Y(
        n9179) );
  CLKMX2X2 U10363 ( .A(\I_cache/cache[0][123] ), .B(n7203), .S0(n3265), .Y(
        n9180) );
  CLKMX2X2 U10364 ( .A(\I_cache/cache[7][122] ), .B(n7179), .S0(n3490), .Y(
        n9181) );
  CLKMX2X2 U10365 ( .A(\I_cache/cache[6][122] ), .B(n7179), .S0(n3534), .Y(
        n9182) );
  CLKMX2X2 U10366 ( .A(\I_cache/cache[5][122] ), .B(n7179), .S0(n3400), .Y(
        n9183) );
  CLKMX2X2 U10367 ( .A(\I_cache/cache[4][122] ), .B(n7179), .S0(n3444), .Y(
        n9184) );
  CLKMX2X2 U10368 ( .A(\I_cache/cache[3][122] ), .B(n7179), .S0(n3312), .Y(
        n9185) );
  CLKMX2X2 U10369 ( .A(\I_cache/cache[2][122] ), .B(n7179), .S0(n3355), .Y(
        n9186) );
  CLKMX2X2 U10370 ( .A(\I_cache/cache[1][122] ), .B(n7179), .S0(n3222), .Y(
        n9187) );
  CLKMX2X2 U10371 ( .A(\I_cache/cache[0][122] ), .B(n7179), .S0(n3265), .Y(
        n9188) );
  CLKMX2X2 U10372 ( .A(\I_cache/cache[7][121] ), .B(n7651), .S0(n3493), .Y(
        n9189) );
  CLKMX2X2 U10373 ( .A(\I_cache/cache[6][121] ), .B(n7651), .S0(n3536), .Y(
        n9190) );
  CLKMX2X2 U10374 ( .A(\I_cache/cache[5][121] ), .B(n7651), .S0(n3401), .Y(
        n9191) );
  CLKMX2X2 U10375 ( .A(\I_cache/cache[4][121] ), .B(n7651), .S0(n3446), .Y(
        n9192) );
  CLKMX2X2 U10376 ( .A(\I_cache/cache[3][121] ), .B(n7651), .S0(n3310), .Y(
        n9193) );
  CLKMX2X2 U10377 ( .A(\I_cache/cache[2][121] ), .B(n7651), .S0(n3353), .Y(
        n9194) );
  CLKMX2X2 U10378 ( .A(\I_cache/cache[1][121] ), .B(n7651), .S0(n3220), .Y(
        n9195) );
  CLKMX2X2 U10379 ( .A(\I_cache/cache[0][121] ), .B(n7651), .S0(n3269), .Y(
        n9196) );
  CLKMX2X2 U10380 ( .A(\I_cache/cache[7][120] ), .B(n7429), .S0(n3489), .Y(
        n9197) );
  CLKMX2X2 U10381 ( .A(\I_cache/cache[6][120] ), .B(n7429), .S0(n3533), .Y(
        n9198) );
  CLKMX2X2 U10382 ( .A(\I_cache/cache[5][120] ), .B(n7429), .S0(n3399), .Y(
        n9199) );
  CLKMX2X2 U10383 ( .A(\I_cache/cache[4][120] ), .B(n7429), .S0(n3448), .Y(
        n9200) );
  CLKMX2X2 U10384 ( .A(\I_cache/cache[3][120] ), .B(n7429), .S0(n3311), .Y(
        n9201) );
  CLKMX2X2 U10385 ( .A(\I_cache/cache[2][120] ), .B(n7429), .S0(n3354), .Y(
        n9202) );
  CLKMX2X2 U10386 ( .A(\I_cache/cache[1][120] ), .B(n7429), .S0(n3221), .Y(
        n9203) );
  CLKMX2X2 U10387 ( .A(\I_cache/cache[0][120] ), .B(n7429), .S0(n3266), .Y(
        n9204) );
  CLKMX2X2 U10388 ( .A(\I_cache/cache[7][119] ), .B(n7453), .S0(n3493), .Y(
        n9205) );
  CLKMX2X2 U10389 ( .A(\I_cache/cache[6][119] ), .B(n7453), .S0(n3538), .Y(
        n9206) );
  CLKMX2X2 U10390 ( .A(\I_cache/cache[5][119] ), .B(n7453), .S0(n3403), .Y(
        n9207) );
  CLKMX2X2 U10391 ( .A(\I_cache/cache[4][119] ), .B(n7453), .S0(n3448), .Y(
        n9208) );
  CLKMX2X2 U10392 ( .A(\I_cache/cache[3][119] ), .B(n7453), .S0(n3315), .Y(
        n9209) );
  CLKMX2X2 U10393 ( .A(\I_cache/cache[2][119] ), .B(n7453), .S0(n3358), .Y(
        n9210) );
  CLKMX2X2 U10394 ( .A(\I_cache/cache[1][119] ), .B(n7453), .S0(n3225), .Y(
        n9211) );
  CLKMX2X2 U10395 ( .A(\I_cache/cache[0][119] ), .B(n7453), .S0(n3271), .Y(
        n9212) );
  CLKMX2X2 U10396 ( .A(\I_cache/cache[7][118] ), .B(n8113), .S0(n3497), .Y(
        n9213) );
  CLKMX2X2 U10397 ( .A(\I_cache/cache[6][118] ), .B(n8113), .S0(n3541), .Y(
        n9214) );
  CLKMX2X2 U10398 ( .A(\I_cache/cache[5][118] ), .B(n8113), .S0(n3406), .Y(
        n9215) );
  CLKMX2X2 U10399 ( .A(\I_cache/cache[4][118] ), .B(n8113), .S0(n3452), .Y(
        n9216) );
  CLKMX2X2 U10400 ( .A(\I_cache/cache[3][118] ), .B(n8113), .S0(n3319), .Y(
        n9217) );
  CLKMX2X2 U10401 ( .A(\I_cache/cache[2][118] ), .B(n8113), .S0(n3362), .Y(
        n9218) );
  CLKMX2X2 U10402 ( .A(\I_cache/cache[1][118] ), .B(n8113), .S0(n3229), .Y(
        n9219) );
  CLKMX2X2 U10403 ( .A(\I_cache/cache[0][118] ), .B(n8113), .S0(n3274), .Y(
        n9220) );
  CLKMX2X2 U10404 ( .A(\I_cache/cache[7][117] ), .B(n7477), .S0(n3493), .Y(
        n9221) );
  CLKMX2X2 U10405 ( .A(\I_cache/cache[6][117] ), .B(n7477), .S0(n3538), .Y(
        n9222) );
  CLKMX2X2 U10406 ( .A(\I_cache/cache[5][117] ), .B(n7477), .S0(n3403), .Y(
        n9223) );
  CLKMX2X2 U10407 ( .A(\I_cache/cache[4][117] ), .B(n7477), .S0(n3448), .Y(
        n9224) );
  CLKMX2X2 U10408 ( .A(\I_cache/cache[3][117] ), .B(n7477), .S0(n3315), .Y(
        n9225) );
  CLKMX2X2 U10409 ( .A(\I_cache/cache[2][117] ), .B(n7477), .S0(n3358), .Y(
        n9226) );
  CLKMX2X2 U10410 ( .A(\I_cache/cache[1][117] ), .B(n7477), .S0(n3225), .Y(
        n9227) );
  CLKMX2X2 U10411 ( .A(\I_cache/cache[0][117] ), .B(n7477), .S0(n3271), .Y(
        n9228) );
  CLKMX2X2 U10412 ( .A(\I_cache/cache[7][116] ), .B(n7501), .S0(n3493), .Y(
        n9229) );
  CLKMX2X2 U10413 ( .A(\I_cache/cache[6][116] ), .B(n7501), .S0(n3538), .Y(
        n9230) );
  CLKMX2X2 U10414 ( .A(\I_cache/cache[5][116] ), .B(n7501), .S0(n3403), .Y(
        n9231) );
  CLKMX2X2 U10415 ( .A(\I_cache/cache[4][116] ), .B(n7501), .S0(n3448), .Y(
        n9232) );
  CLKMX2X2 U10416 ( .A(\I_cache/cache[3][116] ), .B(n7501), .S0(n3315), .Y(
        n9233) );
  CLKMX2X2 U10417 ( .A(\I_cache/cache[2][116] ), .B(n7501), .S0(n3358), .Y(
        n9234) );
  CLKMX2X2 U10418 ( .A(\I_cache/cache[1][116] ), .B(n7501), .S0(n3225), .Y(
        n9235) );
  CLKMX2X2 U10419 ( .A(\I_cache/cache[0][116] ), .B(n7501), .S0(n3271), .Y(
        n9236) );
  CLKMX2X2 U10420 ( .A(\I_cache/cache[7][115] ), .B(n7130), .S0(n3491), .Y(
        n9237) );
  CLKMX2X2 U10421 ( .A(\I_cache/cache[6][115] ), .B(n7130), .S0(n3535), .Y(
        n9238) );
  CLKMX2X2 U10422 ( .A(\I_cache/cache[5][115] ), .B(n7130), .S0(n3406), .Y(
        n9239) );
  CLKMX2X2 U10423 ( .A(\I_cache/cache[4][115] ), .B(n7130), .S0(n3445), .Y(
        n9240) );
  CLKMX2X2 U10424 ( .A(\I_cache/cache[3][115] ), .B(n7130), .S0(n3313), .Y(
        n9241) );
  CLKMX2X2 U10425 ( .A(\I_cache/cache[2][115] ), .B(n7130), .S0(n3356), .Y(
        n9242) );
  CLKMX2X2 U10426 ( .A(\I_cache/cache[1][115] ), .B(n7130), .S0(n3223), .Y(
        n9243) );
  CLKMX2X2 U10427 ( .A(\I_cache/cache[0][115] ), .B(n7130), .S0(n3268), .Y(
        n9244) );
  CLKMX2X2 U10428 ( .A(\I_cache/cache[7][114] ), .B(n7154), .S0(n3491), .Y(
        n9245) );
  CLKMX2X2 U10429 ( .A(\I_cache/cache[6][114] ), .B(n7154), .S0(n3535), .Y(
        n9246) );
  CLKMX2X2 U10430 ( .A(\I_cache/cache[5][114] ), .B(n7154), .S0(n3400), .Y(
        n9247) );
  CLKMX2X2 U10431 ( .A(\I_cache/cache[4][114] ), .B(n7154), .S0(n3445), .Y(
        n9248) );
  CLKMX2X2 U10432 ( .A(\I_cache/cache[3][114] ), .B(n7154), .S0(n3313), .Y(
        n9249) );
  CLKMX2X2 U10433 ( .A(\I_cache/cache[2][114] ), .B(n7154), .S0(n3356), .Y(
        n9250) );
  CLKMX2X2 U10434 ( .A(\I_cache/cache[1][114] ), .B(n7154), .S0(n3223), .Y(
        n9251) );
  CLKMX2X2 U10435 ( .A(\I_cache/cache[0][114] ), .B(n7154), .S0(n3268), .Y(
        n9252) );
  CLKMX2X2 U10436 ( .A(\I_cache/cache[7][113] ), .B(n4583), .S0(n3490), .Y(
        n9253) );
  CLKMX2X2 U10437 ( .A(\I_cache/cache[6][113] ), .B(n4583), .S0(n3534), .Y(
        n9254) );
  CLKMX2X2 U10438 ( .A(\I_cache/cache[5][113] ), .B(n4583), .S0(n3400), .Y(
        n9255) );
  CLKMX2X2 U10439 ( .A(\I_cache/cache[4][113] ), .B(n4583), .S0(n3444), .Y(
        n9256) );
  CLKMX2X2 U10440 ( .A(\I_cache/cache[3][113] ), .B(n4583), .S0(n3312), .Y(
        n9257) );
  CLKMX2X2 U10441 ( .A(\I_cache/cache[2][113] ), .B(n4583), .S0(n3355), .Y(
        n9258) );
  CLKMX2X2 U10442 ( .A(\I_cache/cache[1][113] ), .B(n4583), .S0(n3222), .Y(
        n9259) );
  CLKMX2X2 U10443 ( .A(\I_cache/cache[0][113] ), .B(n4583), .S0(n3267), .Y(
        n9260) );
  CLKMX2X2 U10444 ( .A(\I_cache/cache[7][112] ), .B(n7106), .S0(n3491), .Y(
        n9261) );
  CLKMX2X2 U10445 ( .A(\I_cache/cache[6][112] ), .B(n7106), .S0(n3535), .Y(
        n9262) );
  CLKMX2X2 U10446 ( .A(\I_cache/cache[5][112] ), .B(n7106), .S0(n3406), .Y(
        n9263) );
  CLKMX2X2 U10447 ( .A(\I_cache/cache[4][112] ), .B(n7106), .S0(n3445), .Y(
        n9264) );
  CLKMX2X2 U10448 ( .A(\I_cache/cache[3][112] ), .B(n7106), .S0(n3313), .Y(
        n9265) );
  CLKMX2X2 U10449 ( .A(\I_cache/cache[2][112] ), .B(n7106), .S0(n3356), .Y(
        n9266) );
  CLKMX2X2 U10450 ( .A(\I_cache/cache[1][112] ), .B(n7106), .S0(n3222), .Y(
        n9267) );
  CLKMX2X2 U10451 ( .A(\I_cache/cache[0][112] ), .B(n7106), .S0(n3268), .Y(
        n9268) );
  CLKMX2X2 U10452 ( .A(\I_cache/cache[7][111] ), .B(n7549), .S0(n3494), .Y(
        n9269) );
  CLKMX2X2 U10453 ( .A(\I_cache/cache[6][111] ), .B(n7549), .S0(n3539), .Y(
        n9270) );
  CLKMX2X2 U10454 ( .A(\I_cache/cache[5][111] ), .B(n7549), .S0(n3404), .Y(
        n9271) );
  CLKMX2X2 U10455 ( .A(\I_cache/cache[4][111] ), .B(n7549), .S0(n3449), .Y(
        n9272) );
  CLKMX2X2 U10456 ( .A(\I_cache/cache[3][111] ), .B(n7549), .S0(n3316), .Y(
        n9273) );
  CLKMX2X2 U10457 ( .A(\I_cache/cache[2][111] ), .B(n7549), .S0(n3359), .Y(
        n9274) );
  CLKMX2X2 U10458 ( .A(\I_cache/cache[1][111] ), .B(n7549), .S0(n3226), .Y(
        n9275) );
  CLKMX2X2 U10459 ( .A(\I_cache/cache[0][111] ), .B(n7549), .S0(n3272), .Y(
        n9276) );
  CLKMX2X2 U10460 ( .A(\I_cache/cache[7][110] ), .B(n7525), .S0(n3492), .Y(
        n9277) );
  CLKMX2X2 U10461 ( .A(\I_cache/cache[6][110] ), .B(n7525), .S0(n3537), .Y(
        n9278) );
  CLKMX2X2 U10462 ( .A(\I_cache/cache[5][110] ), .B(n7525), .S0(n3402), .Y(
        n9279) );
  CLKMX2X2 U10463 ( .A(\I_cache/cache[4][110] ), .B(n7525), .S0(n3447), .Y(
        n9280) );
  CLKMX2X2 U10464 ( .A(\I_cache/cache[3][110] ), .B(n7525), .S0(n3314), .Y(
        n9281) );
  CLKMX2X2 U10465 ( .A(\I_cache/cache[2][110] ), .B(n7525), .S0(n3357), .Y(
        n9282) );
  CLKMX2X2 U10466 ( .A(\I_cache/cache[1][110] ), .B(n7525), .S0(n3226), .Y(
        n9283) );
  CLKMX2X2 U10467 ( .A(\I_cache/cache[0][110] ), .B(n7525), .S0(n3272), .Y(
        n9284) );
  CLKMX2X2 U10468 ( .A(\I_cache/cache[7][109] ), .B(n7574), .S0(n3494), .Y(
        n9285) );
  CLKMX2X2 U10469 ( .A(\I_cache/cache[6][109] ), .B(n7574), .S0(n3539), .Y(
        n9286) );
  CLKMX2X2 U10470 ( .A(\I_cache/cache[5][109] ), .B(n7574), .S0(n3404), .Y(
        n9287) );
  CLKMX2X2 U10471 ( .A(\I_cache/cache[4][109] ), .B(n7574), .S0(n3449), .Y(
        n9288) );
  CLKMX2X2 U10472 ( .A(\I_cache/cache[3][109] ), .B(n7574), .S0(n3316), .Y(
        n9289) );
  CLKMX2X2 U10473 ( .A(\I_cache/cache[2][109] ), .B(n7574), .S0(n3359), .Y(
        n9290) );
  CLKMX2X2 U10474 ( .A(\I_cache/cache[1][109] ), .B(n7574), .S0(n3226), .Y(
        n9291) );
  CLKMX2X2 U10475 ( .A(\I_cache/cache[0][109] ), .B(n7574), .S0(n3272), .Y(
        n9292) );
  CLKMX2X2 U10476 ( .A(\I_cache/cache[7][108] ), .B(n7622), .S0(n3492), .Y(
        n9293) );
  CLKMX2X2 U10477 ( .A(\I_cache/cache[6][108] ), .B(n7622), .S0(n3536), .Y(
        n9294) );
  CLKMX2X2 U10478 ( .A(\I_cache/cache[5][108] ), .B(n7622), .S0(n3401), .Y(
        n9295) );
  CLKMX2X2 U10479 ( .A(\I_cache/cache[4][108] ), .B(n7622), .S0(n3446), .Y(
        n9296) );
  CLKMX2X2 U10480 ( .A(\I_cache/cache[3][108] ), .B(n7622), .S0(n3311), .Y(
        n9297) );
  CLKMX2X2 U10481 ( .A(\I_cache/cache[2][108] ), .B(n7622), .S0(n3354), .Y(
        n9298) );
  CLKMX2X2 U10482 ( .A(\I_cache/cache[1][108] ), .B(n7622), .S0(n3221), .Y(
        n9299) );
  CLKMX2X2 U10483 ( .A(\I_cache/cache[0][108] ), .B(n7622), .S0(n3269), .Y(
        n9300) );
  CLKMX2X2 U10484 ( .A(\I_cache/cache[7][107] ), .B(n7598), .S0(n3494), .Y(
        n9301) );
  CLKMX2X2 U10485 ( .A(\I_cache/cache[6][107] ), .B(n7598), .S0(n3539), .Y(
        n9302) );
  CLKMX2X2 U10486 ( .A(\I_cache/cache[5][107] ), .B(n7598), .S0(n3404), .Y(
        n9303) );
  CLKMX2X2 U10487 ( .A(\I_cache/cache[4][107] ), .B(n7598), .S0(n3449), .Y(
        n9304) );
  CLKMX2X2 U10488 ( .A(\I_cache/cache[3][107] ), .B(n7598), .S0(n3316), .Y(
        n9305) );
  CLKMX2X2 U10489 ( .A(\I_cache/cache[2][107] ), .B(n7598), .S0(n3359), .Y(
        n9306) );
  CLKMX2X2 U10490 ( .A(\I_cache/cache[1][107] ), .B(n7598), .S0(n3225), .Y(
        n9307) );
  CLKMX2X2 U10491 ( .A(\I_cache/cache[0][107] ), .B(n7598), .S0(n3269), .Y(
        n9308) );
  CLKMX2X2 U10492 ( .A(\I_cache/cache[7][106] ), .B(n7676), .S0(n3491), .Y(
        n9309) );
  CLKMX2X2 U10493 ( .A(\I_cache/cache[6][106] ), .B(n7676), .S0(n3535), .Y(
        n9310) );
  CLKMX2X2 U10494 ( .A(\I_cache/cache[5][106] ), .B(n7676), .S0(n3400), .Y(
        n9311) );
  CLKMX2X2 U10495 ( .A(\I_cache/cache[4][106] ), .B(n7676), .S0(n3445), .Y(
        n9312) );
  CLKMX2X2 U10496 ( .A(\I_cache/cache[3][106] ), .B(n7676), .S0(n3313), .Y(
        n9313) );
  CLKMX2X2 U10497 ( .A(\I_cache/cache[2][106] ), .B(n7676), .S0(n3356), .Y(
        n9314) );
  CLKMX2X2 U10498 ( .A(\I_cache/cache[1][106] ), .B(n7676), .S0(n3223), .Y(
        n9315) );
  CLKMX2X2 U10499 ( .A(\I_cache/cache[0][106] ), .B(n7676), .S0(n3268), .Y(
        n9316) );
  CLKMX2X2 U10500 ( .A(\I_cache/cache[7][105] ), .B(n7699), .S0(n3492), .Y(
        n9317) );
  CLKMX2X2 U10501 ( .A(\I_cache/cache[6][105] ), .B(n7699), .S0(n3537), .Y(
        n9318) );
  CLKMX2X2 U10502 ( .A(\I_cache/cache[5][105] ), .B(n7699), .S0(n3402), .Y(
        n9319) );
  CLKMX2X2 U10503 ( .A(\I_cache/cache[4][105] ), .B(n7699), .S0(n3447), .Y(
        n9320) );
  CLKMX2X2 U10504 ( .A(\I_cache/cache[3][105] ), .B(n7699), .S0(n3314), .Y(
        n9321) );
  CLKMX2X2 U10505 ( .A(\I_cache/cache[2][105] ), .B(n7699), .S0(n3357), .Y(
        n9322) );
  CLKMX2X2 U10506 ( .A(\I_cache/cache[1][105] ), .B(n7699), .S0(n3224), .Y(
        n9323) );
  CLKMX2X2 U10507 ( .A(\I_cache/cache[0][105] ), .B(n7699), .S0(n3270), .Y(
        n9324) );
  CLKMX2X2 U10508 ( .A(\I_cache/cache[7][104] ), .B(n7723), .S0(n3492), .Y(
        n9325) );
  CLKMX2X2 U10509 ( .A(\I_cache/cache[6][104] ), .B(n7723), .S0(n3537), .Y(
        n9326) );
  CLKMX2X2 U10510 ( .A(\I_cache/cache[5][104] ), .B(n7723), .S0(n3402), .Y(
        n9327) );
  CLKMX2X2 U10511 ( .A(\I_cache/cache[4][104] ), .B(n7723), .S0(n3447), .Y(
        n9328) );
  CLKMX2X2 U10512 ( .A(\I_cache/cache[3][104] ), .B(n7723), .S0(n3314), .Y(
        n9329) );
  CLKMX2X2 U10513 ( .A(\I_cache/cache[2][104] ), .B(n7723), .S0(n3357), .Y(
        n9330) );
  CLKMX2X2 U10514 ( .A(\I_cache/cache[1][104] ), .B(n7723), .S0(n3224), .Y(
        n9331) );
  CLKMX2X2 U10515 ( .A(\I_cache/cache[0][104] ), .B(n7723), .S0(n3270), .Y(
        n9332) );
  CLKMX2X2 U10516 ( .A(\I_cache/cache[7][103] ), .B(n7749), .S0(n3492), .Y(
        n9333) );
  CLKMX2X2 U10517 ( .A(\I_cache/cache[6][103] ), .B(n7749), .S0(n3537), .Y(
        n9334) );
  CLKMX2X2 U10518 ( .A(\I_cache/cache[5][103] ), .B(n7749), .S0(n3402), .Y(
        n9335) );
  CLKMX2X2 U10519 ( .A(\I_cache/cache[4][103] ), .B(n7749), .S0(n3447), .Y(
        n9336) );
  CLKMX2X2 U10520 ( .A(\I_cache/cache[3][103] ), .B(n7749), .S0(n3314), .Y(
        n9337) );
  CLKMX2X2 U10521 ( .A(\I_cache/cache[2][103] ), .B(n7749), .S0(n3357), .Y(
        n9338) );
  CLKMX2X2 U10522 ( .A(\I_cache/cache[1][103] ), .B(n7749), .S0(n3222), .Y(
        n9339) );
  CLKMX2X2 U10523 ( .A(\I_cache/cache[0][103] ), .B(n7749), .S0(n3269), .Y(
        n9340) );
  CLKMX2X2 U10524 ( .A(\I_cache/cache[7][102] ), .B(n7772), .S0(n3497), .Y(
        n9341) );
  CLKMX2X2 U10525 ( .A(\I_cache/cache[6][102] ), .B(n7772), .S0(n3541), .Y(
        n9342) );
  CLKMX2X2 U10526 ( .A(\I_cache/cache[5][102] ), .B(n7772), .S0(n3406), .Y(
        n9343) );
  CLKMX2X2 U10527 ( .A(\I_cache/cache[4][102] ), .B(n7772), .S0(n3452), .Y(
        n9344) );
  CLKMX2X2 U10528 ( .A(\I_cache/cache[3][102] ), .B(n7772), .S0(n3319), .Y(
        n9345) );
  CLKMX2X2 U10529 ( .A(\I_cache/cache[2][102] ), .B(n7772), .S0(n3362), .Y(
        n9346) );
  CLKMX2X2 U10530 ( .A(\I_cache/cache[1][102] ), .B(n7772), .S0(n3229), .Y(
        n9347) );
  CLKMX2X2 U10531 ( .A(\I_cache/cache[0][102] ), .B(n7772), .S0(n3274), .Y(
        n9348) );
  CLKMX2X2 U10532 ( .A(\I_cache/cache[7][101] ), .B(n7401), .S0(n3489), .Y(
        n9349) );
  CLKMX2X2 U10533 ( .A(\I_cache/cache[6][101] ), .B(n7401), .S0(n3533), .Y(
        n9350) );
  CLKMX2X2 U10534 ( .A(\I_cache/cache[5][101] ), .B(n7401), .S0(n3399), .Y(
        n9351) );
  CLKMX2X2 U10535 ( .A(\I_cache/cache[4][101] ), .B(n7401), .S0(n3447), .Y(
        n9352) );
  CLKMX2X2 U10536 ( .A(\I_cache/cache[3][101] ), .B(n7401), .S0(n3311), .Y(
        n9353) );
  CLKMX2X2 U10537 ( .A(\I_cache/cache[2][101] ), .B(n7401), .S0(n3354), .Y(
        n9354) );
  CLKMX2X2 U10538 ( .A(\I_cache/cache[1][101] ), .B(n7401), .S0(n3221), .Y(
        n9355) );
  CLKMX2X2 U10539 ( .A(\I_cache/cache[0][101] ), .B(n7401), .S0(n3266), .Y(
        n9356) );
  CLKMX2X2 U10540 ( .A(\I_cache/cache[7][100] ), .B(n8346), .S0(n3497), .Y(
        n9357) );
  CLKMX2X2 U10541 ( .A(\I_cache/cache[6][100] ), .B(n8346), .S0(n3541), .Y(
        n9358) );
  CLKMX2X2 U10542 ( .A(\I_cache/cache[5][100] ), .B(n8346), .S0(n3406), .Y(
        n9359) );
  CLKMX2X2 U10543 ( .A(\I_cache/cache[4][100] ), .B(n8346), .S0(n3452), .Y(
        n9360) );
  CLKMX2X2 U10544 ( .A(\I_cache/cache[3][100] ), .B(n8346), .S0(n3319), .Y(
        n9361) );
  CLKMX2X2 U10545 ( .A(\I_cache/cache[2][100] ), .B(n8346), .S0(n3362), .Y(
        n9362) );
  CLKMX2X2 U10546 ( .A(\I_cache/cache[1][100] ), .B(n8346), .S0(n3229), .Y(
        n9363) );
  CLKMX2X2 U10547 ( .A(\I_cache/cache[0][100] ), .B(n8346), .S0(n3274), .Y(
        n9364) );
  CLKMX2X2 U10548 ( .A(\I_cache/cache[7][99] ), .B(n8365), .S0(n3496), .Y(
        n9365) );
  CLKMX2X2 U10549 ( .A(\I_cache/cache[6][99] ), .B(n8365), .S0(n3540), .Y(
        n9366) );
  CLKMX2X2 U10550 ( .A(\I_cache/cache[5][99] ), .B(n8365), .S0(n3405), .Y(
        n9367) );
  CLKMX2X2 U10551 ( .A(\I_cache/cache[4][99] ), .B(n8365), .S0(n3451), .Y(
        n9368) );
  CLKMX2X2 U10552 ( .A(\I_cache/cache[3][99] ), .B(n8365), .S0(n3318), .Y(
        n9369) );
  CLKMX2X2 U10553 ( .A(\I_cache/cache[2][99] ), .B(n8365), .S0(n3361), .Y(
        n9370) );
  CLKMX2X2 U10554 ( .A(\I_cache/cache[1][99] ), .B(n8365), .S0(n3228), .Y(
        n9371) );
  CLKMX2X2 U10555 ( .A(\I_cache/cache[0][99] ), .B(n8365), .S0(n3273), .Y(
        n9372) );
  CLKMX2X2 U10556 ( .A(\I_cache/cache[7][98] ), .B(n8379), .S0(n3491), .Y(
        n9373) );
  CLKMX2X2 U10557 ( .A(\I_cache/cache[6][98] ), .B(n8379), .S0(n3538), .Y(
        n9374) );
  CLKMX2X2 U10558 ( .A(\I_cache/cache[5][98] ), .B(n8379), .S0(n3407), .Y(
        n9375) );
  CLKMX2X2 U10559 ( .A(\I_cache/cache[4][98] ), .B(n8379), .S0(n3444), .Y(
        n9376) );
  CLKMX2X2 U10560 ( .A(\I_cache/cache[3][98] ), .B(n8379), .S0(n3319), .Y(
        n9377) );
  CLKMX2X2 U10561 ( .A(\I_cache/cache[2][98] ), .B(n8379), .S0(n3362), .Y(
        n9378) );
  CLKMX2X2 U10562 ( .A(\I_cache/cache[1][98] ), .B(n8379), .S0(n3229), .Y(
        n9379) );
  CLKMX2X2 U10563 ( .A(\I_cache/cache[0][98] ), .B(n8379), .S0(n3274), .Y(
        n9380) );
  CLKMX2X2 U10564 ( .A(\I_cache/cache[7][97] ), .B(n4563), .S0(n3490), .Y(
        n9381) );
  CLKMX2X2 U10565 ( .A(\I_cache/cache[6][97] ), .B(n4563), .S0(n3534), .Y(
        n9382) );
  CLKMX2X2 U10566 ( .A(\I_cache/cache[5][97] ), .B(n4563), .S0(n3400), .Y(
        n9383) );
  CLKMX2X2 U10567 ( .A(\I_cache/cache[4][97] ), .B(n4563), .S0(n3444), .Y(
        n9384) );
  CLKMX2X2 U10568 ( .A(\I_cache/cache[3][97] ), .B(n4563), .S0(n3312), .Y(
        n9385) );
  CLKMX2X2 U10569 ( .A(\I_cache/cache[2][97] ), .B(n4563), .S0(n3355), .Y(
        n9386) );
  CLKMX2X2 U10570 ( .A(\I_cache/cache[1][97] ), .B(n4563), .S0(n3222), .Y(
        n9387) );
  CLKMX2X2 U10571 ( .A(\I_cache/cache[0][97] ), .B(n4563), .S0(n3267), .Y(
        n9388) );
  CLKMX2X2 U10572 ( .A(\I_cache/cache[7][95] ), .B(n8411), .S0(n3495), .Y(
        n9397) );
  CLKMX2X2 U10573 ( .A(\I_cache/cache[6][95] ), .B(n8411), .S0(n3538), .Y(
        n9398) );
  CLKMX2X2 U10574 ( .A(\I_cache/cache[5][95] ), .B(n8411), .S0(n3406), .Y(
        n9399) );
  CLKMX2X2 U10575 ( .A(\I_cache/cache[4][95] ), .B(n8411), .S0(n3450), .Y(
        n9400) );
  CLKMX2X2 U10576 ( .A(\I_cache/cache[3][95] ), .B(n8411), .S0(n3317), .Y(
        n9401) );
  CLKMX2X2 U10577 ( .A(\I_cache/cache[2][95] ), .B(n8411), .S0(n3360), .Y(
        n9402) );
  CLKMX2X2 U10578 ( .A(\I_cache/cache[1][95] ), .B(n8411), .S0(n3227), .Y(
        n9403) );
  CLKMX2X2 U10579 ( .A(\I_cache/cache[0][95] ), .B(n8411), .S0(n3274), .Y(
        n9404) );
  CLKMX2X2 U10580 ( .A(\I_cache/cache[7][94] ), .B(n7280), .S0(n3489), .Y(
        n9405) );
  CLKMX2X2 U10581 ( .A(\I_cache/cache[6][94] ), .B(n7280), .S0(n3533), .Y(
        n9406) );
  CLKMX2X2 U10582 ( .A(\I_cache/cache[5][94] ), .B(n7280), .S0(n3399), .Y(
        n9407) );
  CLKMX2X2 U10583 ( .A(\I_cache/cache[4][94] ), .B(n7280), .S0(n3443), .Y(
        n9408) );
  CLKMX2X2 U10584 ( .A(\I_cache/cache[3][94] ), .B(n7280), .S0(n3311), .Y(
        n9409) );
  CLKMX2X2 U10585 ( .A(\I_cache/cache[2][94] ), .B(n7280), .S0(n3354), .Y(
        n9410) );
  CLKMX2X2 U10586 ( .A(\I_cache/cache[1][94] ), .B(n7280), .S0(n3221), .Y(
        n9411) );
  CLKMX2X2 U10587 ( .A(\I_cache/cache[0][94] ), .B(n7280), .S0(n3266), .Y(
        n9412) );
  CLKMX2X2 U10588 ( .A(\I_cache/cache[7][93] ), .B(n7256), .S0(n3488), .Y(
        n9413) );
  CLKMX2X2 U10589 ( .A(\I_cache/cache[6][93] ), .B(n7256), .S0(n3532), .Y(
        n9414) );
  CLKMX2X2 U10590 ( .A(\I_cache/cache[5][93] ), .B(n7256), .S0(n3398), .Y(
        n9415) );
  CLKMX2X2 U10591 ( .A(\I_cache/cache[4][93] ), .B(n7256), .S0(n3443), .Y(
        n9416) );
  CLKMX2X2 U10592 ( .A(\I_cache/cache[3][93] ), .B(n7256), .S0(n3310), .Y(
        n9417) );
  CLKMX2X2 U10593 ( .A(\I_cache/cache[2][93] ), .B(n7256), .S0(n3353), .Y(
        n9418) );
  CLKMX2X2 U10594 ( .A(\I_cache/cache[1][93] ), .B(n7256), .S0(n3221), .Y(
        n9419) );
  CLKMX2X2 U10595 ( .A(\I_cache/cache[0][93] ), .B(n7256), .S0(n3266), .Y(
        n9420) );
  CLKMX2X2 U10596 ( .A(\I_cache/cache[7][92] ), .B(n7232), .S0(n3488), .Y(
        n9421) );
  CLKMX2X2 U10597 ( .A(\I_cache/cache[6][92] ), .B(n7232), .S0(n3532), .Y(
        n9422) );
  CLKMX2X2 U10598 ( .A(\I_cache/cache[5][92] ), .B(n7232), .S0(n3398), .Y(
        n9423) );
  CLKMX2X2 U10599 ( .A(\I_cache/cache[4][92] ), .B(n7232), .S0(n3443), .Y(
        n9424) );
  CLKMX2X2 U10600 ( .A(\I_cache/cache[3][92] ), .B(n7232), .S0(n3310), .Y(
        n9425) );
  CLKMX2X2 U10601 ( .A(\I_cache/cache[2][92] ), .B(n7232), .S0(n3353), .Y(
        n9426) );
  CLKMX2X2 U10602 ( .A(\I_cache/cache[1][92] ), .B(n7232), .S0(n3220), .Y(
        n9427) );
  CLKMX2X2 U10603 ( .A(\I_cache/cache[0][92] ), .B(n7232), .S0(n3265), .Y(
        n9428) );
  CLKMX2X2 U10604 ( .A(\I_cache/cache[7][91] ), .B(n7208), .S0(n3488), .Y(
        n9429) );
  CLKMX2X2 U10605 ( .A(\I_cache/cache[6][91] ), .B(n7208), .S0(n3532), .Y(
        n9430) );
  CLKMX2X2 U10606 ( .A(\I_cache/cache[5][91] ), .B(n7208), .S0(n3398), .Y(
        n9431) );
  CLKMX2X2 U10607 ( .A(\I_cache/cache[4][91] ), .B(n7208), .S0(n3443), .Y(
        n9432) );
  CLKMX2X2 U10608 ( .A(\I_cache/cache[3][91] ), .B(n7208), .S0(n3310), .Y(
        n9433) );
  CLKMX2X2 U10609 ( .A(\I_cache/cache[2][91] ), .B(n7208), .S0(n3353), .Y(
        n9434) );
  CLKMX2X2 U10610 ( .A(\I_cache/cache[1][91] ), .B(n7208), .S0(n3220), .Y(
        n9435) );
  CLKMX2X2 U10611 ( .A(\I_cache/cache[0][91] ), .B(n7208), .S0(n3265), .Y(
        n9436) );
  CLKMX2X2 U10612 ( .A(\I_cache/cache[7][90] ), .B(n7184), .S0(n3490), .Y(
        n9437) );
  CLKMX2X2 U10613 ( .A(\I_cache/cache[6][90] ), .B(n7184), .S0(n3534), .Y(
        n9438) );
  CLKMX2X2 U10614 ( .A(\I_cache/cache[5][90] ), .B(n7184), .S0(n3400), .Y(
        n9439) );
  CLKMX2X2 U10615 ( .A(\I_cache/cache[4][90] ), .B(n7184), .S0(n3444), .Y(
        n9440) );
  CLKMX2X2 U10616 ( .A(\I_cache/cache[3][90] ), .B(n7184), .S0(n3312), .Y(
        n9441) );
  CLKMX2X2 U10617 ( .A(\I_cache/cache[2][90] ), .B(n7184), .S0(n3355), .Y(
        n9442) );
  CLKMX2X2 U10618 ( .A(\I_cache/cache[1][90] ), .B(n7184), .S0(n3220), .Y(
        n9443) );
  CLKMX2X2 U10619 ( .A(\I_cache/cache[0][90] ), .B(n7184), .S0(n3265), .Y(
        n9444) );
  CLKMX2X2 U10620 ( .A(\I_cache/cache[7][89] ), .B(n7656), .S0(n3490), .Y(
        n9445) );
  CLKMX2X2 U10621 ( .A(\I_cache/cache[6][89] ), .B(n7656), .S0(n3536), .Y(
        n9446) );
  CLKMX2X2 U10622 ( .A(\I_cache/cache[5][89] ), .B(n7656), .S0(n3401), .Y(
        n9447) );
  CLKMX2X2 U10623 ( .A(\I_cache/cache[4][89] ), .B(n7656), .S0(n3446), .Y(
        n9448) );
  CLKMX2X2 U10624 ( .A(\I_cache/cache[3][89] ), .B(n7656), .S0(n3312), .Y(
        n9449) );
  CLKMX2X2 U10625 ( .A(\I_cache/cache[2][89] ), .B(n7656), .S0(n3355), .Y(
        n9450) );
  CLKMX2X2 U10626 ( .A(\I_cache/cache[1][89] ), .B(n7656), .S0(n3223), .Y(
        n9451) );
  CLKMX2X2 U10627 ( .A(\I_cache/cache[0][89] ), .B(n7656), .S0(n3269), .Y(
        n9452) );
  CLKMX2X2 U10628 ( .A(\I_cache/cache[7][88] ), .B(n7434), .S0(n3489), .Y(
        n9453) );
  CLKMX2X2 U10629 ( .A(\I_cache/cache[6][88] ), .B(n7434), .S0(n3533), .Y(
        n9454) );
  CLKMX2X2 U10630 ( .A(\I_cache/cache[5][88] ), .B(n7434), .S0(n3399), .Y(
        n9455) );
  CLKMX2X2 U10631 ( .A(\I_cache/cache[4][88] ), .B(n7434), .S0(n3448), .Y(
        n9456) );
  CLKMX2X2 U10632 ( .A(\I_cache/cache[3][88] ), .B(n7434), .S0(n3311), .Y(
        n9457) );
  CLKMX2X2 U10633 ( .A(\I_cache/cache[2][88] ), .B(n7434), .S0(n3354), .Y(
        n9458) );
  CLKMX2X2 U10634 ( .A(\I_cache/cache[1][88] ), .B(n7434), .S0(n3221), .Y(
        n9459) );
  CLKMX2X2 U10635 ( .A(\I_cache/cache[0][88] ), .B(n7434), .S0(n3266), .Y(
        n9460) );
  CLKMX2X2 U10636 ( .A(\I_cache/cache[7][87] ), .B(n7458), .S0(n3493), .Y(
        n9461) );
  CLKMX2X2 U10637 ( .A(\I_cache/cache[6][87] ), .B(n7458), .S0(n3538), .Y(
        n9462) );
  CLKMX2X2 U10638 ( .A(\I_cache/cache[5][87] ), .B(n7458), .S0(n3403), .Y(
        n9463) );
  CLKMX2X2 U10639 ( .A(\I_cache/cache[4][87] ), .B(n7458), .S0(n3448), .Y(
        n9464) );
  CLKMX2X2 U10640 ( .A(\I_cache/cache[3][87] ), .B(n7458), .S0(n3315), .Y(
        n9465) );
  CLKMX2X2 U10641 ( .A(\I_cache/cache[2][87] ), .B(n7458), .S0(n3358), .Y(
        n9466) );
  CLKMX2X2 U10642 ( .A(\I_cache/cache[1][87] ), .B(n7458), .S0(n3225), .Y(
        n9467) );
  CLKMX2X2 U10643 ( .A(\I_cache/cache[0][87] ), .B(n7458), .S0(n3271), .Y(
        n9468) );
  CLKMX2X2 U10644 ( .A(\I_cache/cache[7][86] ), .B(n8119), .S0(n3497), .Y(
        n9469) );
  CLKMX2X2 U10645 ( .A(\I_cache/cache[6][86] ), .B(n8119), .S0(n3541), .Y(
        n9470) );
  CLKMX2X2 U10646 ( .A(\I_cache/cache[5][86] ), .B(n8119), .S0(n3406), .Y(
        n9471) );
  CLKMX2X2 U10647 ( .A(\I_cache/cache[4][86] ), .B(n8119), .S0(n3452), .Y(
        n9472) );
  CLKMX2X2 U10648 ( .A(\I_cache/cache[3][86] ), .B(n8119), .S0(n3319), .Y(
        n9473) );
  CLKMX2X2 U10649 ( .A(\I_cache/cache[2][86] ), .B(n8119), .S0(n3362), .Y(
        n9474) );
  CLKMX2X2 U10650 ( .A(\I_cache/cache[1][86] ), .B(n8119), .S0(n3229), .Y(
        n9475) );
  CLKMX2X2 U10651 ( .A(\I_cache/cache[0][86] ), .B(n8119), .S0(n3274), .Y(
        n9476) );
  CLKMX2X2 U10652 ( .A(\I_cache/cache[7][85] ), .B(n7482), .S0(n3493), .Y(
        n9477) );
  CLKMX2X2 U10653 ( .A(\I_cache/cache[6][85] ), .B(n7482), .S0(n3538), .Y(
        n9478) );
  CLKMX2X2 U10654 ( .A(\I_cache/cache[5][85] ), .B(n7482), .S0(n3403), .Y(
        n9479) );
  CLKMX2X2 U10655 ( .A(\I_cache/cache[4][85] ), .B(n7482), .S0(n3448), .Y(
        n9480) );
  CLKMX2X2 U10656 ( .A(\I_cache/cache[3][85] ), .B(n7482), .S0(n3315), .Y(
        n9481) );
  CLKMX2X2 U10657 ( .A(\I_cache/cache[2][85] ), .B(n7482), .S0(n3358), .Y(
        n9482) );
  CLKMX2X2 U10658 ( .A(\I_cache/cache[1][85] ), .B(n7482), .S0(n3225), .Y(
        n9483) );
  CLKMX2X2 U10659 ( .A(\I_cache/cache[0][85] ), .B(n7482), .S0(n3271), .Y(
        n9484) );
  CLKMX2X2 U10660 ( .A(\I_cache/cache[7][84] ), .B(n7506), .S0(n3493), .Y(
        n9485) );
  CLKMX2X2 U10661 ( .A(\I_cache/cache[6][84] ), .B(n7506), .S0(n3538), .Y(
        n9486) );
  CLKMX2X2 U10662 ( .A(\I_cache/cache[5][84] ), .B(n7506), .S0(n3403), .Y(
        n9487) );
  CLKMX2X2 U10663 ( .A(\I_cache/cache[4][84] ), .B(n7506), .S0(n3448), .Y(
        n9488) );
  CLKMX2X2 U10664 ( .A(\I_cache/cache[3][84] ), .B(n7506), .S0(n3315), .Y(
        n9489) );
  CLKMX2X2 U10665 ( .A(\I_cache/cache[2][84] ), .B(n7506), .S0(n3358), .Y(
        n9490) );
  CLKMX2X2 U10666 ( .A(\I_cache/cache[1][84] ), .B(n7506), .S0(n3225), .Y(
        n9491) );
  CLKMX2X2 U10667 ( .A(\I_cache/cache[0][84] ), .B(n7506), .S0(n3271), .Y(
        n9492) );
  CLKMX2X2 U10668 ( .A(\I_cache/cache[7][83] ), .B(n7135), .S0(n3491), .Y(
        n9493) );
  CLKMX2X2 U10669 ( .A(\I_cache/cache[6][83] ), .B(n7135), .S0(n3535), .Y(
        n9494) );
  CLKMX2X2 U10670 ( .A(\I_cache/cache[5][83] ), .B(n7135), .S0(n3407), .Y(
        n9495) );
  CLKMX2X2 U10671 ( .A(\I_cache/cache[4][83] ), .B(n7135), .S0(n3445), .Y(
        n9496) );
  CLKMX2X2 U10672 ( .A(\I_cache/cache[3][83] ), .B(n7135), .S0(n3313), .Y(
        n9497) );
  CLKMX2X2 U10673 ( .A(\I_cache/cache[2][83] ), .B(n7135), .S0(n3356), .Y(
        n9498) );
  CLKMX2X2 U10674 ( .A(\I_cache/cache[1][83] ), .B(n7135), .S0(n3223), .Y(
        n9499) );
  CLKMX2X2 U10675 ( .A(\I_cache/cache[0][83] ), .B(n7135), .S0(n3268), .Y(
        n9500) );
  CLKMX2X2 U10676 ( .A(\I_cache/cache[7][82] ), .B(n7159), .S0(n3491), .Y(
        n9501) );
  CLKMX2X2 U10677 ( .A(\I_cache/cache[6][82] ), .B(n7159), .S0(n3535), .Y(
        n9502) );
  CLKMX2X2 U10678 ( .A(\I_cache/cache[5][82] ), .B(n7159), .S0(n3404), .Y(
        n9503) );
  CLKMX2X2 U10679 ( .A(\I_cache/cache[4][82] ), .B(n7159), .S0(n3445), .Y(
        n9504) );
  CLKMX2X2 U10680 ( .A(\I_cache/cache[3][82] ), .B(n7159), .S0(n3313), .Y(
        n9505) );
  CLKMX2X2 U10681 ( .A(\I_cache/cache[2][82] ), .B(n7159), .S0(n3356), .Y(
        n9506) );
  CLKMX2X2 U10682 ( .A(\I_cache/cache[1][82] ), .B(n7159), .S0(n3223), .Y(
        n9507) );
  CLKMX2X2 U10683 ( .A(\I_cache/cache[0][82] ), .B(n7159), .S0(n3268), .Y(
        n9508) );
  CLKMX2X2 U10684 ( .A(\I_cache/cache[7][81] ), .B(n4588), .S0(n3490), .Y(
        n9509) );
  CLKMX2X2 U10685 ( .A(\I_cache/cache[6][81] ), .B(n4588), .S0(n3534), .Y(
        n9510) );
  CLKMX2X2 U10686 ( .A(\I_cache/cache[5][81] ), .B(n4588), .S0(n3400), .Y(
        n9511) );
  CLKMX2X2 U10687 ( .A(\I_cache/cache[4][81] ), .B(n4588), .S0(n3444), .Y(
        n9512) );
  CLKMX2X2 U10688 ( .A(\I_cache/cache[3][81] ), .B(n4588), .S0(n3312), .Y(
        n9513) );
  CLKMX2X2 U10689 ( .A(\I_cache/cache[2][81] ), .B(n4588), .S0(n3355), .Y(
        n9514) );
  CLKMX2X2 U10690 ( .A(\I_cache/cache[1][81] ), .B(n4588), .S0(n3222), .Y(
        n9515) );
  CLKMX2X2 U10691 ( .A(\I_cache/cache[0][81] ), .B(n4588), .S0(n3267), .Y(
        n9516) );
  CLKMX2X2 U10692 ( .A(\I_cache/cache[7][80] ), .B(n7111), .S0(n3490), .Y(
        n9517) );
  CLKMX2X2 U10693 ( .A(\I_cache/cache[6][80] ), .B(n7111), .S0(n3534), .Y(
        n9518) );
  CLKMX2X2 U10694 ( .A(\I_cache/cache[5][80] ), .B(n7111), .S0(n3400), .Y(
        n9519) );
  CLKMX2X2 U10695 ( .A(\I_cache/cache[4][80] ), .B(n7111), .S0(n3444), .Y(
        n9520) );
  CLKMX2X2 U10696 ( .A(\I_cache/cache[3][80] ), .B(n7111), .S0(n3312), .Y(
        n9521) );
  CLKMX2X2 U10697 ( .A(\I_cache/cache[2][80] ), .B(n7111), .S0(n3355), .Y(
        n9522) );
  CLKMX2X2 U10698 ( .A(\I_cache/cache[1][80] ), .B(n7111), .S0(n3223), .Y(
        n9523) );
  CLKMX2X2 U10699 ( .A(\I_cache/cache[0][80] ), .B(n7111), .S0(n3268), .Y(
        n9524) );
  CLKMX2X2 U10700 ( .A(\I_cache/cache[7][79] ), .B(n7554), .S0(n3494), .Y(
        n9525) );
  CLKMX2X2 U10701 ( .A(\I_cache/cache[6][79] ), .B(n7554), .S0(n3539), .Y(
        n9526) );
  CLKMX2X2 U10702 ( .A(\I_cache/cache[5][79] ), .B(n7554), .S0(n3404), .Y(
        n9527) );
  CLKMX2X2 U10703 ( .A(\I_cache/cache[4][79] ), .B(n7554), .S0(n3449), .Y(
        n9528) );
  CLKMX2X2 U10704 ( .A(\I_cache/cache[3][79] ), .B(n7554), .S0(n3316), .Y(
        n9529) );
  CLKMX2X2 U10705 ( .A(\I_cache/cache[2][79] ), .B(n7554), .S0(n3359), .Y(
        n9530) );
  CLKMX2X2 U10706 ( .A(\I_cache/cache[1][79] ), .B(n7554), .S0(n3226), .Y(
        n9531) );
  CLKMX2X2 U10707 ( .A(\I_cache/cache[0][79] ), .B(n7554), .S0(n3272), .Y(
        n9532) );
  CLKMX2X2 U10708 ( .A(\I_cache/cache[7][78] ), .B(n7530), .S0(n3494), .Y(
        n9533) );
  CLKMX2X2 U10709 ( .A(\I_cache/cache[6][78] ), .B(n7530), .S0(n3539), .Y(
        n9534) );
  CLKMX2X2 U10710 ( .A(\I_cache/cache[5][78] ), .B(n7530), .S0(n3404), .Y(
        n9535) );
  CLKMX2X2 U10711 ( .A(\I_cache/cache[4][78] ), .B(n7530), .S0(n3449), .Y(
        n9536) );
  CLKMX2X2 U10712 ( .A(\I_cache/cache[3][78] ), .B(n7530), .S0(n3316), .Y(
        n9537) );
  CLKMX2X2 U10713 ( .A(\I_cache/cache[2][78] ), .B(n7530), .S0(n3359), .Y(
        n9538) );
  CLKMX2X2 U10714 ( .A(\I_cache/cache[1][78] ), .B(n7530), .S0(n3226), .Y(
        n9539) );
  CLKMX2X2 U10715 ( .A(\I_cache/cache[0][78] ), .B(n7530), .S0(n3272), .Y(
        n9540) );
  CLKMX2X2 U10716 ( .A(\I_cache/cache[7][77] ), .B(n7579), .S0(n3494), .Y(
        n9541) );
  CLKMX2X2 U10717 ( .A(\I_cache/cache[6][77] ), .B(n7579), .S0(n3539), .Y(
        n9542) );
  CLKMX2X2 U10718 ( .A(\I_cache/cache[5][77] ), .B(n7579), .S0(n3404), .Y(
        n9543) );
  CLKMX2X2 U10719 ( .A(\I_cache/cache[4][77] ), .B(n7579), .S0(n3449), .Y(
        n9544) );
  CLKMX2X2 U10720 ( .A(\I_cache/cache[3][77] ), .B(n7579), .S0(n3316), .Y(
        n9545) );
  CLKMX2X2 U10721 ( .A(\I_cache/cache[2][77] ), .B(n7579), .S0(n3359), .Y(
        n9546) );
  CLKMX2X2 U10722 ( .A(\I_cache/cache[1][77] ), .B(n7579), .S0(n3226), .Y(
        n9547) );
  CLKMX2X2 U10723 ( .A(\I_cache/cache[0][77] ), .B(n7579), .S0(n3272), .Y(
        n9548) );
  CLKMX2X2 U10724 ( .A(\I_cache/cache[7][76] ), .B(n7627), .S0(n3488), .Y(
        n9549) );
  CLKMX2X2 U10725 ( .A(\I_cache/cache[6][76] ), .B(n7627), .S0(n3536), .Y(
        n9550) );
  CLKMX2X2 U10726 ( .A(\I_cache/cache[5][76] ), .B(n7627), .S0(n3401), .Y(
        n9551) );
  CLKMX2X2 U10727 ( .A(\I_cache/cache[4][76] ), .B(n7627), .S0(n3446), .Y(
        n9552) );
  CLKMX2X2 U10728 ( .A(\I_cache/cache[3][76] ), .B(n7627), .S0(n3313), .Y(
        n9553) );
  CLKMX2X2 U10729 ( .A(\I_cache/cache[2][76] ), .B(n7627), .S0(n3356), .Y(
        n9554) );
  CLKMX2X2 U10730 ( .A(\I_cache/cache[1][76] ), .B(n7627), .S0(n3227), .Y(
        n9555) );
  CLKMX2X2 U10731 ( .A(\I_cache/cache[0][76] ), .B(n7627), .S0(n3269), .Y(
        n9556) );
  CLKMX2X2 U10732 ( .A(\I_cache/cache[7][75] ), .B(n7603), .S0(n3493), .Y(
        n9557) );
  CLKMX2X2 U10733 ( .A(\I_cache/cache[6][75] ), .B(n7603), .S0(n3538), .Y(
        n9558) );
  CLKMX2X2 U10734 ( .A(\I_cache/cache[5][75] ), .B(n7603), .S0(n3403), .Y(
        n9559) );
  CLKMX2X2 U10735 ( .A(\I_cache/cache[4][75] ), .B(n7603), .S0(n3448), .Y(
        n9560) );
  CLKMX2X2 U10736 ( .A(\I_cache/cache[3][75] ), .B(n7603), .S0(n3315), .Y(
        n9561) );
  CLKMX2X2 U10737 ( .A(\I_cache/cache[2][75] ), .B(n7603), .S0(n3358), .Y(
        n9562) );
  CLKMX2X2 U10738 ( .A(\I_cache/cache[1][75] ), .B(n7603), .S0(n3226), .Y(
        n9563) );
  CLKMX2X2 U10739 ( .A(\I_cache/cache[0][75] ), .B(n7603), .S0(n3269), .Y(
        n9564) );
  CLKMX2X2 U10740 ( .A(\I_cache/cache[7][74] ), .B(n7681), .S0(n3491), .Y(
        n9565) );
  CLKMX2X2 U10741 ( .A(\I_cache/cache[6][74] ), .B(n7681), .S0(n3535), .Y(
        n9566) );
  CLKMX2X2 U10742 ( .A(\I_cache/cache[5][74] ), .B(n7681), .S0(n3401), .Y(
        n9567) );
  CLKMX2X2 U10743 ( .A(\I_cache/cache[4][74] ), .B(n7681), .S0(n3445), .Y(
        n9568) );
  CLKMX2X2 U10744 ( .A(\I_cache/cache[3][74] ), .B(n7681), .S0(n3313), .Y(
        n9569) );
  CLKMX2X2 U10745 ( .A(\I_cache/cache[2][74] ), .B(n7681), .S0(n3356), .Y(
        n9570) );
  CLKMX2X2 U10746 ( .A(\I_cache/cache[1][74] ), .B(n7681), .S0(n3224), .Y(
        n9571) );
  CLKMX2X2 U10747 ( .A(\I_cache/cache[0][74] ), .B(n7681), .S0(n3270), .Y(
        n9572) );
  CLKMX2X2 U10748 ( .A(\I_cache/cache[7][73] ), .B(n7704), .S0(n3492), .Y(
        n9573) );
  CLKMX2X2 U10749 ( .A(\I_cache/cache[6][73] ), .B(n7704), .S0(n3537), .Y(
        n9574) );
  CLKMX2X2 U10750 ( .A(\I_cache/cache[5][73] ), .B(n7704), .S0(n3402), .Y(
        n9575) );
  CLKMX2X2 U10751 ( .A(\I_cache/cache[4][73] ), .B(n7704), .S0(n3447), .Y(
        n9576) );
  CLKMX2X2 U10752 ( .A(\I_cache/cache[3][73] ), .B(n7704), .S0(n3314), .Y(
        n9577) );
  CLKMX2X2 U10753 ( .A(\I_cache/cache[2][73] ), .B(n7704), .S0(n3357), .Y(
        n9578) );
  CLKMX2X2 U10754 ( .A(\I_cache/cache[1][73] ), .B(n7704), .S0(n3224), .Y(
        n9579) );
  CLKMX2X2 U10755 ( .A(\I_cache/cache[0][73] ), .B(n7704), .S0(n3270), .Y(
        n9580) );
  CLKMX2X2 U10756 ( .A(\I_cache/cache[7][72] ), .B(n7727), .S0(n3492), .Y(
        n9581) );
  CLKMX2X2 U10757 ( .A(\I_cache/cache[6][72] ), .B(n7727), .S0(n3537), .Y(
        n9582) );
  CLKMX2X2 U10758 ( .A(\I_cache/cache[5][72] ), .B(n7727), .S0(n3402), .Y(
        n9583) );
  CLKMX2X2 U10759 ( .A(\I_cache/cache[4][72] ), .B(n7727), .S0(n3447), .Y(
        n9584) );
  CLKMX2X2 U10760 ( .A(\I_cache/cache[3][72] ), .B(n7727), .S0(n3314), .Y(
        n9585) );
  CLKMX2X2 U10761 ( .A(\I_cache/cache[2][72] ), .B(n7727), .S0(n3357), .Y(
        n9586) );
  CLKMX2X2 U10762 ( .A(\I_cache/cache[1][72] ), .B(n7727), .S0(n3224), .Y(
        n9587) );
  CLKMX2X2 U10763 ( .A(\I_cache/cache[0][72] ), .B(n7727), .S0(n3270), .Y(
        n9588) );
  CLKMX2X2 U10764 ( .A(\I_cache/cache[7][71] ), .B(n7754), .S0(n3489), .Y(
        n9589) );
  CLKMX2X2 U10765 ( .A(\I_cache/cache[6][71] ), .B(n7754), .S0(n3536), .Y(
        n9590) );
  CLKMX2X2 U10766 ( .A(\I_cache/cache[5][71] ), .B(n7754), .S0(n3401), .Y(
        n9591) );
  CLKMX2X2 U10767 ( .A(\I_cache/cache[4][71] ), .B(n7754), .S0(n3446), .Y(
        n9592) );
  CLKMX2X2 U10768 ( .A(\I_cache/cache[3][71] ), .B(n7754), .S0(n3310), .Y(
        n9593) );
  CLKMX2X2 U10769 ( .A(\I_cache/cache[2][71] ), .B(n7754), .S0(n3358), .Y(
        n9594) );
  CLKMX2X2 U10770 ( .A(\I_cache/cache[1][71] ), .B(n7754), .S0(n3224), .Y(
        n9595) );
  CLKMX2X2 U10771 ( .A(\I_cache/cache[0][71] ), .B(n7754), .S0(n3269), .Y(
        n9596) );
  CLKMX2X2 U10772 ( .A(\I_cache/cache[7][70] ), .B(n7777), .S0(n3497), .Y(
        n9597) );
  CLKMX2X2 U10773 ( .A(\I_cache/cache[6][70] ), .B(n7777), .S0(n3541), .Y(
        n9598) );
  CLKMX2X2 U10774 ( .A(\I_cache/cache[5][70] ), .B(n7777), .S0(n3406), .Y(
        n9599) );
  CLKMX2X2 U10775 ( .A(\I_cache/cache[4][70] ), .B(n7777), .S0(n3452), .Y(
        n9600) );
  CLKMX2X2 U10776 ( .A(\I_cache/cache[3][70] ), .B(n7777), .S0(n3319), .Y(
        n9601) );
  CLKMX2X2 U10777 ( .A(\I_cache/cache[2][70] ), .B(n7777), .S0(n3362), .Y(
        n9602) );
  CLKMX2X2 U10778 ( .A(\I_cache/cache[1][70] ), .B(n7777), .S0(n3229), .Y(
        n9603) );
  CLKMX2X2 U10779 ( .A(\I_cache/cache[0][70] ), .B(n7777), .S0(n3274), .Y(
        n9604) );
  CLKMX2X2 U10780 ( .A(\I_cache/cache[7][69] ), .B(n7406), .S0(n3489), .Y(
        n9605) );
  CLKMX2X2 U10781 ( .A(\I_cache/cache[6][69] ), .B(n7406), .S0(n3533), .Y(
        n9606) );
  CLKMX2X2 U10782 ( .A(\I_cache/cache[5][69] ), .B(n7406), .S0(n3399), .Y(
        n9607) );
  CLKMX2X2 U10783 ( .A(\I_cache/cache[4][69] ), .B(n7406), .S0(n3447), .Y(
        n9608) );
  CLKMX2X2 U10784 ( .A(\I_cache/cache[3][69] ), .B(n7406), .S0(n3311), .Y(
        n9609) );
  CLKMX2X2 U10785 ( .A(\I_cache/cache[2][69] ), .B(n7406), .S0(n3354), .Y(
        n9610) );
  CLKMX2X2 U10786 ( .A(\I_cache/cache[1][69] ), .B(n7406), .S0(n3221), .Y(
        n9611) );
  CLKMX2X2 U10787 ( .A(\I_cache/cache[0][69] ), .B(n7406), .S0(n3266), .Y(
        n9612) );
  CLKMX2X2 U10788 ( .A(\I_cache/cache[7][68] ), .B(n8347), .S0(n3497), .Y(
        n9613) );
  CLKMX2X2 U10789 ( .A(\I_cache/cache[6][68] ), .B(n8347), .S0(n3541), .Y(
        n9614) );
  CLKMX2X2 U10790 ( .A(\I_cache/cache[5][68] ), .B(n8347), .S0(n3406), .Y(
        n9615) );
  CLKMX2X2 U10791 ( .A(\I_cache/cache[4][68] ), .B(n8347), .S0(n3452), .Y(
        n9616) );
  CLKMX2X2 U10792 ( .A(\I_cache/cache[3][68] ), .B(n8347), .S0(n3319), .Y(
        n9617) );
  CLKMX2X2 U10793 ( .A(\I_cache/cache[2][68] ), .B(n8347), .S0(n3362), .Y(
        n9618) );
  CLKMX2X2 U10794 ( .A(\I_cache/cache[1][68] ), .B(n8347), .S0(n3229), .Y(
        n9619) );
  CLKMX2X2 U10795 ( .A(\I_cache/cache[0][68] ), .B(n8347), .S0(n3274), .Y(
        n9620) );
  CLKMX2X2 U10796 ( .A(\I_cache/cache[7][67] ), .B(n8366), .S0(n3488), .Y(
        n9621) );
  CLKMX2X2 U10797 ( .A(\I_cache/cache[6][67] ), .B(n8366), .S0(n3532), .Y(
        n9622) );
  CLKMX2X2 U10798 ( .A(\I_cache/cache[5][67] ), .B(n8366), .S0(n3398), .Y(
        n9623) );
  CLKMX2X2 U10799 ( .A(\I_cache/cache[4][67] ), .B(n8366), .S0(n3443), .Y(
        n9624) );
  CLKMX2X2 U10800 ( .A(\I_cache/cache[3][67] ), .B(n8366), .S0(n3310), .Y(
        n9625) );
  CLKMX2X2 U10801 ( .A(\I_cache/cache[2][67] ), .B(n8366), .S0(n3353), .Y(
        n9626) );
  CLKMX2X2 U10802 ( .A(\I_cache/cache[1][67] ), .B(n8366), .S0(n3220), .Y(
        n9627) );
  CLKMX2X2 U10803 ( .A(\I_cache/cache[0][67] ), .B(n8366), .S0(n3265), .Y(
        n9628) );
  CLKMX2X2 U10804 ( .A(\I_cache/cache[7][66] ), .B(n8380), .S0(n3489), .Y(
        n9629) );
  CLKMX2X2 U10805 ( .A(\I_cache/cache[6][66] ), .B(n8380), .S0(n3537), .Y(
        n9630) );
  CLKMX2X2 U10806 ( .A(\I_cache/cache[5][66] ), .B(n8380), .S0(n3407), .Y(
        n9631) );
  CLKMX2X2 U10807 ( .A(\I_cache/cache[4][66] ), .B(n8380), .S0(n3445), .Y(
        n9632) );
  CLKMX2X2 U10808 ( .A(\I_cache/cache[3][66] ), .B(n8380), .S0(n3319), .Y(
        n9633) );
  CLKMX2X2 U10809 ( .A(\I_cache/cache[2][66] ), .B(n8380), .S0(n3362), .Y(
        n9634) );
  CLKMX2X2 U10810 ( .A(\I_cache/cache[1][66] ), .B(n8380), .S0(n3229), .Y(
        n9635) );
  CLKMX2X2 U10811 ( .A(\I_cache/cache[0][66] ), .B(n8380), .S0(n3265), .Y(
        n9636) );
  CLKMX2X2 U10812 ( .A(\I_cache/cache[7][65] ), .B(n4568), .S0(n3490), .Y(
        n9637) );
  CLKMX2X2 U10813 ( .A(\I_cache/cache[6][65] ), .B(n4568), .S0(n3534), .Y(
        n9638) );
  CLKMX2X2 U10814 ( .A(\I_cache/cache[5][65] ), .B(n4568), .S0(n3400), .Y(
        n9639) );
  CLKMX2X2 U10815 ( .A(\I_cache/cache[4][65] ), .B(n4568), .S0(n3444), .Y(
        n9640) );
  CLKMX2X2 U10816 ( .A(\I_cache/cache[3][65] ), .B(n4568), .S0(n3312), .Y(
        n9641) );
  CLKMX2X2 U10817 ( .A(\I_cache/cache[2][65] ), .B(n4568), .S0(n3355), .Y(
        n9642) );
  CLKMX2X2 U10818 ( .A(\I_cache/cache[1][65] ), .B(n4568), .S0(n3222), .Y(
        n9643) );
  CLKMX2X2 U10819 ( .A(\I_cache/cache[0][65] ), .B(n4568), .S0(n3267), .Y(
        n9644) );
  CLKMX2X2 U10820 ( .A(\I_cache/cache[7][63] ), .B(n8408), .S0(n3490), .Y(
        n9653) );
  CLKMX2X2 U10821 ( .A(\I_cache/cache[6][63] ), .B(n8408), .S0(n3538), .Y(
        n9654) );
  CLKMX2X2 U10822 ( .A(\I_cache/cache[5][63] ), .B(n8408), .S0(n3407), .Y(
        n9655) );
  CLKMX2X2 U10823 ( .A(\I_cache/cache[4][63] ), .B(n8408), .S0(n3452), .Y(
        n9656) );
  CLKMX2X2 U10824 ( .A(\I_cache/cache[3][63] ), .B(n8408), .S0(n3310), .Y(
        n9657) );
  CLKMX2X2 U10825 ( .A(\I_cache/cache[2][63] ), .B(n8408), .S0(n3358), .Y(
        n9658) );
  CLKMX2X2 U10826 ( .A(\I_cache/cache[1][63] ), .B(n8408), .S0(n3220), .Y(
        n9659) );
  CLKMX2X2 U10827 ( .A(\I_cache/cache[0][63] ), .B(n8408), .S0(n3266), .Y(
        n9660) );
  CLKMX2X2 U10828 ( .A(\I_cache/cache[7][62] ), .B(n7270), .S0(n3492), .Y(
        n9661) );
  CLKMX2X2 U10829 ( .A(\I_cache/cache[6][62] ), .B(n7270), .S0(n3537), .Y(
        n9662) );
  CLKMX2X2 U10830 ( .A(\I_cache/cache[5][62] ), .B(n7270), .S0(n3402), .Y(
        n9663) );
  CLKMX2X2 U10831 ( .A(\I_cache/cache[4][62] ), .B(n7270), .S0(n3447), .Y(
        n9664) );
  CLKMX2X2 U10832 ( .A(\I_cache/cache[3][62] ), .B(n7270), .S0(n3314), .Y(
        n9665) );
  CLKMX2X2 U10833 ( .A(\I_cache/cache[2][62] ), .B(n7270), .S0(n3357), .Y(
        n9666) );
  CLKMX2X2 U10834 ( .A(\I_cache/cache[1][62] ), .B(n7270), .S0(n3221), .Y(
        n9667) );
  CLKMX2X2 U10835 ( .A(\I_cache/cache[0][62] ), .B(n7270), .S0(n3266), .Y(
        n9668) );
  CLKMX2X2 U10836 ( .A(\I_cache/cache[7][61] ), .B(n7246), .S0(n3488), .Y(
        n9669) );
  CLKMX2X2 U10837 ( .A(\I_cache/cache[6][61] ), .B(n7246), .S0(n3532), .Y(
        n9670) );
  CLKMX2X2 U10838 ( .A(\I_cache/cache[5][61] ), .B(n7246), .S0(n3398), .Y(
        n9671) );
  CLKMX2X2 U10839 ( .A(\I_cache/cache[4][61] ), .B(n7246), .S0(n3443), .Y(
        n9672) );
  CLKMX2X2 U10840 ( .A(\I_cache/cache[3][61] ), .B(n7246), .S0(n3310), .Y(
        n9673) );
  CLKMX2X2 U10841 ( .A(\I_cache/cache[2][61] ), .B(n7246), .S0(n3353), .Y(
        n9674) );
  CLKMX2X2 U10842 ( .A(\I_cache/cache[1][61] ), .B(n7246), .S0(n3220), .Y(
        n9675) );
  CLKMX2X2 U10843 ( .A(\I_cache/cache[0][61] ), .B(n7246), .S0(n3265), .Y(
        n9676) );
  CLKMX2X2 U10844 ( .A(\I_cache/cache[7][60] ), .B(n7222), .S0(n3488), .Y(
        n9677) );
  CLKMX2X2 U10845 ( .A(\I_cache/cache[6][60] ), .B(n7222), .S0(n3532), .Y(
        n9678) );
  CLKMX2X2 U10846 ( .A(\I_cache/cache[5][60] ), .B(n7222), .S0(n3398), .Y(
        n9679) );
  CLKMX2X2 U10847 ( .A(\I_cache/cache[4][60] ), .B(n7222), .S0(n3443), .Y(
        n9680) );
  CLKMX2X2 U10848 ( .A(\I_cache/cache[3][60] ), .B(n7222), .S0(n3310), .Y(
        n9681) );
  CLKMX2X2 U10849 ( .A(\I_cache/cache[2][60] ), .B(n7222), .S0(n3353), .Y(
        n9682) );
  CLKMX2X2 U10850 ( .A(\I_cache/cache[1][60] ), .B(n7222), .S0(n3220), .Y(
        n9683) );
  CLKMX2X2 U10851 ( .A(\I_cache/cache[0][60] ), .B(n7222), .S0(n3265), .Y(
        n9684) );
  CLKMX2X2 U10852 ( .A(\I_cache/cache[7][59] ), .B(n7198), .S0(n3488), .Y(
        n9685) );
  CLKMX2X2 U10853 ( .A(\I_cache/cache[6][59] ), .B(n7198), .S0(n3532), .Y(
        n9686) );
  CLKMX2X2 U10854 ( .A(\I_cache/cache[5][59] ), .B(n7198), .S0(n3398), .Y(
        n9687) );
  CLKMX2X2 U10855 ( .A(\I_cache/cache[4][59] ), .B(n7198), .S0(n3443), .Y(
        n9688) );
  CLKMX2X2 U10856 ( .A(\I_cache/cache[3][59] ), .B(n7198), .S0(n3310), .Y(
        n9689) );
  CLKMX2X2 U10857 ( .A(\I_cache/cache[2][59] ), .B(n7198), .S0(n3353), .Y(
        n9690) );
  CLKMX2X2 U10858 ( .A(\I_cache/cache[1][59] ), .B(n7198), .S0(n3220), .Y(
        n9691) );
  CLKMX2X2 U10859 ( .A(\I_cache/cache[0][59] ), .B(n7198), .S0(n3265), .Y(
        n9692) );
  CLKMX2X2 U10860 ( .A(\I_cache/cache[7][58] ), .B(n7174), .S0(n3491), .Y(
        n9693) );
  CLKMX2X2 U10861 ( .A(\I_cache/cache[6][58] ), .B(n7174), .S0(n3535), .Y(
        n9694) );
  CLKMX2X2 U10862 ( .A(\I_cache/cache[5][58] ), .B(n7174), .S0(n3399), .Y(
        n9695) );
  CLKMX2X2 U10863 ( .A(\I_cache/cache[4][58] ), .B(n7174), .S0(n3445), .Y(
        n9696) );
  CLKMX2X2 U10864 ( .A(\I_cache/cache[3][58] ), .B(n7174), .S0(n3313), .Y(
        n9697) );
  CLKMX2X2 U10865 ( .A(\I_cache/cache[2][58] ), .B(n7174), .S0(n3356), .Y(
        n9698) );
  CLKMX2X2 U10866 ( .A(\I_cache/cache[1][58] ), .B(n7174), .S0(n3222), .Y(
        n9699) );
  CLKMX2X2 U10867 ( .A(\I_cache/cache[0][58] ), .B(n7174), .S0(n3267), .Y(
        n9700) );
  CLKMX2X2 U10868 ( .A(\I_cache/cache[7][57] ), .B(n7646), .S0(n3492), .Y(
        n9701) );
  CLKMX2X2 U10869 ( .A(\I_cache/cache[6][57] ), .B(n7646), .S0(n3536), .Y(
        n9702) );
  CLKMX2X2 U10870 ( .A(\I_cache/cache[5][57] ), .B(n7646), .S0(n3401), .Y(
        n9703) );
  CLKMX2X2 U10871 ( .A(\I_cache/cache[4][57] ), .B(n7646), .S0(n3446), .Y(
        n9704) );
  CLKMX2X2 U10872 ( .A(\I_cache/cache[3][57] ), .B(n7646), .S0(n3311), .Y(
        n9705) );
  CLKMX2X2 U10873 ( .A(\I_cache/cache[2][57] ), .B(n7646), .S0(n3353), .Y(
        n9706) );
  CLKMX2X2 U10874 ( .A(\I_cache/cache[1][57] ), .B(n7646), .S0(n3220), .Y(
        n9707) );
  CLKMX2X2 U10875 ( .A(\I_cache/cache[0][57] ), .B(n7646), .S0(n3269), .Y(
        n9708) );
  CLKMX2X2 U10876 ( .A(\I_cache/cache[7][56] ), .B(n7424), .S0(n3489), .Y(
        n9709) );
  CLKMX2X2 U10877 ( .A(\I_cache/cache[6][56] ), .B(n7424), .S0(n3533), .Y(
        n9710) );
  CLKMX2X2 U10878 ( .A(\I_cache/cache[5][56] ), .B(n7424), .S0(n3399), .Y(
        n9711) );
  CLKMX2X2 U10879 ( .A(\I_cache/cache[4][56] ), .B(n7424), .S0(n3452), .Y(
        n9712) );
  CLKMX2X2 U10880 ( .A(\I_cache/cache[3][56] ), .B(n7424), .S0(n3311), .Y(
        n9713) );
  CLKMX2X2 U10881 ( .A(\I_cache/cache[2][56] ), .B(n7424), .S0(n3354), .Y(
        n9714) );
  CLKMX2X2 U10882 ( .A(\I_cache/cache[1][56] ), .B(n7424), .S0(n3221), .Y(
        n9715) );
  CLKMX2X2 U10883 ( .A(\I_cache/cache[0][56] ), .B(n7424), .S0(n3266), .Y(
        n9716) );
  CLKMX2X2 U10884 ( .A(\I_cache/cache[7][55] ), .B(n7448), .S0(n3489), .Y(
        n9717) );
  CLKMX2X2 U10885 ( .A(\I_cache/cache[6][55] ), .B(n7448), .S0(n3533), .Y(
        n9718) );
  CLKMX2X2 U10886 ( .A(\I_cache/cache[5][55] ), .B(n7448), .S0(n3399), .Y(
        n9719) );
  CLKMX2X2 U10887 ( .A(\I_cache/cache[4][55] ), .B(n7448), .S0(n3444), .Y(
        n9720) );
  CLKMX2X2 U10888 ( .A(\I_cache/cache[3][55] ), .B(n7448), .S0(n3311), .Y(
        n9721) );
  CLKMX2X2 U10889 ( .A(\I_cache/cache[2][55] ), .B(n7448), .S0(n3354), .Y(
        n9722) );
  CLKMX2X2 U10890 ( .A(\I_cache/cache[1][55] ), .B(n7448), .S0(n3225), .Y(
        n9723) );
  CLKMX2X2 U10891 ( .A(\I_cache/cache[0][55] ), .B(n7448), .S0(n3271), .Y(
        n9724) );
  CLKMX2X2 U10892 ( .A(\I_cache/cache[7][54] ), .B(n8108), .S0(n3497), .Y(
        n9725) );
  CLKMX2X2 U10893 ( .A(\I_cache/cache[6][54] ), .B(n8108), .S0(n3541), .Y(
        n9726) );
  CLKMX2X2 U10894 ( .A(\I_cache/cache[5][54] ), .B(n8108), .S0(n3406), .Y(
        n9727) );
  CLKMX2X2 U10895 ( .A(\I_cache/cache[4][54] ), .B(n8108), .S0(n3452), .Y(
        n9728) );
  CLKMX2X2 U10896 ( .A(\I_cache/cache[3][54] ), .B(n8108), .S0(n3319), .Y(
        n9729) );
  CLKMX2X2 U10897 ( .A(\I_cache/cache[2][54] ), .B(n8108), .S0(n3362), .Y(
        n9730) );
  CLKMX2X2 U10898 ( .A(\I_cache/cache[1][54] ), .B(n8108), .S0(n3229), .Y(
        n9731) );
  CLKMX2X2 U10899 ( .A(\I_cache/cache[0][54] ), .B(n8108), .S0(n3274), .Y(
        n9732) );
  CLKMX2X2 U10900 ( .A(\I_cache/cache[7][53] ), .B(n7472), .S0(n3493), .Y(
        n9733) );
  CLKMX2X2 U10901 ( .A(\I_cache/cache[6][53] ), .B(n7472), .S0(n3538), .Y(
        n9734) );
  CLKMX2X2 U10902 ( .A(\I_cache/cache[5][53] ), .B(n7472), .S0(n3403), .Y(
        n9735) );
  CLKMX2X2 U10903 ( .A(\I_cache/cache[4][53] ), .B(n7472), .S0(n3448), .Y(
        n9736) );
  CLKMX2X2 U10904 ( .A(\I_cache/cache[3][53] ), .B(n7472), .S0(n3315), .Y(
        n9737) );
  CLKMX2X2 U10905 ( .A(\I_cache/cache[2][53] ), .B(n7472), .S0(n3358), .Y(
        n9738) );
  CLKMX2X2 U10906 ( .A(\I_cache/cache[1][53] ), .B(n7472), .S0(n3225), .Y(
        n9739) );
  CLKMX2X2 U10907 ( .A(\I_cache/cache[0][53] ), .B(n7472), .S0(n3271), .Y(
        n9740) );
  CLKMX2X2 U10908 ( .A(\I_cache/cache[7][52] ), .B(n7496), .S0(n3493), .Y(
        n9741) );
  CLKMX2X2 U10909 ( .A(\I_cache/cache[6][52] ), .B(n7496), .S0(n3538), .Y(
        n9742) );
  CLKMX2X2 U10910 ( .A(\I_cache/cache[5][52] ), .B(n7496), .S0(n3403), .Y(
        n9743) );
  CLKMX2X2 U10911 ( .A(\I_cache/cache[4][52] ), .B(n7496), .S0(n3448), .Y(
        n9744) );
  CLKMX2X2 U10912 ( .A(\I_cache/cache[3][52] ), .B(n7496), .S0(n3315), .Y(
        n9745) );
  CLKMX2X2 U10913 ( .A(\I_cache/cache[2][52] ), .B(n7496), .S0(n3358), .Y(
        n9746) );
  CLKMX2X2 U10914 ( .A(\I_cache/cache[1][52] ), .B(n7496), .S0(n3225), .Y(
        n9747) );
  CLKMX2X2 U10915 ( .A(\I_cache/cache[0][52] ), .B(n7496), .S0(n3271), .Y(
        n9748) );
  CLKMX2X2 U10916 ( .A(\I_cache/cache[7][51] ), .B(n7125), .S0(n3491), .Y(
        n9749) );
  CLKMX2X2 U10917 ( .A(\I_cache/cache[6][51] ), .B(n7125), .S0(n3535), .Y(
        n9750) );
  CLKMX2X2 U10918 ( .A(\I_cache/cache[5][51] ), .B(n7125), .S0(n3403), .Y(
        n9751) );
  CLKMX2X2 U10919 ( .A(\I_cache/cache[4][51] ), .B(n7125), .S0(n3445), .Y(
        n9752) );
  CLKMX2X2 U10920 ( .A(\I_cache/cache[3][51] ), .B(n7125), .S0(n3313), .Y(
        n9753) );
  CLKMX2X2 U10921 ( .A(\I_cache/cache[2][51] ), .B(n7125), .S0(n3356), .Y(
        n9754) );
  CLKMX2X2 U10922 ( .A(\I_cache/cache[1][51] ), .B(n7125), .S0(n3223), .Y(
        n9755) );
  CLKMX2X2 U10923 ( .A(\I_cache/cache[0][51] ), .B(n7125), .S0(n3268), .Y(
        n9756) );
  CLKMX2X2 U10924 ( .A(\I_cache/cache[7][50] ), .B(n7149), .S0(n3491), .Y(
        n9757) );
  CLKMX2X2 U10925 ( .A(\I_cache/cache[6][50] ), .B(n7149), .S0(n3535), .Y(
        n9758) );
  CLKMX2X2 U10926 ( .A(\I_cache/cache[5][50] ), .B(n7149), .S0(n3402), .Y(
        n9759) );
  CLKMX2X2 U10927 ( .A(\I_cache/cache[4][50] ), .B(n7149), .S0(n3445), .Y(
        n9760) );
  CLKMX2X2 U10928 ( .A(\I_cache/cache[3][50] ), .B(n7149), .S0(n3313), .Y(
        n9761) );
  CLKMX2X2 U10929 ( .A(\I_cache/cache[2][50] ), .B(n7149), .S0(n3356), .Y(
        n9762) );
  CLKMX2X2 U10930 ( .A(\I_cache/cache[1][50] ), .B(n7149), .S0(n3223), .Y(
        n9763) );
  CLKMX2X2 U10931 ( .A(\I_cache/cache[0][50] ), .B(n7149), .S0(n3268), .Y(
        n9764) );
  CLKMX2X2 U10932 ( .A(\I_cache/cache[7][49] ), .B(n4578), .S0(n3490), .Y(
        n9765) );
  CLKMX2X2 U10933 ( .A(\I_cache/cache[6][49] ), .B(n4578), .S0(n3534), .Y(
        n9766) );
  CLKMX2X2 U10934 ( .A(\I_cache/cache[5][49] ), .B(n4578), .S0(n3400), .Y(
        n9767) );
  CLKMX2X2 U10935 ( .A(\I_cache/cache[4][49] ), .B(n4578), .S0(n3444), .Y(
        n9768) );
  CLKMX2X2 U10936 ( .A(\I_cache/cache[3][49] ), .B(n4578), .S0(n3312), .Y(
        n9769) );
  CLKMX2X2 U10937 ( .A(\I_cache/cache[2][49] ), .B(n4578), .S0(n3355), .Y(
        n9770) );
  CLKMX2X2 U10938 ( .A(\I_cache/cache[1][49] ), .B(n4578), .S0(n3222), .Y(
        n9771) );
  CLKMX2X2 U10939 ( .A(\I_cache/cache[0][49] ), .B(n4578), .S0(n3267), .Y(
        n9772) );
  CLKMX2X2 U10940 ( .A(\I_cache/cache[7][48] ), .B(n7101), .S0(n3490), .Y(
        n9773) );
  CLKMX2X2 U10941 ( .A(\I_cache/cache[6][48] ), .B(n7101), .S0(n3534), .Y(
        n9774) );
  CLKMX2X2 U10942 ( .A(\I_cache/cache[5][48] ), .B(n7101), .S0(n3400), .Y(
        n9775) );
  CLKMX2X2 U10943 ( .A(\I_cache/cache[4][48] ), .B(n7101), .S0(n3444), .Y(
        n9776) );
  CLKMX2X2 U10944 ( .A(\I_cache/cache[3][48] ), .B(n7101), .S0(n3312), .Y(
        n9777) );
  CLKMX2X2 U10945 ( .A(\I_cache/cache[2][48] ), .B(n7101), .S0(n3355), .Y(
        n9778) );
  CLKMX2X2 U10946 ( .A(\I_cache/cache[1][48] ), .B(n7101), .S0(n3223), .Y(
        n9779) );
  CLKMX2X2 U10947 ( .A(\I_cache/cache[0][48] ), .B(n7101), .S0(n3268), .Y(
        n9780) );
  CLKMX2X2 U10948 ( .A(\I_cache/cache[7][47] ), .B(n7544), .S0(n3494), .Y(
        n9781) );
  CLKMX2X2 U10949 ( .A(\I_cache/cache[6][47] ), .B(n7544), .S0(n3539), .Y(
        n9782) );
  CLKMX2X2 U10950 ( .A(\I_cache/cache[5][47] ), .B(n7544), .S0(n3404), .Y(
        n9783) );
  CLKMX2X2 U10951 ( .A(\I_cache/cache[4][47] ), .B(n7544), .S0(n3449), .Y(
        n9784) );
  CLKMX2X2 U10952 ( .A(\I_cache/cache[3][47] ), .B(n7544), .S0(n3316), .Y(
        n9785) );
  CLKMX2X2 U10953 ( .A(\I_cache/cache[2][47] ), .B(n7544), .S0(n3359), .Y(
        n9786) );
  CLKMX2X2 U10954 ( .A(\I_cache/cache[1][47] ), .B(n7544), .S0(n3226), .Y(
        n9787) );
  CLKMX2X2 U10955 ( .A(\I_cache/cache[0][47] ), .B(n7544), .S0(n3272), .Y(
        n9788) );
  CLKMX2X2 U10956 ( .A(\I_cache/cache[7][46] ), .B(n7520), .S0(n3493), .Y(
        n9789) );
  CLKMX2X2 U10957 ( .A(\I_cache/cache[6][46] ), .B(n7520), .S0(n3538), .Y(
        n9790) );
  CLKMX2X2 U10958 ( .A(\I_cache/cache[5][46] ), .B(n7520), .S0(n3403), .Y(
        n9791) );
  CLKMX2X2 U10959 ( .A(\I_cache/cache[4][46] ), .B(n7520), .S0(n3448), .Y(
        n9792) );
  CLKMX2X2 U10960 ( .A(\I_cache/cache[3][46] ), .B(n7520), .S0(n3315), .Y(
        n9793) );
  CLKMX2X2 U10961 ( .A(\I_cache/cache[2][46] ), .B(n7520), .S0(n3358), .Y(
        n9794) );
  CLKMX2X2 U10962 ( .A(\I_cache/cache[1][46] ), .B(n7520), .S0(n3224), .Y(
        n9795) );
  CLKMX2X2 U10963 ( .A(\I_cache/cache[0][46] ), .B(n7520), .S0(n3272), .Y(
        n9796) );
  CLKMX2X2 U10964 ( .A(\I_cache/cache[7][45] ), .B(n7569), .S0(n3494), .Y(
        n9797) );
  CLKMX2X2 U10965 ( .A(\I_cache/cache[6][45] ), .B(n7569), .S0(n3539), .Y(
        n9798) );
  CLKMX2X2 U10966 ( .A(\I_cache/cache[5][45] ), .B(n7569), .S0(n3404), .Y(
        n9799) );
  CLKMX2X2 U10967 ( .A(\I_cache/cache[4][45] ), .B(n7569), .S0(n3449), .Y(
        n9800) );
  CLKMX2X2 U10968 ( .A(\I_cache/cache[3][45] ), .B(n7569), .S0(n3316), .Y(
        n9801) );
  CLKMX2X2 U10969 ( .A(\I_cache/cache[2][45] ), .B(n7569), .S0(n3359), .Y(
        n9802) );
  CLKMX2X2 U10970 ( .A(\I_cache/cache[1][45] ), .B(n7569), .S0(n3226), .Y(
        n9803) );
  CLKMX2X2 U10971 ( .A(\I_cache/cache[0][45] ), .B(n7569), .S0(n3272), .Y(
        n9804) );
  CLKMX2X2 U10972 ( .A(\I_cache/cache[7][44] ), .B(n7618), .S0(n3488), .Y(
        n9805) );
  CLKMX2X2 U10973 ( .A(\I_cache/cache[6][44] ), .B(n7618), .S0(n3536), .Y(
        n9806) );
  CLKMX2X2 U10974 ( .A(\I_cache/cache[5][44] ), .B(n7618), .S0(n3401), .Y(
        n9807) );
  CLKMX2X2 U10975 ( .A(\I_cache/cache[4][44] ), .B(n7618), .S0(n3446), .Y(
        n9808) );
  CLKMX2X2 U10976 ( .A(\I_cache/cache[3][44] ), .B(n7618), .S0(n3312), .Y(
        n9809) );
  CLKMX2X2 U10977 ( .A(\I_cache/cache[2][44] ), .B(n7618), .S0(n3354), .Y(
        n9810) );
  CLKMX2X2 U10978 ( .A(\I_cache/cache[1][44] ), .B(n7618), .S0(n3221), .Y(
        n9811) );
  CLKMX2X2 U10979 ( .A(\I_cache/cache[0][44] ), .B(n7618), .S0(n3269), .Y(
        n9812) );
  CLKMX2X2 U10980 ( .A(\I_cache/cache[7][43] ), .B(n7593), .S0(n3494), .Y(
        n9813) );
  CLKMX2X2 U10981 ( .A(\I_cache/cache[6][43] ), .B(n7593), .S0(n3539), .Y(
        n9814) );
  CLKMX2X2 U10982 ( .A(\I_cache/cache[5][43] ), .B(n7593), .S0(n3404), .Y(
        n9815) );
  CLKMX2X2 U10983 ( .A(\I_cache/cache[4][43] ), .B(n7593), .S0(n3449), .Y(
        n9816) );
  CLKMX2X2 U10984 ( .A(\I_cache/cache[3][43] ), .B(n7593), .S0(n3316), .Y(
        n9817) );
  CLKMX2X2 U10985 ( .A(\I_cache/cache[2][43] ), .B(n7593), .S0(n3359), .Y(
        n9818) );
  CLKMX2X2 U10986 ( .A(\I_cache/cache[1][43] ), .B(n7593), .S0(n3226), .Y(
        n9819) );
  CLKMX2X2 U10987 ( .A(\I_cache/cache[0][43] ), .B(n7593), .S0(n3271), .Y(
        n9820) );
  CLKMX2X2 U10988 ( .A(\I_cache/cache[7][42] ), .B(n7671), .S0(n3489), .Y(
        n9821) );
  CLKMX2X2 U10989 ( .A(\I_cache/cache[6][42] ), .B(n7671), .S0(n3536), .Y(
        n9822) );
  CLKMX2X2 U10990 ( .A(\I_cache/cache[5][42] ), .B(n7671), .S0(n3401), .Y(
        n9823) );
  CLKMX2X2 U10991 ( .A(\I_cache/cache[4][42] ), .B(n7671), .S0(n3446), .Y(
        n9824) );
  CLKMX2X2 U10992 ( .A(\I_cache/cache[3][42] ), .B(n7671), .S0(n3313), .Y(
        n9825) );
  CLKMX2X2 U10993 ( .A(\I_cache/cache[2][42] ), .B(n7671), .S0(n3355), .Y(
        n9826) );
  CLKMX2X2 U10994 ( .A(\I_cache/cache[1][42] ), .B(n7671), .S0(n3223), .Y(
        n9827) );
  CLKMX2X2 U10995 ( .A(\I_cache/cache[0][42] ), .B(n7671), .S0(n3268), .Y(
        n9828) );
  CLKMX2X2 U10996 ( .A(\I_cache/cache[7][41] ), .B(n7695), .S0(n3492), .Y(
        n9829) );
  CLKMX2X2 U10997 ( .A(\I_cache/cache[6][41] ), .B(n7695), .S0(n3537), .Y(
        n9830) );
  CLKMX2X2 U10998 ( .A(\I_cache/cache[5][41] ), .B(n7695), .S0(n3402), .Y(
        n9831) );
  CLKMX2X2 U10999 ( .A(\I_cache/cache[4][41] ), .B(n7695), .S0(n3447), .Y(
        n9832) );
  CLKMX2X2 U11000 ( .A(\I_cache/cache[3][41] ), .B(n7695), .S0(n3314), .Y(
        n9833) );
  CLKMX2X2 U11001 ( .A(\I_cache/cache[2][41] ), .B(n7695), .S0(n3357), .Y(
        n9834) );
  CLKMX2X2 U11002 ( .A(\I_cache/cache[1][41] ), .B(n7695), .S0(n3224), .Y(
        n9835) );
  CLKMX2X2 U11003 ( .A(\I_cache/cache[0][41] ), .B(n7695), .S0(n3270), .Y(
        n9836) );
  CLKMX2X2 U11004 ( .A(\I_cache/cache[7][40] ), .B(n7718), .S0(n3492), .Y(
        n9837) );
  CLKMX2X2 U11005 ( .A(\I_cache/cache[6][40] ), .B(n7718), .S0(n3537), .Y(
        n9838) );
  CLKMX2X2 U11006 ( .A(\I_cache/cache[5][40] ), .B(n7718), .S0(n3402), .Y(
        n9839) );
  CLKMX2X2 U11007 ( .A(\I_cache/cache[4][40] ), .B(n7718), .S0(n3447), .Y(
        n9840) );
  CLKMX2X2 U11008 ( .A(\I_cache/cache[3][40] ), .B(n7718), .S0(n3314), .Y(
        n9841) );
  CLKMX2X2 U11009 ( .A(\I_cache/cache[2][40] ), .B(n7718), .S0(n3357), .Y(
        n9842) );
  CLKMX2X2 U11010 ( .A(\I_cache/cache[1][40] ), .B(n7718), .S0(n3224), .Y(
        n9843) );
  CLKMX2X2 U11011 ( .A(\I_cache/cache[0][40] ), .B(n7718), .S0(n3270), .Y(
        n9844) );
  CLKMX2X2 U11012 ( .A(\I_cache/cache[7][39] ), .B(n7744), .S0(n3492), .Y(
        n9845) );
  CLKMX2X2 U11013 ( .A(\I_cache/cache[6][39] ), .B(n7744), .S0(n3537), .Y(
        n9846) );
  CLKMX2X2 U11014 ( .A(\I_cache/cache[5][39] ), .B(n7744), .S0(n3402), .Y(
        n9847) );
  CLKMX2X2 U11015 ( .A(\I_cache/cache[4][39] ), .B(n7744), .S0(n3447), .Y(
        n9848) );
  CLKMX2X2 U11016 ( .A(\I_cache/cache[3][39] ), .B(n7744), .S0(n3314), .Y(
        n9849) );
  CLKMX2X2 U11017 ( .A(\I_cache/cache[2][39] ), .B(n7744), .S0(n3357), .Y(
        n9850) );
  CLKMX2X2 U11018 ( .A(\I_cache/cache[1][39] ), .B(n7744), .S0(n3224), .Y(
        n9851) );
  CLKMX2X2 U11019 ( .A(\I_cache/cache[0][39] ), .B(n7744), .S0(n3270), .Y(
        n9852) );
  CLKMX2X2 U11020 ( .A(\I_cache/cache[7][38] ), .B(n7768), .S0(n3497), .Y(
        n9853) );
  CLKMX2X2 U11021 ( .A(\I_cache/cache[6][38] ), .B(n7768), .S0(n3541), .Y(
        n9854) );
  CLKMX2X2 U11022 ( .A(\I_cache/cache[5][38] ), .B(n7768), .S0(n3406), .Y(
        n9855) );
  CLKMX2X2 U11023 ( .A(\I_cache/cache[4][38] ), .B(n7768), .S0(n3452), .Y(
        n9856) );
  CLKMX2X2 U11024 ( .A(\I_cache/cache[3][38] ), .B(n7768), .S0(n3319), .Y(
        n9857) );
  CLKMX2X2 U11025 ( .A(\I_cache/cache[2][38] ), .B(n7768), .S0(n3362), .Y(
        n9858) );
  CLKMX2X2 U11026 ( .A(\I_cache/cache[1][38] ), .B(n7768), .S0(n3229), .Y(
        n9859) );
  CLKMX2X2 U11027 ( .A(\I_cache/cache[0][38] ), .B(n7768), .S0(n3274), .Y(
        n9860) );
  CLKMX2X2 U11028 ( .A(\I_cache/cache[7][37] ), .B(n7396), .S0(n3489), .Y(
        n9861) );
  CLKMX2X2 U11029 ( .A(\I_cache/cache[6][37] ), .B(n7396), .S0(n3533), .Y(
        n9862) );
  CLKMX2X2 U11030 ( .A(\I_cache/cache[5][37] ), .B(n7396), .S0(n3399), .Y(
        n9863) );
  CLKMX2X2 U11031 ( .A(\I_cache/cache[4][37] ), .B(n7396), .S0(n3445), .Y(
        n9864) );
  CLKMX2X2 U11032 ( .A(\I_cache/cache[3][37] ), .B(n7396), .S0(n3311), .Y(
        n9865) );
  CLKMX2X2 U11033 ( .A(\I_cache/cache[2][37] ), .B(n7396), .S0(n3354), .Y(
        n9866) );
  CLKMX2X2 U11034 ( .A(\I_cache/cache[1][37] ), .B(n7396), .S0(n3221), .Y(
        n9867) );
  CLKMX2X2 U11035 ( .A(\I_cache/cache[0][37] ), .B(n7396), .S0(n3266), .Y(
        n9868) );
  CLKMX2X2 U11036 ( .A(\I_cache/cache[7][36] ), .B(n8345), .S0(n3497), .Y(
        n9869) );
  CLKMX2X2 U11037 ( .A(\I_cache/cache[6][36] ), .B(n8345), .S0(n3541), .Y(
        n9870) );
  CLKMX2X2 U11038 ( .A(\I_cache/cache[5][36] ), .B(n8345), .S0(n3406), .Y(
        n9871) );
  CLKMX2X2 U11039 ( .A(\I_cache/cache[4][36] ), .B(n8345), .S0(n3452), .Y(
        n9872) );
  CLKMX2X2 U11040 ( .A(\I_cache/cache[3][36] ), .B(n8345), .S0(n3319), .Y(
        n9873) );
  CLKMX2X2 U11041 ( .A(\I_cache/cache[2][36] ), .B(n8345), .S0(n3362), .Y(
        n9874) );
  CLKMX2X2 U11042 ( .A(\I_cache/cache[1][36] ), .B(n8345), .S0(n3229), .Y(
        n9875) );
  CLKMX2X2 U11043 ( .A(\I_cache/cache[0][36] ), .B(n8345), .S0(n3274), .Y(
        n9876) );
  CLKMX2X2 U11044 ( .A(\I_cache/cache[7][35] ), .B(n8364), .S0(n3497), .Y(
        n9877) );
  CLKMX2X2 U11045 ( .A(\I_cache/cache[6][35] ), .B(n8364), .S0(n3541), .Y(
        n9878) );
  CLKMX2X2 U11046 ( .A(\I_cache/cache[5][35] ), .B(n8364), .S0(n3406), .Y(
        n9879) );
  CLKMX2X2 U11047 ( .A(\I_cache/cache[4][35] ), .B(n8364), .S0(n3452), .Y(
        n9880) );
  CLKMX2X2 U11048 ( .A(\I_cache/cache[3][35] ), .B(n8364), .S0(n3319), .Y(
        n9881) );
  CLKMX2X2 U11049 ( .A(\I_cache/cache[2][35] ), .B(n8364), .S0(n3362), .Y(
        n9882) );
  CLKMX2X2 U11050 ( .A(\I_cache/cache[1][35] ), .B(n8364), .S0(n3229), .Y(
        n9883) );
  CLKMX2X2 U11051 ( .A(\I_cache/cache[0][35] ), .B(n8364), .S0(n3274), .Y(
        n9884) );
  CLKMX2X2 U11052 ( .A(\I_cache/cache[7][34] ), .B(n8378), .S0(n3497), .Y(
        n9885) );
  CLKMX2X2 U11053 ( .A(\I_cache/cache[6][34] ), .B(n8378), .S0(n3537), .Y(
        n9886) );
  CLKMX2X2 U11054 ( .A(\I_cache/cache[5][34] ), .B(n8378), .S0(n3407), .Y(
        n9887) );
  CLKMX2X2 U11055 ( .A(\I_cache/cache[4][34] ), .B(n8378), .S0(n3444), .Y(
        n9888) );
  CLKMX2X2 U11056 ( .A(\I_cache/cache[3][34] ), .B(n8378), .S0(n3311), .Y(
        n9889) );
  CLKMX2X2 U11057 ( .A(\I_cache/cache[2][34] ), .B(n8378), .S0(n3353), .Y(
        n9890) );
  CLKMX2X2 U11058 ( .A(\I_cache/cache[1][34] ), .B(n8378), .S0(n3221), .Y(
        n9891) );
  CLKMX2X2 U11059 ( .A(\I_cache/cache[0][34] ), .B(n8378), .S0(n3267), .Y(
        n9892) );
  CLKMX2X2 U11060 ( .A(\I_cache/cache[7][33] ), .B(n4558), .S0(n3490), .Y(
        n9893) );
  CLKMX2X2 U11061 ( .A(\I_cache/cache[6][33] ), .B(n4558), .S0(n3534), .Y(
        n9894) );
  CLKMX2X2 U11062 ( .A(\I_cache/cache[5][33] ), .B(n4558), .S0(n3400), .Y(
        n9895) );
  CLKMX2X2 U11063 ( .A(\I_cache/cache[4][33] ), .B(n4558), .S0(n3444), .Y(
        n9896) );
  CLKMX2X2 U11064 ( .A(\I_cache/cache[3][33] ), .B(n4558), .S0(n3312), .Y(
        n9897) );
  CLKMX2X2 U11065 ( .A(\I_cache/cache[2][33] ), .B(n4558), .S0(n3355), .Y(
        n9898) );
  CLKMX2X2 U11066 ( .A(\I_cache/cache[1][33] ), .B(n4558), .S0(n3222), .Y(
        n9899) );
  CLKMX2X2 U11067 ( .A(\I_cache/cache[0][33] ), .B(n4558), .S0(n3267), .Y(
        n9900) );
  CLKMX2X2 U11068 ( .A(\I_cache/cache[7][31] ), .B(n8407), .S0(n3497), .Y(
        n9909) );
  CLKMX2X2 U11069 ( .A(\I_cache/cache[6][31] ), .B(n8407), .S0(n3532), .Y(
        n9910) );
  CLKMX2X2 U11070 ( .A(\I_cache/cache[5][31] ), .B(n8407), .S0(n3407), .Y(
        n9911) );
  CLKMX2X2 U11071 ( .A(\I_cache/cache[4][31] ), .B(n8407), .S0(n3445), .Y(
        n9912) );
  CLKMX2X2 U11072 ( .A(\I_cache/cache[3][31] ), .B(n8407), .S0(n3312), .Y(
        n9913) );
  CLKMX2X2 U11073 ( .A(\I_cache/cache[2][31] ), .B(n8407), .S0(n3354), .Y(
        n9914) );
  CLKMX2X2 U11074 ( .A(\I_cache/cache[1][31] ), .B(n8407), .S0(n3222), .Y(
        n9915) );
  CLKMX2X2 U11075 ( .A(\I_cache/cache[0][31] ), .B(n8407), .S0(n3268), .Y(
        n9916) );
  CLKMX2X2 U11076 ( .A(\I_cache/cache[7][30] ), .B(n7265), .S0(n3489), .Y(
        n9917) );
  CLKMX2X2 U11077 ( .A(\I_cache/cache[6][30] ), .B(n7265), .S0(n3533), .Y(
        n9918) );
  CLKMX2X2 U11078 ( .A(\I_cache/cache[5][30] ), .B(n7265), .S0(n3399), .Y(
        n9919) );
  CLKMX2X2 U11079 ( .A(\I_cache/cache[4][30] ), .B(n7265), .S0(n3443), .Y(
        n9920) );
  CLKMX2X2 U11080 ( .A(\I_cache/cache[3][30] ), .B(n7265), .S0(n3311), .Y(
        n9921) );
  CLKMX2X2 U11081 ( .A(\I_cache/cache[2][30] ), .B(n7265), .S0(n3354), .Y(
        n9922) );
  CLKMX2X2 U11082 ( .A(\I_cache/cache[1][30] ), .B(n7265), .S0(n3224), .Y(
        n9923) );
  CLKMX2X2 U11083 ( .A(\I_cache/cache[0][30] ), .B(n7265), .S0(n3266), .Y(
        n9924) );
  CLKMX2X2 U11084 ( .A(\I_cache/cache[7][29] ), .B(n7241), .S0(n3488), .Y(
        n9925) );
  CLKMX2X2 U11085 ( .A(\I_cache/cache[6][29] ), .B(n7241), .S0(n3532), .Y(
        n9926) );
  CLKMX2X2 U11086 ( .A(\I_cache/cache[5][29] ), .B(n7241), .S0(n3398), .Y(
        n9927) );
  CLKMX2X2 U11087 ( .A(\I_cache/cache[4][29] ), .B(n7241), .S0(n3443), .Y(
        n9928) );
  CLKMX2X2 U11088 ( .A(\I_cache/cache[3][29] ), .B(n7241), .S0(n3310), .Y(
        n9929) );
  CLKMX2X2 U11089 ( .A(\I_cache/cache[2][29] ), .B(n7241), .S0(n3353), .Y(
        n9930) );
  CLKMX2X2 U11090 ( .A(\I_cache/cache[1][29] ), .B(n7241), .S0(n3220), .Y(
        n9931) );
  CLKMX2X2 U11091 ( .A(\I_cache/cache[0][29] ), .B(n7241), .S0(n3265), .Y(
        n9932) );
  CLKMX2X2 U11092 ( .A(\I_cache/cache[7][28] ), .B(n7217), .S0(n3488), .Y(
        n9933) );
  CLKMX2X2 U11093 ( .A(\I_cache/cache[6][28] ), .B(n7217), .S0(n3532), .Y(
        n9934) );
  CLKMX2X2 U11094 ( .A(\I_cache/cache[5][28] ), .B(n7217), .S0(n3398), .Y(
        n9935) );
  CLKMX2X2 U11095 ( .A(\I_cache/cache[4][28] ), .B(n7217), .S0(n3443), .Y(
        n9936) );
  CLKMX2X2 U11096 ( .A(\I_cache/cache[3][28] ), .B(n7217), .S0(n3310), .Y(
        n9937) );
  CLKMX2X2 U11097 ( .A(\I_cache/cache[2][28] ), .B(n7217), .S0(n3353), .Y(
        n9938) );
  CLKMX2X2 U11098 ( .A(\I_cache/cache[1][28] ), .B(n7217), .S0(n3220), .Y(
        n9939) );
  CLKMX2X2 U11099 ( .A(\I_cache/cache[0][28] ), .B(n7217), .S0(n3265), .Y(
        n9940) );
  CLKMX2X2 U11100 ( .A(\I_cache/cache[7][27] ), .B(n7193), .S0(n3488), .Y(
        n9941) );
  CLKMX2X2 U11101 ( .A(\I_cache/cache[6][27] ), .B(n7193), .S0(n3532), .Y(
        n9942) );
  CLKMX2X2 U11102 ( .A(\I_cache/cache[5][27] ), .B(n7193), .S0(n3398), .Y(
        n9943) );
  CLKMX2X2 U11103 ( .A(\I_cache/cache[4][27] ), .B(n7193), .S0(n3443), .Y(
        n9944) );
  CLKMX2X2 U11104 ( .A(\I_cache/cache[3][27] ), .B(n7193), .S0(n3310), .Y(
        n9945) );
  CLKMX2X2 U11105 ( .A(\I_cache/cache[2][27] ), .B(n7193), .S0(n3353), .Y(
        n9946) );
  CLKMX2X2 U11106 ( .A(\I_cache/cache[1][27] ), .B(n7193), .S0(n3220), .Y(
        n9947) );
  CLKMX2X2 U11107 ( .A(\I_cache/cache[0][27] ), .B(n7193), .S0(n3265), .Y(
        n9948) );
  CLKMX2X2 U11108 ( .A(\I_cache/cache[7][26] ), .B(n7169), .S0(n3491), .Y(
        n9949) );
  CLKMX2X2 U11109 ( .A(\I_cache/cache[6][26] ), .B(n7169), .S0(n3535), .Y(
        n9950) );
  CLKMX2X2 U11110 ( .A(\I_cache/cache[5][26] ), .B(n7169), .S0(n3405), .Y(
        n9951) );
  CLKMX2X2 U11111 ( .A(\I_cache/cache[4][26] ), .B(n7169), .S0(n3445), .Y(
        n9952) );
  CLKMX2X2 U11112 ( .A(\I_cache/cache[3][26] ), .B(n7169), .S0(n3313), .Y(
        n9953) );
  CLKMX2X2 U11113 ( .A(\I_cache/cache[2][26] ), .B(n7169), .S0(n3356), .Y(
        n9954) );
  CLKMX2X2 U11114 ( .A(\I_cache/cache[1][26] ), .B(n7169), .S0(n3223), .Y(
        n9955) );
  CLKMX2X2 U11115 ( .A(\I_cache/cache[0][26] ), .B(n7169), .S0(n3267), .Y(
        n9956) );
  CLKMX2X2 U11116 ( .A(\I_cache/cache[7][25] ), .B(n7641), .S0(n3490), .Y(
        n9957) );
  CLKMX2X2 U11117 ( .A(\I_cache/cache[6][25] ), .B(n7641), .S0(n3536), .Y(
        n9958) );
  CLKMX2X2 U11118 ( .A(\I_cache/cache[5][25] ), .B(n7641), .S0(n3401), .Y(
        n9959) );
  CLKMX2X2 U11119 ( .A(\I_cache/cache[4][25] ), .B(n7641), .S0(n3446), .Y(
        n9960) );
  CLKMX2X2 U11120 ( .A(\I_cache/cache[3][25] ), .B(n7641), .S0(n3314), .Y(
        n9961) );
  CLKMX2X2 U11121 ( .A(\I_cache/cache[2][25] ), .B(n7641), .S0(n3356), .Y(
        n9962) );
  CLKMX2X2 U11122 ( .A(\I_cache/cache[1][25] ), .B(n7641), .S0(n3222), .Y(
        n9963) );
  CLKMX2X2 U11123 ( .A(\I_cache/cache[0][25] ), .B(n7641), .S0(n3269), .Y(
        n9964) );
  CLKMX2X2 U11124 ( .A(\I_cache/cache[7][24] ), .B(n7419), .S0(n3489), .Y(
        n9965) );
  CLKMX2X2 U11125 ( .A(\I_cache/cache[6][24] ), .B(n7419), .S0(n3533), .Y(
        n9966) );
  CLKMX2X2 U11126 ( .A(\I_cache/cache[5][24] ), .B(n7419), .S0(n3399), .Y(
        n9967) );
  CLKMX2X2 U11127 ( .A(\I_cache/cache[4][24] ), .B(n7419), .S0(n3448), .Y(
        n9968) );
  CLKMX2X2 U11128 ( .A(\I_cache/cache[3][24] ), .B(n7419), .S0(n3311), .Y(
        n9969) );
  CLKMX2X2 U11129 ( .A(\I_cache/cache[2][24] ), .B(n7419), .S0(n3354), .Y(
        n9970) );
  CLKMX2X2 U11130 ( .A(\I_cache/cache[1][24] ), .B(n7419), .S0(n3221), .Y(
        n9971) );
  CLKMX2X2 U11131 ( .A(\I_cache/cache[0][24] ), .B(n7419), .S0(n3266), .Y(
        n9972) );
  CLKMX2X2 U11132 ( .A(\I_cache/cache[7][23] ), .B(n7443), .S0(n3489), .Y(
        n9973) );
  CLKMX2X2 U11133 ( .A(\I_cache/cache[6][23] ), .B(n7443), .S0(n3533), .Y(
        n9974) );
  CLKMX2X2 U11134 ( .A(\I_cache/cache[5][23] ), .B(n7443), .S0(n3399), .Y(
        n9975) );
  CLKMX2X2 U11135 ( .A(\I_cache/cache[4][23] ), .B(n7443), .S0(n3447), .Y(
        n9976) );
  CLKMX2X2 U11136 ( .A(\I_cache/cache[3][23] ), .B(n7443), .S0(n3311), .Y(
        n9977) );
  CLKMX2X2 U11137 ( .A(\I_cache/cache[2][23] ), .B(n7443), .S0(n3354), .Y(
        n9978) );
  CLKMX2X2 U11138 ( .A(\I_cache/cache[1][23] ), .B(n7443), .S0(n3221), .Y(
        n9979) );
  CLKMX2X2 U11139 ( .A(\I_cache/cache[0][23] ), .B(n7443), .S0(n3271), .Y(
        n9980) );
  CLKMX2X2 U11140 ( .A(\I_cache/cache[7][22] ), .B(n8103), .S0(n3497), .Y(
        n9981) );
  CLKMX2X2 U11141 ( .A(\I_cache/cache[6][22] ), .B(n8103), .S0(n3541), .Y(
        n9982) );
  CLKMX2X2 U11142 ( .A(\I_cache/cache[5][22] ), .B(n8103), .S0(n3406), .Y(
        n9983) );
  CLKMX2X2 U11143 ( .A(\I_cache/cache[4][22] ), .B(n8103), .S0(n3452), .Y(
        n9984) );
  CLKMX2X2 U11144 ( .A(\I_cache/cache[3][22] ), .B(n8103), .S0(n3319), .Y(
        n9985) );
  CLKMX2X2 U11145 ( .A(\I_cache/cache[2][22] ), .B(n8103), .S0(n3362), .Y(
        n9986) );
  CLKMX2X2 U11146 ( .A(\I_cache/cache[1][22] ), .B(n8103), .S0(n3229), .Y(
        n9987) );
  CLKMX2X2 U11147 ( .A(\I_cache/cache[0][22] ), .B(n8103), .S0(n3274), .Y(
        n9988) );
  CLKMX2X2 U11148 ( .A(\I_cache/cache[7][21] ), .B(n7467), .S0(n3493), .Y(
        n9989) );
  CLKMX2X2 U11149 ( .A(\I_cache/cache[6][21] ), .B(n7467), .S0(n3538), .Y(
        n9990) );
  CLKMX2X2 U11150 ( .A(\I_cache/cache[5][21] ), .B(n7467), .S0(n3403), .Y(
        n9991) );
  CLKMX2X2 U11151 ( .A(\I_cache/cache[4][21] ), .B(n7467), .S0(n3448), .Y(
        n9992) );
  CLKMX2X2 U11152 ( .A(\I_cache/cache[3][21] ), .B(n7467), .S0(n3315), .Y(
        n9993) );
  CLKMX2X2 U11153 ( .A(\I_cache/cache[2][21] ), .B(n7467), .S0(n3358), .Y(
        n9994) );
  CLKMX2X2 U11154 ( .A(\I_cache/cache[1][21] ), .B(n7467), .S0(n3225), .Y(
        n9995) );
  CLKMX2X2 U11155 ( .A(\I_cache/cache[0][21] ), .B(n7467), .S0(n3271), .Y(
        n9996) );
  CLKMX2X2 U11156 ( .A(\I_cache/cache[7][20] ), .B(n7491), .S0(n3493), .Y(
        n9997) );
  CLKMX2X2 U11157 ( .A(\I_cache/cache[6][20] ), .B(n7491), .S0(n3538), .Y(
        n9998) );
  CLKMX2X2 U11158 ( .A(\I_cache/cache[5][20] ), .B(n7491), .S0(n3403), .Y(
        n9999) );
  CLKMX2X2 U11159 ( .A(\I_cache/cache[4][20] ), .B(n7491), .S0(n3448), .Y(
        n10000) );
  CLKMX2X2 U11160 ( .A(\I_cache/cache[3][20] ), .B(n7491), .S0(n3315), .Y(
        n10001) );
  CLKMX2X2 U11161 ( .A(\I_cache/cache[2][20] ), .B(n7491), .S0(n3358), .Y(
        n10002) );
  CLKMX2X2 U11162 ( .A(\I_cache/cache[1][20] ), .B(n7491), .S0(n3225), .Y(
        n10003) );
  CLKMX2X2 U11163 ( .A(\I_cache/cache[0][20] ), .B(n7491), .S0(n3271), .Y(
        n10004) );
  CLKMX2X2 U11164 ( .A(\I_cache/cache[7][19] ), .B(n7120), .S0(n3491), .Y(
        n10005) );
  CLKMX2X2 U11165 ( .A(\I_cache/cache[6][19] ), .B(n7120), .S0(n3535), .Y(
        n10006) );
  CLKMX2X2 U11166 ( .A(\I_cache/cache[5][19] ), .B(n7120), .S0(n3407), .Y(
        n10007) );
  CLKMX2X2 U11167 ( .A(\I_cache/cache[4][19] ), .B(n7120), .S0(n3445), .Y(
        n10008) );
  CLKMX2X2 U11168 ( .A(\I_cache/cache[3][19] ), .B(n7120), .S0(n3313), .Y(
        n10009) );
  CLKMX2X2 U11169 ( .A(\I_cache/cache[2][19] ), .B(n7120), .S0(n3356), .Y(
        n10010) );
  CLKMX2X2 U11170 ( .A(\I_cache/cache[1][19] ), .B(n7120), .S0(n3223), .Y(
        n10011) );
  CLKMX2X2 U11171 ( .A(\I_cache/cache[0][19] ), .B(n7120), .S0(n3268), .Y(
        n10012) );
  CLKMX2X2 U11172 ( .A(\I_cache/cache[7][18] ), .B(n7144), .S0(n3491), .Y(
        n10013) );
  CLKMX2X2 U11173 ( .A(\I_cache/cache[6][18] ), .B(n7144), .S0(n3535), .Y(
        n10014) );
  CLKMX2X2 U11174 ( .A(\I_cache/cache[5][18] ), .B(n7144), .S0(n3404), .Y(
        n10015) );
  CLKMX2X2 U11175 ( .A(\I_cache/cache[4][18] ), .B(n7144), .S0(n3445), .Y(
        n10016) );
  CLKMX2X2 U11176 ( .A(\I_cache/cache[3][18] ), .B(n7144), .S0(n3313), .Y(
        n10017) );
  CLKMX2X2 U11177 ( .A(\I_cache/cache[2][18] ), .B(n7144), .S0(n3356), .Y(
        n10018) );
  CLKMX2X2 U11178 ( .A(\I_cache/cache[1][18] ), .B(n7144), .S0(n3223), .Y(
        n10019) );
  CLKMX2X2 U11179 ( .A(\I_cache/cache[0][18] ), .B(n7144), .S0(n3268), .Y(
        n10020) );
  CLKMX2X2 U11180 ( .A(\I_cache/cache[7][17] ), .B(n4573), .S0(n3490), .Y(
        n10021) );
  CLKMX2X2 U11181 ( .A(\I_cache/cache[6][17] ), .B(n4573), .S0(n3534), .Y(
        n10022) );
  CLKMX2X2 U11182 ( .A(\I_cache/cache[5][17] ), .B(n4573), .S0(n3400), .Y(
        n10023) );
  CLKMX2X2 U11183 ( .A(\I_cache/cache[4][17] ), .B(n4573), .S0(n3444), .Y(
        n10024) );
  CLKMX2X2 U11184 ( .A(\I_cache/cache[3][17] ), .B(n4573), .S0(n3312), .Y(
        n10025) );
  CLKMX2X2 U11185 ( .A(\I_cache/cache[2][17] ), .B(n4573), .S0(n3355), .Y(
        n10026) );
  CLKMX2X2 U11186 ( .A(\I_cache/cache[1][17] ), .B(n4573), .S0(n3222), .Y(
        n10027) );
  CLKMX2X2 U11187 ( .A(\I_cache/cache[0][17] ), .B(n4573), .S0(n3267), .Y(
        n10028) );
  CLKMX2X2 U11188 ( .A(\I_cache/cache[7][16] ), .B(n7096), .S0(n3490), .Y(
        n10029) );
  CLKMX2X2 U11189 ( .A(\I_cache/cache[6][16] ), .B(n7096), .S0(n3534), .Y(
        n10030) );
  CLKMX2X2 U11190 ( .A(\I_cache/cache[5][16] ), .B(n7096), .S0(n3400), .Y(
        n10031) );
  CLKMX2X2 U11191 ( .A(\I_cache/cache[4][16] ), .B(n7096), .S0(n3444), .Y(
        n10032) );
  CLKMX2X2 U11192 ( .A(\I_cache/cache[3][16] ), .B(n7096), .S0(n3312), .Y(
        n10033) );
  CLKMX2X2 U11193 ( .A(\I_cache/cache[2][16] ), .B(n7096), .S0(n3355), .Y(
        n10034) );
  CLKMX2X2 U11194 ( .A(\I_cache/cache[1][16] ), .B(n7096), .S0(n3222), .Y(
        n10035) );
  CLKMX2X2 U11195 ( .A(\I_cache/cache[0][16] ), .B(n7096), .S0(n3267), .Y(
        n10036) );
  CLKMX2X2 U11196 ( .A(\I_cache/cache[7][15] ), .B(n7539), .S0(n3494), .Y(
        n10037) );
  CLKMX2X2 U11197 ( .A(\I_cache/cache[6][15] ), .B(n7539), .S0(n3539), .Y(
        n10038) );
  CLKMX2X2 U11198 ( .A(\I_cache/cache[5][15] ), .B(n7539), .S0(n3404), .Y(
        n10039) );
  CLKMX2X2 U11199 ( .A(\I_cache/cache[4][15] ), .B(n7539), .S0(n3449), .Y(
        n10040) );
  CLKMX2X2 U11200 ( .A(\I_cache/cache[3][15] ), .B(n7539), .S0(n3316), .Y(
        n10041) );
  CLKMX2X2 U11201 ( .A(\I_cache/cache[2][15] ), .B(n7539), .S0(n3359), .Y(
        n10042) );
  CLKMX2X2 U11202 ( .A(\I_cache/cache[1][15] ), .B(n7539), .S0(n3226), .Y(
        n10043) );
  CLKMX2X2 U11203 ( .A(\I_cache/cache[0][15] ), .B(n7539), .S0(n3272), .Y(
        n10044) );
  CLKMX2X2 U11204 ( .A(\I_cache/cache[7][14] ), .B(n7515), .S0(n3493), .Y(
        n10045) );
  CLKMX2X2 U11205 ( .A(\I_cache/cache[6][14] ), .B(n7515), .S0(n3538), .Y(
        n10046) );
  CLKMX2X2 U11206 ( .A(\I_cache/cache[5][14] ), .B(n7515), .S0(n3403), .Y(
        n10047) );
  CLKMX2X2 U11207 ( .A(\I_cache/cache[4][14] ), .B(n7515), .S0(n3448), .Y(
        n10048) );
  CLKMX2X2 U11208 ( .A(\I_cache/cache[3][14] ), .B(n7515), .S0(n3315), .Y(
        n10049) );
  CLKMX2X2 U11209 ( .A(\I_cache/cache[2][14] ), .B(n7515), .S0(n3358), .Y(
        n10050) );
  CLKMX2X2 U11210 ( .A(\I_cache/cache[1][14] ), .B(n7515), .S0(n3225), .Y(
        n10051) );
  CLKMX2X2 U11211 ( .A(\I_cache/cache[0][14] ), .B(n7515), .S0(n3270), .Y(
        n10052) );
  CLKMX2X2 U11212 ( .A(\I_cache/cache[7][13] ), .B(n7564), .S0(n3494), .Y(
        n10053) );
  CLKMX2X2 U11213 ( .A(\I_cache/cache[6][13] ), .B(n7564), .S0(n3539), .Y(
        n10054) );
  CLKMX2X2 U11214 ( .A(\I_cache/cache[5][13] ), .B(n7564), .S0(n3404), .Y(
        n10055) );
  CLKMX2X2 U11215 ( .A(\I_cache/cache[4][13] ), .B(n7564), .S0(n3449), .Y(
        n10056) );
  CLKMX2X2 U11216 ( .A(\I_cache/cache[3][13] ), .B(n7564), .S0(n3316), .Y(
        n10057) );
  CLKMX2X2 U11217 ( .A(\I_cache/cache[2][13] ), .B(n7564), .S0(n3359), .Y(
        n10058) );
  CLKMX2X2 U11218 ( .A(\I_cache/cache[1][13] ), .B(n7564), .S0(n3226), .Y(
        n10059) );
  CLKMX2X2 U11219 ( .A(\I_cache/cache[0][13] ), .B(n7564), .S0(n3272), .Y(
        n10060) );
  CLKMX2X2 U11220 ( .A(\I_cache/cache[7][12] ), .B(n7613), .S0(n3491), .Y(
        n10061) );
  CLKMX2X2 U11221 ( .A(\I_cache/cache[6][12] ), .B(n7613), .S0(n3536), .Y(
        n10062) );
  CLKMX2X2 U11222 ( .A(\I_cache/cache[5][12] ), .B(n7613), .S0(n3401), .Y(
        n10063) );
  CLKMX2X2 U11223 ( .A(\I_cache/cache[4][12] ), .B(n7613), .S0(n3446), .Y(
        n10064) );
  CLKMX2X2 U11224 ( .A(\I_cache/cache[3][12] ), .B(n7613), .S0(n3315), .Y(
        n10065) );
  CLKMX2X2 U11225 ( .A(\I_cache/cache[2][12] ), .B(n7613), .S0(n3357), .Y(
        n10066) );
  CLKMX2X2 U11226 ( .A(\I_cache/cache[1][12] ), .B(n7613), .S0(n3223), .Y(
        n10067) );
  CLKMX2X2 U11227 ( .A(\I_cache/cache[0][12] ), .B(n7613), .S0(n3269), .Y(
        n10068) );
  CLKMX2X2 U11228 ( .A(\I_cache/cache[7][11] ), .B(n7588), .S0(n3494), .Y(
        n10069) );
  CLKMX2X2 U11229 ( .A(\I_cache/cache[6][11] ), .B(n7588), .S0(n3539), .Y(
        n10070) );
  CLKMX2X2 U11230 ( .A(\I_cache/cache[5][11] ), .B(n7588), .S0(n3404), .Y(
        n10071) );
  CLKMX2X2 U11231 ( .A(\I_cache/cache[4][11] ), .B(n7588), .S0(n3449), .Y(
        n10072) );
  CLKMX2X2 U11232 ( .A(\I_cache/cache[3][11] ), .B(n7588), .S0(n3316), .Y(
        n10073) );
  CLKMX2X2 U11233 ( .A(\I_cache/cache[2][11] ), .B(n7588), .S0(n3359), .Y(
        n10074) );
  CLKMX2X2 U11234 ( .A(\I_cache/cache[1][11] ), .B(n7588), .S0(n3226), .Y(
        n10075) );
  CLKMX2X2 U11235 ( .A(\I_cache/cache[0][11] ), .B(n7588), .S0(n3272), .Y(
        n10076) );
  CLKMX2X2 U11236 ( .A(\I_cache/cache[7][10] ), .B(n7666), .S0(n3491), .Y(
        n10077) );
  CLKMX2X2 U11237 ( .A(\I_cache/cache[6][10] ), .B(n7666), .S0(n3536), .Y(
        n10078) );
  CLKMX2X2 U11238 ( .A(\I_cache/cache[5][10] ), .B(n7666), .S0(n3401), .Y(
        n10079) );
  CLKMX2X2 U11239 ( .A(\I_cache/cache[4][10] ), .B(n7666), .S0(n3446), .Y(
        n10080) );
  CLKMX2X2 U11240 ( .A(\I_cache/cache[3][10] ), .B(n7666), .S0(n3317), .Y(
        n10081) );
  CLKMX2X2 U11241 ( .A(\I_cache/cache[2][10] ), .B(n7666), .S0(n3360), .Y(
        n10082) );
  CLKMX2X2 U11242 ( .A(\I_cache/cache[1][10] ), .B(n7666), .S0(n3225), .Y(
        n10083) );
  CLKMX2X2 U11243 ( .A(\I_cache/cache[0][10] ), .B(n7666), .S0(n3269), .Y(
        n10084) );
  CLKMX2X2 U11244 ( .A(\I_cache/cache[7][9] ), .B(n7690), .S0(n3492), .Y(
        n10085) );
  CLKMX2X2 U11245 ( .A(\I_cache/cache[6][9] ), .B(n7690), .S0(n3537), .Y(
        n10086) );
  CLKMX2X2 U11246 ( .A(\I_cache/cache[5][9] ), .B(n7690), .S0(n3402), .Y(
        n10087) );
  CLKMX2X2 U11247 ( .A(\I_cache/cache[4][9] ), .B(n7690), .S0(n3447), .Y(
        n10088) );
  CLKMX2X2 U11248 ( .A(\I_cache/cache[3][9] ), .B(n7690), .S0(n3314), .Y(
        n10089) );
  CLKMX2X2 U11249 ( .A(\I_cache/cache[2][9] ), .B(n7690), .S0(n3357), .Y(
        n10090) );
  CLKMX2X2 U11250 ( .A(\I_cache/cache[1][9] ), .B(n7690), .S0(n3224), .Y(
        n10091) );
  CLKMX2X2 U11251 ( .A(\I_cache/cache[0][9] ), .B(n7690), .S0(n3270), .Y(
        n10092) );
  CLKMX2X2 U11252 ( .A(\I_cache/cache[7][8] ), .B(n7713), .S0(n3492), .Y(
        n10093) );
  CLKMX2X2 U11253 ( .A(\I_cache/cache[6][8] ), .B(n7713), .S0(n3537), .Y(
        n10094) );
  CLKMX2X2 U11254 ( .A(\I_cache/cache[5][8] ), .B(n7713), .S0(n3402), .Y(
        n10095) );
  CLKMX2X2 U11255 ( .A(\I_cache/cache[4][8] ), .B(n7713), .S0(n3447), .Y(
        n10096) );
  CLKMX2X2 U11256 ( .A(\I_cache/cache[3][8] ), .B(n7713), .S0(n3314), .Y(
        n10097) );
  CLKMX2X2 U11257 ( .A(\I_cache/cache[2][8] ), .B(n7713), .S0(n3357), .Y(
        n10098) );
  CLKMX2X2 U11258 ( .A(\I_cache/cache[1][8] ), .B(n7713), .S0(n3224), .Y(
        n10099) );
  CLKMX2X2 U11259 ( .A(\I_cache/cache[0][8] ), .B(n7713), .S0(n3270), .Y(
        n10100) );
  CLKMX2X2 U11260 ( .A(\I_cache/cache[7][7] ), .B(n7739), .S0(n3492), .Y(
        n10101) );
  CLKMX2X2 U11261 ( .A(\I_cache/cache[6][7] ), .B(n7739), .S0(n3537), .Y(
        n10102) );
  CLKMX2X2 U11262 ( .A(\I_cache/cache[5][7] ), .B(n7739), .S0(n3402), .Y(
        n10103) );
  CLKMX2X2 U11263 ( .A(\I_cache/cache[4][7] ), .B(n7739), .S0(n3447), .Y(
        n10104) );
  CLKMX2X2 U11264 ( .A(\I_cache/cache[3][7] ), .B(n7739), .S0(n3314), .Y(
        n10105) );
  CLKMX2X2 U11265 ( .A(\I_cache/cache[2][7] ), .B(n7739), .S0(n3357), .Y(
        n10106) );
  CLKMX2X2 U11266 ( .A(\I_cache/cache[1][7] ), .B(n7739), .S0(n3224), .Y(
        n10107) );
  CLKMX2X2 U11267 ( .A(\I_cache/cache[0][7] ), .B(n7739), .S0(n3270), .Y(
        n10108) );
  CLKMX2X2 U11268 ( .A(\I_cache/cache[7][6] ), .B(n7763), .S0(n3495), .Y(
        n10109) );
  CLKMX2X2 U11269 ( .A(\I_cache/cache[6][6] ), .B(n7763), .S0(n3536), .Y(
        n10110) );
  CLKMX2X2 U11270 ( .A(\I_cache/cache[5][6] ), .B(n7763), .S0(n3401), .Y(
        n10111) );
  CLKMX2X2 U11271 ( .A(\I_cache/cache[4][6] ), .B(n7763), .S0(n3446), .Y(
        n10112) );
  CLKMX2X2 U11272 ( .A(\I_cache/cache[3][6] ), .B(n7763), .S0(n3316), .Y(
        n10113) );
  CLKMX2X2 U11273 ( .A(\I_cache/cache[2][6] ), .B(n7763), .S0(n3357), .Y(
        n10114) );
  CLKMX2X2 U11274 ( .A(\I_cache/cache[1][6] ), .B(n7763), .S0(n3229), .Y(
        n10115) );
  CLKMX2X2 U11275 ( .A(\I_cache/cache[0][6] ), .B(n7763), .S0(n3274), .Y(
        n10116) );
  CLKMX2X2 U11276 ( .A(\I_cache/cache[7][5] ), .B(n7391), .S0(n3489), .Y(
        n10117) );
  CLKMX2X2 U11277 ( .A(\I_cache/cache[6][5] ), .B(n7391), .S0(n3533), .Y(
        n10118) );
  CLKMX2X2 U11278 ( .A(\I_cache/cache[5][5] ), .B(n7391), .S0(n3399), .Y(
        n10119) );
  CLKMX2X2 U11279 ( .A(\I_cache/cache[4][5] ), .B(n7391), .S0(n3450), .Y(
        n10120) );
  CLKMX2X2 U11280 ( .A(\I_cache/cache[3][5] ), .B(n7391), .S0(n3311), .Y(
        n10121) );
  CLKMX2X2 U11281 ( .A(\I_cache/cache[2][5] ), .B(n7391), .S0(n3354), .Y(
        n10122) );
  CLKMX2X2 U11282 ( .A(\I_cache/cache[1][5] ), .B(n7391), .S0(n3221), .Y(
        n10123) );
  CLKMX2X2 U11283 ( .A(\I_cache/cache[0][5] ), .B(n7391), .S0(n3266), .Y(
        n10124) );
  CLKMX2X2 U11284 ( .A(\I_cache/cache[7][4] ), .B(n4548), .S0(n3495), .Y(
        n10125) );
  CLKMX2X2 U11285 ( .A(\I_cache/cache[6][4] ), .B(n4548), .S0(n3537), .Y(
        n10126) );
  CLKMX2X2 U11286 ( .A(\I_cache/cache[5][4] ), .B(n4548), .S0(n3400), .Y(
        n10127) );
  CLKMX2X2 U11287 ( .A(\I_cache/cache[4][4] ), .B(n4548), .S0(n3450), .Y(
        n10128) );
  CLKMX2X2 U11288 ( .A(\I_cache/cache[3][4] ), .B(n4548), .S0(n3317), .Y(
        n10129) );
  CLKMX2X2 U11289 ( .A(\I_cache/cache[2][4] ), .B(n4548), .S0(n3360), .Y(
        n10130) );
  CLKMX2X2 U11290 ( .A(\I_cache/cache[1][4] ), .B(n4548), .S0(n3222), .Y(
        n10131) );
  CLKMX2X2 U11291 ( .A(\I_cache/cache[0][4] ), .B(n4548), .S0(n3267), .Y(
        n10132) );
  CLKMX2X2 U11292 ( .A(\I_cache/cache[7][3] ), .B(n8363), .S0(n3497), .Y(
        n10133) );
  CLKMX2X2 U11293 ( .A(\I_cache/cache[6][3] ), .B(n8363), .S0(n3541), .Y(
        n10134) );
  CLKMX2X2 U11294 ( .A(\I_cache/cache[5][3] ), .B(n8363), .S0(n3406), .Y(
        n10135) );
  CLKMX2X2 U11295 ( .A(\I_cache/cache[4][3] ), .B(n8363), .S0(n3452), .Y(
        n10136) );
  CLKMX2X2 U11296 ( .A(\I_cache/cache[3][3] ), .B(n8363), .S0(n3319), .Y(
        n10137) );
  CLKMX2X2 U11297 ( .A(\I_cache/cache[2][3] ), .B(n8363), .S0(n3362), .Y(
        n10138) );
  CLKMX2X2 U11298 ( .A(\I_cache/cache[1][3] ), .B(n8363), .S0(n3227), .Y(
        n10139) );
  CLKMX2X2 U11299 ( .A(\I_cache/cache[0][3] ), .B(n8363), .S0(n3267), .Y(
        n10140) );
  CLKMX2X2 U11300 ( .A(\I_cache/cache[7][2] ), .B(n8377), .S0(n3497), .Y(
        n10141) );
  CLKMX2X2 U11301 ( .A(\I_cache/cache[6][2] ), .B(n8377), .S0(n3533), .Y(
        n10142) );
  CLKMX2X2 U11302 ( .A(\I_cache/cache[5][2] ), .B(n8377), .S0(n3407), .Y(
        n10143) );
  CLKMX2X2 U11303 ( .A(\I_cache/cache[4][2] ), .B(n8377), .S0(n3446), .Y(
        n10144) );
  CLKMX2X2 U11304 ( .A(\I_cache/cache[3][2] ), .B(n8377), .S0(n3313), .Y(
        n10145) );
  CLKMX2X2 U11305 ( .A(\I_cache/cache[2][2] ), .B(n8377), .S0(n3355), .Y(
        n10146) );
  CLKMX2X2 U11306 ( .A(\I_cache/cache[1][2] ), .B(n8377), .S0(n3223), .Y(
        n10147) );
  CLKMX2X2 U11307 ( .A(\I_cache/cache[0][2] ), .B(n8377), .S0(n3274), .Y(
        n10148) );
  CLKMX2X2 U11308 ( .A(\I_cache/cache[7][1] ), .B(n4553), .S0(n3490), .Y(
        n10149) );
  CLKMX2X2 U11309 ( .A(\I_cache/cache[6][1] ), .B(n4553), .S0(n3534), .Y(
        n10150) );
  CLKMX2X2 U11310 ( .A(\I_cache/cache[5][1] ), .B(n4553), .S0(n3400), .Y(
        n10151) );
  CLKMX2X2 U11311 ( .A(\I_cache/cache[4][1] ), .B(n4553), .S0(n3444), .Y(
        n10152) );
  CLKMX2X2 U11312 ( .A(\I_cache/cache[3][1] ), .B(n4553), .S0(n3312), .Y(
        n10153) );
  CLKMX2X2 U11313 ( .A(\I_cache/cache[2][1] ), .B(n4553), .S0(n3355), .Y(
        n10154) );
  CLKMX2X2 U11314 ( .A(\I_cache/cache[1][1] ), .B(n4553), .S0(n3222), .Y(
        n10155) );
  CLKMX2X2 U11315 ( .A(\I_cache/cache[0][1] ), .B(n4553), .S0(n3267), .Y(
        n10156) );
  CLKINVX1 U11316 ( .A(\i_MIPS/n297 ), .Y(n7802) );
  AO22X1 U11317 ( .A0(n13), .A1(n7314), .B0(n3630), .B1(\i_MIPS/ALUOp[0] ), 
        .Y(\i_MIPS/n472 ) );
  OAI31XL U11318 ( .A0(n7313), .A1(\i_MIPS/IR_ID[30] ), .A2(\i_MIPS/IR_ID[27] ), .B0(\i_MIPS/Control_ID/n15 ), .Y(n7314) );
  AO22X1 U11319 ( .A0(\i_MIPS/control_out[0] ), .A1(n3614), .B0(n3629), .B1(
        \i_MIPS/ID_EX_0 ), .Y(\i_MIPS/n528 ) );
  NAND3BX1 U11320 ( .AN(\i_MIPS/control_out[7] ), .B(n3688), .C(
        \i_MIPS/Control_ID/n12 ), .Y(\i_MIPS/control_out[0] ) );
  AO21X1 U11321 ( .A0(\i_MIPS/ID_EX[88] ), .A1(n3629), .B0(n2804), .Y(
        \i_MIPS/n497 ) );
  AO21X1 U11322 ( .A0(\i_MIPS/ID_EX[104] ), .A1(n3628), .B0(n2804), .Y(
        \i_MIPS/n481 ) );
  AO21X1 U11323 ( .A0(n3629), .A1(n1893), .B0(n8455), .Y(\i_MIPS/n527 ) );
  AO21X1 U11324 ( .A0(n3628), .A1(\i_MIPS/ID_EX_3 ), .B0(n8455), .Y(
        \i_MIPS/n525 ) );
  AO21X1 U11325 ( .A0(n3629), .A1(n1894), .B0(n2803), .Y(\i_MIPS/n480 ) );
  AND3X2 U11326 ( .A(\i_MIPS/Register/n120 ), .B(\i_MIPS/Reg_W[3] ), .C(
        \i_MIPS/Reg_W[4] ), .Y(\i_MIPS/Register/n104 ) );
  AO22X2 U11327 ( .A0(n3603), .A1(ICACHE_addr[29]), .B0(n3601), .B1(n8712), 
        .Y(n8449) );
  AO22X2 U11328 ( .A0(n3609), .A1(ICACHE_addr[25]), .B0(n3601), .B1(n8708), 
        .Y(n8443) );
  AO22X2 U11329 ( .A0(n3603), .A1(ICACHE_addr[20]), .B0(n3600), .B1(n8703), 
        .Y(n8430) );
  NOR2BX1 U11330 ( .AN(\i_MIPS/EX_MEM_0 ), .B(\i_MIPS/EX_MEM_74 ), .Y(
        \i_MIPS/Register/n120 ) );
  NAND3BX1 U11331 ( .AN(\i_MIPS/IR_ID[29] ), .B(\i_MIPS/n326 ), .C(
        \i_MIPS/n330 ), .Y(n7305) );
  OAI2BB2XL U11332 ( .B0(\D_cache/n205 ), .B1(n3784), .A0N(
        \D_cache/cache[7][154] ), .A1N(n3797), .Y(\D_cache/n557 ) );
  OAI2BB2XL U11333 ( .B0(\D_cache/n205 ), .B1(n3804), .A0N(
        \D_cache/cache[6][154] ), .A1N(n3817), .Y(\D_cache/n558 ) );
  OAI2BB2XL U11334 ( .B0(\D_cache/n205 ), .B1(n3830), .A0N(
        \D_cache/cache[5][154] ), .A1N(n3835), .Y(\D_cache/n559 ) );
  OAI2BB2XL U11335 ( .B0(\D_cache/n205 ), .B1(n3852), .A0N(
        \D_cache/cache[4][154] ), .A1N(n3857), .Y(\D_cache/n560 ) );
  OAI2BB2XL U11336 ( .B0(\D_cache/n205 ), .B1(n3869), .A0N(
        \D_cache/cache[3][154] ), .A1N(n3876), .Y(\D_cache/n561 ) );
  OAI2BB2XL U11337 ( .B0(\D_cache/n205 ), .B1(n3884), .A0N(
        \D_cache/cache[2][154] ), .A1N(n3897), .Y(\D_cache/n562 ) );
  OAI2BB2XL U11338 ( .B0(\D_cache/n205 ), .B1(n3904), .A0N(
        \D_cache/cache[1][154] ), .A1N(n3918), .Y(\D_cache/n563 ) );
  OAI2BB2XL U11339 ( .B0(\D_cache/n205 ), .B1(n3927), .A0N(
        \D_cache/cache[0][154] ), .A1N(n3939), .Y(\D_cache/n564 ) );
  NOR3X1 U11340 ( .A(\i_MIPS/Hazard_detection/n8 ), .B(
        \i_MIPS/Hazard_detection/n9 ), .C(\i_MIPS/Hazard_detection/n10 ), .Y(
        \i_MIPS/Hazard_detection/n7 ) );
  NOR3X1 U11341 ( .A(\i_MIPS/Hazard_detection/n11 ), .B(
        \i_MIPS/Hazard_detection/n12 ), .C(\i_MIPS/Hazard_detection/n13 ), .Y(
        \i_MIPS/Hazard_detection/n4 ) );
  AND2X2 U11342 ( .A(\i_MIPS/IR_ID[27] ), .B(\i_MIPS/IR_ID[26] ), .Y(n2995) );
  NOR2X1 U11343 ( .A(n7077), .B(n7076), .Y(n7833) );
  OR2X1 U11344 ( .A(\i_MIPS/Sign_Extend_ID[4] ), .B(\i_MIPS/Sign_Extend_ID[2] ), .Y(n7076) );
  NAND4X1 U11345 ( .A(\i_MIPS/Sign_Extend_ID[3] ), .B(n7075), .C(n7074), .D(
        \i_MIPS/n213 ), .Y(n7077) );
  CLKINVX1 U11346 ( .A(mem_ready_D), .Y(n8772) );
  CLKBUFX3 U11347 ( .A(\i_MIPS/IR_ID[25] ), .Y(n4012) );
  CLKMX2X2 U11348 ( .A(\I_cache/cache[7][153] ), .B(n8394), .S0(n3488), .Y(
        n8933) );
  CLKMX2X2 U11349 ( .A(\I_cache/cache[6][153] ), .B(n8394), .S0(n3534), .Y(
        n8934) );
  CLKMX2X2 U11350 ( .A(\I_cache/cache[5][153] ), .B(n8394), .S0(n3407), .Y(
        n8935) );
  CLKMX2X2 U11351 ( .A(\I_cache/cache[4][153] ), .B(n8394), .S0(n3452), .Y(
        n8936) );
  CLKMX2X2 U11352 ( .A(\I_cache/cache[3][153] ), .B(n8394), .S0(n3319), .Y(
        n8937) );
  CLKMX2X2 U11353 ( .A(\I_cache/cache[2][153] ), .B(n8394), .S0(n3356), .Y(
        n8938) );
  CLKMX2X2 U11354 ( .A(\I_cache/cache[1][153] ), .B(n8394), .S0(n3229), .Y(
        n8939) );
  CLKMX2X2 U11355 ( .A(\I_cache/cache[0][153] ), .B(n8394), .S0(n3265), .Y(
        n8940) );
  CLKBUFX3 U11356 ( .A(mem_ready_I), .Y(n3051) );
  AND3X2 U11357 ( .A(\i_MIPS/Register/n120 ), .B(n2996), .C(\i_MIPS/Reg_W[3] ), 
        .Y(\i_MIPS/Register/n131 ) );
  AND3X2 U11358 ( .A(\i_MIPS/Register/n120 ), .B(n2997), .C(\i_MIPS/Reg_W[4] ), 
        .Y(\i_MIPS/Register/n122 ) );
  NAND3BX1 U11359 ( .AN(n7311), .B(\i_MIPS/IR_ID[29] ), .C(n7310), .Y(
        \i_MIPS/Control_ID/n15 ) );
  AOI2BB1X1 U11360 ( .A0N(\i_MIPS/n322 ), .A1N(\i_MIPS/n332 ), .B0(
        \i_MIPS/IR_ID[30] ), .Y(n7310) );
  XOR2X1 U11361 ( .A(n7309), .B(n7308), .Y(n7311) );
  NAND2X1 U11362 ( .A(\i_MIPS/IR_ID[28] ), .B(\i_MIPS/n324 ), .Y(n7309) );
  NAND2X1 U11363 ( .A(n2882), .B(\i_MIPS/IR_ID[31] ), .Y(
        \i_MIPS/Control_ID/n12 ) );
  NAND2X1 U11364 ( .A(\i_MIPS/IF_ID[64] ), .B(\i_MIPS/IF_ID[97] ), .Y(n7081)
         );
  NOR2X1 U11365 ( .A(\i_MIPS/Sign_Extend_ID[5] ), .B(
        \i_MIPS/Sign_Extend_ID[0] ), .Y(n7074) );
  OAI222XL U11366 ( .A0(n3070), .A1(n4971), .B0(n6402), .B1(n6677), .C0(n6341), 
        .C1(n5548), .Y(n4922) );
  AO22X2 U11367 ( .A0(n3609), .A1(ICACHE_addr[7]), .B0(n3600), .B1(n8690), .Y(
        n8433) );
  AOI2BB1X1 U11368 ( .A0N(n3078), .A1N(n6610), .B0(n5108), .Y(n5109) );
  OA22X1 U11369 ( .A0(n5046), .A1(n6610), .B0(n5045), .B1(n5044), .Y(n5058) );
  CLKINVX1 U11370 ( .A(n6610), .Y(n5402) );
  NAND2BX1 U11371 ( .AN(n3577), .B(n8286), .Y(n8292) );
  AO22X2 U11372 ( .A0(n3602), .A1(ICACHE_addr[8]), .B0(n3600), .B1(n8691), .Y(
        n8432) );
  XNOR2X1 U11373 ( .A(ICACHE_addr[8]), .B(n8691), .Y(n4428) );
  AO22X2 U11374 ( .A0(n3609), .A1(ICACHE_addr[23]), .B0(n3600), .B1(n8706), 
        .Y(n8434) );
  NAND2X1 U11375 ( .A(n3579), .B(n8042), .Y(n8062) );
  AO22X2 U11376 ( .A0(n3609), .A1(ICACHE_addr[22]), .B0(n3600), .B1(n8705), 
        .Y(n8436) );
  XNOR2X1 U11377 ( .A(ICACHE_addr[22]), .B(n8705), .Y(n4461) );
  NAND2X1 U11378 ( .A(n4972), .B(n4971), .Y(n4905) );
  AO22X2 U11379 ( .A0(n3609), .A1(ICACHE_addr[27]), .B0(n3600), .B1(n8710), 
        .Y(n8435) );
  AO22X2 U11380 ( .A0(n3609), .A1(ICACHE_addr[24]), .B0(n3601), .B1(n8707), 
        .Y(n8442) );
  AO22X2 U11381 ( .A0(n3606), .A1(ICACHE_addr[18]), .B0(n3600), .B1(n8701), 
        .Y(n8429) );
  AO22X2 U11382 ( .A0(n3609), .A1(ICACHE_addr[11]), .B0(n3600), .B1(n8694), 
        .Y(n8439) );
  INVX2 U11383 ( .A(n21), .Y(n5986) );
  AO22X2 U11384 ( .A0(n3609), .A1(ICACHE_addr[26]), .B0(n3601), .B1(n8709), 
        .Y(n8441) );
  NAND4XL U11385 ( .A(n4725), .B(n5048), .C(n4724), .D(n4726), .Y(n7004) );
  AO22X2 U11386 ( .A0(n3607), .A1(ICACHE_addr[5]), .B0(n3601), .B1(n8688), .Y(
        n8448) );
  AO22X2 U11387 ( .A0(n3609), .A1(ICACHE_addr[12]), .B0(n3601), .B1(n8695), 
        .Y(n8445) );
  AO22X2 U11388 ( .A0(n3608), .A1(ICACHE_addr[6]), .B0(n3600), .B1(n8689), .Y(
        n8431) );
  AO22X2 U11389 ( .A0(n3602), .A1(ICACHE_addr[19]), .B0(n3600), .B1(n8702), 
        .Y(n8428) );
  AO22X2 U11390 ( .A0(n3609), .A1(ICACHE_addr[10]), .B0(n3600), .B1(n8693), 
        .Y(n8438) );
  AO22X2 U11391 ( .A0(n3608), .A1(ICACHE_addr[28]), .B0(n3601), .B1(n8711), 
        .Y(n8447) );
  AO22X2 U11392 ( .A0(n3607), .A1(ICACHE_addr[21]), .B0(n3601), .B1(n8704), 
        .Y(n8451) );
  AO22X2 U11393 ( .A0(n3609), .A1(ICACHE_addr[14]), .B0(n3601), .B1(n8697), 
        .Y(n8444) );
  AO22X2 U11394 ( .A0(n3609), .A1(ICACHE_addr[9]), .B0(n3601), .B1(n8692), .Y(
        n8440) );
  AO22X2 U11395 ( .A0(n3607), .A1(ICACHE_addr[13]), .B0(n3601), .B1(n8696), 
        .Y(n8446) );
  AO22X2 U11396 ( .A0(n3609), .A1(ICACHE_addr[15]), .B0(n3600), .B1(n8698), 
        .Y(n8437) );
  BUFX16 U11397 ( .A(n10312), .Y(DCACHE_addr[14]) );
  MX2XL U11398 ( .A(DCACHE_addr[13]), .B(n8253), .S0(n3626), .Y(\i_MIPS/n454 )
         );
  BUFX16 U11399 ( .A(n10314), .Y(DCACHE_addr[12]) );
  OA22X2 U11400 ( .A0(n3547), .A1(n139), .B0(n3506), .B1(n1029), .Y(n4476) );
  OA22X2 U11401 ( .A0(n3548), .A1(n140), .B0(n3507), .B1(n1030), .Y(n4508) );
  NAND2XL U11402 ( .A(n3579), .B(n8301), .Y(n8322) );
  MX2XL U11403 ( .A(DCACHE_addr[16]), .B(n7977), .S0(n3624), .Y(\i_MIPS/n451 )
         );
  MX2XL U11404 ( .A(DCACHE_addr[5]), .B(n8009), .S0(n3626), .Y(\i_MIPS/n462 )
         );
  AND3X2 U11405 ( .A(n4975), .B(n3076), .C(n6614), .Y(n4976) );
  NAND2X1 U11406 ( .A(n6614), .B(n2826), .Y(n6625) );
  BUFX16 U11407 ( .A(n10306), .Y(DCACHE_addr[20]) );
  BUFX16 U11408 ( .A(n10319), .Y(DCACHE_addr[7]) );
  BUFX16 U11409 ( .A(n10304), .Y(DCACHE_addr[22]) );
  BUFX16 U11410 ( .A(n10308), .Y(DCACHE_addr[18]) );
  BUFX16 U11411 ( .A(n10320), .Y(DCACHE_addr[6]) );
  BUFX16 U11412 ( .A(n10299), .Y(DCACHE_addr[27]) );
  BUFX16 U11413 ( .A(n10307), .Y(DCACHE_addr[19]) );
  CLKBUFX3 U11414 ( .A(\D_cache/n314 ), .Y(n3010) );
  BUFX16 U11415 ( .A(n10318), .Y(DCACHE_addr[8]) );
  BUFX16 U11416 ( .A(n10303), .Y(DCACHE_addr[23]) );
  BUFX16 U11417 ( .A(n10317), .Y(DCACHE_addr[9]) );
  NAND2XL U11418 ( .A(n5107), .B(n5106), .Y(n5110) );
  BUFX16 U11419 ( .A(n10311), .Y(DCACHE_addr[15]) );
  INVX12 U11420 ( .A(n1621), .Y(DCACHE_addr[11]) );
  MX2XL U11421 ( .A(DCACHE_addr[9]), .B(n8246), .S0(n3626), .Y(\i_MIPS/n458 )
         );
  MX2XL U11422 ( .A(\i_MIPS/ID_EX[50] ), .B(n7805), .S0(n3625), .Y(
        \i_MIPS/n419 ) );
  CLKBUFX2 U11423 ( .A(n8728), .Y(n3657) );
  OAI2BB2XL U11424 ( .B0(n3652), .B1(n3694), .A0N(
        \i_MIPS/Register/register[29][0] ), .A1N(n3694), .Y(
        \i_MIPS/Register/n180 ) );
  OAI2BB2XL U11425 ( .B0(n3652), .B1(n3697), .A0N(
        \i_MIPS/Register/register[28][0] ), .A1N(n3697), .Y(
        \i_MIPS/Register/n212 ) );
  OAI2BB2XL U11426 ( .B0(n3652), .B1(n3700), .A0N(
        \i_MIPS/Register/register[27][0] ), .A1N(n3700), .Y(
        \i_MIPS/Register/n244 ) );
  OAI2BB2XL U11427 ( .B0(n3652), .B1(n3703), .A0N(
        \i_MIPS/Register/register[26][0] ), .A1N(n3703), .Y(
        \i_MIPS/Register/n276 ) );
  OAI2BB2XL U11428 ( .B0(n3652), .B1(n3706), .A0N(
        \i_MIPS/Register/register[25][0] ), .A1N(n3706), .Y(
        \i_MIPS/Register/n308 ) );
  OAI2BB2XL U11429 ( .B0(n3652), .B1(n3709), .A0N(
        \i_MIPS/Register/register[24][0] ), .A1N(n3709), .Y(
        \i_MIPS/Register/n340 ) );
  OAI2BB2XL U11430 ( .B0(n3652), .B1(n3712), .A0N(
        \i_MIPS/Register/register[23][0] ), .A1N(n3711), .Y(
        \i_MIPS/Register/n372 ) );
  OAI2BB2XL U11431 ( .B0(n3652), .B1(n3715), .A0N(
        \i_MIPS/Register/register[22][0] ), .A1N(n3714), .Y(
        \i_MIPS/Register/n404 ) );
  OAI2BB2XL U11432 ( .B0(n3652), .B1(n3718), .A0N(
        \i_MIPS/Register/register[21][0] ), .A1N(n3718), .Y(
        \i_MIPS/Register/n436 ) );
  OAI2BB2XL U11433 ( .B0(n3652), .B1(n3721), .A0N(
        \i_MIPS/Register/register[20][0] ), .A1N(n3720), .Y(
        \i_MIPS/Register/n468 ) );
  OAI2BB2XL U11434 ( .B0(n3652), .B1(n3724), .A0N(
        \i_MIPS/Register/register[19][0] ), .A1N(n3724), .Y(
        \i_MIPS/Register/n500 ) );
  OAI2BB2XL U11435 ( .B0(n3652), .B1(n3727), .A0N(
        \i_MIPS/Register/register[18][0] ), .A1N(n3726), .Y(
        \i_MIPS/Register/n532 ) );
  OAI2BB2XL U11436 ( .B0(n3653), .B1(n3730), .A0N(
        \i_MIPS/Register/register[17][0] ), .A1N(n3730), .Y(
        \i_MIPS/Register/n564 ) );
  OAI2BB2XL U11437 ( .B0(n3653), .B1(n3733), .A0N(
        \i_MIPS/Register/register[16][0] ), .A1N(n3733), .Y(
        \i_MIPS/Register/n596 ) );
  OAI2BB2XL U11438 ( .B0(n3653), .B1(n3736), .A0N(
        \i_MIPS/Register/register[15][0] ), .A1N(n3736), .Y(
        \i_MIPS/Register/n628 ) );
  OAI2BB2XL U11439 ( .B0(n3653), .B1(n3739), .A0N(
        \i_MIPS/Register/register[14][0] ), .A1N(n3739), .Y(
        \i_MIPS/Register/n660 ) );
  OAI2BB2XL U11440 ( .B0(n3653), .B1(n3691), .A0N(
        \i_MIPS/Register/register[30][0] ), .A1N(n3690), .Y(
        \i_MIPS/Register/n148 ) );
  OAI2BB2XL U11441 ( .B0(n3653), .B1(n3742), .A0N(
        \i_MIPS/Register/register[13][0] ), .A1N(n3741), .Y(
        \i_MIPS/Register/n692 ) );
  OAI2BB2XL U11442 ( .B0(n3653), .B1(n3745), .A0N(
        \i_MIPS/Register/register[12][0] ), .A1N(n3745), .Y(
        \i_MIPS/Register/n724 ) );
  OAI2BB2XL U11443 ( .B0(n3653), .B1(n3748), .A0N(
        \i_MIPS/Register/register[11][0] ), .A1N(n3747), .Y(
        \i_MIPS/Register/n756 ) );
  OAI2BB2XL U11444 ( .B0(n3653), .B1(n3751), .A0N(
        \i_MIPS/Register/register[10][0] ), .A1N(n3751), .Y(
        \i_MIPS/Register/n788 ) );
  OAI2BB2XL U11445 ( .B0(n3653), .B1(n3754), .A0N(
        \i_MIPS/Register/register[9][0] ), .A1N(n3753), .Y(
        \i_MIPS/Register/n820 ) );
  OAI2BB2XL U11446 ( .B0(n3653), .B1(n3757), .A0N(
        \i_MIPS/Register/register[8][0] ), .A1N(n3756), .Y(
        \i_MIPS/Register/n852 ) );
  OAI2BB2XL U11447 ( .B0(n3653), .B1(n3760), .A0N(
        \i_MIPS/Register/register[7][0] ), .A1N(n3759), .Y(
        \i_MIPS/Register/n884 ) );
  OAI2BB2XL U11448 ( .B0(n3654), .B1(n3763), .A0N(
        \i_MIPS/Register/register[6][0] ), .A1N(n3763), .Y(
        \i_MIPS/Register/n916 ) );
  OAI2BB2XL U11449 ( .B0(n3654), .B1(n3766), .A0N(
        \i_MIPS/Register/register[5][0] ), .A1N(n3766), .Y(
        \i_MIPS/Register/n948 ) );
  OAI2BB2XL U11450 ( .B0(n3654), .B1(n3769), .A0N(
        \i_MIPS/Register/register[4][0] ), .A1N(n3769), .Y(
        \i_MIPS/Register/n980 ) );
  OAI2BB2XL U11451 ( .B0(n3654), .B1(n3772), .A0N(
        \i_MIPS/Register/register[3][0] ), .A1N(n3772), .Y(
        \i_MIPS/Register/n1012 ) );
  OAI2BB2XL U11452 ( .B0(n3654), .B1(n3775), .A0N(
        \i_MIPS/Register/register[2][0] ), .A1N(n3775), .Y(
        \i_MIPS/Register/n1044 ) );
  OAI2BB2XL U11453 ( .B0(n3654), .B1(n3778), .A0N(
        \i_MIPS/Register/register[1][0] ), .A1N(n3778), .Y(
        \i_MIPS/Register/n1076 ) );
  OAI2BB2XL U11454 ( .B0(n3654), .B1(n3781), .A0N(
        \i_MIPS/Register/register[0][0] ), .A1N(n3781), .Y(
        \i_MIPS/Register/n1108 ) );
  OAI222XL U11455 ( .A0(n8334), .A1(n70), .B0(n3654), .B1(n8333), .C0(n3688), 
        .C1(\i_MIPS/n180 ), .Y(n8804) );
  CLKBUFX2 U11456 ( .A(n8723), .Y(n3645) );
  OAI222XL U11457 ( .A0(n6971), .A1(n7071), .B0(n6949), .B1(n3217), .C0(n3657), 
        .C1(n3214), .Y(n3021) );
  NAND2X2 U11458 ( .A(n3010), .B(\D_cache/n519 ), .Y(\D_cache/n454 ) );
  NAND2X2 U11459 ( .A(n3010), .B(\D_cache/n383 ), .Y(\D_cache/n319 ) );
  CLKBUFX2 U11460 ( .A(n8724), .Y(n3646) );
  AOI221X4 U11461 ( .A0(\D_cache/N98 ), .A1(n3026), .B0(\D_cache/N66 ), .B1(
        n3023), .C0(n3024), .Y(n3022) );
  MX2XL U11462 ( .A(n1883), .B(n7812), .S0(n3626), .Y(\i_MIPS/n409 ) );
  CLKBUFX2 U11463 ( .A(n8737), .Y(n3672) );
  AOI2BB2X2 U11464 ( .B0(\D_cache/N149 ), .B1(n2153), .A0N(n23), .A1N(n8899), 
        .Y(\D_cache/n174 ) );
  AOI2BB2X1 U11465 ( .B0(\D_cache/N133 ), .B1(n2153), .A0N(n24), .A1N(n8883), 
        .Y(\D_cache/n189 ) );
  AOI2BB2X2 U11466 ( .B0(\D_cache/N151 ), .B1(n2153), .A0N(n3040), .A1N(n8901), 
        .Y(\D_cache/n188 ) );
  CLKBUFX2 U11467 ( .A(n8731), .Y(n3661) );
  MXI2XL U11468 ( .A(n2219), .B(DCACHE_rdata[5]), .S0(n4021), .Y(n8741) );
  CLKBUFX2 U11469 ( .A(n8735), .Y(n3668) );
  AOI2BB2X2 U11470 ( .B0(\D_cache/N123 ), .B1(n2153), .A0N(n23), .A1N(n8873), 
        .Y(\D_cache/n178 ) );
  AOI2BB2X2 U11471 ( .B0(\D_cache/N127 ), .B1(n2153), .A0N(n24), .A1N(n8877), 
        .Y(\D_cache/n182 ) );
  MX2XL U11472 ( .A(DCACHE_addr[6]), .B(n8231), .S0(n3625), .Y(\i_MIPS/n461 )
         );
  INVXL U11473 ( .A(n8241), .Y(n8338) );
  NAND3BX4 U11474 ( .AN(n4702), .B(n6064), .C(n4701), .Y(n6765) );
  OAI222XL U11475 ( .A0(n5598), .A1(n3164), .B0(n5576), .B1(n2761), .C0(n3646), 
        .C1(n3163), .Y(n3028) );
  INVXL U11476 ( .A(n2748), .Y(n3029) );
  INVX3 U11477 ( .A(n3029), .Y(n3030) );
  CLKBUFX2 U11478 ( .A(n8734), .Y(n3667) );
  CLKBUFX2 U11479 ( .A(n8717), .Y(n3636) );
  CLKBUFX2 U11480 ( .A(n8739), .Y(n3676) );
  OAI2BB2XL U11481 ( .B0(n3662), .B1(n3693), .A0N(
        \i_MIPS/Register/register[29][1] ), .A1N(n3693), .Y(
        \i_MIPS/Register/n181 ) );
  OAI2BB2XL U11482 ( .B0(n3662), .B1(n3696), .A0N(
        \i_MIPS/Register/register[28][1] ), .A1N(n3696), .Y(
        \i_MIPS/Register/n213 ) );
  OAI2BB2XL U11483 ( .B0(n3662), .B1(n3699), .A0N(
        \i_MIPS/Register/register[27][1] ), .A1N(n3699), .Y(
        \i_MIPS/Register/n245 ) );
  OAI2BB2XL U11484 ( .B0(n8732), .B1(n3702), .A0N(
        \i_MIPS/Register/register[26][1] ), .A1N(n3702), .Y(
        \i_MIPS/Register/n277 ) );
  OAI2BB2XL U11485 ( .B0(n3662), .B1(n3705), .A0N(
        \i_MIPS/Register/register[25][1] ), .A1N(n3705), .Y(
        \i_MIPS/Register/n309 ) );
  OAI2BB2XL U11486 ( .B0(n3662), .B1(n3708), .A0N(
        \i_MIPS/Register/register[24][1] ), .A1N(n3708), .Y(
        \i_MIPS/Register/n341 ) );
  OAI2BB2XL U11487 ( .B0(n3662), .B1(n3711), .A0N(
        \i_MIPS/Register/register[23][1] ), .A1N(n3712), .Y(
        \i_MIPS/Register/n373 ) );
  OAI2BB2XL U11488 ( .B0(n3015), .B1(n3714), .A0N(
        \i_MIPS/Register/register[22][1] ), .A1N(n3714), .Y(
        \i_MIPS/Register/n405 ) );
  OAI2BB2XL U11489 ( .B0(n3015), .B1(n3717), .A0N(
        \i_MIPS/Register/register[21][1] ), .A1N(n3718), .Y(
        \i_MIPS/Register/n437 ) );
  OAI2BB2XL U11490 ( .B0(n3015), .B1(n3720), .A0N(
        \i_MIPS/Register/register[20][1] ), .A1N(n3720), .Y(
        \i_MIPS/Register/n469 ) );
  OAI2BB2XL U11491 ( .B0(n3015), .B1(n3723), .A0N(
        \i_MIPS/Register/register[19][1] ), .A1N(n3724), .Y(
        \i_MIPS/Register/n501 ) );
  OAI2BB2XL U11492 ( .B0(n3015), .B1(n3726), .A0N(
        \i_MIPS/Register/register[18][1] ), .A1N(n3726), .Y(
        \i_MIPS/Register/n533 ) );
  OAI2BB2XL U11493 ( .B0(n3015), .B1(n3729), .A0N(
        \i_MIPS/Register/register[17][1] ), .A1N(n3730), .Y(
        \i_MIPS/Register/n565 ) );
  OAI2BB2XL U11494 ( .B0(n3662), .B1(n3732), .A0N(
        \i_MIPS/Register/register[16][1] ), .A1N(n3732), .Y(
        \i_MIPS/Register/n597 ) );
  OAI2BB2XL U11495 ( .B0(n3015), .B1(n3735), .A0N(
        \i_MIPS/Register/register[15][1] ), .A1N(n3736), .Y(
        \i_MIPS/Register/n629 ) );
  OAI2BB2XL U11496 ( .B0(n3662), .B1(n3738), .A0N(
        \i_MIPS/Register/register[14][1] ), .A1N(n3738), .Y(
        \i_MIPS/Register/n661 ) );
  OAI2BB2XL U11497 ( .B0(n3662), .B1(n3690), .A0N(
        \i_MIPS/Register/register[30][1] ), .A1N(n3691), .Y(
        \i_MIPS/Register/n149 ) );
  OAI2BB2XL U11498 ( .B0(n3662), .B1(n3741), .A0N(
        \i_MIPS/Register/register[13][1] ), .A1N(n3742), .Y(
        \i_MIPS/Register/n693 ) );
  OAI2BB2XL U11499 ( .B0(n3662), .B1(n3744), .A0N(
        \i_MIPS/Register/register[12][1] ), .A1N(n3744), .Y(
        \i_MIPS/Register/n725 ) );
  OAI2BB2XL U11500 ( .B0(n3662), .B1(n3747), .A0N(
        \i_MIPS/Register/register[11][1] ), .A1N(n3748), .Y(
        \i_MIPS/Register/n757 ) );
  OAI2BB2XL U11501 ( .B0(n3662), .B1(n3750), .A0N(
        \i_MIPS/Register/register[10][1] ), .A1N(n3750), .Y(
        \i_MIPS/Register/n789 ) );
  OAI2BB2XL U11502 ( .B0(n3662), .B1(n3753), .A0N(
        \i_MIPS/Register/register[9][1] ), .A1N(n3754), .Y(
        \i_MIPS/Register/n821 ) );
  OAI2BB2XL U11503 ( .B0(n3662), .B1(n3756), .A0N(
        \i_MIPS/Register/register[8][1] ), .A1N(n3757), .Y(
        \i_MIPS/Register/n853 ) );
  OAI2BB2XL U11504 ( .B0(n3662), .B1(n3759), .A0N(
        \i_MIPS/Register/register[7][1] ), .A1N(n3760), .Y(
        \i_MIPS/Register/n885 ) );
  OAI2BB2XL U11505 ( .B0(n3662), .B1(n3762), .A0N(
        \i_MIPS/Register/register[6][1] ), .A1N(n3763), .Y(
        \i_MIPS/Register/n917 ) );
  OAI2BB2XL U11506 ( .B0(n3015), .B1(n3765), .A0N(
        \i_MIPS/Register/register[5][1] ), .A1N(n3765), .Y(
        \i_MIPS/Register/n949 ) );
  OAI2BB2XL U11507 ( .B0(n3015), .B1(n3768), .A0N(
        \i_MIPS/Register/register[4][1] ), .A1N(n3768), .Y(
        \i_MIPS/Register/n981 ) );
  OAI2BB2XL U11508 ( .B0(n3015), .B1(n3771), .A0N(
        \i_MIPS/Register/register[3][1] ), .A1N(n3771), .Y(
        \i_MIPS/Register/n1013 ) );
  OAI2BB2XL U11509 ( .B0(n3015), .B1(n3774), .A0N(
        \i_MIPS/Register/register[2][1] ), .A1N(n3775), .Y(
        \i_MIPS/Register/n1045 ) );
  OAI2BB2XL U11510 ( .B0(n3015), .B1(n3777), .A0N(
        \i_MIPS/Register/register[1][1] ), .A1N(n3777), .Y(
        \i_MIPS/Register/n1077 ) );
  OAI2BB2XL U11511 ( .B0(n3015), .B1(n3780), .A0N(
        \i_MIPS/Register/register[0][1] ), .A1N(n3781), .Y(
        \i_MIPS/Register/n1109 ) );
  OAI222XL U11512 ( .A0(n3584), .A1(n206), .B0(n3015), .B1(n3583), .C0(n3689), 
        .C1(\i_MIPS/n181 ), .Y(n8803) );
  NAND3BXL U11513 ( .AN(n4726), .B(n4725), .C(n5048), .Y(n6842) );
  INVX4 U11514 ( .A(n6985), .Y(n7021) );
  NAND2XL U11515 ( .A(n5185), .B(n5184), .Y(n6128) );
  AO22XL U11516 ( .A0(n5892), .A1(n3102), .B0(n3109), .B1(n5893), .Y(n5897) );
  OAI221XL U11517 ( .A0(n3106), .A1(n5893), .B0(n5892), .B1(n3098), .C0(n3097), 
        .Y(n5894) );
  OAI222XL U11518 ( .A0(n5598), .A1(n3218), .B0(n5597), .B1(n3216), .C0(n3646), 
        .C1(n3215), .Y(n3034) );
  OAI221X4 U11519 ( .A0(n8769), .A1(n7044), .B0(n8756), .B1(n7043), .C0(n6502), 
        .Y(n6503) );
  CLKBUFX2 U11520 ( .A(n8743), .Y(n3685) );
  OAI221X4 U11521 ( .A0(n8770), .A1(n7044), .B0(n8757), .B1(n7043), .C0(n4866), 
        .Y(n4867) );
  OAI2BB2XL U11522 ( .B0(n3030), .B1(n3780), .A0N(
        \i_MIPS/Register/register[0][5] ), .A1N(n3782), .Y(
        \i_MIPS/Register/n1113 ) );
  OAI2BB2XL U11523 ( .B0(n3030), .B1(n3777), .A0N(
        \i_MIPS/Register/register[1][5] ), .A1N(n3779), .Y(
        \i_MIPS/Register/n1081 ) );
  OAI2BB2XL U11524 ( .B0(n3030), .B1(n3774), .A0N(
        \i_MIPS/Register/register[2][5] ), .A1N(n3776), .Y(
        \i_MIPS/Register/n1049 ) );
  OAI2BB2XL U11525 ( .B0(n3030), .B1(n3771), .A0N(
        \i_MIPS/Register/register[3][5] ), .A1N(n3773), .Y(
        \i_MIPS/Register/n1017 ) );
  OAI2BB2XL U11526 ( .B0(n3030), .B1(n3768), .A0N(
        \i_MIPS/Register/register[4][5] ), .A1N(n3770), .Y(
        \i_MIPS/Register/n985 ) );
  OAI2BB2XL U11527 ( .B0(n3030), .B1(n3765), .A0N(
        \i_MIPS/Register/register[5][5] ), .A1N(n3767), .Y(
        \i_MIPS/Register/n953 ) );
  OAI2BB2XL U11528 ( .B0(n3030), .B1(n3762), .A0N(
        \i_MIPS/Register/register[6][5] ), .A1N(n3764), .Y(
        \i_MIPS/Register/n921 ) );
  OAI222XL U11529 ( .A0(n3584), .A1(n207), .B0(n3030), .B1(n3583), .C0(n3688), 
        .C1(\i_MIPS/n185 ), .Y(n8799) );
  CLKBUFX2 U11530 ( .A(n8720), .Y(n3642) );
  OAI221X4 U11531 ( .A0(n8761), .A1(n7044), .B0(n8748), .B1(n7043), .C0(n5859), 
        .Y(n5860) );
  INVX12 U11532 ( .A(n1847), .Y(DCACHE_addr[29]) );
  OAI222XL U11533 ( .A0(n5379), .A1(n3218), .B0(n5378), .B1(n3216), .C0(n8735), 
        .C1(n3215), .Y(n3036) );
  AOI2BB2X2 U11534 ( .B0(\D_cache/N121 ), .B1(n2153), .A0N(n23), .A1N(n8871), 
        .Y(\D_cache/n175 ) );
  CLKBUFX2 U11535 ( .A(n8736), .Y(n3669) );
  NAND2X1 U11536 ( .A(n5398), .B(n5390), .Y(n5391) );
  CLKBUFX2 U11537 ( .A(n8740), .Y(n3677) );
  CLKBUFX2 U11538 ( .A(n8742), .Y(n3682) );
  AOI2BB2X2 U11539 ( .B0(\D_cache/N131 ), .B1(n2153), .A0N(n23), .A1N(n8881), 
        .Y(\D_cache/n186 ) );
  AOI2BB2X2 U11540 ( .B0(\D_cache/N132 ), .B1(n2153), .A0N(n24), .A1N(n8882), 
        .Y(\D_cache/n187 ) );
  OAI2BB2XL U11541 ( .B0(n3673), .B1(n3763), .A0N(
        \i_MIPS/Register/register[6][24] ), .A1N(n3764), .Y(
        \i_MIPS/Register/n940 ) );
  OAI2BB2XL U11542 ( .B0(n3674), .B1(n3766), .A0N(
        \i_MIPS/Register/register[5][24] ), .A1N(n3767), .Y(
        \i_MIPS/Register/n972 ) );
  OAI2BB2XL U11543 ( .B0(n3674), .B1(n3769), .A0N(
        \i_MIPS/Register/register[4][24] ), .A1N(n3770), .Y(
        \i_MIPS/Register/n1004 ) );
  OAI2BB2XL U11544 ( .B0(n3673), .B1(n3772), .A0N(
        \i_MIPS/Register/register[3][24] ), .A1N(n3773), .Y(
        \i_MIPS/Register/n1036 ) );
  OAI2BB2XL U11545 ( .B0(n3673), .B1(n3775), .A0N(
        \i_MIPS/Register/register[2][24] ), .A1N(n3776), .Y(
        \i_MIPS/Register/n1068 ) );
  OAI2BB2XL U11546 ( .B0(n3674), .B1(n3778), .A0N(
        \i_MIPS/Register/register[1][24] ), .A1N(n3779), .Y(
        \i_MIPS/Register/n1100 ) );
  OAI2BB2XL U11547 ( .B0(n3674), .B1(n3781), .A0N(
        \i_MIPS/Register/register[0][24] ), .A1N(n3782), .Y(
        \i_MIPS/Register/n1132 ) );
  OAI222XL U11548 ( .A0(n3584), .A1(n208), .B0(n3673), .B1(n3582), .C0(n3689), 
        .C1(\i_MIPS/n204 ), .Y(n8780) );
  CLKBUFX2 U11549 ( .A(n8745), .Y(n3687) );
  OAI2BB2XL U11550 ( .B0(n3671), .B1(n45), .A0N(
        \i_MIPS/Register/register[6][26] ), .A1N(n3764), .Y(
        \i_MIPS/Register/n942 ) );
  OAI2BB2XL U11551 ( .B0(n3671), .B1(n3765), .A0N(
        \i_MIPS/Register/register[5][26] ), .A1N(n3767), .Y(
        \i_MIPS/Register/n974 ) );
  OAI2BB2XL U11552 ( .B0(n3671), .B1(n47), .A0N(
        \i_MIPS/Register/register[4][26] ), .A1N(n3770), .Y(
        \i_MIPS/Register/n1006 ) );
  OAI2BB2XL U11553 ( .B0(n3672), .B1(n48), .A0N(
        \i_MIPS/Register/register[3][26] ), .A1N(n3773), .Y(
        \i_MIPS/Register/n1038 ) );
  OAI2BB2XL U11554 ( .B0(n3671), .B1(n49), .A0N(
        \i_MIPS/Register/register[2][26] ), .A1N(n3776), .Y(
        \i_MIPS/Register/n1070 ) );
  OAI2BB2XL U11555 ( .B0(n3671), .B1(n3777), .A0N(
        \i_MIPS/Register/register[1][26] ), .A1N(n3779), .Y(
        \i_MIPS/Register/n1102 ) );
  OAI2BB2XL U11556 ( .B0(n3671), .B1(n51), .A0N(
        \i_MIPS/Register/register[0][26] ), .A1N(n3782), .Y(
        \i_MIPS/Register/n1134 ) );
  OAI222XL U11557 ( .A0(n3584), .A1(n71), .B0(n3672), .B1(n3582), .C0(n3688), 
        .C1(\i_MIPS/n206 ), .Y(n8778) );
  MX2XL U11558 ( .A(n1886), .B(n7783), .S0(n3626), .Y(\i_MIPS/n431 ) );
  CLKBUFX2 U11559 ( .A(n8719), .Y(n3640) );
  CLKBUFX2 U11560 ( .A(n8725), .Y(n3648) );
  INVXL U11561 ( .A(n8214), .Y(n8248) );
  AND4X4 U11562 ( .A(n3042), .B(n3043), .C(n3044), .D(n3045), .Y(
        \D_cache/n525 ) );
  MX2XL U11563 ( .A(DCACHE_addr[8]), .B(n8012), .S0(n3625), .Y(\i_MIPS/n459 )
         );
  MX2XL U11564 ( .A(n1891), .B(n8222), .S0(n3625), .Y(\i_MIPS/n413 ) );
  MX2XL U11565 ( .A(DCACHE_addr[15]), .B(n8255), .S0(n3626), .Y(\i_MIPS/n452 )
         );
  MX2XL U11566 ( .A(n1888), .B(n7807), .S0(n3625), .Y(\i_MIPS/n423 ) );
  CLKBUFX2 U11567 ( .A(n2795), .Y(n3680) );
  MX2XL U11568 ( .A(\i_MIPS/ID_EX[58] ), .B(n7809), .S0(n3626), .Y(
        \i_MIPS/n403 ) );
  MXI2XL U11569 ( .A(\i_MIPS/n351 ), .B(n8224), .S0(n3617), .Y(\i_MIPS/n542 )
         );
  CLKBUFX2 U11570 ( .A(n3019), .Y(n3650) );
  NAND3BX4 U11571 ( .AN(n4700), .B(n5473), .C(n5472), .Y(n4701) );
  NAND3BX4 U11572 ( .AN(n5985), .B(n4699), .C(n21), .Y(n5472) );
  OAI211X4 U11573 ( .A0(n4694), .A1(n4693), .B0(n5256), .C0(n5270), .Y(n6257)
         );
  CLKBUFX2 U11574 ( .A(n3020), .Y(n3664) );
  OAI2BB1XL U11575 ( .A0N(n8809), .A1N(\D_cache/n520 ), .B0(\D_cache/N30 ), 
        .Y(\D_cache/n518 ) );
  MX2XL U11576 ( .A(n10316), .B(n7786), .S0(n3627), .Y(\i_MIPS/n457 ) );
  OAI21XL U11577 ( .A0(\D_cache/n203 ), .A1(\D_cache/n384 ), .B0(
        \D_cache/n204 ), .Y(\D_cache/n451 ) );
  OAI21XL U11578 ( .A0(\D_cache/n201 ), .A1(\D_cache/n384 ), .B0(
        \D_cache/n204 ), .Y(\D_cache/n383 ) );
  OAI31XL U11579 ( .A0(\D_cache/n201 ), .A1(\D_cache/n202 ), .A2(
        \D_cache/n203 ), .B0(\D_cache/n204 ), .Y(\D_cache/n519 ) );
  OAI31XL U11580 ( .A0(\D_cache/n201 ), .A1(n8903), .A2(\D_cache/n203 ), .B0(
        \D_cache/n204 ), .Y(\D_cache/n315 ) );
  AOI222XL U11581 ( .A0(\D_cache/n520 ), .A1(\D_cache/n247 ), .B0(
        \D_cache/n204 ), .B1(DCACHE_ren), .C0(n8772), .C1(n8808), .Y(
        \D_cache/n314 ) );
  OAI2BB2XL U11582 ( .B0(n8729), .B1(n3762), .A0N(
        \i_MIPS/Register/register[6][12] ), .A1N(n3764), .Y(
        \i_MIPS/Register/n928 ) );
  OAI2BB2XL U11583 ( .B0(n8729), .B1(n3765), .A0N(
        \i_MIPS/Register/register[5][12] ), .A1N(n3767), .Y(
        \i_MIPS/Register/n960 ) );
  OAI2BB2XL U11584 ( .B0(n8729), .B1(n3768), .A0N(
        \i_MIPS/Register/register[4][12] ), .A1N(n3770), .Y(
        \i_MIPS/Register/n992 ) );
  OAI2BB2XL U11585 ( .B0(n8729), .B1(n3771), .A0N(
        \i_MIPS/Register/register[3][12] ), .A1N(n3773), .Y(
        \i_MIPS/Register/n1024 ) );
  OAI2BB2XL U11586 ( .B0(n8729), .B1(n3774), .A0N(
        \i_MIPS/Register/register[2][12] ), .A1N(n3776), .Y(
        \i_MIPS/Register/n1056 ) );
  OAI2BB2XL U11587 ( .B0(n8729), .B1(n3777), .A0N(
        \i_MIPS/Register/register[1][12] ), .A1N(n3779), .Y(
        \i_MIPS/Register/n1088 ) );
  OAI2BB2XL U11588 ( .B0(n8729), .B1(n3780), .A0N(
        \i_MIPS/Register/register[0][12] ), .A1N(n3782), .Y(
        \i_MIPS/Register/n1120 ) );
  OAI222XL U11589 ( .A0(n3584), .A1(n209), .B0(n8729), .B1(n3582), .C0(n3689), 
        .C1(\i_MIPS/n192 ), .Y(n8792) );
  MX2XL U11590 ( .A(n10315), .B(n8249), .S0(n3626), .Y(\i_MIPS/n456 ) );
  OAI31X4 U11591 ( .A0(n7873), .A1(n7872), .A2(n7871), .B0(n7870), .Y(n7952)
         );
  NAND2X1 U11592 ( .A(n7788), .B(\i_MIPS/n233 ), .Y(n7791) );
  AOI221X2 U11593 ( .A0(n7078), .A1(n7788), .B0(n7078), .B1(n7789), .C0(n7833), 
        .Y(n7079) );
  NAND2X1 U11594 ( .A(n6993), .B(n2892), .Y(n5061) );
  OAI221XL U11595 ( .A0(n6765), .A1(n3106), .B0(n6764), .B1(n3098), .C0(n3096), 
        .Y(n6767) );
  AO22XL U11596 ( .A0(n2839), .A1(n3104), .B0(n3111), .B1(n2892), .Y(n5126) );
  NAND2X1 U11597 ( .A(n6533), .B(n6532), .Y(n6601) );
  MX2XL U11598 ( .A(\i_MIPS/ID_EX[62] ), .B(n8161), .S0(n3624), .Y(
        \i_MIPS/n395 ) );
  MX2XL U11599 ( .A(\i_MIPS/ID_EX[66] ), .B(n8038), .S0(n3624), .Y(
        \i_MIPS/n387 ) );
  OA22X4 U11600 ( .A0(n3280), .A1(n1007), .B0(n3264), .B1(n119), .Y(n4427) );
  OA22X4 U11601 ( .A0(n3285), .A1(n1008), .B0(n3237), .B1(n120), .Y(n4455) );
  OA22X4 U11602 ( .A0(n3547), .A1(n1009), .B0(n3506), .B1(n121), .Y(n4452) );
  OA22X4 U11603 ( .A0(n3285), .A1(n1010), .B0(n3237), .B1(n122), .Y(n4459) );
  CLKINVX3 U11604 ( .A(n4667), .Y(n4687) );
  NAND2X2 U11605 ( .A(n4687), .B(\i_MIPS/n363 ), .Y(n8467) );
  OAI211X2 U11606 ( .A0(n4596), .A1(n5192), .B0(n8466), .C0(n7), .Y(n6260) );
  OAI31X2 U11607 ( .A0(n2758), .A1(n8479), .A2(n4822), .B0(n4600), .Y(n5976)
         );
  OAI211X2 U11608 ( .A0(n4604), .A1(n4603), .B0(n4602), .C0(n4601), .Y(n5470)
         );
  OAI211X2 U11609 ( .A0(n4605), .A1(n8462), .B0(n8517), .C0(n8522), .Y(n4606)
         );
  NAND2X2 U11610 ( .A(n4606), .B(n8461), .Y(n6761) );
  CLKINVX3 U11611 ( .A(\i_MIPS/ALUin1[28] ), .Y(n5900) );
  CLKINVX3 U11612 ( .A(n4617), .Y(n4622) );
  NAND4BX2 U11613 ( .AN(n4621), .B(n4620), .C(\i_MIPS/ALU_Control/n20 ), .D(
        n4619), .Y(n4724) );
  CLKINVX3 U11614 ( .A(n4724), .Y(n4728) );
  NAND2X2 U11615 ( .A(\i_MIPS/ALUin1[15] ), .B(n4647), .Y(n5545) );
  NAND2X2 U11616 ( .A(\i_MIPS/ALUin1[6] ), .B(n4672), .Y(n4971) );
  NAND2X2 U11617 ( .A(\i_MIPS/ALUin1[3] ), .B(n4677), .Y(n6537) );
  NAND2X2 U11618 ( .A(\i_MIPS/ALUin1[1] ), .B(n5106), .Y(n6533) );
  NAND2X2 U11619 ( .A(\i_MIPS/ALUin1[2] ), .B(n2716), .Y(n6603) );
  AND3X4 U11620 ( .A(n4685), .B(n5185), .C(n5184), .Y(n4694) );
  NAND2X2 U11621 ( .A(\i_MIPS/ALUin1[8] ), .B(n4687), .Y(n6188) );
  OAI211X2 U11622 ( .A0(n4698), .A1(n4697), .B0(n5621), .C0(n4696), .Y(n6467)
         );
  NAND2X2 U11623 ( .A(n2834), .B(\i_MIPS/ID_EX[83] ), .Y(n7009) );
  OAI222X2 U11624 ( .A0(n4810), .A1(n3165), .B0(n4773), .B1(n2761), .C0(n8718), 
        .C1(n3163), .Y(n7661) );
  OAI222X2 U11625 ( .A0(n4810), .A1(n3219), .B0(n4809), .B1(n3216), .C0(n8718), 
        .C1(n3214), .Y(n8313) );
  NAND2BX2 U11626 ( .AN(n4823), .B(n6389), .Y(n6323) );
  CLKMX2X4 U11627 ( .A(n1087), .B(\D_cache/n187 ), .S0(n4021), .Y(n4866) );
  OAI221X2 U11628 ( .A0(\i_MIPS/n371 ), .A1(n3087), .B0(n5381), .B1(n3077), 
        .C0(n5042), .Y(n6619) );
  CLKINVX3 U11629 ( .A(n5396), .Y(n5121) );
  AO21X4 U11630 ( .A0(n2825), .A1(n6324), .B0(n5675), .Y(n6911) );
  AO21X4 U11631 ( .A0(n6911), .A1(n6913), .B0(n6917), .Y(n5735) );
  AO21X4 U11632 ( .A0(n5735), .A1(n5734), .B0(n5733), .Y(n5737) );
  NAND4BX2 U11633 ( .AN(n5760), .B(n7014), .C(n5759), .D(n5758), .Y(n7977) );
  OAI222X2 U11634 ( .A0(n5883), .A1(n3218), .B0(n5882), .B1(n3217), .C0(n8720), 
        .C1(n3215), .Y(n8283) );
  NOR3BX4 U11635 ( .AN(n5886), .B(n5885), .C(n5884), .Y(n6981) );
  NAND3BX2 U11636 ( .AN(n5911), .B(n5910), .C(n5909), .Y(n8266) );
  OAI222X2 U11637 ( .A0(n5956), .A1(n3218), .B0(n5955), .B1(n3217), .C0(n8721), 
        .C1(n3215), .Y(n8265) );
  AOI2BB1X2 U11638 ( .A0N(n5986), .A1N(n5985), .B0(n5984), .Y(n5987) );
  OAI222X2 U11639 ( .A0(n6045), .A1(n3218), .B0(n6044), .B1(n3217), .C0(n3), 
        .C1(n3215), .Y(n8037) );
  NAND3BX2 U11640 ( .AN(n6144), .B(n6143), .C(n6142), .Y(n8231) );
  CLKMX2X4 U11641 ( .A(n1088), .B(\D_cache/n186 ), .S0(n4022), .Y(n6502) );
  OAI222X2 U11642 ( .A0(n6823), .A1(n3166), .B0(n6801), .B1(n2761), .C0(n8723), 
        .C1(n3162), .Y(n8199) );
  OAI222X2 U11643 ( .A0(n6823), .A1(n3219), .B0(n6822), .B1(n3217), .C0(n8723), 
        .C1(n3214), .Y(n8166) );
  NOR4BX4 U11644 ( .AN(n6978), .B(n6977), .C(n6976), .D(n6975), .Y(n6979) );
  OAI222X2 U11645 ( .A0(n7072), .A1(n3164), .B0(n7047), .B1(n2761), .C0(n8719), 
        .C1(n3163), .Y(n8308) );
  OAI222X2 U11646 ( .A0(n7072), .A1(n3219), .B0(n7070), .B1(n3216), .C0(n8719), 
        .C1(n3214), .Y(n7633) );
  OAI221X2 U11647 ( .A0(n7787), .A1(n7081), .B0(n7080), .B1(n7832), .C0(n7079), 
        .Y(n7840) );
  OAI211X2 U11648 ( .A0(n1627), .A1(n7834), .B0(n7833), .C0(n3611), .Y(n8415)
         );
  NAND2X2 U11649 ( .A(n7865), .B(n7864), .Y(n7871) );
  AO22X4 U11650 ( .A0(n7950), .A1(n7949), .B0(n2861), .B1(n7951), .Y(n8017) );
  NAND2X2 U11651 ( .A(n8016), .B(ICACHE_addr[15]), .Y(n7995) );
  CLKINVX3 U11652 ( .A(n8023), .Y(n8019) );
  NAND2X2 U11653 ( .A(n8056), .B(ICACHE_addr[17]), .Y(n8041) );
  NAND2X2 U11654 ( .A(n8080), .B(ICACHE_addr[19]), .Y(n8057) );
  NAND2X2 U11655 ( .A(n8142), .B(ICACHE_addr[21]), .Y(n8121) );
  NAND3BX2 U11656 ( .AN(n8362), .B(n8361), .C(n8360), .Y(\i_MIPS/PC/n40 ) );
  CLKINVX3 U11657 ( .A(n8393), .Y(n8394) );
endmodule

