
module CHIP ( clk, rst_n, mem_read_D, mem_write_D, mem_addr_D, mem_wdata_D, 
        mem_rdata_D, mem_ready_D, mem_read_I, mem_write_I, mem_addr_I, 
        mem_wdata_I, mem_rdata_I, mem_ready_I, DCACHE_addr, DCACHE_wdata, 
        DCACHE_wen );
  output [31:4] mem_addr_D;
  output [127:0] mem_wdata_D;
  input [127:0] mem_rdata_D;
  output [31:4] mem_addr_I;
  output [127:0] mem_wdata_I;
  input [127:0] mem_rdata_I;
  output [29:0] DCACHE_addr;
  output [31:0] DCACHE_wdata;
  input clk, rst_n, mem_ready_D, mem_ready_I;
  output mem_read_D, mem_write_D, mem_read_I, mem_write_I, DCACHE_wen;
  wire   n12788, n12789, n12790, n12791, n12792, n12793, n12794, n12795,
         n12796, n12797, n12798, n12799, n12800, n12801, n12802, n12803,
         n12804, n12805, n12806, n12807, n12808, n12809, n12810, n12811,
         n12812, n12813, n12814, n12815, n12816, n12817, n12818, n12819,
         n12820, n12821, n12822, n12823, n12824, n12825, n12826, n12827,
         n12828, n12829, n12830, n12831, n12832, n12833, n12834, n12835,
         n12836, n12837, n12838, n12839, n12840, n12841, n12842, n12843,
         n12844, n12845, n12846, n12847, n12848, n12849, n12850, n12851,
         n12852, n12853, n12854, n12855, n12856, n12857, n12858, n12859,
         n12860, n12861, n12862, n12863, n12864, n12865, n12866, n12867,
         n12868, n12869, n12870, n12871, n12872, n12873, n12874, n12875,
         n12876, n12877, n12878, n12879, n12880, n12881, n12882, n12883,
         n12884, n12885, n12886, n12887, n12888, n12889, n12890, n12891,
         n12892, n12893, n12894, n12895, n12896, n12897, n12898, n12899,
         n12900, n12901, n12902, n12903, n12904, n12905, n12906, n12907,
         n12908, n12909, n12910, n12911, n12912, n12913, n12914, n12915,
         n12916, n12917, n12918, n12919, n12920, n12921, n12922, n12923,
         n12924, n12925, n12926, n12927, n12928, n12929, n12930, n12931,
         n12932, n12933, n12934, n12935, n12936, n12937, n12938, n12939,
         n12940, n12941, n12942, n12943, n12944, n12945, n12946, n12947,
         n12948, n12949, n12950, n12951, n12952, n12953, n12954, n12955,
         n12956, n12957, n12958, n12959, n12960, n12961, n12962, n12963,
         n12964, n12965, n12966, n12967, n12968, n12969, n12970, n12971,
         n12972, n12973, n12974, n12975, n12976, n12977, n12978, n12979,
         n12980, n12981, n12982, n12983, n12984, n12985, n12986, n12987,
         n12988, DCACHE_ren, \i_MIPS/n567 , \i_MIPS/n563 , \i_MIPS/n562 ,
         \i_MIPS/n561 , \i_MIPS/n560 , \i_MIPS/n559 , \i_MIPS/n558 ,
         \i_MIPS/n557 , \i_MIPS/n556 , \i_MIPS/n555 , \i_MIPS/n554 ,
         \i_MIPS/n553 , \i_MIPS/n552 , \i_MIPS/n551 , \i_MIPS/n550 ,
         \i_MIPS/n549 , \i_MIPS/n548 , \i_MIPS/n547 , \i_MIPS/n546 ,
         \i_MIPS/n545 , \i_MIPS/n544 , \i_MIPS/n543 , \i_MIPS/n542 ,
         \i_MIPS/n541 , \i_MIPS/n540 , \i_MIPS/n539 , \i_MIPS/n538 ,
         \i_MIPS/n537 , \i_MIPS/n536 , \i_MIPS/n535 , \i_MIPS/n534 ,
         \i_MIPS/n533 , \i_MIPS/n532 , \i_MIPS/n531 , \i_MIPS/n530 ,
         \i_MIPS/n529 , \i_MIPS/n528 , \i_MIPS/n527 , \i_MIPS/n526 ,
         \i_MIPS/n525 , \i_MIPS/n524 , \i_MIPS/n523 , \i_MIPS/n522 ,
         \i_MIPS/n521 , \i_MIPS/n520 , \i_MIPS/n519 , \i_MIPS/n518 ,
         \i_MIPS/n517 , \i_MIPS/n516 , \i_MIPS/n515 , \i_MIPS/n514 ,
         \i_MIPS/n513 , \i_MIPS/n512 , \i_MIPS/n511 , \i_MIPS/n510 ,
         \i_MIPS/n509 , \i_MIPS/n508 , \i_MIPS/n507 , \i_MIPS/n506 ,
         \i_MIPS/n505 , \i_MIPS/n504 , \i_MIPS/n503 , \i_MIPS/n502 ,
         \i_MIPS/n501 , \i_MIPS/n500 , \i_MIPS/n499 , \i_MIPS/n498 ,
         \i_MIPS/n497 , \i_MIPS/n496 , \i_MIPS/n495 , \i_MIPS/n494 ,
         \i_MIPS/n493 , \i_MIPS/n492 , \i_MIPS/n491 , \i_MIPS/n490 ,
         \i_MIPS/n489 , \i_MIPS/n488 , \i_MIPS/n487 , \i_MIPS/n486 ,
         \i_MIPS/n485 , \i_MIPS/n484 , \i_MIPS/n483 , \i_MIPS/n482 ,
         \i_MIPS/n481 , \i_MIPS/n480 , \i_MIPS/n479 , \i_MIPS/n478 ,
         \i_MIPS/n477 , \i_MIPS/n476 , \i_MIPS/n475 , \i_MIPS/n474 ,
         \i_MIPS/n473 , \i_MIPS/n472 , \i_MIPS/n471 , \i_MIPS/n470 ,
         \i_MIPS/n469 , \i_MIPS/n468 , \i_MIPS/n467 , \i_MIPS/n466 ,
         \i_MIPS/n465 , \i_MIPS/n464 , \i_MIPS/n463 , \i_MIPS/n462 ,
         \i_MIPS/n461 , \i_MIPS/n460 , \i_MIPS/n459 , \i_MIPS/n458 ,
         \i_MIPS/n457 , \i_MIPS/n456 , \i_MIPS/n455 , \i_MIPS/n454 ,
         \i_MIPS/n453 , \i_MIPS/n452 , \i_MIPS/n451 , \i_MIPS/n450 ,
         \i_MIPS/n449 , \i_MIPS/n448 , \i_MIPS/n447 , \i_MIPS/n446 ,
         \i_MIPS/n445 , \i_MIPS/n444 , \i_MIPS/n443 , \i_MIPS/n442 ,
         \i_MIPS/n441 , \i_MIPS/n440 , \i_MIPS/n439 , \i_MIPS/n438 ,
         \i_MIPS/n437 , \i_MIPS/n436 , \i_MIPS/n435 , \i_MIPS/n434 ,
         \i_MIPS/n433 , \i_MIPS/n432 , \i_MIPS/n431 , \i_MIPS/n430 ,
         \i_MIPS/n429 , \i_MIPS/n428 , \i_MIPS/n427 , \i_MIPS/n426 ,
         \i_MIPS/n425 , \i_MIPS/n424 , \i_MIPS/n423 , \i_MIPS/n422 ,
         \i_MIPS/n421 , \i_MIPS/n420 , \i_MIPS/n419 , \i_MIPS/n418 ,
         \i_MIPS/n417 , \i_MIPS/n416 , \i_MIPS/n415 , \i_MIPS/n414 ,
         \i_MIPS/n413 , \i_MIPS/n412 , \i_MIPS/n411 , \i_MIPS/n410 ,
         \i_MIPS/n409 , \i_MIPS/n408 , \i_MIPS/n407 , \i_MIPS/n406 ,
         \i_MIPS/n405 , \i_MIPS/n404 , \i_MIPS/n403 , \i_MIPS/n402 ,
         \i_MIPS/n401 , \i_MIPS/n400 , \i_MIPS/n399 , \i_MIPS/n398 ,
         \i_MIPS/n397 , \i_MIPS/n396 , \i_MIPS/n395 , \i_MIPS/n394 ,
         \i_MIPS/n393 , \i_MIPS/n392 , \i_MIPS/n391 , \i_MIPS/n390 ,
         \i_MIPS/n389 , \i_MIPS/n388 , \i_MIPS/n387 , \i_MIPS/n386 ,
         \i_MIPS/n385 , \i_MIPS/n384 , \i_MIPS/n383 , \i_MIPS/n382 ,
         \i_MIPS/n381 , \i_MIPS/n380 , \i_MIPS/n379 , \i_MIPS/n378 ,
         \i_MIPS/n377 , \i_MIPS/n376 , \i_MIPS/n375 , \i_MIPS/n374 ,
         \i_MIPS/n373 , \i_MIPS/n372 , \i_MIPS/n371 , \i_MIPS/n370 ,
         \i_MIPS/n369 , \i_MIPS/n368 , \i_MIPS/n367 , \i_MIPS/n366 ,
         \i_MIPS/n365 , \i_MIPS/n364 , \i_MIPS/n363 , \i_MIPS/n362 ,
         \i_MIPS/n361 , \i_MIPS/n360 , \i_MIPS/n359 , \i_MIPS/n358 ,
         \i_MIPS/n357 , \i_MIPS/n356 , \i_MIPS/n355 , \i_MIPS/n354 ,
         \i_MIPS/n353 , \i_MIPS/n352 , \i_MIPS/n351 , \i_MIPS/n350 ,
         \i_MIPS/n349 , \i_MIPS/n348 , \i_MIPS/n347 , \i_MIPS/n346 ,
         \i_MIPS/n345 , \i_MIPS/n344 , \i_MIPS/n343 , \i_MIPS/n341 ,
         \i_MIPS/n340 , \i_MIPS/n339 , \i_MIPS/n338 , \i_MIPS/n337 ,
         \i_MIPS/n336 , \i_MIPS/n335 , \i_MIPS/n334 , \i_MIPS/n333 ,
         \i_MIPS/n332 , \i_MIPS/n331 , \i_MIPS/n330 , \i_MIPS/n329 ,
         \i_MIPS/n328 , \i_MIPS/n327 , \i_MIPS/n326 , \i_MIPS/n325 ,
         \i_MIPS/n324 , \i_MIPS/n323 , \i_MIPS/n322 , \i_MIPS/n321 ,
         \i_MIPS/n320 , \i_MIPS/n319 , \i_MIPS/n318 , \i_MIPS/n317 ,
         \i_MIPS/n316 , \i_MIPS/n315 , \i_MIPS/n314 , \i_MIPS/n313 ,
         \i_MIPS/n312 , \i_MIPS/n311 , \i_MIPS/n310 , \i_MIPS/n309 ,
         \i_MIPS/n308 , \i_MIPS/n307 , \i_MIPS/n306 , \i_MIPS/n305 ,
         \i_MIPS/n304 , \i_MIPS/n303 , \i_MIPS/n302 , \i_MIPS/n301 ,
         \i_MIPS/n300 , \i_MIPS/n299 , \i_MIPS/n298 , \i_MIPS/n297 ,
         \i_MIPS/n296 , \i_MIPS/n295 , \i_MIPS/n294 , \i_MIPS/n293 ,
         \i_MIPS/n292 , \i_MIPS/n291 , \i_MIPS/n290 , \i_MIPS/n289 ,
         \i_MIPS/n288 , \i_MIPS/n287 , \i_MIPS/n286 , \i_MIPS/n285 ,
         \i_MIPS/n284 , \i_MIPS/n283 , \i_MIPS/n282 , \i_MIPS/n281 ,
         \i_MIPS/n280 , \i_MIPS/n279 , \i_MIPS/n278 , \i_MIPS/n277 ,
         \i_MIPS/n276 , \i_MIPS/n275 , \i_MIPS/n274 , \i_MIPS/n273 ,
         \i_MIPS/n272 , \i_MIPS/n271 , \i_MIPS/n270 , \i_MIPS/n269 ,
         \i_MIPS/n268 , \i_MIPS/n267 , \i_MIPS/n266 , \i_MIPS/n265 ,
         \i_MIPS/n264 , \i_MIPS/n263 , \i_MIPS/n262 , \i_MIPS/n261 ,
         \i_MIPS/n260 , \i_MIPS/n259 , \i_MIPS/n258 , \i_MIPS/n257 ,
         \i_MIPS/n256 , \i_MIPS/n255 , \i_MIPS/n254 , \i_MIPS/n253 ,
         \i_MIPS/n252 , \i_MIPS/n251 , \i_MIPS/n250 , \i_MIPS/n249 ,
         \i_MIPS/n248 , \i_MIPS/n247 , \i_MIPS/n246 , \i_MIPS/n245 ,
         \i_MIPS/n244 , \i_MIPS/n243 , \i_MIPS/n242 , \i_MIPS/n241 ,
         \i_MIPS/n240 , \i_MIPS/n239 , \i_MIPS/n238 , \i_MIPS/n237 ,
         \i_MIPS/n236 , \i_MIPS/n235 , \i_MIPS/n234 , \i_MIPS/n233 ,
         \i_MIPS/n232 , \i_MIPS/n231 , \i_MIPS/n230 , \i_MIPS/n229 ,
         \i_MIPS/n228 , \i_MIPS/n227 , \i_MIPS/n226 , \i_MIPS/n225 ,
         \i_MIPS/n224 , \i_MIPS/n223 , \i_MIPS/n222 , \i_MIPS/n221 ,
         \i_MIPS/n220 , \i_MIPS/n219 , \i_MIPS/n218 , \i_MIPS/n217 ,
         \i_MIPS/n216 , \i_MIPS/n215 , \i_MIPS/n214 , \i_MIPS/n213 ,
         \i_MIPS/n212 , \i_MIPS/n211 , \i_MIPS/n210 , \i_MIPS/n209 ,
         \i_MIPS/n208 , \i_MIPS/n207 , \i_MIPS/n206 , \i_MIPS/n205 ,
         \i_MIPS/n204 , \i_MIPS/n203 , \i_MIPS/n202 , \i_MIPS/n201 ,
         \i_MIPS/n200 , \i_MIPS/n199 , \i_MIPS/n198 , \i_MIPS/n197 ,
         \i_MIPS/n196 , \i_MIPS/n195 , \i_MIPS/n194 , \i_MIPS/n193 ,
         \i_MIPS/n192 , \i_MIPS/n191 , \i_MIPS/n190 , \i_MIPS/n189 ,
         \i_MIPS/n188 , \i_MIPS/n187 , \i_MIPS/n186 , \i_MIPS/n185 ,
         \i_MIPS/n184 , \i_MIPS/n183 , \i_MIPS/n182 , \i_MIPS/n181 ,
         \i_MIPS/n180 , \i_MIPS/n179 , \i_MIPS/n178 , \i_MIPS/n177 ,
         \i_MIPS/n176 , \i_MIPS/n175 , \i_MIPS/n174 , \i_MIPS/n173 ,
         \i_MIPS/n172 , \i_MIPS/n171 , \i_MIPS/n170 , \i_MIPS/n169 ,
         \i_MIPS/n168 , \i_MIPS/n167 , \i_MIPS/n166 , \i_MIPS/n165 ,
         \i_MIPS/n164 , \i_MIPS/n163 , \i_MIPS/n162 , \i_MIPS/n161 ,
         \i_MIPS/n160 , \i_MIPS/N123 , \i_MIPS/N122 , \i_MIPS/N121 ,
         \i_MIPS/N120 , \i_MIPS/N119 , \i_MIPS/N118 , \i_MIPS/N117 ,
         \i_MIPS/N116 , \i_MIPS/N115 , \i_MIPS/N114 , \i_MIPS/N113 ,
         \i_MIPS/N112 , \i_MIPS/N111 , \i_MIPS/N110 , \i_MIPS/N109 ,
         \i_MIPS/N108 , \i_MIPS/N107 , \i_MIPS/N106 , \i_MIPS/N105 ,
         \i_MIPS/N104 , \i_MIPS/N103 , \i_MIPS/N102 , \i_MIPS/N101 ,
         \i_MIPS/N100 , \i_MIPS/N99 , \i_MIPS/N98 , \i_MIPS/N97 , \i_MIPS/N96 ,
         \i_MIPS/N95 , \i_MIPS/N94 , \i_MIPS/N93 , \i_MIPS/N92 , \i_MIPS/N91 ,
         \i_MIPS/N90 , \i_MIPS/N89 , \i_MIPS/N88 , \i_MIPS/N87 , \i_MIPS/N86 ,
         \i_MIPS/N85 , \i_MIPS/N84 , \i_MIPS/N83 , \i_MIPS/N82 , \i_MIPS/N81 ,
         \i_MIPS/N80 , \i_MIPS/N79 , \i_MIPS/N78 , \i_MIPS/N77 , \i_MIPS/N76 ,
         \i_MIPS/N75 , \i_MIPS/N74 , \i_MIPS/N73 , \i_MIPS/N72 , \i_MIPS/N71 ,
         \i_MIPS/N70 , \i_MIPS/N69 , \i_MIPS/N68 , \i_MIPS/N67 , \i_MIPS/N66 ,
         \i_MIPS/N65 , \i_MIPS/N64 , \i_MIPS/N63 , \i_MIPS/N62 , \i_MIPS/N61 ,
         \i_MIPS/N60 , \i_MIPS/N59 , \i_MIPS/N58 , \i_MIPS/N57 , \i_MIPS/N56 ,
         \i_MIPS/N55 , \i_MIPS/N54 , \i_MIPS/N53 , \i_MIPS/N52 , \i_MIPS/N51 ,
         \i_MIPS/N50 , \i_MIPS/N49 , \i_MIPS/N48 , \i_MIPS/N47 , \i_MIPS/N46 ,
         \i_MIPS/N45 , \i_MIPS/N44 , \i_MIPS/N43 , \i_MIPS/N42 , \i_MIPS/N41 ,
         \i_MIPS/N40 , \i_MIPS/N39 , \i_MIPS/N38 , \i_MIPS/N37 , \i_MIPS/N36 ,
         \i_MIPS/N35 , \i_MIPS/N34 , \i_MIPS/N33 , \i_MIPS/N32 , \i_MIPS/N31 ,
         \i_MIPS/N30 , \i_MIPS/N29 , \i_MIPS/N28 , \i_MIPS/N27 , \i_MIPS/N26 ,
         \i_MIPS/ALUin1[30] , \i_MIPS/ALUin1[29] , \i_MIPS/ALUin1[28] ,
         \i_MIPS/ALUin1[27] , \i_MIPS/ALUin1[26] , \i_MIPS/ALUin1[25] ,
         \i_MIPS/ALUin1[24] , \i_MIPS/ALUin1[23] , \i_MIPS/ALUin1[22] ,
         \i_MIPS/ALUin1[21] , \i_MIPS/ALUin1[20] , \i_MIPS/ALUin1[19] ,
         \i_MIPS/ALUin1[18] , \i_MIPS/ALUin1[17] , \i_MIPS/ALUin1[16] ,
         \i_MIPS/ALUin1[15] , \i_MIPS/ALUin1[14] , \i_MIPS/ALUin1[13] ,
         \i_MIPS/ALUin1[12] , \i_MIPS/ALUin1[11] , \i_MIPS/ALUin1[10] ,
         \i_MIPS/ALUin1[9] , \i_MIPS/ALUin1[8] , \i_MIPS/ALUin1[7] ,
         \i_MIPS/ALUin1[6] , \i_MIPS/ALUin1[5] , \i_MIPS/ALUin1[4] ,
         \i_MIPS/ALUin1[3] , \i_MIPS/ALUin1[2] , \i_MIPS/ALUin1[1] ,
         \i_MIPS/ALUin1[0] , \i_MIPS/ALUOp[1] , \i_MIPS/EX_MEM_0 ,
         \i_MIPS/EX_MEM_1 , \i_MIPS/EX_MEM[5] , \i_MIPS/EX_MEM[6] ,
         \i_MIPS/EX_MEM_74 , \i_MIPS/Sign_Extend_ID[31] ,
         \i_MIPS/Sign_Extend_ID[8] , \i_MIPS/Sign_Extend_ID[6] ,
         \i_MIPS/Sign_Extend_ID[5] , \i_MIPS/Sign_Extend_ID[4] ,
         \i_MIPS/Sign_Extend_ID[3] , \i_MIPS/Sign_Extend_ID[2] ,
         \i_MIPS/Sign_Extend_ID[1] , \i_MIPS/Sign_Extend_ID[0] ,
         \i_MIPS/ID_EX_0 , \i_MIPS/ID_EX_3 , \i_MIPS/ID_EX_5 ,
         \i_MIPS/ID_EX[42] , \i_MIPS/ID_EX[43] , \i_MIPS/ID_EX[49] ,
         \i_MIPS/ID_EX[50] , \i_MIPS/ID_EX[64] , \i_MIPS/ID_EX[66] ,
         \i_MIPS/ID_EX[67] , \i_MIPS/ID_EX[68] , \i_MIPS/ID_EX[69] ,
         \i_MIPS/ID_EX[70] , \i_MIPS/ID_EX[73] , \i_MIPS/ID_EX[75] ,
         \i_MIPS/ID_EX[77] , \i_MIPS/ID_EX[78] , \i_MIPS/ID_EX[79] ,
         \i_MIPS/ID_EX[80] , \i_MIPS/ID_EX[81] , \i_MIPS/ID_EX[82] ,
         \i_MIPS/ID_EX[83] , \i_MIPS/ID_EX[84] , \i_MIPS/ID_EX[85] ,
         \i_MIPS/ID_EX[86] , \i_MIPS/ID_EX[88] , \i_MIPS/ID_EX[89] ,
         \i_MIPS/ID_EX[90] , \i_MIPS/ID_EX[91] , \i_MIPS/ID_EX[92] ,
         \i_MIPS/ID_EX[93] , \i_MIPS/ID_EX[94] , \i_MIPS/ID_EX[95] ,
         \i_MIPS/ID_EX[96] , \i_MIPS/ID_EX[97] , \i_MIPS/ID_EX[98] ,
         \i_MIPS/ID_EX[99] , \i_MIPS/ID_EX[100] , \i_MIPS/ID_EX[101] ,
         \i_MIPS/ID_EX[102] , \i_MIPS/ID_EX[103] , \i_MIPS/ID_EX[104] ,
         \i_MIPS/ID_EX[105] , \i_MIPS/ID_EX[106] , \i_MIPS/ID_EX[107] ,
         \i_MIPS/ID_EX[112] , \i_MIPS/ID_EX[114] , \i_MIPS/ID_EX[115] ,
         \i_MIPS/control_out[7] , \i_MIPS/control_out[0] , \i_MIPS/Reg_W[0] ,
         \i_MIPS/Reg_W[1] , \i_MIPS/Reg_W[2] , \i_MIPS/Reg_W[3] ,
         \i_MIPS/Reg_W[4] , \i_MIPS/IR_ID[16] , \i_MIPS/IR_ID[17] ,
         \i_MIPS/IR_ID[18] , \i_MIPS/IR_ID[19] , \i_MIPS/IR_ID[20] ,
         \i_MIPS/IR_ID[21] , \i_MIPS/IR_ID[22] , \i_MIPS/IR_ID[23] ,
         \i_MIPS/IR_ID[24] , \i_MIPS/IR_ID[25] , \i_MIPS/IR_ID[26] ,
         \i_MIPS/IR_ID[27] , \i_MIPS/IR_ID[28] , \i_MIPS/IR_ID[29] ,
         \i_MIPS/IR_ID[30] , \i_MIPS/IR_ID[31] , \i_MIPS/PC_o[1] ,
         \i_MIPS/IF_ID_28 , \i_MIPS/IF_ID_29 , \i_MIPS/IF_ID_30 ,
         \i_MIPS/IF_ID_31 , \i_MIPS/IF_ID[64] , \i_MIPS/IF_ID[65] ,
         \i_MIPS/IF_ID[66] , \i_MIPS/IF_ID[67] , \i_MIPS/IF_ID[68] ,
         \i_MIPS/IF_ID[69] , \i_MIPS/IF_ID[70] , \i_MIPS/IF_ID[71] ,
         \i_MIPS/IF_ID[72] , \i_MIPS/IF_ID[73] , \i_MIPS/IF_ID[74] ,
         \i_MIPS/IF_ID[75] , \i_MIPS/IF_ID[76] , \i_MIPS/IF_ID[77] ,
         \i_MIPS/IF_ID[78] , \i_MIPS/IF_ID[79] , \i_MIPS/IF_ID[80] ,
         \i_MIPS/IF_ID[81] , \i_MIPS/IF_ID[82] , \i_MIPS/IF_ID[83] ,
         \i_MIPS/IF_ID[84] , \i_MIPS/IF_ID[85] , \i_MIPS/IF_ID[86] ,
         \i_MIPS/IF_ID[87] , \i_MIPS/IF_ID[88] , \i_MIPS/IF_ID[89] ,
         \i_MIPS/IF_ID[90] , \i_MIPS/IF_ID[91] , \i_MIPS/IF_ID[92] ,
         \i_MIPS/IF_ID[93] , \i_MIPS/IF_ID[94] , \i_MIPS/IF_ID[95] ,
         \i_MIPS/IF_ID[96] , \i_MIPS/IF_ID[97] , \i_MIPS/BranchAddr[0] ,
         \D_cache/n1796 , \D_cache/n1795 , \D_cache/n1794 , \D_cache/n1793 ,
         \D_cache/n1792 , \D_cache/n1791 , \D_cache/n1790 , \D_cache/n1789 ,
         \D_cache/n1788 , \D_cache/n1787 , \D_cache/n1786 , \D_cache/n1785 ,
         \D_cache/n1784 , \D_cache/n1783 , \D_cache/n1782 , \D_cache/n1781 ,
         \D_cache/n1780 , \D_cache/n1779 , \D_cache/n1778 , \D_cache/n1777 ,
         \D_cache/n1776 , \D_cache/n1775 , \D_cache/n1774 , \D_cache/n1773 ,
         \D_cache/n1772 , \D_cache/n1771 , \D_cache/n1770 , \D_cache/n1769 ,
         \D_cache/n1768 , \D_cache/n1767 , \D_cache/n1766 , \D_cache/n1765 ,
         \D_cache/n1764 , \D_cache/n1763 , \D_cache/n1762 , \D_cache/n1761 ,
         \D_cache/n1760 , \D_cache/n1759 , \D_cache/n1758 , \D_cache/n1757 ,
         \D_cache/n1756 , \D_cache/n1755 , \D_cache/n1754 , \D_cache/n1753 ,
         \D_cache/n1752 , \D_cache/n1751 , \D_cache/n1750 , \D_cache/n1749 ,
         \D_cache/n1748 , \D_cache/n1747 , \D_cache/n1746 , \D_cache/n1745 ,
         \D_cache/n1744 , \D_cache/n1743 , \D_cache/n1742 , \D_cache/n1741 ,
         \D_cache/n1740 , \D_cache/n1739 , \D_cache/n1738 , \D_cache/n1737 ,
         \D_cache/n1736 , \D_cache/n1735 , \D_cache/n1734 , \D_cache/n1733 ,
         \D_cache/n1732 , \D_cache/n1731 , \D_cache/n1730 , \D_cache/n1729 ,
         \D_cache/n1728 , \D_cache/n1727 , \D_cache/n1726 , \D_cache/n1725 ,
         \D_cache/n1724 , \D_cache/n1723 , \D_cache/n1722 , \D_cache/n1721 ,
         \D_cache/n1720 , \D_cache/n1719 , \D_cache/n1718 , \D_cache/n1717 ,
         \D_cache/n1716 , \D_cache/n1715 , \D_cache/n1714 , \D_cache/n1713 ,
         \D_cache/n1712 , \D_cache/n1711 , \D_cache/n1710 , \D_cache/n1709 ,
         \D_cache/n1708 , \D_cache/n1707 , \D_cache/n1706 , \D_cache/n1705 ,
         \D_cache/n1704 , \D_cache/n1703 , \D_cache/n1702 , \D_cache/n1701 ,
         \D_cache/n1700 , \D_cache/n1699 , \D_cache/n1698 , \D_cache/n1697 ,
         \D_cache/n1696 , \D_cache/n1695 , \D_cache/n1694 , \D_cache/n1693 ,
         \D_cache/n1692 , \D_cache/n1691 , \D_cache/n1690 , \D_cache/n1689 ,
         \D_cache/n1688 , \D_cache/n1687 , \D_cache/n1686 , \D_cache/n1685 ,
         \D_cache/n1684 , \D_cache/n1683 , \D_cache/n1682 , \D_cache/n1681 ,
         \D_cache/n1680 , \D_cache/n1679 , \D_cache/n1678 , \D_cache/n1677 ,
         \D_cache/n1676 , \D_cache/n1675 , \D_cache/n1674 , \D_cache/n1673 ,
         \D_cache/n1672 , \D_cache/n1671 , \D_cache/n1670 , \D_cache/n1669 ,
         \D_cache/n1668 , \D_cache/n1667 , \D_cache/n1666 , \D_cache/n1665 ,
         \D_cache/n1664 , \D_cache/n1663 , \D_cache/n1662 , \D_cache/n1661 ,
         \D_cache/n1660 , \D_cache/n1659 , \D_cache/n1658 , \D_cache/n1657 ,
         \D_cache/n1656 , \D_cache/n1655 , \D_cache/n1654 , \D_cache/n1653 ,
         \D_cache/n1652 , \D_cache/n1651 , \D_cache/n1650 , \D_cache/n1649 ,
         \D_cache/n1648 , \D_cache/n1647 , \D_cache/n1646 , \D_cache/n1645 ,
         \D_cache/n1644 , \D_cache/n1643 , \D_cache/n1642 , \D_cache/n1641 ,
         \D_cache/n1640 , \D_cache/n1639 , \D_cache/n1638 , \D_cache/n1637 ,
         \D_cache/n1636 , \D_cache/n1635 , \D_cache/n1634 , \D_cache/n1633 ,
         \D_cache/n1632 , \D_cache/n1631 , \D_cache/n1630 , \D_cache/n1629 ,
         \D_cache/n1628 , \D_cache/n1627 , \D_cache/n1626 , \D_cache/n1625 ,
         \D_cache/n1624 , \D_cache/n1623 , \D_cache/n1622 , \D_cache/n1621 ,
         \D_cache/n1620 , \D_cache/n1619 , \D_cache/n1618 , \D_cache/n1617 ,
         \D_cache/n1616 , \D_cache/n1615 , \D_cache/n1614 , \D_cache/n1613 ,
         \D_cache/n1612 , \D_cache/n1611 , \D_cache/n1610 , \D_cache/n1609 ,
         \D_cache/n1608 , \D_cache/n1607 , \D_cache/n1606 , \D_cache/n1605 ,
         \D_cache/n1604 , \D_cache/n1603 , \D_cache/n1602 , \D_cache/n1601 ,
         \D_cache/n1600 , \D_cache/n1599 , \D_cache/n1598 , \D_cache/n1597 ,
         \D_cache/n1596 , \D_cache/n1595 , \D_cache/n1594 , \D_cache/n1593 ,
         \D_cache/n1592 , \D_cache/n1591 , \D_cache/n1590 , \D_cache/n1589 ,
         \D_cache/n1588 , \D_cache/n1587 , \D_cache/n1586 , \D_cache/n1585 ,
         \D_cache/n1584 , \D_cache/n1583 , \D_cache/n1582 , \D_cache/n1581 ,
         \D_cache/n1580 , \D_cache/n1579 , \D_cache/n1578 , \D_cache/n1577 ,
         \D_cache/n1576 , \D_cache/n1575 , \D_cache/n1574 , \D_cache/n1573 ,
         \D_cache/n1572 , \D_cache/n1571 , \D_cache/n1570 , \D_cache/n1569 ,
         \D_cache/n1568 , \D_cache/n1567 , \D_cache/n1566 , \D_cache/n1565 ,
         \D_cache/n1564 , \D_cache/n1563 , \D_cache/n1562 , \D_cache/n1561 ,
         \D_cache/n1560 , \D_cache/n1559 , \D_cache/n1558 , \D_cache/n1557 ,
         \D_cache/n1556 , \D_cache/n1555 , \D_cache/n1554 , \D_cache/n1553 ,
         \D_cache/n1552 , \D_cache/n1551 , \D_cache/n1550 , \D_cache/n1549 ,
         \D_cache/n1548 , \D_cache/n1547 , \D_cache/n1546 , \D_cache/n1545 ,
         \D_cache/n1544 , \D_cache/n1543 , \D_cache/n1542 , \D_cache/n1541 ,
         \D_cache/n1540 , \D_cache/n1539 , \D_cache/n1538 , \D_cache/n1537 ,
         \D_cache/n1536 , \D_cache/n1535 , \D_cache/n1534 , \D_cache/n1533 ,
         \D_cache/n1532 , \D_cache/n1531 , \D_cache/n1530 , \D_cache/n1529 ,
         \D_cache/n1528 , \D_cache/n1527 , \D_cache/n1526 , \D_cache/n1525 ,
         \D_cache/n1524 , \D_cache/n1523 , \D_cache/n1522 , \D_cache/n1521 ,
         \D_cache/n1520 , \D_cache/n1519 , \D_cache/n1518 , \D_cache/n1517 ,
         \D_cache/n1516 , \D_cache/n1515 , \D_cache/n1514 , \D_cache/n1513 ,
         \D_cache/n1512 , \D_cache/n1511 , \D_cache/n1510 , \D_cache/n1509 ,
         \D_cache/n1508 , \D_cache/n1507 , \D_cache/n1506 , \D_cache/n1505 ,
         \D_cache/n1504 , \D_cache/n1503 , \D_cache/n1502 , \D_cache/n1501 ,
         \D_cache/n1500 , \D_cache/n1499 , \D_cache/n1498 , \D_cache/n1497 ,
         \D_cache/n1496 , \D_cache/n1495 , \D_cache/n1494 , \D_cache/n1493 ,
         \D_cache/n1492 , \D_cache/n1491 , \D_cache/n1490 , \D_cache/n1489 ,
         \D_cache/n1488 , \D_cache/n1487 , \D_cache/n1486 , \D_cache/n1485 ,
         \D_cache/n1484 , \D_cache/n1483 , \D_cache/n1482 , \D_cache/n1481 ,
         \D_cache/n1480 , \D_cache/n1479 , \D_cache/n1478 , \D_cache/n1477 ,
         \D_cache/n1476 , \D_cache/n1475 , \D_cache/n1474 , \D_cache/n1473 ,
         \D_cache/n1472 , \D_cache/n1471 , \D_cache/n1470 , \D_cache/n1469 ,
         \D_cache/n1468 , \D_cache/n1467 , \D_cache/n1466 , \D_cache/n1465 ,
         \D_cache/n1464 , \D_cache/n1463 , \D_cache/n1462 , \D_cache/n1461 ,
         \D_cache/n1460 , \D_cache/n1459 , \D_cache/n1458 , \D_cache/n1457 ,
         \D_cache/n1456 , \D_cache/n1455 , \D_cache/n1454 , \D_cache/n1453 ,
         \D_cache/n1452 , \D_cache/n1451 , \D_cache/n1450 , \D_cache/n1449 ,
         \D_cache/n1448 , \D_cache/n1447 , \D_cache/n1446 , \D_cache/n1445 ,
         \D_cache/n1444 , \D_cache/n1443 , \D_cache/n1442 , \D_cache/n1441 ,
         \D_cache/n1440 , \D_cache/n1439 , \D_cache/n1438 , \D_cache/n1437 ,
         \D_cache/n1436 , \D_cache/n1435 , \D_cache/n1434 , \D_cache/n1433 ,
         \D_cache/n1432 , \D_cache/n1431 , \D_cache/n1430 , \D_cache/n1429 ,
         \D_cache/n1428 , \D_cache/n1427 , \D_cache/n1426 , \D_cache/n1425 ,
         \D_cache/n1424 , \D_cache/n1423 , \D_cache/n1422 , \D_cache/n1421 ,
         \D_cache/n1420 , \D_cache/n1419 , \D_cache/n1418 , \D_cache/n1417 ,
         \D_cache/n1416 , \D_cache/n1415 , \D_cache/n1414 , \D_cache/n1413 ,
         \D_cache/n1412 , \D_cache/n1411 , \D_cache/n1410 , \D_cache/n1409 ,
         \D_cache/n1408 , \D_cache/n1407 , \D_cache/n1406 , \D_cache/n1405 ,
         \D_cache/n1404 , \D_cache/n1403 , \D_cache/n1402 , \D_cache/n1401 ,
         \D_cache/n1400 , \D_cache/n1399 , \D_cache/n1398 , \D_cache/n1397 ,
         \D_cache/n1396 , \D_cache/n1395 , \D_cache/n1394 , \D_cache/n1393 ,
         \D_cache/n1392 , \D_cache/n1391 , \D_cache/n1390 , \D_cache/n1389 ,
         \D_cache/n1388 , \D_cache/n1387 , \D_cache/n1386 , \D_cache/n1385 ,
         \D_cache/n1384 , \D_cache/n1383 , \D_cache/n1382 , \D_cache/n1381 ,
         \D_cache/n1380 , \D_cache/n1379 , \D_cache/n1378 , \D_cache/n1377 ,
         \D_cache/n1376 , \D_cache/n1375 , \D_cache/n1374 , \D_cache/n1373 ,
         \D_cache/n1372 , \D_cache/n1371 , \D_cache/n1370 , \D_cache/n1369 ,
         \D_cache/n1368 , \D_cache/n1367 , \D_cache/n1366 , \D_cache/n1365 ,
         \D_cache/n1364 , \D_cache/n1363 , \D_cache/n1362 , \D_cache/n1361 ,
         \D_cache/n1360 , \D_cache/n1359 , \D_cache/n1358 , \D_cache/n1357 ,
         \D_cache/n1356 , \D_cache/n1355 , \D_cache/n1354 , \D_cache/n1353 ,
         \D_cache/n1352 , \D_cache/n1351 , \D_cache/n1350 , \D_cache/n1349 ,
         \D_cache/n1348 , \D_cache/n1347 , \D_cache/n1346 , \D_cache/n1345 ,
         \D_cache/n1344 , \D_cache/n1343 , \D_cache/n1342 , \D_cache/n1341 ,
         \D_cache/n1340 , \D_cache/n1339 , \D_cache/n1338 , \D_cache/n1337 ,
         \D_cache/n1336 , \D_cache/n1335 , \D_cache/n1334 , \D_cache/n1333 ,
         \D_cache/n1332 , \D_cache/n1331 , \D_cache/n1330 , \D_cache/n1329 ,
         \D_cache/n1328 , \D_cache/n1327 , \D_cache/n1326 , \D_cache/n1325 ,
         \D_cache/n1324 , \D_cache/n1323 , \D_cache/n1322 , \D_cache/n1321 ,
         \D_cache/n1320 , \D_cache/n1319 , \D_cache/n1318 , \D_cache/n1317 ,
         \D_cache/n1316 , \D_cache/n1315 , \D_cache/n1314 , \D_cache/n1313 ,
         \D_cache/n1312 , \D_cache/n1311 , \D_cache/n1310 , \D_cache/n1309 ,
         \D_cache/n1308 , \D_cache/n1307 , \D_cache/n1306 , \D_cache/n1305 ,
         \D_cache/n1304 , \D_cache/n1303 , \D_cache/n1302 , \D_cache/n1301 ,
         \D_cache/n1300 , \D_cache/n1299 , \D_cache/n1298 , \D_cache/n1297 ,
         \D_cache/n1296 , \D_cache/n1295 , \D_cache/n1294 , \D_cache/n1293 ,
         \D_cache/n1292 , \D_cache/n1291 , \D_cache/n1290 , \D_cache/n1289 ,
         \D_cache/n1288 , \D_cache/n1287 , \D_cache/n1286 , \D_cache/n1285 ,
         \D_cache/n1284 , \D_cache/n1283 , \D_cache/n1282 , \D_cache/n1281 ,
         \D_cache/n1280 , \D_cache/n1279 , \D_cache/n1278 , \D_cache/n1277 ,
         \D_cache/n1276 , \D_cache/n1275 , \D_cache/n1274 , \D_cache/n1273 ,
         \D_cache/n1272 , \D_cache/n1271 , \D_cache/n1270 , \D_cache/n1269 ,
         \D_cache/n1268 , \D_cache/n1267 , \D_cache/n1266 , \D_cache/n1265 ,
         \D_cache/n1264 , \D_cache/n1263 , \D_cache/n1262 , \D_cache/n1261 ,
         \D_cache/n1260 , \D_cache/n1259 , \D_cache/n1258 , \D_cache/n1257 ,
         \D_cache/n1256 , \D_cache/n1255 , \D_cache/n1254 , \D_cache/n1253 ,
         \D_cache/n1252 , \D_cache/n1251 , \D_cache/n1250 , \D_cache/n1249 ,
         \D_cache/n1248 , \D_cache/n1247 , \D_cache/n1246 , \D_cache/n1245 ,
         \D_cache/n1244 , \D_cache/n1243 , \D_cache/n1242 , \D_cache/n1241 ,
         \D_cache/n1240 , \D_cache/n1239 , \D_cache/n1238 , \D_cache/n1237 ,
         \D_cache/n1236 , \D_cache/n1235 , \D_cache/n1234 , \D_cache/n1233 ,
         \D_cache/n1232 , \D_cache/n1231 , \D_cache/n1230 , \D_cache/n1229 ,
         \D_cache/n1228 , \D_cache/n1227 , \D_cache/n1226 , \D_cache/n1225 ,
         \D_cache/n1224 , \D_cache/n1223 , \D_cache/n1222 , \D_cache/n1221 ,
         \D_cache/n1220 , \D_cache/n1219 , \D_cache/n1218 , \D_cache/n1217 ,
         \D_cache/n1216 , \D_cache/n1215 , \D_cache/n1214 , \D_cache/n1213 ,
         \D_cache/n1212 , \D_cache/n1211 , \D_cache/n1210 , \D_cache/n1209 ,
         \D_cache/n1208 , \D_cache/n1207 , \D_cache/n1206 , \D_cache/n1205 ,
         \D_cache/n1204 , \D_cache/n1203 , \D_cache/n1202 , \D_cache/n1201 ,
         \D_cache/n1200 , \D_cache/n1199 , \D_cache/n1198 , \D_cache/n1197 ,
         \D_cache/n1196 , \D_cache/n1195 , \D_cache/n1194 , \D_cache/n1193 ,
         \D_cache/n1192 , \D_cache/n1191 , \D_cache/n1190 , \D_cache/n1189 ,
         \D_cache/n1188 , \D_cache/n1187 , \D_cache/n1186 , \D_cache/n1185 ,
         \D_cache/n1184 , \D_cache/n1183 , \D_cache/n1182 , \D_cache/n1181 ,
         \D_cache/n1180 , \D_cache/n1179 , \D_cache/n1178 , \D_cache/n1177 ,
         \D_cache/n1176 , \D_cache/n1175 , \D_cache/n1174 , \D_cache/n1173 ,
         \D_cache/n1172 , \D_cache/n1171 , \D_cache/n1170 , \D_cache/n1169 ,
         \D_cache/n1168 , \D_cache/n1167 , \D_cache/n1166 , \D_cache/n1165 ,
         \D_cache/n1164 , \D_cache/n1163 , \D_cache/n1162 , \D_cache/n1161 ,
         \D_cache/n1160 , \D_cache/n1159 , \D_cache/n1158 , \D_cache/n1157 ,
         \D_cache/n1156 , \D_cache/n1155 , \D_cache/n1154 , \D_cache/n1153 ,
         \D_cache/n1152 , \D_cache/n1151 , \D_cache/n1150 , \D_cache/n1149 ,
         \D_cache/n1148 , \D_cache/n1147 , \D_cache/n1146 , \D_cache/n1145 ,
         \D_cache/n1144 , \D_cache/n1143 , \D_cache/n1142 , \D_cache/n1141 ,
         \D_cache/n1140 , \D_cache/n1139 , \D_cache/n1138 , \D_cache/n1137 ,
         \D_cache/n1136 , \D_cache/n1135 , \D_cache/n1134 , \D_cache/n1133 ,
         \D_cache/n1132 , \D_cache/n1131 , \D_cache/n1130 , \D_cache/n1129 ,
         \D_cache/n1128 , \D_cache/n1127 , \D_cache/n1126 , \D_cache/n1125 ,
         \D_cache/n1124 , \D_cache/n1123 , \D_cache/n1122 , \D_cache/n1121 ,
         \D_cache/n1120 , \D_cache/n1119 , \D_cache/n1118 , \D_cache/n1117 ,
         \D_cache/n1116 , \D_cache/n1115 , \D_cache/n1114 , \D_cache/n1113 ,
         \D_cache/n1112 , \D_cache/n1111 , \D_cache/n1110 , \D_cache/n1109 ,
         \D_cache/n1108 , \D_cache/n1107 , \D_cache/n1106 , \D_cache/n1105 ,
         \D_cache/n1104 , \D_cache/n1103 , \D_cache/n1102 , \D_cache/n1101 ,
         \D_cache/n1100 , \D_cache/n1099 , \D_cache/n1098 , \D_cache/n1097 ,
         \D_cache/n1096 , \D_cache/n1095 , \D_cache/n1094 , \D_cache/n1093 ,
         \D_cache/n1092 , \D_cache/n1091 , \D_cache/n1090 , \D_cache/n1089 ,
         \D_cache/n1088 , \D_cache/n1087 , \D_cache/n1086 , \D_cache/n1085 ,
         \D_cache/n1084 , \D_cache/n1083 , \D_cache/n1082 , \D_cache/n1081 ,
         \D_cache/n1080 , \D_cache/n1079 , \D_cache/n1078 , \D_cache/n1077 ,
         \D_cache/n1076 , \D_cache/n1075 , \D_cache/n1074 , \D_cache/n1073 ,
         \D_cache/n1072 , \D_cache/n1071 , \D_cache/n1070 , \D_cache/n1069 ,
         \D_cache/n1068 , \D_cache/n1067 , \D_cache/n1066 , \D_cache/n1065 ,
         \D_cache/n1064 , \D_cache/n1063 , \D_cache/n1062 , \D_cache/n1061 ,
         \D_cache/n1060 , \D_cache/n1059 , \D_cache/n1058 , \D_cache/n1057 ,
         \D_cache/n1056 , \D_cache/n1055 , \D_cache/n1054 , \D_cache/n1053 ,
         \D_cache/n1052 , \D_cache/n1051 , \D_cache/n1050 , \D_cache/n1049 ,
         \D_cache/n1048 , \D_cache/n1047 , \D_cache/n1046 , \D_cache/n1045 ,
         \D_cache/n1044 , \D_cache/n1043 , \D_cache/n1042 , \D_cache/n1041 ,
         \D_cache/n1040 , \D_cache/n1039 , \D_cache/n1038 , \D_cache/n1037 ,
         \D_cache/n1036 , \D_cache/n1035 , \D_cache/n1034 , \D_cache/n1033 ,
         \D_cache/n1032 , \D_cache/n1031 , \D_cache/n1030 , \D_cache/n1029 ,
         \D_cache/n1028 , \D_cache/n1027 , \D_cache/n1026 , \D_cache/n1025 ,
         \D_cache/n1024 , \D_cache/n1023 , \D_cache/n1022 , \D_cache/n1021 ,
         \D_cache/n1020 , \D_cache/n1019 , \D_cache/n1018 , \D_cache/n1017 ,
         \D_cache/n1016 , \D_cache/n1015 , \D_cache/n1014 , \D_cache/n1013 ,
         \D_cache/n1012 , \D_cache/n1011 , \D_cache/n1010 , \D_cache/n1009 ,
         \D_cache/n1008 , \D_cache/n1007 , \D_cache/n1006 , \D_cache/n1005 ,
         \D_cache/n1004 , \D_cache/n1003 , \D_cache/n1002 , \D_cache/n1001 ,
         \D_cache/n1000 , \D_cache/n999 , \D_cache/n998 , \D_cache/n997 ,
         \D_cache/n996 , \D_cache/n995 , \D_cache/n994 , \D_cache/n993 ,
         \D_cache/n992 , \D_cache/n991 , \D_cache/n990 , \D_cache/n989 ,
         \D_cache/n988 , \D_cache/n987 , \D_cache/n986 , \D_cache/n985 ,
         \D_cache/n984 , \D_cache/n983 , \D_cache/n982 , \D_cache/n981 ,
         \D_cache/n980 , \D_cache/n979 , \D_cache/n978 , \D_cache/n977 ,
         \D_cache/n976 , \D_cache/n975 , \D_cache/n974 , \D_cache/n973 ,
         \D_cache/n972 , \D_cache/n971 , \D_cache/n970 , \D_cache/n969 ,
         \D_cache/n968 , \D_cache/n967 , \D_cache/n966 , \D_cache/n965 ,
         \D_cache/n964 , \D_cache/n963 , \D_cache/n962 , \D_cache/n961 ,
         \D_cache/n960 , \D_cache/n959 , \D_cache/n958 , \D_cache/n957 ,
         \D_cache/n956 , \D_cache/n955 , \D_cache/n954 , \D_cache/n953 ,
         \D_cache/n952 , \D_cache/n951 , \D_cache/n950 , \D_cache/n949 ,
         \D_cache/n948 , \D_cache/n947 , \D_cache/n946 , \D_cache/n945 ,
         \D_cache/n944 , \D_cache/n943 , \D_cache/n942 , \D_cache/n941 ,
         \D_cache/n940 , \D_cache/n939 , \D_cache/n938 , \D_cache/n937 ,
         \D_cache/n936 , \D_cache/n935 , \D_cache/n934 , \D_cache/n933 ,
         \D_cache/n932 , \D_cache/n931 , \D_cache/n930 , \D_cache/n929 ,
         \D_cache/n928 , \D_cache/n927 , \D_cache/n926 , \D_cache/n925 ,
         \D_cache/n924 , \D_cache/n923 , \D_cache/n922 , \D_cache/n921 ,
         \D_cache/n920 , \D_cache/n919 , \D_cache/n918 , \D_cache/n917 ,
         \D_cache/n916 , \D_cache/n915 , \D_cache/n914 , \D_cache/n913 ,
         \D_cache/n912 , \D_cache/n911 , \D_cache/n910 , \D_cache/n909 ,
         \D_cache/n908 , \D_cache/n907 , \D_cache/n906 , \D_cache/n905 ,
         \D_cache/n904 , \D_cache/n903 , \D_cache/n902 , \D_cache/n901 ,
         \D_cache/n900 , \D_cache/n899 , \D_cache/n898 , \D_cache/n897 ,
         \D_cache/n896 , \D_cache/n895 , \D_cache/n894 , \D_cache/n893 ,
         \D_cache/n892 , \D_cache/n891 , \D_cache/n890 , \D_cache/n889 ,
         \D_cache/n888 , \D_cache/n887 , \D_cache/n886 , \D_cache/n885 ,
         \D_cache/n884 , \D_cache/n883 , \D_cache/n882 , \D_cache/n881 ,
         \D_cache/n880 , \D_cache/n879 , \D_cache/n878 , \D_cache/n877 ,
         \D_cache/n876 , \D_cache/n875 , \D_cache/n874 , \D_cache/n873 ,
         \D_cache/n872 , \D_cache/n871 , \D_cache/n870 , \D_cache/n869 ,
         \D_cache/n868 , \D_cache/n867 , \D_cache/n866 , \D_cache/n865 ,
         \D_cache/n864 , \D_cache/n863 , \D_cache/n862 , \D_cache/n861 ,
         \D_cache/n860 , \D_cache/n859 , \D_cache/n858 , \D_cache/n857 ,
         \D_cache/n856 , \D_cache/n855 , \D_cache/n854 , \D_cache/n853 ,
         \D_cache/n852 , \D_cache/n851 , \D_cache/n850 , \D_cache/n849 ,
         \D_cache/n848 , \D_cache/n847 , \D_cache/n846 , \D_cache/n845 ,
         \D_cache/n844 , \D_cache/n843 , \D_cache/n842 , \D_cache/n841 ,
         \D_cache/n840 , \D_cache/n839 , \D_cache/n838 , \D_cache/n837 ,
         \D_cache/n836 , \D_cache/n835 , \D_cache/n834 , \D_cache/n833 ,
         \D_cache/n832 , \D_cache/n831 , \D_cache/n830 , \D_cache/n829 ,
         \D_cache/n828 , \D_cache/n827 , \D_cache/n826 , \D_cache/n825 ,
         \D_cache/n824 , \D_cache/n823 , \D_cache/n822 , \D_cache/n821 ,
         \D_cache/n820 , \D_cache/n819 , \D_cache/n818 , \D_cache/n817 ,
         \D_cache/n816 , \D_cache/n815 , \D_cache/n814 , \D_cache/n813 ,
         \D_cache/n812 , \D_cache/n811 , \D_cache/n810 , \D_cache/n809 ,
         \D_cache/n808 , \D_cache/n807 , \D_cache/n806 , \D_cache/n805 ,
         \D_cache/n804 , \D_cache/n803 , \D_cache/n802 , \D_cache/n801 ,
         \D_cache/n800 , \D_cache/n799 , \D_cache/n798 , \D_cache/n797 ,
         \D_cache/n796 , \D_cache/n795 , \D_cache/n794 , \D_cache/n793 ,
         \D_cache/n792 , \D_cache/n791 , \D_cache/n790 , \D_cache/n789 ,
         \D_cache/n788 , \D_cache/n787 , \D_cache/n786 , \D_cache/n785 ,
         \D_cache/n784 , \D_cache/n783 , \D_cache/n782 , \D_cache/n781 ,
         \D_cache/n780 , \D_cache/n779 , \D_cache/n778 , \D_cache/n777 ,
         \D_cache/n776 , \D_cache/n775 , \D_cache/n774 , \D_cache/n773 ,
         \D_cache/n772 , \D_cache/n771 , \D_cache/n770 , \D_cache/n769 ,
         \D_cache/n768 , \D_cache/n767 , \D_cache/n766 , \D_cache/n765 ,
         \D_cache/n764 , \D_cache/n763 , \D_cache/n762 , \D_cache/n761 ,
         \D_cache/n760 , \D_cache/n759 , \D_cache/n758 , \D_cache/n757 ,
         \D_cache/n756 , \D_cache/n755 , \D_cache/n754 , \D_cache/n753 ,
         \D_cache/n752 , \D_cache/n751 , \D_cache/n750 , \D_cache/n749 ,
         \D_cache/n748 , \D_cache/n747 , \D_cache/n746 , \D_cache/n745 ,
         \D_cache/n744 , \D_cache/n743 , \D_cache/n742 , \D_cache/n741 ,
         \D_cache/n740 , \D_cache/n739 , \D_cache/n738 , \D_cache/n737 ,
         \D_cache/n736 , \D_cache/n735 , \D_cache/n734 , \D_cache/n733 ,
         \D_cache/n732 , \D_cache/n731 , \D_cache/n730 , \D_cache/n729 ,
         \D_cache/n728 , \D_cache/n727 , \D_cache/n726 , \D_cache/n725 ,
         \D_cache/n724 , \D_cache/n723 , \D_cache/n722 , \D_cache/n721 ,
         \D_cache/n720 , \D_cache/n719 , \D_cache/n718 , \D_cache/n717 ,
         \D_cache/n716 , \D_cache/n715 , \D_cache/n714 , \D_cache/n713 ,
         \D_cache/n712 , \D_cache/n711 , \D_cache/n710 , \D_cache/n709 ,
         \D_cache/n708 , \D_cache/n707 , \D_cache/n706 , \D_cache/n705 ,
         \D_cache/n704 , \D_cache/n703 , \D_cache/n702 , \D_cache/n701 ,
         \D_cache/n700 , \D_cache/n699 , \D_cache/n698 , \D_cache/n697 ,
         \D_cache/n696 , \D_cache/n695 , \D_cache/n694 , \D_cache/n693 ,
         \D_cache/n692 , \D_cache/n691 , \D_cache/n690 , \D_cache/n689 ,
         \D_cache/n688 , \D_cache/n687 , \D_cache/n686 , \D_cache/n685 ,
         \D_cache/n684 , \D_cache/n683 , \D_cache/n682 , \D_cache/n681 ,
         \D_cache/n680 , \D_cache/n679 , \D_cache/n678 , \D_cache/n677 ,
         \D_cache/n676 , \D_cache/n675 , \D_cache/n674 , \D_cache/n673 ,
         \D_cache/n672 , \D_cache/n671 , \D_cache/n670 , \D_cache/n669 ,
         \D_cache/n668 , \D_cache/n667 , \D_cache/n666 , \D_cache/n665 ,
         \D_cache/n664 , \D_cache/n663 , \D_cache/n662 , \D_cache/n661 ,
         \D_cache/n660 , \D_cache/n659 , \D_cache/n658 , \D_cache/n657 ,
         \D_cache/n656 , \D_cache/n655 , \D_cache/n654 , \D_cache/n653 ,
         \D_cache/n652 , \D_cache/n651 , \D_cache/n650 , \D_cache/n649 ,
         \D_cache/n648 , \D_cache/n647 , \D_cache/n646 , \D_cache/n645 ,
         \D_cache/n644 , \D_cache/n643 , \D_cache/n642 , \D_cache/n641 ,
         \D_cache/n640 , \D_cache/n639 , \D_cache/n638 , \D_cache/n637 ,
         \D_cache/n636 , \D_cache/n635 , \D_cache/n634 , \D_cache/n633 ,
         \D_cache/n632 , \D_cache/n631 , \D_cache/n630 , \D_cache/n629 ,
         \D_cache/n628 , \D_cache/n627 , \D_cache/n626 , \D_cache/n625 ,
         \D_cache/n624 , \D_cache/n623 , \D_cache/n622 , \D_cache/n621 ,
         \D_cache/n620 , \D_cache/n619 , \D_cache/n618 , \D_cache/n617 ,
         \D_cache/n616 , \D_cache/n615 , \D_cache/n614 , \D_cache/n613 ,
         \D_cache/n612 , \D_cache/n611 , \D_cache/n610 , \D_cache/n609 ,
         \D_cache/n608 , \D_cache/n607 , \D_cache/n606 , \D_cache/n605 ,
         \D_cache/n604 , \D_cache/n603 , \D_cache/n602 , \D_cache/n601 ,
         \D_cache/n600 , \D_cache/n599 , \D_cache/n598 , \D_cache/n597 ,
         \D_cache/n596 , \D_cache/n595 , \D_cache/n594 , \D_cache/n593 ,
         \D_cache/n592 , \D_cache/n591 , \D_cache/n590 , \D_cache/n589 ,
         \D_cache/n588 , \D_cache/n587 , \D_cache/n586 , \D_cache/n585 ,
         \D_cache/n584 , \D_cache/n583 , \D_cache/n582 , \D_cache/n581 ,
         \D_cache/n580 , \D_cache/n579 , \D_cache/n578 , \D_cache/n577 ,
         \D_cache/n576 , \D_cache/n575 , \D_cache/n574 , \D_cache/n573 ,
         \D_cache/n572 , \D_cache/n571 , \D_cache/n570 , \D_cache/n569 ,
         \D_cache/n568 , \D_cache/n567 , \D_cache/n566 , \D_cache/n565 ,
         \D_cache/n564 , \D_cache/n563 , \D_cache/n562 , \D_cache/n561 ,
         \D_cache/n560 , \D_cache/n559 , \D_cache/n558 , \D_cache/n557 ,
         \D_cache/cache[7][0] , \D_cache/cache[7][1] , \D_cache/cache[7][2] ,
         \D_cache/cache[7][3] , \D_cache/cache[7][4] , \D_cache/cache[7][5] ,
         \D_cache/cache[7][6] , \D_cache/cache[7][7] , \D_cache/cache[7][8] ,
         \D_cache/cache[7][9] , \D_cache/cache[7][10] , \D_cache/cache[7][11] ,
         \D_cache/cache[7][12] , \D_cache/cache[7][13] ,
         \D_cache/cache[7][14] , \D_cache/cache[7][15] ,
         \D_cache/cache[7][16] , \D_cache/cache[7][17] ,
         \D_cache/cache[7][18] , \D_cache/cache[7][19] ,
         \D_cache/cache[7][20] , \D_cache/cache[7][21] ,
         \D_cache/cache[7][22] , \D_cache/cache[7][23] ,
         \D_cache/cache[7][24] , \D_cache/cache[7][25] ,
         \D_cache/cache[7][26] , \D_cache/cache[7][27] ,
         \D_cache/cache[7][28] , \D_cache/cache[7][29] ,
         \D_cache/cache[7][30] , \D_cache/cache[7][31] ,
         \D_cache/cache[7][32] , \D_cache/cache[7][33] ,
         \D_cache/cache[7][34] , \D_cache/cache[7][35] ,
         \D_cache/cache[7][36] , \D_cache/cache[7][37] ,
         \D_cache/cache[7][38] , \D_cache/cache[7][39] ,
         \D_cache/cache[7][40] , \D_cache/cache[7][41] ,
         \D_cache/cache[7][42] , \D_cache/cache[7][43] ,
         \D_cache/cache[7][44] , \D_cache/cache[7][45] ,
         \D_cache/cache[7][46] , \D_cache/cache[7][47] ,
         \D_cache/cache[7][48] , \D_cache/cache[7][49] ,
         \D_cache/cache[7][50] , \D_cache/cache[7][51] ,
         \D_cache/cache[7][52] , \D_cache/cache[7][53] ,
         \D_cache/cache[7][54] , \D_cache/cache[7][55] ,
         \D_cache/cache[7][56] , \D_cache/cache[7][57] ,
         \D_cache/cache[7][58] , \D_cache/cache[7][59] ,
         \D_cache/cache[7][60] , \D_cache/cache[7][61] ,
         \D_cache/cache[7][62] , \D_cache/cache[7][63] ,
         \D_cache/cache[7][64] , \D_cache/cache[7][65] ,
         \D_cache/cache[7][66] , \D_cache/cache[7][67] ,
         \D_cache/cache[7][68] , \D_cache/cache[7][69] ,
         \D_cache/cache[7][70] , \D_cache/cache[7][71] ,
         \D_cache/cache[7][72] , \D_cache/cache[7][73] ,
         \D_cache/cache[7][74] , \D_cache/cache[7][75] ,
         \D_cache/cache[7][76] , \D_cache/cache[7][77] ,
         \D_cache/cache[7][78] , \D_cache/cache[7][79] ,
         \D_cache/cache[7][80] , \D_cache/cache[7][81] ,
         \D_cache/cache[7][82] , \D_cache/cache[7][83] ,
         \D_cache/cache[7][84] , \D_cache/cache[7][85] ,
         \D_cache/cache[7][86] , \D_cache/cache[7][87] ,
         \D_cache/cache[7][88] , \D_cache/cache[7][89] ,
         \D_cache/cache[7][90] , \D_cache/cache[7][91] ,
         \D_cache/cache[7][92] , \D_cache/cache[7][93] ,
         \D_cache/cache[7][94] , \D_cache/cache[7][95] ,
         \D_cache/cache[7][96] , \D_cache/cache[7][97] ,
         \D_cache/cache[7][98] , \D_cache/cache[7][99] ,
         \D_cache/cache[7][100] , \D_cache/cache[7][101] ,
         \D_cache/cache[7][102] , \D_cache/cache[7][103] ,
         \D_cache/cache[7][104] , \D_cache/cache[7][105] ,
         \D_cache/cache[7][106] , \D_cache/cache[7][107] ,
         \D_cache/cache[7][108] , \D_cache/cache[7][109] ,
         \D_cache/cache[7][110] , \D_cache/cache[7][111] ,
         \D_cache/cache[7][112] , \D_cache/cache[7][113] ,
         \D_cache/cache[7][114] , \D_cache/cache[7][115] ,
         \D_cache/cache[7][116] , \D_cache/cache[7][117] ,
         \D_cache/cache[7][118] , \D_cache/cache[7][119] ,
         \D_cache/cache[7][120] , \D_cache/cache[7][121] ,
         \D_cache/cache[7][122] , \D_cache/cache[7][123] ,
         \D_cache/cache[7][124] , \D_cache/cache[7][125] ,
         \D_cache/cache[7][126] , \D_cache/cache[7][127] ,
         \D_cache/cache[7][128] , \D_cache/cache[7][129] ,
         \D_cache/cache[7][130] , \D_cache/cache[7][131] ,
         \D_cache/cache[7][132] , \D_cache/cache[7][133] ,
         \D_cache/cache[7][134] , \D_cache/cache[7][135] ,
         \D_cache/cache[7][136] , \D_cache/cache[7][137] ,
         \D_cache/cache[7][138] , \D_cache/cache[7][139] ,
         \D_cache/cache[7][140] , \D_cache/cache[7][141] ,
         \D_cache/cache[7][142] , \D_cache/cache[7][143] ,
         \D_cache/cache[7][144] , \D_cache/cache[7][145] ,
         \D_cache/cache[7][146] , \D_cache/cache[7][147] ,
         \D_cache/cache[7][148] , \D_cache/cache[7][149] ,
         \D_cache/cache[7][150] , \D_cache/cache[7][151] ,
         \D_cache/cache[7][152] , \D_cache/cache[7][153] ,
         \D_cache/cache[7][154] , \D_cache/cache[6][0] , \D_cache/cache[6][1] ,
         \D_cache/cache[6][2] , \D_cache/cache[6][3] , \D_cache/cache[6][4] ,
         \D_cache/cache[6][5] , \D_cache/cache[6][6] , \D_cache/cache[6][7] ,
         \D_cache/cache[6][8] , \D_cache/cache[6][9] , \D_cache/cache[6][10] ,
         \D_cache/cache[6][11] , \D_cache/cache[6][12] ,
         \D_cache/cache[6][13] , \D_cache/cache[6][14] ,
         \D_cache/cache[6][15] , \D_cache/cache[6][16] ,
         \D_cache/cache[6][17] , \D_cache/cache[6][18] ,
         \D_cache/cache[6][19] , \D_cache/cache[6][20] ,
         \D_cache/cache[6][21] , \D_cache/cache[6][22] ,
         \D_cache/cache[6][23] , \D_cache/cache[6][24] ,
         \D_cache/cache[6][25] , \D_cache/cache[6][26] ,
         \D_cache/cache[6][27] , \D_cache/cache[6][28] ,
         \D_cache/cache[6][29] , \D_cache/cache[6][30] ,
         \D_cache/cache[6][31] , \D_cache/cache[6][32] ,
         \D_cache/cache[6][33] , \D_cache/cache[6][34] ,
         \D_cache/cache[6][35] , \D_cache/cache[6][36] ,
         \D_cache/cache[6][37] , \D_cache/cache[6][38] ,
         \D_cache/cache[6][39] , \D_cache/cache[6][40] ,
         \D_cache/cache[6][41] , \D_cache/cache[6][42] ,
         \D_cache/cache[6][43] , \D_cache/cache[6][44] ,
         \D_cache/cache[6][45] , \D_cache/cache[6][46] ,
         \D_cache/cache[6][47] , \D_cache/cache[6][48] ,
         \D_cache/cache[6][49] , \D_cache/cache[6][50] ,
         \D_cache/cache[6][51] , \D_cache/cache[6][52] ,
         \D_cache/cache[6][53] , \D_cache/cache[6][54] ,
         \D_cache/cache[6][55] , \D_cache/cache[6][56] ,
         \D_cache/cache[6][57] , \D_cache/cache[6][58] ,
         \D_cache/cache[6][59] , \D_cache/cache[6][60] ,
         \D_cache/cache[6][61] , \D_cache/cache[6][62] ,
         \D_cache/cache[6][63] , \D_cache/cache[6][64] ,
         \D_cache/cache[6][65] , \D_cache/cache[6][66] ,
         \D_cache/cache[6][67] , \D_cache/cache[6][68] ,
         \D_cache/cache[6][69] , \D_cache/cache[6][70] ,
         \D_cache/cache[6][71] , \D_cache/cache[6][72] ,
         \D_cache/cache[6][73] , \D_cache/cache[6][74] ,
         \D_cache/cache[6][75] , \D_cache/cache[6][76] ,
         \D_cache/cache[6][77] , \D_cache/cache[6][78] ,
         \D_cache/cache[6][79] , \D_cache/cache[6][80] ,
         \D_cache/cache[6][81] , \D_cache/cache[6][82] ,
         \D_cache/cache[6][83] , \D_cache/cache[6][84] ,
         \D_cache/cache[6][85] , \D_cache/cache[6][86] ,
         \D_cache/cache[6][87] , \D_cache/cache[6][88] ,
         \D_cache/cache[6][89] , \D_cache/cache[6][90] ,
         \D_cache/cache[6][91] , \D_cache/cache[6][92] ,
         \D_cache/cache[6][93] , \D_cache/cache[6][94] ,
         \D_cache/cache[6][95] , \D_cache/cache[6][96] ,
         \D_cache/cache[6][97] , \D_cache/cache[6][98] ,
         \D_cache/cache[6][99] , \D_cache/cache[6][100] ,
         \D_cache/cache[6][101] , \D_cache/cache[6][102] ,
         \D_cache/cache[6][103] , \D_cache/cache[6][104] ,
         \D_cache/cache[6][105] , \D_cache/cache[6][106] ,
         \D_cache/cache[6][107] , \D_cache/cache[6][108] ,
         \D_cache/cache[6][109] , \D_cache/cache[6][110] ,
         \D_cache/cache[6][111] , \D_cache/cache[6][112] ,
         \D_cache/cache[6][113] , \D_cache/cache[6][114] ,
         \D_cache/cache[6][115] , \D_cache/cache[6][116] ,
         \D_cache/cache[6][117] , \D_cache/cache[6][118] ,
         \D_cache/cache[6][119] , \D_cache/cache[6][120] ,
         \D_cache/cache[6][121] , \D_cache/cache[6][122] ,
         \D_cache/cache[6][123] , \D_cache/cache[6][124] ,
         \D_cache/cache[6][125] , \D_cache/cache[6][126] ,
         \D_cache/cache[6][127] , \D_cache/cache[6][128] ,
         \D_cache/cache[6][129] , \D_cache/cache[6][130] ,
         \D_cache/cache[6][131] , \D_cache/cache[6][132] ,
         \D_cache/cache[6][133] , \D_cache/cache[6][134] ,
         \D_cache/cache[6][135] , \D_cache/cache[6][136] ,
         \D_cache/cache[6][137] , \D_cache/cache[6][138] ,
         \D_cache/cache[6][139] , \D_cache/cache[6][140] ,
         \D_cache/cache[6][141] , \D_cache/cache[6][142] ,
         \D_cache/cache[6][143] , \D_cache/cache[6][144] ,
         \D_cache/cache[6][145] , \D_cache/cache[6][146] ,
         \D_cache/cache[6][147] , \D_cache/cache[6][148] ,
         \D_cache/cache[6][149] , \D_cache/cache[6][150] ,
         \D_cache/cache[6][151] , \D_cache/cache[6][152] ,
         \D_cache/cache[6][153] , \D_cache/cache[6][154] ,
         \D_cache/cache[5][0] , \D_cache/cache[5][1] , \D_cache/cache[5][2] ,
         \D_cache/cache[5][3] , \D_cache/cache[5][4] , \D_cache/cache[5][5] ,
         \D_cache/cache[5][6] , \D_cache/cache[5][7] , \D_cache/cache[5][8] ,
         \D_cache/cache[5][9] , \D_cache/cache[5][10] , \D_cache/cache[5][11] ,
         \D_cache/cache[5][12] , \D_cache/cache[5][13] ,
         \D_cache/cache[5][14] , \D_cache/cache[5][15] ,
         \D_cache/cache[5][16] , \D_cache/cache[5][17] ,
         \D_cache/cache[5][18] , \D_cache/cache[5][19] ,
         \D_cache/cache[5][20] , \D_cache/cache[5][21] ,
         \D_cache/cache[5][22] , \D_cache/cache[5][23] ,
         \D_cache/cache[5][24] , \D_cache/cache[5][25] ,
         \D_cache/cache[5][26] , \D_cache/cache[5][27] ,
         \D_cache/cache[5][28] , \D_cache/cache[5][29] ,
         \D_cache/cache[5][30] , \D_cache/cache[5][31] ,
         \D_cache/cache[5][32] , \D_cache/cache[5][33] ,
         \D_cache/cache[5][34] , \D_cache/cache[5][35] ,
         \D_cache/cache[5][36] , \D_cache/cache[5][37] ,
         \D_cache/cache[5][38] , \D_cache/cache[5][39] ,
         \D_cache/cache[5][40] , \D_cache/cache[5][41] ,
         \D_cache/cache[5][42] , \D_cache/cache[5][43] ,
         \D_cache/cache[5][44] , \D_cache/cache[5][45] ,
         \D_cache/cache[5][46] , \D_cache/cache[5][47] ,
         \D_cache/cache[5][48] , \D_cache/cache[5][49] ,
         \D_cache/cache[5][50] , \D_cache/cache[5][51] ,
         \D_cache/cache[5][52] , \D_cache/cache[5][53] ,
         \D_cache/cache[5][54] , \D_cache/cache[5][55] ,
         \D_cache/cache[5][56] , \D_cache/cache[5][57] ,
         \D_cache/cache[5][58] , \D_cache/cache[5][59] ,
         \D_cache/cache[5][60] , \D_cache/cache[5][61] ,
         \D_cache/cache[5][62] , \D_cache/cache[5][63] ,
         \D_cache/cache[5][64] , \D_cache/cache[5][65] ,
         \D_cache/cache[5][66] , \D_cache/cache[5][67] ,
         \D_cache/cache[5][68] , \D_cache/cache[5][69] ,
         \D_cache/cache[5][70] , \D_cache/cache[5][71] ,
         \D_cache/cache[5][72] , \D_cache/cache[5][73] ,
         \D_cache/cache[5][74] , \D_cache/cache[5][75] ,
         \D_cache/cache[5][76] , \D_cache/cache[5][77] ,
         \D_cache/cache[5][78] , \D_cache/cache[5][79] ,
         \D_cache/cache[5][80] , \D_cache/cache[5][81] ,
         \D_cache/cache[5][82] , \D_cache/cache[5][83] ,
         \D_cache/cache[5][84] , \D_cache/cache[5][85] ,
         \D_cache/cache[5][86] , \D_cache/cache[5][87] ,
         \D_cache/cache[5][88] , \D_cache/cache[5][89] ,
         \D_cache/cache[5][90] , \D_cache/cache[5][91] ,
         \D_cache/cache[5][92] , \D_cache/cache[5][93] ,
         \D_cache/cache[5][94] , \D_cache/cache[5][95] ,
         \D_cache/cache[5][96] , \D_cache/cache[5][97] ,
         \D_cache/cache[5][98] , \D_cache/cache[5][99] ,
         \D_cache/cache[5][100] , \D_cache/cache[5][101] ,
         \D_cache/cache[5][102] , \D_cache/cache[5][103] ,
         \D_cache/cache[5][104] , \D_cache/cache[5][105] ,
         \D_cache/cache[5][106] , \D_cache/cache[5][107] ,
         \D_cache/cache[5][108] , \D_cache/cache[5][109] ,
         \D_cache/cache[5][110] , \D_cache/cache[5][111] ,
         \D_cache/cache[5][112] , \D_cache/cache[5][113] ,
         \D_cache/cache[5][114] , \D_cache/cache[5][115] ,
         \D_cache/cache[5][116] , \D_cache/cache[5][117] ,
         \D_cache/cache[5][118] , \D_cache/cache[5][119] ,
         \D_cache/cache[5][120] , \D_cache/cache[5][121] ,
         \D_cache/cache[5][122] , \D_cache/cache[5][123] ,
         \D_cache/cache[5][124] , \D_cache/cache[5][125] ,
         \D_cache/cache[5][126] , \D_cache/cache[5][127] ,
         \D_cache/cache[5][128] , \D_cache/cache[5][129] ,
         \D_cache/cache[5][130] , \D_cache/cache[5][131] ,
         \D_cache/cache[5][132] , \D_cache/cache[5][133] ,
         \D_cache/cache[5][134] , \D_cache/cache[5][135] ,
         \D_cache/cache[5][136] , \D_cache/cache[5][137] ,
         \D_cache/cache[5][138] , \D_cache/cache[5][139] ,
         \D_cache/cache[5][140] , \D_cache/cache[5][141] ,
         \D_cache/cache[5][142] , \D_cache/cache[5][143] ,
         \D_cache/cache[5][144] , \D_cache/cache[5][145] ,
         \D_cache/cache[5][146] , \D_cache/cache[5][147] ,
         \D_cache/cache[5][148] , \D_cache/cache[5][149] ,
         \D_cache/cache[5][150] , \D_cache/cache[5][151] ,
         \D_cache/cache[5][152] , \D_cache/cache[5][153] ,
         \D_cache/cache[5][154] , \D_cache/cache[4][0] , \D_cache/cache[4][1] ,
         \D_cache/cache[4][2] , \D_cache/cache[4][3] , \D_cache/cache[4][4] ,
         \D_cache/cache[4][5] , \D_cache/cache[4][6] , \D_cache/cache[4][7] ,
         \D_cache/cache[4][8] , \D_cache/cache[4][9] , \D_cache/cache[4][10] ,
         \D_cache/cache[4][11] , \D_cache/cache[4][12] ,
         \D_cache/cache[4][13] , \D_cache/cache[4][14] ,
         \D_cache/cache[4][15] , \D_cache/cache[4][16] ,
         \D_cache/cache[4][17] , \D_cache/cache[4][18] ,
         \D_cache/cache[4][19] , \D_cache/cache[4][20] ,
         \D_cache/cache[4][21] , \D_cache/cache[4][22] ,
         \D_cache/cache[4][23] , \D_cache/cache[4][24] ,
         \D_cache/cache[4][25] , \D_cache/cache[4][26] ,
         \D_cache/cache[4][27] , \D_cache/cache[4][28] ,
         \D_cache/cache[4][29] , \D_cache/cache[4][30] ,
         \D_cache/cache[4][31] , \D_cache/cache[4][32] ,
         \D_cache/cache[4][33] , \D_cache/cache[4][34] ,
         \D_cache/cache[4][35] , \D_cache/cache[4][36] ,
         \D_cache/cache[4][37] , \D_cache/cache[4][38] ,
         \D_cache/cache[4][39] , \D_cache/cache[4][40] ,
         \D_cache/cache[4][41] , \D_cache/cache[4][42] ,
         \D_cache/cache[4][43] , \D_cache/cache[4][44] ,
         \D_cache/cache[4][45] , \D_cache/cache[4][46] ,
         \D_cache/cache[4][47] , \D_cache/cache[4][48] ,
         \D_cache/cache[4][49] , \D_cache/cache[4][50] ,
         \D_cache/cache[4][51] , \D_cache/cache[4][52] ,
         \D_cache/cache[4][53] , \D_cache/cache[4][54] ,
         \D_cache/cache[4][55] , \D_cache/cache[4][56] ,
         \D_cache/cache[4][57] , \D_cache/cache[4][58] ,
         \D_cache/cache[4][59] , \D_cache/cache[4][60] ,
         \D_cache/cache[4][61] , \D_cache/cache[4][62] ,
         \D_cache/cache[4][63] , \D_cache/cache[4][64] ,
         \D_cache/cache[4][65] , \D_cache/cache[4][66] ,
         \D_cache/cache[4][67] , \D_cache/cache[4][68] ,
         \D_cache/cache[4][69] , \D_cache/cache[4][70] ,
         \D_cache/cache[4][71] , \D_cache/cache[4][72] ,
         \D_cache/cache[4][73] , \D_cache/cache[4][74] ,
         \D_cache/cache[4][75] , \D_cache/cache[4][76] ,
         \D_cache/cache[4][77] , \D_cache/cache[4][78] ,
         \D_cache/cache[4][79] , \D_cache/cache[4][80] ,
         \D_cache/cache[4][81] , \D_cache/cache[4][82] ,
         \D_cache/cache[4][83] , \D_cache/cache[4][84] ,
         \D_cache/cache[4][85] , \D_cache/cache[4][86] ,
         \D_cache/cache[4][87] , \D_cache/cache[4][88] ,
         \D_cache/cache[4][89] , \D_cache/cache[4][90] ,
         \D_cache/cache[4][91] , \D_cache/cache[4][92] ,
         \D_cache/cache[4][93] , \D_cache/cache[4][94] ,
         \D_cache/cache[4][95] , \D_cache/cache[4][96] ,
         \D_cache/cache[4][97] , \D_cache/cache[4][98] ,
         \D_cache/cache[4][99] , \D_cache/cache[4][100] ,
         \D_cache/cache[4][101] , \D_cache/cache[4][102] ,
         \D_cache/cache[4][103] , \D_cache/cache[4][104] ,
         \D_cache/cache[4][105] , \D_cache/cache[4][106] ,
         \D_cache/cache[4][107] , \D_cache/cache[4][108] ,
         \D_cache/cache[4][109] , \D_cache/cache[4][110] ,
         \D_cache/cache[4][111] , \D_cache/cache[4][112] ,
         \D_cache/cache[4][113] , \D_cache/cache[4][114] ,
         \D_cache/cache[4][115] , \D_cache/cache[4][116] ,
         \D_cache/cache[4][117] , \D_cache/cache[4][118] ,
         \D_cache/cache[4][119] , \D_cache/cache[4][120] ,
         \D_cache/cache[4][121] , \D_cache/cache[4][122] ,
         \D_cache/cache[4][123] , \D_cache/cache[4][124] ,
         \D_cache/cache[4][125] , \D_cache/cache[4][126] ,
         \D_cache/cache[4][127] , \D_cache/cache[4][128] ,
         \D_cache/cache[4][129] , \D_cache/cache[4][130] ,
         \D_cache/cache[4][131] , \D_cache/cache[4][132] ,
         \D_cache/cache[4][133] , \D_cache/cache[4][134] ,
         \D_cache/cache[4][135] , \D_cache/cache[4][136] ,
         \D_cache/cache[4][137] , \D_cache/cache[4][138] ,
         \D_cache/cache[4][139] , \D_cache/cache[4][140] ,
         \D_cache/cache[4][141] , \D_cache/cache[4][142] ,
         \D_cache/cache[4][143] , \D_cache/cache[4][144] ,
         \D_cache/cache[4][145] , \D_cache/cache[4][146] ,
         \D_cache/cache[4][147] , \D_cache/cache[4][148] ,
         \D_cache/cache[4][149] , \D_cache/cache[4][150] ,
         \D_cache/cache[4][151] , \D_cache/cache[4][152] ,
         \D_cache/cache[4][153] , \D_cache/cache[4][154] ,
         \D_cache/cache[3][0] , \D_cache/cache[3][1] , \D_cache/cache[3][2] ,
         \D_cache/cache[3][3] , \D_cache/cache[3][4] , \D_cache/cache[3][5] ,
         \D_cache/cache[3][6] , \D_cache/cache[3][7] , \D_cache/cache[3][8] ,
         \D_cache/cache[3][9] , \D_cache/cache[3][10] , \D_cache/cache[3][11] ,
         \D_cache/cache[3][12] , \D_cache/cache[3][13] ,
         \D_cache/cache[3][14] , \D_cache/cache[3][15] ,
         \D_cache/cache[3][16] , \D_cache/cache[3][17] ,
         \D_cache/cache[3][18] , \D_cache/cache[3][19] ,
         \D_cache/cache[3][20] , \D_cache/cache[3][21] ,
         \D_cache/cache[3][22] , \D_cache/cache[3][23] ,
         \D_cache/cache[3][24] , \D_cache/cache[3][25] ,
         \D_cache/cache[3][26] , \D_cache/cache[3][27] ,
         \D_cache/cache[3][28] , \D_cache/cache[3][29] ,
         \D_cache/cache[3][30] , \D_cache/cache[3][31] ,
         \D_cache/cache[3][32] , \D_cache/cache[3][33] ,
         \D_cache/cache[3][34] , \D_cache/cache[3][35] ,
         \D_cache/cache[3][36] , \D_cache/cache[3][37] ,
         \D_cache/cache[3][38] , \D_cache/cache[3][39] ,
         \D_cache/cache[3][40] , \D_cache/cache[3][41] ,
         \D_cache/cache[3][42] , \D_cache/cache[3][43] ,
         \D_cache/cache[3][44] , \D_cache/cache[3][45] ,
         \D_cache/cache[3][46] , \D_cache/cache[3][47] ,
         \D_cache/cache[3][48] , \D_cache/cache[3][49] ,
         \D_cache/cache[3][50] , \D_cache/cache[3][51] ,
         \D_cache/cache[3][52] , \D_cache/cache[3][53] ,
         \D_cache/cache[3][54] , \D_cache/cache[3][55] ,
         \D_cache/cache[3][56] , \D_cache/cache[3][57] ,
         \D_cache/cache[3][58] , \D_cache/cache[3][59] ,
         \D_cache/cache[3][60] , \D_cache/cache[3][61] ,
         \D_cache/cache[3][62] , \D_cache/cache[3][63] ,
         \D_cache/cache[3][64] , \D_cache/cache[3][65] ,
         \D_cache/cache[3][66] , \D_cache/cache[3][67] ,
         \D_cache/cache[3][68] , \D_cache/cache[3][69] ,
         \D_cache/cache[3][70] , \D_cache/cache[3][71] ,
         \D_cache/cache[3][72] , \D_cache/cache[3][73] ,
         \D_cache/cache[3][74] , \D_cache/cache[3][75] ,
         \D_cache/cache[3][76] , \D_cache/cache[3][77] ,
         \D_cache/cache[3][78] , \D_cache/cache[3][79] ,
         \D_cache/cache[3][80] , \D_cache/cache[3][81] ,
         \D_cache/cache[3][82] , \D_cache/cache[3][83] ,
         \D_cache/cache[3][84] , \D_cache/cache[3][85] ,
         \D_cache/cache[3][86] , \D_cache/cache[3][87] ,
         \D_cache/cache[3][88] , \D_cache/cache[3][89] ,
         \D_cache/cache[3][90] , \D_cache/cache[3][91] ,
         \D_cache/cache[3][92] , \D_cache/cache[3][93] ,
         \D_cache/cache[3][94] , \D_cache/cache[3][95] ,
         \D_cache/cache[3][96] , \D_cache/cache[3][97] ,
         \D_cache/cache[3][98] , \D_cache/cache[3][99] ,
         \D_cache/cache[3][100] , \D_cache/cache[3][101] ,
         \D_cache/cache[3][102] , \D_cache/cache[3][103] ,
         \D_cache/cache[3][104] , \D_cache/cache[3][105] ,
         \D_cache/cache[3][106] , \D_cache/cache[3][107] ,
         \D_cache/cache[3][108] , \D_cache/cache[3][109] ,
         \D_cache/cache[3][110] , \D_cache/cache[3][111] ,
         \D_cache/cache[3][112] , \D_cache/cache[3][113] ,
         \D_cache/cache[3][114] , \D_cache/cache[3][115] ,
         \D_cache/cache[3][116] , \D_cache/cache[3][117] ,
         \D_cache/cache[3][118] , \D_cache/cache[3][119] ,
         \D_cache/cache[3][120] , \D_cache/cache[3][121] ,
         \D_cache/cache[3][122] , \D_cache/cache[3][123] ,
         \D_cache/cache[3][124] , \D_cache/cache[3][125] ,
         \D_cache/cache[3][126] , \D_cache/cache[3][127] ,
         \D_cache/cache[3][128] , \D_cache/cache[3][129] ,
         \D_cache/cache[3][130] , \D_cache/cache[3][131] ,
         \D_cache/cache[3][132] , \D_cache/cache[3][133] ,
         \D_cache/cache[3][134] , \D_cache/cache[3][135] ,
         \D_cache/cache[3][136] , \D_cache/cache[3][137] ,
         \D_cache/cache[3][138] , \D_cache/cache[3][139] ,
         \D_cache/cache[3][140] , \D_cache/cache[3][141] ,
         \D_cache/cache[3][142] , \D_cache/cache[3][143] ,
         \D_cache/cache[3][144] , \D_cache/cache[3][145] ,
         \D_cache/cache[3][146] , \D_cache/cache[3][147] ,
         \D_cache/cache[3][148] , \D_cache/cache[3][149] ,
         \D_cache/cache[3][150] , \D_cache/cache[3][151] ,
         \D_cache/cache[3][152] , \D_cache/cache[3][153] ,
         \D_cache/cache[3][154] , \D_cache/cache[2][0] , \D_cache/cache[2][1] ,
         \D_cache/cache[2][2] , \D_cache/cache[2][3] , \D_cache/cache[2][4] ,
         \D_cache/cache[2][5] , \D_cache/cache[2][6] , \D_cache/cache[2][7] ,
         \D_cache/cache[2][8] , \D_cache/cache[2][9] , \D_cache/cache[2][10] ,
         \D_cache/cache[2][11] , \D_cache/cache[2][12] ,
         \D_cache/cache[2][13] , \D_cache/cache[2][14] ,
         \D_cache/cache[2][15] , \D_cache/cache[2][16] ,
         \D_cache/cache[2][17] , \D_cache/cache[2][18] ,
         \D_cache/cache[2][19] , \D_cache/cache[2][20] ,
         \D_cache/cache[2][21] , \D_cache/cache[2][22] ,
         \D_cache/cache[2][23] , \D_cache/cache[2][24] ,
         \D_cache/cache[2][25] , \D_cache/cache[2][26] ,
         \D_cache/cache[2][27] , \D_cache/cache[2][28] ,
         \D_cache/cache[2][29] , \D_cache/cache[2][30] ,
         \D_cache/cache[2][31] , \D_cache/cache[2][32] ,
         \D_cache/cache[2][33] , \D_cache/cache[2][34] ,
         \D_cache/cache[2][35] , \D_cache/cache[2][36] ,
         \D_cache/cache[2][37] , \D_cache/cache[2][38] ,
         \D_cache/cache[2][39] , \D_cache/cache[2][40] ,
         \D_cache/cache[2][41] , \D_cache/cache[2][42] ,
         \D_cache/cache[2][43] , \D_cache/cache[2][44] ,
         \D_cache/cache[2][45] , \D_cache/cache[2][46] ,
         \D_cache/cache[2][47] , \D_cache/cache[2][48] ,
         \D_cache/cache[2][49] , \D_cache/cache[2][50] ,
         \D_cache/cache[2][51] , \D_cache/cache[2][52] ,
         \D_cache/cache[2][53] , \D_cache/cache[2][54] ,
         \D_cache/cache[2][55] , \D_cache/cache[2][56] ,
         \D_cache/cache[2][57] , \D_cache/cache[2][58] ,
         \D_cache/cache[2][59] , \D_cache/cache[2][60] ,
         \D_cache/cache[2][61] , \D_cache/cache[2][62] ,
         \D_cache/cache[2][63] , \D_cache/cache[2][64] ,
         \D_cache/cache[2][65] , \D_cache/cache[2][66] ,
         \D_cache/cache[2][67] , \D_cache/cache[2][68] ,
         \D_cache/cache[2][69] , \D_cache/cache[2][70] ,
         \D_cache/cache[2][71] , \D_cache/cache[2][72] ,
         \D_cache/cache[2][73] , \D_cache/cache[2][74] ,
         \D_cache/cache[2][75] , \D_cache/cache[2][76] ,
         \D_cache/cache[2][77] , \D_cache/cache[2][78] ,
         \D_cache/cache[2][79] , \D_cache/cache[2][80] ,
         \D_cache/cache[2][81] , \D_cache/cache[2][82] ,
         \D_cache/cache[2][83] , \D_cache/cache[2][84] ,
         \D_cache/cache[2][85] , \D_cache/cache[2][86] ,
         \D_cache/cache[2][87] , \D_cache/cache[2][88] ,
         \D_cache/cache[2][89] , \D_cache/cache[2][90] ,
         \D_cache/cache[2][91] , \D_cache/cache[2][92] ,
         \D_cache/cache[2][93] , \D_cache/cache[2][94] ,
         \D_cache/cache[2][95] , \D_cache/cache[2][96] ,
         \D_cache/cache[2][97] , \D_cache/cache[2][98] ,
         \D_cache/cache[2][99] , \D_cache/cache[2][100] ,
         \D_cache/cache[2][101] , \D_cache/cache[2][102] ,
         \D_cache/cache[2][103] , \D_cache/cache[2][104] ,
         \D_cache/cache[2][105] , \D_cache/cache[2][106] ,
         \D_cache/cache[2][107] , \D_cache/cache[2][108] ,
         \D_cache/cache[2][109] , \D_cache/cache[2][110] ,
         \D_cache/cache[2][111] , \D_cache/cache[2][112] ,
         \D_cache/cache[2][113] , \D_cache/cache[2][114] ,
         \D_cache/cache[2][115] , \D_cache/cache[2][116] ,
         \D_cache/cache[2][117] , \D_cache/cache[2][118] ,
         \D_cache/cache[2][119] , \D_cache/cache[2][120] ,
         \D_cache/cache[2][121] , \D_cache/cache[2][122] ,
         \D_cache/cache[2][123] , \D_cache/cache[2][124] ,
         \D_cache/cache[2][125] , \D_cache/cache[2][126] ,
         \D_cache/cache[2][127] , \D_cache/cache[2][128] ,
         \D_cache/cache[2][129] , \D_cache/cache[2][130] ,
         \D_cache/cache[2][131] , \D_cache/cache[2][132] ,
         \D_cache/cache[2][133] , \D_cache/cache[2][134] ,
         \D_cache/cache[2][135] , \D_cache/cache[2][136] ,
         \D_cache/cache[2][137] , \D_cache/cache[2][138] ,
         \D_cache/cache[2][139] , \D_cache/cache[2][140] ,
         \D_cache/cache[2][141] , \D_cache/cache[2][142] ,
         \D_cache/cache[2][143] , \D_cache/cache[2][144] ,
         \D_cache/cache[2][145] , \D_cache/cache[2][146] ,
         \D_cache/cache[2][147] , \D_cache/cache[2][148] ,
         \D_cache/cache[2][149] , \D_cache/cache[2][150] ,
         \D_cache/cache[2][151] , \D_cache/cache[2][152] ,
         \D_cache/cache[2][153] , \D_cache/cache[2][154] ,
         \D_cache/cache[1][0] , \D_cache/cache[1][1] , \D_cache/cache[1][2] ,
         \D_cache/cache[1][3] , \D_cache/cache[1][4] , \D_cache/cache[1][5] ,
         \D_cache/cache[1][6] , \D_cache/cache[1][7] , \D_cache/cache[1][8] ,
         \D_cache/cache[1][9] , \D_cache/cache[1][10] , \D_cache/cache[1][11] ,
         \D_cache/cache[1][12] , \D_cache/cache[1][13] ,
         \D_cache/cache[1][14] , \D_cache/cache[1][15] ,
         \D_cache/cache[1][16] , \D_cache/cache[1][17] ,
         \D_cache/cache[1][18] , \D_cache/cache[1][19] ,
         \D_cache/cache[1][20] , \D_cache/cache[1][21] ,
         \D_cache/cache[1][22] , \D_cache/cache[1][23] ,
         \D_cache/cache[1][24] , \D_cache/cache[1][25] ,
         \D_cache/cache[1][26] , \D_cache/cache[1][27] ,
         \D_cache/cache[1][28] , \D_cache/cache[1][29] ,
         \D_cache/cache[1][30] , \D_cache/cache[1][31] ,
         \D_cache/cache[1][32] , \D_cache/cache[1][33] ,
         \D_cache/cache[1][34] , \D_cache/cache[1][35] ,
         \D_cache/cache[1][36] , \D_cache/cache[1][37] ,
         \D_cache/cache[1][38] , \D_cache/cache[1][39] ,
         \D_cache/cache[1][40] , \D_cache/cache[1][41] ,
         \D_cache/cache[1][42] , \D_cache/cache[1][43] ,
         \D_cache/cache[1][44] , \D_cache/cache[1][45] ,
         \D_cache/cache[1][46] , \D_cache/cache[1][47] ,
         \D_cache/cache[1][48] , \D_cache/cache[1][49] ,
         \D_cache/cache[1][50] , \D_cache/cache[1][51] ,
         \D_cache/cache[1][52] , \D_cache/cache[1][53] ,
         \D_cache/cache[1][54] , \D_cache/cache[1][55] ,
         \D_cache/cache[1][56] , \D_cache/cache[1][57] ,
         \D_cache/cache[1][58] , \D_cache/cache[1][59] ,
         \D_cache/cache[1][60] , \D_cache/cache[1][61] ,
         \D_cache/cache[1][62] , \D_cache/cache[1][63] ,
         \D_cache/cache[1][64] , \D_cache/cache[1][65] ,
         \D_cache/cache[1][66] , \D_cache/cache[1][67] ,
         \D_cache/cache[1][68] , \D_cache/cache[1][69] ,
         \D_cache/cache[1][70] , \D_cache/cache[1][71] ,
         \D_cache/cache[1][72] , \D_cache/cache[1][73] ,
         \D_cache/cache[1][74] , \D_cache/cache[1][75] ,
         \D_cache/cache[1][76] , \D_cache/cache[1][77] ,
         \D_cache/cache[1][78] , \D_cache/cache[1][79] ,
         \D_cache/cache[1][80] , \D_cache/cache[1][81] ,
         \D_cache/cache[1][82] , \D_cache/cache[1][83] ,
         \D_cache/cache[1][84] , \D_cache/cache[1][85] ,
         \D_cache/cache[1][86] , \D_cache/cache[1][87] ,
         \D_cache/cache[1][88] , \D_cache/cache[1][89] ,
         \D_cache/cache[1][90] , \D_cache/cache[1][91] ,
         \D_cache/cache[1][92] , \D_cache/cache[1][93] ,
         \D_cache/cache[1][94] , \D_cache/cache[1][95] ,
         \D_cache/cache[1][96] , \D_cache/cache[1][97] ,
         \D_cache/cache[1][98] , \D_cache/cache[1][99] ,
         \D_cache/cache[1][100] , \D_cache/cache[1][101] ,
         \D_cache/cache[1][102] , \D_cache/cache[1][103] ,
         \D_cache/cache[1][104] , \D_cache/cache[1][105] ,
         \D_cache/cache[1][106] , \D_cache/cache[1][107] ,
         \D_cache/cache[1][108] , \D_cache/cache[1][109] ,
         \D_cache/cache[1][110] , \D_cache/cache[1][111] ,
         \D_cache/cache[1][112] , \D_cache/cache[1][113] ,
         \D_cache/cache[1][114] , \D_cache/cache[1][115] ,
         \D_cache/cache[1][116] , \D_cache/cache[1][117] ,
         \D_cache/cache[1][118] , \D_cache/cache[1][119] ,
         \D_cache/cache[1][120] , \D_cache/cache[1][121] ,
         \D_cache/cache[1][122] , \D_cache/cache[1][123] ,
         \D_cache/cache[1][124] , \D_cache/cache[1][125] ,
         \D_cache/cache[1][126] , \D_cache/cache[1][127] ,
         \D_cache/cache[1][128] , \D_cache/cache[1][129] ,
         \D_cache/cache[1][130] , \D_cache/cache[1][131] ,
         \D_cache/cache[1][132] , \D_cache/cache[1][133] ,
         \D_cache/cache[1][134] , \D_cache/cache[1][135] ,
         \D_cache/cache[1][136] , \D_cache/cache[1][137] ,
         \D_cache/cache[1][138] , \D_cache/cache[1][139] ,
         \D_cache/cache[1][140] , \D_cache/cache[1][141] ,
         \D_cache/cache[1][142] , \D_cache/cache[1][143] ,
         \D_cache/cache[1][144] , \D_cache/cache[1][145] ,
         \D_cache/cache[1][146] , \D_cache/cache[1][147] ,
         \D_cache/cache[1][148] , \D_cache/cache[1][149] ,
         \D_cache/cache[1][150] , \D_cache/cache[1][151] ,
         \D_cache/cache[1][152] , \D_cache/cache[1][153] ,
         \D_cache/cache[1][154] , \D_cache/cache[0][0] , \D_cache/cache[0][1] ,
         \D_cache/cache[0][2] , \D_cache/cache[0][3] , \D_cache/cache[0][4] ,
         \D_cache/cache[0][5] , \D_cache/cache[0][6] , \D_cache/cache[0][7] ,
         \D_cache/cache[0][8] , \D_cache/cache[0][9] , \D_cache/cache[0][10] ,
         \D_cache/cache[0][11] , \D_cache/cache[0][12] ,
         \D_cache/cache[0][13] , \D_cache/cache[0][14] ,
         \D_cache/cache[0][15] , \D_cache/cache[0][16] ,
         \D_cache/cache[0][17] , \D_cache/cache[0][18] ,
         \D_cache/cache[0][19] , \D_cache/cache[0][20] ,
         \D_cache/cache[0][21] , \D_cache/cache[0][22] ,
         \D_cache/cache[0][23] , \D_cache/cache[0][24] ,
         \D_cache/cache[0][25] , \D_cache/cache[0][26] ,
         \D_cache/cache[0][27] , \D_cache/cache[0][28] ,
         \D_cache/cache[0][29] , \D_cache/cache[0][30] ,
         \D_cache/cache[0][31] , \D_cache/cache[0][32] ,
         \D_cache/cache[0][33] , \D_cache/cache[0][34] ,
         \D_cache/cache[0][35] , \D_cache/cache[0][36] ,
         \D_cache/cache[0][37] , \D_cache/cache[0][38] ,
         \D_cache/cache[0][39] , \D_cache/cache[0][40] ,
         \D_cache/cache[0][41] , \D_cache/cache[0][42] ,
         \D_cache/cache[0][43] , \D_cache/cache[0][44] ,
         \D_cache/cache[0][45] , \D_cache/cache[0][46] ,
         \D_cache/cache[0][47] , \D_cache/cache[0][48] ,
         \D_cache/cache[0][49] , \D_cache/cache[0][50] ,
         \D_cache/cache[0][51] , \D_cache/cache[0][52] ,
         \D_cache/cache[0][53] , \D_cache/cache[0][54] ,
         \D_cache/cache[0][55] , \D_cache/cache[0][56] ,
         \D_cache/cache[0][57] , \D_cache/cache[0][58] ,
         \D_cache/cache[0][59] , \D_cache/cache[0][60] ,
         \D_cache/cache[0][61] , \D_cache/cache[0][62] ,
         \D_cache/cache[0][63] , \D_cache/cache[0][64] ,
         \D_cache/cache[0][65] , \D_cache/cache[0][66] ,
         \D_cache/cache[0][67] , \D_cache/cache[0][68] ,
         \D_cache/cache[0][69] , \D_cache/cache[0][70] ,
         \D_cache/cache[0][71] , \D_cache/cache[0][72] ,
         \D_cache/cache[0][73] , \D_cache/cache[0][74] ,
         \D_cache/cache[0][75] , \D_cache/cache[0][76] ,
         \D_cache/cache[0][77] , \D_cache/cache[0][78] ,
         \D_cache/cache[0][79] , \D_cache/cache[0][80] ,
         \D_cache/cache[0][81] , \D_cache/cache[0][82] ,
         \D_cache/cache[0][83] , \D_cache/cache[0][84] ,
         \D_cache/cache[0][85] , \D_cache/cache[0][86] ,
         \D_cache/cache[0][87] , \D_cache/cache[0][88] ,
         \D_cache/cache[0][89] , \D_cache/cache[0][90] ,
         \D_cache/cache[0][91] , \D_cache/cache[0][92] ,
         \D_cache/cache[0][93] , \D_cache/cache[0][94] ,
         \D_cache/cache[0][95] , \D_cache/cache[0][96] ,
         \D_cache/cache[0][97] , \D_cache/cache[0][98] ,
         \D_cache/cache[0][99] , \D_cache/cache[0][100] ,
         \D_cache/cache[0][101] , \D_cache/cache[0][102] ,
         \D_cache/cache[0][103] , \D_cache/cache[0][104] ,
         \D_cache/cache[0][105] , \D_cache/cache[0][106] ,
         \D_cache/cache[0][107] , \D_cache/cache[0][108] ,
         \D_cache/cache[0][109] , \D_cache/cache[0][110] ,
         \D_cache/cache[0][111] , \D_cache/cache[0][112] ,
         \D_cache/cache[0][113] , \D_cache/cache[0][114] ,
         \D_cache/cache[0][115] , \D_cache/cache[0][116] ,
         \D_cache/cache[0][117] , \D_cache/cache[0][118] ,
         \D_cache/cache[0][119] , \D_cache/cache[0][120] ,
         \D_cache/cache[0][121] , \D_cache/cache[0][122] ,
         \D_cache/cache[0][123] , \D_cache/cache[0][124] ,
         \D_cache/cache[0][125] , \D_cache/cache[0][126] ,
         \D_cache/cache[0][127] , \D_cache/cache[0][128] ,
         \D_cache/cache[0][129] , \D_cache/cache[0][130] ,
         \D_cache/cache[0][131] , \D_cache/cache[0][132] ,
         \D_cache/cache[0][133] , \D_cache/cache[0][134] ,
         \D_cache/cache[0][135] , \D_cache/cache[0][136] ,
         \D_cache/cache[0][137] , \D_cache/cache[0][138] ,
         \D_cache/cache[0][139] , \D_cache/cache[0][140] ,
         \D_cache/cache[0][141] , \D_cache/cache[0][142] ,
         \D_cache/cache[0][143] , \D_cache/cache[0][144] ,
         \D_cache/cache[0][145] , \D_cache/cache[0][146] ,
         \D_cache/cache[0][147] , \D_cache/cache[0][148] ,
         \D_cache/cache[0][149] , \D_cache/cache[0][150] ,
         \D_cache/cache[0][151] , \D_cache/cache[0][152] ,
         \D_cache/cache[0][153] , \D_cache/cache[0][154] , \i_MIPS/PHT_2/n54 ,
         \i_MIPS/PHT_2/n53 , \i_MIPS/PHT_2/n52 , \i_MIPS/PHT_2/n50 ,
         \i_MIPS/PHT_2/n48 , \i_MIPS/PHT_2/n47 , \i_MIPS/PHT_2/n46 ,
         \i_MIPS/PHT_2/n45 , \i_MIPS/PHT_2/n44 , \i_MIPS/PHT_2/n13 ,
         \i_MIPS/PHT_2/n12 , \i_MIPS/PHT_2/n8 , \i_MIPS/PHT_2/n7 ,
         \i_MIPS/PHT_2/n6 , \i_MIPS/PHT_2/n5 , \i_MIPS/PHT_2/n4 ,
         \i_MIPS/PHT_2/n3 , \i_MIPS/PHT_2/n2 , \i_MIPS/PHT_2/counter ,
         \i_MIPS/PHT_2/history_state[1] , \i_MIPS/PHT_2/history_state[0] ,
         \i_MIPS/PHT_2/current_state_3[0] , \i_MIPS/PHT_2/current_state_2[1] ,
         \i_MIPS/PHT_2/current_state_2[0] , \i_MIPS/PHT_2/current_state_1[1] ,
         \i_MIPS/PHT_2/current_state_0[1] , \i_MIPS/PC/n65 , \i_MIPS/PC/n64 ,
         \i_MIPS/PC/n63 , \i_MIPS/PC/n62 , \i_MIPS/PC/n61 , \i_MIPS/PC/n60 ,
         \i_MIPS/PC/n59 , \i_MIPS/PC/n58 , \i_MIPS/PC/n57 , \i_MIPS/PC/n56 ,
         \i_MIPS/PC/n55 , \i_MIPS/PC/n54 , \i_MIPS/PC/n53 , \i_MIPS/PC/n52 ,
         \i_MIPS/PC/n51 , \i_MIPS/PC/n50 , \i_MIPS/PC/n49 , \i_MIPS/PC/n48 ,
         \i_MIPS/PC/n47 , \i_MIPS/PC/n46 , \i_MIPS/PC/n45 , \i_MIPS/PC/n44 ,
         \i_MIPS/PC/n43 , \i_MIPS/PC/n42 , \i_MIPS/PC/n41 , \i_MIPS/PC/n40 ,
         \i_MIPS/PC/n39 , \i_MIPS/PC/n38 , \i_MIPS/PC/n37 , \i_MIPS/PC/n36 ,
         \i_MIPS/PC/n35 , \i_MIPS/PC/n34 , \i_MIPS/PC/n33 , \i_MIPS/PC/n32 ,
         \i_MIPS/PC/n31 , \i_MIPS/PC/n30 , \i_MIPS/PC/n29 , \i_MIPS/PC/n28 ,
         \i_MIPS/PC/n27 , \i_MIPS/PC/n26 , \i_MIPS/PC/n25 , \i_MIPS/PC/n24 ,
         \i_MIPS/PC/n23 , \i_MIPS/PC/n22 , \i_MIPS/PC/n21 , \i_MIPS/PC/n20 ,
         \i_MIPS/PC/n19 , \i_MIPS/PC/n18 , \i_MIPS/PC/n17 , \i_MIPS/PC/n16 ,
         \i_MIPS/PC/n15 , \i_MIPS/PC/n14 , \i_MIPS/PC/n13 , \i_MIPS/PC/n12 ,
         \i_MIPS/PC/n11 , \i_MIPS/PC/n9 , \i_MIPS/PC/n7 , \i_MIPS/PC/n5 ,
         \i_MIPS/PC/n3 , \i_MIPS/PC/n2 , \i_MIPS/Register/n1139 ,
         \i_MIPS/Register/n1138 , \i_MIPS/Register/n1137 ,
         \i_MIPS/Register/n1136 , \i_MIPS/Register/n1135 ,
         \i_MIPS/Register/n1134 , \i_MIPS/Register/n1133 ,
         \i_MIPS/Register/n1132 , \i_MIPS/Register/n1131 ,
         \i_MIPS/Register/n1130 , \i_MIPS/Register/n1129 ,
         \i_MIPS/Register/n1128 , \i_MIPS/Register/n1127 ,
         \i_MIPS/Register/n1126 , \i_MIPS/Register/n1125 ,
         \i_MIPS/Register/n1124 , \i_MIPS/Register/n1123 ,
         \i_MIPS/Register/n1122 , \i_MIPS/Register/n1121 ,
         \i_MIPS/Register/n1120 , \i_MIPS/Register/n1119 ,
         \i_MIPS/Register/n1118 , \i_MIPS/Register/n1117 ,
         \i_MIPS/Register/n1116 , \i_MIPS/Register/n1115 ,
         \i_MIPS/Register/n1114 , \i_MIPS/Register/n1113 ,
         \i_MIPS/Register/n1112 , \i_MIPS/Register/n1111 ,
         \i_MIPS/Register/n1110 , \i_MIPS/Register/n1109 ,
         \i_MIPS/Register/n1108 , \i_MIPS/Register/n1107 ,
         \i_MIPS/Register/n1106 , \i_MIPS/Register/n1105 ,
         \i_MIPS/Register/n1104 , \i_MIPS/Register/n1103 ,
         \i_MIPS/Register/n1102 , \i_MIPS/Register/n1101 ,
         \i_MIPS/Register/n1100 , \i_MIPS/Register/n1099 ,
         \i_MIPS/Register/n1098 , \i_MIPS/Register/n1097 ,
         \i_MIPS/Register/n1096 , \i_MIPS/Register/n1095 ,
         \i_MIPS/Register/n1094 , \i_MIPS/Register/n1093 ,
         \i_MIPS/Register/n1092 , \i_MIPS/Register/n1091 ,
         \i_MIPS/Register/n1090 , \i_MIPS/Register/n1089 ,
         \i_MIPS/Register/n1088 , \i_MIPS/Register/n1087 ,
         \i_MIPS/Register/n1086 , \i_MIPS/Register/n1085 ,
         \i_MIPS/Register/n1084 , \i_MIPS/Register/n1083 ,
         \i_MIPS/Register/n1082 , \i_MIPS/Register/n1081 ,
         \i_MIPS/Register/n1080 , \i_MIPS/Register/n1079 ,
         \i_MIPS/Register/n1078 , \i_MIPS/Register/n1077 ,
         \i_MIPS/Register/n1076 , \i_MIPS/Register/n1075 ,
         \i_MIPS/Register/n1074 , \i_MIPS/Register/n1073 ,
         \i_MIPS/Register/n1072 , \i_MIPS/Register/n1071 ,
         \i_MIPS/Register/n1070 , \i_MIPS/Register/n1069 ,
         \i_MIPS/Register/n1068 , \i_MIPS/Register/n1067 ,
         \i_MIPS/Register/n1066 , \i_MIPS/Register/n1065 ,
         \i_MIPS/Register/n1064 , \i_MIPS/Register/n1063 ,
         \i_MIPS/Register/n1062 , \i_MIPS/Register/n1061 ,
         \i_MIPS/Register/n1060 , \i_MIPS/Register/n1059 ,
         \i_MIPS/Register/n1058 , \i_MIPS/Register/n1057 ,
         \i_MIPS/Register/n1056 , \i_MIPS/Register/n1055 ,
         \i_MIPS/Register/n1054 , \i_MIPS/Register/n1053 ,
         \i_MIPS/Register/n1052 , \i_MIPS/Register/n1051 ,
         \i_MIPS/Register/n1050 , \i_MIPS/Register/n1049 ,
         \i_MIPS/Register/n1048 , \i_MIPS/Register/n1047 ,
         \i_MIPS/Register/n1046 , \i_MIPS/Register/n1045 ,
         \i_MIPS/Register/n1044 , \i_MIPS/Register/n1043 ,
         \i_MIPS/Register/n1042 , \i_MIPS/Register/n1041 ,
         \i_MIPS/Register/n1040 , \i_MIPS/Register/n1039 ,
         \i_MIPS/Register/n1038 , \i_MIPS/Register/n1037 ,
         \i_MIPS/Register/n1036 , \i_MIPS/Register/n1035 ,
         \i_MIPS/Register/n1034 , \i_MIPS/Register/n1033 ,
         \i_MIPS/Register/n1032 , \i_MIPS/Register/n1031 ,
         \i_MIPS/Register/n1030 , \i_MIPS/Register/n1029 ,
         \i_MIPS/Register/n1028 , \i_MIPS/Register/n1027 ,
         \i_MIPS/Register/n1026 , \i_MIPS/Register/n1025 ,
         \i_MIPS/Register/n1024 , \i_MIPS/Register/n1023 ,
         \i_MIPS/Register/n1022 , \i_MIPS/Register/n1021 ,
         \i_MIPS/Register/n1020 , \i_MIPS/Register/n1019 ,
         \i_MIPS/Register/n1018 , \i_MIPS/Register/n1017 ,
         \i_MIPS/Register/n1016 , \i_MIPS/Register/n1015 ,
         \i_MIPS/Register/n1014 , \i_MIPS/Register/n1013 ,
         \i_MIPS/Register/n1012 , \i_MIPS/Register/n1011 ,
         \i_MIPS/Register/n1010 , \i_MIPS/Register/n1009 ,
         \i_MIPS/Register/n1008 , \i_MIPS/Register/n1007 ,
         \i_MIPS/Register/n1006 , \i_MIPS/Register/n1005 ,
         \i_MIPS/Register/n1004 , \i_MIPS/Register/n1003 ,
         \i_MIPS/Register/n1002 , \i_MIPS/Register/n1001 ,
         \i_MIPS/Register/n1000 , \i_MIPS/Register/n999 ,
         \i_MIPS/Register/n998 , \i_MIPS/Register/n997 ,
         \i_MIPS/Register/n996 , \i_MIPS/Register/n995 ,
         \i_MIPS/Register/n994 , \i_MIPS/Register/n993 ,
         \i_MIPS/Register/n992 , \i_MIPS/Register/n991 ,
         \i_MIPS/Register/n990 , \i_MIPS/Register/n989 ,
         \i_MIPS/Register/n988 , \i_MIPS/Register/n987 ,
         \i_MIPS/Register/n986 , \i_MIPS/Register/n985 ,
         \i_MIPS/Register/n984 , \i_MIPS/Register/n983 ,
         \i_MIPS/Register/n982 , \i_MIPS/Register/n981 ,
         \i_MIPS/Register/n980 , \i_MIPS/Register/n979 ,
         \i_MIPS/Register/n978 , \i_MIPS/Register/n977 ,
         \i_MIPS/Register/n976 , \i_MIPS/Register/n975 ,
         \i_MIPS/Register/n974 , \i_MIPS/Register/n973 ,
         \i_MIPS/Register/n972 , \i_MIPS/Register/n971 ,
         \i_MIPS/Register/n970 , \i_MIPS/Register/n969 ,
         \i_MIPS/Register/n968 , \i_MIPS/Register/n967 ,
         \i_MIPS/Register/n966 , \i_MIPS/Register/n965 ,
         \i_MIPS/Register/n964 , \i_MIPS/Register/n963 ,
         \i_MIPS/Register/n962 , \i_MIPS/Register/n961 ,
         \i_MIPS/Register/n960 , \i_MIPS/Register/n959 ,
         \i_MIPS/Register/n958 , \i_MIPS/Register/n957 ,
         \i_MIPS/Register/n956 , \i_MIPS/Register/n955 ,
         \i_MIPS/Register/n954 , \i_MIPS/Register/n953 ,
         \i_MIPS/Register/n952 , \i_MIPS/Register/n951 ,
         \i_MIPS/Register/n950 , \i_MIPS/Register/n949 ,
         \i_MIPS/Register/n948 , \i_MIPS/Register/n947 ,
         \i_MIPS/Register/n946 , \i_MIPS/Register/n945 ,
         \i_MIPS/Register/n944 , \i_MIPS/Register/n943 ,
         \i_MIPS/Register/n942 , \i_MIPS/Register/n941 ,
         \i_MIPS/Register/n940 , \i_MIPS/Register/n939 ,
         \i_MIPS/Register/n938 , \i_MIPS/Register/n937 ,
         \i_MIPS/Register/n936 , \i_MIPS/Register/n935 ,
         \i_MIPS/Register/n934 , \i_MIPS/Register/n933 ,
         \i_MIPS/Register/n932 , \i_MIPS/Register/n931 ,
         \i_MIPS/Register/n930 , \i_MIPS/Register/n929 ,
         \i_MIPS/Register/n928 , \i_MIPS/Register/n927 ,
         \i_MIPS/Register/n926 , \i_MIPS/Register/n925 ,
         \i_MIPS/Register/n924 , \i_MIPS/Register/n923 ,
         \i_MIPS/Register/n922 , \i_MIPS/Register/n921 ,
         \i_MIPS/Register/n920 , \i_MIPS/Register/n919 ,
         \i_MIPS/Register/n918 , \i_MIPS/Register/n917 ,
         \i_MIPS/Register/n916 , \i_MIPS/Register/n915 ,
         \i_MIPS/Register/n914 , \i_MIPS/Register/n913 ,
         \i_MIPS/Register/n912 , \i_MIPS/Register/n911 ,
         \i_MIPS/Register/n910 , \i_MIPS/Register/n909 ,
         \i_MIPS/Register/n908 , \i_MIPS/Register/n907 ,
         \i_MIPS/Register/n906 , \i_MIPS/Register/n905 ,
         \i_MIPS/Register/n904 , \i_MIPS/Register/n903 ,
         \i_MIPS/Register/n902 , \i_MIPS/Register/n901 ,
         \i_MIPS/Register/n900 , \i_MIPS/Register/n899 ,
         \i_MIPS/Register/n898 , \i_MIPS/Register/n897 ,
         \i_MIPS/Register/n896 , \i_MIPS/Register/n895 ,
         \i_MIPS/Register/n894 , \i_MIPS/Register/n893 ,
         \i_MIPS/Register/n892 , \i_MIPS/Register/n891 ,
         \i_MIPS/Register/n890 , \i_MIPS/Register/n889 ,
         \i_MIPS/Register/n888 , \i_MIPS/Register/n887 ,
         \i_MIPS/Register/n886 , \i_MIPS/Register/n885 ,
         \i_MIPS/Register/n884 , \i_MIPS/Register/n883 ,
         \i_MIPS/Register/n882 , \i_MIPS/Register/n881 ,
         \i_MIPS/Register/n880 , \i_MIPS/Register/n879 ,
         \i_MIPS/Register/n878 , \i_MIPS/Register/n877 ,
         \i_MIPS/Register/n876 , \i_MIPS/Register/n875 ,
         \i_MIPS/Register/n874 , \i_MIPS/Register/n873 ,
         \i_MIPS/Register/n872 , \i_MIPS/Register/n871 ,
         \i_MIPS/Register/n870 , \i_MIPS/Register/n869 ,
         \i_MIPS/Register/n868 , \i_MIPS/Register/n867 ,
         \i_MIPS/Register/n866 , \i_MIPS/Register/n865 ,
         \i_MIPS/Register/n864 , \i_MIPS/Register/n863 ,
         \i_MIPS/Register/n862 , \i_MIPS/Register/n861 ,
         \i_MIPS/Register/n860 , \i_MIPS/Register/n859 ,
         \i_MIPS/Register/n858 , \i_MIPS/Register/n857 ,
         \i_MIPS/Register/n856 , \i_MIPS/Register/n855 ,
         \i_MIPS/Register/n854 , \i_MIPS/Register/n853 ,
         \i_MIPS/Register/n852 , \i_MIPS/Register/n851 ,
         \i_MIPS/Register/n850 , \i_MIPS/Register/n849 ,
         \i_MIPS/Register/n848 , \i_MIPS/Register/n847 ,
         \i_MIPS/Register/n846 , \i_MIPS/Register/n845 ,
         \i_MIPS/Register/n844 , \i_MIPS/Register/n843 ,
         \i_MIPS/Register/n842 , \i_MIPS/Register/n841 ,
         \i_MIPS/Register/n840 , \i_MIPS/Register/n839 ,
         \i_MIPS/Register/n838 , \i_MIPS/Register/n837 ,
         \i_MIPS/Register/n836 , \i_MIPS/Register/n835 ,
         \i_MIPS/Register/n834 , \i_MIPS/Register/n833 ,
         \i_MIPS/Register/n832 , \i_MIPS/Register/n831 ,
         \i_MIPS/Register/n830 , \i_MIPS/Register/n829 ,
         \i_MIPS/Register/n828 , \i_MIPS/Register/n827 ,
         \i_MIPS/Register/n826 , \i_MIPS/Register/n825 ,
         \i_MIPS/Register/n824 , \i_MIPS/Register/n823 ,
         \i_MIPS/Register/n822 , \i_MIPS/Register/n821 ,
         \i_MIPS/Register/n820 , \i_MIPS/Register/n819 ,
         \i_MIPS/Register/n818 , \i_MIPS/Register/n817 ,
         \i_MIPS/Register/n816 , \i_MIPS/Register/n815 ,
         \i_MIPS/Register/n814 , \i_MIPS/Register/n813 ,
         \i_MIPS/Register/n812 , \i_MIPS/Register/n811 ,
         \i_MIPS/Register/n810 , \i_MIPS/Register/n809 ,
         \i_MIPS/Register/n808 , \i_MIPS/Register/n807 ,
         \i_MIPS/Register/n806 , \i_MIPS/Register/n805 ,
         \i_MIPS/Register/n804 , \i_MIPS/Register/n803 ,
         \i_MIPS/Register/n802 , \i_MIPS/Register/n801 ,
         \i_MIPS/Register/n800 , \i_MIPS/Register/n799 ,
         \i_MIPS/Register/n798 , \i_MIPS/Register/n797 ,
         \i_MIPS/Register/n796 , \i_MIPS/Register/n795 ,
         \i_MIPS/Register/n794 , \i_MIPS/Register/n793 ,
         \i_MIPS/Register/n792 , \i_MIPS/Register/n791 ,
         \i_MIPS/Register/n790 , \i_MIPS/Register/n789 ,
         \i_MIPS/Register/n788 , \i_MIPS/Register/n787 ,
         \i_MIPS/Register/n786 , \i_MIPS/Register/n785 ,
         \i_MIPS/Register/n784 , \i_MIPS/Register/n783 ,
         \i_MIPS/Register/n782 , \i_MIPS/Register/n781 ,
         \i_MIPS/Register/n780 , \i_MIPS/Register/n779 ,
         \i_MIPS/Register/n778 , \i_MIPS/Register/n777 ,
         \i_MIPS/Register/n776 , \i_MIPS/Register/n775 ,
         \i_MIPS/Register/n774 , \i_MIPS/Register/n773 ,
         \i_MIPS/Register/n772 , \i_MIPS/Register/n771 ,
         \i_MIPS/Register/n770 , \i_MIPS/Register/n769 ,
         \i_MIPS/Register/n768 , \i_MIPS/Register/n767 ,
         \i_MIPS/Register/n766 , \i_MIPS/Register/n765 ,
         \i_MIPS/Register/n764 , \i_MIPS/Register/n763 ,
         \i_MIPS/Register/n762 , \i_MIPS/Register/n761 ,
         \i_MIPS/Register/n760 , \i_MIPS/Register/n759 ,
         \i_MIPS/Register/n758 , \i_MIPS/Register/n757 ,
         \i_MIPS/Register/n756 , \i_MIPS/Register/n755 ,
         \i_MIPS/Register/n754 , \i_MIPS/Register/n753 ,
         \i_MIPS/Register/n752 , \i_MIPS/Register/n751 ,
         \i_MIPS/Register/n750 , \i_MIPS/Register/n749 ,
         \i_MIPS/Register/n748 , \i_MIPS/Register/n747 ,
         \i_MIPS/Register/n746 , \i_MIPS/Register/n745 ,
         \i_MIPS/Register/n744 , \i_MIPS/Register/n743 ,
         \i_MIPS/Register/n742 , \i_MIPS/Register/n741 ,
         \i_MIPS/Register/n740 , \i_MIPS/Register/n739 ,
         \i_MIPS/Register/n738 , \i_MIPS/Register/n737 ,
         \i_MIPS/Register/n736 , \i_MIPS/Register/n735 ,
         \i_MIPS/Register/n734 , \i_MIPS/Register/n733 ,
         \i_MIPS/Register/n732 , \i_MIPS/Register/n731 ,
         \i_MIPS/Register/n730 , \i_MIPS/Register/n729 ,
         \i_MIPS/Register/n728 , \i_MIPS/Register/n727 ,
         \i_MIPS/Register/n726 , \i_MIPS/Register/n725 ,
         \i_MIPS/Register/n724 , \i_MIPS/Register/n723 ,
         \i_MIPS/Register/n722 , \i_MIPS/Register/n721 ,
         \i_MIPS/Register/n720 , \i_MIPS/Register/n719 ,
         \i_MIPS/Register/n718 , \i_MIPS/Register/n717 ,
         \i_MIPS/Register/n716 , \i_MIPS/Register/n715 ,
         \i_MIPS/Register/n714 , \i_MIPS/Register/n713 ,
         \i_MIPS/Register/n712 , \i_MIPS/Register/n711 ,
         \i_MIPS/Register/n710 , \i_MIPS/Register/n709 ,
         \i_MIPS/Register/n708 , \i_MIPS/Register/n707 ,
         \i_MIPS/Register/n706 , \i_MIPS/Register/n705 ,
         \i_MIPS/Register/n704 , \i_MIPS/Register/n703 ,
         \i_MIPS/Register/n702 , \i_MIPS/Register/n701 ,
         \i_MIPS/Register/n700 , \i_MIPS/Register/n699 ,
         \i_MIPS/Register/n698 , \i_MIPS/Register/n697 ,
         \i_MIPS/Register/n696 , \i_MIPS/Register/n695 ,
         \i_MIPS/Register/n694 , \i_MIPS/Register/n693 ,
         \i_MIPS/Register/n692 , \i_MIPS/Register/n691 ,
         \i_MIPS/Register/n690 , \i_MIPS/Register/n689 ,
         \i_MIPS/Register/n688 , \i_MIPS/Register/n687 ,
         \i_MIPS/Register/n686 , \i_MIPS/Register/n685 ,
         \i_MIPS/Register/n684 , \i_MIPS/Register/n683 ,
         \i_MIPS/Register/n682 , \i_MIPS/Register/n681 ,
         \i_MIPS/Register/n680 , \i_MIPS/Register/n679 ,
         \i_MIPS/Register/n678 , \i_MIPS/Register/n677 ,
         \i_MIPS/Register/n676 , \i_MIPS/Register/n675 ,
         \i_MIPS/Register/n674 , \i_MIPS/Register/n673 ,
         \i_MIPS/Register/n672 , \i_MIPS/Register/n671 ,
         \i_MIPS/Register/n670 , \i_MIPS/Register/n669 ,
         \i_MIPS/Register/n668 , \i_MIPS/Register/n667 ,
         \i_MIPS/Register/n666 , \i_MIPS/Register/n665 ,
         \i_MIPS/Register/n664 , \i_MIPS/Register/n663 ,
         \i_MIPS/Register/n662 , \i_MIPS/Register/n661 ,
         \i_MIPS/Register/n660 , \i_MIPS/Register/n659 ,
         \i_MIPS/Register/n658 , \i_MIPS/Register/n657 ,
         \i_MIPS/Register/n656 , \i_MIPS/Register/n655 ,
         \i_MIPS/Register/n654 , \i_MIPS/Register/n653 ,
         \i_MIPS/Register/n652 , \i_MIPS/Register/n651 ,
         \i_MIPS/Register/n650 , \i_MIPS/Register/n649 ,
         \i_MIPS/Register/n648 , \i_MIPS/Register/n647 ,
         \i_MIPS/Register/n646 , \i_MIPS/Register/n645 ,
         \i_MIPS/Register/n644 , \i_MIPS/Register/n643 ,
         \i_MIPS/Register/n642 , \i_MIPS/Register/n641 ,
         \i_MIPS/Register/n640 , \i_MIPS/Register/n639 ,
         \i_MIPS/Register/n638 , \i_MIPS/Register/n637 ,
         \i_MIPS/Register/n636 , \i_MIPS/Register/n635 ,
         \i_MIPS/Register/n634 , \i_MIPS/Register/n633 ,
         \i_MIPS/Register/n632 , \i_MIPS/Register/n631 ,
         \i_MIPS/Register/n630 , \i_MIPS/Register/n629 ,
         \i_MIPS/Register/n628 , \i_MIPS/Register/n627 ,
         \i_MIPS/Register/n626 , \i_MIPS/Register/n625 ,
         \i_MIPS/Register/n624 , \i_MIPS/Register/n623 ,
         \i_MIPS/Register/n622 , \i_MIPS/Register/n621 ,
         \i_MIPS/Register/n620 , \i_MIPS/Register/n619 ,
         \i_MIPS/Register/n618 , \i_MIPS/Register/n617 ,
         \i_MIPS/Register/n616 , \i_MIPS/Register/n615 ,
         \i_MIPS/Register/n614 , \i_MIPS/Register/n613 ,
         \i_MIPS/Register/n612 , \i_MIPS/Register/n611 ,
         \i_MIPS/Register/n610 , \i_MIPS/Register/n609 ,
         \i_MIPS/Register/n608 , \i_MIPS/Register/n607 ,
         \i_MIPS/Register/n606 , \i_MIPS/Register/n605 ,
         \i_MIPS/Register/n604 , \i_MIPS/Register/n603 ,
         \i_MIPS/Register/n602 , \i_MIPS/Register/n601 ,
         \i_MIPS/Register/n600 , \i_MIPS/Register/n599 ,
         \i_MIPS/Register/n598 , \i_MIPS/Register/n597 ,
         \i_MIPS/Register/n596 , \i_MIPS/Register/n595 ,
         \i_MIPS/Register/n594 , \i_MIPS/Register/n593 ,
         \i_MIPS/Register/n592 , \i_MIPS/Register/n591 ,
         \i_MIPS/Register/n590 , \i_MIPS/Register/n589 ,
         \i_MIPS/Register/n588 , \i_MIPS/Register/n587 ,
         \i_MIPS/Register/n586 , \i_MIPS/Register/n585 ,
         \i_MIPS/Register/n584 , \i_MIPS/Register/n583 ,
         \i_MIPS/Register/n582 , \i_MIPS/Register/n581 ,
         \i_MIPS/Register/n580 , \i_MIPS/Register/n579 ,
         \i_MIPS/Register/n578 , \i_MIPS/Register/n577 ,
         \i_MIPS/Register/n576 , \i_MIPS/Register/n575 ,
         \i_MIPS/Register/n574 , \i_MIPS/Register/n573 ,
         \i_MIPS/Register/n572 , \i_MIPS/Register/n571 ,
         \i_MIPS/Register/n570 , \i_MIPS/Register/n569 ,
         \i_MIPS/Register/n568 , \i_MIPS/Register/n567 ,
         \i_MIPS/Register/n566 , \i_MIPS/Register/n565 ,
         \i_MIPS/Register/n564 , \i_MIPS/Register/n563 ,
         \i_MIPS/Register/n562 , \i_MIPS/Register/n561 ,
         \i_MIPS/Register/n560 , \i_MIPS/Register/n559 ,
         \i_MIPS/Register/n558 , \i_MIPS/Register/n557 ,
         \i_MIPS/Register/n556 , \i_MIPS/Register/n555 ,
         \i_MIPS/Register/n554 , \i_MIPS/Register/n553 ,
         \i_MIPS/Register/n552 , \i_MIPS/Register/n551 ,
         \i_MIPS/Register/n550 , \i_MIPS/Register/n549 ,
         \i_MIPS/Register/n548 , \i_MIPS/Register/n547 ,
         \i_MIPS/Register/n546 , \i_MIPS/Register/n545 ,
         \i_MIPS/Register/n544 , \i_MIPS/Register/n543 ,
         \i_MIPS/Register/n542 , \i_MIPS/Register/n541 ,
         \i_MIPS/Register/n540 , \i_MIPS/Register/n539 ,
         \i_MIPS/Register/n538 , \i_MIPS/Register/n537 ,
         \i_MIPS/Register/n536 , \i_MIPS/Register/n535 ,
         \i_MIPS/Register/n534 , \i_MIPS/Register/n533 ,
         \i_MIPS/Register/n532 , \i_MIPS/Register/n531 ,
         \i_MIPS/Register/n530 , \i_MIPS/Register/n529 ,
         \i_MIPS/Register/n528 , \i_MIPS/Register/n527 ,
         \i_MIPS/Register/n526 , \i_MIPS/Register/n525 ,
         \i_MIPS/Register/n524 , \i_MIPS/Register/n523 ,
         \i_MIPS/Register/n522 , \i_MIPS/Register/n521 ,
         \i_MIPS/Register/n520 , \i_MIPS/Register/n519 ,
         \i_MIPS/Register/n518 , \i_MIPS/Register/n517 ,
         \i_MIPS/Register/n516 , \i_MIPS/Register/n515 ,
         \i_MIPS/Register/n514 , \i_MIPS/Register/n513 ,
         \i_MIPS/Register/n512 , \i_MIPS/Register/n511 ,
         \i_MIPS/Register/n510 , \i_MIPS/Register/n509 ,
         \i_MIPS/Register/n508 , \i_MIPS/Register/n507 ,
         \i_MIPS/Register/n506 , \i_MIPS/Register/n505 ,
         \i_MIPS/Register/n504 , \i_MIPS/Register/n503 ,
         \i_MIPS/Register/n502 , \i_MIPS/Register/n501 ,
         \i_MIPS/Register/n500 , \i_MIPS/Register/n499 ,
         \i_MIPS/Register/n498 , \i_MIPS/Register/n497 ,
         \i_MIPS/Register/n496 , \i_MIPS/Register/n495 ,
         \i_MIPS/Register/n494 , \i_MIPS/Register/n493 ,
         \i_MIPS/Register/n492 , \i_MIPS/Register/n491 ,
         \i_MIPS/Register/n490 , \i_MIPS/Register/n489 ,
         \i_MIPS/Register/n488 , \i_MIPS/Register/n487 ,
         \i_MIPS/Register/n486 , \i_MIPS/Register/n485 ,
         \i_MIPS/Register/n484 , \i_MIPS/Register/n483 ,
         \i_MIPS/Register/n482 , \i_MIPS/Register/n481 ,
         \i_MIPS/Register/n480 , \i_MIPS/Register/n479 ,
         \i_MIPS/Register/n478 , \i_MIPS/Register/n477 ,
         \i_MIPS/Register/n476 , \i_MIPS/Register/n475 ,
         \i_MIPS/Register/n474 , \i_MIPS/Register/n473 ,
         \i_MIPS/Register/n472 , \i_MIPS/Register/n471 ,
         \i_MIPS/Register/n470 , \i_MIPS/Register/n469 ,
         \i_MIPS/Register/n468 , \i_MIPS/Register/n467 ,
         \i_MIPS/Register/n466 , \i_MIPS/Register/n465 ,
         \i_MIPS/Register/n464 , \i_MIPS/Register/n463 ,
         \i_MIPS/Register/n462 , \i_MIPS/Register/n461 ,
         \i_MIPS/Register/n460 , \i_MIPS/Register/n459 ,
         \i_MIPS/Register/n458 , \i_MIPS/Register/n457 ,
         \i_MIPS/Register/n456 , \i_MIPS/Register/n455 ,
         \i_MIPS/Register/n454 , \i_MIPS/Register/n453 ,
         \i_MIPS/Register/n452 , \i_MIPS/Register/n451 ,
         \i_MIPS/Register/n450 , \i_MIPS/Register/n449 ,
         \i_MIPS/Register/n448 , \i_MIPS/Register/n447 ,
         \i_MIPS/Register/n446 , \i_MIPS/Register/n445 ,
         \i_MIPS/Register/n444 , \i_MIPS/Register/n443 ,
         \i_MIPS/Register/n442 , \i_MIPS/Register/n441 ,
         \i_MIPS/Register/n440 , \i_MIPS/Register/n439 ,
         \i_MIPS/Register/n438 , \i_MIPS/Register/n437 ,
         \i_MIPS/Register/n436 , \i_MIPS/Register/n435 ,
         \i_MIPS/Register/n434 , \i_MIPS/Register/n433 ,
         \i_MIPS/Register/n432 , \i_MIPS/Register/n431 ,
         \i_MIPS/Register/n430 , \i_MIPS/Register/n429 ,
         \i_MIPS/Register/n428 , \i_MIPS/Register/n427 ,
         \i_MIPS/Register/n426 , \i_MIPS/Register/n425 ,
         \i_MIPS/Register/n424 , \i_MIPS/Register/n423 ,
         \i_MIPS/Register/n422 , \i_MIPS/Register/n421 ,
         \i_MIPS/Register/n420 , \i_MIPS/Register/n419 ,
         \i_MIPS/Register/n418 , \i_MIPS/Register/n417 ,
         \i_MIPS/Register/n416 , \i_MIPS/Register/n415 ,
         \i_MIPS/Register/n414 , \i_MIPS/Register/n413 ,
         \i_MIPS/Register/n412 , \i_MIPS/Register/n411 ,
         \i_MIPS/Register/n410 , \i_MIPS/Register/n409 ,
         \i_MIPS/Register/n408 , \i_MIPS/Register/n407 ,
         \i_MIPS/Register/n406 , \i_MIPS/Register/n405 ,
         \i_MIPS/Register/n404 , \i_MIPS/Register/n403 ,
         \i_MIPS/Register/n402 , \i_MIPS/Register/n401 ,
         \i_MIPS/Register/n400 , \i_MIPS/Register/n399 ,
         \i_MIPS/Register/n398 , \i_MIPS/Register/n397 ,
         \i_MIPS/Register/n396 , \i_MIPS/Register/n395 ,
         \i_MIPS/Register/n394 , \i_MIPS/Register/n393 ,
         \i_MIPS/Register/n392 , \i_MIPS/Register/n391 ,
         \i_MIPS/Register/n390 , \i_MIPS/Register/n389 ,
         \i_MIPS/Register/n388 , \i_MIPS/Register/n387 ,
         \i_MIPS/Register/n386 , \i_MIPS/Register/n385 ,
         \i_MIPS/Register/n384 , \i_MIPS/Register/n383 ,
         \i_MIPS/Register/n382 , \i_MIPS/Register/n381 ,
         \i_MIPS/Register/n380 , \i_MIPS/Register/n379 ,
         \i_MIPS/Register/n378 , \i_MIPS/Register/n377 ,
         \i_MIPS/Register/n376 , \i_MIPS/Register/n375 ,
         \i_MIPS/Register/n374 , \i_MIPS/Register/n373 ,
         \i_MIPS/Register/n372 , \i_MIPS/Register/n371 ,
         \i_MIPS/Register/n370 , \i_MIPS/Register/n369 ,
         \i_MIPS/Register/n368 , \i_MIPS/Register/n367 ,
         \i_MIPS/Register/n366 , \i_MIPS/Register/n365 ,
         \i_MIPS/Register/n364 , \i_MIPS/Register/n363 ,
         \i_MIPS/Register/n362 , \i_MIPS/Register/n361 ,
         \i_MIPS/Register/n360 , \i_MIPS/Register/n359 ,
         \i_MIPS/Register/n358 , \i_MIPS/Register/n357 ,
         \i_MIPS/Register/n356 , \i_MIPS/Register/n355 ,
         \i_MIPS/Register/n354 , \i_MIPS/Register/n353 ,
         \i_MIPS/Register/n352 , \i_MIPS/Register/n351 ,
         \i_MIPS/Register/n350 , \i_MIPS/Register/n349 ,
         \i_MIPS/Register/n348 , \i_MIPS/Register/n347 ,
         \i_MIPS/Register/n346 , \i_MIPS/Register/n345 ,
         \i_MIPS/Register/n344 , \i_MIPS/Register/n343 ,
         \i_MIPS/Register/n342 , \i_MIPS/Register/n341 ,
         \i_MIPS/Register/n340 , \i_MIPS/Register/n339 ,
         \i_MIPS/Register/n338 , \i_MIPS/Register/n337 ,
         \i_MIPS/Register/n336 , \i_MIPS/Register/n335 ,
         \i_MIPS/Register/n334 , \i_MIPS/Register/n333 ,
         \i_MIPS/Register/n332 , \i_MIPS/Register/n331 ,
         \i_MIPS/Register/n330 , \i_MIPS/Register/n329 ,
         \i_MIPS/Register/n328 , \i_MIPS/Register/n327 ,
         \i_MIPS/Register/n326 , \i_MIPS/Register/n325 ,
         \i_MIPS/Register/n324 , \i_MIPS/Register/n323 ,
         \i_MIPS/Register/n322 , \i_MIPS/Register/n321 ,
         \i_MIPS/Register/n320 , \i_MIPS/Register/n319 ,
         \i_MIPS/Register/n318 , \i_MIPS/Register/n317 ,
         \i_MIPS/Register/n316 , \i_MIPS/Register/n315 ,
         \i_MIPS/Register/n314 , \i_MIPS/Register/n313 ,
         \i_MIPS/Register/n312 , \i_MIPS/Register/n311 ,
         \i_MIPS/Register/n310 , \i_MIPS/Register/n309 ,
         \i_MIPS/Register/n308 , \i_MIPS/Register/n307 ,
         \i_MIPS/Register/n306 , \i_MIPS/Register/n305 ,
         \i_MIPS/Register/n304 , \i_MIPS/Register/n303 ,
         \i_MIPS/Register/n302 , \i_MIPS/Register/n301 ,
         \i_MIPS/Register/n300 , \i_MIPS/Register/n299 ,
         \i_MIPS/Register/n298 , \i_MIPS/Register/n297 ,
         \i_MIPS/Register/n296 , \i_MIPS/Register/n295 ,
         \i_MIPS/Register/n294 , \i_MIPS/Register/n293 ,
         \i_MIPS/Register/n292 , \i_MIPS/Register/n291 ,
         \i_MIPS/Register/n290 , \i_MIPS/Register/n289 ,
         \i_MIPS/Register/n288 , \i_MIPS/Register/n287 ,
         \i_MIPS/Register/n286 , \i_MIPS/Register/n285 ,
         \i_MIPS/Register/n284 , \i_MIPS/Register/n283 ,
         \i_MIPS/Register/n282 , \i_MIPS/Register/n281 ,
         \i_MIPS/Register/n280 , \i_MIPS/Register/n279 ,
         \i_MIPS/Register/n278 , \i_MIPS/Register/n277 ,
         \i_MIPS/Register/n276 , \i_MIPS/Register/n275 ,
         \i_MIPS/Register/n274 , \i_MIPS/Register/n273 ,
         \i_MIPS/Register/n272 , \i_MIPS/Register/n271 ,
         \i_MIPS/Register/n270 , \i_MIPS/Register/n269 ,
         \i_MIPS/Register/n268 , \i_MIPS/Register/n267 ,
         \i_MIPS/Register/n266 , \i_MIPS/Register/n265 ,
         \i_MIPS/Register/n264 , \i_MIPS/Register/n263 ,
         \i_MIPS/Register/n262 , \i_MIPS/Register/n261 ,
         \i_MIPS/Register/n260 , \i_MIPS/Register/n259 ,
         \i_MIPS/Register/n258 , \i_MIPS/Register/n257 ,
         \i_MIPS/Register/n256 , \i_MIPS/Register/n255 ,
         \i_MIPS/Register/n254 , \i_MIPS/Register/n253 ,
         \i_MIPS/Register/n252 , \i_MIPS/Register/n251 ,
         \i_MIPS/Register/n250 , \i_MIPS/Register/n249 ,
         \i_MIPS/Register/n248 , \i_MIPS/Register/n247 ,
         \i_MIPS/Register/n246 , \i_MIPS/Register/n245 ,
         \i_MIPS/Register/n244 , \i_MIPS/Register/n243 ,
         \i_MIPS/Register/n242 , \i_MIPS/Register/n241 ,
         \i_MIPS/Register/n240 , \i_MIPS/Register/n239 ,
         \i_MIPS/Register/n238 , \i_MIPS/Register/n237 ,
         \i_MIPS/Register/n236 , \i_MIPS/Register/n235 ,
         \i_MIPS/Register/n234 , \i_MIPS/Register/n233 ,
         \i_MIPS/Register/n232 , \i_MIPS/Register/n231 ,
         \i_MIPS/Register/n230 , \i_MIPS/Register/n229 ,
         \i_MIPS/Register/n228 , \i_MIPS/Register/n227 ,
         \i_MIPS/Register/n226 , \i_MIPS/Register/n225 ,
         \i_MIPS/Register/n224 , \i_MIPS/Register/n223 ,
         \i_MIPS/Register/n222 , \i_MIPS/Register/n221 ,
         \i_MIPS/Register/n220 , \i_MIPS/Register/n219 ,
         \i_MIPS/Register/n218 , \i_MIPS/Register/n217 ,
         \i_MIPS/Register/n216 , \i_MIPS/Register/n215 ,
         \i_MIPS/Register/n214 , \i_MIPS/Register/n213 ,
         \i_MIPS/Register/n212 , \i_MIPS/Register/n211 ,
         \i_MIPS/Register/n210 , \i_MIPS/Register/n209 ,
         \i_MIPS/Register/n208 , \i_MIPS/Register/n207 ,
         \i_MIPS/Register/n206 , \i_MIPS/Register/n205 ,
         \i_MIPS/Register/n204 , \i_MIPS/Register/n203 ,
         \i_MIPS/Register/n202 , \i_MIPS/Register/n201 ,
         \i_MIPS/Register/n200 , \i_MIPS/Register/n199 ,
         \i_MIPS/Register/n198 , \i_MIPS/Register/n197 ,
         \i_MIPS/Register/n196 , \i_MIPS/Register/n195 ,
         \i_MIPS/Register/n194 , \i_MIPS/Register/n193 ,
         \i_MIPS/Register/n192 , \i_MIPS/Register/n191 ,
         \i_MIPS/Register/n190 , \i_MIPS/Register/n189 ,
         \i_MIPS/Register/n188 , \i_MIPS/Register/n187 ,
         \i_MIPS/Register/n186 , \i_MIPS/Register/n185 ,
         \i_MIPS/Register/n184 , \i_MIPS/Register/n183 ,
         \i_MIPS/Register/n182 , \i_MIPS/Register/n181 ,
         \i_MIPS/Register/n180 , \i_MIPS/Register/n179 ,
         \i_MIPS/Register/n178 , \i_MIPS/Register/n177 ,
         \i_MIPS/Register/n176 , \i_MIPS/Register/n175 ,
         \i_MIPS/Register/n174 , \i_MIPS/Register/n173 ,
         \i_MIPS/Register/n172 , \i_MIPS/Register/n171 ,
         \i_MIPS/Register/n170 , \i_MIPS/Register/n169 ,
         \i_MIPS/Register/n168 , \i_MIPS/Register/n167 ,
         \i_MIPS/Register/n166 , \i_MIPS/Register/n165 ,
         \i_MIPS/Register/n164 , \i_MIPS/Register/n163 ,
         \i_MIPS/Register/n162 , \i_MIPS/Register/n161 ,
         \i_MIPS/Register/n160 , \i_MIPS/Register/n159 ,
         \i_MIPS/Register/n158 , \i_MIPS/Register/n157 ,
         \i_MIPS/Register/n156 , \i_MIPS/Register/n155 ,
         \i_MIPS/Register/n154 , \i_MIPS/Register/n153 ,
         \i_MIPS/Register/n152 , \i_MIPS/Register/n151 ,
         \i_MIPS/Register/n150 , \i_MIPS/Register/n149 ,
         \i_MIPS/Register/n148 , \i_MIPS/Register/n147 ,
         \i_MIPS/Register/n146 , \i_MIPS/Register/n145 ,
         \i_MIPS/Register/n144 , \i_MIPS/Register/n143 ,
         \i_MIPS/Register/n142 , \i_MIPS/Register/n141 ,
         \i_MIPS/Register/n140 , \i_MIPS/Register/n139 ,
         \i_MIPS/Register/n138 , \i_MIPS/Register/n137 ,
         \i_MIPS/Register/n136 , \i_MIPS/Register/n135 ,
         \i_MIPS/Register/n134 , \i_MIPS/Register/n133 ,
         \i_MIPS/Register/n132 , \i_MIPS/Register/n131 ,
         \i_MIPS/Register/n130 , \i_MIPS/Register/n129 ,
         \i_MIPS/Register/n128 , \i_MIPS/Register/n127 ,
         \i_MIPS/Register/n126 , \i_MIPS/Register/n125 ,
         \i_MIPS/Register/n124 , \i_MIPS/Register/n123 ,
         \i_MIPS/Register/n122 , \i_MIPS/Register/n121 ,
         \i_MIPS/Register/n120 , \i_MIPS/Register/n119 ,
         \i_MIPS/Register/n118 , \i_MIPS/Register/n117 ,
         \i_MIPS/Register/n116 , \i_MIPS/Register/n115 ,
         \i_MIPS/Register/n114 , \i_MIPS/Register/n113 ,
         \i_MIPS/Register/n112 , \i_MIPS/Register/n111 ,
         \i_MIPS/Register/n110 , \i_MIPS/Register/n109 ,
         \i_MIPS/Register/n108 , \i_MIPS/Register/n107 ,
         \i_MIPS/Register/n106 , \i_MIPS/Register/n105 ,
         \i_MIPS/Register/n104 , \i_MIPS/Register/register[31][0] ,
         \i_MIPS/Register/register[31][1] , \i_MIPS/Register/register[31][2] ,
         \i_MIPS/Register/register[31][3] , \i_MIPS/Register/register[31][4] ,
         \i_MIPS/Register/register[31][5] , \i_MIPS/Register/register[31][6] ,
         \i_MIPS/Register/register[31][7] , \i_MIPS/Register/register[31][8] ,
         \i_MIPS/Register/register[31][9] , \i_MIPS/Register/register[31][10] ,
         \i_MIPS/Register/register[31][11] ,
         \i_MIPS/Register/register[31][12] ,
         \i_MIPS/Register/register[31][13] ,
         \i_MIPS/Register/register[31][14] ,
         \i_MIPS/Register/register[31][15] ,
         \i_MIPS/Register/register[31][16] ,
         \i_MIPS/Register/register[31][17] ,
         \i_MIPS/Register/register[31][18] ,
         \i_MIPS/Register/register[31][20] ,
         \i_MIPS/Register/register[31][21] ,
         \i_MIPS/Register/register[31][22] ,
         \i_MIPS/Register/register[31][23] ,
         \i_MIPS/Register/register[31][24] ,
         \i_MIPS/Register/register[31][25] ,
         \i_MIPS/Register/register[31][26] ,
         \i_MIPS/Register/register[31][27] ,
         \i_MIPS/Register/register[31][28] ,
         \i_MIPS/Register/register[31][29] ,
         \i_MIPS/Register/register[31][31] , \i_MIPS/Register/register[30][0] ,
         \i_MIPS/Register/register[30][1] , \i_MIPS/Register/register[30][2] ,
         \i_MIPS/Register/register[30][3] , \i_MIPS/Register/register[30][4] ,
         \i_MIPS/Register/register[30][5] , \i_MIPS/Register/register[30][6] ,
         \i_MIPS/Register/register[30][7] , \i_MIPS/Register/register[30][8] ,
         \i_MIPS/Register/register[30][9] , \i_MIPS/Register/register[30][10] ,
         \i_MIPS/Register/register[30][11] ,
         \i_MIPS/Register/register[30][12] ,
         \i_MIPS/Register/register[30][13] ,
         \i_MIPS/Register/register[30][14] ,
         \i_MIPS/Register/register[30][15] ,
         \i_MIPS/Register/register[30][16] ,
         \i_MIPS/Register/register[30][17] ,
         \i_MIPS/Register/register[30][18] ,
         \i_MIPS/Register/register[30][19] ,
         \i_MIPS/Register/register[30][20] ,
         \i_MIPS/Register/register[30][21] ,
         \i_MIPS/Register/register[30][22] ,
         \i_MIPS/Register/register[30][23] ,
         \i_MIPS/Register/register[30][24] ,
         \i_MIPS/Register/register[30][25] ,
         \i_MIPS/Register/register[30][26] ,
         \i_MIPS/Register/register[30][27] ,
         \i_MIPS/Register/register[30][28] ,
         \i_MIPS/Register/register[30][29] ,
         \i_MIPS/Register/register[30][30] ,
         \i_MIPS/Register/register[30][31] , \i_MIPS/Register/register[29][0] ,
         \i_MIPS/Register/register[29][1] , \i_MIPS/Register/register[29][2] ,
         \i_MIPS/Register/register[29][3] , \i_MIPS/Register/register[29][4] ,
         \i_MIPS/Register/register[29][5] , \i_MIPS/Register/register[29][6] ,
         \i_MIPS/Register/register[29][7] , \i_MIPS/Register/register[29][8] ,
         \i_MIPS/Register/register[29][9] , \i_MIPS/Register/register[29][10] ,
         \i_MIPS/Register/register[29][11] ,
         \i_MIPS/Register/register[29][12] ,
         \i_MIPS/Register/register[29][13] ,
         \i_MIPS/Register/register[29][14] ,
         \i_MIPS/Register/register[29][15] ,
         \i_MIPS/Register/register[29][16] ,
         \i_MIPS/Register/register[29][17] ,
         \i_MIPS/Register/register[29][18] ,
         \i_MIPS/Register/register[29][19] ,
         \i_MIPS/Register/register[29][20] ,
         \i_MIPS/Register/register[29][21] ,
         \i_MIPS/Register/register[29][22] ,
         \i_MIPS/Register/register[29][23] ,
         \i_MIPS/Register/register[29][24] ,
         \i_MIPS/Register/register[29][25] ,
         \i_MIPS/Register/register[29][26] ,
         \i_MIPS/Register/register[29][27] ,
         \i_MIPS/Register/register[29][28] ,
         \i_MIPS/Register/register[29][29] ,
         \i_MIPS/Register/register[29][30] ,
         \i_MIPS/Register/register[29][31] , \i_MIPS/Register/register[28][0] ,
         \i_MIPS/Register/register[28][1] , \i_MIPS/Register/register[28][2] ,
         \i_MIPS/Register/register[28][3] , \i_MIPS/Register/register[28][4] ,
         \i_MIPS/Register/register[28][5] , \i_MIPS/Register/register[28][6] ,
         \i_MIPS/Register/register[28][7] , \i_MIPS/Register/register[28][8] ,
         \i_MIPS/Register/register[28][9] , \i_MIPS/Register/register[28][10] ,
         \i_MIPS/Register/register[28][11] ,
         \i_MIPS/Register/register[28][12] ,
         \i_MIPS/Register/register[28][13] ,
         \i_MIPS/Register/register[28][14] ,
         \i_MIPS/Register/register[28][15] ,
         \i_MIPS/Register/register[28][16] ,
         \i_MIPS/Register/register[28][17] ,
         \i_MIPS/Register/register[28][18] ,
         \i_MIPS/Register/register[28][19] ,
         \i_MIPS/Register/register[28][20] ,
         \i_MIPS/Register/register[28][21] ,
         \i_MIPS/Register/register[28][22] ,
         \i_MIPS/Register/register[28][23] ,
         \i_MIPS/Register/register[28][24] ,
         \i_MIPS/Register/register[28][25] ,
         \i_MIPS/Register/register[28][26] ,
         \i_MIPS/Register/register[28][27] ,
         \i_MIPS/Register/register[28][28] ,
         \i_MIPS/Register/register[28][29] ,
         \i_MIPS/Register/register[28][30] ,
         \i_MIPS/Register/register[28][31] , \i_MIPS/Register/register[27][0] ,
         \i_MIPS/Register/register[27][1] , \i_MIPS/Register/register[27][2] ,
         \i_MIPS/Register/register[27][3] , \i_MIPS/Register/register[27][4] ,
         \i_MIPS/Register/register[27][5] , \i_MIPS/Register/register[27][6] ,
         \i_MIPS/Register/register[27][7] , \i_MIPS/Register/register[27][8] ,
         \i_MIPS/Register/register[27][9] , \i_MIPS/Register/register[27][10] ,
         \i_MIPS/Register/register[27][11] ,
         \i_MIPS/Register/register[27][12] ,
         \i_MIPS/Register/register[27][13] ,
         \i_MIPS/Register/register[27][14] ,
         \i_MIPS/Register/register[27][15] ,
         \i_MIPS/Register/register[27][16] ,
         \i_MIPS/Register/register[27][17] ,
         \i_MIPS/Register/register[27][18] ,
         \i_MIPS/Register/register[27][19] ,
         \i_MIPS/Register/register[27][20] ,
         \i_MIPS/Register/register[27][21] ,
         \i_MIPS/Register/register[27][22] ,
         \i_MIPS/Register/register[27][23] ,
         \i_MIPS/Register/register[27][24] ,
         \i_MIPS/Register/register[27][25] ,
         \i_MIPS/Register/register[27][26] ,
         \i_MIPS/Register/register[27][27] ,
         \i_MIPS/Register/register[27][28] ,
         \i_MIPS/Register/register[27][29] ,
         \i_MIPS/Register/register[27][30] ,
         \i_MIPS/Register/register[27][31] , \i_MIPS/Register/register[26][0] ,
         \i_MIPS/Register/register[26][1] , \i_MIPS/Register/register[26][2] ,
         \i_MIPS/Register/register[26][3] , \i_MIPS/Register/register[26][4] ,
         \i_MIPS/Register/register[26][5] , \i_MIPS/Register/register[26][6] ,
         \i_MIPS/Register/register[26][7] , \i_MIPS/Register/register[26][8] ,
         \i_MIPS/Register/register[26][9] , \i_MIPS/Register/register[26][10] ,
         \i_MIPS/Register/register[26][11] ,
         \i_MIPS/Register/register[26][12] ,
         \i_MIPS/Register/register[26][13] ,
         \i_MIPS/Register/register[26][14] ,
         \i_MIPS/Register/register[26][15] ,
         \i_MIPS/Register/register[26][16] ,
         \i_MIPS/Register/register[26][17] ,
         \i_MIPS/Register/register[26][18] ,
         \i_MIPS/Register/register[26][19] ,
         \i_MIPS/Register/register[26][20] ,
         \i_MIPS/Register/register[26][21] ,
         \i_MIPS/Register/register[26][22] ,
         \i_MIPS/Register/register[26][23] ,
         \i_MIPS/Register/register[26][24] ,
         \i_MIPS/Register/register[26][25] ,
         \i_MIPS/Register/register[26][26] ,
         \i_MIPS/Register/register[26][27] ,
         \i_MIPS/Register/register[26][28] ,
         \i_MIPS/Register/register[26][29] ,
         \i_MIPS/Register/register[26][30] ,
         \i_MIPS/Register/register[26][31] , \i_MIPS/Register/register[25][0] ,
         \i_MIPS/Register/register[25][1] , \i_MIPS/Register/register[25][2] ,
         \i_MIPS/Register/register[25][3] , \i_MIPS/Register/register[25][4] ,
         \i_MIPS/Register/register[25][5] , \i_MIPS/Register/register[25][6] ,
         \i_MIPS/Register/register[25][7] , \i_MIPS/Register/register[25][8] ,
         \i_MIPS/Register/register[25][9] , \i_MIPS/Register/register[25][10] ,
         \i_MIPS/Register/register[25][11] ,
         \i_MIPS/Register/register[25][12] ,
         \i_MIPS/Register/register[25][13] ,
         \i_MIPS/Register/register[25][14] ,
         \i_MIPS/Register/register[25][15] ,
         \i_MIPS/Register/register[25][16] ,
         \i_MIPS/Register/register[25][17] ,
         \i_MIPS/Register/register[25][18] ,
         \i_MIPS/Register/register[25][19] ,
         \i_MIPS/Register/register[25][20] ,
         \i_MIPS/Register/register[25][21] ,
         \i_MIPS/Register/register[25][22] ,
         \i_MIPS/Register/register[25][23] ,
         \i_MIPS/Register/register[25][24] ,
         \i_MIPS/Register/register[25][25] ,
         \i_MIPS/Register/register[25][26] ,
         \i_MIPS/Register/register[25][27] ,
         \i_MIPS/Register/register[25][28] ,
         \i_MIPS/Register/register[25][29] ,
         \i_MIPS/Register/register[25][30] ,
         \i_MIPS/Register/register[25][31] , \i_MIPS/Register/register[24][0] ,
         \i_MIPS/Register/register[24][1] , \i_MIPS/Register/register[24][2] ,
         \i_MIPS/Register/register[24][3] , \i_MIPS/Register/register[24][4] ,
         \i_MIPS/Register/register[24][5] , \i_MIPS/Register/register[24][6] ,
         \i_MIPS/Register/register[24][7] , \i_MIPS/Register/register[24][8] ,
         \i_MIPS/Register/register[24][9] , \i_MIPS/Register/register[24][10] ,
         \i_MIPS/Register/register[24][11] ,
         \i_MIPS/Register/register[24][12] ,
         \i_MIPS/Register/register[24][13] ,
         \i_MIPS/Register/register[24][14] ,
         \i_MIPS/Register/register[24][15] ,
         \i_MIPS/Register/register[24][16] ,
         \i_MIPS/Register/register[24][17] ,
         \i_MIPS/Register/register[24][18] ,
         \i_MIPS/Register/register[24][19] ,
         \i_MIPS/Register/register[24][20] ,
         \i_MIPS/Register/register[24][21] ,
         \i_MIPS/Register/register[24][22] ,
         \i_MIPS/Register/register[24][23] ,
         \i_MIPS/Register/register[24][24] ,
         \i_MIPS/Register/register[24][25] ,
         \i_MIPS/Register/register[24][26] ,
         \i_MIPS/Register/register[24][27] ,
         \i_MIPS/Register/register[24][28] ,
         \i_MIPS/Register/register[24][29] ,
         \i_MIPS/Register/register[24][30] ,
         \i_MIPS/Register/register[24][31] , \i_MIPS/Register/register[23][0] ,
         \i_MIPS/Register/register[23][1] , \i_MIPS/Register/register[23][2] ,
         \i_MIPS/Register/register[23][3] , \i_MIPS/Register/register[23][4] ,
         \i_MIPS/Register/register[23][5] , \i_MIPS/Register/register[23][6] ,
         \i_MIPS/Register/register[23][7] , \i_MIPS/Register/register[23][8] ,
         \i_MIPS/Register/register[23][9] , \i_MIPS/Register/register[23][10] ,
         \i_MIPS/Register/register[23][11] ,
         \i_MIPS/Register/register[23][12] ,
         \i_MIPS/Register/register[23][13] ,
         \i_MIPS/Register/register[23][14] ,
         \i_MIPS/Register/register[23][15] ,
         \i_MIPS/Register/register[23][16] ,
         \i_MIPS/Register/register[23][17] ,
         \i_MIPS/Register/register[23][18] ,
         \i_MIPS/Register/register[23][19] ,
         \i_MIPS/Register/register[23][20] ,
         \i_MIPS/Register/register[23][21] ,
         \i_MIPS/Register/register[23][22] ,
         \i_MIPS/Register/register[23][23] ,
         \i_MIPS/Register/register[23][24] ,
         \i_MIPS/Register/register[23][25] ,
         \i_MIPS/Register/register[23][26] ,
         \i_MIPS/Register/register[23][27] ,
         \i_MIPS/Register/register[23][28] ,
         \i_MIPS/Register/register[23][29] ,
         \i_MIPS/Register/register[23][30] ,
         \i_MIPS/Register/register[23][31] , \i_MIPS/Register/register[22][0] ,
         \i_MIPS/Register/register[22][1] , \i_MIPS/Register/register[22][2] ,
         \i_MIPS/Register/register[22][3] , \i_MIPS/Register/register[22][4] ,
         \i_MIPS/Register/register[22][5] , \i_MIPS/Register/register[22][6] ,
         \i_MIPS/Register/register[22][7] , \i_MIPS/Register/register[22][8] ,
         \i_MIPS/Register/register[22][9] , \i_MIPS/Register/register[22][10] ,
         \i_MIPS/Register/register[22][11] ,
         \i_MIPS/Register/register[22][12] ,
         \i_MIPS/Register/register[22][13] ,
         \i_MIPS/Register/register[22][14] ,
         \i_MIPS/Register/register[22][15] ,
         \i_MIPS/Register/register[22][16] ,
         \i_MIPS/Register/register[22][17] ,
         \i_MIPS/Register/register[22][18] ,
         \i_MIPS/Register/register[22][19] ,
         \i_MIPS/Register/register[22][20] ,
         \i_MIPS/Register/register[22][21] ,
         \i_MIPS/Register/register[22][22] ,
         \i_MIPS/Register/register[22][23] ,
         \i_MIPS/Register/register[22][24] ,
         \i_MIPS/Register/register[22][25] ,
         \i_MIPS/Register/register[22][26] ,
         \i_MIPS/Register/register[22][27] ,
         \i_MIPS/Register/register[22][28] ,
         \i_MIPS/Register/register[22][29] ,
         \i_MIPS/Register/register[22][30] ,
         \i_MIPS/Register/register[22][31] , \i_MIPS/Register/register[21][0] ,
         \i_MIPS/Register/register[21][1] , \i_MIPS/Register/register[21][2] ,
         \i_MIPS/Register/register[21][3] , \i_MIPS/Register/register[21][4] ,
         \i_MIPS/Register/register[21][5] , \i_MIPS/Register/register[21][6] ,
         \i_MIPS/Register/register[21][7] , \i_MIPS/Register/register[21][8] ,
         \i_MIPS/Register/register[21][9] , \i_MIPS/Register/register[21][10] ,
         \i_MIPS/Register/register[21][11] ,
         \i_MIPS/Register/register[21][12] ,
         \i_MIPS/Register/register[21][13] ,
         \i_MIPS/Register/register[21][14] ,
         \i_MIPS/Register/register[21][15] ,
         \i_MIPS/Register/register[21][16] ,
         \i_MIPS/Register/register[21][17] ,
         \i_MIPS/Register/register[21][18] ,
         \i_MIPS/Register/register[21][19] ,
         \i_MIPS/Register/register[21][20] ,
         \i_MIPS/Register/register[21][21] ,
         \i_MIPS/Register/register[21][22] ,
         \i_MIPS/Register/register[21][23] ,
         \i_MIPS/Register/register[21][24] ,
         \i_MIPS/Register/register[21][25] ,
         \i_MIPS/Register/register[21][26] ,
         \i_MIPS/Register/register[21][27] ,
         \i_MIPS/Register/register[21][28] ,
         \i_MIPS/Register/register[21][29] ,
         \i_MIPS/Register/register[21][30] ,
         \i_MIPS/Register/register[21][31] , \i_MIPS/Register/register[20][0] ,
         \i_MIPS/Register/register[20][1] , \i_MIPS/Register/register[20][2] ,
         \i_MIPS/Register/register[20][3] , \i_MIPS/Register/register[20][4] ,
         \i_MIPS/Register/register[20][5] , \i_MIPS/Register/register[20][6] ,
         \i_MIPS/Register/register[20][7] , \i_MIPS/Register/register[20][8] ,
         \i_MIPS/Register/register[20][9] , \i_MIPS/Register/register[20][10] ,
         \i_MIPS/Register/register[20][11] ,
         \i_MIPS/Register/register[20][12] ,
         \i_MIPS/Register/register[20][13] ,
         \i_MIPS/Register/register[20][14] ,
         \i_MIPS/Register/register[20][15] ,
         \i_MIPS/Register/register[20][16] ,
         \i_MIPS/Register/register[20][17] ,
         \i_MIPS/Register/register[20][18] ,
         \i_MIPS/Register/register[20][19] ,
         \i_MIPS/Register/register[20][20] ,
         \i_MIPS/Register/register[20][21] ,
         \i_MIPS/Register/register[20][22] ,
         \i_MIPS/Register/register[20][23] ,
         \i_MIPS/Register/register[20][24] ,
         \i_MIPS/Register/register[20][25] ,
         \i_MIPS/Register/register[20][26] ,
         \i_MIPS/Register/register[20][27] ,
         \i_MIPS/Register/register[20][28] ,
         \i_MIPS/Register/register[20][29] ,
         \i_MIPS/Register/register[20][30] ,
         \i_MIPS/Register/register[20][31] , \i_MIPS/Register/register[19][0] ,
         \i_MIPS/Register/register[19][1] , \i_MIPS/Register/register[19][2] ,
         \i_MIPS/Register/register[19][3] , \i_MIPS/Register/register[19][4] ,
         \i_MIPS/Register/register[19][5] , \i_MIPS/Register/register[19][6] ,
         \i_MIPS/Register/register[19][7] , \i_MIPS/Register/register[19][8] ,
         \i_MIPS/Register/register[19][9] , \i_MIPS/Register/register[19][10] ,
         \i_MIPS/Register/register[19][11] ,
         \i_MIPS/Register/register[19][12] ,
         \i_MIPS/Register/register[19][13] ,
         \i_MIPS/Register/register[19][14] ,
         \i_MIPS/Register/register[19][15] ,
         \i_MIPS/Register/register[19][16] ,
         \i_MIPS/Register/register[19][17] ,
         \i_MIPS/Register/register[19][18] ,
         \i_MIPS/Register/register[19][19] ,
         \i_MIPS/Register/register[19][20] ,
         \i_MIPS/Register/register[19][21] ,
         \i_MIPS/Register/register[19][22] ,
         \i_MIPS/Register/register[19][23] ,
         \i_MIPS/Register/register[19][24] ,
         \i_MIPS/Register/register[19][25] ,
         \i_MIPS/Register/register[19][26] ,
         \i_MIPS/Register/register[19][27] ,
         \i_MIPS/Register/register[19][28] ,
         \i_MIPS/Register/register[19][29] ,
         \i_MIPS/Register/register[19][30] ,
         \i_MIPS/Register/register[19][31] , \i_MIPS/Register/register[18][0] ,
         \i_MIPS/Register/register[18][1] , \i_MIPS/Register/register[18][2] ,
         \i_MIPS/Register/register[18][3] , \i_MIPS/Register/register[18][4] ,
         \i_MIPS/Register/register[18][5] , \i_MIPS/Register/register[18][6] ,
         \i_MIPS/Register/register[18][7] , \i_MIPS/Register/register[18][8] ,
         \i_MIPS/Register/register[18][9] , \i_MIPS/Register/register[18][10] ,
         \i_MIPS/Register/register[18][11] ,
         \i_MIPS/Register/register[18][12] ,
         \i_MIPS/Register/register[18][13] ,
         \i_MIPS/Register/register[18][14] ,
         \i_MIPS/Register/register[18][15] ,
         \i_MIPS/Register/register[18][16] ,
         \i_MIPS/Register/register[18][17] ,
         \i_MIPS/Register/register[18][18] ,
         \i_MIPS/Register/register[18][19] ,
         \i_MIPS/Register/register[18][20] ,
         \i_MIPS/Register/register[18][21] ,
         \i_MIPS/Register/register[18][22] ,
         \i_MIPS/Register/register[18][23] ,
         \i_MIPS/Register/register[18][24] ,
         \i_MIPS/Register/register[18][25] ,
         \i_MIPS/Register/register[18][26] ,
         \i_MIPS/Register/register[18][27] ,
         \i_MIPS/Register/register[18][28] ,
         \i_MIPS/Register/register[18][29] ,
         \i_MIPS/Register/register[18][30] ,
         \i_MIPS/Register/register[18][31] , \i_MIPS/Register/register[17][0] ,
         \i_MIPS/Register/register[17][1] , \i_MIPS/Register/register[17][2] ,
         \i_MIPS/Register/register[17][3] , \i_MIPS/Register/register[17][4] ,
         \i_MIPS/Register/register[17][5] , \i_MIPS/Register/register[17][6] ,
         \i_MIPS/Register/register[17][7] , \i_MIPS/Register/register[17][8] ,
         \i_MIPS/Register/register[17][9] , \i_MIPS/Register/register[17][10] ,
         \i_MIPS/Register/register[17][11] ,
         \i_MIPS/Register/register[17][12] ,
         \i_MIPS/Register/register[17][13] ,
         \i_MIPS/Register/register[17][14] ,
         \i_MIPS/Register/register[17][15] ,
         \i_MIPS/Register/register[17][16] ,
         \i_MIPS/Register/register[17][17] ,
         \i_MIPS/Register/register[17][18] ,
         \i_MIPS/Register/register[17][19] ,
         \i_MIPS/Register/register[17][20] ,
         \i_MIPS/Register/register[17][21] ,
         \i_MIPS/Register/register[17][22] ,
         \i_MIPS/Register/register[17][23] ,
         \i_MIPS/Register/register[17][24] ,
         \i_MIPS/Register/register[17][25] ,
         \i_MIPS/Register/register[17][26] ,
         \i_MIPS/Register/register[17][27] ,
         \i_MIPS/Register/register[17][28] ,
         \i_MIPS/Register/register[17][29] ,
         \i_MIPS/Register/register[17][30] ,
         \i_MIPS/Register/register[17][31] , \i_MIPS/Register/register[16][0] ,
         \i_MIPS/Register/register[16][1] , \i_MIPS/Register/register[16][2] ,
         \i_MIPS/Register/register[16][3] , \i_MIPS/Register/register[16][4] ,
         \i_MIPS/Register/register[16][5] , \i_MIPS/Register/register[16][6] ,
         \i_MIPS/Register/register[16][7] , \i_MIPS/Register/register[16][8] ,
         \i_MIPS/Register/register[16][9] , \i_MIPS/Register/register[16][10] ,
         \i_MIPS/Register/register[16][11] ,
         \i_MIPS/Register/register[16][12] ,
         \i_MIPS/Register/register[16][13] ,
         \i_MIPS/Register/register[16][14] ,
         \i_MIPS/Register/register[16][15] ,
         \i_MIPS/Register/register[16][16] ,
         \i_MIPS/Register/register[16][17] ,
         \i_MIPS/Register/register[16][18] ,
         \i_MIPS/Register/register[16][19] ,
         \i_MIPS/Register/register[16][20] ,
         \i_MIPS/Register/register[16][21] ,
         \i_MIPS/Register/register[16][22] ,
         \i_MIPS/Register/register[16][23] ,
         \i_MIPS/Register/register[16][24] ,
         \i_MIPS/Register/register[16][25] ,
         \i_MIPS/Register/register[16][26] ,
         \i_MIPS/Register/register[16][27] ,
         \i_MIPS/Register/register[16][28] ,
         \i_MIPS/Register/register[16][29] ,
         \i_MIPS/Register/register[16][30] ,
         \i_MIPS/Register/register[16][31] , \i_MIPS/Register/register[15][0] ,
         \i_MIPS/Register/register[15][1] , \i_MIPS/Register/register[15][2] ,
         \i_MIPS/Register/register[15][3] , \i_MIPS/Register/register[15][4] ,
         \i_MIPS/Register/register[15][5] , \i_MIPS/Register/register[15][6] ,
         \i_MIPS/Register/register[15][7] , \i_MIPS/Register/register[15][8] ,
         \i_MIPS/Register/register[15][9] , \i_MIPS/Register/register[15][10] ,
         \i_MIPS/Register/register[15][11] ,
         \i_MIPS/Register/register[15][12] ,
         \i_MIPS/Register/register[15][13] ,
         \i_MIPS/Register/register[15][14] ,
         \i_MIPS/Register/register[15][15] ,
         \i_MIPS/Register/register[15][16] ,
         \i_MIPS/Register/register[15][17] ,
         \i_MIPS/Register/register[15][18] ,
         \i_MIPS/Register/register[15][19] ,
         \i_MIPS/Register/register[15][20] ,
         \i_MIPS/Register/register[15][21] ,
         \i_MIPS/Register/register[15][22] ,
         \i_MIPS/Register/register[15][23] ,
         \i_MIPS/Register/register[15][24] ,
         \i_MIPS/Register/register[15][25] ,
         \i_MIPS/Register/register[15][26] ,
         \i_MIPS/Register/register[15][27] ,
         \i_MIPS/Register/register[15][28] ,
         \i_MIPS/Register/register[15][29] ,
         \i_MIPS/Register/register[15][30] ,
         \i_MIPS/Register/register[15][31] , \i_MIPS/Register/register[14][0] ,
         \i_MIPS/Register/register[14][1] , \i_MIPS/Register/register[14][2] ,
         \i_MIPS/Register/register[14][3] , \i_MIPS/Register/register[14][4] ,
         \i_MIPS/Register/register[14][5] , \i_MIPS/Register/register[14][6] ,
         \i_MIPS/Register/register[14][7] , \i_MIPS/Register/register[14][8] ,
         \i_MIPS/Register/register[14][9] , \i_MIPS/Register/register[14][10] ,
         \i_MIPS/Register/register[14][11] ,
         \i_MIPS/Register/register[14][12] ,
         \i_MIPS/Register/register[14][13] ,
         \i_MIPS/Register/register[14][14] ,
         \i_MIPS/Register/register[14][15] ,
         \i_MIPS/Register/register[14][16] ,
         \i_MIPS/Register/register[14][17] ,
         \i_MIPS/Register/register[14][18] ,
         \i_MIPS/Register/register[14][19] ,
         \i_MIPS/Register/register[14][20] ,
         \i_MIPS/Register/register[14][21] ,
         \i_MIPS/Register/register[14][22] ,
         \i_MIPS/Register/register[14][23] ,
         \i_MIPS/Register/register[14][24] ,
         \i_MIPS/Register/register[14][25] ,
         \i_MIPS/Register/register[14][26] ,
         \i_MIPS/Register/register[14][27] ,
         \i_MIPS/Register/register[14][28] ,
         \i_MIPS/Register/register[14][29] ,
         \i_MIPS/Register/register[14][30] ,
         \i_MIPS/Register/register[14][31] , \i_MIPS/Register/register[13][0] ,
         \i_MIPS/Register/register[13][1] , \i_MIPS/Register/register[13][2] ,
         \i_MIPS/Register/register[13][3] , \i_MIPS/Register/register[13][4] ,
         \i_MIPS/Register/register[13][5] , \i_MIPS/Register/register[13][6] ,
         \i_MIPS/Register/register[13][7] , \i_MIPS/Register/register[13][8] ,
         \i_MIPS/Register/register[13][9] , \i_MIPS/Register/register[13][10] ,
         \i_MIPS/Register/register[13][11] ,
         \i_MIPS/Register/register[13][12] ,
         \i_MIPS/Register/register[13][13] ,
         \i_MIPS/Register/register[13][14] ,
         \i_MIPS/Register/register[13][15] ,
         \i_MIPS/Register/register[13][16] ,
         \i_MIPS/Register/register[13][17] ,
         \i_MIPS/Register/register[13][18] ,
         \i_MIPS/Register/register[13][19] ,
         \i_MIPS/Register/register[13][20] ,
         \i_MIPS/Register/register[13][21] ,
         \i_MIPS/Register/register[13][22] ,
         \i_MIPS/Register/register[13][23] ,
         \i_MIPS/Register/register[13][24] ,
         \i_MIPS/Register/register[13][25] ,
         \i_MIPS/Register/register[13][26] ,
         \i_MIPS/Register/register[13][27] ,
         \i_MIPS/Register/register[13][28] ,
         \i_MIPS/Register/register[13][29] ,
         \i_MIPS/Register/register[13][30] ,
         \i_MIPS/Register/register[13][31] , \i_MIPS/Register/register[12][0] ,
         \i_MIPS/Register/register[12][1] , \i_MIPS/Register/register[12][2] ,
         \i_MIPS/Register/register[12][3] , \i_MIPS/Register/register[12][4] ,
         \i_MIPS/Register/register[12][5] , \i_MIPS/Register/register[12][6] ,
         \i_MIPS/Register/register[12][7] , \i_MIPS/Register/register[12][8] ,
         \i_MIPS/Register/register[12][9] , \i_MIPS/Register/register[12][10] ,
         \i_MIPS/Register/register[12][11] ,
         \i_MIPS/Register/register[12][12] ,
         \i_MIPS/Register/register[12][13] ,
         \i_MIPS/Register/register[12][14] ,
         \i_MIPS/Register/register[12][15] ,
         \i_MIPS/Register/register[12][16] ,
         \i_MIPS/Register/register[12][17] ,
         \i_MIPS/Register/register[12][18] ,
         \i_MIPS/Register/register[12][19] ,
         \i_MIPS/Register/register[12][20] ,
         \i_MIPS/Register/register[12][21] ,
         \i_MIPS/Register/register[12][22] ,
         \i_MIPS/Register/register[12][23] ,
         \i_MIPS/Register/register[12][24] ,
         \i_MIPS/Register/register[12][25] ,
         \i_MIPS/Register/register[12][26] ,
         \i_MIPS/Register/register[12][27] ,
         \i_MIPS/Register/register[12][28] ,
         \i_MIPS/Register/register[12][29] ,
         \i_MIPS/Register/register[12][30] ,
         \i_MIPS/Register/register[12][31] , \i_MIPS/Register/register[11][0] ,
         \i_MIPS/Register/register[11][1] , \i_MIPS/Register/register[11][2] ,
         \i_MIPS/Register/register[11][3] , \i_MIPS/Register/register[11][4] ,
         \i_MIPS/Register/register[11][5] , \i_MIPS/Register/register[11][6] ,
         \i_MIPS/Register/register[11][7] , \i_MIPS/Register/register[11][8] ,
         \i_MIPS/Register/register[11][9] , \i_MIPS/Register/register[11][10] ,
         \i_MIPS/Register/register[11][11] ,
         \i_MIPS/Register/register[11][12] ,
         \i_MIPS/Register/register[11][13] ,
         \i_MIPS/Register/register[11][14] ,
         \i_MIPS/Register/register[11][15] ,
         \i_MIPS/Register/register[11][16] ,
         \i_MIPS/Register/register[11][17] ,
         \i_MIPS/Register/register[11][18] ,
         \i_MIPS/Register/register[11][19] ,
         \i_MIPS/Register/register[11][20] ,
         \i_MIPS/Register/register[11][21] ,
         \i_MIPS/Register/register[11][22] ,
         \i_MIPS/Register/register[11][23] ,
         \i_MIPS/Register/register[11][24] ,
         \i_MIPS/Register/register[11][25] ,
         \i_MIPS/Register/register[11][26] ,
         \i_MIPS/Register/register[11][27] ,
         \i_MIPS/Register/register[11][28] ,
         \i_MIPS/Register/register[11][29] ,
         \i_MIPS/Register/register[11][30] ,
         \i_MIPS/Register/register[11][31] , \i_MIPS/Register/register[10][0] ,
         \i_MIPS/Register/register[10][1] , \i_MIPS/Register/register[10][2] ,
         \i_MIPS/Register/register[10][3] , \i_MIPS/Register/register[10][4] ,
         \i_MIPS/Register/register[10][5] , \i_MIPS/Register/register[10][6] ,
         \i_MIPS/Register/register[10][7] , \i_MIPS/Register/register[10][8] ,
         \i_MIPS/Register/register[10][9] , \i_MIPS/Register/register[10][10] ,
         \i_MIPS/Register/register[10][11] ,
         \i_MIPS/Register/register[10][12] ,
         \i_MIPS/Register/register[10][13] ,
         \i_MIPS/Register/register[10][14] ,
         \i_MIPS/Register/register[10][15] ,
         \i_MIPS/Register/register[10][16] ,
         \i_MIPS/Register/register[10][17] ,
         \i_MIPS/Register/register[10][18] ,
         \i_MIPS/Register/register[10][19] ,
         \i_MIPS/Register/register[10][20] ,
         \i_MIPS/Register/register[10][21] ,
         \i_MIPS/Register/register[10][22] ,
         \i_MIPS/Register/register[10][23] ,
         \i_MIPS/Register/register[10][24] ,
         \i_MIPS/Register/register[10][25] ,
         \i_MIPS/Register/register[10][26] ,
         \i_MIPS/Register/register[10][27] ,
         \i_MIPS/Register/register[10][28] ,
         \i_MIPS/Register/register[10][29] ,
         \i_MIPS/Register/register[10][30] ,
         \i_MIPS/Register/register[10][31] , \i_MIPS/Register/register[9][0] ,
         \i_MIPS/Register/register[9][1] , \i_MIPS/Register/register[9][2] ,
         \i_MIPS/Register/register[9][3] , \i_MIPS/Register/register[9][4] ,
         \i_MIPS/Register/register[9][5] , \i_MIPS/Register/register[9][6] ,
         \i_MIPS/Register/register[9][7] , \i_MIPS/Register/register[9][8] ,
         \i_MIPS/Register/register[9][9] , \i_MIPS/Register/register[9][10] ,
         \i_MIPS/Register/register[9][11] , \i_MIPS/Register/register[9][12] ,
         \i_MIPS/Register/register[9][13] , \i_MIPS/Register/register[9][14] ,
         \i_MIPS/Register/register[9][15] , \i_MIPS/Register/register[9][16] ,
         \i_MIPS/Register/register[9][17] , \i_MIPS/Register/register[9][18] ,
         \i_MIPS/Register/register[9][19] , \i_MIPS/Register/register[9][20] ,
         \i_MIPS/Register/register[9][21] , \i_MIPS/Register/register[9][22] ,
         \i_MIPS/Register/register[9][23] , \i_MIPS/Register/register[9][24] ,
         \i_MIPS/Register/register[9][25] , \i_MIPS/Register/register[9][26] ,
         \i_MIPS/Register/register[9][27] , \i_MIPS/Register/register[9][28] ,
         \i_MIPS/Register/register[9][29] , \i_MIPS/Register/register[9][30] ,
         \i_MIPS/Register/register[9][31] , \i_MIPS/Register/register[8][0] ,
         \i_MIPS/Register/register[8][1] , \i_MIPS/Register/register[8][2] ,
         \i_MIPS/Register/register[8][3] , \i_MIPS/Register/register[8][4] ,
         \i_MIPS/Register/register[8][5] , \i_MIPS/Register/register[8][6] ,
         \i_MIPS/Register/register[8][7] , \i_MIPS/Register/register[8][8] ,
         \i_MIPS/Register/register[8][9] , \i_MIPS/Register/register[8][10] ,
         \i_MIPS/Register/register[8][11] , \i_MIPS/Register/register[8][12] ,
         \i_MIPS/Register/register[8][13] , \i_MIPS/Register/register[8][14] ,
         \i_MIPS/Register/register[8][15] , \i_MIPS/Register/register[8][16] ,
         \i_MIPS/Register/register[8][17] , \i_MIPS/Register/register[8][18] ,
         \i_MIPS/Register/register[8][19] , \i_MIPS/Register/register[8][20] ,
         \i_MIPS/Register/register[8][21] , \i_MIPS/Register/register[8][22] ,
         \i_MIPS/Register/register[8][23] , \i_MIPS/Register/register[8][24] ,
         \i_MIPS/Register/register[8][25] , \i_MIPS/Register/register[8][26] ,
         \i_MIPS/Register/register[8][27] , \i_MIPS/Register/register[8][28] ,
         \i_MIPS/Register/register[8][29] , \i_MIPS/Register/register[8][30] ,
         \i_MIPS/Register/register[8][31] , \i_MIPS/Register/register[7][0] ,
         \i_MIPS/Register/register[7][1] , \i_MIPS/Register/register[7][2] ,
         \i_MIPS/Register/register[7][3] , \i_MIPS/Register/register[7][4] ,
         \i_MIPS/Register/register[7][5] , \i_MIPS/Register/register[7][6] ,
         \i_MIPS/Register/register[7][7] , \i_MIPS/Register/register[7][8] ,
         \i_MIPS/Register/register[7][9] , \i_MIPS/Register/register[7][10] ,
         \i_MIPS/Register/register[7][11] , \i_MIPS/Register/register[7][12] ,
         \i_MIPS/Register/register[7][13] , \i_MIPS/Register/register[7][14] ,
         \i_MIPS/Register/register[7][15] , \i_MIPS/Register/register[7][16] ,
         \i_MIPS/Register/register[7][17] , \i_MIPS/Register/register[7][18] ,
         \i_MIPS/Register/register[7][19] , \i_MIPS/Register/register[7][20] ,
         \i_MIPS/Register/register[7][21] , \i_MIPS/Register/register[7][22] ,
         \i_MIPS/Register/register[7][23] , \i_MIPS/Register/register[7][24] ,
         \i_MIPS/Register/register[7][25] , \i_MIPS/Register/register[7][26] ,
         \i_MIPS/Register/register[7][27] , \i_MIPS/Register/register[7][28] ,
         \i_MIPS/Register/register[7][29] , \i_MIPS/Register/register[7][30] ,
         \i_MIPS/Register/register[7][31] , \i_MIPS/Register/register[6][0] ,
         \i_MIPS/Register/register[6][1] , \i_MIPS/Register/register[6][2] ,
         \i_MIPS/Register/register[6][3] , \i_MIPS/Register/register[6][4] ,
         \i_MIPS/Register/register[6][5] , \i_MIPS/Register/register[6][6] ,
         \i_MIPS/Register/register[6][7] , \i_MIPS/Register/register[6][8] ,
         \i_MIPS/Register/register[6][9] , \i_MIPS/Register/register[6][10] ,
         \i_MIPS/Register/register[6][11] , \i_MIPS/Register/register[6][12] ,
         \i_MIPS/Register/register[6][13] , \i_MIPS/Register/register[6][14] ,
         \i_MIPS/Register/register[6][15] , \i_MIPS/Register/register[6][16] ,
         \i_MIPS/Register/register[6][17] , \i_MIPS/Register/register[6][18] ,
         \i_MIPS/Register/register[6][19] , \i_MIPS/Register/register[6][20] ,
         \i_MIPS/Register/register[6][21] , \i_MIPS/Register/register[6][22] ,
         \i_MIPS/Register/register[6][23] , \i_MIPS/Register/register[6][24] ,
         \i_MIPS/Register/register[6][25] , \i_MIPS/Register/register[6][26] ,
         \i_MIPS/Register/register[6][27] , \i_MIPS/Register/register[6][28] ,
         \i_MIPS/Register/register[6][29] , \i_MIPS/Register/register[6][30] ,
         \i_MIPS/Register/register[6][31] , \i_MIPS/Register/register[5][0] ,
         \i_MIPS/Register/register[5][1] , \i_MIPS/Register/register[5][2] ,
         \i_MIPS/Register/register[5][3] , \i_MIPS/Register/register[5][4] ,
         \i_MIPS/Register/register[5][5] , \i_MIPS/Register/register[5][6] ,
         \i_MIPS/Register/register[5][7] , \i_MIPS/Register/register[5][8] ,
         \i_MIPS/Register/register[5][9] , \i_MIPS/Register/register[5][10] ,
         \i_MIPS/Register/register[5][11] , \i_MIPS/Register/register[5][12] ,
         \i_MIPS/Register/register[5][13] , \i_MIPS/Register/register[5][14] ,
         \i_MIPS/Register/register[5][15] , \i_MIPS/Register/register[5][16] ,
         \i_MIPS/Register/register[5][17] , \i_MIPS/Register/register[5][18] ,
         \i_MIPS/Register/register[5][19] , \i_MIPS/Register/register[5][20] ,
         \i_MIPS/Register/register[5][21] , \i_MIPS/Register/register[5][22] ,
         \i_MIPS/Register/register[5][23] , \i_MIPS/Register/register[5][24] ,
         \i_MIPS/Register/register[5][25] , \i_MIPS/Register/register[5][26] ,
         \i_MIPS/Register/register[5][27] , \i_MIPS/Register/register[5][28] ,
         \i_MIPS/Register/register[5][29] , \i_MIPS/Register/register[5][30] ,
         \i_MIPS/Register/register[5][31] , \i_MIPS/Register/register[4][0] ,
         \i_MIPS/Register/register[4][1] , \i_MIPS/Register/register[4][2] ,
         \i_MIPS/Register/register[4][3] , \i_MIPS/Register/register[4][4] ,
         \i_MIPS/Register/register[4][5] , \i_MIPS/Register/register[4][6] ,
         \i_MIPS/Register/register[4][7] , \i_MIPS/Register/register[4][8] ,
         \i_MIPS/Register/register[4][9] , \i_MIPS/Register/register[4][10] ,
         \i_MIPS/Register/register[4][11] , \i_MIPS/Register/register[4][12] ,
         \i_MIPS/Register/register[4][13] , \i_MIPS/Register/register[4][14] ,
         \i_MIPS/Register/register[4][15] , \i_MIPS/Register/register[4][16] ,
         \i_MIPS/Register/register[4][17] , \i_MIPS/Register/register[4][18] ,
         \i_MIPS/Register/register[4][19] , \i_MIPS/Register/register[4][20] ,
         \i_MIPS/Register/register[4][21] , \i_MIPS/Register/register[4][22] ,
         \i_MIPS/Register/register[4][23] , \i_MIPS/Register/register[4][24] ,
         \i_MIPS/Register/register[4][25] , \i_MIPS/Register/register[4][26] ,
         \i_MIPS/Register/register[4][27] , \i_MIPS/Register/register[4][28] ,
         \i_MIPS/Register/register[4][29] , \i_MIPS/Register/register[4][30] ,
         \i_MIPS/Register/register[4][31] , \i_MIPS/Register/register[3][0] ,
         \i_MIPS/Register/register[3][1] , \i_MIPS/Register/register[3][2] ,
         \i_MIPS/Register/register[3][3] , \i_MIPS/Register/register[3][4] ,
         \i_MIPS/Register/register[3][5] , \i_MIPS/Register/register[3][6] ,
         \i_MIPS/Register/register[3][7] , \i_MIPS/Register/register[3][8] ,
         \i_MIPS/Register/register[3][9] , \i_MIPS/Register/register[3][10] ,
         \i_MIPS/Register/register[3][11] , \i_MIPS/Register/register[3][12] ,
         \i_MIPS/Register/register[3][13] , \i_MIPS/Register/register[3][14] ,
         \i_MIPS/Register/register[3][15] , \i_MIPS/Register/register[3][16] ,
         \i_MIPS/Register/register[3][17] , \i_MIPS/Register/register[3][18] ,
         \i_MIPS/Register/register[3][19] , \i_MIPS/Register/register[3][20] ,
         \i_MIPS/Register/register[3][21] , \i_MIPS/Register/register[3][22] ,
         \i_MIPS/Register/register[3][23] , \i_MIPS/Register/register[3][24] ,
         \i_MIPS/Register/register[3][25] , \i_MIPS/Register/register[3][26] ,
         \i_MIPS/Register/register[3][27] , \i_MIPS/Register/register[3][28] ,
         \i_MIPS/Register/register[3][29] , \i_MIPS/Register/register[3][30] ,
         \i_MIPS/Register/register[3][31] , \i_MIPS/Register/register[2][0] ,
         \i_MIPS/Register/register[2][1] , \i_MIPS/Register/register[2][2] ,
         \i_MIPS/Register/register[2][3] , \i_MIPS/Register/register[2][4] ,
         \i_MIPS/Register/register[2][5] , \i_MIPS/Register/register[2][6] ,
         \i_MIPS/Register/register[2][7] , \i_MIPS/Register/register[2][8] ,
         \i_MIPS/Register/register[2][9] , \i_MIPS/Register/register[2][10] ,
         \i_MIPS/Register/register[2][11] , \i_MIPS/Register/register[2][12] ,
         \i_MIPS/Register/register[2][13] , \i_MIPS/Register/register[2][14] ,
         \i_MIPS/Register/register[2][15] , \i_MIPS/Register/register[2][16] ,
         \i_MIPS/Register/register[2][17] , \i_MIPS/Register/register[2][18] ,
         \i_MIPS/Register/register[2][19] , \i_MIPS/Register/register[2][20] ,
         \i_MIPS/Register/register[2][21] , \i_MIPS/Register/register[2][22] ,
         \i_MIPS/Register/register[2][23] , \i_MIPS/Register/register[2][24] ,
         \i_MIPS/Register/register[2][25] , \i_MIPS/Register/register[2][26] ,
         \i_MIPS/Register/register[2][27] , \i_MIPS/Register/register[2][28] ,
         \i_MIPS/Register/register[2][29] , \i_MIPS/Register/register[2][30] ,
         \i_MIPS/Register/register[2][31] , \i_MIPS/Register/register[1][0] ,
         \i_MIPS/Register/register[1][1] , \i_MIPS/Register/register[1][2] ,
         \i_MIPS/Register/register[1][3] , \i_MIPS/Register/register[1][4] ,
         \i_MIPS/Register/register[1][5] , \i_MIPS/Register/register[1][6] ,
         \i_MIPS/Register/register[1][7] , \i_MIPS/Register/register[1][8] ,
         \i_MIPS/Register/register[1][9] , \i_MIPS/Register/register[1][10] ,
         \i_MIPS/Register/register[1][11] , \i_MIPS/Register/register[1][12] ,
         \i_MIPS/Register/register[1][13] , \i_MIPS/Register/register[1][14] ,
         \i_MIPS/Register/register[1][15] , \i_MIPS/Register/register[1][16] ,
         \i_MIPS/Register/register[1][17] , \i_MIPS/Register/register[1][18] ,
         \i_MIPS/Register/register[1][19] , \i_MIPS/Register/register[1][20] ,
         \i_MIPS/Register/register[1][21] , \i_MIPS/Register/register[1][22] ,
         \i_MIPS/Register/register[1][23] , \i_MIPS/Register/register[1][24] ,
         \i_MIPS/Register/register[1][25] , \i_MIPS/Register/register[1][26] ,
         \i_MIPS/Register/register[1][27] , \i_MIPS/Register/register[1][28] ,
         \i_MIPS/Register/register[1][29] , \i_MIPS/Register/register[1][30] ,
         \i_MIPS/Register/register[1][31] , \i_MIPS/Register/register[0][0] ,
         \i_MIPS/Register/register[0][1] , \i_MIPS/Register/register[0][2] ,
         \i_MIPS/Register/register[0][3] , \i_MIPS/Register/register[0][4] ,
         \i_MIPS/Register/register[0][5] , \i_MIPS/Register/register[0][6] ,
         \i_MIPS/Register/register[0][7] , \i_MIPS/Register/register[0][8] ,
         \i_MIPS/Register/register[0][9] , \i_MIPS/Register/register[0][10] ,
         \i_MIPS/Register/register[0][11] , \i_MIPS/Register/register[0][12] ,
         \i_MIPS/Register/register[0][13] , \i_MIPS/Register/register[0][14] ,
         \i_MIPS/Register/register[0][15] , \i_MIPS/Register/register[0][16] ,
         \i_MIPS/Register/register[0][17] , \i_MIPS/Register/register[0][18] ,
         \i_MIPS/Register/register[0][19] , \i_MIPS/Register/register[0][20] ,
         \i_MIPS/Register/register[0][21] , \i_MIPS/Register/register[0][22] ,
         \i_MIPS/Register/register[0][23] , \i_MIPS/Register/register[0][24] ,
         \i_MIPS/Register/register[0][25] , \i_MIPS/Register/register[0][26] ,
         \i_MIPS/Register/register[0][27] , \i_MIPS/Register/register[0][28] ,
         \i_MIPS/Register/register[0][29] , \i_MIPS/Register/register[0][30] ,
         \i_MIPS/Register/register[0][31] , \i_MIPS/Control_ID/n15 ,
         \i_MIPS/Control_ID/n12 , \i_MIPS/Control_ID/n10 ,
         \i_MIPS/Hazard_detection/n13 , \i_MIPS/Hazard_detection/n12 ,
         \i_MIPS/Hazard_detection/n11 , \i_MIPS/Hazard_detection/n10 ,
         \i_MIPS/Hazard_detection/n9 , \i_MIPS/Hazard_detection/n8 ,
         \i_MIPS/Hazard_detection/n7 , \i_MIPS/Hazard_detection/n4 ,
         \i_MIPS/forward_unit/n25 , \i_MIPS/forward_unit/n10 ,
         \i_MIPS/ALU_Control/n20 , \i_MIPS/ALU_Control/n18 ,
         \i_MIPS/ALU_Control/n11 , \i_MIPS/ALU/N303 , \I_cache/cache[7][0] ,
         \I_cache/cache[7][1] , \I_cache/cache[7][2] , \I_cache/cache[7][3] ,
         \I_cache/cache[7][4] , \I_cache/cache[7][5] , \I_cache/cache[7][6] ,
         \I_cache/cache[7][7] , \I_cache/cache[7][8] , \I_cache/cache[7][9] ,
         \I_cache/cache[7][10] , \I_cache/cache[7][11] ,
         \I_cache/cache[7][12] , \I_cache/cache[7][13] ,
         \I_cache/cache[7][14] , \I_cache/cache[7][15] ,
         \I_cache/cache[7][16] , \I_cache/cache[7][17] ,
         \I_cache/cache[7][18] , \I_cache/cache[7][19] ,
         \I_cache/cache[7][20] , \I_cache/cache[7][21] ,
         \I_cache/cache[7][22] , \I_cache/cache[7][23] ,
         \I_cache/cache[7][24] , \I_cache/cache[7][25] ,
         \I_cache/cache[7][26] , \I_cache/cache[7][27] ,
         \I_cache/cache[7][28] , \I_cache/cache[7][29] ,
         \I_cache/cache[7][30] , \I_cache/cache[7][31] ,
         \I_cache/cache[7][32] , \I_cache/cache[7][33] ,
         \I_cache/cache[7][34] , \I_cache/cache[7][35] ,
         \I_cache/cache[7][36] , \I_cache/cache[7][37] ,
         \I_cache/cache[7][38] , \I_cache/cache[7][39] ,
         \I_cache/cache[7][40] , \I_cache/cache[7][41] ,
         \I_cache/cache[7][42] , \I_cache/cache[7][43] ,
         \I_cache/cache[7][44] , \I_cache/cache[7][45] ,
         \I_cache/cache[7][46] , \I_cache/cache[7][47] ,
         \I_cache/cache[7][48] , \I_cache/cache[7][49] ,
         \I_cache/cache[7][50] , \I_cache/cache[7][51] ,
         \I_cache/cache[7][52] , \I_cache/cache[7][53] ,
         \I_cache/cache[7][54] , \I_cache/cache[7][55] ,
         \I_cache/cache[7][56] , \I_cache/cache[7][57] ,
         \I_cache/cache[7][58] , \I_cache/cache[7][59] ,
         \I_cache/cache[7][60] , \I_cache/cache[7][61] ,
         \I_cache/cache[7][62] , \I_cache/cache[7][63] ,
         \I_cache/cache[7][64] , \I_cache/cache[7][65] ,
         \I_cache/cache[7][66] , \I_cache/cache[7][67] ,
         \I_cache/cache[7][68] , \I_cache/cache[7][69] ,
         \I_cache/cache[7][70] , \I_cache/cache[7][71] ,
         \I_cache/cache[7][72] , \I_cache/cache[7][73] ,
         \I_cache/cache[7][74] , \I_cache/cache[7][75] ,
         \I_cache/cache[7][76] , \I_cache/cache[7][77] ,
         \I_cache/cache[7][78] , \I_cache/cache[7][79] ,
         \I_cache/cache[7][80] , \I_cache/cache[7][81] ,
         \I_cache/cache[7][82] , \I_cache/cache[7][83] ,
         \I_cache/cache[7][84] , \I_cache/cache[7][85] ,
         \I_cache/cache[7][86] , \I_cache/cache[7][87] ,
         \I_cache/cache[7][88] , \I_cache/cache[7][89] ,
         \I_cache/cache[7][90] , \I_cache/cache[7][91] ,
         \I_cache/cache[7][92] , \I_cache/cache[7][93] ,
         \I_cache/cache[7][94] , \I_cache/cache[7][95] ,
         \I_cache/cache[7][96] , \I_cache/cache[7][97] ,
         \I_cache/cache[7][98] , \I_cache/cache[7][99] ,
         \I_cache/cache[7][100] , \I_cache/cache[7][101] ,
         \I_cache/cache[7][102] , \I_cache/cache[7][103] ,
         \I_cache/cache[7][104] , \I_cache/cache[7][105] ,
         \I_cache/cache[7][106] , \I_cache/cache[7][107] ,
         \I_cache/cache[7][108] , \I_cache/cache[7][109] ,
         \I_cache/cache[7][110] , \I_cache/cache[7][111] ,
         \I_cache/cache[7][112] , \I_cache/cache[7][113] ,
         \I_cache/cache[7][114] , \I_cache/cache[7][115] ,
         \I_cache/cache[7][116] , \I_cache/cache[7][117] ,
         \I_cache/cache[7][118] , \I_cache/cache[7][119] ,
         \I_cache/cache[7][120] , \I_cache/cache[7][121] ,
         \I_cache/cache[7][122] , \I_cache/cache[7][123] ,
         \I_cache/cache[7][124] , \I_cache/cache[7][125] ,
         \I_cache/cache[7][126] , \I_cache/cache[7][127] ,
         \I_cache/cache[7][128] , \I_cache/cache[7][129] ,
         \I_cache/cache[7][130] , \I_cache/cache[7][131] ,
         \I_cache/cache[7][132] , \I_cache/cache[7][133] ,
         \I_cache/cache[7][134] , \I_cache/cache[7][135] ,
         \I_cache/cache[7][136] , \I_cache/cache[7][137] ,
         \I_cache/cache[7][138] , \I_cache/cache[7][139] ,
         \I_cache/cache[7][140] , \I_cache/cache[7][141] ,
         \I_cache/cache[7][142] , \I_cache/cache[7][143] ,
         \I_cache/cache[7][144] , \I_cache/cache[7][145] ,
         \I_cache/cache[7][146] , \I_cache/cache[7][147] ,
         \I_cache/cache[7][148] , \I_cache/cache[7][149] ,
         \I_cache/cache[7][150] , \I_cache/cache[7][151] ,
         \I_cache/cache[7][152] , \I_cache/cache[7][153] ,
         \I_cache/cache[7][154] , \I_cache/cache[6][0] , \I_cache/cache[6][1] ,
         \I_cache/cache[6][2] , \I_cache/cache[6][3] , \I_cache/cache[6][4] ,
         \I_cache/cache[6][5] , \I_cache/cache[6][6] , \I_cache/cache[6][7] ,
         \I_cache/cache[6][8] , \I_cache/cache[6][9] , \I_cache/cache[6][10] ,
         \I_cache/cache[6][11] , \I_cache/cache[6][12] ,
         \I_cache/cache[6][13] , \I_cache/cache[6][14] ,
         \I_cache/cache[6][15] , \I_cache/cache[6][16] ,
         \I_cache/cache[6][17] , \I_cache/cache[6][18] ,
         \I_cache/cache[6][19] , \I_cache/cache[6][20] ,
         \I_cache/cache[6][21] , \I_cache/cache[6][22] ,
         \I_cache/cache[6][23] , \I_cache/cache[6][24] ,
         \I_cache/cache[6][25] , \I_cache/cache[6][26] ,
         \I_cache/cache[6][27] , \I_cache/cache[6][28] ,
         \I_cache/cache[6][29] , \I_cache/cache[6][30] ,
         \I_cache/cache[6][31] , \I_cache/cache[6][32] ,
         \I_cache/cache[6][33] , \I_cache/cache[6][34] ,
         \I_cache/cache[6][35] , \I_cache/cache[6][36] ,
         \I_cache/cache[6][37] , \I_cache/cache[6][38] ,
         \I_cache/cache[6][39] , \I_cache/cache[6][40] ,
         \I_cache/cache[6][41] , \I_cache/cache[6][42] ,
         \I_cache/cache[6][43] , \I_cache/cache[6][44] ,
         \I_cache/cache[6][45] , \I_cache/cache[6][46] ,
         \I_cache/cache[6][47] , \I_cache/cache[6][48] ,
         \I_cache/cache[6][49] , \I_cache/cache[6][50] ,
         \I_cache/cache[6][51] , \I_cache/cache[6][52] ,
         \I_cache/cache[6][53] , \I_cache/cache[6][54] ,
         \I_cache/cache[6][55] , \I_cache/cache[6][56] ,
         \I_cache/cache[6][57] , \I_cache/cache[6][58] ,
         \I_cache/cache[6][59] , \I_cache/cache[6][60] ,
         \I_cache/cache[6][61] , \I_cache/cache[6][62] ,
         \I_cache/cache[6][63] , \I_cache/cache[6][64] ,
         \I_cache/cache[6][65] , \I_cache/cache[6][66] ,
         \I_cache/cache[6][67] , \I_cache/cache[6][68] ,
         \I_cache/cache[6][69] , \I_cache/cache[6][70] ,
         \I_cache/cache[6][71] , \I_cache/cache[6][72] ,
         \I_cache/cache[6][73] , \I_cache/cache[6][74] ,
         \I_cache/cache[6][75] , \I_cache/cache[6][76] ,
         \I_cache/cache[6][77] , \I_cache/cache[6][78] ,
         \I_cache/cache[6][79] , \I_cache/cache[6][80] ,
         \I_cache/cache[6][81] , \I_cache/cache[6][82] ,
         \I_cache/cache[6][83] , \I_cache/cache[6][84] ,
         \I_cache/cache[6][85] , \I_cache/cache[6][86] ,
         \I_cache/cache[6][87] , \I_cache/cache[6][88] ,
         \I_cache/cache[6][89] , \I_cache/cache[6][90] ,
         \I_cache/cache[6][91] , \I_cache/cache[6][92] ,
         \I_cache/cache[6][93] , \I_cache/cache[6][94] ,
         \I_cache/cache[6][95] , \I_cache/cache[6][96] ,
         \I_cache/cache[6][97] , \I_cache/cache[6][98] ,
         \I_cache/cache[6][99] , \I_cache/cache[6][100] ,
         \I_cache/cache[6][101] , \I_cache/cache[6][102] ,
         \I_cache/cache[6][103] , \I_cache/cache[6][104] ,
         \I_cache/cache[6][105] , \I_cache/cache[6][106] ,
         \I_cache/cache[6][107] , \I_cache/cache[6][108] ,
         \I_cache/cache[6][109] , \I_cache/cache[6][110] ,
         \I_cache/cache[6][111] , \I_cache/cache[6][112] ,
         \I_cache/cache[6][113] , \I_cache/cache[6][114] ,
         \I_cache/cache[6][115] , \I_cache/cache[6][116] ,
         \I_cache/cache[6][117] , \I_cache/cache[6][118] ,
         \I_cache/cache[6][119] , \I_cache/cache[6][120] ,
         \I_cache/cache[6][121] , \I_cache/cache[6][122] ,
         \I_cache/cache[6][123] , \I_cache/cache[6][124] ,
         \I_cache/cache[6][125] , \I_cache/cache[6][126] ,
         \I_cache/cache[6][127] , \I_cache/cache[6][128] ,
         \I_cache/cache[6][129] , \I_cache/cache[6][130] ,
         \I_cache/cache[6][131] , \I_cache/cache[6][132] ,
         \I_cache/cache[6][133] , \I_cache/cache[6][134] ,
         \I_cache/cache[6][135] , \I_cache/cache[6][136] ,
         \I_cache/cache[6][137] , \I_cache/cache[6][138] ,
         \I_cache/cache[6][139] , \I_cache/cache[6][140] ,
         \I_cache/cache[6][141] , \I_cache/cache[6][142] ,
         \I_cache/cache[6][143] , \I_cache/cache[6][144] ,
         \I_cache/cache[6][145] , \I_cache/cache[6][146] ,
         \I_cache/cache[6][147] , \I_cache/cache[6][148] ,
         \I_cache/cache[6][149] , \I_cache/cache[6][150] ,
         \I_cache/cache[6][151] , \I_cache/cache[6][152] ,
         \I_cache/cache[6][153] , \I_cache/cache[6][154] ,
         \I_cache/cache[5][0] , \I_cache/cache[5][1] , \I_cache/cache[5][2] ,
         \I_cache/cache[5][3] , \I_cache/cache[5][4] , \I_cache/cache[5][5] ,
         \I_cache/cache[5][6] , \I_cache/cache[5][7] , \I_cache/cache[5][8] ,
         \I_cache/cache[5][9] , \I_cache/cache[5][10] , \I_cache/cache[5][11] ,
         \I_cache/cache[5][12] , \I_cache/cache[5][13] ,
         \I_cache/cache[5][14] , \I_cache/cache[5][15] ,
         \I_cache/cache[5][16] , \I_cache/cache[5][17] ,
         \I_cache/cache[5][18] , \I_cache/cache[5][19] ,
         \I_cache/cache[5][20] , \I_cache/cache[5][21] ,
         \I_cache/cache[5][22] , \I_cache/cache[5][23] ,
         \I_cache/cache[5][24] , \I_cache/cache[5][25] ,
         \I_cache/cache[5][26] , \I_cache/cache[5][27] ,
         \I_cache/cache[5][28] , \I_cache/cache[5][29] ,
         \I_cache/cache[5][30] , \I_cache/cache[5][31] ,
         \I_cache/cache[5][32] , \I_cache/cache[5][33] ,
         \I_cache/cache[5][34] , \I_cache/cache[5][35] ,
         \I_cache/cache[5][36] , \I_cache/cache[5][37] ,
         \I_cache/cache[5][38] , \I_cache/cache[5][39] ,
         \I_cache/cache[5][40] , \I_cache/cache[5][41] ,
         \I_cache/cache[5][42] , \I_cache/cache[5][43] ,
         \I_cache/cache[5][44] , \I_cache/cache[5][45] ,
         \I_cache/cache[5][46] , \I_cache/cache[5][47] ,
         \I_cache/cache[5][48] , \I_cache/cache[5][49] ,
         \I_cache/cache[5][50] , \I_cache/cache[5][51] ,
         \I_cache/cache[5][52] , \I_cache/cache[5][53] ,
         \I_cache/cache[5][54] , \I_cache/cache[5][55] ,
         \I_cache/cache[5][56] , \I_cache/cache[5][57] ,
         \I_cache/cache[5][58] , \I_cache/cache[5][59] ,
         \I_cache/cache[5][60] , \I_cache/cache[5][61] ,
         \I_cache/cache[5][62] , \I_cache/cache[5][63] ,
         \I_cache/cache[5][64] , \I_cache/cache[5][65] ,
         \I_cache/cache[5][66] , \I_cache/cache[5][67] ,
         \I_cache/cache[5][68] , \I_cache/cache[5][69] ,
         \I_cache/cache[5][70] , \I_cache/cache[5][71] ,
         \I_cache/cache[5][72] , \I_cache/cache[5][73] ,
         \I_cache/cache[5][74] , \I_cache/cache[5][75] ,
         \I_cache/cache[5][76] , \I_cache/cache[5][77] ,
         \I_cache/cache[5][78] , \I_cache/cache[5][79] ,
         \I_cache/cache[5][80] , \I_cache/cache[5][81] ,
         \I_cache/cache[5][82] , \I_cache/cache[5][83] ,
         \I_cache/cache[5][84] , \I_cache/cache[5][85] ,
         \I_cache/cache[5][86] , \I_cache/cache[5][87] ,
         \I_cache/cache[5][88] , \I_cache/cache[5][89] ,
         \I_cache/cache[5][90] , \I_cache/cache[5][91] ,
         \I_cache/cache[5][92] , \I_cache/cache[5][93] ,
         \I_cache/cache[5][94] , \I_cache/cache[5][95] ,
         \I_cache/cache[5][96] , \I_cache/cache[5][97] ,
         \I_cache/cache[5][98] , \I_cache/cache[5][99] ,
         \I_cache/cache[5][100] , \I_cache/cache[5][101] ,
         \I_cache/cache[5][102] , \I_cache/cache[5][103] ,
         \I_cache/cache[5][104] , \I_cache/cache[5][105] ,
         \I_cache/cache[5][106] , \I_cache/cache[5][107] ,
         \I_cache/cache[5][108] , \I_cache/cache[5][109] ,
         \I_cache/cache[5][110] , \I_cache/cache[5][111] ,
         \I_cache/cache[5][112] , \I_cache/cache[5][113] ,
         \I_cache/cache[5][114] , \I_cache/cache[5][115] ,
         \I_cache/cache[5][116] , \I_cache/cache[5][117] ,
         \I_cache/cache[5][118] , \I_cache/cache[5][119] ,
         \I_cache/cache[5][120] , \I_cache/cache[5][121] ,
         \I_cache/cache[5][122] , \I_cache/cache[5][123] ,
         \I_cache/cache[5][124] , \I_cache/cache[5][125] ,
         \I_cache/cache[5][126] , \I_cache/cache[5][127] ,
         \I_cache/cache[5][128] , \I_cache/cache[5][129] ,
         \I_cache/cache[5][130] , \I_cache/cache[5][131] ,
         \I_cache/cache[5][132] , \I_cache/cache[5][133] ,
         \I_cache/cache[5][134] , \I_cache/cache[5][135] ,
         \I_cache/cache[5][136] , \I_cache/cache[5][137] ,
         \I_cache/cache[5][138] , \I_cache/cache[5][139] ,
         \I_cache/cache[5][140] , \I_cache/cache[5][141] ,
         \I_cache/cache[5][142] , \I_cache/cache[5][143] ,
         \I_cache/cache[5][144] , \I_cache/cache[5][145] ,
         \I_cache/cache[5][146] , \I_cache/cache[5][147] ,
         \I_cache/cache[5][148] , \I_cache/cache[5][149] ,
         \I_cache/cache[5][150] , \I_cache/cache[5][151] ,
         \I_cache/cache[5][152] , \I_cache/cache[5][153] ,
         \I_cache/cache[5][154] , \I_cache/cache[4][0] , \I_cache/cache[4][1] ,
         \I_cache/cache[4][2] , \I_cache/cache[4][3] , \I_cache/cache[4][4] ,
         \I_cache/cache[4][5] , \I_cache/cache[4][6] , \I_cache/cache[4][7] ,
         \I_cache/cache[4][8] , \I_cache/cache[4][9] , \I_cache/cache[4][10] ,
         \I_cache/cache[4][11] , \I_cache/cache[4][12] ,
         \I_cache/cache[4][13] , \I_cache/cache[4][14] ,
         \I_cache/cache[4][15] , \I_cache/cache[4][16] ,
         \I_cache/cache[4][17] , \I_cache/cache[4][18] ,
         \I_cache/cache[4][19] , \I_cache/cache[4][20] ,
         \I_cache/cache[4][21] , \I_cache/cache[4][22] ,
         \I_cache/cache[4][23] , \I_cache/cache[4][24] ,
         \I_cache/cache[4][25] , \I_cache/cache[4][26] ,
         \I_cache/cache[4][27] , \I_cache/cache[4][28] ,
         \I_cache/cache[4][29] , \I_cache/cache[4][30] ,
         \I_cache/cache[4][31] , \I_cache/cache[4][32] ,
         \I_cache/cache[4][33] , \I_cache/cache[4][34] ,
         \I_cache/cache[4][35] , \I_cache/cache[4][36] ,
         \I_cache/cache[4][37] , \I_cache/cache[4][38] ,
         \I_cache/cache[4][39] , \I_cache/cache[4][40] ,
         \I_cache/cache[4][41] , \I_cache/cache[4][42] ,
         \I_cache/cache[4][43] , \I_cache/cache[4][44] ,
         \I_cache/cache[4][45] , \I_cache/cache[4][46] ,
         \I_cache/cache[4][47] , \I_cache/cache[4][48] ,
         \I_cache/cache[4][49] , \I_cache/cache[4][50] ,
         \I_cache/cache[4][51] , \I_cache/cache[4][52] ,
         \I_cache/cache[4][53] , \I_cache/cache[4][54] ,
         \I_cache/cache[4][55] , \I_cache/cache[4][56] ,
         \I_cache/cache[4][57] , \I_cache/cache[4][58] ,
         \I_cache/cache[4][59] , \I_cache/cache[4][60] ,
         \I_cache/cache[4][61] , \I_cache/cache[4][62] ,
         \I_cache/cache[4][63] , \I_cache/cache[4][64] ,
         \I_cache/cache[4][65] , \I_cache/cache[4][66] ,
         \I_cache/cache[4][67] , \I_cache/cache[4][68] ,
         \I_cache/cache[4][69] , \I_cache/cache[4][70] ,
         \I_cache/cache[4][71] , \I_cache/cache[4][72] ,
         \I_cache/cache[4][73] , \I_cache/cache[4][74] ,
         \I_cache/cache[4][75] , \I_cache/cache[4][76] ,
         \I_cache/cache[4][77] , \I_cache/cache[4][78] ,
         \I_cache/cache[4][79] , \I_cache/cache[4][80] ,
         \I_cache/cache[4][81] , \I_cache/cache[4][82] ,
         \I_cache/cache[4][83] , \I_cache/cache[4][84] ,
         \I_cache/cache[4][85] , \I_cache/cache[4][86] ,
         \I_cache/cache[4][87] , \I_cache/cache[4][88] ,
         \I_cache/cache[4][89] , \I_cache/cache[4][90] ,
         \I_cache/cache[4][91] , \I_cache/cache[4][92] ,
         \I_cache/cache[4][93] , \I_cache/cache[4][94] ,
         \I_cache/cache[4][95] , \I_cache/cache[4][96] ,
         \I_cache/cache[4][97] , \I_cache/cache[4][98] ,
         \I_cache/cache[4][99] , \I_cache/cache[4][100] ,
         \I_cache/cache[4][101] , \I_cache/cache[4][102] ,
         \I_cache/cache[4][103] , \I_cache/cache[4][104] ,
         \I_cache/cache[4][105] , \I_cache/cache[4][106] ,
         \I_cache/cache[4][107] , \I_cache/cache[4][108] ,
         \I_cache/cache[4][109] , \I_cache/cache[4][110] ,
         \I_cache/cache[4][111] , \I_cache/cache[4][112] ,
         \I_cache/cache[4][113] , \I_cache/cache[4][114] ,
         \I_cache/cache[4][115] , \I_cache/cache[4][116] ,
         \I_cache/cache[4][117] , \I_cache/cache[4][118] ,
         \I_cache/cache[4][119] , \I_cache/cache[4][120] ,
         \I_cache/cache[4][121] , \I_cache/cache[4][122] ,
         \I_cache/cache[4][123] , \I_cache/cache[4][124] ,
         \I_cache/cache[4][125] , \I_cache/cache[4][126] ,
         \I_cache/cache[4][127] , \I_cache/cache[4][128] ,
         \I_cache/cache[4][129] , \I_cache/cache[4][130] ,
         \I_cache/cache[4][131] , \I_cache/cache[4][132] ,
         \I_cache/cache[4][133] , \I_cache/cache[4][134] ,
         \I_cache/cache[4][135] , \I_cache/cache[4][136] ,
         \I_cache/cache[4][137] , \I_cache/cache[4][138] ,
         \I_cache/cache[4][139] , \I_cache/cache[4][140] ,
         \I_cache/cache[4][141] , \I_cache/cache[4][142] ,
         \I_cache/cache[4][143] , \I_cache/cache[4][144] ,
         \I_cache/cache[4][145] , \I_cache/cache[4][146] ,
         \I_cache/cache[4][147] , \I_cache/cache[4][148] ,
         \I_cache/cache[4][149] , \I_cache/cache[4][150] ,
         \I_cache/cache[4][151] , \I_cache/cache[4][152] ,
         \I_cache/cache[4][153] , \I_cache/cache[4][154] ,
         \I_cache/cache[3][0] , \I_cache/cache[3][1] , \I_cache/cache[3][2] ,
         \I_cache/cache[3][3] , \I_cache/cache[3][4] , \I_cache/cache[3][5] ,
         \I_cache/cache[3][6] , \I_cache/cache[3][7] , \I_cache/cache[3][8] ,
         \I_cache/cache[3][9] , \I_cache/cache[3][10] , \I_cache/cache[3][11] ,
         \I_cache/cache[3][12] , \I_cache/cache[3][13] ,
         \I_cache/cache[3][14] , \I_cache/cache[3][15] ,
         \I_cache/cache[3][16] , \I_cache/cache[3][17] ,
         \I_cache/cache[3][18] , \I_cache/cache[3][19] ,
         \I_cache/cache[3][20] , \I_cache/cache[3][21] ,
         \I_cache/cache[3][22] , \I_cache/cache[3][23] ,
         \I_cache/cache[3][24] , \I_cache/cache[3][25] ,
         \I_cache/cache[3][26] , \I_cache/cache[3][27] ,
         \I_cache/cache[3][28] , \I_cache/cache[3][29] ,
         \I_cache/cache[3][30] , \I_cache/cache[3][31] ,
         \I_cache/cache[3][32] , \I_cache/cache[3][33] ,
         \I_cache/cache[3][34] , \I_cache/cache[3][35] ,
         \I_cache/cache[3][36] , \I_cache/cache[3][37] ,
         \I_cache/cache[3][38] , \I_cache/cache[3][39] ,
         \I_cache/cache[3][40] , \I_cache/cache[3][41] ,
         \I_cache/cache[3][42] , \I_cache/cache[3][43] ,
         \I_cache/cache[3][44] , \I_cache/cache[3][45] ,
         \I_cache/cache[3][46] , \I_cache/cache[3][47] ,
         \I_cache/cache[3][48] , \I_cache/cache[3][49] ,
         \I_cache/cache[3][50] , \I_cache/cache[3][51] ,
         \I_cache/cache[3][52] , \I_cache/cache[3][53] ,
         \I_cache/cache[3][54] , \I_cache/cache[3][55] ,
         \I_cache/cache[3][56] , \I_cache/cache[3][57] ,
         \I_cache/cache[3][58] , \I_cache/cache[3][59] ,
         \I_cache/cache[3][60] , \I_cache/cache[3][61] ,
         \I_cache/cache[3][62] , \I_cache/cache[3][63] ,
         \I_cache/cache[3][64] , \I_cache/cache[3][65] ,
         \I_cache/cache[3][66] , \I_cache/cache[3][67] ,
         \I_cache/cache[3][68] , \I_cache/cache[3][69] ,
         \I_cache/cache[3][70] , \I_cache/cache[3][71] ,
         \I_cache/cache[3][72] , \I_cache/cache[3][73] ,
         \I_cache/cache[3][74] , \I_cache/cache[3][75] ,
         \I_cache/cache[3][76] , \I_cache/cache[3][77] ,
         \I_cache/cache[3][78] , \I_cache/cache[3][79] ,
         \I_cache/cache[3][80] , \I_cache/cache[3][81] ,
         \I_cache/cache[3][82] , \I_cache/cache[3][83] ,
         \I_cache/cache[3][84] , \I_cache/cache[3][85] ,
         \I_cache/cache[3][86] , \I_cache/cache[3][87] ,
         \I_cache/cache[3][88] , \I_cache/cache[3][89] ,
         \I_cache/cache[3][90] , \I_cache/cache[3][91] ,
         \I_cache/cache[3][92] , \I_cache/cache[3][93] ,
         \I_cache/cache[3][94] , \I_cache/cache[3][95] ,
         \I_cache/cache[3][96] , \I_cache/cache[3][97] ,
         \I_cache/cache[3][98] , \I_cache/cache[3][99] ,
         \I_cache/cache[3][100] , \I_cache/cache[3][101] ,
         \I_cache/cache[3][102] , \I_cache/cache[3][103] ,
         \I_cache/cache[3][104] , \I_cache/cache[3][105] ,
         \I_cache/cache[3][106] , \I_cache/cache[3][107] ,
         \I_cache/cache[3][108] , \I_cache/cache[3][109] ,
         \I_cache/cache[3][110] , \I_cache/cache[3][111] ,
         \I_cache/cache[3][112] , \I_cache/cache[3][113] ,
         \I_cache/cache[3][114] , \I_cache/cache[3][115] ,
         \I_cache/cache[3][116] , \I_cache/cache[3][117] ,
         \I_cache/cache[3][118] , \I_cache/cache[3][119] ,
         \I_cache/cache[3][120] , \I_cache/cache[3][121] ,
         \I_cache/cache[3][122] , \I_cache/cache[3][123] ,
         \I_cache/cache[3][124] , \I_cache/cache[3][125] ,
         \I_cache/cache[3][126] , \I_cache/cache[3][127] ,
         \I_cache/cache[3][128] , \I_cache/cache[3][129] ,
         \I_cache/cache[3][130] , \I_cache/cache[3][131] ,
         \I_cache/cache[3][132] , \I_cache/cache[3][133] ,
         \I_cache/cache[3][134] , \I_cache/cache[3][135] ,
         \I_cache/cache[3][136] , \I_cache/cache[3][137] ,
         \I_cache/cache[3][138] , \I_cache/cache[3][139] ,
         \I_cache/cache[3][140] , \I_cache/cache[3][141] ,
         \I_cache/cache[3][142] , \I_cache/cache[3][143] ,
         \I_cache/cache[3][144] , \I_cache/cache[3][145] ,
         \I_cache/cache[3][146] , \I_cache/cache[3][147] ,
         \I_cache/cache[3][148] , \I_cache/cache[3][149] ,
         \I_cache/cache[3][150] , \I_cache/cache[3][151] ,
         \I_cache/cache[3][152] , \I_cache/cache[3][153] ,
         \I_cache/cache[3][154] , \I_cache/cache[2][0] , \I_cache/cache[2][1] ,
         \I_cache/cache[2][2] , \I_cache/cache[2][3] , \I_cache/cache[2][4] ,
         \I_cache/cache[2][5] , \I_cache/cache[2][6] , \I_cache/cache[2][7] ,
         \I_cache/cache[2][8] , \I_cache/cache[2][9] , \I_cache/cache[2][10] ,
         \I_cache/cache[2][11] , \I_cache/cache[2][12] ,
         \I_cache/cache[2][13] , \I_cache/cache[2][14] ,
         \I_cache/cache[2][15] , \I_cache/cache[2][16] ,
         \I_cache/cache[2][17] , \I_cache/cache[2][18] ,
         \I_cache/cache[2][19] , \I_cache/cache[2][20] ,
         \I_cache/cache[2][21] , \I_cache/cache[2][22] ,
         \I_cache/cache[2][23] , \I_cache/cache[2][24] ,
         \I_cache/cache[2][25] , \I_cache/cache[2][26] ,
         \I_cache/cache[2][27] , \I_cache/cache[2][28] ,
         \I_cache/cache[2][29] , \I_cache/cache[2][30] ,
         \I_cache/cache[2][31] , \I_cache/cache[2][32] ,
         \I_cache/cache[2][33] , \I_cache/cache[2][34] ,
         \I_cache/cache[2][35] , \I_cache/cache[2][36] ,
         \I_cache/cache[2][37] , \I_cache/cache[2][38] ,
         \I_cache/cache[2][39] , \I_cache/cache[2][40] ,
         \I_cache/cache[2][41] , \I_cache/cache[2][42] ,
         \I_cache/cache[2][43] , \I_cache/cache[2][44] ,
         \I_cache/cache[2][45] , \I_cache/cache[2][46] ,
         \I_cache/cache[2][47] , \I_cache/cache[2][48] ,
         \I_cache/cache[2][49] , \I_cache/cache[2][50] ,
         \I_cache/cache[2][51] , \I_cache/cache[2][52] ,
         \I_cache/cache[2][53] , \I_cache/cache[2][54] ,
         \I_cache/cache[2][55] , \I_cache/cache[2][56] ,
         \I_cache/cache[2][57] , \I_cache/cache[2][58] ,
         \I_cache/cache[2][59] , \I_cache/cache[2][60] ,
         \I_cache/cache[2][61] , \I_cache/cache[2][62] ,
         \I_cache/cache[2][63] , \I_cache/cache[2][64] ,
         \I_cache/cache[2][65] , \I_cache/cache[2][66] ,
         \I_cache/cache[2][67] , \I_cache/cache[2][68] ,
         \I_cache/cache[2][69] , \I_cache/cache[2][70] ,
         \I_cache/cache[2][71] , \I_cache/cache[2][72] ,
         \I_cache/cache[2][73] , \I_cache/cache[2][74] ,
         \I_cache/cache[2][75] , \I_cache/cache[2][76] ,
         \I_cache/cache[2][77] , \I_cache/cache[2][78] ,
         \I_cache/cache[2][79] , \I_cache/cache[2][80] ,
         \I_cache/cache[2][81] , \I_cache/cache[2][82] ,
         \I_cache/cache[2][83] , \I_cache/cache[2][84] ,
         \I_cache/cache[2][85] , \I_cache/cache[2][86] ,
         \I_cache/cache[2][87] , \I_cache/cache[2][88] ,
         \I_cache/cache[2][89] , \I_cache/cache[2][90] ,
         \I_cache/cache[2][91] , \I_cache/cache[2][92] ,
         \I_cache/cache[2][93] , \I_cache/cache[2][94] ,
         \I_cache/cache[2][95] , \I_cache/cache[2][96] ,
         \I_cache/cache[2][97] , \I_cache/cache[2][98] ,
         \I_cache/cache[2][99] , \I_cache/cache[2][100] ,
         \I_cache/cache[2][101] , \I_cache/cache[2][102] ,
         \I_cache/cache[2][103] , \I_cache/cache[2][104] ,
         \I_cache/cache[2][105] , \I_cache/cache[2][106] ,
         \I_cache/cache[2][107] , \I_cache/cache[2][108] ,
         \I_cache/cache[2][109] , \I_cache/cache[2][110] ,
         \I_cache/cache[2][111] , \I_cache/cache[2][112] ,
         \I_cache/cache[2][113] , \I_cache/cache[2][114] ,
         \I_cache/cache[2][115] , \I_cache/cache[2][116] ,
         \I_cache/cache[2][117] , \I_cache/cache[2][118] ,
         \I_cache/cache[2][119] , \I_cache/cache[2][120] ,
         \I_cache/cache[2][121] , \I_cache/cache[2][122] ,
         \I_cache/cache[2][123] , \I_cache/cache[2][124] ,
         \I_cache/cache[2][125] , \I_cache/cache[2][126] ,
         \I_cache/cache[2][127] , \I_cache/cache[2][128] ,
         \I_cache/cache[2][129] , \I_cache/cache[2][130] ,
         \I_cache/cache[2][131] , \I_cache/cache[2][132] ,
         \I_cache/cache[2][133] , \I_cache/cache[2][134] ,
         \I_cache/cache[2][135] , \I_cache/cache[2][136] ,
         \I_cache/cache[2][137] , \I_cache/cache[2][138] ,
         \I_cache/cache[2][139] , \I_cache/cache[2][140] ,
         \I_cache/cache[2][141] , \I_cache/cache[2][142] ,
         \I_cache/cache[2][143] , \I_cache/cache[2][144] ,
         \I_cache/cache[2][145] , \I_cache/cache[2][146] ,
         \I_cache/cache[2][147] , \I_cache/cache[2][148] ,
         \I_cache/cache[2][149] , \I_cache/cache[2][150] ,
         \I_cache/cache[2][151] , \I_cache/cache[2][152] ,
         \I_cache/cache[2][153] , \I_cache/cache[2][154] ,
         \I_cache/cache[1][0] , \I_cache/cache[1][1] , \I_cache/cache[1][2] ,
         \I_cache/cache[1][3] , \I_cache/cache[1][4] , \I_cache/cache[1][5] ,
         \I_cache/cache[1][6] , \I_cache/cache[1][7] , \I_cache/cache[1][8] ,
         \I_cache/cache[1][9] , \I_cache/cache[1][10] , \I_cache/cache[1][11] ,
         \I_cache/cache[1][12] , \I_cache/cache[1][13] ,
         \I_cache/cache[1][14] , \I_cache/cache[1][15] ,
         \I_cache/cache[1][16] , \I_cache/cache[1][17] ,
         \I_cache/cache[1][18] , \I_cache/cache[1][19] ,
         \I_cache/cache[1][20] , \I_cache/cache[1][21] ,
         \I_cache/cache[1][22] , \I_cache/cache[1][23] ,
         \I_cache/cache[1][24] , \I_cache/cache[1][25] ,
         \I_cache/cache[1][26] , \I_cache/cache[1][27] ,
         \I_cache/cache[1][28] , \I_cache/cache[1][29] ,
         \I_cache/cache[1][30] , \I_cache/cache[1][31] ,
         \I_cache/cache[1][32] , \I_cache/cache[1][33] ,
         \I_cache/cache[1][34] , \I_cache/cache[1][35] ,
         \I_cache/cache[1][36] , \I_cache/cache[1][37] ,
         \I_cache/cache[1][38] , \I_cache/cache[1][39] ,
         \I_cache/cache[1][40] , \I_cache/cache[1][41] ,
         \I_cache/cache[1][42] , \I_cache/cache[1][43] ,
         \I_cache/cache[1][44] , \I_cache/cache[1][45] ,
         \I_cache/cache[1][46] , \I_cache/cache[1][47] ,
         \I_cache/cache[1][48] , \I_cache/cache[1][49] ,
         \I_cache/cache[1][50] , \I_cache/cache[1][51] ,
         \I_cache/cache[1][52] , \I_cache/cache[1][53] ,
         \I_cache/cache[1][54] , \I_cache/cache[1][55] ,
         \I_cache/cache[1][56] , \I_cache/cache[1][57] ,
         \I_cache/cache[1][58] , \I_cache/cache[1][59] ,
         \I_cache/cache[1][60] , \I_cache/cache[1][61] ,
         \I_cache/cache[1][62] , \I_cache/cache[1][63] ,
         \I_cache/cache[1][64] , \I_cache/cache[1][65] ,
         \I_cache/cache[1][66] , \I_cache/cache[1][67] ,
         \I_cache/cache[1][68] , \I_cache/cache[1][69] ,
         \I_cache/cache[1][70] , \I_cache/cache[1][71] ,
         \I_cache/cache[1][72] , \I_cache/cache[1][73] ,
         \I_cache/cache[1][74] , \I_cache/cache[1][75] ,
         \I_cache/cache[1][76] , \I_cache/cache[1][77] ,
         \I_cache/cache[1][78] , \I_cache/cache[1][79] ,
         \I_cache/cache[1][80] , \I_cache/cache[1][81] ,
         \I_cache/cache[1][82] , \I_cache/cache[1][83] ,
         \I_cache/cache[1][84] , \I_cache/cache[1][85] ,
         \I_cache/cache[1][86] , \I_cache/cache[1][87] ,
         \I_cache/cache[1][88] , \I_cache/cache[1][89] ,
         \I_cache/cache[1][90] , \I_cache/cache[1][91] ,
         \I_cache/cache[1][92] , \I_cache/cache[1][93] ,
         \I_cache/cache[1][94] , \I_cache/cache[1][95] ,
         \I_cache/cache[1][96] , \I_cache/cache[1][97] ,
         \I_cache/cache[1][98] , \I_cache/cache[1][99] ,
         \I_cache/cache[1][100] , \I_cache/cache[1][101] ,
         \I_cache/cache[1][102] , \I_cache/cache[1][103] ,
         \I_cache/cache[1][104] , \I_cache/cache[1][105] ,
         \I_cache/cache[1][106] , \I_cache/cache[1][107] ,
         \I_cache/cache[1][108] , \I_cache/cache[1][109] ,
         \I_cache/cache[1][110] , \I_cache/cache[1][111] ,
         \I_cache/cache[1][112] , \I_cache/cache[1][113] ,
         \I_cache/cache[1][114] , \I_cache/cache[1][115] ,
         \I_cache/cache[1][116] , \I_cache/cache[1][117] ,
         \I_cache/cache[1][118] , \I_cache/cache[1][119] ,
         \I_cache/cache[1][120] , \I_cache/cache[1][121] ,
         \I_cache/cache[1][122] , \I_cache/cache[1][123] ,
         \I_cache/cache[1][124] , \I_cache/cache[1][125] ,
         \I_cache/cache[1][126] , \I_cache/cache[1][127] ,
         \I_cache/cache[1][128] , \I_cache/cache[1][129] ,
         \I_cache/cache[1][130] , \I_cache/cache[1][131] ,
         \I_cache/cache[1][132] , \I_cache/cache[1][133] ,
         \I_cache/cache[1][134] , \I_cache/cache[1][135] ,
         \I_cache/cache[1][136] , \I_cache/cache[1][137] ,
         \I_cache/cache[1][138] , \I_cache/cache[1][139] ,
         \I_cache/cache[1][140] , \I_cache/cache[1][141] ,
         \I_cache/cache[1][142] , \I_cache/cache[1][143] ,
         \I_cache/cache[1][144] , \I_cache/cache[1][145] ,
         \I_cache/cache[1][146] , \I_cache/cache[1][147] ,
         \I_cache/cache[1][148] , \I_cache/cache[1][149] ,
         \I_cache/cache[1][150] , \I_cache/cache[1][151] ,
         \I_cache/cache[1][152] , \I_cache/cache[1][153] ,
         \I_cache/cache[1][154] , \I_cache/cache[0][0] , \I_cache/cache[0][1] ,
         \I_cache/cache[0][2] , \I_cache/cache[0][3] , \I_cache/cache[0][4] ,
         \I_cache/cache[0][5] , \I_cache/cache[0][6] , \I_cache/cache[0][7] ,
         \I_cache/cache[0][8] , \I_cache/cache[0][9] , \I_cache/cache[0][10] ,
         \I_cache/cache[0][11] , \I_cache/cache[0][12] ,
         \I_cache/cache[0][13] , \I_cache/cache[0][14] ,
         \I_cache/cache[0][15] , \I_cache/cache[0][16] ,
         \I_cache/cache[0][17] , \I_cache/cache[0][18] ,
         \I_cache/cache[0][19] , \I_cache/cache[0][20] ,
         \I_cache/cache[0][21] , \I_cache/cache[0][22] ,
         \I_cache/cache[0][23] , \I_cache/cache[0][24] ,
         \I_cache/cache[0][25] , \I_cache/cache[0][26] ,
         \I_cache/cache[0][27] , \I_cache/cache[0][28] ,
         \I_cache/cache[0][29] , \I_cache/cache[0][30] ,
         \I_cache/cache[0][31] , \I_cache/cache[0][32] ,
         \I_cache/cache[0][33] , \I_cache/cache[0][34] ,
         \I_cache/cache[0][35] , \I_cache/cache[0][36] ,
         \I_cache/cache[0][37] , \I_cache/cache[0][38] ,
         \I_cache/cache[0][39] , \I_cache/cache[0][40] ,
         \I_cache/cache[0][41] , \I_cache/cache[0][42] ,
         \I_cache/cache[0][43] , \I_cache/cache[0][44] ,
         \I_cache/cache[0][45] , \I_cache/cache[0][46] ,
         \I_cache/cache[0][47] , \I_cache/cache[0][48] ,
         \I_cache/cache[0][49] , \I_cache/cache[0][50] ,
         \I_cache/cache[0][51] , \I_cache/cache[0][52] ,
         \I_cache/cache[0][53] , \I_cache/cache[0][54] ,
         \I_cache/cache[0][55] , \I_cache/cache[0][56] ,
         \I_cache/cache[0][57] , \I_cache/cache[0][58] ,
         \I_cache/cache[0][59] , \I_cache/cache[0][60] ,
         \I_cache/cache[0][61] , \I_cache/cache[0][62] ,
         \I_cache/cache[0][63] , \I_cache/cache[0][64] ,
         \I_cache/cache[0][65] , \I_cache/cache[0][66] ,
         \I_cache/cache[0][67] , \I_cache/cache[0][68] ,
         \I_cache/cache[0][69] , \I_cache/cache[0][70] ,
         \I_cache/cache[0][71] , \I_cache/cache[0][72] ,
         \I_cache/cache[0][73] , \I_cache/cache[0][74] ,
         \I_cache/cache[0][75] , \I_cache/cache[0][76] ,
         \I_cache/cache[0][77] , \I_cache/cache[0][78] ,
         \I_cache/cache[0][79] , \I_cache/cache[0][80] ,
         \I_cache/cache[0][81] , \I_cache/cache[0][82] ,
         \I_cache/cache[0][83] , \I_cache/cache[0][84] ,
         \I_cache/cache[0][85] , \I_cache/cache[0][86] ,
         \I_cache/cache[0][87] , \I_cache/cache[0][88] ,
         \I_cache/cache[0][89] , \I_cache/cache[0][90] ,
         \I_cache/cache[0][91] , \I_cache/cache[0][92] ,
         \I_cache/cache[0][93] , \I_cache/cache[0][94] ,
         \I_cache/cache[0][95] , \I_cache/cache[0][96] ,
         \I_cache/cache[0][97] , \I_cache/cache[0][98] ,
         \I_cache/cache[0][99] , \I_cache/cache[0][100] ,
         \I_cache/cache[0][101] , \I_cache/cache[0][102] ,
         \I_cache/cache[0][103] , \I_cache/cache[0][104] ,
         \I_cache/cache[0][105] , \I_cache/cache[0][106] ,
         \I_cache/cache[0][107] , \I_cache/cache[0][108] ,
         \I_cache/cache[0][109] , \I_cache/cache[0][110] ,
         \I_cache/cache[0][111] , \I_cache/cache[0][112] ,
         \I_cache/cache[0][113] , \I_cache/cache[0][114] ,
         \I_cache/cache[0][115] , \I_cache/cache[0][116] ,
         \I_cache/cache[0][117] , \I_cache/cache[0][118] ,
         \I_cache/cache[0][119] , \I_cache/cache[0][120] ,
         \I_cache/cache[0][121] , \I_cache/cache[0][122] ,
         \I_cache/cache[0][123] , \I_cache/cache[0][124] ,
         \I_cache/cache[0][125] , \I_cache/cache[0][126] ,
         \I_cache/cache[0][127] , \I_cache/cache[0][128] ,
         \I_cache/cache[0][129] , \I_cache/cache[0][130] ,
         \I_cache/cache[0][131] , \I_cache/cache[0][132] ,
         \I_cache/cache[0][133] , \I_cache/cache[0][134] ,
         \I_cache/cache[0][135] , \I_cache/cache[0][136] ,
         \I_cache/cache[0][137] , \I_cache/cache[0][138] ,
         \I_cache/cache[0][139] , \I_cache/cache[0][140] ,
         \I_cache/cache[0][141] , \I_cache/cache[0][142] ,
         \I_cache/cache[0][143] , \I_cache/cache[0][144] ,
         \I_cache/cache[0][145] , \I_cache/cache[0][146] ,
         \I_cache/cache[0][147] , \I_cache/cache[0][148] ,
         \I_cache/cache[0][149] , \I_cache/cache[0][150] ,
         \I_cache/cache[0][151] , \I_cache/cache[0][152] ,
         \I_cache/cache[0][153] , \I_cache/cache[0][154] , net97410, net97416,
         net97418, net97444, net97445, net97452, net97496, net97574, net97592,
         net97684, net97686, net97687, net97701, net97703, net97736, net97753,
         net97755, net97770, net97798, net97800, net97815, net97817, net97834,
         net97874, net97936, net97937, net97995, net98012, net98027, net98029,
         net98044, net98046, net98061, net98063, net98080, net98216, net98217,
         net98231, net98335, net98336, net98340, net98341, net98351, net98352,
         net98363, net98364, net98366, net98367, net98371, net98372, net98375,
         net98380, net98385, net98386, net98390, net98391, net98393, net98487,
         net98495, net98496, net98497, net98499, net98500, net98501, net98502,
         net98514, net98530, net98531, net98550, net98571, net98572, net98598,
         net98630, net98662, net98663, net98707, net98708, net98722, net98728,
         net98755, net98758, net98759, net98776, net98777, net98780, net98781,
         net99002, net99003, net99118, net99151, net99157, net99161, net99164,
         net99165, net99633, net99634, net99635, net99636, net100396,
         net100397, net100398, net100400, net100401, net100415, net100416,
         net100417, net100424, net100426, net100478, net100535, net100537,
         net100573, net100574, net100581, net100583, net100585, net100597,
         net100599, net100601, net100603, net100682, net100791, net101082,
         net101257, net101401, net101402, net101465, net101552, net101554,
         net101555, net101556, net101771, net101906, net101908, net101910,
         net101914, net101978, net102048, net102049, net102050, net102051,
         net102253, net102393, net102404, net102405, net102426, net102427,
         net102428, net102429, net102430, net102431, net102554, net102555,
         net102573, net102790, net102791, net102792, net102878, net102937,
         net102938, net102939, net103025, net103060, net103070, net103076,
         net103079, net103089, net103090, net103091, net103092, net103093,
         net103177, net103224, net103249, net103250, net103251, net103252,
         net103253, net103354, net103416, net103417, net103418, net103504,
         net103548, net103552, net103561, net103581, net103582, net103583,
         net103710, net103718, net103719, net103720, net103721, net103722,
         net103806, net103840, net103889, net103891, net103907, net103910,
         net103911, net103913, net103914, net103917, net103919, net103923,
         net103924, net103954, net103955, net103956, net104042, net104105,
         net104106, net104107, net104108, net104109, net104229, net104230,
         net104248, net104251, net104252, net104253, net104254, net104255,
         net104407, net104408, net104409, net104410, net104411, net104495,
         net104582, net104583, net104584, net104739, net104740, net104741,
         net104864, net104866, net104868, net104885, net104887, net104889,
         net105012, net105034, net105038, net105043, net105045, net105046,
         net105047, net105048, net105049, net105194, net105195, net105196,
         net105282, net105349, net105350, net105600, net105677, net105777,
         net105781, net105783, net105787, net107808, net107804, net107802,
         net107798, net107796, net107794, net107812, net107810, net107816,
         net108156, net108154, net108150, net108132, net108128, net108126,
         net108118, net108116, net108114, net108112, net108110, net108108,
         net108098, net108160, net108200, net108198, net108194, net108192,
         net108190, net108664, net108662, net108660, net108658, net108670,
         net108682, net108680, net108678, net108676, net108674, net108690,
         net108688, net108686, net108710, net108708, net108704, net108702,
         net111630, net111628, net111624, net111622, net111636, net111634,
         net111646, net111644, net111642, net111640, net111910, net111906,
         net111904, net111902, net111964, net111962, net111960, net111968,
         net111966, net111992, net111996, net111994, net112008, net112006,
         net112004, net112002, net112000, net112014, net112026, net112020,
         net112018, net112034, net112032, net112030, net112038, net112036,
         net112050, net112046, net112078, net112076, net112072, net112084,
         net112104, net112100, net112098, net112096, net112090, net112116,
         net112112, net112110, net112134, net112132, net112128, net112142,
         net112138, net112160, net112158, net112152, net112150, net112148,
         net112178, net112176, net112172, net112170, net112166, net112164,
         net112196, net112188, net112182, net112214, net112232, net112228,
         net112224, net112222, net112218, net112250, net112248, net112246,
         net112244, net112242, net112240, net112236, net112268, net112266,
         net112264, net112260, net112258, net112254, net112286, net112306,
         net112304, net112300, net112296, net112294, net112292, net112340,
         net112338, net112336, net112334, net112332, net112330, net112356,
         net112350, net112348, net112346, net112376, net112374, net112372,
         net112370, net112368, net112366, net112364, net112400, net112404,
         net112406, net112415, net112420, net112438, net112676, net112691,
         net112736, net112764, net112782, net112786, net112799, net112962,
         net112999, net127703, net127702, net127709, net127710, net127829,
         net127833, net127930, net127933, net128151, net128154, net128155,
         net128156, net128157, net128158, net128159, net128160, net128161,
         net128301, net128830, net128955, net128963, net129005, net129017,
         net129024, net129200, net133317, net133411, net133414, net133468,
         net133469, net133470, net133471, net133496, net133585, net133688,
         net137684, net137891, net137952, net137951, net138001, net138000,
         net138213, net98620, net100404, net100403, net100402, net97783,
         net105676, net105008, net105007, net105006, net104888, net102784,
         net102783, net102782, net102781, net100399, net101413,
         \i_MIPS/ALU_Control/n10 , n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n169, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n244, n246, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
         n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
         n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
         n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
         n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
         n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
         n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531,
         n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541,
         n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551,
         n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
         n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571,
         n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
         n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591,
         n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
         n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
         n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
         n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
         n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
         n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651,
         n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661,
         n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671,
         n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681,
         n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691,
         n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701,
         n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711,
         n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721,
         n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731,
         n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741,
         n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751,
         n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761,
         n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771,
         n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781,
         n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791,
         n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801,
         n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811,
         n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821,
         n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831,
         n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841,
         n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851,
         n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861,
         n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
         n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881,
         n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891,
         n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901,
         n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911,
         n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921,
         n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931,
         n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941,
         n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951,
         n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961,
         n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971,
         n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981,
         n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991,
         n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001,
         n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011,
         n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021,
         n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031,
         n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041,
         n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051,
         n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061,
         n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071,
         n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081,
         n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091,
         n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101,
         n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111,
         n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121,
         n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131,
         n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141,
         n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151,
         n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161,
         n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171,
         n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181,
         n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191,
         n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201,
         n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211,
         n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221,
         n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231,
         n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241,
         n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251,
         n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261,
         n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271,
         n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281,
         n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291,
         n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301,
         n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311,
         n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321,
         n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331,
         n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341,
         n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351,
         n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361,
         n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371,
         n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381,
         n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391,
         n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401,
         n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411,
         n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421,
         n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431,
         n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441,
         n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451,
         n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461,
         n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471,
         n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481,
         n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491,
         n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501,
         n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511,
         n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521,
         n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531,
         n2532, n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541,
         n2542, n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551,
         n2552, n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561,
         n2562, n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571,
         n2572, n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581,
         n2582, n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591,
         n2592, n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601,
         n2602, n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611,
         n2612, n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621,
         n2622, n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631,
         n2632, n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641,
         n2642, n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651,
         n2652, n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661,
         n2662, n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671,
         n2672, n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681,
         n2682, n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691,
         n2692, n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701,
         n2702, n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711,
         n2712, n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721,
         n2722, n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731,
         n2732, n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741,
         n2742, n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751,
         n2752, n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761,
         n2762, n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771,
         n2772, n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781,
         n2782, n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791,
         n2792, n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801,
         n2802, n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811,
         n2812, n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821,
         n2822, n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831,
         n2832, n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841,
         n2842, n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851,
         n2852, n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861,
         n2862, n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871,
         n2872, n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881,
         n2882, n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891,
         n2892, n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901,
         n2902, n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911,
         n2912, n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921,
         n2922, n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931,
         n2932, n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941,
         n2942, n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951,
         n2952, n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961,
         n2962, n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971,
         n2972, n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981,
         n2982, n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991,
         n2992, n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001,
         n3002, n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011,
         n3012, n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021,
         n3022, n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031,
         n3032, n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041,
         n3042, n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051,
         n3052, n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061,
         n3062, n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071,
         n3072, n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081,
         n3082, n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091,
         n3092, n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101,
         n3102, n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111,
         n3112, n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121,
         n3122, n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131,
         n3132, n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141,
         n3142, n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151,
         n3152, n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161,
         n3162, n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171,
         n3172, n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181,
         n3182, n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191,
         n3192, n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201,
         n3202, n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211,
         n3212, n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221,
         n3222, n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231,
         n3232, n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241,
         n3242, n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251,
         n3252, n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261,
         n3262, n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271,
         n3272, n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281,
         n3282, n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291,
         n3292, n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301,
         n3302, n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311,
         n3312, n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321,
         n3322, n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331,
         n3332, n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341,
         n3342, n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3619, n3621, n3634, n3635, n3636, n3637, n3638,
         n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3683, n3684, n3685, n3686, n3687, n3688, n3689,
         n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699,
         n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709,
         n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719,
         n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729,
         n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739,
         n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749,
         n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759,
         n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769,
         n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779,
         n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789,
         n3790, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3858, n3860, n3865, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3880, n3881, n3882, n3883, n3884, n3889, n3890, n3891, n3892, n3893,
         n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
         n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913, n3914,
         n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923, n3924,
         n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933, n3934,
         n3935, n3936, n3945, n3946, n3947, n3948, n3952, n3953, n3954, n3955,
         n3956, n3957, n3958, n3959, n3960, n4002, n4009, n4015, n4018, n4027,
         n4033, n4036, n4042, n4045, n4048, n4057, n4059, n4060, n4062, n4064,
         n4066, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077,
         n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087,
         n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097,
         n4098, n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107,
         n4108, n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117,
         n4118, n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127,
         n4128, n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137,
         n4138, n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147,
         n4148, n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157,
         n4158, n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167,
         n4168, n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177,
         n4178, n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187,
         n4188, n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197,
         n4198, n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207,
         n4208, n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217,
         n4218, n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227,
         n4228, n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237,
         n4238, n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247,
         n4248, n4249, n4250, n4251, n4289, n4291, n4293, n4295, n4296, n4297,
         n4298, n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307,
         n4308, n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317,
         n4318, n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327,
         n4328, n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337,
         n4338, n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347,
         n4348, n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357,
         n4358, n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367,
         n4368, n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377,
         n4378, n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387,
         n4388, n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397,
         n4398, n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407,
         n4408, n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417,
         n4418, n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427,
         n4428, n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437,
         n4438, n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447,
         n4448, n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457,
         n4458, n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467,
         n4468, n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477,
         n4478, n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487,
         n4488, n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497,
         n4498, n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507,
         n4508, n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517,
         n4518, n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527,
         n4528, n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537,
         n4538, n4539, n4540, n4541, n4542, n4543, n4544, n4570, n4571, n4587,
         n4592, n4593, n4594, n4596, n4598, n4600, n4601, n4602, n4603, n4604,
         n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613, n4614,
         n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623, n4624,
         n4625, n4626, n4627, n4628, n4629, n4631, n4633, n4636, n4637, n4638,
         n4639, n4640, n4641, n4648, n4649, n4650, n4651, n4652, n4653, n4654,
         n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663, n4664,
         n4665, n4666, n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675,
         n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685,
         n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695,
         n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705,
         n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715,
         n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725,
         n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735,
         n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745,
         n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755,
         n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765,
         n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775,
         n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785,
         n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795,
         n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805,
         n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815,
         n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825,
         n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835,
         n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845,
         n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855,
         n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865,
         n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875,
         n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885,
         n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895,
         n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905,
         n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915,
         n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925,
         n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935,
         n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945,
         n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955,
         n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965,
         n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975,
         n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985,
         n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995,
         n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005,
         n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015,
         n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025,
         n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035,
         n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045,
         n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055,
         n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065,
         n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075,
         n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085,
         n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095,
         n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105,
         n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115,
         n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125,
         n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135,
         n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145,
         n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155,
         n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165,
         n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175,
         n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185,
         n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195,
         n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205,
         n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215,
         n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225,
         n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235,
         n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245,
         n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255,
         n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265,
         n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275,
         n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285,
         n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295,
         n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305,
         n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315,
         n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325,
         n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335,
         n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345,
         n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355,
         n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365,
         n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375,
         n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385,
         n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395,
         n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405,
         n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415,
         n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425,
         n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435,
         n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445,
         n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455,
         n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465,
         n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475,
         n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485,
         n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495,
         n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505,
         n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515,
         n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523, n5524, n5525,
         n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533, n5534, n5535,
         n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543, n5544, n5545,
         n5546, n5547, n5548, n5549, n5551, n5554, n5556, n5557, n5558, n5559,
         n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569,
         n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579,
         n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589,
         n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599,
         n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609,
         n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619,
         n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629,
         n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639,
         n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649,
         n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659,
         n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669,
         n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679,
         n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689,
         n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699,
         n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709,
         n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719,
         n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729,
         n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739,
         n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749,
         n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759,
         n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769,
         n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779,
         n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789,
         n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799,
         n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809,
         n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819,
         n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829,
         n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839,
         n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849,
         n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859,
         n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869,
         n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879,
         n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889,
         n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899,
         n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909,
         n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919,
         n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929,
         n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939,
         n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949,
         n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959,
         n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969,
         n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979,
         n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989,
         n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999,
         n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009,
         n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019,
         n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029,
         n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039,
         n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049,
         n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059,
         n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069,
         n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079,
         n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089,
         n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099,
         n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109,
         n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119,
         n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129,
         n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139,
         n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149,
         n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159,
         n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169,
         n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179,
         n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189,
         n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199,
         n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209,
         n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219,
         n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229,
         n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239,
         n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249,
         n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259,
         n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269,
         n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279,
         n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289,
         n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299,
         n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309,
         n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319,
         n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329,
         n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339,
         n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349,
         n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359,
         n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369,
         n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379,
         n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389,
         n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399,
         n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409,
         n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419,
         n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429,
         n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439,
         n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449,
         n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459,
         n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469,
         n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479,
         n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489,
         n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499,
         n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509,
         n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519,
         n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529,
         n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539,
         n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549,
         n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559,
         n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569,
         n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579,
         n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589,
         n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599,
         n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609,
         n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619,
         n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629,
         n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639,
         n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649,
         n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659,
         n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669,
         n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679,
         n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689,
         n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699,
         n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709,
         n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719,
         n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729,
         n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739,
         n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749,
         n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759,
         n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769,
         n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779,
         n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789,
         n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799,
         n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809,
         n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819,
         n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829,
         n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839,
         n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849,
         n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859,
         n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869,
         n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879,
         n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889,
         n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899,
         n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909,
         n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919,
         n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929,
         n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939,
         n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949,
         n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959,
         n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969,
         n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979,
         n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989,
         n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999,
         n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009,
         n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019,
         n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029,
         n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039,
         n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049,
         n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059,
         n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069,
         n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079,
         n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089,
         n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099,
         n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109,
         n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119,
         n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129,
         n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139,
         n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149,
         n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159,
         n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169,
         n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179,
         n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189,
         n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199,
         n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209,
         n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219,
         n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229,
         n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239,
         n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249,
         n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259,
         n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269,
         n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279,
         n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289,
         n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299,
         n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309,
         n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319,
         n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329,
         n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339,
         n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349,
         n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359,
         n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369,
         n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379,
         n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389,
         n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399,
         n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409,
         n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419,
         n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429,
         n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439,
         n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449,
         n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459,
         n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469,
         n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479,
         n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489,
         n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499,
         n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509,
         n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519,
         n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529,
         n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539,
         n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549,
         n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559,
         n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569,
         n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579,
         n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589,
         n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599,
         n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609,
         n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619,
         n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629,
         n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639,
         n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649,
         n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659,
         n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669,
         n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679,
         n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689,
         n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699,
         n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709,
         n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719,
         n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729,
         n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739,
         n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749,
         n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759,
         n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769,
         n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779,
         n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789,
         n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799,
         n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809,
         n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819,
         n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829,
         n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839,
         n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849,
         n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859,
         n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869,
         n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879,
         n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889,
         n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899,
         n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909,
         n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919,
         n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929,
         n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939,
         n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949,
         n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959,
         n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969,
         n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979,
         n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989,
         n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999,
         n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009,
         n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019,
         n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029,
         n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039,
         n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049,
         n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059,
         n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069,
         n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079,
         n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089,
         n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099,
         n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109,
         n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119,
         n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129,
         n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139,
         n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149,
         n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159,
         n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169,
         n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179,
         n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189,
         n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199,
         n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209,
         n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219,
         n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229,
         n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239,
         n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249,
         n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259,
         n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269,
         n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279,
         n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289,
         n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299,
         n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309,
         n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319,
         n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329,
         n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339,
         n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349,
         n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359,
         n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369,
         n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379,
         n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389,
         n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399,
         n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409,
         n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419,
         n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429,
         n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439,
         n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449,
         n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459,
         n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469,
         n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479,
         n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489,
         n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499,
         n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509,
         n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519,
         n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529,
         n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539,
         n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549,
         n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559,
         n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569,
         n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579,
         n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589,
         n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599,
         n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609,
         n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619,
         n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629,
         n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639,
         n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649,
         n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659,
         n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669,
         n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679,
         n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689,
         n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699,
         n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709,
         n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719,
         n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729,
         n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739,
         n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749,
         n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759,
         n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769,
         n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779,
         n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789,
         n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799,
         n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809,
         n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819,
         n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829,
         n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839,
         n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849,
         n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859,
         n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869,
         n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879,
         n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889,
         n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899,
         n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909,
         n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919,
         n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929,
         n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939,
         n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949,
         n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959,
         n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969,
         n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979,
         n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989,
         n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999,
         n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009,
         n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019,
         n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029,
         n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039,
         n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049,
         n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059,
         n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069,
         n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079,
         n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089,
         n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099,
         n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109,
         n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119,
         n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129,
         n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139,
         n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149,
         n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159,
         n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169,
         n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179,
         n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189,
         n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199,
         n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209,
         n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219,
         n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229,
         n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239,
         n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249,
         n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259,
         n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269,
         n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279,
         n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289,
         n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299,
         n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309,
         n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319,
         n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329,
         n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339,
         n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349,
         n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359,
         n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369,
         n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379,
         n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389,
         n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399,
         n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409,
         n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419,
         n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429,
         n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439,
         n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449,
         n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459,
         n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469,
         n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479,
         n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489,
         n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499,
         n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509,
         n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519,
         n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529,
         n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539,
         n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549,
         n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559,
         n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569,
         n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579,
         n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589,
         n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599,
         n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609,
         n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619,
         n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629,
         n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639,
         n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649,
         n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659,
         n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669,
         n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679,
         n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689,
         n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699,
         n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709,
         n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719,
         n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729,
         n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739,
         n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749,
         n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759,
         n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769,
         n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779,
         n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789,
         n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799,
         n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809,
         n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819,
         n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829,
         n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839,
         n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849,
         n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859,
         n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869,
         n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879,
         n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889,
         n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899,
         n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909,
         n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919,
         n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929,
         n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939,
         n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949,
         n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959,
         n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969,
         n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979,
         n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989,
         n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999,
         n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
         n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567,
         n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
         n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
         n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591,
         n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
         n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
         n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
         n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
         n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
         n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
         n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
         n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
         n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
         n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
         n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
         n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
         n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
         n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
         n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
         n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
         n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
         n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759,
         n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767,
         n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
         n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783,
         n12784, n12785, n12786, n12787;
  wire   [29:0] ICACHE_addr;
  assign DCACHE_addr[0] = net112962;

  DFFRX4 \i_MIPS/EX_MEM_reg[9]  ( .D(\i_MIPS/n465 ), .CK(clk), .RN(n5744), .Q(
        n12953), .QN(n4295) );
  DFFRX4 \i_MIPS/ID_EX_reg[7]  ( .D(\i_MIPS/n471 ), .CK(clk), .RN(n5743), .Q(
        \i_MIPS/ALUOp[1] ), .QN(n3820) );
  DFFRX4 \i_MIPS/ID_EX_reg[5]  ( .D(\i_MIPS/n478 ), .CK(clk), .RN(n5742), .Q(
        \i_MIPS/ID_EX_5 ) );
  DFFRX4 \i_MIPS/ID_EX_reg[83]  ( .D(\i_MIPS/n502 ), .CK(clk), .RN(n5740), .Q(
        \i_MIPS/ID_EX[83] ), .QN(n4535) );
  DFFRX4 \i_MIPS/ID_EX_reg[82]  ( .D(\i_MIPS/n503 ), .CK(clk), .RN(n5740), .Q(
        \i_MIPS/ID_EX[82] ), .QN(n4536) );
  DFFRX4 \i_MIPS/ID_EX_reg[81]  ( .D(\i_MIPS/n504 ), .CK(clk), .RN(n5740), .Q(
        \i_MIPS/ID_EX[81] ), .QN(n3837) );
  DFFRX4 \i_MIPS/ID_EX_reg[80]  ( .D(\i_MIPS/n505 ), .CK(clk), .RN(n5740), .Q(
        \i_MIPS/ID_EX[80] ), .QN(net112764) );
  DFFRX4 \i_MIPS/ID_EX_reg[79]  ( .D(\i_MIPS/n506 ), .CK(clk), .RN(n5740), .Q(
        \i_MIPS/ID_EX[79] ), .QN(n3839) );
  DFFRX4 \i_MIPS/ID_EX_reg[78]  ( .D(\i_MIPS/n507 ), .CK(clk), .RN(n5740), .Q(
        \i_MIPS/ID_EX[78] ), .QN(net127930) );
  DFFRX4 \i_MIPS/ID_EX_reg[77]  ( .D(\i_MIPS/n508 ), .CK(clk), .RN(n5740), .Q(
        \i_MIPS/ID_EX[77] ), .QN(net127933) );
  DFFRX4 \i_MIPS/ID_EX_reg[75]  ( .D(\i_MIPS/n510 ), .CK(clk), .RN(n5740), .Q(
        \i_MIPS/ID_EX[75] ), .QN(n3836) );
  DFFRX4 \i_MIPS/ID_EX_reg[73]  ( .D(\i_MIPS/n512 ), .CK(clk), .RN(n5739), .Q(
        \i_MIPS/ID_EX[73] ), .QN(net137684) );
  DFFRX4 \i_MIPS/IF_ID_reg[48]  ( .D(\i_MIPS/N74 ), .CK(clk), .RN(n5738), .Q(
        \i_MIPS/IR_ID[16] ), .QN(\i_MIPS/n312 ) );
  DFFRX4 \i_MIPS/IF_ID_reg[50]  ( .D(\i_MIPS/N76 ), .CK(clk), .RN(n5738), .Q(
        \i_MIPS/IR_ID[18] ), .QN(\i_MIPS/n316 ) );
  DFFRX4 \i_MIPS/IF_ID_reg[51]  ( .D(\i_MIPS/N77 ), .CK(clk), .RN(n5737), .Q(
        \i_MIPS/IR_ID[19] ), .QN(\i_MIPS/n318 ) );
  DFFRX4 \i_MIPS/IF_ID_reg[53]  ( .D(\i_MIPS/N79 ), .CK(clk), .RN(n5737), .Q(
        \i_MIPS/IR_ID[21] ), .QN(\i_MIPS/n231 ) );
  DFFRX4 \i_MIPS/IF_ID_reg[54]  ( .D(\i_MIPS/N80 ), .CK(clk), .RN(n5737), .Q(
        \i_MIPS/IR_ID[22] ), .QN(\i_MIPS/n232 ) );
  DFFRX4 \i_MIPS/IF_ID_reg[55]  ( .D(\i_MIPS/N81 ), .CK(clk), .RN(n5737), .Q(
        \i_MIPS/IR_ID[23] ), .QN(\i_MIPS/n233 ) );
  DFFRX4 \i_MIPS/ID_EX_reg[28]  ( .D(\i_MIPS/n543 ), .CK(clk), .RN(n5714), .Q(
        \i_MIPS/ALUin1[19] ), .QN(\i_MIPS/n352 ) );
  DFFRX4 \i_MIPS/ID_EX_reg[25]  ( .D(\i_MIPS/n546 ), .CK(clk), .RN(n5714), .Q(
        \i_MIPS/ALUin1[16] ), .QN(\i_MIPS/n355 ) );
  DFFRX4 \i_MIPS/ID_EX_reg[20]  ( .D(\i_MIPS/n551 ), .CK(clk), .RN(n5714), .Q(
        \i_MIPS/ALUin1[11] ), .QN(\i_MIPS/n360 ) );
  DFFRX4 \i_MIPS/ID_EX_reg[18]  ( .D(\i_MIPS/n553 ), .CK(clk), .RN(n5713), .Q(
        \i_MIPS/ALUin1[9] ), .QN(\i_MIPS/n362 ) );
  DFFRX4 \i_MIPS/ID_EX_reg[17]  ( .D(\i_MIPS/n554 ), .CK(clk), .RN(n5713), .Q(
        \i_MIPS/ALUin1[8] ), .QN(\i_MIPS/n363 ) );
  DFFRX4 \i_MIPS/ID_EX_reg[16]  ( .D(\i_MIPS/n555 ), .CK(clk), .RN(n5713), .Q(
        \i_MIPS/ALUin1[7] ), .QN(\i_MIPS/n364 ) );
  DFFRX4 \i_MIPS/ID_EX_reg[15]  ( .D(\i_MIPS/n556 ), .CK(clk), .RN(n5713), .Q(
        \i_MIPS/ALUin1[6] ), .QN(\i_MIPS/n365 ) );
  DFFRX4 \i_MIPS/PC/PC_o_reg[3]  ( .D(\i_MIPS/PC/n37 ), .CK(clk), .RN(n5712), 
        .Q(ICACHE_addr[1]), .QN(\i_MIPS/PC/n5 ) );
  DFFRX4 \i_MIPS/PC/PC_o_reg[5]  ( .D(\i_MIPS/PC/n39 ), .CK(clk), .RN(n5711), 
        .Q(ICACHE_addr[3]), .QN(\i_MIPS/PC/n7 ) );
  DFFRX1 \i_MIPS/PHT_2/current_state_2_reg[0]  ( .D(\i_MIPS/PHT_2/n47 ), .CK(
        clk), .RN(n5712), .Q(\i_MIPS/PHT_2/current_state_2[0] ), .QN(
        \i_MIPS/PHT_2/n6 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[13]  ( .D(\i_MIPS/N39 ), .CK(clk), .RN(n5732), .QN(
        \i_MIPS/n196 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[1]  ( .D(\i_MIPS/N27 ), .CK(clk), .RN(n5731), .QN(
        \i_MIPS/n184 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[0]  ( .D(\i_MIPS/N26 ), .CK(clk), .RN(n5731), .QN(
        \i_MIPS/n183 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[65]  ( .D(\i_MIPS/N91 ), .CK(clk), .RN(n5734), .Q(
        \i_MIPS/IF_ID[65] ), .QN(\i_MIPS/n237 ) );
  DFFSX1 \i_MIPS/PHT_2/current_state_3_reg[1]  ( .D(\i_MIPS/PHT_2/n44 ), .CK(
        clk), .SN(n5950), .Q(n406) );
  DFFRX1 \i_MIPS/PHT_2/counter_reg  ( .D(\i_MIPS/PHT_2/n54 ), .CK(clk), .RN(
        n5712), .Q(\i_MIPS/PHT_2/counter ) );
  DFFRX1 \i_MIPS/IF_ID_reg[30]  ( .D(\i_MIPS/N56 ), .CK(clk), .RN(n5734), .Q(
        \i_MIPS/IF_ID_30 ), .QN(\i_MIPS/n213 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[4]  ( .D(\i_MIPS/n480 ), .CK(clk), .RN(n5742), .Q(
        n3614), .QN(\i_MIPS/n311 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[1]  ( .D(\i_MIPS/n527 ), .CK(clk), .RN(n5716), .Q(
        n3609), .QN(\i_MIPS/n337 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[116]  ( .D(\i_MIPS/n530 ), .CK(clk), .RN(n5715), 
        .Q(n3608), .QN(\i_MIPS/n339 ) );
  DFFRX1 \i_MIPS/PHT_2/current_state_3_reg[0]  ( .D(\i_MIPS/PHT_2/n45 ), .CK(
        clk), .RN(n5712), .Q(\i_MIPS/PHT_2/current_state_3[0] ), .QN(
        \i_MIPS/PHT_2/n2 ) );
  DFFSX1 \i_MIPS/PHT_2/current_state_1_reg[1]  ( .D(\i_MIPS/PHT_2/n48 ), .CK(
        clk), .SN(n5949), .Q(\i_MIPS/PHT_2/current_state_1[1] ), .QN(
        \i_MIPS/PHT_2/n7 ) );
  DFFSX1 \i_MIPS/PHT_2/current_state_0_reg[1]  ( .D(\i_MIPS/PHT_2/n50 ), .CK(
        clk), .SN(n5950), .Q(\i_MIPS/PHT_2/current_state_0[1] ), .QN(
        \i_MIPS/PHT_2/n3 ) );
  DFFSX1 \i_MIPS/PHT_2/current_state_2_reg[1]  ( .D(\i_MIPS/PHT_2/n46 ), .CK(
        clk), .SN(n5949), .Q(\i_MIPS/PHT_2/current_state_2[1] ), .QN(
        \i_MIPS/PHT_2/n5 ) );
  DFFRX1 \i_MIPS/PHT_2/current_state_0_reg[0]  ( .D(n11509), .CK(clk), .RN(
        n5712), .Q(n3605), .QN(\i_MIPS/PHT_2/n4 ) );
  DFFRX1 \i_MIPS/PHT_2/history_state_reg[1]  ( .D(\i_MIPS/PHT_2/n53 ), .CK(clk), .RN(n5712), .Q(\i_MIPS/PHT_2/history_state[1] ), .QN(\i_MIPS/PHT_2/n12 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[3]  ( .D(\i_MIPS/n525 ), .CK(clk), .RN(n5716), .Q(
        \i_MIPS/ID_EX_3 ), .QN(\i_MIPS/n335 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[74]  ( .D(\i_MIPS/n529 ), .CK(clk), .RN(n5715), 
        .Q(\i_MIPS/EX_MEM_74 ), .QN(\i_MIPS/n338 ) );
  DFFRX1 \i_MIPS/Register/register_reg[12][27]  ( .D(\i_MIPS/Register/n751 ), 
        .CK(clk), .RN(n5656), .Q(\i_MIPS/Register/register[12][27] ), .QN(n285) );
  DFFRX1 \i_MIPS/EX_MEM_reg[6]  ( .D(\i_MIPS/n468 ), .CK(clk), .RN(n5743), .Q(
        \i_MIPS/EX_MEM[6] ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[5]  ( .D(\i_MIPS/n469 ), .CK(clk), .RN(n5743), .Q(
        \i_MIPS/EX_MEM[5] ) );
  DFFRX1 \I_cache/cache_reg[0][16]  ( .D(n12659), .CK(clk), .RN(n5909), .Q(
        \I_cache/cache[0][16] ), .QN(n1907) );
  DFFRX1 \I_cache/cache_reg[1][16]  ( .D(n12658), .CK(clk), .RN(n5909), .Q(
        \I_cache/cache[1][16] ), .QN(n3562) );
  DFFRX1 \I_cache/cache_reg[2][16]  ( .D(n12657), .CK(clk), .RN(n5909), .Q(
        \I_cache/cache[2][16] ), .QN(n1908) );
  DFFRX1 \I_cache/cache_reg[3][16]  ( .D(n12656), .CK(clk), .RN(n5908), .Q(
        \I_cache/cache[3][16] ), .QN(n3563) );
  DFFRX1 \I_cache/cache_reg[4][16]  ( .D(n12655), .CK(clk), .RN(n5908), .Q(
        \I_cache/cache[4][16] ), .QN(n1849) );
  DFFRX1 \I_cache/cache_reg[5][16]  ( .D(n12654), .CK(clk), .RN(n5908), .Q(
        \I_cache/cache[5][16] ), .QN(n3505) );
  DFFRX1 \I_cache/cache_reg[6][16]  ( .D(n12653), .CK(clk), .RN(n5908), .Q(
        \I_cache/cache[6][16] ), .QN(n1931) );
  DFFRX1 \I_cache/cache_reg[7][16]  ( .D(n12652), .CK(clk), .RN(n5908), .Q(
        \I_cache/cache[7][16] ), .QN(n3585) );
  DFFRX1 \I_cache/cache_reg[0][17]  ( .D(n12651), .CK(clk), .RN(n5908), .Q(
        \I_cache/cache[0][17] ), .QN(n1898) );
  DFFRX1 \I_cache/cache_reg[1][17]  ( .D(n12650), .CK(clk), .RN(n5908), .Q(
        \I_cache/cache[1][17] ), .QN(n3553) );
  DFFRX1 \I_cache/cache_reg[2][17]  ( .D(n12649), .CK(clk), .RN(n5908), .Q(
        \I_cache/cache[2][17] ), .QN(n1899) );
  DFFRX1 \I_cache/cache_reg[3][17]  ( .D(n12648), .CK(clk), .RN(n5908), .Q(
        \I_cache/cache[3][17] ), .QN(n3554) );
  DFFRX1 \I_cache/cache_reg[4][17]  ( .D(n12647), .CK(clk), .RN(n5908), .Q(
        \I_cache/cache[4][17] ), .QN(n1829) );
  DFFRX1 \I_cache/cache_reg[5][17]  ( .D(n12646), .CK(clk), .RN(n5908), .Q(
        \I_cache/cache[5][17] ), .QN(n3485) );
  DFFRX1 \I_cache/cache_reg[6][17]  ( .D(n12645), .CK(clk), .RN(n5908), .Q(
        \I_cache/cache[6][17] ), .QN(n1927) );
  DFFRX1 \I_cache/cache_reg[7][17]  ( .D(n12644), .CK(clk), .RN(n5907), .Q(
        \I_cache/cache[7][17] ), .QN(n3581) );
  DFFRX1 \I_cache/cache_reg[0][18]  ( .D(n12643), .CK(clk), .RN(n5907), .Q(
        \I_cache/cache[0][18] ), .QN(n1893) );
  DFFRX1 \I_cache/cache_reg[1][18]  ( .D(n12642), .CK(clk), .RN(n5907), .Q(
        \I_cache/cache[1][18] ), .QN(n3548) );
  DFFRX1 \I_cache/cache_reg[2][18]  ( .D(n12641), .CK(clk), .RN(n5907), .Q(
        \I_cache/cache[2][18] ), .QN(n1862) );
  DFFRX1 \I_cache/cache_reg[3][18]  ( .D(n12640), .CK(clk), .RN(n5907), .Q(
        \I_cache/cache[3][18] ), .QN(n3518) );
  DFFRX1 \I_cache/cache_reg[4][18]  ( .D(n12639), .CK(clk), .RN(n5907), .Q(
        \I_cache/cache[4][18] ), .QN(n1861) );
  DFFRX1 \I_cache/cache_reg[5][18]  ( .D(n12638), .CK(clk), .RN(n5907), .Q(
        \I_cache/cache[5][18] ), .QN(n3517) );
  DFFRX1 \I_cache/cache_reg[6][18]  ( .D(n12637), .CK(clk), .RN(n5907), .Q(
        \I_cache/cache[6][18] ), .QN(n1923) );
  DFFRX1 \I_cache/cache_reg[7][18]  ( .D(n12636), .CK(clk), .RN(n5907), .Q(
        \I_cache/cache[7][18] ), .QN(n3577) );
  DFFRX1 \I_cache/cache_reg[0][19]  ( .D(n12635), .CK(clk), .RN(n5907), .Q(
        \I_cache/cache[0][19] ), .QN(n1864) );
  DFFRX1 \I_cache/cache_reg[1][19]  ( .D(n12634), .CK(clk), .RN(n5907), .Q(
        \I_cache/cache[1][19] ), .QN(n3520) );
  DFFRX1 \I_cache/cache_reg[2][19]  ( .D(n12633), .CK(clk), .RN(n5907), .Q(
        \I_cache/cache[2][19] ), .QN(n1866) );
  DFFRX1 \I_cache/cache_reg[3][19]  ( .D(n12632), .CK(clk), .RN(n5906), .Q(
        \I_cache/cache[3][19] ), .QN(n3522) );
  DFFRX1 \I_cache/cache_reg[4][19]  ( .D(n12631), .CK(clk), .RN(n5906), .Q(
        \I_cache/cache[4][19] ), .QN(n1865) );
  DFFRX1 \I_cache/cache_reg[5][19]  ( .D(n12630), .CK(clk), .RN(n5906), .Q(
        \I_cache/cache[5][19] ), .QN(n3521) );
  DFFRX1 \I_cache/cache_reg[6][19]  ( .D(n12629), .CK(clk), .RN(n5906), .Q(
        \I_cache/cache[6][19] ), .QN(n1869) );
  DFFRX1 \I_cache/cache_reg[7][19]  ( .D(n12628), .CK(clk), .RN(n5906), .Q(
        \I_cache/cache[7][19] ), .QN(n3525) );
  DFFRX1 \I_cache/cache_reg[0][20]  ( .D(n12627), .CK(clk), .RN(n5906), .Q(
        \I_cache/cache[0][20] ), .QN(n1879) );
  DFFRX1 \I_cache/cache_reg[1][20]  ( .D(n12626), .CK(clk), .RN(n5906), .Q(
        \I_cache/cache[1][20] ), .QN(n3534) );
  DFFRX1 \I_cache/cache_reg[2][20]  ( .D(n12625), .CK(clk), .RN(n5911), .Q(
        \I_cache/cache[2][20] ), .QN(n1881) );
  DFFRX1 \I_cache/cache_reg[3][20]  ( .D(n12624), .CK(clk), .RN(n5926), .Q(
        \I_cache/cache[3][20] ), .QN(n3536) );
  DFFRX1 \I_cache/cache_reg[4][20]  ( .D(n12623), .CK(clk), .RN(n5926), .Q(
        \I_cache/cache[4][20] ), .QN(n1880) );
  DFFRX1 \I_cache/cache_reg[5][20]  ( .D(n12622), .CK(clk), .RN(n5926), .Q(
        \I_cache/cache[5][20] ), .QN(n3535) );
  DFFRX1 \I_cache/cache_reg[6][20]  ( .D(n12621), .CK(clk), .RN(n5926), .Q(
        \I_cache/cache[6][20] ), .QN(n1917) );
  DFFRX1 \I_cache/cache_reg[7][20]  ( .D(n12620), .CK(clk), .RN(n5925), .Q(
        \I_cache/cache[7][20] ), .QN(n3571) );
  DFFRX1 \I_cache/cache_reg[0][21]  ( .D(n12619), .CK(clk), .RN(n5925), .Q(
        \I_cache/cache[0][21] ), .QN(n1793) );
  DFFRX1 \I_cache/cache_reg[1][21]  ( .D(n12618), .CK(clk), .RN(n5925), .Q(
        \I_cache/cache[1][21] ), .QN(n3449) );
  DFFRX1 \I_cache/cache_reg[2][21]  ( .D(n12617), .CK(clk), .RN(n5925), .Q(
        \I_cache/cache[2][21] ), .QN(n1822) );
  DFFRX1 \I_cache/cache_reg[3][21]  ( .D(n12616), .CK(clk), .RN(n5925), .Q(
        \I_cache/cache[3][21] ), .QN(n3478) );
  DFFRX1 \I_cache/cache_reg[4][21]  ( .D(n12615), .CK(clk), .RN(n5925), .Q(
        \I_cache/cache[4][21] ), .QN(n1821) );
  DFFRX1 \I_cache/cache_reg[5][21]  ( .D(n12614), .CK(clk), .RN(n5925), .Q(
        \I_cache/cache[5][21] ), .QN(n3477) );
  DFFRX1 \I_cache/cache_reg[6][21]  ( .D(n12613), .CK(clk), .RN(n5925), .Q(
        \I_cache/cache[6][21] ), .QN(n1845) );
  DFFRX1 \I_cache/cache_reg[7][21]  ( .D(n12612), .CK(clk), .RN(n5925), .Q(
        \I_cache/cache[7][21] ), .QN(n3501) );
  DFFRX1 \I_cache/cache_reg[7][22]  ( .D(n12604), .CK(clk), .RN(n5924), .Q(
        \I_cache/cache[7][22] ), .QN(n1915) );
  DFFRX1 \I_cache/cache_reg[0][23]  ( .D(n12603), .CK(clk), .RN(n5924), .Q(
        \I_cache/cache[0][23] ), .QN(n1790) );
  DFFRX1 \I_cache/cache_reg[1][23]  ( .D(n12602), .CK(clk), .RN(n5924), .Q(
        \I_cache/cache[1][23] ), .QN(n3446) );
  DFFRX1 \I_cache/cache_reg[2][23]  ( .D(n12601), .CK(clk), .RN(n5924), .Q(
        \I_cache/cache[2][23] ), .QN(n1809) );
  DFFRX1 \I_cache/cache_reg[3][23]  ( .D(n12600), .CK(clk), .RN(n5924), .Q(
        \I_cache/cache[3][23] ), .QN(n3465) );
  DFFRX1 \I_cache/cache_reg[4][23]  ( .D(n12599), .CK(clk), .RN(n5924), .Q(
        \I_cache/cache[4][23] ), .QN(n1808) );
  DFFRX1 \I_cache/cache_reg[5][23]  ( .D(n12598), .CK(clk), .RN(n5924), .Q(
        \I_cache/cache[5][23] ), .QN(n3464) );
  DFFRX1 \I_cache/cache_reg[6][23]  ( .D(n12597), .CK(clk), .RN(n5924), .Q(
        \I_cache/cache[6][23] ), .QN(n1838) );
  DFFRX1 \I_cache/cache_reg[7][23]  ( .D(n12596), .CK(clk), .RN(n5923), .Q(
        \I_cache/cache[7][23] ), .QN(n3494) );
  DFFRX1 \I_cache/cache_reg[0][24]  ( .D(n12595), .CK(clk), .RN(n5923), .Q(
        \I_cache/cache[0][24] ), .QN(n1871) );
  DFFRX1 \I_cache/cache_reg[1][24]  ( .D(n12594), .CK(clk), .RN(n5923), .Q(
        \I_cache/cache[1][24] ), .QN(n3527) );
  DFFRX1 \I_cache/cache_reg[2][24]  ( .D(n12593), .CK(clk), .RN(n5923), .Q(
        \I_cache/cache[2][24] ), .QN(n1872) );
  DFFRX1 \I_cache/cache_reg[3][24]  ( .D(n12592), .CK(clk), .RN(n5923), .Q(
        \I_cache/cache[3][24] ), .QN(n3528) );
  DFFRX1 \I_cache/cache_reg[4][24]  ( .D(n12591), .CK(clk), .RN(n5923), .Q(
        \I_cache/cache[4][24] ), .QN(n1867) );
  DFFRX1 \I_cache/cache_reg[5][24]  ( .D(n12590), .CK(clk), .RN(n5923), .Q(
        \I_cache/cache[5][24] ), .QN(n3523) );
  DFFRX1 \I_cache/cache_reg[6][24]  ( .D(n12589), .CK(clk), .RN(n5923), .Q(
        \I_cache/cache[6][24] ), .QN(n1913) );
  DFFRX1 \I_cache/cache_reg[7][24]  ( .D(n12588), .CK(clk), .RN(n5923), .Q(
        \I_cache/cache[7][24] ), .QN(n3568) );
  DFFRX1 \I_cache/cache_reg[0][25]  ( .D(n12587), .CK(clk), .RN(n5923), .Q(
        \I_cache/cache[0][25] ), .QN(n1787) );
  DFFRX1 \I_cache/cache_reg[1][25]  ( .D(n12586), .CK(clk), .RN(n5923), .Q(
        \I_cache/cache[1][25] ), .QN(n3443) );
  DFFRX1 \I_cache/cache_reg[2][25]  ( .D(n12585), .CK(clk), .RN(n5923), .Q(
        \I_cache/cache[2][25] ), .QN(n1797) );
  DFFRX1 \I_cache/cache_reg[3][25]  ( .D(n12584), .CK(clk), .RN(n5922), .Q(
        \I_cache/cache[3][25] ), .QN(n3453) );
  DFFRX1 \I_cache/cache_reg[4][25]  ( .D(n12583), .CK(clk), .RN(n5922), .Q(
        \I_cache/cache[4][25] ), .QN(n1796) );
  DFFRX1 \I_cache/cache_reg[5][25]  ( .D(n12582), .CK(clk), .RN(n5922), .Q(
        \I_cache/cache[5][25] ), .QN(n3452) );
  DFFRX1 \I_cache/cache_reg[6][25]  ( .D(n12581), .CK(clk), .RN(n5922), .Q(
        \I_cache/cache[6][25] ), .QN(n1832) );
  DFFRX1 \I_cache/cache_reg[7][25]  ( .D(n12580), .CK(clk), .RN(n5922), .Q(
        \I_cache/cache[7][25] ), .QN(n3488) );
  DFFRX1 \I_cache/cache_reg[0][26]  ( .D(n12579), .CK(clk), .RN(n5922), .Q(
        \I_cache/cache[0][26] ), .QN(n1559) );
  DFFRX1 \I_cache/cache_reg[1][26]  ( .D(n12578), .CK(clk), .RN(n5922), .Q(
        \I_cache/cache[1][26] ), .QN(n3142) );
  DFFRX1 \I_cache/cache_reg[2][26]  ( .D(n12577), .CK(clk), .RN(n5922), .Q(
        \I_cache/cache[2][26] ), .QN(n1455) );
  DFFRX1 \I_cache/cache_reg[3][26]  ( .D(n12576), .CK(clk), .RN(n5922), .Q(
        \I_cache/cache[3][26] ), .QN(n3141) );
  DFFRX1 \I_cache/cache_reg[4][26]  ( .D(n12575), .CK(clk), .RN(n5922), .Q(
        \I_cache/cache[4][26] ), .QN(n1571) );
  DFFRX1 \I_cache/cache_reg[5][26]  ( .D(n12574), .CK(clk), .RN(n5922), .Q(
        \I_cache/cache[5][26] ), .QN(n3153) );
  DFFRX1 \I_cache/cache_reg[6][26]  ( .D(n12573), .CK(clk), .RN(n5922), .Q(
        \I_cache/cache[6][26] ), .QN(n1560) );
  DFFRX1 \I_cache/cache_reg[7][26]  ( .D(n12572), .CK(clk), .RN(n5921), .Q(
        \I_cache/cache[7][26] ), .QN(n3143) );
  DFFRX1 \I_cache/cache_reg[0][27]  ( .D(n12571), .CK(clk), .RN(n5921), .Q(
        \I_cache/cache[0][27] ), .QN(n1536) );
  DFFRX1 \I_cache/cache_reg[1][27]  ( .D(n12570), .CK(clk), .RN(n5921), .Q(
        \I_cache/cache[1][27] ), .QN(n3118) );
  DFFRX1 \I_cache/cache_reg[2][27]  ( .D(n12569), .CK(clk), .RN(n5921), .Q(
        \I_cache/cache[2][27] ), .QN(n1535) );
  DFFRX1 \I_cache/cache_reg[3][27]  ( .D(n12568), .CK(clk), .RN(n5921), .Q(
        \I_cache/cache[3][27] ), .QN(n3117) );
  DFFRX1 \I_cache/cache_reg[4][27]  ( .D(n12567), .CK(clk), .RN(n5921), .Q(
        \I_cache/cache[4][27] ), .QN(n1604) );
  DFFRX1 \I_cache/cache_reg[5][27]  ( .D(n12566), .CK(clk), .RN(n5921), .Q(
        \I_cache/cache[5][27] ), .QN(n3181) );
  DFFRX1 \I_cache/cache_reg[6][27]  ( .D(n12565), .CK(clk), .RN(n5921), .Q(
        \I_cache/cache[6][27] ), .QN(n1537) );
  DFFRX1 \I_cache/cache_reg[7][27]  ( .D(n12564), .CK(clk), .RN(n5921), .Q(
        \I_cache/cache[7][27] ), .QN(n3119) );
  DFFRX1 \I_cache/cache_reg[0][31]  ( .D(n12539), .CK(clk), .RN(n5919), .Q(
        \I_cache/cache[0][31] ), .QN(n1548) );
  DFFRX1 \I_cache/cache_reg[1][31]  ( .D(n12538), .CK(clk), .RN(n5919), .Q(
        \I_cache/cache[1][31] ), .QN(n3130) );
  DFFRX1 \I_cache/cache_reg[2][31]  ( .D(n12537), .CK(clk), .RN(n5918), .Q(
        \I_cache/cache[2][31] ), .QN(n1547) );
  DFFRX1 \I_cache/cache_reg[3][31]  ( .D(n12536), .CK(clk), .RN(n5918), .Q(
        \I_cache/cache[3][31] ), .QN(n3129) );
  DFFRX1 \I_cache/cache_reg[4][31]  ( .D(n12535), .CK(clk), .RN(n5918), .Q(
        \I_cache/cache[4][31] ), .QN(n1605) );
  DFFRX1 \I_cache/cache_reg[6][31]  ( .D(n12533), .CK(clk), .RN(n5918), .Q(
        \I_cache/cache[6][31] ), .QN(n1549) );
  DFFRX1 \I_cache/cache_reg[0][48]  ( .D(n12403), .CK(clk), .RN(n5808), .Q(
        \I_cache/cache[0][48] ), .QN(n1911) );
  DFFRX1 \I_cache/cache_reg[1][48]  ( .D(n12402), .CK(clk), .RN(n5808), .Q(
        \I_cache/cache[1][48] ), .QN(n3566) );
  DFFRX1 \I_cache/cache_reg[2][48]  ( .D(n12401), .CK(clk), .RN(n5807), .Q(
        \I_cache/cache[2][48] ), .QN(n1912) );
  DFFRX1 \I_cache/cache_reg[3][48]  ( .D(n12400), .CK(clk), .RN(n5807), .Q(
        \I_cache/cache[3][48] ), .QN(n3567) );
  DFFRX1 \I_cache/cache_reg[4][48]  ( .D(n12399), .CK(clk), .RN(n5807), .Q(
        \I_cache/cache[4][48] ), .QN(n1850) );
  DFFRX1 \I_cache/cache_reg[5][48]  ( .D(n12398), .CK(clk), .RN(n5807), .Q(
        \I_cache/cache[5][48] ), .QN(n3506) );
  DFFRX1 \I_cache/cache_reg[6][48]  ( .D(n12397), .CK(clk), .RN(n5807), .Q(
        \I_cache/cache[6][48] ), .QN(n1933) );
  DFFRX1 \I_cache/cache_reg[7][48]  ( .D(n12396), .CK(clk), .RN(n5807), .Q(
        \I_cache/cache[7][48] ), .QN(n3587) );
  DFFRX1 \I_cache/cache_reg[0][49]  ( .D(n12395), .CK(clk), .RN(n5807), .Q(
        \I_cache/cache[0][49] ), .QN(n1903) );
  DFFRX1 \I_cache/cache_reg[1][49]  ( .D(n12394), .CK(clk), .RN(n5807), .Q(
        \I_cache/cache[1][49] ), .QN(n3558) );
  DFFRX1 \I_cache/cache_reg[2][49]  ( .D(n12393), .CK(clk), .RN(n5807), .Q(
        \I_cache/cache[2][49] ), .QN(n1904) );
  DFFRX1 \I_cache/cache_reg[3][49]  ( .D(n12392), .CK(clk), .RN(n5807), .Q(
        \I_cache/cache[3][49] ), .QN(n3559) );
  DFFRX1 \I_cache/cache_reg[4][49]  ( .D(n12391), .CK(clk), .RN(n5807), .Q(
        \I_cache/cache[4][49] ), .QN(n1830) );
  DFFRX1 \I_cache/cache_reg[5][49]  ( .D(n12390), .CK(clk), .RN(n5807), .Q(
        \I_cache/cache[5][49] ), .QN(n3486) );
  DFFRX1 \I_cache/cache_reg[6][49]  ( .D(n12389), .CK(clk), .RN(n5806), .Q(
        \I_cache/cache[6][49] ), .QN(n1929) );
  DFFRX1 \I_cache/cache_reg[7][49]  ( .D(n12388), .CK(clk), .RN(n5806), .Q(
        \I_cache/cache[7][49] ), .QN(n3583) );
  DFFRX1 \I_cache/cache_reg[0][50]  ( .D(n12387), .CK(clk), .RN(n5806), .Q(
        \I_cache/cache[0][50] ), .QN(n1895) );
  DFFRX1 \I_cache/cache_reg[1][50]  ( .D(n12386), .CK(clk), .RN(n5806), .Q(
        \I_cache/cache[1][50] ), .QN(n3550) );
  DFFRX1 \I_cache/cache_reg[2][50]  ( .D(n12385), .CK(clk), .RN(n5811), .Q(
        \I_cache/cache[2][50] ), .QN(n1827) );
  DFFRX1 \I_cache/cache_reg[3][50]  ( .D(n12384), .CK(clk), .RN(n5826), .Q(
        \I_cache/cache[3][50] ), .QN(n3483) );
  DFFRX1 \I_cache/cache_reg[4][50]  ( .D(n12383), .CK(clk), .RN(n5826), .Q(
        \I_cache/cache[4][50] ), .QN(n1852) );
  DFFRX1 \I_cache/cache_reg[5][50]  ( .D(n12382), .CK(clk), .RN(n5826), .Q(
        \I_cache/cache[5][50] ), .QN(n3508) );
  DFFRX1 \I_cache/cache_reg[6][50]  ( .D(n12381), .CK(clk), .RN(n5826), .Q(
        \I_cache/cache[6][50] ), .QN(n1925) );
  DFFRX1 \I_cache/cache_reg[7][50]  ( .D(n12380), .CK(clk), .RN(n5826), .Q(
        \I_cache/cache[7][50] ), .QN(n3579) );
  DFFRX1 \I_cache/cache_reg[0][51]  ( .D(n12379), .CK(clk), .RN(n5826), .Q(
        \I_cache/cache[0][51] ), .QN(n1854) );
  DFFRX1 \I_cache/cache_reg[1][51]  ( .D(n12378), .CK(clk), .RN(n5825), .Q(
        \I_cache/cache[1][51] ), .QN(n3510) );
  DFFRX1 \I_cache/cache_reg[2][51]  ( .D(n12377), .CK(clk), .RN(n5825), .Q(
        \I_cache/cache[2][51] ), .QN(n1856) );
  DFFRX1 \I_cache/cache_reg[3][51]  ( .D(n12376), .CK(clk), .RN(n5825), .Q(
        \I_cache/cache[3][51] ), .QN(n3512) );
  DFFRX1 \I_cache/cache_reg[4][51]  ( .D(n12375), .CK(clk), .RN(n5825), .Q(
        \I_cache/cache[4][51] ), .QN(n1855) );
  DFFRX1 \I_cache/cache_reg[5][51]  ( .D(n12374), .CK(clk), .RN(n5825), .Q(
        \I_cache/cache[5][51] ), .QN(n3511) );
  DFFRX1 \I_cache/cache_reg[6][51]  ( .D(n12373), .CK(clk), .RN(n5825), .Q(
        \I_cache/cache[6][51] ), .QN(n1870) );
  DFFRX1 \I_cache/cache_reg[7][51]  ( .D(n12372), .CK(clk), .RN(n5825), .Q(
        \I_cache/cache[7][51] ), .QN(n3526) );
  DFFRX1 \I_cache/cache_reg[0][52]  ( .D(n12371), .CK(clk), .RN(n5825), .Q(
        \I_cache/cache[0][52] ), .QN(n1885) );
  DFFRX1 \I_cache/cache_reg[1][52]  ( .D(n12370), .CK(clk), .RN(n5825), .Q(
        \I_cache/cache[1][52] ), .QN(n3540) );
  DFFRX1 \I_cache/cache_reg[2][52]  ( .D(n12369), .CK(clk), .RN(n5825), .Q(
        \I_cache/cache[2][52] ), .QN(n1887) );
  DFFRX1 \I_cache/cache_reg[3][52]  ( .D(n12368), .CK(clk), .RN(n5825), .Q(
        \I_cache/cache[3][52] ), .QN(n3542) );
  DFFRX1 \I_cache/cache_reg[4][52]  ( .D(n12367), .CK(clk), .RN(n5825), .Q(
        \I_cache/cache[4][52] ), .QN(n1886) );
  DFFRX1 \I_cache/cache_reg[5][52]  ( .D(n12366), .CK(clk), .RN(n5824), .Q(
        \I_cache/cache[5][52] ), .QN(n3541) );
  DFFRX1 \I_cache/cache_reg[6][52]  ( .D(n12365), .CK(clk), .RN(n5824), .Q(
        \I_cache/cache[6][52] ), .QN(n1919) );
  DFFRX1 \I_cache/cache_reg[7][52]  ( .D(n12364), .CK(clk), .RN(n5824), .Q(
        \I_cache/cache[7][52] ), .QN(n3573) );
  DFFRX1 \I_cache/cache_reg[0][53]  ( .D(n12363), .CK(clk), .RN(n5824), .Q(
        \I_cache/cache[0][53] ), .QN(n1785) );
  DFFRX1 \I_cache/cache_reg[1][53]  ( .D(n12362), .CK(clk), .RN(n5824), .Q(
        \I_cache/cache[1][53] ), .QN(n3441) );
  DFFRX1 \I_cache/cache_reg[2][53]  ( .D(n12361), .CK(clk), .RN(n5824), .Q(
        \I_cache/cache[2][53] ), .QN(n1826) );
  DFFRX1 \I_cache/cache_reg[3][53]  ( .D(n12360), .CK(clk), .RN(n5824), .Q(
        \I_cache/cache[3][53] ), .QN(n3482) );
  DFFRX1 \I_cache/cache_reg[4][53]  ( .D(n12359), .CK(clk), .RN(n5824), .Q(
        \I_cache/cache[4][53] ), .QN(n1825) );
  DFFRX1 \I_cache/cache_reg[5][53]  ( .D(n12358), .CK(clk), .RN(n5824), .Q(
        \I_cache/cache[5][53] ), .QN(n3481) );
  DFFRX1 \I_cache/cache_reg[6][53]  ( .D(n12357), .CK(clk), .RN(n5824), .Q(
        \I_cache/cache[6][53] ), .QN(n1847) );
  DFFRX1 \I_cache/cache_reg[7][53]  ( .D(n12356), .CK(clk), .RN(n5824), .Q(
        \I_cache/cache[7][53] ), .QN(n3503) );
  DFFRX1 \I_cache/cache_reg[0][54]  ( .D(n12355), .CK(clk), .RN(n5824), .Q(
        \I_cache/cache[0][54] ), .QN(n1783) );
  DFFRX1 \I_cache/cache_reg[1][54]  ( .D(n12354), .CK(clk), .RN(n5823), .Q(
        \I_cache/cache[1][54] ), .QN(n3439) );
  DFFRX1 \I_cache/cache_reg[2][54]  ( .D(n12353), .CK(clk), .RN(n5823), .Q(
        \I_cache/cache[2][54] ), .QN(n1818) );
  DFFRX1 \I_cache/cache_reg[3][54]  ( .D(n12352), .CK(clk), .RN(n5823), .Q(
        \I_cache/cache[3][54] ), .QN(n3474) );
  DFFRX1 \I_cache/cache_reg[4][54]  ( .D(n12351), .CK(clk), .RN(n5823), .Q(
        \I_cache/cache[4][54] ), .QN(n1817) );
  DFFRX1 \I_cache/cache_reg[5][54]  ( .D(n12350), .CK(clk), .RN(n5823), .Q(
        \I_cache/cache[5][54] ), .QN(n3473) );
  DFFRX1 \I_cache/cache_reg[6][54]  ( .D(n12349), .CK(clk), .RN(n5823), .Q(
        \I_cache/cache[6][54] ), .QN(n1843) );
  DFFRX1 \I_cache/cache_reg[7][54]  ( .D(n12348), .CK(clk), .RN(n5823), .Q(
        \I_cache/cache[7][54] ), .QN(n3499) );
  DFFRX1 \I_cache/cache_reg[0][55]  ( .D(n12347), .CK(clk), .RN(n5823), .Q(
        \I_cache/cache[0][55] ), .QN(n1781) );
  DFFRX1 \I_cache/cache_reg[1][55]  ( .D(n12346), .CK(clk), .RN(n5823), .Q(
        \I_cache/cache[1][55] ), .QN(n3437) );
  DFFRX1 \I_cache/cache_reg[2][55]  ( .D(n12345), .CK(clk), .RN(n5823), .Q(
        \I_cache/cache[2][55] ), .QN(n1813) );
  DFFRX1 \I_cache/cache_reg[3][55]  ( .D(n12344), .CK(clk), .RN(n5823), .Q(
        \I_cache/cache[3][55] ), .QN(n3469) );
  DFFRX1 \I_cache/cache_reg[4][55]  ( .D(n12343), .CK(clk), .RN(n5823), .Q(
        \I_cache/cache[4][55] ), .QN(n1812) );
  DFFRX1 \I_cache/cache_reg[5][55]  ( .D(n12342), .CK(clk), .RN(n5822), .Q(
        \I_cache/cache[5][55] ), .QN(n3468) );
  DFFRX1 \I_cache/cache_reg[6][55]  ( .D(n12341), .CK(clk), .RN(n5822), .Q(
        \I_cache/cache[6][55] ), .QN(n1840) );
  DFFRX1 \I_cache/cache_reg[7][55]  ( .D(n12340), .CK(clk), .RN(n5822), .Q(
        \I_cache/cache[7][55] ), .QN(n3496) );
  DFFRX1 \I_cache/cache_reg[0][56]  ( .D(n12339), .CK(clk), .RN(n5822), .Q(
        \I_cache/cache[0][56] ), .QN(n1873) );
  DFFRX1 \I_cache/cache_reg[1][56]  ( .D(n12338), .CK(clk), .RN(n5822), .Q(
        \I_cache/cache[1][56] ), .QN(n3529) );
  DFFRX1 \I_cache/cache_reg[2][56]  ( .D(n12337), .CK(clk), .RN(n5822), .Q(
        \I_cache/cache[2][56] ), .QN(n1874) );
  DFFRX1 \I_cache/cache_reg[3][56]  ( .D(n12336), .CK(clk), .RN(n5822), .Q(
        \I_cache/cache[3][56] ), .QN(n3530) );
  DFFRX1 \I_cache/cache_reg[4][56]  ( .D(n12335), .CK(clk), .RN(n5822), .Q(
        \I_cache/cache[4][56] ), .QN(n1857) );
  DFFRX1 \I_cache/cache_reg[5][56]  ( .D(n12334), .CK(clk), .RN(n5822), .Q(
        \I_cache/cache[5][56] ), .QN(n3513) );
  DFFRX1 \I_cache/cache_reg[6][56]  ( .D(n12333), .CK(clk), .RN(n5822), .Q(
        \I_cache/cache[6][56] ), .QN(n1914) );
  DFFRX1 \I_cache/cache_reg[7][56]  ( .D(n12332), .CK(clk), .RN(n5822), .Q(
        \I_cache/cache[7][56] ), .QN(n3569) );
  DFFRX1 \I_cache/cache_reg[0][57]  ( .D(n12331), .CK(clk), .RN(n5822), .Q(
        \I_cache/cache[0][57] ), .QN(n1778) );
  DFFRX1 \I_cache/cache_reg[1][57]  ( .D(n12330), .CK(clk), .RN(n5821), .Q(
        \I_cache/cache[1][57] ), .QN(n3434) );
  DFFRX1 \I_cache/cache_reg[2][57]  ( .D(n12329), .CK(clk), .RN(n5821), .Q(
        \I_cache/cache[2][57] ), .QN(n1801) );
  DFFRX1 \I_cache/cache_reg[3][57]  ( .D(n12328), .CK(clk), .RN(n5821), .Q(
        \I_cache/cache[3][57] ), .QN(n3457) );
  DFFRX1 \I_cache/cache_reg[4][57]  ( .D(n12327), .CK(clk), .RN(n5821), .Q(
        \I_cache/cache[4][57] ), .QN(n1800) );
  DFFRX1 \I_cache/cache_reg[5][57]  ( .D(n12326), .CK(clk), .RN(n5821), .Q(
        \I_cache/cache[5][57] ), .QN(n3456) );
  DFFRX1 \I_cache/cache_reg[6][57]  ( .D(n12325), .CK(clk), .RN(n5821), .Q(
        \I_cache/cache[6][57] ), .QN(n1834) );
  DFFRX1 \I_cache/cache_reg[7][57]  ( .D(n12324), .CK(clk), .RN(n5821), .Q(
        \I_cache/cache[7][57] ), .QN(n3490) );
  DFFRX1 \I_cache/cache_reg[0][58]  ( .D(n12323), .CK(clk), .RN(n5821), .Q(
        \I_cache/cache[0][58] ), .QN(n1565) );
  DFFRX1 \I_cache/cache_reg[1][58]  ( .D(n12322), .CK(clk), .RN(n5821), .Q(
        \I_cache/cache[1][58] ), .QN(n3148) );
  DFFRX1 \I_cache/cache_reg[2][58]  ( .D(n12321), .CK(clk), .RN(n5821), .Q(
        \I_cache/cache[2][58] ), .QN(n1564) );
  DFFRX1 \I_cache/cache_reg[3][58]  ( .D(n12320), .CK(clk), .RN(n5821), .Q(
        \I_cache/cache[3][58] ), .QN(n3147) );
  DFFRX1 \I_cache/cache_reg[4][58]  ( .D(n12319), .CK(clk), .RN(n5820), .Q(
        \I_cache/cache[4][58] ), .QN(n1573) );
  DFFRX1 \I_cache/cache_reg[5][58]  ( .D(n12318), .CK(clk), .RN(n5820), .Q(
        \I_cache/cache[5][58] ), .QN(n3155) );
  DFFRX1 \I_cache/cache_reg[6][58]  ( .D(n12317), .CK(clk), .RN(n5820), .Q(
        \I_cache/cache[6][58] ), .QN(n1566) );
  DFFRX1 \I_cache/cache_reg[7][58]  ( .D(n12316), .CK(clk), .RN(n5820), .Q(
        \I_cache/cache[7][58] ), .QN(n3149) );
  DFFRX1 \I_cache/cache_reg[0][59]  ( .D(n12315), .CK(clk), .RN(n5820), .Q(
        \I_cache/cache[0][59] ), .QN(n1542) );
  DFFRX1 \I_cache/cache_reg[1][59]  ( .D(n12314), .CK(clk), .RN(n5820), .Q(
        \I_cache/cache[1][59] ), .QN(n3124) );
  DFFRX1 \I_cache/cache_reg[2][59]  ( .D(n12313), .CK(clk), .RN(n5820), .Q(
        \I_cache/cache[2][59] ), .QN(n1541) );
  DFFRX1 \I_cache/cache_reg[3][59]  ( .D(n12312), .CK(clk), .RN(n5820), .Q(
        \I_cache/cache[3][59] ), .QN(n3123) );
  DFFRX1 \I_cache/cache_reg[4][59]  ( .D(n12311), .CK(clk), .RN(n5820), .Q(
        \I_cache/cache[4][59] ), .QN(n1608) );
  DFFRX1 \I_cache/cache_reg[5][59]  ( .D(n12310), .CK(clk), .RN(n5820), .Q(
        \I_cache/cache[5][59] ), .QN(n3185) );
  DFFRX1 \I_cache/cache_reg[6][59]  ( .D(n12309), .CK(clk), .RN(n5820), .Q(
        \I_cache/cache[6][59] ), .QN(n1543) );
  DFFRX1 \I_cache/cache_reg[7][59]  ( .D(n12308), .CK(clk), .RN(n5820), .Q(
        \I_cache/cache[7][59] ), .QN(n3125) );
  DFFRX1 \I_cache/cache_reg[0][63]  ( .D(n12283), .CK(clk), .RN(n5817), .Q(
        \I_cache/cache[0][63] ), .QN(n1554) );
  DFFRX1 \I_cache/cache_reg[1][63]  ( .D(n12282), .CK(clk), .RN(n5817), .Q(
        \I_cache/cache[1][63] ), .QN(n3136) );
  DFFRX1 \I_cache/cache_reg[2][63]  ( .D(n12281), .CK(clk), .RN(n5817), .Q(
        \I_cache/cache[2][63] ), .QN(n1553) );
  DFFRX1 \I_cache/cache_reg[4][63]  ( .D(n12279), .CK(clk), .RN(n5817), .Q(
        \I_cache/cache[4][63] ), .QN(n1603) );
  DFFRX1 \I_cache/cache_reg[6][63]  ( .D(n12277), .CK(clk), .RN(n5817), .Q(
        \I_cache/cache[6][63] ), .QN(n1555) );
  DFFRX1 \I_cache/cache_reg[0][80]  ( .D(n12147), .CK(clk), .RN(n5791), .Q(
        \I_cache/cache[0][80] ), .QN(n1909) );
  DFFRX1 \I_cache/cache_reg[1][80]  ( .D(n12146), .CK(clk), .RN(n5806), .Q(
        \I_cache/cache[1][80] ), .QN(n3564) );
  DFFRX1 \I_cache/cache_reg[2][80]  ( .D(n12145), .CK(clk), .RN(n5806), .Q(
        \I_cache/cache[2][80] ), .QN(n1910) );
  DFFRX1 \I_cache/cache_reg[3][80]  ( .D(n12144), .CK(clk), .RN(n5806), .Q(
        \I_cache/cache[3][80] ), .QN(n3565) );
  DFFRX1 \I_cache/cache_reg[4][80]  ( .D(n12143), .CK(clk), .RN(n5806), .Q(
        \I_cache/cache[4][80] ), .QN(n1858) );
  DFFRX1 \I_cache/cache_reg[5][80]  ( .D(n12142), .CK(clk), .RN(n5806), .Q(
        \I_cache/cache[5][80] ), .QN(n3514) );
  DFFRX1 \I_cache/cache_reg[6][80]  ( .D(n12141), .CK(clk), .RN(n5806), .Q(
        \I_cache/cache[6][80] ), .QN(n1932) );
  DFFRX1 \I_cache/cache_reg[7][80]  ( .D(n12140), .CK(clk), .RN(n5806), .Q(
        \I_cache/cache[7][80] ), .QN(n3586) );
  DFFRX1 \I_cache/cache_reg[0][81]  ( .D(n12139), .CK(clk), .RN(n5805), .Q(
        \I_cache/cache[0][81] ), .QN(n1900) );
  DFFRX1 \I_cache/cache_reg[1][81]  ( .D(n12138), .CK(clk), .RN(n5805), .Q(
        \I_cache/cache[1][81] ), .QN(n3555) );
  DFFRX1 \I_cache/cache_reg[2][81]  ( .D(n12137), .CK(clk), .RN(n5805), .Q(
        \I_cache/cache[2][81] ), .QN(n1902) );
  DFFRX1 \I_cache/cache_reg[3][81]  ( .D(n12136), .CK(clk), .RN(n5805), .Q(
        \I_cache/cache[3][81] ), .QN(n3557) );
  DFFRX1 \I_cache/cache_reg[4][81]  ( .D(n12135), .CK(clk), .RN(n5805), .Q(
        \I_cache/cache[4][81] ), .QN(n1901) );
  DFFRX1 \I_cache/cache_reg[5][81]  ( .D(n12134), .CK(clk), .RN(n5805), .Q(
        \I_cache/cache[5][81] ), .QN(n3556) );
  DFFRX1 \I_cache/cache_reg[6][81]  ( .D(n12133), .CK(clk), .RN(n5805), .Q(
        \I_cache/cache[6][81] ), .QN(n1928) );
  DFFRX1 \I_cache/cache_reg[7][81]  ( .D(n12132), .CK(clk), .RN(n5805), .Q(
        \I_cache/cache[7][81] ), .QN(n3582) );
  DFFRX1 \I_cache/cache_reg[0][82]  ( .D(n12131), .CK(clk), .RN(n5805), .Q(
        \I_cache/cache[0][82] ), .QN(n1894) );
  DFFRX1 \I_cache/cache_reg[1][82]  ( .D(n12130), .CK(clk), .RN(n5805), .Q(
        \I_cache/cache[1][82] ), .QN(n3549) );
  DFFRX1 \I_cache/cache_reg[2][82]  ( .D(n12129), .CK(clk), .RN(n5805), .Q(
        \I_cache/cache[2][82] ), .QN(n1848) );
  DFFRX1 \I_cache/cache_reg[3][82]  ( .D(n12128), .CK(clk), .RN(n5805), .Q(
        \I_cache/cache[3][82] ), .QN(n3504) );
  DFFRX1 \I_cache/cache_reg[4][82]  ( .D(n12127), .CK(clk), .RN(n5804), .Q(
        \I_cache/cache[4][82] ), .QN(n1851) );
  DFFRX1 \I_cache/cache_reg[5][82]  ( .D(n12126), .CK(clk), .RN(n5804), .Q(
        \I_cache/cache[5][82] ), .QN(n3507) );
  DFFRX1 \I_cache/cache_reg[6][82]  ( .D(n12125), .CK(clk), .RN(n5804), .Q(
        \I_cache/cache[6][82] ), .QN(n1924) );
  DFFRX1 \I_cache/cache_reg[7][82]  ( .D(n12124), .CK(clk), .RN(n5804), .Q(
        \I_cache/cache[7][82] ), .QN(n3578) );
  DFFRX1 \I_cache/cache_reg[0][83]  ( .D(n12123), .CK(clk), .RN(n5804), .Q(
        \I_cache/cache[0][83] ), .QN(n1890) );
  DFFRX1 \I_cache/cache_reg[1][83]  ( .D(n12122), .CK(clk), .RN(n5804), .Q(
        \I_cache/cache[1][83] ), .QN(n3545) );
  DFFRX1 \I_cache/cache_reg[2][83]  ( .D(n12121), .CK(clk), .RN(n5804), .Q(
        \I_cache/cache[2][83] ), .QN(n1891) );
  DFFRX1 \I_cache/cache_reg[3][83]  ( .D(n12120), .CK(clk), .RN(n5804), .Q(
        \I_cache/cache[3][83] ), .QN(n3546) );
  DFFRX1 \I_cache/cache_reg[4][83]  ( .D(n12119), .CK(clk), .RN(n5804), .Q(
        \I_cache/cache[4][83] ), .QN(n1853) );
  DFFRX1 \I_cache/cache_reg[5][83]  ( .D(n12118), .CK(clk), .RN(n5804), .Q(
        \I_cache/cache[5][83] ), .QN(n3509) );
  DFFRX1 \I_cache/cache_reg[6][83]  ( .D(n12117), .CK(clk), .RN(n5804), .Q(
        \I_cache/cache[6][83] ), .QN(n1921) );
  DFFRX1 \I_cache/cache_reg[7][83]  ( .D(n12116), .CK(clk), .RN(n5804), .Q(
        \I_cache/cache[7][83] ), .QN(n3575) );
  DFFRX1 \I_cache/cache_reg[0][84]  ( .D(n12115), .CK(clk), .RN(n5803), .Q(
        \I_cache/cache[0][84] ), .QN(n1882) );
  DFFRX1 \I_cache/cache_reg[1][84]  ( .D(n12114), .CK(clk), .RN(n5803), .Q(
        \I_cache/cache[1][84] ), .QN(n3537) );
  DFFRX1 \I_cache/cache_reg[2][84]  ( .D(n12113), .CK(clk), .RN(n5803), .Q(
        \I_cache/cache[2][84] ), .QN(n1884) );
  DFFRX1 \I_cache/cache_reg[3][84]  ( .D(n12112), .CK(clk), .RN(n5803), .Q(
        \I_cache/cache[3][84] ), .QN(n3539) );
  DFFRX1 \I_cache/cache_reg[4][84]  ( .D(n12111), .CK(clk), .RN(n5803), .Q(
        \I_cache/cache[4][84] ), .QN(n1883) );
  DFFRX1 \I_cache/cache_reg[5][84]  ( .D(n12110), .CK(clk), .RN(n5803), .Q(
        \I_cache/cache[5][84] ), .QN(n3538) );
  DFFRX1 \I_cache/cache_reg[6][84]  ( .D(n12109), .CK(clk), .RN(n5803), .Q(
        \I_cache/cache[6][84] ), .QN(n1918) );
  DFFRX1 \I_cache/cache_reg[7][84]  ( .D(n12108), .CK(clk), .RN(n5803), .Q(
        \I_cache/cache[7][84] ), .QN(n3572) );
  DFFRX1 \I_cache/cache_reg[0][85]  ( .D(n12107), .CK(clk), .RN(n5803), .Q(
        \I_cache/cache[0][85] ), .QN(n1784) );
  DFFRX1 \I_cache/cache_reg[1][85]  ( .D(n12106), .CK(clk), .RN(n5803), .Q(
        \I_cache/cache[1][85] ), .QN(n3440) );
  DFFRX1 \I_cache/cache_reg[2][85]  ( .D(n12105), .CK(clk), .RN(n5803), .Q(
        \I_cache/cache[2][85] ), .QN(n1824) );
  DFFRX1 \I_cache/cache_reg[3][85]  ( .D(n12104), .CK(clk), .RN(n5803), .Q(
        \I_cache/cache[3][85] ), .QN(n3480) );
  DFFRX1 \I_cache/cache_reg[4][85]  ( .D(n12103), .CK(clk), .RN(n5802), .Q(
        \I_cache/cache[4][85] ), .QN(n1823) );
  DFFRX1 \I_cache/cache_reg[5][85]  ( .D(n12102), .CK(clk), .RN(n5802), .Q(
        \I_cache/cache[5][85] ), .QN(n3479) );
  DFFRX1 \I_cache/cache_reg[6][85]  ( .D(n12101), .CK(clk), .RN(n5802), .Q(
        \I_cache/cache[6][85] ), .QN(n1846) );
  DFFRX1 \I_cache/cache_reg[7][85]  ( .D(n12100), .CK(clk), .RN(n5802), .Q(
        \I_cache/cache[7][85] ), .QN(n3502) );
  DFFRX1 \I_cache/cache_reg[0][86]  ( .D(n12099), .CK(clk), .RN(n5802), .Q(
        \I_cache/cache[0][86] ), .QN(n1782) );
  DFFRX1 \I_cache/cache_reg[1][86]  ( .D(n12098), .CK(clk), .RN(n5802), .Q(
        \I_cache/cache[1][86] ), .QN(n3438) );
  DFFRX1 \I_cache/cache_reg[2][86]  ( .D(n12097), .CK(clk), .RN(n5802), .Q(
        \I_cache/cache[2][86] ), .QN(n1816) );
  DFFRX1 \I_cache/cache_reg[3][86]  ( .D(n12096), .CK(clk), .RN(n5802), .Q(
        \I_cache/cache[3][86] ), .QN(n3472) );
  DFFRX1 \I_cache/cache_reg[4][86]  ( .D(n12095), .CK(clk), .RN(n5802), .Q(
        \I_cache/cache[4][86] ), .QN(n1815) );
  DFFRX1 \I_cache/cache_reg[5][86]  ( .D(n12094), .CK(clk), .RN(n5802), .Q(
        \I_cache/cache[5][86] ), .QN(n3471) );
  DFFRX1 \I_cache/cache_reg[6][86]  ( .D(n12093), .CK(clk), .RN(n5802), .Q(
        \I_cache/cache[6][86] ), .QN(n1842) );
  DFFRX1 \I_cache/cache_reg[7][86]  ( .D(n12092), .CK(clk), .RN(n5802), .Q(
        \I_cache/cache[7][86] ), .QN(n3498) );
  DFFRX1 \I_cache/cache_reg[0][87]  ( .D(n12091), .CK(clk), .RN(n5801), .Q(
        \I_cache/cache[0][87] ), .QN(n1780) );
  DFFRX1 \I_cache/cache_reg[1][87]  ( .D(n12090), .CK(clk), .RN(n5801), .Q(
        \I_cache/cache[1][87] ), .QN(n3436) );
  DFFRX1 \I_cache/cache_reg[2][87]  ( .D(n12089), .CK(clk), .RN(n5801), .Q(
        \I_cache/cache[2][87] ), .QN(n1811) );
  DFFRX1 \I_cache/cache_reg[3][87]  ( .D(n12088), .CK(clk), .RN(n5801), .Q(
        \I_cache/cache[3][87] ), .QN(n3467) );
  DFFRX1 \I_cache/cache_reg[4][87]  ( .D(n12087), .CK(clk), .RN(n5801), .Q(
        \I_cache/cache[4][87] ), .QN(n1810) );
  DFFRX1 \I_cache/cache_reg[5][87]  ( .D(n12086), .CK(clk), .RN(n5801), .Q(
        \I_cache/cache[5][87] ), .QN(n3466) );
  DFFRX1 \I_cache/cache_reg[6][87]  ( .D(n12085), .CK(clk), .RN(n5801), .Q(
        \I_cache/cache[6][87] ), .QN(n1839) );
  DFFRX1 \I_cache/cache_reg[7][87]  ( .D(n12084), .CK(clk), .RN(n5801), .Q(
        \I_cache/cache[7][87] ), .QN(n3495) );
  DFFRX1 \I_cache/cache_reg[0][88]  ( .D(n12083), .CK(clk), .RN(n5801), .Q(
        \I_cache/cache[0][88] ), .QN(n1779) );
  DFFRX1 \I_cache/cache_reg[1][88]  ( .D(n12082), .CK(clk), .RN(n5801), .Q(
        \I_cache/cache[1][88] ), .QN(n3435) );
  DFFRX1 \I_cache/cache_reg[2][88]  ( .D(n12081), .CK(clk), .RN(n5801), .Q(
        \I_cache/cache[2][88] ), .QN(n1805) );
  DFFRX1 \I_cache/cache_reg[3][88]  ( .D(n12080), .CK(clk), .RN(n5800), .Q(
        \I_cache/cache[3][88] ), .QN(n3461) );
  DFFRX1 \I_cache/cache_reg[4][88]  ( .D(n12079), .CK(clk), .RN(n5800), .Q(
        \I_cache/cache[4][88] ), .QN(n1804) );
  DFFRX1 \I_cache/cache_reg[5][88]  ( .D(n12078), .CK(clk), .RN(n5800), .Q(
        \I_cache/cache[5][88] ), .QN(n3460) );
  DFFRX1 \I_cache/cache_reg[6][88]  ( .D(n12077), .CK(clk), .RN(n5800), .Q(
        \I_cache/cache[6][88] ), .QN(n1836) );
  DFFRX1 \I_cache/cache_reg[7][88]  ( .D(n12076), .CK(clk), .RN(n5800), .Q(
        \I_cache/cache[7][88] ), .QN(n3492) );
  DFFRX1 \I_cache/cache_reg[0][89]  ( .D(n12075), .CK(clk), .RN(n5800), .Q(
        \I_cache/cache[0][89] ), .QN(n1777) );
  DFFRX1 \I_cache/cache_reg[1][89]  ( .D(n12074), .CK(clk), .RN(n5800), .Q(
        \I_cache/cache[1][89] ), .QN(n3433) );
  DFFRX1 \I_cache/cache_reg[2][89]  ( .D(n12073), .CK(clk), .RN(n5800), .Q(
        \I_cache/cache[2][89] ), .QN(n1799) );
  DFFRX1 \I_cache/cache_reg[3][89]  ( .D(n12072), .CK(clk), .RN(n5800), .Q(
        \I_cache/cache[3][89] ), .QN(n3455) );
  DFFRX1 \I_cache/cache_reg[4][89]  ( .D(n12071), .CK(clk), .RN(n5800), .Q(
        \I_cache/cache[4][89] ), .QN(n1798) );
  DFFRX1 \I_cache/cache_reg[5][89]  ( .D(n12070), .CK(clk), .RN(n5800), .Q(
        \I_cache/cache[5][89] ), .QN(n3454) );
  DFFRX1 \I_cache/cache_reg[6][89]  ( .D(n12069), .CK(clk), .RN(n5800), .Q(
        \I_cache/cache[6][89] ), .QN(n1833) );
  DFFRX1 \I_cache/cache_reg[7][89]  ( .D(n12068), .CK(clk), .RN(n5799), .Q(
        \I_cache/cache[7][89] ), .QN(n3489) );
  DFFRX1 \I_cache/cache_reg[0][90]  ( .D(n12067), .CK(clk), .RN(n5799), .Q(
        \I_cache/cache[0][90] ), .QN(n1562) );
  DFFRX1 \I_cache/cache_reg[1][90]  ( .D(n12066), .CK(clk), .RN(n5799), .Q(
        \I_cache/cache[1][90] ), .QN(n3145) );
  DFFRX1 \I_cache/cache_reg[2][90]  ( .D(n12065), .CK(clk), .RN(n5799), .Q(
        \I_cache/cache[2][90] ), .QN(n1561) );
  DFFRX1 \I_cache/cache_reg[3][90]  ( .D(n12064), .CK(clk), .RN(n5799), .Q(
        \I_cache/cache[3][90] ), .QN(n3144) );
  DFFRX1 \I_cache/cache_reg[4][90]  ( .D(n12063), .CK(clk), .RN(n5799), .Q(
        \I_cache/cache[4][90] ), .QN(n1572) );
  DFFRX1 \I_cache/cache_reg[5][90]  ( .D(n12062), .CK(clk), .RN(n5799), .Q(
        \I_cache/cache[5][90] ), .QN(n3154) );
  DFFRX1 \I_cache/cache_reg[6][90]  ( .D(n12061), .CK(clk), .RN(n5799), .Q(
        \I_cache/cache[6][90] ), .QN(n1563) );
  DFFRX1 \I_cache/cache_reg[7][90]  ( .D(n12060), .CK(clk), .RN(n5799), .Q(
        \I_cache/cache[7][90] ), .QN(n3146) );
  DFFRX1 \I_cache/cache_reg[0][91]  ( .D(n12059), .CK(clk), .RN(n5799), .Q(
        \I_cache/cache[0][91] ), .QN(n1539) );
  DFFRX1 \I_cache/cache_reg[1][91]  ( .D(n12058), .CK(clk), .RN(n5799), .Q(
        \I_cache/cache[1][91] ), .QN(n3121) );
  DFFRX1 \I_cache/cache_reg[2][91]  ( .D(n12057), .CK(clk), .RN(n5799), .Q(
        \I_cache/cache[2][91] ), .QN(n1538) );
  DFFRX1 \I_cache/cache_reg[3][91]  ( .D(n12056), .CK(clk), .RN(n5798), .Q(
        \I_cache/cache[3][91] ), .QN(n3120) );
  DFFRX1 \I_cache/cache_reg[4][91]  ( .D(n12055), .CK(clk), .RN(n5798), .Q(
        \I_cache/cache[4][91] ), .QN(n1607) );
  DFFRX1 \I_cache/cache_reg[5][91]  ( .D(n12054), .CK(clk), .RN(n5798), .Q(
        \I_cache/cache[5][91] ), .QN(n3184) );
  DFFRX1 \I_cache/cache_reg[6][91]  ( .D(n12053), .CK(clk), .RN(n5798), .Q(
        \I_cache/cache[6][91] ), .QN(n1540) );
  DFFRX1 \I_cache/cache_reg[0][95]  ( .D(n12027), .CK(clk), .RN(n5806), .Q(
        \I_cache/cache[0][95] ), .QN(n1551) );
  DFFRX1 \I_cache/cache_reg[2][95]  ( .D(n12025), .CK(clk), .RN(n5856), .Q(
        \I_cache/cache[2][95] ), .QN(n1550) );
  DFFRX1 \I_cache/cache_reg[0][112]  ( .D(n11891), .CK(clk), .RN(n5865), .Q(
        \I_cache/cache[0][112] ), .QN(n1905) );
  DFFRX1 \I_cache/cache_reg[1][112]  ( .D(n11890), .CK(clk), .RN(n5865), .Q(
        \I_cache/cache[1][112] ), .QN(n3560) );
  DFFRX1 \I_cache/cache_reg[2][112]  ( .D(n11889), .CK(clk), .RN(n5865), .Q(
        \I_cache/cache[2][112] ), .QN(n1906) );
  DFFRX1 \I_cache/cache_reg[3][112]  ( .D(n11888), .CK(clk), .RN(n5864), .Q(
        \I_cache/cache[3][112] ), .QN(n3561) );
  DFFRX1 \I_cache/cache_reg[4][112]  ( .D(n11887), .CK(clk), .RN(n5864), .Q(
        \I_cache/cache[4][112] ), .QN(n1868) );
  DFFRX1 \I_cache/cache_reg[5][112]  ( .D(n11886), .CK(clk), .RN(n5864), .Q(
        \I_cache/cache[5][112] ), .QN(n3524) );
  DFFRX1 \I_cache/cache_reg[6][112]  ( .D(n11885), .CK(clk), .RN(n5864), .Q(
        \I_cache/cache[6][112] ), .QN(n1930) );
  DFFRX1 \I_cache/cache_reg[7][112]  ( .D(n11884), .CK(clk), .RN(n5864), .Q(
        \I_cache/cache[7][112] ), .QN(n3584) );
  DFFRX1 \I_cache/cache_reg[0][113]  ( .D(n11883), .CK(clk), .RN(n5864), .Q(
        \I_cache/cache[0][113] ), .QN(n1896) );
  DFFRX1 \I_cache/cache_reg[1][113]  ( .D(n11882), .CK(clk), .RN(n5864), .Q(
        \I_cache/cache[1][113] ), .QN(n3551) );
  DFFRX1 \I_cache/cache_reg[2][113]  ( .D(n11881), .CK(clk), .RN(n5864), .Q(
        \I_cache/cache[2][113] ), .QN(n1897) );
  DFFRX1 \I_cache/cache_reg[3][113]  ( .D(n11880), .CK(clk), .RN(n5864), .Q(
        \I_cache/cache[3][113] ), .QN(n3552) );
  DFFRX1 \I_cache/cache_reg[4][113]  ( .D(n11879), .CK(clk), .RN(n5864), .Q(
        \I_cache/cache[4][113] ), .QN(n1828) );
  DFFRX1 \I_cache/cache_reg[5][113]  ( .D(n11878), .CK(clk), .RN(n5864), .Q(
        \I_cache/cache[5][113] ), .QN(n3484) );
  DFFRX1 \I_cache/cache_reg[6][113]  ( .D(n11877), .CK(clk), .RN(n5864), .Q(
        \I_cache/cache[6][113] ), .QN(n1926) );
  DFFRX1 \I_cache/cache_reg[7][113]  ( .D(n11876), .CK(clk), .RN(n5863), .Q(
        \I_cache/cache[7][113] ), .QN(n3580) );
  DFFRX1 \I_cache/cache_reg[0][114]  ( .D(n11875), .CK(clk), .RN(n5863), .Q(
        \I_cache/cache[0][114] ), .QN(n1892) );
  DFFRX1 \I_cache/cache_reg[1][114]  ( .D(n11874), .CK(clk), .RN(n5863), .Q(
        \I_cache/cache[1][114] ), .QN(n3547) );
  DFFRX1 \I_cache/cache_reg[2][114]  ( .D(n11873), .CK(clk), .RN(n5863), .Q(
        \I_cache/cache[2][114] ), .QN(n1860) );
  DFFRX1 \I_cache/cache_reg[3][114]  ( .D(n11872), .CK(clk), .RN(n5863), .Q(
        \I_cache/cache[3][114] ), .QN(n3516) );
  DFFRX1 \I_cache/cache_reg[4][114]  ( .D(n11871), .CK(clk), .RN(n5863), .Q(
        \I_cache/cache[4][114] ), .QN(n1859) );
  DFFRX1 \I_cache/cache_reg[5][114]  ( .D(n11870), .CK(clk), .RN(n5863), .Q(
        \I_cache/cache[5][114] ), .QN(n3515) );
  DFFRX1 \I_cache/cache_reg[6][114]  ( .D(n11869), .CK(clk), .RN(n5863), .Q(
        \I_cache/cache[6][114] ), .QN(n1922) );
  DFFRX1 \I_cache/cache_reg[7][114]  ( .D(n11868), .CK(clk), .RN(n5863), .Q(
        \I_cache/cache[7][114] ), .QN(n3576) );
  DFFRX1 \I_cache/cache_reg[0][115]  ( .D(n11867), .CK(clk), .RN(n5863), .Q(
        \I_cache/cache[0][115] ), .QN(n1888) );
  DFFRX1 \I_cache/cache_reg[1][115]  ( .D(n11866), .CK(clk), .RN(n5863), .Q(
        \I_cache/cache[1][115] ), .QN(n3543) );
  DFFRX1 \I_cache/cache_reg[2][115]  ( .D(n11865), .CK(clk), .RN(n5863), .Q(
        \I_cache/cache[2][115] ), .QN(n1889) );
  DFFRX1 \I_cache/cache_reg[3][115]  ( .D(n11864), .CK(clk), .RN(n5862), .Q(
        \I_cache/cache[3][115] ), .QN(n3544) );
  DFFRX1 \I_cache/cache_reg[4][115]  ( .D(n11863), .CK(clk), .RN(n5862), .Q(
        \I_cache/cache[4][115] ), .QN(n1863) );
  DFFRX1 \I_cache/cache_reg[5][115]  ( .D(n11862), .CK(clk), .RN(n5862), .Q(
        \I_cache/cache[5][115] ), .QN(n3519) );
  DFFRX1 \I_cache/cache_reg[6][115]  ( .D(n11861), .CK(clk), .RN(n5862), .Q(
        \I_cache/cache[6][115] ), .QN(n1920) );
  DFFRX1 \I_cache/cache_reg[7][115]  ( .D(n11860), .CK(clk), .RN(n5862), .Q(
        \I_cache/cache[7][115] ), .QN(n3574) );
  DFFRX1 \I_cache/cache_reg[0][116]  ( .D(n11859), .CK(clk), .RN(n5862), .Q(
        \I_cache/cache[0][116] ), .QN(n1876) );
  DFFRX1 \I_cache/cache_reg[1][116]  ( .D(n11858), .CK(clk), .RN(n5862), .Q(
        \I_cache/cache[1][116] ), .QN(n3531) );
  DFFRX1 \I_cache/cache_reg[2][116]  ( .D(n11857), .CK(clk), .RN(n5862), .Q(
        \I_cache/cache[2][116] ), .QN(n1878) );
  DFFRX1 \I_cache/cache_reg[3][116]  ( .D(n11856), .CK(clk), .RN(n5862), .Q(
        \I_cache/cache[3][116] ), .QN(n3533) );
  DFFRX1 \I_cache/cache_reg[4][116]  ( .D(n11855), .CK(clk), .RN(n5862), .Q(
        \I_cache/cache[4][116] ), .QN(n1877) );
  DFFRX1 \I_cache/cache_reg[5][116]  ( .D(n11854), .CK(clk), .RN(n5862), .Q(
        \I_cache/cache[5][116] ), .QN(n3532) );
  DFFRX1 \I_cache/cache_reg[6][116]  ( .D(n11853), .CK(clk), .RN(n5862), .Q(
        \I_cache/cache[6][116] ), .QN(n1916) );
  DFFRX1 \I_cache/cache_reg[7][116]  ( .D(n11852), .CK(clk), .RN(n5861), .Q(
        \I_cache/cache[7][116] ), .QN(n3570) );
  DFFRX1 \I_cache/cache_reg[0][117]  ( .D(n11851), .CK(clk), .RN(n5861), .Q(
        \I_cache/cache[0][117] ), .QN(n1792) );
  DFFRX1 \I_cache/cache_reg[1][117]  ( .D(n11850), .CK(clk), .RN(n5861), .Q(
        \I_cache/cache[1][117] ), .QN(n3448) );
  DFFRX1 \I_cache/cache_reg[2][117]  ( .D(n11849), .CK(clk), .RN(n5861), .Q(
        \I_cache/cache[2][117] ), .QN(n1820) );
  DFFRX1 \I_cache/cache_reg[3][117]  ( .D(n11848), .CK(clk), .RN(n5861), .Q(
        \I_cache/cache[3][117] ), .QN(n3476) );
  DFFRX1 \I_cache/cache_reg[4][117]  ( .D(n11847), .CK(clk), .RN(n5861), .Q(
        \I_cache/cache[4][117] ), .QN(n1819) );
  DFFRX1 \I_cache/cache_reg[5][117]  ( .D(n11846), .CK(clk), .RN(n5861), .Q(
        \I_cache/cache[5][117] ), .QN(n3475) );
  DFFRX1 \I_cache/cache_reg[6][117]  ( .D(n11845), .CK(clk), .RN(n5861), .Q(
        \I_cache/cache[6][117] ), .QN(n1844) );
  DFFRX1 \I_cache/cache_reg[7][117]  ( .D(n11844), .CK(clk), .RN(n5861), .Q(
        \I_cache/cache[7][117] ), .QN(n3500) );
  DFFRX1 \I_cache/cache_reg[0][118]  ( .D(n11843), .CK(clk), .RN(n5861), .Q(
        \I_cache/cache[0][118] ), .QN(n1791) );
  DFFRX1 \I_cache/cache_reg[1][118]  ( .D(n11842), .CK(clk), .RN(n5861), .Q(
        \I_cache/cache[1][118] ), .QN(n3447) );
  DFFRX1 \I_cache/cache_reg[3][118]  ( .D(n11840), .CK(clk), .RN(n5860), .Q(
        \I_cache/cache[3][118] ), .QN(n1875) );
  DFFRX1 \I_cache/cache_reg[4][118]  ( .D(n11839), .CK(clk), .RN(n5860), .Q(
        \I_cache/cache[4][118] ), .QN(n1814) );
  DFFRX1 \I_cache/cache_reg[5][118]  ( .D(n11838), .CK(clk), .RN(n5860), .Q(
        \I_cache/cache[5][118] ), .QN(n3470) );
  DFFRX1 \I_cache/cache_reg[6][118]  ( .D(n11837), .CK(clk), .RN(n5860), .Q(
        \I_cache/cache[6][118] ), .QN(n1841) );
  DFFRX1 \I_cache/cache_reg[7][118]  ( .D(n11836), .CK(clk), .RN(n5860), .Q(
        \I_cache/cache[7][118] ), .QN(n3497) );
  DFFRX1 \I_cache/cache_reg[0][119]  ( .D(n11835), .CK(clk), .RN(n5860), .Q(
        \I_cache/cache[0][119] ), .QN(n1789) );
  DFFRX1 \I_cache/cache_reg[1][119]  ( .D(n11834), .CK(clk), .RN(n5860), .Q(
        \I_cache/cache[1][119] ), .QN(n3445) );
  DFFRX1 \I_cache/cache_reg[2][119]  ( .D(n11833), .CK(clk), .RN(n5860), .Q(
        \I_cache/cache[2][119] ), .QN(n1807) );
  DFFRX1 \I_cache/cache_reg[3][119]  ( .D(n11832), .CK(clk), .RN(n5860), .Q(
        \I_cache/cache[3][119] ), .QN(n3463) );
  DFFRX1 \I_cache/cache_reg[4][119]  ( .D(n11831), .CK(clk), .RN(n5860), .Q(
        \I_cache/cache[4][119] ), .QN(n1806) );
  DFFRX1 \I_cache/cache_reg[5][119]  ( .D(n11830), .CK(clk), .RN(n5860), .Q(
        \I_cache/cache[5][119] ), .QN(n3462) );
  DFFRX1 \I_cache/cache_reg[6][119]  ( .D(n11829), .CK(clk), .RN(n5859), .Q(
        \I_cache/cache[6][119] ), .QN(n1837) );
  DFFRX1 \I_cache/cache_reg[7][119]  ( .D(n11828), .CK(clk), .RN(n5859), .Q(
        \I_cache/cache[7][119] ), .QN(n3493) );
  DFFRX1 \I_cache/cache_reg[0][120]  ( .D(n11827), .CK(clk), .RN(n5859), .Q(
        \I_cache/cache[0][120] ), .QN(n1788) );
  DFFRX1 \I_cache/cache_reg[1][120]  ( .D(n11826), .CK(clk), .RN(n5859), .Q(
        \I_cache/cache[1][120] ), .QN(n3444) );
  DFFRX1 \I_cache/cache_reg[2][120]  ( .D(n11825), .CK(clk), .RN(n5859), .Q(
        \I_cache/cache[2][120] ), .QN(n1803) );
  DFFRX1 \I_cache/cache_reg[3][120]  ( .D(n11824), .CK(clk), .RN(n5859), .Q(
        \I_cache/cache[3][120] ), .QN(n3459) );
  DFFRX1 \I_cache/cache_reg[4][120]  ( .D(n11823), .CK(clk), .RN(n5859), .Q(
        \I_cache/cache[4][120] ), .QN(n1802) );
  DFFRX1 \I_cache/cache_reg[5][120]  ( .D(n11822), .CK(clk), .RN(n5859), .Q(
        \I_cache/cache[5][120] ), .QN(n3458) );
  DFFRX1 \I_cache/cache_reg[6][120]  ( .D(n11821), .CK(clk), .RN(n5859), .Q(
        \I_cache/cache[6][120] ), .QN(n1835) );
  DFFRX1 \I_cache/cache_reg[7][120]  ( .D(n11820), .CK(clk), .RN(n5859), .Q(
        \I_cache/cache[7][120] ), .QN(n3491) );
  DFFRX1 \I_cache/cache_reg[0][121]  ( .D(n11819), .CK(clk), .RN(n5859), .Q(
        \I_cache/cache[0][121] ), .QN(n1786) );
  DFFRX1 \I_cache/cache_reg[1][121]  ( .D(n11818), .CK(clk), .RN(n5859), .Q(
        \I_cache/cache[1][121] ), .QN(n3442) );
  DFFRX1 \I_cache/cache_reg[2][121]  ( .D(n11817), .CK(clk), .RN(n5858), .Q(
        \I_cache/cache[2][121] ), .QN(n1795) );
  DFFRX1 \I_cache/cache_reg[3][121]  ( .D(n11816), .CK(clk), .RN(n5858), .Q(
        \I_cache/cache[3][121] ), .QN(n3451) );
  DFFRX1 \I_cache/cache_reg[4][121]  ( .D(n11815), .CK(clk), .RN(n5858), .Q(
        \I_cache/cache[4][121] ), .QN(n1794) );
  DFFRX1 \I_cache/cache_reg[5][121]  ( .D(n11814), .CK(clk), .RN(n5858), .Q(
        \I_cache/cache[5][121] ), .QN(n3450) );
  DFFRX1 \I_cache/cache_reg[6][121]  ( .D(n11813), .CK(clk), .RN(n5858), .Q(
        \I_cache/cache[6][121] ), .QN(n1831) );
  DFFRX1 \I_cache/cache_reg[7][121]  ( .D(n11812), .CK(clk), .RN(n5858), .Q(
        \I_cache/cache[7][121] ), .QN(n3487) );
  DFFRX1 \I_cache/cache_reg[0][122]  ( .D(n11811), .CK(clk), .RN(n5858), .Q(
        \I_cache/cache[0][122] ), .QN(n1557) );
  DFFRX1 \I_cache/cache_reg[1][122]  ( .D(n11810), .CK(clk), .RN(n5858), .Q(
        \I_cache/cache[1][122] ), .QN(n3139) );
  DFFRX1 \I_cache/cache_reg[2][122]  ( .D(n11809), .CK(clk), .RN(n5858), .Q(
        \I_cache/cache[2][122] ), .QN(n1556) );
  DFFRX1 \I_cache/cache_reg[3][122]  ( .D(n11808), .CK(clk), .RN(n5858), .Q(
        \I_cache/cache[3][122] ), .QN(n3138) );
  DFFRX1 \I_cache/cache_reg[4][122]  ( .D(n11807), .CK(clk), .RN(n5858), .Q(
        \I_cache/cache[4][122] ), .QN(n1570) );
  DFFRX1 \I_cache/cache_reg[5][122]  ( .D(n11806), .CK(clk), .RN(n5858), .Q(
        \I_cache/cache[5][122] ), .QN(n3152) );
  DFFRX1 \I_cache/cache_reg[6][122]  ( .D(n11805), .CK(clk), .RN(n5857), .Q(
        \I_cache/cache[6][122] ), .QN(n1558) );
  DFFRX1 \I_cache/cache_reg[7][122]  ( .D(n11804), .CK(clk), .RN(n5857), .Q(
        \I_cache/cache[7][122] ), .QN(n3140) );
  DFFRX1 \I_cache/cache_reg[0][123]  ( .D(n11803), .CK(clk), .RN(n5857), .Q(
        \I_cache/cache[0][123] ), .QN(n1533) );
  DFFRX1 \I_cache/cache_reg[1][123]  ( .D(n11802), .CK(clk), .RN(n5857), .Q(
        \I_cache/cache[1][123] ), .QN(n3115) );
  DFFRX1 \I_cache/cache_reg[2][123]  ( .D(n11801), .CK(clk), .RN(n5857), .Q(
        \I_cache/cache[2][123] ), .QN(n1532) );
  DFFRX1 \I_cache/cache_reg[3][123]  ( .D(n11800), .CK(clk), .RN(n5857), .Q(
        \I_cache/cache[3][123] ), .QN(n3114) );
  DFFRX1 \I_cache/cache_reg[4][123]  ( .D(n11799), .CK(clk), .RN(n5857), .Q(
        \I_cache/cache[4][123] ), .QN(n1606) );
  DFFRX1 \I_cache/cache_reg[5][123]  ( .D(n11798), .CK(clk), .RN(n5857), .Q(
        \I_cache/cache[5][123] ), .QN(n3183) );
  DFFRX1 \I_cache/cache_reg[6][123]  ( .D(n11797), .CK(clk), .RN(n5857), .Q(
        \I_cache/cache[6][123] ), .QN(n1534) );
  DFFRX1 \I_cache/cache_reg[7][123]  ( .D(n11796), .CK(clk), .RN(n5857), .Q(
        \I_cache/cache[7][123] ), .QN(n3116) );
  DFFRX1 \I_cache/cache_reg[0][127]  ( .D(n11771), .CK(clk), .RN(n5835), .Q(
        \I_cache/cache[0][127] ), .QN(n1545) );
  DFFRX1 \I_cache/cache_reg[2][127]  ( .D(n11769), .CK(clk), .RN(n5835), .Q(
        \I_cache/cache[2][127] ), .QN(n1544) );
  DFFRX1 \I_cache/cache_reg[4][127]  ( .D(n11767), .CK(clk), .RN(n5834), .Q(
        \I_cache/cache[4][127] ), .QN(n1602) );
  DFFRX1 \i_MIPS/Register/register_reg[30][19]  ( .D(\i_MIPS/Register/n167 ), 
        .CK(clk), .RN(n5725), .Q(\i_MIPS/Register/register[30][19] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][30]  ( .D(\i_MIPS/Register/n178 ), 
        .CK(clk), .RN(n5724), .Q(\i_MIPS/Register/register[30][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[28][19]  ( .D(\i_MIPS/Register/n231 ), 
        .CK(clk), .RN(n5719), .Q(\i_MIPS/Register/register[28][19] ) );
  DFFRX1 \i_MIPS/Register/register_reg[28][30]  ( .D(\i_MIPS/Register/n242 ), 
        .CK(clk), .RN(n5718), .Q(\i_MIPS/Register/register[28][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[24][19]  ( .D(\i_MIPS/Register/n359 ), 
        .CK(clk), .RN(n5769), .Q(\i_MIPS/Register/register[24][19] ) );
  DFFRX1 \i_MIPS/Register/register_reg[24][30]  ( .D(\i_MIPS/Register/n370 ), 
        .CK(clk), .RN(n5768), .Q(\i_MIPS/Register/register[24][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][19]  ( .D(\i_MIPS/Register/n679 ), 
        .CK(clk), .RN(n5762), .Q(\i_MIPS/Register/register[14][19] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][30]  ( .D(\i_MIPS/Register/n690 ), 
        .CK(clk), .RN(n5761), .Q(\i_MIPS/Register/register[14][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[12][19]  ( .D(\i_MIPS/Register/n743 ), 
        .CK(clk), .RN(n5756), .Q(\i_MIPS/Register/register[12][19] ) );
  DFFRX1 \i_MIPS/Register/register_reg[12][30]  ( .D(\i_MIPS/Register/n754 ), 
        .CK(clk), .RN(n5656), .Q(\i_MIPS/Register/register[12][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[8][19]  ( .D(\i_MIPS/Register/n871 ), 
        .CK(clk), .RN(n5666), .Q(\i_MIPS/Register/register[8][19] ) );
  DFFRX1 \i_MIPS/Register/register_reg[8][30]  ( .D(\i_MIPS/Register/n882 ), 
        .CK(clk), .RN(n5665), .Q(\i_MIPS/Register/register[8][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][19]  ( .D(\i_MIPS/Register/n423 ), 
        .CK(clk), .RN(n5783), .Q(\i_MIPS/Register/register[22][19] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][22]  ( .D(\i_MIPS/Register/n426 ), 
        .CK(clk), .RN(n5783), .Q(\i_MIPS/Register/register[22][22] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][30]  ( .D(\i_MIPS/Register/n434 ), 
        .CK(clk), .RN(n5782), .Q(\i_MIPS/Register/register[22][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[20][19]  ( .D(\i_MIPS/Register/n487 ), 
        .CK(clk), .RN(n5778), .Q(\i_MIPS/Register/register[20][19] ) );
  DFFRX1 \i_MIPS/Register/register_reg[20][30]  ( .D(\i_MIPS/Register/n498 ), 
        .CK(clk), .RN(n5777), .Q(\i_MIPS/Register/register[20][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[16][19]  ( .D(\i_MIPS/Register/n615 ), 
        .CK(clk), .RN(n5747), .Q(\i_MIPS/Register/register[16][19] ) );
  DFFRX1 \i_MIPS/Register/register_reg[16][30]  ( .D(\i_MIPS/Register/n626 ), 
        .CK(clk), .RN(n5746), .Q(\i_MIPS/Register/register[16][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][12]  ( .D(\i_MIPS/Register/n928 ), 
        .CK(clk), .RN(n5661), .Q(\i_MIPS/Register/register[6][12] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][17]  ( .D(\i_MIPS/Register/n933 ), 
        .CK(clk), .RN(n5661), .Q(\i_MIPS/Register/register[6][17] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][19]  ( .D(\i_MIPS/Register/n935 ), 
        .CK(clk), .RN(n5661), .Q(\i_MIPS/Register/register[6][19] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][22]  ( .D(\i_MIPS/Register/n938 ), 
        .CK(clk), .RN(n5661), .Q(\i_MIPS/Register/register[6][22] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][29]  ( .D(\i_MIPS/Register/n945 ), 
        .CK(clk), .RN(n5660), .Q(\i_MIPS/Register/register[6][29] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][30]  ( .D(\i_MIPS/Register/n946 ), 
        .CK(clk), .RN(n5660), .Q(\i_MIPS/Register/register[6][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[4][19]  ( .D(\i_MIPS/Register/n999 ), 
        .CK(clk), .RN(n5636), .Q(\i_MIPS/Register/register[4][19] ) );
  DFFRX1 \i_MIPS/Register/register_reg[4][30]  ( .D(\i_MIPS/Register/n1010 ), 
        .CK(clk), .RN(n5635), .Q(\i_MIPS/Register/register[4][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[0][19]  ( .D(\i_MIPS/Register/n1127 ), 
        .CK(clk), .RN(n5645), .Q(\i_MIPS/Register/register[0][19] ) );
  DFFRX1 \i_MIPS/Register/register_reg[0][30]  ( .D(\i_MIPS/Register/n1138 ), 
        .CK(clk), .RN(n5644), .Q(\i_MIPS/Register/register[0][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[28][5]  ( .D(\i_MIPS/Register/n217 ), 
        .CK(clk), .RN(n5721), .Q(\i_MIPS/Register/register[28][5] ), .QN(n1017) );
  DFFRX1 \i_MIPS/Register/register_reg[28][8]  ( .D(\i_MIPS/Register/n220 ), 
        .CK(clk), .RN(n5720), .Q(\i_MIPS/Register/register[28][8] ), .QN(n961)
         );
  DFFRX1 \i_MIPS/Register/register_reg[28][11]  ( .D(\i_MIPS/Register/n223 ), 
        .CK(clk), .RN(n5720), .Q(\i_MIPS/Register/register[28][11] ), .QN(n398) );
  DFFRX1 \i_MIPS/Register/register_reg[28][12]  ( .D(\i_MIPS/Register/n224 ), 
        .CK(clk), .RN(n5720), .Q(\i_MIPS/Register/register[28][12] ), .QN(n399) );
  DFFRX1 \i_MIPS/Register/register_reg[28][17]  ( .D(\i_MIPS/Register/n229 ), 
        .CK(clk), .RN(n5720), .Q(\i_MIPS/Register/register[28][17] ), .QN(
        n1018) );
  DFFRX1 \i_MIPS/Register/register_reg[28][22]  ( .D(\i_MIPS/Register/n234 ), 
        .CK(clk), .RN(n5719), .Q(\i_MIPS/Register/register[28][22] ), .QN(n957) );
  DFFRX1 \i_MIPS/Register/register_reg[28][24]  ( .D(\i_MIPS/Register/n236 ), 
        .CK(clk), .RN(n5719), .Q(\i_MIPS/Register/register[28][24] ), .QN(
        n1016) );
  DFFRX1 \i_MIPS/Register/register_reg[28][29]  ( .D(\i_MIPS/Register/n241 ), 
        .CK(clk), .RN(n5719), .Q(\i_MIPS/Register/register[28][29] ), .QN(n888) );
  DFFRX1 \i_MIPS/Register/register_reg[24][5]  ( .D(\i_MIPS/Register/n345 ), 
        .CK(clk), .RN(n5770), .Q(\i_MIPS/Register/register[24][5] ), .QN(n466)
         );
  DFFRX1 \i_MIPS/Register/register_reg[24][12]  ( .D(\i_MIPS/Register/n352 ), 
        .CK(clk), .RN(n5769), .Q(\i_MIPS/Register/register[24][12] ), .QN(n992) );
  DFFRX1 \i_MIPS/Register/register_reg[24][17]  ( .D(\i_MIPS/Register/n357 ), 
        .CK(clk), .RN(n5769), .Q(\i_MIPS/Register/register[24][17] ), .QN(n359) );
  DFFRX1 \i_MIPS/Register/register_reg[24][22]  ( .D(\i_MIPS/Register/n362 ), 
        .CK(clk), .RN(n5768), .Q(\i_MIPS/Register/register[24][22] ), .QN(n945) );
  DFFRX1 \i_MIPS/Register/register_reg[24][29]  ( .D(\i_MIPS/Register/n369 ), 
        .CK(clk), .RN(n5768), .Q(\i_MIPS/Register/register[24][29] ), .QN(n400) );
  DFFRX1 \i_MIPS/Register/register_reg[12][5]  ( .D(\i_MIPS/Register/n729 ), 
        .CK(clk), .RN(n5758), .Q(\i_MIPS/Register/register[12][5] ), .QN(n968)
         );
  DFFRX1 \i_MIPS/Register/register_reg[12][8]  ( .D(\i_MIPS/Register/n732 ), 
        .CK(clk), .RN(n5757), .Q(\i_MIPS/Register/register[12][8] ), .QN(n1021) );
  DFFRX1 \i_MIPS/Register/register_reg[12][11]  ( .D(\i_MIPS/Register/n735 ), 
        .CK(clk), .RN(n5757), .Q(\i_MIPS/Register/register[12][11] ), .QN(n336) );
  DFFRX1 \i_MIPS/Register/register_reg[12][12]  ( .D(\i_MIPS/Register/n736 ), 
        .CK(clk), .RN(n5757), .Q(\i_MIPS/Register/register[12][12] ), .QN(n380) );
  DFFRX1 \i_MIPS/Register/register_reg[12][17]  ( .D(\i_MIPS/Register/n741 ), 
        .CK(clk), .RN(n5757), .Q(\i_MIPS/Register/register[12][17] ), .QN(n859) );
  DFFRX1 \i_MIPS/Register/register_reg[12][22]  ( .D(\i_MIPS/Register/n746 ), 
        .CK(clk), .RN(n5761), .Q(\i_MIPS/Register/register[12][22] ), .QN(
        n1019) );
  DFFRX1 \i_MIPS/Register/register_reg[12][24]  ( .D(\i_MIPS/Register/n748 ), 
        .CK(clk), .RN(n5666), .Q(\i_MIPS/Register/register[12][24] ), .QN(n977) );
  DFFRX1 \i_MIPS/Register/register_reg[12][29]  ( .D(\i_MIPS/Register/n753 ), 
        .CK(clk), .RN(n5656), .Q(\i_MIPS/Register/register[12][29] ), .QN(n866) );
  DFFRX1 \i_MIPS/Register/register_reg[8][5]  ( .D(\i_MIPS/Register/n857 ), 
        .CK(clk), .RN(n5647), .Q(\i_MIPS/Register/register[8][5] ), .QN(n445)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][11]  ( .D(\i_MIPS/Register/n863 ), 
        .CK(clk), .RN(n5647), .Q(\i_MIPS/Register/register[8][11] ), .QN(n895)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][12]  ( .D(\i_MIPS/Register/n864 ), 
        .CK(clk), .RN(n5647), .Q(\i_MIPS/Register/register[8][12] ), .QN(n944)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][17]  ( .D(\i_MIPS/Register/n869 ), 
        .CK(clk), .RN(n5666), .Q(\i_MIPS/Register/register[8][17] ), .QN(n328)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][22]  ( .D(\i_MIPS/Register/n874 ), 
        .CK(clk), .RN(n5666), .Q(\i_MIPS/Register/register[8][22] ), .QN(n993)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][29]  ( .D(\i_MIPS/Register/n881 ), 
        .CK(clk), .RN(n5665), .Q(\i_MIPS/Register/register[8][29] ), .QN(n379)
         );
  DFFRX1 \i_MIPS/Register/register_reg[20][22]  ( .D(\i_MIPS/Register/n490 ), 
        .CK(clk), .RN(n5778), .Q(\i_MIPS/Register/register[20][22] ), .QN(
        n2473) );
  DFFRX1 \i_MIPS/Register/register_reg[16][22]  ( .D(\i_MIPS/Register/n618 ), 
        .CK(clk), .RN(n5747), .Q(\i_MIPS/Register/register[16][22] ), .QN(
        n2457) );
  DFFRX1 \i_MIPS/Register/register_reg[4][22]  ( .D(\i_MIPS/Register/n1002 ), 
        .CK(clk), .RN(n5635), .Q(\i_MIPS/Register/register[4][22] ), .QN(n2545) );
  DFFRX1 \i_MIPS/Register/register_reg[0][22]  ( .D(\i_MIPS/Register/n1130 ), 
        .CK(clk), .RN(n5644), .Q(\i_MIPS/Register/register[0][22] ), .QN(n2517) );
  DFFRX1 \i_MIPS/Register/register_reg[18][0]  ( .D(\i_MIPS/Register/n532 ), 
        .CK(clk), .RN(n5754), .Q(\i_MIPS/Register/register[18][0] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][2]  ( .D(\i_MIPS/Register/n534 ), 
        .CK(clk), .RN(n5754), .Q(\i_MIPS/Register/register[18][2] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][3]  ( .D(\i_MIPS/Register/n535 ), 
        .CK(clk), .RN(n5754), .Q(\i_MIPS/Register/register[18][3] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][4]  ( .D(\i_MIPS/Register/n536 ), 
        .CK(clk), .RN(n5754), .Q(\i_MIPS/Register/register[18][4] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][5]  ( .D(\i_MIPS/Register/n537 ), 
        .CK(clk), .RN(n5754), .Q(\i_MIPS/Register/register[18][5] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][6]  ( .D(\i_MIPS/Register/n538 ), 
        .CK(clk), .RN(n5754), .Q(\i_MIPS/Register/register[18][6] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][7]  ( .D(\i_MIPS/Register/n539 ), 
        .CK(clk), .RN(n5754), .Q(\i_MIPS/Register/register[18][7] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][8]  ( .D(\i_MIPS/Register/n540 ), 
        .CK(clk), .RN(n5754), .Q(\i_MIPS/Register/register[18][8] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][9]  ( .D(\i_MIPS/Register/n541 ), 
        .CK(clk), .RN(n5754), .Q(\i_MIPS/Register/register[18][9] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][11]  ( .D(\i_MIPS/Register/n543 ), 
        .CK(clk), .RN(n5753), .Q(\i_MIPS/Register/register[18][11] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][12]  ( .D(\i_MIPS/Register/n544 ), 
        .CK(clk), .RN(n5753), .Q(\i_MIPS/Register/register[18][12] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][14]  ( .D(\i_MIPS/Register/n546 ), 
        .CK(clk), .RN(n5753), .Q(\i_MIPS/Register/register[18][14] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][15]  ( .D(\i_MIPS/Register/n547 ), 
        .CK(clk), .RN(n5753), .Q(\i_MIPS/Register/register[18][15] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][16]  ( .D(\i_MIPS/Register/n548 ), 
        .CK(clk), .RN(n5753), .Q(\i_MIPS/Register/register[18][16] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][17]  ( .D(\i_MIPS/Register/n549 ), 
        .CK(clk), .RN(n5753), .Q(\i_MIPS/Register/register[18][17] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][19]  ( .D(\i_MIPS/Register/n551 ), 
        .CK(clk), .RN(n5753), .Q(\i_MIPS/Register/register[18][19] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][20]  ( .D(\i_MIPS/Register/n552 ), 
        .CK(clk), .RN(n5753), .Q(\i_MIPS/Register/register[18][20] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][21]  ( .D(\i_MIPS/Register/n553 ), 
        .CK(clk), .RN(n5753), .Q(\i_MIPS/Register/register[18][21] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][22]  ( .D(\i_MIPS/Register/n554 ), 
        .CK(clk), .RN(n5752), .Q(\i_MIPS/Register/register[18][22] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][23]  ( .D(\i_MIPS/Register/n555 ), 
        .CK(clk), .RN(n5752), .Q(\i_MIPS/Register/register[18][23] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][25]  ( .D(\i_MIPS/Register/n557 ), 
        .CK(clk), .RN(n5752), .Q(\i_MIPS/Register/register[18][25] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][26]  ( .D(\i_MIPS/Register/n558 ), 
        .CK(clk), .RN(n5752), .Q(\i_MIPS/Register/register[18][26] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][27]  ( .D(\i_MIPS/Register/n559 ), 
        .CK(clk), .RN(n5752), .Q(\i_MIPS/Register/register[18][27] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][28]  ( .D(\i_MIPS/Register/n560 ), 
        .CK(clk), .RN(n5752), .Q(\i_MIPS/Register/register[18][28] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][29]  ( .D(\i_MIPS/Register/n561 ), 
        .CK(clk), .RN(n5752), .Q(\i_MIPS/Register/register[18][29] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][30]  ( .D(\i_MIPS/Register/n562 ), 
        .CK(clk), .RN(n5752), .Q(\i_MIPS/Register/register[18][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][0]  ( .D(\i_MIPS/Register/n1044 ), 
        .CK(clk), .RN(n5632), .Q(\i_MIPS/Register/register[2][0] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][2]  ( .D(\i_MIPS/Register/n1046 ), 
        .CK(clk), .RN(n5632), .Q(\i_MIPS/Register/register[2][2] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][3]  ( .D(\i_MIPS/Register/n1047 ), 
        .CK(clk), .RN(n5632), .Q(\i_MIPS/Register/register[2][3] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][4]  ( .D(\i_MIPS/Register/n1048 ), 
        .CK(clk), .RN(n5631), .Q(\i_MIPS/Register/register[2][4] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][5]  ( .D(\i_MIPS/Register/n1049 ), 
        .CK(clk), .RN(n5631), .Q(\i_MIPS/Register/register[2][5] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][6]  ( .D(\i_MIPS/Register/n1050 ), 
        .CK(clk), .RN(n5631), .Q(\i_MIPS/Register/register[2][6] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][7]  ( .D(\i_MIPS/Register/n1051 ), 
        .CK(clk), .RN(n5631), .Q(\i_MIPS/Register/register[2][7] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][8]  ( .D(\i_MIPS/Register/n1052 ), 
        .CK(clk), .RN(n5631), .Q(\i_MIPS/Register/register[2][8] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][9]  ( .D(\i_MIPS/Register/n1053 ), 
        .CK(clk), .RN(n5631), .Q(\i_MIPS/Register/register[2][9] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][11]  ( .D(\i_MIPS/Register/n1055 ), 
        .CK(clk), .RN(n5631), .Q(\i_MIPS/Register/register[2][11] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][12]  ( .D(\i_MIPS/Register/n1056 ), 
        .CK(clk), .RN(n5631), .Q(\i_MIPS/Register/register[2][12] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][14]  ( .D(\i_MIPS/Register/n1058 ), 
        .CK(clk), .RN(n5631), .Q(\i_MIPS/Register/register[2][14] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][15]  ( .D(\i_MIPS/Register/n1059 ), 
        .CK(clk), .RN(n5630), .Q(\i_MIPS/Register/register[2][15] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][16]  ( .D(\i_MIPS/Register/n1060 ), 
        .CK(clk), .RN(n5630), .Q(\i_MIPS/Register/register[2][16] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][17]  ( .D(\i_MIPS/Register/n1061 ), 
        .CK(clk), .RN(n5630), .Q(\i_MIPS/Register/register[2][17] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][19]  ( .D(\i_MIPS/Register/n1063 ), 
        .CK(clk), .RN(n5630), .Q(\i_MIPS/Register/register[2][19] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][20]  ( .D(\i_MIPS/Register/n1064 ), 
        .CK(clk), .RN(n5630), .Q(\i_MIPS/Register/register[2][20] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][21]  ( .D(\i_MIPS/Register/n1065 ), 
        .CK(clk), .RN(n5630), .Q(\i_MIPS/Register/register[2][21] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][22]  ( .D(\i_MIPS/Register/n1066 ), 
        .CK(clk), .RN(n5630), .Q(\i_MIPS/Register/register[2][22] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][23]  ( .D(\i_MIPS/Register/n1067 ), 
        .CK(clk), .RN(n5630), .Q(\i_MIPS/Register/register[2][23] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][25]  ( .D(\i_MIPS/Register/n1069 ), 
        .CK(clk), .RN(n5630), .Q(\i_MIPS/Register/register[2][25] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][26]  ( .D(\i_MIPS/Register/n1070 ), 
        .CK(clk), .RN(n5630), .Q(\i_MIPS/Register/register[2][26] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][27]  ( .D(\i_MIPS/Register/n1071 ), 
        .CK(clk), .RN(n5629), .Q(\i_MIPS/Register/register[2][27] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][28]  ( .D(\i_MIPS/Register/n1072 ), 
        .CK(clk), .RN(n5629), .Q(\i_MIPS/Register/register[2][28] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][29]  ( .D(\i_MIPS/Register/n1073 ), 
        .CK(clk), .RN(n5629), .Q(\i_MIPS/Register/register[2][29] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][30]  ( .D(\i_MIPS/Register/n1074 ), 
        .CK(clk), .RN(n5629), .Q(\i_MIPS/Register/register[2][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][3]  ( .D(\i_MIPS/Register/n279 ), 
        .CK(clk), .RN(n5775), .Q(\i_MIPS/Register/register[26][3] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][4]  ( .D(\i_MIPS/Register/n280 ), 
        .CK(clk), .RN(n5775), .Q(\i_MIPS/Register/register[26][4] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][5]  ( .D(\i_MIPS/Register/n281 ), 
        .CK(clk), .RN(n5775), .Q(\i_MIPS/Register/register[26][5] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][8]  ( .D(\i_MIPS/Register/n284 ), 
        .CK(clk), .RN(n5775), .Q(\i_MIPS/Register/register[26][8] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][11]  ( .D(\i_MIPS/Register/n287 ), 
        .CK(clk), .RN(n5775), .Q(\i_MIPS/Register/register[26][11] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][12]  ( .D(\i_MIPS/Register/n288 ), 
        .CK(clk), .RN(n5775), .Q(\i_MIPS/Register/register[26][12] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][15]  ( .D(\i_MIPS/Register/n291 ), 
        .CK(clk), .RN(n5774), .Q(\i_MIPS/Register/register[26][15] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][17]  ( .D(\i_MIPS/Register/n293 ), 
        .CK(clk), .RN(n5774), .Q(\i_MIPS/Register/register[26][17] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][19]  ( .D(\i_MIPS/Register/n295 ), 
        .CK(clk), .RN(n5774), .Q(\i_MIPS/Register/register[26][19] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][22]  ( .D(\i_MIPS/Register/n298 ), 
        .CK(clk), .RN(n5774), .Q(\i_MIPS/Register/register[26][22] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][25]  ( .D(\i_MIPS/Register/n301 ), 
        .CK(clk), .RN(n5774), .Q(\i_MIPS/Register/register[26][25] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][26]  ( .D(\i_MIPS/Register/n302 ), 
        .CK(clk), .RN(n5774), .Q(\i_MIPS/Register/register[26][26] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][27]  ( .D(\i_MIPS/Register/n303 ), 
        .CK(clk), .RN(n5773), .Q(\i_MIPS/Register/register[26][27] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][29]  ( .D(\i_MIPS/Register/n305 ), 
        .CK(clk), .RN(n5773), .Q(\i_MIPS/Register/register[26][29] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][30]  ( .D(\i_MIPS/Register/n306 ), 
        .CK(clk), .RN(n5773), .Q(\i_MIPS/Register/register[26][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][0]  ( .D(\i_MIPS/Register/n788 ), 
        .CK(clk), .RN(n5653), .Q(\i_MIPS/Register/register[10][0] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][3]  ( .D(\i_MIPS/Register/n791 ), 
        .CK(clk), .RN(n5653), .Q(\i_MIPS/Register/register[10][3] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][4]  ( .D(\i_MIPS/Register/n792 ), 
        .CK(clk), .RN(n5653), .Q(\i_MIPS/Register/register[10][4] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][5]  ( .D(\i_MIPS/Register/n793 ), 
        .CK(clk), .RN(n5653), .Q(\i_MIPS/Register/register[10][5] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][7]  ( .D(\i_MIPS/Register/n795 ), 
        .CK(clk), .RN(n5653), .Q(\i_MIPS/Register/register[10][7] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][8]  ( .D(\i_MIPS/Register/n796 ), 
        .CK(clk), .RN(n5653), .Q(\i_MIPS/Register/register[10][8] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][11]  ( .D(\i_MIPS/Register/n799 ), 
        .CK(clk), .RN(n5652), .Q(\i_MIPS/Register/register[10][11] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][12]  ( .D(\i_MIPS/Register/n800 ), 
        .CK(clk), .RN(n5652), .Q(\i_MIPS/Register/register[10][12] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][15]  ( .D(\i_MIPS/Register/n803 ), 
        .CK(clk), .RN(n5652), .Q(\i_MIPS/Register/register[10][15] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][17]  ( .D(\i_MIPS/Register/n805 ), 
        .CK(clk), .RN(n5652), .Q(\i_MIPS/Register/register[10][17] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][19]  ( .D(\i_MIPS/Register/n807 ), 
        .CK(clk), .RN(n5652), .Q(\i_MIPS/Register/register[10][19] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][22]  ( .D(\i_MIPS/Register/n810 ), 
        .CK(clk), .RN(n5651), .Q(\i_MIPS/Register/register[10][22] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][25]  ( .D(\i_MIPS/Register/n813 ), 
        .CK(clk), .RN(n5651), .Q(\i_MIPS/Register/register[10][25] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][26]  ( .D(\i_MIPS/Register/n814 ), 
        .CK(clk), .RN(n5651), .Q(\i_MIPS/Register/register[10][26] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][27]  ( .D(\i_MIPS/Register/n815 ), 
        .CK(clk), .RN(n5651), .Q(\i_MIPS/Register/register[10][27] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][29]  ( .D(\i_MIPS/Register/n817 ), 
        .CK(clk), .RN(n5651), .Q(\i_MIPS/Register/register[10][29] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][30]  ( .D(\i_MIPS/Register/n818 ), 
        .CK(clk), .RN(n5651), .Q(\i_MIPS/Register/register[10][30] ) );
  DFFRX1 \i_MIPS/IF_ID_reg[62]  ( .D(\i_MIPS/N88 ), .CK(clk), .RN(n5716), .Q(
        \i_MIPS/IR_ID[30] ), .QN(\i_MIPS/n330 ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][31]  ( .D(\i_MIPS/Register/n179 ), 
        .CK(clk), .RN(n5724), .Q(\i_MIPS/Register/register[30][31] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][31]  ( .D(\i_MIPS/Register/n691 ), 
        .CK(clk), .RN(n5761), .Q(\i_MIPS/Register/register[14][31] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][31]  ( .D(\i_MIPS/Register/n435 ), 
        .CK(clk), .RN(n5782), .Q(\i_MIPS/Register/register[22][31] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][31]  ( .D(\i_MIPS/Register/n947 ), 
        .CK(clk), .RN(n5660), .Q(\i_MIPS/Register/register[6][31] ) );
  DFFRX1 \i_MIPS/Register/register_reg[23][31]  ( .D(\i_MIPS/Register/n403 ), 
        .CK(clk), .RN(n5785), .Q(\i_MIPS/Register/register[23][31] ) );
  DFFRX1 \i_MIPS/Register/register_reg[21][31]  ( .D(\i_MIPS/Register/n467 ), 
        .CK(clk), .RN(n5780), .Q(\i_MIPS/Register/register[21][31] ) );
  DFFRX1 \i_MIPS/Register/register_reg[19][31]  ( .D(\i_MIPS/Register/n531 ), 
        .CK(clk), .RN(n5754), .Q(\i_MIPS/Register/register[19][31] ) );
  DFFRX1 \i_MIPS/Register/register_reg[17][31]  ( .D(\i_MIPS/Register/n595 ), 
        .CK(clk), .RN(n5749), .Q(\i_MIPS/Register/register[17][31] ) );
  DFFRX1 \i_MIPS/Register/register_reg[7][31]  ( .D(\i_MIPS/Register/n915 ), 
        .CK(clk), .RN(n5663), .Q(\i_MIPS/Register/register[7][31] ) );
  DFFRX1 \i_MIPS/Register/register_reg[5][31]  ( .D(\i_MIPS/Register/n979 ), 
        .CK(clk), .RN(n5657), .Q(\i_MIPS/Register/register[5][31] ) );
  DFFRX1 \i_MIPS/Register/register_reg[3][31]  ( .D(\i_MIPS/Register/n1043 ), 
        .CK(clk), .RN(n5632), .Q(\i_MIPS/Register/register[3][31] ) );
  DFFRX1 \i_MIPS/Register/register_reg[1][31]  ( .D(\i_MIPS/Register/n1107 ), 
        .CK(clk), .RN(n5646), .Q(\i_MIPS/Register/register[1][31] ) );
  DFFRX1 \i_MIPS/Register/register_reg[29][31]  ( .D(\i_MIPS/Register/n211 ), 
        .CK(clk), .RN(n5721), .Q(\i_MIPS/Register/register[29][31] ) );
  DFFRX1 \i_MIPS/Register/register_reg[27][31]  ( .D(\i_MIPS/Register/n275 ), 
        .CK(clk), .RN(n5776), .Q(\i_MIPS/Register/register[27][31] ) );
  DFFRX1 \i_MIPS/Register/register_reg[25][31]  ( .D(\i_MIPS/Register/n339 ), 
        .CK(clk), .RN(n5770), .Q(\i_MIPS/Register/register[25][31] ) );
  DFFRX1 \i_MIPS/Register/register_reg[15][31]  ( .D(\i_MIPS/Register/n659 ), 
        .CK(clk), .RN(n5764), .Q(\i_MIPS/Register/register[15][31] ) );
  DFFRX1 \i_MIPS/Register/register_reg[13][31]  ( .D(\i_MIPS/Register/n723 ), 
        .CK(clk), .RN(n5758), .Q(\i_MIPS/Register/register[13][31] ) );
  DFFRX1 \i_MIPS/Register/register_reg[11][31]  ( .D(\i_MIPS/Register/n787 ), 
        .CK(clk), .RN(n5653), .Q(\i_MIPS/Register/register[11][31] ) );
  DFFRX1 \i_MIPS/Register/register_reg[9][31]  ( .D(\i_MIPS/Register/n851 ), 
        .CK(clk), .RN(n5648), .Q(\i_MIPS/Register/register[9][31] ) );
  DFFRX1 \i_MIPS/Register/register_reg[28][31]  ( .D(\i_MIPS/Register/n243 ), 
        .CK(clk), .RN(n5718), .Q(\i_MIPS/Register/register[28][31] ), .QN(n434) );
  DFFRX1 \i_MIPS/Register/register_reg[12][31]  ( .D(\i_MIPS/Register/n755 ), 
        .CK(clk), .RN(n5656), .Q(\i_MIPS/Register/register[12][31] ), .QN(n435) );
  DFFRX1 \i_MIPS/Register/register_reg[20][31]  ( .D(\i_MIPS/Register/n499 ), 
        .CK(clk), .RN(n5777), .Q(\i_MIPS/Register/register[20][31] ), .QN(
        n2014) );
  DFFRX1 \i_MIPS/Register/register_reg[4][31]  ( .D(\i_MIPS/Register/n1011 ), 
        .CK(clk), .RN(n5635), .Q(\i_MIPS/Register/register[4][31] ), .QN(n2015) );
  DFFRX1 \i_MIPS/Register/register_reg[31][31]  ( .D(n11514), .CK(clk), .RN(
        n5707), .Q(\i_MIPS/Register/register[31][31] ), .QN(n1937) );
  DFFRX1 \i_MIPS/Register/register_reg[26][31]  ( .D(\i_MIPS/Register/n307 ), 
        .CK(clk), .RN(n5773), .Q(\i_MIPS/Register/register[26][31] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][31]  ( .D(\i_MIPS/Register/n819 ), 
        .CK(clk), .RN(n5651), .Q(\i_MIPS/Register/register[10][31] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][31]  ( .D(\i_MIPS/Register/n563 ), 
        .CK(clk), .RN(n5752), .Q(\i_MIPS/Register/register[18][31] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][31]  ( .D(\i_MIPS/Register/n1075 ), 
        .CK(clk), .RN(n5629), .Q(\i_MIPS/Register/register[2][31] ) );
  DFFRX1 \i_MIPS/Register/register_reg[24][31]  ( .D(\i_MIPS/Register/n371 ), 
        .CK(clk), .RN(n5768), .Q(\i_MIPS/Register/register[24][31] ), .QN(n936) );
  DFFRX1 \i_MIPS/Register/register_reg[16][31]  ( .D(\i_MIPS/Register/n627 ), 
        .CK(clk), .RN(n5751), .Q(\i_MIPS/Register/register[16][31] ), .QN(
        n2645) );
  DFFRX1 \i_MIPS/Register/register_reg[8][31]  ( .D(\i_MIPS/Register/n883 ), 
        .CK(clk), .RN(n5665), .Q(\i_MIPS/Register/register[8][31] ), .QN(n433)
         );
  DFFRX1 \i_MIPS/Register/register_reg[0][31]  ( .D(\i_MIPS/Register/n1139 ), 
        .CK(clk), .RN(n5644), .Q(\i_MIPS/Register/register[0][31] ), .QN(n2644) );
  DFFRX1 \i_MIPS/PHT_2/history_state_reg[0]  ( .D(\i_MIPS/PHT_2/n52 ), .CK(clk), .RN(n5712), .Q(\i_MIPS/PHT_2/history_state[0] ), .QN(\i_MIPS/PHT_2/n13 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[62]  ( .D(\i_MIPS/n395 ), .CK(clk), .RN(n5729), .Q(
        n3597), .QN(\i_MIPS/n267 ) );
  DFFRX1 \i_MIPS/Register/register_reg[31][19]  ( .D(n11526), .CK(clk), .RN(
        n5708), .QN(n272) );
  DFFRX1 \i_MIPS/Register/register_reg[31][30]  ( .D(n11515), .CK(clk), .RN(
        n5707), .QN(n265) );
  DFFRX1 \i_MIPS/ID_EX_reg[0]  ( .D(\i_MIPS/n528 ), .CK(clk), .RN(n5716), .Q(
        \i_MIPS/ID_EX_0 ), .QN(\i_MIPS/n372 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[68]  ( .D(\i_MIPS/n383 ), .CK(clk), .RN(n5730), .Q(
        \i_MIPS/ID_EX[68] ), .QN(\i_MIPS/n255 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[70]  ( .D(\i_MIPS/n379 ), .CK(clk), .RN(n5731), .Q(
        \i_MIPS/ID_EX[70] ), .QN(\i_MIPS/n251 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[66]  ( .D(\i_MIPS/n387 ), .CK(clk), .RN(n5730), .Q(
        \i_MIPS/ID_EX[66] ), .QN(\i_MIPS/n259 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[69]  ( .D(\i_MIPS/n381 ), .CK(clk), .RN(n5731), .Q(
        \i_MIPS/ID_EX[69] ), .QN(\i_MIPS/n253 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[71]  ( .D(\i_MIPS/n377 ), .CK(clk), .RN(n5731), .Q(
        n3598), .QN(\i_MIPS/n249 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[67]  ( .D(\i_MIPS/n385 ), .CK(clk), .RN(n5730), .Q(
        \i_MIPS/ID_EX[67] ), .QN(\i_MIPS/n257 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[104]  ( .D(\i_MIPS/n481 ), .CK(clk), .RN(n5742), 
        .Q(\i_MIPS/ID_EX[104] ), .QN(n4490) );
  DFFRX1 \i_MIPS/ID_EX_reg[97]  ( .D(\i_MIPS/n488 ), .CK(clk), .RN(n5741), .Q(
        \i_MIPS/ID_EX[97] ), .QN(n4489) );
  DFFRX1 \i_MIPS/ID_EX_reg[95]  ( .D(\i_MIPS/n490 ), .CK(clk), .RN(n5741), .Q(
        \i_MIPS/ID_EX[95] ), .QN(n4375) );
  DFFRX1 \i_MIPS/ID_EX_reg[94]  ( .D(\i_MIPS/n491 ), .CK(clk), .RN(n5741), .Q(
        \i_MIPS/ID_EX[94] ), .QN(n4491) );
  DFFRX1 \I_cache/cache_reg[4][154]  ( .D(n11551), .CK(clk), .RN(n5836), .Q(
        \I_cache/cache[4][154] ), .QN(n3334) );
  DFFRX1 \I_cache/cache_reg[5][154]  ( .D(n11550), .CK(clk), .RN(n5836), .Q(
        \I_cache/cache[5][154] ), .QN(n1727) );
  DFFRX1 \I_cache/cache_reg[0][154]  ( .D(n11555), .CK(clk), .RN(n5836), .Q(
        \I_cache/cache[0][154] ), .QN(n1724) );
  DFFRX1 \I_cache/cache_reg[2][154]  ( .D(n11553), .CK(clk), .RN(n5836), .Q(
        \I_cache/cache[2][154] ), .QN(n1725) );
  DFFRX1 \i_MIPS/Register/register_reg[29][19]  ( .D(\i_MIPS/Register/n199 ), 
        .CK(clk), .RN(n5722), .Q(\i_MIPS/Register/register[29][19] ), .QN(n417) );
  DFFRX1 \i_MIPS/Register/register_reg[29][30]  ( .D(\i_MIPS/Register/n210 ), 
        .CK(clk), .RN(n5721), .Q(\i_MIPS/Register/register[29][30] ), .QN(n423) );
  DFFRX1 \i_MIPS/Register/register_reg[28][27]  ( .D(\i_MIPS/Register/n239 ), 
        .CK(clk), .RN(n5719), .Q(\i_MIPS/Register/register[28][27] ), .QN(n286) );
  DFFRX1 \i_MIPS/Register/register_reg[27][19]  ( .D(\i_MIPS/Register/n263 ), 
        .CK(clk), .RN(n5717), .Q(\i_MIPS/Register/register[27][19] ), .QN(n318) );
  DFFRX1 \i_MIPS/Register/register_reg[27][30]  ( .D(\i_MIPS/Register/n274 ), 
        .CK(clk), .RN(n5776), .Q(\i_MIPS/Register/register[27][30] ), .QN(n421) );
  DFFRX1 \i_MIPS/Register/register_reg[25][19]  ( .D(\i_MIPS/Register/n327 ), 
        .CK(clk), .RN(n5771), .Q(\i_MIPS/Register/register[25][19] ), .QN(n320) );
  DFFRX1 \i_MIPS/Register/register_reg[25][30]  ( .D(\i_MIPS/Register/n338 ), 
        .CK(clk), .RN(n5770), .Q(\i_MIPS/Register/register[25][30] ), .QN(n426) );
  DFFRX1 \i_MIPS/Register/register_reg[24][27]  ( .D(\i_MIPS/Register/n367 ), 
        .CK(clk), .RN(n5768), .Q(\i_MIPS/Register/register[24][27] ), .QN(n275) );
  DFFRX1 \i_MIPS/Register/register_reg[23][19]  ( .D(\i_MIPS/Register/n391 ), 
        .CK(clk), .RN(n5786), .Q(\i_MIPS/Register/register[23][19] ), .QN(
        n2004) );
  DFFRX1 \i_MIPS/Register/register_reg[23][30]  ( .D(\i_MIPS/Register/n402 ), 
        .CK(clk), .RN(n5785), .Q(\i_MIPS/Register/register[23][30] ), .QN(
        n2011) );
  DFFRX1 \i_MIPS/Register/register_reg[21][19]  ( .D(\i_MIPS/Register/n455 ), 
        .CK(clk), .RN(n5781), .Q(\i_MIPS/Register/register[21][19] ), .QN(
        n2001) );
  DFFRX1 \i_MIPS/Register/register_reg[21][30]  ( .D(\i_MIPS/Register/n466 ), 
        .CK(clk), .RN(n5780), .Q(\i_MIPS/Register/register[21][30] ), .QN(
        n2002) );
  DFFRX1 \i_MIPS/Register/register_reg[20][27]  ( .D(\i_MIPS/Register/n495 ), 
        .CK(clk), .RN(n5777), .Q(\i_MIPS/Register/register[20][27] ), .QN(n431) );
  DFFRX1 \i_MIPS/Register/register_reg[19][19]  ( .D(\i_MIPS/Register/n519 ), 
        .CK(clk), .RN(n5755), .Q(\i_MIPS/Register/register[19][19] ), .QN(
        n2005) );
  DFFRX1 \i_MIPS/Register/register_reg[19][30]  ( .D(\i_MIPS/Register/n530 ), 
        .CK(clk), .RN(n5754), .Q(\i_MIPS/Register/register[19][30] ), .QN(
        n2012) );
  DFFRX1 \i_MIPS/Register/register_reg[17][19]  ( .D(\i_MIPS/Register/n583 ), 
        .CK(clk), .RN(n5750), .Q(\i_MIPS/Register/register[17][19] ), .QN(n428) );
  DFFRX1 \i_MIPS/Register/register_reg[17][30]  ( .D(\i_MIPS/Register/n594 ), 
        .CK(clk), .RN(n5749), .Q(\i_MIPS/Register/register[17][30] ), .QN(
        n2008) );
  DFFRX1 \i_MIPS/Register/register_reg[16][27]  ( .D(\i_MIPS/Register/n623 ), 
        .CK(clk), .RN(n5747), .Q(\i_MIPS/Register/register[16][27] ), .QN(n307) );
  DFFRX1 \i_MIPS/Register/register_reg[15][19]  ( .D(\i_MIPS/Register/n647 ), 
        .CK(clk), .RN(n5765), .Q(\i_MIPS/Register/register[15][19] ), .QN(n425) );
  DFFRX1 \i_MIPS/Register/register_reg[15][30]  ( .D(\i_MIPS/Register/n658 ), 
        .CK(clk), .RN(n5764), .Q(\i_MIPS/Register/register[15][30] ), .QN(n424) );
  DFFRX1 \i_MIPS/Register/register_reg[13][19]  ( .D(\i_MIPS/Register/n711 ), 
        .CK(clk), .RN(n5759), .Q(\i_MIPS/Register/register[13][19] ), .QN(n416) );
  DFFRX1 \i_MIPS/Register/register_reg[13][30]  ( .D(\i_MIPS/Register/n722 ), 
        .CK(clk), .RN(n5758), .Q(\i_MIPS/Register/register[13][30] ), .QN(n420) );
  DFFRX1 \i_MIPS/Register/register_reg[11][19]  ( .D(\i_MIPS/Register/n775 ), 
        .CK(clk), .RN(n5654), .Q(\i_MIPS/Register/register[11][19] ), .QN(n319) );
  DFFRX1 \i_MIPS/Register/register_reg[11][30]  ( .D(\i_MIPS/Register/n786 ), 
        .CK(clk), .RN(n5653), .Q(\i_MIPS/Register/register[11][30] ), .QN(n422) );
  DFFRX1 \i_MIPS/Register/register_reg[9][19]  ( .D(\i_MIPS/Register/n839 ), 
        .CK(clk), .RN(n5649), .Q(\i_MIPS/Register/register[9][19] ), .QN(n321)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][30]  ( .D(\i_MIPS/Register/n850 ), 
        .CK(clk), .RN(n5648), .Q(\i_MIPS/Register/register[9][30] ), .QN(n427)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][27]  ( .D(\i_MIPS/Register/n879 ), 
        .CK(clk), .RN(n5666), .Q(\i_MIPS/Register/register[8][27] ), .QN(n274)
         );
  DFFRX1 \i_MIPS/Register/register_reg[7][19]  ( .D(\i_MIPS/Register/n903 ), 
        .CK(clk), .RN(n5664), .Q(\i_MIPS/Register/register[7][19] ), .QN(n2006) );
  DFFRX1 \i_MIPS/Register/register_reg[7][30]  ( .D(\i_MIPS/Register/n914 ), 
        .CK(clk), .RN(n5663), .Q(\i_MIPS/Register/register[7][30] ), .QN(n2003) );
  DFFRX1 \i_MIPS/Register/register_reg[5][19]  ( .D(\i_MIPS/Register/n967 ), 
        .CK(clk), .RN(n5658), .Q(\i_MIPS/Register/register[5][19] ), .QN(n1977) );
  DFFRX1 \i_MIPS/Register/register_reg[5][30]  ( .D(\i_MIPS/Register/n978 ), 
        .CK(clk), .RN(n5657), .Q(\i_MIPS/Register/register[5][30] ), .QN(n2010) );
  DFFRX1 \i_MIPS/Register/register_reg[4][27]  ( .D(\i_MIPS/Register/n1007 ), 
        .CK(clk), .RN(n5635), .Q(\i_MIPS/Register/register[4][27] ), .QN(n430)
         );
  DFFRX1 \i_MIPS/Register/register_reg[3][19]  ( .D(\i_MIPS/Register/n1031 ), 
        .CK(clk), .RN(n5633), .Q(\i_MIPS/Register/register[3][19] ), .QN(n2007) );
  DFFRX1 \i_MIPS/Register/register_reg[3][30]  ( .D(\i_MIPS/Register/n1042 ), 
        .CK(clk), .RN(n5632), .Q(\i_MIPS/Register/register[3][30] ), .QN(n2013) );
  DFFRX1 \i_MIPS/Register/register_reg[1][19]  ( .D(\i_MIPS/Register/n1095 ), 
        .CK(clk), .RN(n5627), .Q(\i_MIPS/Register/register[1][19] ), .QN(n429)
         );
  DFFRX1 \i_MIPS/Register/register_reg[1][30]  ( .D(\i_MIPS/Register/n1106 ), 
        .CK(clk), .RN(n5631), .Q(\i_MIPS/Register/register[1][30] ), .QN(n2009) );
  DFFRX1 \i_MIPS/Register/register_reg[0][27]  ( .D(\i_MIPS/Register/n1135 ), 
        .CK(clk), .RN(n5644), .Q(\i_MIPS/Register/register[0][27] ), .QN(n306)
         );
  DFFRX1 \i_MIPS/Register/register_reg[31][0]  ( .D(n11545), .CK(clk), .RN(
        n5709), .Q(\i_MIPS/Register/register[31][0] ), .QN(n315) );
  DFFRX1 \i_MIPS/Register/register_reg[31][1]  ( .D(n11544), .CK(clk), .RN(
        n5709), .Q(\i_MIPS/Register/register[31][1] ), .QN(n281) );
  DFFRX1 \i_MIPS/Register/register_reg[31][2]  ( .D(n11543), .CK(clk), .RN(
        n5709), .Q(\i_MIPS/Register/register[31][2] ), .QN(n316) );
  DFFRX1 \i_MIPS/Register/register_reg[31][3]  ( .D(n11542), .CK(clk), .RN(
        n5709), .Q(\i_MIPS/Register/register[31][3] ), .QN(n268) );
  DFFRX1 \i_MIPS/Register/register_reg[31][4]  ( .D(n11541), .CK(clk), .RN(
        n5709), .Q(\i_MIPS/Register/register[31][4] ), .QN(n310) );
  DFFRX1 \i_MIPS/Register/register_reg[31][5]  ( .D(n11540), .CK(clk), .RN(
        n5709), .Q(\i_MIPS/Register/register[31][5] ), .QN(n277) );
  DFFRX1 \i_MIPS/Register/register_reg[31][6]  ( .D(n11539), .CK(clk), .RN(
        n5709), .Q(\i_MIPS/Register/register[31][6] ), .QN(n317) );
  DFFRX1 \i_MIPS/Register/register_reg[31][7]  ( .D(n11538), .CK(clk), .RN(
        n5709), .Q(\i_MIPS/Register/register[31][7] ), .QN(n280) );
  DFFRX1 \i_MIPS/Register/register_reg[31][8]  ( .D(n11537), .CK(clk), .RN(
        n5708), .Q(\i_MIPS/Register/register[31][8] ), .QN(n309) );
  DFFRX1 \i_MIPS/Register/register_reg[31][9]  ( .D(n11536), .CK(clk), .RN(
        n5708), .Q(\i_MIPS/Register/register[31][9] ), .QN(n276) );
  DFFRX1 \i_MIPS/Register/register_reg[31][10]  ( .D(n11535), .CK(clk), .RN(
        n5708), .Q(\i_MIPS/Register/register[31][10] ), .QN(n314) );
  DFFRX1 \i_MIPS/Register/register_reg[31][11]  ( .D(n11534), .CK(clk), .RN(
        n5708), .Q(\i_MIPS/Register/register[31][11] ), .QN(n313) );
  DFFRX1 \i_MIPS/Register/register_reg[31][12]  ( .D(n11533), .CK(clk), .RN(
        n5708), .Q(\i_MIPS/Register/register[31][12] ), .QN(n419) );
  DFFRX1 \i_MIPS/Register/register_reg[31][13]  ( .D(n11532), .CK(clk), .RN(
        n5708), .Q(\i_MIPS/Register/register[31][13] ), .QN(n283) );
  DFFRX1 \i_MIPS/Register/register_reg[31][14]  ( .D(n11531), .CK(clk), .RN(
        n5708), .Q(\i_MIPS/Register/register[31][14] ), .QN(n273) );
  DFFRX1 \i_MIPS/Register/register_reg[31][15]  ( .D(n11530), .CK(clk), .RN(
        n5708), .Q(\i_MIPS/Register/register[31][15] ), .QN(n312) );
  DFFRX1 \i_MIPS/Register/register_reg[31][16]  ( .D(n11529), .CK(clk), .RN(
        n5708), .Q(\i_MIPS/Register/register[31][16] ), .QN(n282) );
  DFFRX1 \i_MIPS/Register/register_reg[31][17]  ( .D(n11528), .CK(clk), .RN(
        n5708), .Q(\i_MIPS/Register/register[31][17] ), .QN(n279) );
  DFFRX1 \i_MIPS/Register/register_reg[31][18]  ( .D(n11527), .CK(clk), .RN(
        n5708), .Q(\i_MIPS/Register/register[31][18] ), .QN(n418) );
  DFFRX1 \i_MIPS/Register/register_reg[31][20]  ( .D(n11525), .CK(clk), .RN(
        n5707), .Q(\i_MIPS/Register/register[31][20] ), .QN(n305) );
  DFFRX1 \i_MIPS/Register/register_reg[31][21]  ( .D(n11524), .CK(clk), .RN(
        n5707), .Q(\i_MIPS/Register/register[31][21] ), .QN(n311) );
  DFFRX1 \i_MIPS/Register/register_reg[31][22]  ( .D(n11523), .CK(clk), .RN(
        n5707), .Q(\i_MIPS/Register/register[31][22] ), .QN(n266) );
  DFFRX1 \i_MIPS/Register/register_reg[31][23]  ( .D(n11522), .CK(clk), .RN(
        n5707), .Q(\i_MIPS/Register/register[31][23] ), .QN(n308) );
  DFFRX1 \i_MIPS/Register/register_reg[31][24]  ( .D(n11521), .CK(clk), .RN(
        n5707), .Q(\i_MIPS/Register/register[31][24] ), .QN(n271) );
  DFFRX1 \i_MIPS/Register/register_reg[31][25]  ( .D(n11520), .CK(clk), .RN(
        n5707), .Q(\i_MIPS/Register/register[31][25] ), .QN(n304) );
  DFFRX1 \i_MIPS/Register/register_reg[31][26]  ( .D(n11519), .CK(clk), .RN(
        n5707), .Q(\i_MIPS/Register/register[31][26] ), .QN(n267) );
  DFFRX1 \i_MIPS/Register/register_reg[31][28]  ( .D(n11517), .CK(clk), .RN(
        n5707), .Q(\i_MIPS/Register/register[31][28] ), .QN(n278) );
  DFFRX1 \i_MIPS/Register/register_reg[31][29]  ( .D(n11516), .CK(clk), .RN(
        n5707), .Q(\i_MIPS/Register/register[31][29] ), .QN(n284) );
  DFFRX1 \D_cache/cache_reg[1][0]  ( .D(\D_cache/n1794 ), .CK(clk), .RN(n5644), 
        .Q(\D_cache/cache[1][0] ), .QN(n1198) );
  DFFRX1 \D_cache/cache_reg[2][0]  ( .D(\D_cache/n1793 ), .CK(clk), .RN(n5643), 
        .Q(\D_cache/cache[2][0] ), .QN(n3078) );
  DFFRX1 \D_cache/cache_reg[4][0]  ( .D(\D_cache/n1791 ), .CK(clk), .RN(n5643), 
        .Q(\D_cache/cache[4][0] ), .QN(n1453) );
  DFFRX1 \D_cache/cache_reg[5][0]  ( .D(\D_cache/n1790 ), .CK(clk), .RN(n5643), 
        .Q(\D_cache/cache[5][0] ), .QN(n3023) );
  DFFRX1 \D_cache/cache_reg[6][0]  ( .D(\D_cache/n1789 ), .CK(clk), .RN(n5643), 
        .Q(\D_cache/cache[6][0] ), .QN(n2092) );
  DFFRX1 \D_cache/cache_reg[7][0]  ( .D(\D_cache/n1796 ), .CK(clk), .RN(n5643), 
        .Q(\D_cache/cache[7][0] ), .QN(n505) );
  DFFRX1 \D_cache/cache_reg[0][1]  ( .D(\D_cache/n1788 ), .CK(clk), .RN(n5643), 
        .Q(\D_cache/cache[0][1] ), .QN(n834) );
  DFFRX1 \D_cache/cache_reg[1][1]  ( .D(\D_cache/n1787 ), .CK(clk), .RN(n5643), 
        .Q(\D_cache/cache[1][1] ), .QN(n2397) );
  DFFRX1 \D_cache/cache_reg[2][1]  ( .D(\D_cache/n1786 ), .CK(clk), .RN(n5643), 
        .Q(\D_cache/cache[2][1] ), .QN(n2116) );
  DFFRX1 \D_cache/cache_reg[3][1]  ( .D(\D_cache/n1785 ), .CK(clk), .RN(n5643), 
        .Q(\D_cache/cache[3][1] ), .QN(n529) );
  DFFRX1 \D_cache/cache_reg[4][1]  ( .D(\D_cache/n1784 ), .CK(clk), .RN(n5643), 
        .Q(\D_cache/cache[4][1] ), .QN(n1377) );
  DFFRX1 \D_cache/cache_reg[5][1]  ( .D(\D_cache/n1783 ), .CK(clk), .RN(n5643), 
        .Q(\D_cache/cache[5][1] ), .QN(n2907) );
  DFFRX1 \D_cache/cache_reg[6][1]  ( .D(\D_cache/n1782 ), .CK(clk), .RN(n5642), 
        .Q(\D_cache/cache[6][1] ), .QN(n833) );
  DFFRX1 \D_cache/cache_reg[7][1]  ( .D(\D_cache/n1781 ), .CK(clk), .RN(n5642), 
        .Q(\D_cache/cache[7][1] ), .QN(n2396) );
  DFFRX1 \D_cache/cache_reg[0][2]  ( .D(\D_cache/n1780 ), .CK(clk), .RN(n5642), 
        .Q(\D_cache/cache[0][2] ), .QN(n1342) );
  DFFRX1 \D_cache/cache_reg[1][2]  ( .D(\D_cache/n1779 ), .CK(clk), .RN(n5642), 
        .Q(\D_cache/cache[1][2] ), .QN(n2871) );
  DFFRX1 \D_cache/cache_reg[2][2]  ( .D(\D_cache/n1778 ), .CK(clk), .RN(n5642), 
        .Q(\D_cache/cache[2][2] ), .QN(n1341) );
  DFFRX1 \D_cache/cache_reg[3][2]  ( .D(\D_cache/n1777 ), .CK(clk), .RN(n5642), 
        .Q(\D_cache/cache[3][2] ), .QN(n2870) );
  DFFRX1 \D_cache/cache_reg[4][2]  ( .D(\D_cache/n1776 ), .CK(clk), .RN(n5642), 
        .Q(\D_cache/cache[4][2] ), .QN(n1359) );
  DFFRX1 \D_cache/cache_reg[5][2]  ( .D(\D_cache/n1775 ), .CK(clk), .RN(n5642), 
        .Q(\D_cache/cache[5][2] ), .QN(n2889) );
  DFFRX1 \D_cache/cache_reg[6][2]  ( .D(\D_cache/n1774 ), .CK(clk), .RN(n5642), 
        .Q(\D_cache/cache[6][2] ), .QN(n1340) );
  DFFRX1 \D_cache/cache_reg[7][2]  ( .D(\D_cache/n1773 ), .CK(clk), .RN(n5642), 
        .Q(\D_cache/cache[7][2] ), .QN(n2869) );
  DFFRX1 \D_cache/cache_reg[0][3]  ( .D(\D_cache/n1772 ), .CK(clk), .RN(n5642), 
        .Q(\D_cache/cache[0][3] ), .QN(n1350) );
  DFFRX1 \D_cache/cache_reg[1][3]  ( .D(\D_cache/n1771 ), .CK(clk), .RN(n5642), 
        .Q(\D_cache/cache[1][3] ), .QN(n2880) );
  DFFRX1 \D_cache/cache_reg[2][3]  ( .D(\D_cache/n1770 ), .CK(clk), .RN(n5641), 
        .Q(\D_cache/cache[2][3] ), .QN(n1351) );
  DFFRX1 \D_cache/cache_reg[3][3]  ( .D(\D_cache/n1769 ), .CK(clk), .RN(n5641), 
        .Q(\D_cache/cache[3][3] ), .QN(n2881) );
  DFFRX1 \D_cache/cache_reg[4][3]  ( .D(\D_cache/n1768 ), .CK(clk), .RN(n5641), 
        .Q(\D_cache/cache[4][3] ), .QN(n3398) );
  DFFRX1 \D_cache/cache_reg[5][3]  ( .D(\D_cache/n1767 ), .CK(clk), .RN(n5641), 
        .Q(\D_cache/cache[5][3] ), .QN(n1769) );
  DFFRX1 \D_cache/cache_reg[6][3]  ( .D(\D_cache/n1766 ), .CK(clk), .RN(n5641), 
        .Q(\D_cache/cache[6][3] ), .QN(n2199) );
  DFFRX1 \D_cache/cache_reg[7][3]  ( .D(\D_cache/n1765 ), .CK(clk), .RN(n5641), 
        .Q(\D_cache/cache[7][3] ), .QN(n625) );
  DFFRX1 \D_cache/cache_reg[1][4]  ( .D(\D_cache/n1763 ), .CK(clk), .RN(n5641), 
        .Q(\D_cache/cache[1][4] ), .QN(n735) );
  DFFRX1 \D_cache/cache_reg[2][4]  ( .D(\D_cache/n1762 ), .CK(clk), .RN(n5641), 
        .Q(\D_cache/cache[2][4] ), .QN(n680) );
  DFFRX1 \D_cache/cache_reg[3][4]  ( .D(\D_cache/n1761 ), .CK(clk), .RN(n5641), 
        .Q(\D_cache/cache[3][4] ), .QN(n2252) );
  DFFRX1 \D_cache/cache_reg[4][4]  ( .D(\D_cache/n1760 ), .CK(clk), .RN(n5641), 
        .Q(\D_cache/cache[4][4] ), .QN(n681) );
  DFFRX1 \D_cache/cache_reg[5][4]  ( .D(\D_cache/n1759 ), .CK(clk), .RN(n5640), 
        .Q(\D_cache/cache[5][4] ), .QN(n2253) );
  DFFRX1 \D_cache/cache_reg[6][4]  ( .D(\D_cache/n1758 ), .CK(clk), .RN(n5640), 
        .Q(\D_cache/cache[6][4] ), .QN(n719) );
  DFFRX1 \D_cache/cache_reg[7][4]  ( .D(\D_cache/n1757 ), .CK(clk), .RN(n5640), 
        .Q(\D_cache/cache[7][4] ), .QN(n2287) );
  DFFRX1 \D_cache/cache_reg[0][5]  ( .D(\D_cache/n1756 ), .CK(clk), .RN(n5640), 
        .Q(\D_cache/cache[0][5] ), .QN(n3266) );
  DFFRX1 \D_cache/cache_reg[1][5]  ( .D(\D_cache/n1755 ), .CK(clk), .RN(n5640), 
        .Q(\D_cache/cache[1][5] ), .QN(n1426) );
  DFFRX1 \D_cache/cache_reg[2][5]  ( .D(\D_cache/n1754 ), .CK(clk), .RN(n5640), 
        .Q(\D_cache/cache[2][5] ), .QN(n1250) );
  DFFRX1 \D_cache/cache_reg[3][5]  ( .D(\D_cache/n1753 ), .CK(clk), .RN(n5640), 
        .Q(\D_cache/cache[3][5] ), .QN(n2792) );
  DFFRX1 \D_cache/cache_reg[4][5]  ( .D(\D_cache/n1752 ), .CK(clk), .RN(n5640), 
        .Q(\D_cache/cache[4][5] ), .QN(n1719) );
  DFFRX1 \D_cache/cache_reg[5][5]  ( .D(\D_cache/n1751 ), .CK(clk), .RN(n5640), 
        .Q(\D_cache/cache[5][5] ), .QN(n3317) );
  DFFRX1 \D_cache/cache_reg[6][5]  ( .D(\D_cache/n1750 ), .CK(clk), .RN(n5640), 
        .Q(\D_cache/cache[6][5] ), .QN(n829) );
  DFFRX1 \D_cache/cache_reg[7][5]  ( .D(\D_cache/n1749 ), .CK(clk), .RN(n5640), 
        .Q(\D_cache/cache[7][5] ), .QN(n2392) );
  DFFRX1 \D_cache/cache_reg[0][6]  ( .D(\D_cache/n1748 ), .CK(clk), .RN(n5640), 
        .Q(\D_cache/cache[0][6] ), .QN(n1353) );
  DFFRX1 \D_cache/cache_reg[1][6]  ( .D(\D_cache/n1747 ), .CK(clk), .RN(n5639), 
        .Q(\D_cache/cache[1][6] ), .QN(n2883) );
  DFFRX1 \D_cache/cache_reg[2][6]  ( .D(\D_cache/n1746 ), .CK(clk), .RN(n5639), 
        .Q(\D_cache/cache[2][6] ), .QN(n2190) );
  DFFRX1 \D_cache/cache_reg[3][6]  ( .D(\D_cache/n1745 ), .CK(clk), .RN(n5639), 
        .Q(\D_cache/cache[3][6] ), .QN(n616) );
  DFFRX1 \D_cache/cache_reg[4][6]  ( .D(\D_cache/n1744 ), .CK(clk), .RN(n5639), 
        .Q(\D_cache/cache[4][6] ), .QN(n3394) );
  DFFRX1 \D_cache/cache_reg[5][6]  ( .D(\D_cache/n1743 ), .CK(clk), .RN(n5639), 
        .Q(\D_cache/cache[5][6] ), .QN(n1765) );
  DFFRX1 \D_cache/cache_reg[6][6]  ( .D(\D_cache/n1742 ), .CK(clk), .RN(n5639), 
        .Q(\D_cache/cache[6][6] ), .QN(n2191) );
  DFFRX1 \D_cache/cache_reg[7][6]  ( .D(\D_cache/n1741 ), .CK(clk), .RN(n5639), 
        .Q(\D_cache/cache[7][6] ), .QN(n617) );
  DFFRX1 \D_cache/cache_reg[0][7]  ( .D(\D_cache/n1740 ), .CK(clk), .RN(n5639), 
        .Q(\D_cache/cache[0][7] ), .QN(n1268) );
  DFFRX1 \D_cache/cache_reg[1][7]  ( .D(\D_cache/n1739 ), .CK(clk), .RN(n5639), 
        .Q(\D_cache/cache[1][7] ), .QN(n2811) );
  DFFRX1 \D_cache/cache_reg[2][7]  ( .D(\D_cache/n1738 ), .CK(clk), .RN(n5639), 
        .Q(\D_cache/cache[2][7] ), .QN(n1267) );
  DFFRX1 \D_cache/cache_reg[3][7]  ( .D(\D_cache/n1737 ), .CK(clk), .RN(n5639), 
        .Q(\D_cache/cache[3][7] ), .QN(n2810) );
  DFFRX1 \D_cache/cache_reg[4][7]  ( .D(\D_cache/n1736 ), .CK(clk), .RN(n5639), 
        .Q(\D_cache/cache[4][7] ), .QN(n757) );
  DFFRX1 \D_cache/cache_reg[5][7]  ( .D(\D_cache/n1735 ), .CK(clk), .RN(n5638), 
        .Q(\D_cache/cache[5][7] ), .QN(n2318) );
  DFFRX1 \D_cache/cache_reg[6][7]  ( .D(\D_cache/n1734 ), .CK(clk), .RN(n5638), 
        .Q(\D_cache/cache[6][7] ), .QN(n2128) );
  DFFRX1 \D_cache/cache_reg[7][7]  ( .D(\D_cache/n1733 ), .CK(clk), .RN(n5638), 
        .Q(\D_cache/cache[7][7] ), .QN(n542) );
  DFFRX1 \D_cache/cache_reg[1][8]  ( .D(\D_cache/n1731 ), .CK(clk), .RN(n5638), 
        .Q(\D_cache/cache[1][8] ), .QN(n734) );
  DFFRX1 \D_cache/cache_reg[2][8]  ( .D(\D_cache/n1730 ), .CK(clk), .RN(n5638), 
        .Q(\D_cache/cache[2][8] ), .QN(n699) );
  DFFRX1 \D_cache/cache_reg[3][8]  ( .D(\D_cache/n1729 ), .CK(clk), .RN(n5638), 
        .Q(\D_cache/cache[3][8] ), .QN(n2268) );
  DFFRX1 \D_cache/cache_reg[4][8]  ( .D(\D_cache/n1728 ), .CK(clk), .RN(n5638), 
        .Q(\D_cache/cache[4][8] ), .QN(n1083) );
  DFFRX1 \D_cache/cache_reg[5][8]  ( .D(\D_cache/n1727 ), .CK(clk), .RN(n5638), 
        .Q(\D_cache/cache[5][8] ), .QN(n2676) );
  DFFRX1 \D_cache/cache_reg[6][8]  ( .D(\D_cache/n1726 ), .CK(clk), .RN(n5638), 
        .Q(\D_cache/cache[6][8] ), .QN(n718) );
  DFFRX1 \D_cache/cache_reg[7][8]  ( .D(\D_cache/n1725 ), .CK(clk), .RN(n5638), 
        .Q(\D_cache/cache[7][8] ), .QN(n2286) );
  DFFRX1 \D_cache/cache_reg[0][9]  ( .D(\D_cache/n1724 ), .CK(clk), .RN(n5638), 
        .Q(\D_cache/cache[0][9] ), .QN(n1293) );
  DFFRX1 \D_cache/cache_reg[1][9]  ( .D(\D_cache/n1723 ), .CK(clk), .RN(n5637), 
        .Q(\D_cache/cache[1][9] ), .QN(n2824) );
  DFFRX1 \D_cache/cache_reg[2][9]  ( .D(\D_cache/n1722 ), .CK(clk), .RN(n5637), 
        .Q(\D_cache/cache[2][9] ), .QN(n1258) );
  DFFRX1 \D_cache/cache_reg[3][9]  ( .D(\D_cache/n1721 ), .CK(clk), .RN(n5637), 
        .Q(\D_cache/cache[3][9] ), .QN(n2800) );
  DFFRX1 \D_cache/cache_reg[4][9]  ( .D(\D_cache/n1720 ), .CK(clk), .RN(n5637), 
        .Q(\D_cache/cache[4][9] ), .QN(n1376) );
  DFFRX1 \D_cache/cache_reg[5][9]  ( .D(\D_cache/n1719 ), .CK(clk), .RN(n5637), 
        .Q(\D_cache/cache[5][9] ), .QN(n2906) );
  DFFRX1 \D_cache/cache_reg[6][9]  ( .D(\D_cache/n1718 ), .CK(clk), .RN(n5637), 
        .Q(\D_cache/cache[6][9] ), .QN(n2133) );
  DFFRX1 \D_cache/cache_reg[7][9]  ( .D(\D_cache/n1717 ), .CK(clk), .RN(n5637), 
        .Q(\D_cache/cache[7][9] ), .QN(n547) );
  DFFRX1 \D_cache/cache_reg[0][10]  ( .D(\D_cache/n1716 ), .CK(clk), .RN(n5637), .Q(\D_cache/cache[0][10] ), .QN(n754) );
  DFFRX1 \D_cache/cache_reg[1][10]  ( .D(\D_cache/n1715 ), .CK(clk), .RN(n5637), .Q(\D_cache/cache[1][10] ), .QN(n2315) );
  DFFRX1 \D_cache/cache_reg[2][10]  ( .D(\D_cache/n1714 ), .CK(clk), .RN(n5637), .Q(\D_cache/cache[2][10] ), .QN(n1272) );
  DFFRX1 \D_cache/cache_reg[3][10]  ( .D(\D_cache/n1713 ), .CK(clk), .RN(n5637), .Q(\D_cache/cache[3][10] ), .QN(n2815) );
  DFFRX1 \D_cache/cache_reg[4][10]  ( .D(\D_cache/n1712 ), .CK(clk), .RN(n5637), .Q(\D_cache/cache[4][10] ), .QN(n2141) );
  DFFRX1 \D_cache/cache_reg[5][10]  ( .D(\D_cache/n1711 ), .CK(clk), .RN(n5641), .Q(\D_cache/cache[5][10] ), .QN(n561) );
  DFFRX1 \D_cache/cache_reg[6][10]  ( .D(\D_cache/n1710 ), .CK(clk), .RN(n5646), .Q(\D_cache/cache[6][10] ), .QN(n1271) );
  DFFRX1 \D_cache/cache_reg[7][10]  ( .D(\D_cache/n1709 ), .CK(clk), .RN(n5696), .Q(\D_cache/cache[7][10] ), .QN(n2814) );
  DFFRX1 \D_cache/cache_reg[0][11]  ( .D(\D_cache/n1708 ), .CK(clk), .RN(n5696), .Q(\D_cache/cache[0][11] ), .QN(n1077) );
  DFFRX1 \D_cache/cache_reg[1][11]  ( .D(\D_cache/n1707 ), .CK(clk), .RN(n5696), .Q(\D_cache/cache[1][11] ), .QN(n2809) );
  DFFRX1 \D_cache/cache_reg[2][11]  ( .D(\D_cache/n1706 ), .CK(clk), .RN(n5696), .Q(\D_cache/cache[2][11] ), .QN(n1266) );
  DFFRX1 \D_cache/cache_reg[3][11]  ( .D(\D_cache/n1705 ), .CK(clk), .RN(n5696), .Q(\D_cache/cache[3][11] ), .QN(n2808) );
  DFFRX1 \D_cache/cache_reg[4][11]  ( .D(\D_cache/n1704 ), .CK(clk), .RN(n5696), .Q(\D_cache/cache[4][11] ), .QN(n1365) );
  DFFRX1 \D_cache/cache_reg[5][11]  ( .D(\D_cache/n1703 ), .CK(clk), .RN(n5696), .Q(\D_cache/cache[5][11] ), .QN(n2895) );
  DFFRX1 \D_cache/cache_reg[6][11]  ( .D(\D_cache/n1702 ), .CK(clk), .RN(n5696), .Q(\D_cache/cache[6][11] ), .QN(n1265) );
  DFFRX1 \D_cache/cache_reg[7][11]  ( .D(\D_cache/n1701 ), .CK(clk), .RN(n5696), .Q(\D_cache/cache[7][11] ), .QN(n2807) );
  DFFRX1 \D_cache/cache_reg[0][12]  ( .D(\D_cache/n1700 ), .CK(clk), .RN(n5696), .Q(\D_cache/cache[0][12] ), .QN(n838) );
  DFFRX1 \D_cache/cache_reg[1][12]  ( .D(\D_cache/n1699 ), .CK(clk), .RN(n5696), .Q(\D_cache/cache[1][12] ), .QN(n2401) );
  DFFRX1 \D_cache/cache_reg[2][12]  ( .D(\D_cache/n1698 ), .CK(clk), .RN(n5695), .Q(\D_cache/cache[2][12] ), .QN(n748) );
  DFFRX1 \D_cache/cache_reg[3][12]  ( .D(\D_cache/n1697 ), .CK(clk), .RN(n5695), .Q(\D_cache/cache[3][12] ), .QN(n2309) );
  DFFRX1 \D_cache/cache_reg[4][12]  ( .D(\D_cache/n1696 ), .CK(clk), .RN(n5695), .Q(\D_cache/cache[4][12] ), .QN(n778) );
  DFFRX1 \D_cache/cache_reg[5][12]  ( .D(\D_cache/n1695 ), .CK(clk), .RN(n5695), .Q(\D_cache/cache[5][12] ), .QN(n2340) );
  DFFRX1 \D_cache/cache_reg[6][12]  ( .D(\D_cache/n1694 ), .CK(clk), .RN(n5695), .Q(\D_cache/cache[6][12] ), .QN(n837) );
  DFFRX1 \D_cache/cache_reg[7][12]  ( .D(\D_cache/n1693 ), .CK(clk), .RN(n5695), .Q(\D_cache/cache[7][12] ), .QN(n2400) );
  DFFRX1 \D_cache/cache_reg[1][13]  ( .D(\D_cache/n1691 ), .CK(clk), .RN(n5695), .Q(\D_cache/cache[1][13] ), .QN(n1278) );
  DFFRX1 \D_cache/cache_reg[2][13]  ( .D(\D_cache/n1690 ), .CK(clk), .RN(n5695), .Q(\D_cache/cache[2][13] ), .QN(n1262) );
  DFFRX1 \D_cache/cache_reg[3][13]  ( .D(\D_cache/n1689 ), .CK(clk), .RN(n5695), .Q(\D_cache/cache[3][13] ), .QN(n2804) );
  DFFRX1 \D_cache/cache_reg[4][13]  ( .D(\D_cache/n1688 ), .CK(clk), .RN(n5695), .Q(\D_cache/cache[4][13] ), .QN(n2106) );
  DFFRX1 \D_cache/cache_reg[5][13]  ( .D(\D_cache/n1687 ), .CK(clk), .RN(n5695), .Q(\D_cache/cache[5][13] ), .QN(n512) );
  DFFRX1 \D_cache/cache_reg[6][13]  ( .D(\D_cache/n1686 ), .CK(clk), .RN(n5694), .Q(\D_cache/cache[6][13] ), .QN(n747) );
  DFFRX1 \D_cache/cache_reg[7][13]  ( .D(\D_cache/n1685 ), .CK(clk), .RN(n5694), .Q(\D_cache/cache[7][13] ), .QN(n2308) );
  DFFRX1 \D_cache/cache_reg[1][14]  ( .D(\D_cache/n1683 ), .CK(clk), .RN(n5694), .Q(\D_cache/cache[1][14] ), .QN(n1181) );
  DFFRX1 \D_cache/cache_reg[2][14]  ( .D(\D_cache/n1682 ), .CK(clk), .RN(n5694), .Q(\D_cache/cache[2][14] ), .QN(n1264) );
  DFFRX1 \D_cache/cache_reg[3][14]  ( .D(\D_cache/n1681 ), .CK(clk), .RN(n5694), .Q(\D_cache/cache[3][14] ), .QN(n2806) );
  DFFRX1 \D_cache/cache_reg[4][14]  ( .D(\D_cache/n1680 ), .CK(clk), .RN(n5694), .Q(\D_cache/cache[4][14] ), .QN(n2772) );
  DFFRX1 \D_cache/cache_reg[5][14]  ( .D(\D_cache/n1679 ), .CK(clk), .RN(n5694), .Q(\D_cache/cache[5][14] ), .QN(n1201) );
  DFFRX1 \D_cache/cache_reg[6][14]  ( .D(\D_cache/n1678 ), .CK(clk), .RN(n5694), .Q(\D_cache/cache[6][14] ), .QN(n1263) );
  DFFRX1 \D_cache/cache_reg[7][14]  ( .D(\D_cache/n1677 ), .CK(clk), .RN(n5694), .Q(\D_cache/cache[7][14] ), .QN(n2805) );
  DFFRX1 \D_cache/cache_reg[0][15]  ( .D(\D_cache/n1676 ), .CK(clk), .RN(n5694), .Q(\D_cache/cache[0][15] ), .QN(n842) );
  DFFRX1 \D_cache/cache_reg[1][15]  ( .D(\D_cache/n1675 ), .CK(clk), .RN(n5694), .Q(\D_cache/cache[1][15] ), .QN(n2405) );
  DFFRX1 \D_cache/cache_reg[2][15]  ( .D(\D_cache/n1674 ), .CK(clk), .RN(n5693), .Q(\D_cache/cache[2][15] ), .QN(n1259) );
  DFFRX1 \D_cache/cache_reg[3][15]  ( .D(\D_cache/n1673 ), .CK(clk), .RN(n5693), .Q(\D_cache/cache[3][15] ), .QN(n2801) );
  DFFRX1 \D_cache/cache_reg[4][15]  ( .D(\D_cache/n1672 ), .CK(clk), .RN(n5693), .Q(\D_cache/cache[4][15] ), .QN(n1364) );
  DFFRX1 \D_cache/cache_reg[5][15]  ( .D(\D_cache/n1671 ), .CK(clk), .RN(n5693), .Q(\D_cache/cache[5][15] ), .QN(n2894) );
  DFFRX1 \D_cache/cache_reg[6][15]  ( .D(\D_cache/n1670 ), .CK(clk), .RN(n5693), .Q(\D_cache/cache[6][15] ), .QN(n841) );
  DFFRX1 \D_cache/cache_reg[7][15]  ( .D(\D_cache/n1669 ), .CK(clk), .RN(n5693), .Q(\D_cache/cache[7][15] ), .QN(n2404) );
  DFFRX1 \D_cache/cache_reg[0][16]  ( .D(\D_cache/n1668 ), .CK(clk), .RN(n5693), .Q(\D_cache/cache[0][16] ), .QN(n1159) );
  DFFRX1 \D_cache/cache_reg[1][16]  ( .D(\D_cache/n1667 ), .CK(clk), .RN(n5693), .Q(\D_cache/cache[1][16] ), .QN(n2879) );
  DFFRX1 \D_cache/cache_reg[2][16]  ( .D(\D_cache/n1666 ), .CK(clk), .RN(n5693), .Q(\D_cache/cache[2][16] ), .QN(n2115) );
  DFFRX1 \D_cache/cache_reg[3][16]  ( .D(\D_cache/n1665 ), .CK(clk), .RN(n5693), .Q(\D_cache/cache[3][16] ), .QN(n528) );
  DFFRX1 \D_cache/cache_reg[4][16]  ( .D(\D_cache/n1664 ), .CK(clk), .RN(n5693), .Q(\D_cache/cache[4][16] ), .QN(n2126) );
  DFFRX1 \D_cache/cache_reg[5][16]  ( .D(\D_cache/n1663 ), .CK(clk), .RN(n5693), .Q(\D_cache/cache[5][16] ), .QN(n539) );
  DFFRX1 \D_cache/cache_reg[6][16]  ( .D(\D_cache/n1662 ), .CK(clk), .RN(n5692), .Q(\D_cache/cache[6][16] ), .QN(n2135) );
  DFFRX1 \D_cache/cache_reg[7][16]  ( .D(\D_cache/n1661 ), .CK(clk), .RN(n5692), .Q(\D_cache/cache[7][16] ), .QN(n550) );
  DFFRX1 \D_cache/cache_reg[0][17]  ( .D(\D_cache/n1660 ), .CK(clk), .RN(n5692), .Q(\D_cache/cache[0][17] ), .QN(n1182) );
  DFFRX1 \D_cache/cache_reg[1][17]  ( .D(\D_cache/n1659 ), .CK(clk), .RN(n5692), .Q(\D_cache/cache[1][17] ), .QN(n2950) );
  DFFRX1 \D_cache/cache_reg[2][17]  ( .D(\D_cache/n1658 ), .CK(clk), .RN(n5692), .Q(\D_cache/cache[2][17] ), .QN(n1418) );
  DFFRX1 \D_cache/cache_reg[3][17]  ( .D(\D_cache/n1657 ), .CK(clk), .RN(n5692), .Q(\D_cache/cache[3][17] ), .QN(n2949) );
  DFFRX1 \D_cache/cache_reg[4][17]  ( .D(\D_cache/n1656 ), .CK(clk), .RN(n5692), .Q(\D_cache/cache[4][17] ), .QN(n1712) );
  DFFRX1 \D_cache/cache_reg[5][17]  ( .D(\D_cache/n1655 ), .CK(clk), .RN(n5692), .Q(\D_cache/cache[5][17] ), .QN(n3309) );
  DFFRX1 \D_cache/cache_reg[6][17]  ( .D(\D_cache/n1654 ), .CK(clk), .RN(n5692), .Q(\D_cache/cache[6][17] ), .QN(n1217) );
  DFFRX1 \D_cache/cache_reg[7][17]  ( .D(\D_cache/n1653 ), .CK(clk), .RN(n5692), .Q(\D_cache/cache[7][17] ), .QN(n2754) );
  DFFRX1 \D_cache/cache_reg[0][18]  ( .D(\D_cache/n1652 ), .CK(clk), .RN(n5692), .Q(\D_cache/cache[0][18] ), .QN(n1292) );
  DFFRX1 \D_cache/cache_reg[1][18]  ( .D(\D_cache/n1651 ), .CK(clk), .RN(n5692), .Q(\D_cache/cache[1][18] ), .QN(n2823) );
  DFFRX1 \D_cache/cache_reg[2][18]  ( .D(\D_cache/n1650 ), .CK(clk), .RN(n5691), .Q(\D_cache/cache[2][18] ), .QN(n1270) );
  DFFRX1 \D_cache/cache_reg[3][18]  ( .D(\D_cache/n1649 ), .CK(clk), .RN(n5691), .Q(\D_cache/cache[3][18] ), .QN(n2813) );
  DFFRX1 \D_cache/cache_reg[4][18]  ( .D(\D_cache/n1648 ), .CK(clk), .RN(n5691), .Q(\D_cache/cache[4][18] ), .QN(n1711) );
  DFFRX1 \D_cache/cache_reg[5][18]  ( .D(\D_cache/n1647 ), .CK(clk), .RN(n5691), .Q(\D_cache/cache[5][18] ), .QN(n3308) );
  DFFRX1 \D_cache/cache_reg[6][18]  ( .D(\D_cache/n1646 ), .CK(clk), .RN(n5691), .Q(\D_cache/cache[6][18] ), .QN(n1269) );
  DFFRX1 \D_cache/cache_reg[7][18]  ( .D(\D_cache/n1645 ), .CK(clk), .RN(n5691), .Q(\D_cache/cache[7][18] ), .QN(n2812) );
  DFFRX1 \D_cache/cache_reg[1][19]  ( .D(\D_cache/n1643 ), .CK(clk), .RN(n5691), .Q(\D_cache/cache[1][19] ), .QN(n725) );
  DFFRX1 \D_cache/cache_reg[2][19]  ( .D(\D_cache/n1642 ), .CK(clk), .RN(n5691), .Q(\D_cache/cache[2][19] ), .QN(n1087) );
  DFFRX1 \D_cache/cache_reg[3][19]  ( .D(\D_cache/n1641 ), .CK(clk), .RN(n5691), .Q(\D_cache/cache[3][19] ), .QN(n2682) );
  DFFRX1 \D_cache/cache_reg[4][19]  ( .D(\D_cache/n1640 ), .CK(clk), .RN(n5691), .Q(\D_cache/cache[4][19] ), .QN(n1160) );
  DFFRX1 \D_cache/cache_reg[5][19]  ( .D(\D_cache/n1639 ), .CK(clk), .RN(n5690), .Q(\D_cache/cache[5][19] ), .QN(n2716) );
  DFFRX1 \D_cache/cache_reg[6][19]  ( .D(\D_cache/n1638 ), .CK(clk), .RN(n5690), .Q(\D_cache/cache[6][19] ), .QN(n2081) );
  DFFRX1 \D_cache/cache_reg[7][19]  ( .D(\D_cache/n1637 ), .CK(clk), .RN(n5690), .Q(\D_cache/cache[7][19] ), .QN(n493) );
  DFFRX1 \D_cache/cache_reg[1][20]  ( .D(\D_cache/n1635 ), .CK(clk), .RN(n5690), .Q(\D_cache/cache[1][20] ), .QN(n1424) );
  DFFRX1 \D_cache/cache_reg[2][20]  ( .D(\D_cache/n1634 ), .CK(clk), .RN(n5690), .Q(\D_cache/cache[2][20] ), .QN(n1349) );
  DFFRX1 \D_cache/cache_reg[3][20]  ( .D(\D_cache/n1633 ), .CK(clk), .RN(n5690), .Q(\D_cache/cache[3][20] ), .QN(n2878) );
  DFFRX1 \D_cache/cache_reg[4][20]  ( .D(\D_cache/n1632 ), .CK(clk), .RN(n5690), .Q(\D_cache/cache[4][20] ), .QN(n3270) );
  DFFRX1 \D_cache/cache_reg[5][20]  ( .D(\D_cache/n1631 ), .CK(clk), .RN(n5690), .Q(\D_cache/cache[5][20] ), .QN(n1635) );
  DFFRX1 \D_cache/cache_reg[6][20]  ( .D(\D_cache/n1630 ), .CK(clk), .RN(n5690), .Q(\D_cache/cache[6][20] ), .QN(n1157) );
  DFFRX1 \D_cache/cache_reg[7][20]  ( .D(\D_cache/n1629 ), .CK(clk), .RN(n5690), .Q(\D_cache/cache[7][20] ), .QN(n2714) );
  DFFRX1 \D_cache/cache_reg[2][21]  ( .D(\D_cache/n1626 ), .CK(clk), .RN(n5689), .Q(\D_cache/cache[2][21] ), .QN(n1112) );
  DFFRX1 \D_cache/cache_reg[3][21]  ( .D(\D_cache/n1625 ), .CK(clk), .RN(n5689), .Q(\D_cache/cache[3][21] ), .QN(n2701) );
  DFFRX1 \D_cache/cache_reg[4][21]  ( .D(\D_cache/n1624 ), .CK(clk), .RN(n5689), .Q(\D_cache/cache[4][21] ), .QN(n1622) );
  DFFRX1 \D_cache/cache_reg[5][21]  ( .D(\D_cache/n1623 ), .CK(clk), .RN(n5689), .Q(\D_cache/cache[5][21] ), .QN(n3199) );
  DFFRX1 \D_cache/cache_reg[6][21]  ( .D(\D_cache/n1622 ), .CK(clk), .RN(n5689), .Q(\D_cache/cache[6][21] ), .QN(n1076) );
  DFFRX1 \D_cache/cache_reg[7][21]  ( .D(\D_cache/n1621 ), .CK(clk), .RN(n5689), .Q(\D_cache/cache[7][21] ), .QN(n2653) );
  DFFRX1 \D_cache/cache_reg[0][22]  ( .D(\D_cache/n1620 ), .CK(clk), .RN(n5689), .Q(\D_cache/cache[0][22] ), .QN(n650) );
  DFFRX1 \D_cache/cache_reg[1][22]  ( .D(\D_cache/n1619 ), .CK(clk), .RN(n5689), .Q(\D_cache/cache[1][22] ), .QN(n2227) );
  DFFRX1 \D_cache/cache_reg[2][22]  ( .D(\D_cache/n1618 ), .CK(clk), .RN(n5689), .Q(\D_cache/cache[2][22] ), .QN(n1260) );
  DFFRX1 \D_cache/cache_reg[3][22]  ( .D(\D_cache/n1617 ), .CK(clk), .RN(n5689), .Q(\D_cache/cache[3][22] ), .QN(n2802) );
  DFFRX1 \D_cache/cache_reg[4][22]  ( .D(\D_cache/n1616 ), .CK(clk), .RN(n5689), .Q(\D_cache/cache[4][22] ), .QN(n1718) );
  DFFRX1 \D_cache/cache_reg[5][22]  ( .D(\D_cache/n1615 ), .CK(clk), .RN(n5688), .Q(\D_cache/cache[5][22] ), .QN(n3316) );
  DFFRX1 \D_cache/cache_reg[6][22]  ( .D(\D_cache/n1614 ), .CK(clk), .RN(n5688), .Q(\D_cache/cache[6][22] ), .QN(n843) );
  DFFRX1 \D_cache/cache_reg[7][22]  ( .D(\D_cache/n1613 ), .CK(clk), .RN(n5688), .Q(\D_cache/cache[7][22] ), .QN(n2406) );
  DFFRX1 \D_cache/cache_reg[1][23]  ( .D(\D_cache/n1611 ), .CK(clk), .RN(n5688), .Q(\D_cache/cache[1][23] ), .QN(n1196) );
  DFFRX1 \D_cache/cache_reg[2][23]  ( .D(\D_cache/n1610 ), .CK(clk), .RN(n5688), .Q(\D_cache/cache[2][23] ), .QN(n697) );
  DFFRX1 \D_cache/cache_reg[3][23]  ( .D(\D_cache/n1609 ), .CK(clk), .RN(n5688), .Q(\D_cache/cache[3][23] ), .QN(n2266) );
  DFFRX1 \D_cache/cache_reg[4][23]  ( .D(\D_cache/n1608 ), .CK(clk), .RN(n5688), .Q(\D_cache/cache[4][23] ), .QN(n2090) );
  DFFRX1 \D_cache/cache_reg[5][23]  ( .D(\D_cache/n1607 ), .CK(clk), .RN(n5688), .Q(\D_cache/cache[5][23] ), .QN(n503) );
  DFFRX1 \D_cache/cache_reg[6][23]  ( .D(\D_cache/n1606 ), .CK(clk), .RN(n5688), .Q(\D_cache/cache[6][23] ), .QN(n696) );
  DFFRX1 \D_cache/cache_reg[7][23]  ( .D(\D_cache/n1605 ), .CK(clk), .RN(n5688), .Q(\D_cache/cache[7][23] ), .QN(n2265) );
  DFFRX1 \D_cache/cache_reg[0][24]  ( .D(\D_cache/n1604 ), .CK(clk), .RN(n5688), .Q(\D_cache/cache[0][24] ), .QN(n836) );
  DFFRX1 \D_cache/cache_reg[1][24]  ( .D(\D_cache/n1603 ), .CK(clk), .RN(n5687), .Q(\D_cache/cache[1][24] ), .QN(n2399) );
  DFFRX1 \D_cache/cache_reg[2][24]  ( .D(\D_cache/n1602 ), .CK(clk), .RN(n5687), .Q(\D_cache/cache[2][24] ), .QN(n1256) );
  DFFRX1 \D_cache/cache_reg[3][24]  ( .D(\D_cache/n1601 ), .CK(clk), .RN(n5687), .Q(\D_cache/cache[3][24] ), .QN(n2798) );
  DFFRX1 \D_cache/cache_reg[4][24]  ( .D(\D_cache/n1600 ), .CK(clk), .RN(n5687), .Q(\D_cache/cache[4][24] ), .QN(n1374) );
  DFFRX1 \D_cache/cache_reg[5][24]  ( .D(\D_cache/n1599 ), .CK(clk), .RN(n5687), .Q(\D_cache/cache[5][24] ), .QN(n2904) );
  DFFRX1 \D_cache/cache_reg[6][24]  ( .D(\D_cache/n1598 ), .CK(clk), .RN(n5687), .Q(\D_cache/cache[6][24] ), .QN(n835) );
  DFFRX1 \D_cache/cache_reg[7][24]  ( .D(\D_cache/n1597 ), .CK(clk), .RN(n5687), .Q(\D_cache/cache[7][24] ), .QN(n2398) );
  DFFRX1 \D_cache/cache_reg[0][25]  ( .D(\D_cache/n1596 ), .CK(clk), .RN(n5687), .Q(\D_cache/cache[0][25] ), .QN(n840) );
  DFFRX1 \D_cache/cache_reg[1][25]  ( .D(\D_cache/n1595 ), .CK(clk), .RN(n5687), .Q(\D_cache/cache[1][25] ), .QN(n2403) );
  DFFRX1 \D_cache/cache_reg[2][25]  ( .D(\D_cache/n1594 ), .CK(clk), .RN(n5687), .Q(\D_cache/cache[2][25] ), .QN(n1257) );
  DFFRX1 \D_cache/cache_reg[3][25]  ( .D(\D_cache/n1593 ), .CK(clk), .RN(n5687), .Q(\D_cache/cache[3][25] ), .QN(n2799) );
  DFFRX1 \D_cache/cache_reg[4][25]  ( .D(\D_cache/n1592 ), .CK(clk), .RN(n5687), .Q(\D_cache/cache[4][25] ), .QN(n1212) );
  DFFRX1 \D_cache/cache_reg[5][25]  ( .D(\D_cache/n1591 ), .CK(clk), .RN(n5686), .Q(\D_cache/cache[5][25] ), .QN(n2749) );
  DFFRX1 \D_cache/cache_reg[6][25]  ( .D(\D_cache/n1590 ), .CK(clk), .RN(n5691), .Q(\D_cache/cache[6][25] ), .QN(n839) );
  DFFRX1 \D_cache/cache_reg[7][25]  ( .D(\D_cache/n1589 ), .CK(clk), .RN(n5706), .Q(\D_cache/cache[7][25] ), .QN(n2402) );
  DFFRX1 \D_cache/cache_reg[0][26]  ( .D(\D_cache/n1588 ), .CK(clk), .RN(n5706), .Q(\D_cache/cache[0][26] ), .QN(n702) );
  DFFRX1 \D_cache/cache_reg[1][26]  ( .D(\D_cache/n1587 ), .CK(clk), .RN(n5706), .Q(\D_cache/cache[1][26] ), .QN(n2357) );
  DFFRX1 \D_cache/cache_reg[2][26]  ( .D(\D_cache/n1586 ), .CK(clk), .RN(n5706), .Q(\D_cache/cache[2][26] ), .QN(n1232) );
  DFFRX1 \D_cache/cache_reg[3][26]  ( .D(\D_cache/n1585 ), .CK(clk), .RN(n5706), .Q(\D_cache/cache[3][26] ), .QN(n2773) );
  DFFRX1 \D_cache/cache_reg[4][26]  ( .D(\D_cache/n1584 ), .CK(clk), .RN(n5706), .Q(\D_cache/cache[4][26] ), .QN(n1363) );
  DFFRX1 \D_cache/cache_reg[5][26]  ( .D(\D_cache/n1583 ), .CK(clk), .RN(n5706), .Q(\D_cache/cache[5][26] ), .QN(n2893) );
  DFFRX1 \D_cache/cache_reg[6][26]  ( .D(\D_cache/n1582 ), .CK(clk), .RN(n5706), .Q(\D_cache/cache[6][26] ), .QN(n2291) );
  DFFRX1 \D_cache/cache_reg[7][26]  ( .D(\D_cache/n1581 ), .CK(clk), .RN(n5706), .Q(\D_cache/cache[7][26] ), .QN(n726) );
  DFFRX1 \D_cache/cache_reg[0][27]  ( .D(\D_cache/n1580 ), .CK(clk), .RN(n5706), .Q(\D_cache/cache[0][27] ), .QN(n832) );
  DFFRX1 \D_cache/cache_reg[1][27]  ( .D(\D_cache/n1579 ), .CK(clk), .RN(n5705), .Q(\D_cache/cache[1][27] ), .QN(n2395) );
  DFFRX1 \D_cache/cache_reg[2][27]  ( .D(\D_cache/n1578 ), .CK(clk), .RN(n5705), .Q(\D_cache/cache[2][27] ), .QN(n831) );
  DFFRX1 \D_cache/cache_reg[3][27]  ( .D(\D_cache/n1577 ), .CK(clk), .RN(n5705), .Q(\D_cache/cache[3][27] ), .QN(n2394) );
  DFFRX1 \D_cache/cache_reg[4][27]  ( .D(\D_cache/n1576 ), .CK(clk), .RN(n5705), .Q(\D_cache/cache[4][27] ), .QN(n1380) );
  DFFRX1 \D_cache/cache_reg[5][27]  ( .D(\D_cache/n1575 ), .CK(clk), .RN(n5705), .Q(\D_cache/cache[5][27] ), .QN(n2910) );
  DFFRX1 \D_cache/cache_reg[6][27]  ( .D(\D_cache/n1574 ), .CK(clk), .RN(n5705), .Q(\D_cache/cache[6][27] ), .QN(n830) );
  DFFRX1 \D_cache/cache_reg[7][27]  ( .D(\D_cache/n1573 ), .CK(clk), .RN(n5705), .Q(\D_cache/cache[7][27] ), .QN(n2393) );
  DFFRX1 \D_cache/cache_reg[1][28]  ( .D(\D_cache/n1571 ), .CK(clk), .RN(n5705), .Q(\D_cache/cache[1][28] ), .QN(n500) );
  DFFRX1 \D_cache/cache_reg[2][28]  ( .D(\D_cache/n1570 ), .CK(clk), .RN(n5705), .Q(\D_cache/cache[2][28] ), .QN(n1158) );
  DFFRX1 \D_cache/cache_reg[3][28]  ( .D(\D_cache/n1569 ), .CK(clk), .RN(n5705), .Q(\D_cache/cache[3][28] ), .QN(n2715) );
  DFFRX1 \D_cache/cache_reg[4][28]  ( .D(\D_cache/n1568 ), .CK(clk), .RN(n5705), .Q(\D_cache/cache[4][28] ), .QN(n2077) );
  DFFRX1 \D_cache/cache_reg[5][28]  ( .D(\D_cache/n1567 ), .CK(clk), .RN(n5704), .Q(\D_cache/cache[5][28] ), .QN(n489) );
  DFFRX1 \D_cache/cache_reg[6][28]  ( .D(\D_cache/n1566 ), .CK(clk), .RN(n5704), .Q(\D_cache/cache[6][28] ), .QN(n686) );
  DFFRX1 \D_cache/cache_reg[7][28]  ( .D(\D_cache/n1565 ), .CK(clk), .RN(n5704), .Q(\D_cache/cache[7][28] ), .QN(n2258) );
  DFFRX1 \D_cache/cache_reg[0][29]  ( .D(\D_cache/n1564 ), .CK(clk), .RN(n5704), .Q(\D_cache/cache[0][29] ), .QN(n796) );
  DFFRX1 \D_cache/cache_reg[1][29]  ( .D(\D_cache/n1563 ), .CK(clk), .RN(n5704), .Q(\D_cache/cache[1][29] ), .QN(n2359) );
  DFFRX1 \D_cache/cache_reg[2][29]  ( .D(\D_cache/n1562 ), .CK(clk), .RN(n5704), .Q(\D_cache/cache[2][29] ), .QN(n1233) );
  DFFRX1 \D_cache/cache_reg[3][29]  ( .D(\D_cache/n1561 ), .CK(clk), .RN(n5704), .Q(\D_cache/cache[3][29] ), .QN(n2774) );
  DFFRX1 \D_cache/cache_reg[4][29]  ( .D(\D_cache/n1560 ), .CK(clk), .RN(n5704), .Q(\D_cache/cache[4][29] ), .QN(n1379) );
  DFFRX1 \D_cache/cache_reg[5][29]  ( .D(\D_cache/n1559 ), .CK(clk), .RN(n5704), .Q(\D_cache/cache[5][29] ), .QN(n2909) );
  DFFRX1 \D_cache/cache_reg[6][29]  ( .D(\D_cache/n1558 ), .CK(clk), .RN(n5704), .Q(\D_cache/cache[6][29] ), .QN(n795) );
  DFFRX1 \D_cache/cache_reg[7][29]  ( .D(\D_cache/n1557 ), .CK(clk), .RN(n5704), .Q(\D_cache/cache[7][29] ), .QN(n2358) );
  DFFRX1 \D_cache/cache_reg[1][30]  ( .D(\D_cache/n1555 ), .CK(clk), .RN(n5703), .Q(\D_cache/cache[1][30] ), .QN(n1180) );
  DFFRX1 \D_cache/cache_reg[2][30]  ( .D(\D_cache/n1554 ), .CK(clk), .RN(n5703), .Q(\D_cache/cache[2][30] ), .QN(n717) );
  DFFRX1 \D_cache/cache_reg[3][30]  ( .D(\D_cache/n1553 ), .CK(clk), .RN(n5703), .Q(\D_cache/cache[3][30] ), .QN(n2285) );
  DFFRX1 \D_cache/cache_reg[4][30]  ( .D(\D_cache/n1552 ), .CK(clk), .RN(n5703), .Q(\D_cache/cache[4][30] ), .QN(n1628) );
  DFFRX1 \D_cache/cache_reg[5][30]  ( .D(\D_cache/n1551 ), .CK(clk), .RN(n5703), .Q(\D_cache/cache[5][30] ), .QN(n3204) );
  DFFRX1 \D_cache/cache_reg[6][30]  ( .D(\D_cache/n1550 ), .CK(clk), .RN(n5703), .Q(\D_cache/cache[6][30] ), .QN(n716) );
  DFFRX1 \D_cache/cache_reg[7][30]  ( .D(\D_cache/n1549 ), .CK(clk), .RN(n5703), .Q(\D_cache/cache[7][30] ), .QN(n2284) );
  DFFRX1 \D_cache/cache_reg[1][31]  ( .D(\D_cache/n1547 ), .CK(clk), .RN(n5703), .Q(\D_cache/cache[1][31] ), .QN(n1207) );
  DFFRX1 \D_cache/cache_reg[2][31]  ( .D(\D_cache/n1546 ), .CK(clk), .RN(n5703), .Q(\D_cache/cache[2][31] ), .QN(n682) );
  DFFRX1 \D_cache/cache_reg[3][31]  ( .D(\D_cache/n1545 ), .CK(clk), .RN(n5703), .Q(\D_cache/cache[3][31] ), .QN(n2254) );
  DFFRX1 \D_cache/cache_reg[4][31]  ( .D(\D_cache/n1544 ), .CK(clk), .RN(n5703), .Q(\D_cache/cache[4][31] ), .QN(n1631) );
  DFFRX1 \D_cache/cache_reg[5][31]  ( .D(\D_cache/n1543 ), .CK(clk), .RN(n5702), .Q(\D_cache/cache[5][31] ), .QN(n3207) );
  DFFRX1 \D_cache/cache_reg[6][31]  ( .D(\D_cache/n1542 ), .CK(clk), .RN(n5702), .Q(\D_cache/cache[6][31] ), .QN(n720) );
  DFFRX1 \D_cache/cache_reg[7][31]  ( .D(\D_cache/n1541 ), .CK(clk), .RN(n5702), .Q(\D_cache/cache[7][31] ), .QN(n2288) );
  DFFRX1 \D_cache/cache_reg[1][32]  ( .D(\D_cache/n1539 ), .CK(clk), .RN(n5702), .Q(\D_cache/cache[1][32] ), .QN(n1191) );
  DFFRX1 \D_cache/cache_reg[2][32]  ( .D(\D_cache/n1538 ), .CK(clk), .RN(n5702), .Q(\D_cache/cache[2][32] ), .QN(n690) );
  DFFRX1 \D_cache/cache_reg[3][32]  ( .D(\D_cache/n1537 ), .CK(clk), .RN(n5702), .Q(\D_cache/cache[3][32] ), .QN(n2259) );
  DFFRX1 \D_cache/cache_reg[4][32]  ( .D(\D_cache/n1536 ), .CK(clk), .RN(n5702), .Q(\D_cache/cache[4][32] ), .QN(n2084) );
  DFFRX1 \D_cache/cache_reg[5][32]  ( .D(\D_cache/n1535 ), .CK(clk), .RN(n5702), .Q(\D_cache/cache[5][32] ), .QN(n496) );
  DFFRX1 \D_cache/cache_reg[6][32]  ( .D(\D_cache/n1534 ), .CK(clk), .RN(n5702), .Q(\D_cache/cache[6][32] ), .QN(n2085) );
  DFFRX1 \D_cache/cache_reg[7][32]  ( .D(\D_cache/n1533 ), .CK(clk), .RN(n5702), .Q(\D_cache/cache[7][32] ), .QN(n497) );
  DFFRX1 \D_cache/cache_reg[0][33]  ( .D(\D_cache/n1532 ), .CK(clk), .RN(n5702), .Q(\D_cache/cache[0][33] ), .QN(n1320) );
  DFFRX1 \D_cache/cache_reg[1][33]  ( .D(\D_cache/n1531 ), .CK(clk), .RN(n5701), .Q(\D_cache/cache[1][33] ), .QN(n2849) );
  DFFRX1 \D_cache/cache_reg[2][33]  ( .D(\D_cache/n1530 ), .CK(clk), .RN(n5701), .Q(\D_cache/cache[2][33] ), .QN(n2118) );
  DFFRX1 \D_cache/cache_reg[3][33]  ( .D(\D_cache/n1529 ), .CK(clk), .RN(n5701), .Q(\D_cache/cache[3][33] ), .QN(n531) );
  DFFRX1 \D_cache/cache_reg[4][33]  ( .D(\D_cache/n1528 ), .CK(clk), .RN(n5701), .Q(\D_cache/cache[4][33] ), .QN(n1373) );
  DFFRX1 \D_cache/cache_reg[5][33]  ( .D(\D_cache/n1527 ), .CK(clk), .RN(n5701), .Q(\D_cache/cache[5][33] ), .QN(n2903) );
  DFFRX1 \D_cache/cache_reg[6][33]  ( .D(\D_cache/n1526 ), .CK(clk), .RN(n5701), .Q(\D_cache/cache[6][33] ), .QN(n1319) );
  DFFRX1 \D_cache/cache_reg[7][33]  ( .D(\D_cache/n1525 ), .CK(clk), .RN(n5701), .Q(\D_cache/cache[7][33] ), .QN(n2848) );
  DFFRX1 \D_cache/cache_reg[0][34]  ( .D(\D_cache/n1524 ), .CK(clk), .RN(n5701), .Q(\D_cache/cache[0][34] ), .QN(n779) );
  DFFRX1 \D_cache/cache_reg[1][34]  ( .D(\D_cache/n1523 ), .CK(clk), .RN(n5701), .Q(\D_cache/cache[1][34] ), .QN(n2341) );
  DFFRX1 \D_cache/cache_reg[2][34]  ( .D(\D_cache/n1522 ), .CK(clk), .RN(n5701), .Q(\D_cache/cache[2][34] ), .QN(n781) );
  DFFRX1 \D_cache/cache_reg[3][34]  ( .D(\D_cache/n1521 ), .CK(clk), .RN(n5701), .Q(\D_cache/cache[3][34] ), .QN(n2343) );
  DFFRX1 \D_cache/cache_reg[4][34]  ( .D(\D_cache/n1520 ), .CK(clk), .RN(n5700), .Q(\D_cache/cache[4][34] ), .QN(n782) );
  DFFRX1 \D_cache/cache_reg[5][34]  ( .D(\D_cache/n1519 ), .CK(clk), .RN(n5700), .Q(\D_cache/cache[5][34] ), .QN(n2344) );
  DFFRX1 \D_cache/cache_reg[6][34]  ( .D(\D_cache/n1518 ), .CK(clk), .RN(n5700), .Q(\D_cache/cache[6][34] ), .QN(n780) );
  DFFRX1 \D_cache/cache_reg[7][34]  ( .D(\D_cache/n1517 ), .CK(clk), .RN(n5700), .Q(\D_cache/cache[7][34] ), .QN(n2342) );
  DFFRX1 \D_cache/cache_reg[0][35]  ( .D(\D_cache/n1516 ), .CK(clk), .RN(n5700), .Q(\D_cache/cache[0][35] ), .QN(n1327) );
  DFFRX1 \D_cache/cache_reg[1][35]  ( .D(\D_cache/n1515 ), .CK(clk), .RN(n5700), .Q(\D_cache/cache[1][35] ), .QN(n2856) );
  DFFRX1 \D_cache/cache_reg[2][35]  ( .D(\D_cache/n1514 ), .CK(clk), .RN(n5700), .Q(\D_cache/cache[2][35] ), .QN(n1326) );
  DFFRX1 \D_cache/cache_reg[3][35]  ( .D(\D_cache/n1513 ), .CK(clk), .RN(n5700), .Q(\D_cache/cache[3][35] ), .QN(n2855) );
  DFFRX1 \D_cache/cache_reg[4][35]  ( .D(\D_cache/n1512 ), .CK(clk), .RN(n5700), .Q(\D_cache/cache[4][35] ), .QN(n1370) );
  DFFRX1 \D_cache/cache_reg[5][35]  ( .D(\D_cache/n1511 ), .CK(clk), .RN(n5700), .Q(\D_cache/cache[5][35] ), .QN(n2900) );
  DFFRX1 \D_cache/cache_reg[6][35]  ( .D(\D_cache/n1510 ), .CK(clk), .RN(n5700), .Q(\D_cache/cache[6][35] ), .QN(n1325) );
  DFFRX1 \D_cache/cache_reg[7][35]  ( .D(\D_cache/n1509 ), .CK(clk), .RN(n5700), .Q(\D_cache/cache[7][35] ), .QN(n2854) );
  DFFRX1 \D_cache/cache_reg[0][36]  ( .D(\D_cache/n1508 ), .CK(clk), .RN(n5699), .Q(\D_cache/cache[0][36] ), .QN(n1311) );
  DFFRX1 \D_cache/cache_reg[1][36]  ( .D(\D_cache/n1507 ), .CK(clk), .RN(n5699), .Q(\D_cache/cache[1][36] ), .QN(n2840) );
  DFFRX1 \D_cache/cache_reg[2][36]  ( .D(\D_cache/n1506 ), .CK(clk), .RN(n5699), .Q(\D_cache/cache[2][36] ), .QN(n1310) );
  DFFRX1 \D_cache/cache_reg[3][36]  ( .D(\D_cache/n1505 ), .CK(clk), .RN(n5699), .Q(\D_cache/cache[3][36] ), .QN(n2839) );
  DFFRX1 \D_cache/cache_reg[4][36]  ( .D(\D_cache/n1504 ), .CK(clk), .RN(n5699), .Q(\D_cache/cache[4][36] ), .QN(n1356) );
  DFFRX1 \D_cache/cache_reg[5][36]  ( .D(\D_cache/n1503 ), .CK(clk), .RN(n5699), .Q(\D_cache/cache[5][36] ), .QN(n2886) );
  DFFRX1 \D_cache/cache_reg[6][36]  ( .D(\D_cache/n1502 ), .CK(clk), .RN(n5699), .Q(\D_cache/cache[6][36] ), .QN(n772) );
  DFFRX1 \D_cache/cache_reg[7][36]  ( .D(\D_cache/n1501 ), .CK(clk), .RN(n5699), .Q(\D_cache/cache[7][36] ), .QN(n2334) );
  DFFRX1 \D_cache/cache_reg[0][37]  ( .D(\D_cache/n1500 ), .CK(clk), .RN(n5699), .Q(\D_cache/cache[0][37] ), .QN(n1394) );
  DFFRX1 \D_cache/cache_reg[1][37]  ( .D(\D_cache/n1499 ), .CK(clk), .RN(n5699), .Q(\D_cache/cache[1][37] ), .QN(n2924) );
  DFFRX1 \D_cache/cache_reg[2][37]  ( .D(\D_cache/n1498 ), .CK(clk), .RN(n5699), .Q(\D_cache/cache[2][37] ), .QN(n1248) );
  DFFRX1 \D_cache/cache_reg[3][37]  ( .D(\D_cache/n1497 ), .CK(clk), .RN(n5699), .Q(\D_cache/cache[3][37] ), .QN(n2790) );
  DFFRX1 \D_cache/cache_reg[4][37]  ( .D(\D_cache/n1496 ), .CK(clk), .RN(n5698), .Q(\D_cache/cache[4][37] ), .QN(n1304) );
  DFFRX1 \D_cache/cache_reg[5][37]  ( .D(\D_cache/n1495 ), .CK(clk), .RN(n5698), .Q(\D_cache/cache[5][37] ), .QN(n2833) );
  DFFRX1 \D_cache/cache_reg[6][37]  ( .D(\D_cache/n1494 ), .CK(clk), .RN(n5698), .Q(\D_cache/cache[6][37] ), .QN(n828) );
  DFFRX1 \D_cache/cache_reg[7][37]  ( .D(\D_cache/n1493 ), .CK(clk), .RN(n5698), .Q(\D_cache/cache[7][37] ), .QN(n2391) );
  DFFRX1 \D_cache/cache_reg[0][38]  ( .D(\D_cache/n1492 ), .CK(clk), .RN(n5698), .Q(\D_cache/cache[0][38] ), .QN(n816) );
  DFFRX1 \D_cache/cache_reg[1][38]  ( .D(\D_cache/n1491 ), .CK(clk), .RN(n5698), .Q(\D_cache/cache[1][38] ), .QN(n2379) );
  DFFRX1 \D_cache/cache_reg[2][38]  ( .D(\D_cache/n1490 ), .CK(clk), .RN(n5698), .Q(\D_cache/cache[2][38] ), .QN(n815) );
  DFFRX1 \D_cache/cache_reg[3][38]  ( .D(\D_cache/n1489 ), .CK(clk), .RN(n5698), .Q(\D_cache/cache[3][38] ), .QN(n2378) );
  DFFRX1 \D_cache/cache_reg[4][38]  ( .D(\D_cache/n1488 ), .CK(clk), .RN(n5698), .Q(\D_cache/cache[4][38] ), .QN(n1355) );
  DFFRX1 \D_cache/cache_reg[5][38]  ( .D(\D_cache/n1487 ), .CK(clk), .RN(n5698), .Q(\D_cache/cache[5][38] ), .QN(n2885) );
  DFFRX1 \D_cache/cache_reg[6][38]  ( .D(\D_cache/n1486 ), .CK(clk), .RN(n5698), .Q(\D_cache/cache[6][38] ), .QN(n814) );
  DFFRX1 \D_cache/cache_reg[7][38]  ( .D(\D_cache/n1485 ), .CK(clk), .RN(n5698), .Q(\D_cache/cache[7][38] ), .QN(n2377) );
  DFFRX1 \D_cache/cache_reg[0][39]  ( .D(\D_cache/n1484 ), .CK(clk), .RN(n5697), .Q(\D_cache/cache[0][39] ), .QN(n1334) );
  DFFRX1 \D_cache/cache_reg[1][39]  ( .D(\D_cache/n1483 ), .CK(clk), .RN(n5697), .Q(\D_cache/cache[1][39] ), .QN(n2863) );
  DFFRX1 \D_cache/cache_reg[2][39]  ( .D(\D_cache/n1482 ), .CK(clk), .RN(n5697), .Q(\D_cache/cache[2][39] ), .QN(n1216) );
  DFFRX1 \D_cache/cache_reg[3][39]  ( .D(\D_cache/n1481 ), .CK(clk), .RN(n5697), .Q(\D_cache/cache[3][39] ), .QN(n2753) );
  DFFRX1 \D_cache/cache_reg[4][39]  ( .D(\D_cache/n1480 ), .CK(clk), .RN(n5697), .Q(\D_cache/cache[4][39] ), .QN(n1372) );
  DFFRX1 \D_cache/cache_reg[5][39]  ( .D(\D_cache/n1479 ), .CK(clk), .RN(n5697), .Q(\D_cache/cache[5][39] ), .QN(n2902) );
  DFFRX1 \D_cache/cache_reg[6][39]  ( .D(\D_cache/n1478 ), .CK(clk), .RN(n5697), .Q(\D_cache/cache[6][39] ), .QN(n1333) );
  DFFRX1 \D_cache/cache_reg[7][39]  ( .D(\D_cache/n1477 ), .CK(clk), .RN(n5697), .Q(\D_cache/cache[7][39] ), .QN(n2862) );
  DFFRX1 \D_cache/cache_reg[0][40]  ( .D(\D_cache/n1476 ), .CK(clk), .RN(n5697), .Q(\D_cache/cache[0][40] ), .QN(n2192) );
  DFFRX1 \D_cache/cache_reg[1][40]  ( .D(\D_cache/n1475 ), .CK(clk), .RN(n5697), .Q(\D_cache/cache[1][40] ), .QN(n618) );
  DFFRX1 \D_cache/cache_reg[2][40]  ( .D(\D_cache/n1474 ), .CK(clk), .RN(n5697), .Q(\D_cache/cache[2][40] ), .QN(n2193) );
  DFFRX1 \D_cache/cache_reg[3][40]  ( .D(\D_cache/n1473 ), .CK(clk), .RN(n5697), .Q(\D_cache/cache[3][40] ), .QN(n619) );
  DFFRX1 \D_cache/cache_reg[4][40]  ( .D(\D_cache/n1472 ), .CK(clk), .RN(n5696), .Q(\D_cache/cache[4][40] ), .QN(n3395) );
  DFFRX1 \D_cache/cache_reg[5][40]  ( .D(\D_cache/n1471 ), .CK(clk), .RN(n5701), .Q(\D_cache/cache[5][40] ), .QN(n1766) );
  DFFRX1 \D_cache/cache_reg[6][40]  ( .D(\D_cache/n1470 ), .CK(clk), .RN(n5676), .Q(\D_cache/cache[6][40] ), .QN(n2194) );
  DFFRX1 \D_cache/cache_reg[7][40]  ( .D(\D_cache/n1469 ), .CK(clk), .RN(n5676), .Q(\D_cache/cache[7][40] ), .QN(n620) );
  DFFRX1 \D_cache/cache_reg[0][41]  ( .D(\D_cache/n1468 ), .CK(clk), .RN(n5676), .Q(\D_cache/cache[0][41] ), .QN(n784) );
  DFFRX1 \D_cache/cache_reg[1][41]  ( .D(\D_cache/n1467 ), .CK(clk), .RN(n5676), .Q(\D_cache/cache[1][41] ), .QN(n2346) );
  DFFRX1 \D_cache/cache_reg[2][41]  ( .D(\D_cache/n1466 ), .CK(clk), .RN(n5676), .Q(\D_cache/cache[2][41] ), .QN(n2143) );
  DFFRX1 \D_cache/cache_reg[3][41]  ( .D(\D_cache/n1465 ), .CK(clk), .RN(n5676), .Q(\D_cache/cache[3][41] ), .QN(n563) );
  DFFRX1 \D_cache/cache_reg[4][41]  ( .D(\D_cache/n1464 ), .CK(clk), .RN(n5676), .Q(\D_cache/cache[4][41] ), .QN(n1300) );
  DFFRX1 \D_cache/cache_reg[6][41]  ( .D(\D_cache/n1462 ), .CK(clk), .RN(n5676), .Q(\D_cache/cache[6][41] ), .QN(n2153) );
  DFFRX1 \D_cache/cache_reg[7][41]  ( .D(\D_cache/n1461 ), .CK(clk), .RN(n5676), .Q(\D_cache/cache[7][41] ), .QN(n574) );
  DFFRX1 \D_cache/cache_reg[0][42]  ( .D(\D_cache/n1460 ), .CK(clk), .RN(n5676), .Q(\D_cache/cache[0][42] ), .QN(n759) );
  DFFRX1 \D_cache/cache_reg[1][42]  ( .D(\D_cache/n1459 ), .CK(clk), .RN(n5675), .Q(\D_cache/cache[1][42] ), .QN(n2320) );
  DFFRX1 \D_cache/cache_reg[2][42]  ( .D(\D_cache/n1458 ), .CK(clk), .RN(n5675), .Q(\D_cache/cache[2][42] ), .QN(n1312) );
  DFFRX1 \D_cache/cache_reg[3][42]  ( .D(\D_cache/n1457 ), .CK(clk), .RN(n5675), .Q(\D_cache/cache[3][42] ), .QN(n2841) );
  DFFRX1 \D_cache/cache_reg[4][42]  ( .D(\D_cache/n1456 ), .CK(clk), .RN(n5675), .Q(\D_cache/cache[4][42] ), .QN(n767) );
  DFFRX1 \D_cache/cache_reg[5][42]  ( .D(\D_cache/n1455 ), .CK(clk), .RN(n5675), .Q(\D_cache/cache[5][42] ), .QN(n2329) );
  DFFRX1 \D_cache/cache_reg[6][42]  ( .D(\D_cache/n1454 ), .CK(clk), .RN(n5675), .Q(\D_cache/cache[6][42] ), .QN(n766) );
  DFFRX1 \D_cache/cache_reg[7][42]  ( .D(\D_cache/n1453 ), .CK(clk), .RN(n5675), .Q(\D_cache/cache[7][42] ), .QN(n2328) );
  DFFRX1 \D_cache/cache_reg[0][43]  ( .D(\D_cache/n1452 ), .CK(clk), .RN(n5675), .Q(\D_cache/cache[0][43] ), .QN(n2195) );
  DFFRX1 \D_cache/cache_reg[1][43]  ( .D(\D_cache/n1451 ), .CK(clk), .RN(n5675), .Q(\D_cache/cache[1][43] ), .QN(n621) );
  DFFRX1 \D_cache/cache_reg[2][43]  ( .D(\D_cache/n1450 ), .CK(clk), .RN(n5675), .Q(\D_cache/cache[2][43] ), .QN(n2196) );
  DFFRX1 \D_cache/cache_reg[3][43]  ( .D(\D_cache/n1449 ), .CK(clk), .RN(n5675), .Q(\D_cache/cache[3][43] ), .QN(n622) );
  DFFRX1 \D_cache/cache_reg[4][43]  ( .D(\D_cache/n1448 ), .CK(clk), .RN(n5675), .Q(\D_cache/cache[4][43] ), .QN(n3396) );
  DFFRX1 \D_cache/cache_reg[5][43]  ( .D(\D_cache/n1447 ), .CK(clk), .RN(n5674), .Q(\D_cache/cache[5][43] ), .QN(n1767) );
  DFFRX1 \D_cache/cache_reg[6][43]  ( .D(\D_cache/n1446 ), .CK(clk), .RN(n5674), .Q(\D_cache/cache[6][43] ), .QN(n2197) );
  DFFRX1 \D_cache/cache_reg[7][43]  ( .D(\D_cache/n1445 ), .CK(clk), .RN(n5674), .Q(\D_cache/cache[7][43] ), .QN(n623) );
  DFFRX1 \D_cache/cache_reg[1][44]  ( .D(\D_cache/n1443 ), .CK(clk), .RN(n5674), .Q(\D_cache/cache[1][44] ), .QN(n1185) );
  DFFRX1 \D_cache/cache_reg[2][44]  ( .D(\D_cache/n1442 ), .CK(clk), .RN(n5674), .Q(\D_cache/cache[2][44] ), .QN(n1148) );
  DFFRX1 \D_cache/cache_reg[3][44]  ( .D(\D_cache/n1441 ), .CK(clk), .RN(n5674), .Q(\D_cache/cache[3][44] ), .QN(n2706) );
  DFFRX1 \D_cache/cache_reg[4][44]  ( .D(\D_cache/n1440 ), .CK(clk), .RN(n5674), .Q(\D_cache/cache[4][44] ), .QN(n2677) );
  DFFRX1 \D_cache/cache_reg[5][44]  ( .D(\D_cache/n1439 ), .CK(clk), .RN(n5674), .Q(\D_cache/cache[5][44] ), .QN(n1120) );
  DFFRX1 \D_cache/cache_reg[6][44]  ( .D(\D_cache/n1438 ), .CK(clk), .RN(n5674), .Q(\D_cache/cache[6][44] ), .QN(n695) );
  DFFRX1 \D_cache/cache_reg[7][44]  ( .D(\D_cache/n1437 ), .CK(clk), .RN(n5674), .Q(\D_cache/cache[7][44] ), .QN(n2264) );
  DFFRX1 \D_cache/cache_reg[1][45]  ( .D(\D_cache/n1435 ), .CK(clk), .RN(n5673), .Q(\D_cache/cache[1][45] ), .QN(n1147) );
  DFFRX1 \D_cache/cache_reg[2][45]  ( .D(\D_cache/n1434 ), .CK(clk), .RN(n5673), .Q(\D_cache/cache[2][45] ), .QN(n1297) );
  DFFRX1 \D_cache/cache_reg[3][45]  ( .D(\D_cache/n1433 ), .CK(clk), .RN(n5673), .Q(\D_cache/cache[3][45] ), .QN(n2828) );
  DFFRX1 \D_cache/cache_reg[4][45]  ( .D(\D_cache/n1432 ), .CK(clk), .RN(n5673), .Q(\D_cache/cache[4][45] ), .QN(n2289) );
  DFFRX1 \D_cache/cache_reg[5][45]  ( .D(\D_cache/n1431 ), .CK(clk), .RN(n5673), .Q(\D_cache/cache[5][45] ), .QN(n724) );
  DFFRX1 \D_cache/cache_reg[6][45]  ( .D(\D_cache/n1430 ), .CK(clk), .RN(n5673), .Q(\D_cache/cache[6][45] ), .QN(n2110) );
  DFFRX1 \D_cache/cache_reg[7][45]  ( .D(\D_cache/n1429 ), .CK(clk), .RN(n5673), .Q(\D_cache/cache[7][45] ), .QN(n523) );
  DFFRX1 \D_cache/cache_reg[1][46]  ( .D(\D_cache/n1427 ), .CK(clk), .RN(n5673), .Q(\D_cache/cache[1][46] ), .QN(n1199) );
  DFFRX1 \D_cache/cache_reg[2][46]  ( .D(\D_cache/n1426 ), .CK(clk), .RN(n5673), .Q(\D_cache/cache[2][46] ), .QN(n2093) );
  DFFRX1 \D_cache/cache_reg[3][46]  ( .D(\D_cache/n1425 ), .CK(clk), .RN(n5673), .Q(\D_cache/cache[3][46] ), .QN(n506) );
  DFFRX1 \D_cache/cache_reg[4][46]  ( .D(\D_cache/n1424 ), .CK(clk), .RN(n5673), .Q(\D_cache/cache[4][46] ), .QN(n3355) );
  DFFRX1 \D_cache/cache_reg[5][46]  ( .D(\D_cache/n1423 ), .CK(clk), .RN(n5672), .Q(\D_cache/cache[5][46] ), .QN(n1735) );
  DFFRX1 \D_cache/cache_reg[6][46]  ( .D(\D_cache/n1422 ), .CK(clk), .RN(n5672), .Q(\D_cache/cache[6][46] ), .QN(n2094) );
  DFFRX1 \D_cache/cache_reg[7][46]  ( .D(\D_cache/n1421 ), .CK(clk), .RN(n5672), .Q(\D_cache/cache[7][46] ), .QN(n507) );
  DFFRX1 \D_cache/cache_reg[0][47]  ( .D(\D_cache/n1420 ), .CK(clk), .RN(n5672), .Q(\D_cache/cache[0][47] ), .QN(n689) );
  DFFRX1 \D_cache/cache_reg[1][47]  ( .D(\D_cache/n1419 ), .CK(clk), .RN(n5672), .Q(\D_cache/cache[1][47] ), .QN(n2323) );
  DFFRX1 \D_cache/cache_reg[2][47]  ( .D(\D_cache/n1418 ), .CK(clk), .RN(n5672), .Q(\D_cache/cache[2][47] ), .QN(n2149) );
  DFFRX1 \D_cache/cache_reg[3][47]  ( .D(\D_cache/n1417 ), .CK(clk), .RN(n5672), .Q(\D_cache/cache[3][47] ), .QN(n569) );
  DFFRX1 \D_cache/cache_reg[4][47]  ( .D(\D_cache/n1416 ), .CK(clk), .RN(n5672), .Q(\D_cache/cache[4][47] ), .QN(n2167) );
  DFFRX1 \D_cache/cache_reg[5][47]  ( .D(\D_cache/n1415 ), .CK(clk), .RN(n5672), .Q(\D_cache/cache[5][47] ), .QN(n593) );
  DFFRX1 \D_cache/cache_reg[6][47]  ( .D(\D_cache/n1414 ), .CK(clk), .RN(n5672), .Q(\D_cache/cache[6][47] ), .QN(n2147) );
  DFFRX1 \D_cache/cache_reg[7][47]  ( .D(\D_cache/n1413 ), .CK(clk), .RN(n5672), .Q(\D_cache/cache[7][47] ), .QN(n567) );
  DFFRX1 \D_cache/cache_reg[1][48]  ( .D(\D_cache/n1411 ), .CK(clk), .RN(n5671), .Q(\D_cache/cache[1][48] ), .QN(n1193) );
  DFFRX1 \D_cache/cache_reg[2][48]  ( .D(\D_cache/n1410 ), .CK(clk), .RN(n5671), .Q(\D_cache/cache[2][48] ), .QN(n691) );
  DFFRX1 \D_cache/cache_reg[3][48]  ( .D(\D_cache/n1409 ), .CK(clk), .RN(n5671), .Q(\D_cache/cache[3][48] ), .QN(n2260) );
  DFFRX1 \D_cache/cache_reg[4][48]  ( .D(\D_cache/n1408 ), .CK(clk), .RN(n5671), .Q(\D_cache/cache[4][48] ), .QN(n1146) );
  DFFRX1 \D_cache/cache_reg[5][48]  ( .D(\D_cache/n1407 ), .CK(clk), .RN(n5671), .Q(\D_cache/cache[5][48] ), .QN(n2705) );
  DFFRX1 \D_cache/cache_reg[6][48]  ( .D(\D_cache/n1406 ), .CK(clk), .RN(n5671), .Q(\D_cache/cache[6][48] ), .QN(n2087) );
  DFFRX1 \D_cache/cache_reg[7][48]  ( .D(\D_cache/n1405 ), .CK(clk), .RN(n5671), .Q(\D_cache/cache[7][48] ), .QN(n499) );
  DFFRX1 \D_cache/cache_reg[1][49]  ( .D(\D_cache/n1403 ), .CK(clk), .RN(n5671), .Q(\D_cache/cache[1][49] ), .QN(n1285) );
  DFFRX1 \D_cache/cache_reg[2][49]  ( .D(\D_cache/n1402 ), .CK(clk), .RN(n5671), .Q(\D_cache/cache[2][49] ), .QN(n737) );
  DFFRX1 \D_cache/cache_reg[3][49]  ( .D(\D_cache/n1401 ), .CK(clk), .RN(n5671), .Q(\D_cache/cache[3][49] ), .QN(n2296) );
  DFFRX1 \D_cache/cache_reg[4][49]  ( .D(\D_cache/n1400 ), .CK(clk), .RN(n5670), .Q(\D_cache/cache[4][49] ), .QN(n1454) );
  DFFRX1 \D_cache/cache_reg[5][49]  ( .D(\D_cache/n1399 ), .CK(clk), .RN(n5670), .Q(\D_cache/cache[5][49] ), .QN(n3025) );
  DFFRX1 \D_cache/cache_reg[6][49]  ( .D(\D_cache/n1398 ), .CK(clk), .RN(n5670), .Q(\D_cache/cache[6][49] ), .QN(n2099) );
  DFFRX1 \D_cache/cache_reg[7][49]  ( .D(\D_cache/n1397 ), .CK(clk), .RN(n5670), .Q(\D_cache/cache[7][49] ), .QN(n514) );
  DFFRX1 \D_cache/cache_reg[1][50]  ( .D(\D_cache/n1395 ), .CK(clk), .RN(n5670), .Q(\D_cache/cache[1][50] ), .QN(n1190) );
  DFFRX1 \D_cache/cache_reg[2][50]  ( .D(\D_cache/n1394 ), .CK(clk), .RN(n5670), .Q(\D_cache/cache[2][50] ), .QN(n1151) );
  DFFRX1 \D_cache/cache_reg[3][50]  ( .D(\D_cache/n1393 ), .CK(clk), .RN(n5670), .Q(\D_cache/cache[3][50] ), .QN(n2708) );
  DFFRX1 \D_cache/cache_reg[4][50]  ( .D(\D_cache/n1392 ), .CK(clk), .RN(n5670), .Q(\D_cache/cache[4][50] ), .QN(n2091) );
  DFFRX1 \D_cache/cache_reg[5][50]  ( .D(\D_cache/n1391 ), .CK(clk), .RN(n5670), .Q(\D_cache/cache[5][50] ), .QN(n504) );
  DFFRX1 \D_cache/cache_reg[6][50]  ( .D(\D_cache/n1390 ), .CK(clk), .RN(n5670), .Q(\D_cache/cache[6][50] ), .QN(n678) );
  DFFRX1 \D_cache/cache_reg[7][50]  ( .D(\D_cache/n1389 ), .CK(clk), .RN(n5670), .Q(\D_cache/cache[7][50] ), .QN(n2249) );
  DFFRX1 \D_cache/cache_reg[2][51]  ( .D(\D_cache/n1386 ), .CK(clk), .RN(n5669), .Q(\D_cache/cache[2][51] ), .QN(n1110) );
  DFFRX1 \D_cache/cache_reg[3][51]  ( .D(\D_cache/n1385 ), .CK(clk), .RN(n5669), .Q(\D_cache/cache[3][51] ), .QN(n2699) );
  DFFRX1 \D_cache/cache_reg[4][51]  ( .D(\D_cache/n1384 ), .CK(clk), .RN(n5669), .Q(\D_cache/cache[4][51] ), .QN(n1161) );
  DFFRX1 \D_cache/cache_reg[5][51]  ( .D(\D_cache/n1383 ), .CK(clk), .RN(n5669), .Q(\D_cache/cache[5][51] ), .QN(n2717) );
  DFFRX1 \D_cache/cache_reg[6][51]  ( .D(\D_cache/n1382 ), .CK(clk), .RN(n5669), .Q(\D_cache/cache[6][51] ), .QN(n2080) );
  DFFRX1 \D_cache/cache_reg[7][51]  ( .D(\D_cache/n1381 ), .CK(clk), .RN(n5669), .Q(\D_cache/cache[7][51] ), .QN(n492) );
  DFFRX1 \D_cache/cache_reg[0][52]  ( .D(\D_cache/n1380 ), .CK(clk), .RN(n5669), .Q(\D_cache/cache[0][52] ), .QN(n1352) );
  DFFRX1 \D_cache/cache_reg[1][52]  ( .D(\D_cache/n1379 ), .CK(clk), .RN(n5669), .Q(\D_cache/cache[1][52] ), .QN(n2882) );
  DFFRX1 \D_cache/cache_reg[2][52]  ( .D(\D_cache/n1378 ), .CK(clk), .RN(n5669), .Q(\D_cache/cache[2][52] ), .QN(n2200) );
  DFFRX1 \D_cache/cache_reg[3][52]  ( .D(\D_cache/n1377 ), .CK(clk), .RN(n5669), .Q(\D_cache/cache[3][52] ), .QN(n626) );
  DFFRX1 \D_cache/cache_reg[4][52]  ( .D(\D_cache/n1376 ), .CK(clk), .RN(n5668), .Q(\D_cache/cache[4][52] ), .QN(n3399) );
  DFFRX1 \D_cache/cache_reg[5][52]  ( .D(\D_cache/n1375 ), .CK(clk), .RN(n5668), .Q(\D_cache/cache[5][52] ), .QN(n1770) );
  DFFRX1 \D_cache/cache_reg[6][52]  ( .D(\D_cache/n1374 ), .CK(clk), .RN(n5668), .Q(\D_cache/cache[6][52] ), .QN(n2201) );
  DFFRX1 \D_cache/cache_reg[7][52]  ( .D(\D_cache/n1373 ), .CK(clk), .RN(n5668), .Q(\D_cache/cache[7][52] ), .QN(n627) );
  DFFRX1 \D_cache/cache_reg[0][53]  ( .D(\D_cache/n1372 ), .CK(clk), .RN(n5668), .Q(\D_cache/cache[0][53] ), .QN(n746) );
  DFFRX1 \D_cache/cache_reg[1][53]  ( .D(\D_cache/n1371 ), .CK(clk), .RN(n5668), .Q(\D_cache/cache[1][53] ), .QN(n2307) );
  DFFRX1 \D_cache/cache_reg[2][53]  ( .D(\D_cache/n1370 ), .CK(clk), .RN(n5668), .Q(\D_cache/cache[2][53] ), .QN(n2140) );
  DFFRX1 \D_cache/cache_reg[3][53]  ( .D(\D_cache/n1369 ), .CK(clk), .RN(n5668), .Q(\D_cache/cache[3][53] ), .QN(n560) );
  DFFRX1 \D_cache/cache_reg[4][53]  ( .D(\D_cache/n1368 ), .CK(clk), .RN(n5668), .Q(\D_cache/cache[4][53] ), .QN(n745) );
  DFFRX1 \D_cache/cache_reg[5][53]  ( .D(\D_cache/n1367 ), .CK(clk), .RN(n5668), .Q(\D_cache/cache[5][53] ), .QN(n2306) );
  DFFRX1 \D_cache/cache_reg[6][53]  ( .D(\D_cache/n1366 ), .CK(clk), .RN(n5668), .Q(\D_cache/cache[6][53] ), .QN(n773) );
  DFFRX1 \D_cache/cache_reg[7][53]  ( .D(\D_cache/n1365 ), .CK(clk), .RN(n5668), .Q(\D_cache/cache[7][53] ), .QN(n2335) );
  DFFRX1 \D_cache/cache_reg[0][54]  ( .D(\D_cache/n1364 ), .CK(clk), .RN(n5667), .Q(\D_cache/cache[0][54] ), .QN(n648) );
  DFFRX1 \D_cache/cache_reg[1][54]  ( .D(\D_cache/n1363 ), .CK(clk), .RN(n5667), .Q(\D_cache/cache[1][54] ), .QN(n2225) );
  DFFRX1 \D_cache/cache_reg[2][54]  ( .D(\D_cache/n1362 ), .CK(clk), .RN(n5667), .Q(\D_cache/cache[2][54] ), .QN(n2114) );
  DFFRX1 \D_cache/cache_reg[3][54]  ( .D(\D_cache/n1361 ), .CK(clk), .RN(n5667), .Q(\D_cache/cache[3][54] ), .QN(n527) );
  DFFRX1 \D_cache/cache_reg[4][54]  ( .D(\D_cache/n1360 ), .CK(clk), .RN(n5667), .Q(\D_cache/cache[4][54] ), .QN(n1302) );
  DFFRX1 \D_cache/cache_reg[5][54]  ( .D(\D_cache/n1359 ), .CK(clk), .RN(n5667), .Q(\D_cache/cache[5][54] ), .QN(n2832) );
  DFFRX1 \D_cache/cache_reg[6][54]  ( .D(\D_cache/n1358 ), .CK(clk), .RN(n5667), .Q(\D_cache/cache[6][54] ), .QN(n2100) );
  DFFRX1 \D_cache/cache_reg[7][54]  ( .D(\D_cache/n1357 ), .CK(clk), .RN(n5667), .Q(\D_cache/cache[7][54] ), .QN(n515) );
  DFFRX1 \D_cache/cache_reg[1][55]  ( .D(\D_cache/n1355 ), .CK(clk), .RN(n5667), .Q(\D_cache/cache[1][55] ), .QN(n1200) );
  DFFRX1 \D_cache/cache_reg[2][55]  ( .D(\D_cache/n1354 ), .CK(clk), .RN(n5667), .Q(\D_cache/cache[2][55] ), .QN(n2095) );
  DFFRX1 \D_cache/cache_reg[3][55]  ( .D(\D_cache/n1353 ), .CK(clk), .RN(n5667), .Q(\D_cache/cache[3][55] ), .QN(n508) );
  DFFRX1 \D_cache/cache_reg[4][55]  ( .D(\D_cache/n1352 ), .CK(clk), .RN(n5671), .Q(\D_cache/cache[4][55] ), .QN(n3356) );
  DFFRX1 \D_cache/cache_reg[5][55]  ( .D(\D_cache/n1351 ), .CK(clk), .RN(n5686), .Q(\D_cache/cache[5][55] ), .QN(n1736) );
  DFFRX1 \D_cache/cache_reg[6][55]  ( .D(\D_cache/n1350 ), .CK(clk), .RN(n5686), .Q(\D_cache/cache[6][55] ), .QN(n2096) );
  DFFRX1 \D_cache/cache_reg[7][55]  ( .D(\D_cache/n1349 ), .CK(clk), .RN(n5686), .Q(\D_cache/cache[7][55] ), .QN(n509) );
  DFFRX1 \D_cache/cache_reg[0][56]  ( .D(\D_cache/n1348 ), .CK(clk), .RN(n5686), .Q(\D_cache/cache[0][56] ), .QN(n817) );
  DFFRX1 \D_cache/cache_reg[1][56]  ( .D(\D_cache/n1347 ), .CK(clk), .RN(n5686), .Q(\D_cache/cache[1][56] ), .QN(n2380) );
  DFFRX1 \D_cache/cache_reg[2][56]  ( .D(\D_cache/n1346 ), .CK(clk), .RN(n5686), .Q(\D_cache/cache[2][56] ), .QN(n1313) );
  DFFRX1 \D_cache/cache_reg[3][56]  ( .D(\D_cache/n1345 ), .CK(clk), .RN(n5686), .Q(\D_cache/cache[3][56] ), .QN(n2842) );
  DFFRX1 \D_cache/cache_reg[4][56]  ( .D(\D_cache/n1344 ), .CK(clk), .RN(n5686), .Q(\D_cache/cache[4][56] ), .QN(n761) );
  DFFRX1 \D_cache/cache_reg[5][56]  ( .D(\D_cache/n1343 ), .CK(clk), .RN(n5686), .Q(\D_cache/cache[5][56] ), .QN(n2322) );
  DFFRX1 \D_cache/cache_reg[6][56]  ( .D(\D_cache/n1342 ), .CK(clk), .RN(n5686), .Q(\D_cache/cache[6][56] ), .QN(n2136) );
  DFFRX1 \D_cache/cache_reg[7][56]  ( .D(\D_cache/n1341 ), .CK(clk), .RN(n5685), .Q(\D_cache/cache[7][56] ), .QN(n551) );
  DFFRX1 \D_cache/cache_reg[1][57]  ( .D(\D_cache/n1339 ), .CK(clk), .RN(n5685), .Q(\D_cache/cache[1][57] ), .QN(n729) );
  DFFRX1 \D_cache/cache_reg[2][57]  ( .D(\D_cache/n1338 ), .CK(clk), .RN(n5685), .Q(\D_cache/cache[2][57] ), .QN(n709) );
  DFFRX1 \D_cache/cache_reg[3][57]  ( .D(\D_cache/n1337 ), .CK(clk), .RN(n5685), .Q(\D_cache/cache[3][57] ), .QN(n2277) );
  DFFRX1 \D_cache/cache_reg[4][57]  ( .D(\D_cache/n1336 ), .CK(clk), .RN(n5685), .Q(\D_cache/cache[4][57] ), .QN(n693) );
  DFFRX1 \D_cache/cache_reg[5][57]  ( .D(\D_cache/n1335 ), .CK(clk), .RN(n5685), .Q(\D_cache/cache[5][57] ), .QN(n2262) );
  DFFRX1 \D_cache/cache_reg[6][57]  ( .D(\D_cache/n1334 ), .CK(clk), .RN(n5685), .Q(\D_cache/cache[6][57] ), .QN(n708) );
  DFFRX1 \D_cache/cache_reg[7][57]  ( .D(\D_cache/n1333 ), .CK(clk), .RN(n5685), .Q(\D_cache/cache[7][57] ), .QN(n2276) );
  DFFRX1 \D_cache/cache_reg[1][58]  ( .D(\D_cache/n1331 ), .CK(clk), .RN(n5685), .Q(\D_cache/cache[1][58] ), .QN(n1197) );
  DFFRX1 \D_cache/cache_reg[2][58]  ( .D(\D_cache/n1330 ), .CK(clk), .RN(n5685), .Q(\D_cache/cache[2][58] ), .QN(n692) );
  DFFRX1 \D_cache/cache_reg[3][58]  ( .D(\D_cache/n1329 ), .CK(clk), .RN(n5684), .Q(\D_cache/cache[3][58] ), .QN(n2261) );
  DFFRX1 \D_cache/cache_reg[4][58]  ( .D(\D_cache/n1328 ), .CK(clk), .RN(n5684), .Q(\D_cache/cache[4][58] ), .QN(n1452) );
  DFFRX1 \D_cache/cache_reg[5][58]  ( .D(\D_cache/n1327 ), .CK(clk), .RN(n5684), .Q(\D_cache/cache[5][58] ), .QN(n3022) );
  DFFRX1 \D_cache/cache_reg[6][58]  ( .D(\D_cache/n1326 ), .CK(clk), .RN(n5684), .Q(\D_cache/cache[6][58] ), .QN(n2097) );
  DFFRX1 \D_cache/cache_reg[7][58]  ( .D(\D_cache/n1325 ), .CK(clk), .RN(n5684), .Q(\D_cache/cache[7][58] ), .QN(n510) );
  DFFRX1 \D_cache/cache_reg[1][59]  ( .D(\D_cache/n1323 ), .CK(clk), .RN(n5684), .Q(\D_cache/cache[1][59] ), .QN(n733) );
  DFFRX1 \D_cache/cache_reg[2][59]  ( .D(\D_cache/n1322 ), .CK(clk), .RN(n5684), .Q(\D_cache/cache[2][59] ), .QN(n715) );
  DFFRX1 \D_cache/cache_reg[3][59]  ( .D(\D_cache/n1321 ), .CK(clk), .RN(n5684), .Q(\D_cache/cache[3][59] ), .QN(n2283) );
  DFFRX1 \D_cache/cache_reg[4][59]  ( .D(\D_cache/n1320 ), .CK(clk), .RN(n5684), .Q(\D_cache/cache[4][59] ), .QN(n1085) );
  DFFRX1 \D_cache/cache_reg[5][59]  ( .D(\D_cache/n1319 ), .CK(clk), .RN(n5684), .Q(\D_cache/cache[5][59] ), .QN(n2679) );
  DFFRX1 \D_cache/cache_reg[6][59]  ( .D(\D_cache/n1318 ), .CK(clk), .RN(n5684), .Q(\D_cache/cache[6][59] ), .QN(n2079) );
  DFFRX1 \D_cache/cache_reg[7][59]  ( .D(\D_cache/n1317 ), .CK(clk), .RN(n5683), .Q(\D_cache/cache[7][59] ), .QN(n491) );
  DFFRX1 \D_cache/cache_reg[0][60]  ( .D(\D_cache/n1316 ), .CK(clk), .RN(n5683), .Q(\D_cache/cache[0][60] ), .QN(n2162) );
  DFFRX1 \D_cache/cache_reg[1][60]  ( .D(\D_cache/n1315 ), .CK(clk), .RN(n5683), .Q(\D_cache/cache[1][60] ), .QN(n586) );
  DFFRX1 \D_cache/cache_reg[2][60]  ( .D(\D_cache/n1314 ), .CK(clk), .RN(n5683), .Q(\D_cache/cache[2][60] ), .QN(n1301) );
  DFFRX1 \D_cache/cache_reg[3][60]  ( .D(\D_cache/n1313 ), .CK(clk), .RN(n5683), .Q(\D_cache/cache[3][60] ), .QN(n2831) );
  DFFRX1 \D_cache/cache_reg[4][60]  ( .D(\D_cache/n1312 ), .CK(clk), .RN(n5683), .Q(\D_cache/cache[4][60] ), .QN(n1367) );
  DFFRX1 \D_cache/cache_reg[5][60]  ( .D(\D_cache/n1311 ), .CK(clk), .RN(n5683), .Q(\D_cache/cache[5][60] ), .QN(n2897) );
  DFFRX1 \D_cache/cache_reg[6][60]  ( .D(\D_cache/n1310 ), .CK(clk), .RN(n5683), .Q(\D_cache/cache[6][60] ), .QN(n2142) );
  DFFRX1 \D_cache/cache_reg[7][60]  ( .D(\D_cache/n1309 ), .CK(clk), .RN(n5683), .Q(\D_cache/cache[7][60] ), .QN(n562) );
  DFFRX1 \D_cache/cache_reg[0][61]  ( .D(\D_cache/n1308 ), .CK(clk), .RN(n5683), .Q(\D_cache/cache[0][61] ), .QN(n1215) );
  DFFRX1 \D_cache/cache_reg[1][61]  ( .D(\D_cache/n1307 ), .CK(clk), .RN(n5683), .Q(\D_cache/cache[1][61] ), .QN(n2752) );
  DFFRX1 \D_cache/cache_reg[2][61]  ( .D(\D_cache/n1306 ), .CK(clk), .RN(n5683), .Q(\D_cache/cache[2][61] ), .QN(n2198) );
  DFFRX1 \D_cache/cache_reg[3][61]  ( .D(\D_cache/n1305 ), .CK(clk), .RN(n5682), .Q(\D_cache/cache[3][61] ), .QN(n624) );
  DFFRX1 \D_cache/cache_reg[4][61]  ( .D(\D_cache/n1304 ), .CK(clk), .RN(n5682), .Q(\D_cache/cache[4][61] ), .QN(n3397) );
  DFFRX1 \D_cache/cache_reg[5][61]  ( .D(\D_cache/n1303 ), .CK(clk), .RN(n5682), .Q(\D_cache/cache[5][61] ), .QN(n1768) );
  DFFRX1 \D_cache/cache_reg[6][61]  ( .D(\D_cache/n1302 ), .CK(clk), .RN(n5682), .Q(\D_cache/cache[6][61] ), .QN(n2072) );
  DFFRX1 \D_cache/cache_reg[7][61]  ( .D(\D_cache/n1301 ), .CK(clk), .RN(n5682), .Q(\D_cache/cache[7][61] ), .QN(n481) );
  DFFRX1 \D_cache/cache_reg[1][62]  ( .D(\D_cache/n1299 ), .CK(clk), .RN(n5682), .Q(\D_cache/cache[1][62] ), .QN(n1206) );
  DFFRX1 \D_cache/cache_reg[2][62]  ( .D(\D_cache/n1298 ), .CK(clk), .RN(n5682), .Q(\D_cache/cache[2][62] ), .QN(n1179) );
  DFFRX1 \D_cache/cache_reg[3][62]  ( .D(\D_cache/n1297 ), .CK(clk), .RN(n5682), .Q(\D_cache/cache[3][62] ), .QN(n2728) );
  DFFRX1 \D_cache/cache_reg[4][62]  ( .D(\D_cache/n1296 ), .CK(clk), .RN(n5682), .Q(\D_cache/cache[4][62] ), .QN(n1574) );
  DFFRX1 \D_cache/cache_reg[5][62]  ( .D(\D_cache/n1295 ), .CK(clk), .RN(n5682), .Q(\D_cache/cache[5][62] ), .QN(n3156) );
  DFFRX1 \D_cache/cache_reg[6][62]  ( .D(\D_cache/n1294 ), .CK(clk), .RN(n5682), .Q(\D_cache/cache[6][62] ), .QN(n2082) );
  DFFRX1 \D_cache/cache_reg[7][62]  ( .D(\D_cache/n1293 ), .CK(clk), .RN(n5681), .Q(\D_cache/cache[7][62] ), .QN(n494) );
  DFFRX1 \D_cache/cache_reg[1][63]  ( .D(\D_cache/n1291 ), .CK(clk), .RN(n5681), .Q(\D_cache/cache[1][63] ), .QN(n1205) );
  DFFRX1 \D_cache/cache_reg[2][63]  ( .D(\D_cache/n1290 ), .CK(clk), .RN(n5681), .Q(\D_cache/cache[2][63] ), .QN(n711) );
  DFFRX1 \D_cache/cache_reg[3][63]  ( .D(\D_cache/n1289 ), .CK(clk), .RN(n5681), .Q(\D_cache/cache[3][63] ), .QN(n2279) );
  DFFRX1 \D_cache/cache_reg[4][63]  ( .D(\D_cache/n1288 ), .CK(clk), .RN(n5681), .Q(\D_cache/cache[4][63] ), .QN(n1630) );
  DFFRX1 \D_cache/cache_reg[5][63]  ( .D(\D_cache/n1287 ), .CK(clk), .RN(n5681), .Q(\D_cache/cache[5][63] ), .QN(n3206) );
  DFFRX1 \D_cache/cache_reg[6][63]  ( .D(\D_cache/n1286 ), .CK(clk), .RN(n5681), .Q(\D_cache/cache[6][63] ), .QN(n710) );
  DFFRX1 \D_cache/cache_reg[7][63]  ( .D(\D_cache/n1285 ), .CK(clk), .RN(n5681), .Q(\D_cache/cache[7][63] ), .QN(n2278) );
  DFFRX1 \D_cache/cache_reg[1][64]  ( .D(\D_cache/n1283 ), .CK(clk), .RN(n5681), .Q(\D_cache/cache[1][64] ), .QN(n849) );
  DFFRX1 \D_cache/cache_reg[2][64]  ( .D(\D_cache/n1282 ), .CK(clk), .RN(n5680), .Q(\D_cache/cache[2][64] ), .QN(n744) );
  DFFRX1 \D_cache/cache_reg[3][64]  ( .D(\D_cache/n1281 ), .CK(clk), .RN(n5680), .Q(\D_cache/cache[3][64] ), .QN(n2305) );
  DFFRX1 \D_cache/cache_reg[4][64]  ( .D(\D_cache/n1280 ), .CK(clk), .RN(n5680), .Q(\D_cache/cache[4][64] ), .QN(n2730) );
  DFFRX1 \D_cache/cache_reg[5][64]  ( .D(\D_cache/n1279 ), .CK(clk), .RN(n5680), .Q(\D_cache/cache[5][64] ), .QN(n1124) );
  DFFRX1 \D_cache/cache_reg[6][64]  ( .D(\D_cache/n1278 ), .CK(clk), .RN(n5680), .Q(\D_cache/cache[6][64] ), .QN(n654) );
  DFFRX1 \D_cache/cache_reg[7][64]  ( .D(\D_cache/n1277 ), .CK(clk), .RN(n5680), .Q(\D_cache/cache[7][64] ), .QN(n2229) );
  DFFRX1 \D_cache/cache_reg[0][65]  ( .D(\D_cache/n1276 ), .CK(clk), .RN(n5680), .Q(\D_cache/cache[0][65] ), .QN(n805) );
  DFFRX1 \D_cache/cache_reg[1][65]  ( .D(\D_cache/n1275 ), .CK(clk), .RN(n5680), .Q(\D_cache/cache[1][65] ), .QN(n2368) );
  DFFRX1 \D_cache/cache_reg[2][65]  ( .D(\D_cache/n1274 ), .CK(clk), .RN(n5680), .Q(\D_cache/cache[2][65] ), .QN(n2120) );
  DFFRX1 \D_cache/cache_reg[3][65]  ( .D(\D_cache/n1273 ), .CK(clk), .RN(n5680), .Q(\D_cache/cache[3][65] ), .QN(n533) );
  DFFRX1 \D_cache/cache_reg[4][65]  ( .D(\D_cache/n1272 ), .CK(clk), .RN(n5680), .Q(\D_cache/cache[4][65] ), .QN(n783) );
  DFFRX1 \D_cache/cache_reg[5][65]  ( .D(\D_cache/n1271 ), .CK(clk), .RN(n5680), .Q(\D_cache/cache[5][65] ), .QN(n2345) );
  DFFRX1 \D_cache/cache_reg[6][65]  ( .D(\D_cache/n1270 ), .CK(clk), .RN(n5679), .Q(\D_cache/cache[6][65] ), .QN(n804) );
  DFFRX1 \D_cache/cache_reg[7][65]  ( .D(\D_cache/n1269 ), .CK(clk), .RN(n5679), .Q(\D_cache/cache[7][65] ), .QN(n2367) );
  DFFRX1 \D_cache/cache_reg[0][66]  ( .D(\D_cache/n1268 ), .CK(clk), .RN(n5679), .Q(\D_cache/cache[0][66] ), .QN(n1294) );
  DFFRX1 \D_cache/cache_reg[1][66]  ( .D(\D_cache/n1267 ), .CK(clk), .RN(n5679), .Q(\D_cache/cache[1][66] ), .QN(n2825) );
  DFFRX1 \D_cache/cache_reg[2][66]  ( .D(\D_cache/n1266 ), .CK(clk), .RN(n5679), .Q(\D_cache/cache[2][66] ), .QN(n1219) );
  DFFRX1 \D_cache/cache_reg[3][66]  ( .D(\D_cache/n1265 ), .CK(clk), .RN(n5679), .Q(\D_cache/cache[3][66] ), .QN(n2756) );
  DFFRX1 \D_cache/cache_reg[4][66]  ( .D(\D_cache/n1264 ), .CK(clk), .RN(n5679), .Q(\D_cache/cache[4][66] ), .QN(n1295) );
  DFFRX1 \D_cache/cache_reg[5][66]  ( .D(\D_cache/n1263 ), .CK(clk), .RN(n5679), .Q(\D_cache/cache[5][66] ), .QN(n2826) );
  DFFRX1 \D_cache/cache_reg[6][66]  ( .D(\D_cache/n1262 ), .CK(clk), .RN(n5679), .Q(\D_cache/cache[6][66] ), .QN(n774) );
  DFFRX1 \D_cache/cache_reg[7][66]  ( .D(\D_cache/n1261 ), .CK(clk), .RN(n5679), .Q(\D_cache/cache[7][66] ), .QN(n2336) );
  DFFRX1 \D_cache/cache_reg[0][67]  ( .D(\D_cache/n1260 ), .CK(clk), .RN(n5679), .Q(\D_cache/cache[0][67] ), .QN(n813) );
  DFFRX1 \D_cache/cache_reg[1][67]  ( .D(\D_cache/n1259 ), .CK(clk), .RN(n5679), .Q(\D_cache/cache[1][67] ), .QN(n2376) );
  DFFRX1 \D_cache/cache_reg[2][67]  ( .D(\D_cache/n1258 ), .CK(clk), .RN(n5678), .Q(\D_cache/cache[2][67] ), .QN(n812) );
  DFFRX1 \D_cache/cache_reg[3][67]  ( .D(\D_cache/n1257 ), .CK(clk), .RN(n5678), .Q(\D_cache/cache[3][67] ), .QN(n2375) );
  DFFRX1 \D_cache/cache_reg[4][67]  ( .D(\D_cache/n1256 ), .CK(clk), .RN(n5678), .Q(\D_cache/cache[4][67] ), .QN(n752) );
  DFFRX1 \D_cache/cache_reg[5][67]  ( .D(\D_cache/n1255 ), .CK(clk), .RN(n5678), .Q(\D_cache/cache[5][67] ), .QN(n2313) );
  DFFRX1 \D_cache/cache_reg[6][67]  ( .D(\D_cache/n1254 ), .CK(clk), .RN(n5678), .Q(\D_cache/cache[6][67] ), .QN(n811) );
  DFFRX1 \D_cache/cache_reg[7][67]  ( .D(\D_cache/n1253 ), .CK(clk), .RN(n5678), .Q(\D_cache/cache[7][67] ), .QN(n2374) );
  DFFRX1 \D_cache/cache_reg[0][68]  ( .D(\D_cache/n1252 ), .CK(clk), .RN(n5678), .Q(\D_cache/cache[0][68] ), .QN(n1306) );
  DFFRX1 \D_cache/cache_reg[1][68]  ( .D(\D_cache/n1251 ), .CK(clk), .RN(n5678), .Q(\D_cache/cache[1][68] ), .QN(n2835) );
  DFFRX1 \D_cache/cache_reg[2][68]  ( .D(\D_cache/n1250 ), .CK(clk), .RN(n5678), .Q(\D_cache/cache[2][68] ), .QN(n2148) );
  DFFRX1 \D_cache/cache_reg[3][68]  ( .D(\D_cache/n1249 ), .CK(clk), .RN(n5678), .Q(\D_cache/cache[3][68] ), .QN(n568) );
  DFFRX1 \D_cache/cache_reg[4][68]  ( .D(\D_cache/n1248 ), .CK(clk), .RN(n5678), .Q(\D_cache/cache[4][68] ), .QN(n1354) );
  DFFRX1 \D_cache/cache_reg[5][68]  ( .D(\D_cache/n1247 ), .CK(clk), .RN(n5678), .Q(\D_cache/cache[5][68] ), .QN(n2884) );
  DFFRX1 \D_cache/cache_reg[6][68]  ( .D(\D_cache/n1246 ), .CK(clk), .RN(n5677), .Q(\D_cache/cache[6][68] ), .QN(n1229) );
  DFFRX1 \D_cache/cache_reg[7][68]  ( .D(\D_cache/n1245 ), .CK(clk), .RN(n5677), .Q(\D_cache/cache[7][68] ), .QN(n2766) );
  DFFRX1 \D_cache/cache_reg[1][69]  ( .D(\D_cache/n1243 ), .CK(clk), .RN(n5677), .Q(\D_cache/cache[1][69] ), .QN(n731) );
  DFFRX1 \D_cache/cache_reg[2][69]  ( .D(\D_cache/n1242 ), .CK(clk), .RN(n5677), .Q(\D_cache/cache[2][69] ), .QN(n700) );
  DFFRX1 \D_cache/cache_reg[3][69]  ( .D(\D_cache/n1241 ), .CK(clk), .RN(n5677), .Q(\D_cache/cache[3][69] ), .QN(n2269) );
  DFFRX1 \D_cache/cache_reg[4][69]  ( .D(\D_cache/n1240 ), .CK(clk), .RN(n5677), .Q(\D_cache/cache[4][69] ), .QN(n2083) );
  DFFRX1 \D_cache/cache_reg[5][69]  ( .D(\D_cache/n1239 ), .CK(clk), .RN(n5677), .Q(\D_cache/cache[5][69] ), .QN(n495) );
  DFFRX1 \D_cache/cache_reg[6][69]  ( .D(\D_cache/n1238 ), .CK(clk), .RN(n5677), .Q(\D_cache/cache[6][69] ), .QN(n713) );
  DFFRX1 \D_cache/cache_reg[7][69]  ( .D(\D_cache/n1237 ), .CK(clk), .RN(n5677), .Q(\D_cache/cache[7][69] ), .QN(n2281) );
  DFFRX1 \D_cache/cache_reg[0][70]  ( .D(\D_cache/n1236 ), .CK(clk), .RN(n5677), .Q(\D_cache/cache[0][70] ), .QN(n2292) );
  DFFRX1 \D_cache/cache_reg[1][70]  ( .D(\D_cache/n1235 ), .CK(clk), .RN(n5677), .Q(\D_cache/cache[1][70] ), .QN(n675) );
  DFFRX1 \D_cache/cache_reg[2][70]  ( .D(\D_cache/n1234 ), .CK(clk), .RN(n5676), .Q(\D_cache/cache[2][70] ), .QN(n668) );
  DFFRX1 \D_cache/cache_reg[3][70]  ( .D(\D_cache/n1233 ), .CK(clk), .RN(n5681), .Q(\D_cache/cache[3][70] ), .QN(n2239) );
  DFFRX1 \D_cache/cache_reg[4][70]  ( .D(\D_cache/n1232 ), .CK(clk), .RN(n5686), .Q(\D_cache/cache[4][70] ), .QN(n1113) );
  DFFRX1 \D_cache/cache_reg[5][70]  ( .D(\D_cache/n1231 ), .CK(clk), .RN(n5706), .Q(\D_cache/cache[5][70] ), .QN(n2659) );
  DFFRX1 \D_cache/cache_reg[6][70]  ( .D(\D_cache/n1230 ), .CK(clk), .RN(n5906), .Q(\D_cache/cache[6][70] ), .QN(n667) );
  DFFRX1 \D_cache/cache_reg[7][70]  ( .D(\D_cache/n1229 ), .CK(clk), .RN(n5896), .Q(\D_cache/cache[7][70] ), .QN(n2238) );
  DFFRX1 \D_cache/cache_reg[0][71]  ( .D(\D_cache/n1228 ), .CK(clk), .RN(n5896), .Q(\D_cache/cache[0][71] ), .QN(n1322) );
  DFFRX1 \D_cache/cache_reg[1][71]  ( .D(\D_cache/n1227 ), .CK(clk), .RN(n5896), .Q(\D_cache/cache[1][71] ), .QN(n2851) );
  DFFRX1 \D_cache/cache_reg[2][71]  ( .D(\D_cache/n1226 ), .CK(clk), .RN(n5896), .Q(\D_cache/cache[2][71] ), .QN(n2119) );
  DFFRX1 \D_cache/cache_reg[3][71]  ( .D(\D_cache/n1225 ), .CK(clk), .RN(n5896), .Q(\D_cache/cache[3][71] ), .QN(n532) );
  DFFRX1 \D_cache/cache_reg[4][71]  ( .D(\D_cache/n1224 ), .CK(clk), .RN(n5895), .Q(\D_cache/cache[4][71] ), .QN(n1369) );
  DFFRX1 \D_cache/cache_reg[5][71]  ( .D(\D_cache/n1223 ), .CK(clk), .RN(n5895), .Q(\D_cache/cache[5][71] ), .QN(n2899) );
  DFFRX1 \D_cache/cache_reg[6][71]  ( .D(\D_cache/n1222 ), .CK(clk), .RN(n5895), .Q(\D_cache/cache[6][71] ), .QN(n1321) );
  DFFRX1 \D_cache/cache_reg[7][71]  ( .D(\D_cache/n1221 ), .CK(clk), .RN(n5895), .Q(\D_cache/cache[7][71] ), .QN(n2850) );
  DFFRX1 \D_cache/cache_reg[0][72]  ( .D(\D_cache/n1220 ), .CK(clk), .RN(n5895), .Q(\D_cache/cache[0][72] ), .QN(n1307) );
  DFFRX1 \D_cache/cache_reg[1][72]  ( .D(\D_cache/n1219 ), .CK(clk), .RN(n5895), .Q(\D_cache/cache[1][72] ), .QN(n2836) );
  DFFRX1 \D_cache/cache_reg[2][72]  ( .D(\D_cache/n1218 ), .CK(clk), .RN(n5895), .Q(\D_cache/cache[2][72] ), .QN(n771) );
  DFFRX1 \D_cache/cache_reg[3][72]  ( .D(\D_cache/n1217 ), .CK(clk), .RN(n5895), .Q(\D_cache/cache[3][72] ), .QN(n2333) );
  DFFRX1 \D_cache/cache_reg[4][72]  ( .D(\D_cache/n1216 ), .CK(clk), .RN(n5895), .Q(\D_cache/cache[4][72] ), .QN(n1358) );
  DFFRX1 \D_cache/cache_reg[5][72]  ( .D(\D_cache/n1215 ), .CK(clk), .RN(n5895), .Q(\D_cache/cache[5][72] ), .QN(n2888) );
  DFFRX1 \D_cache/cache_reg[6][72]  ( .D(\D_cache/n1214 ), .CK(clk), .RN(n5895), .Q(\D_cache/cache[6][72] ), .QN(n775) );
  DFFRX1 \D_cache/cache_reg[7][72]  ( .D(\D_cache/n1213 ), .CK(clk), .RN(n5895), .Q(\D_cache/cache[7][72] ), .QN(n2337) );
  DFFRX1 \D_cache/cache_reg[0][73]  ( .D(\D_cache/n1212 ), .CK(clk), .RN(n5894), .Q(\D_cache/cache[0][73] ), .QN(n810) );
  DFFRX1 \D_cache/cache_reg[1][73]  ( .D(\D_cache/n1211 ), .CK(clk), .RN(n5894), .Q(\D_cache/cache[1][73] ), .QN(n2373) );
  DFFRX1 \D_cache/cache_reg[2][73]  ( .D(\D_cache/n1210 ), .CK(clk), .RN(n5894), .Q(\D_cache/cache[2][73] ), .QN(n809) );
  DFFRX1 \D_cache/cache_reg[3][73]  ( .D(\D_cache/n1209 ), .CK(clk), .RN(n5894), .Q(\D_cache/cache[3][73] ), .QN(n2372) );
  DFFRX1 \D_cache/cache_reg[4][73]  ( .D(\D_cache/n1208 ), .CK(clk), .RN(n5894), .Q(\D_cache/cache[4][73] ), .QN(n2166) );
  DFFRX1 \D_cache/cache_reg[5][73]  ( .D(\D_cache/n1207 ), .CK(clk), .RN(n5894), .Q(\D_cache/cache[5][73] ), .QN(n592) );
  DFFRX1 \D_cache/cache_reg[6][73]  ( .D(\D_cache/n1206 ), .CK(clk), .RN(n5894), .Q(\D_cache/cache[6][73] ), .QN(n808) );
  DFFRX1 \D_cache/cache_reg[7][73]  ( .D(\D_cache/n1205 ), .CK(clk), .RN(n5894), .Q(\D_cache/cache[7][73] ), .QN(n2371) );
  DFFRX1 \D_cache/cache_reg[0][74]  ( .D(\D_cache/n1204 ), .CK(clk), .RN(n5894), .Q(\D_cache/cache[0][74] ), .QN(n1308) );
  DFFRX1 \D_cache/cache_reg[1][74]  ( .D(\D_cache/n1203 ), .CK(clk), .RN(n5894), .Q(\D_cache/cache[1][74] ), .QN(n2837) );
  DFFRX1 \D_cache/cache_reg[2][74]  ( .D(\D_cache/n1202 ), .CK(clk), .RN(n5894), .Q(\D_cache/cache[2][74] ), .QN(n1231) );
  DFFRX1 \D_cache/cache_reg[3][74]  ( .D(\D_cache/n1201 ), .CK(clk), .RN(n5894), .Q(\D_cache/cache[3][74] ), .QN(n2769) );
  DFFRX1 \D_cache/cache_reg[4][74]  ( .D(\D_cache/n1200 ), .CK(clk), .RN(n5893), .Q(\D_cache/cache[4][74] ), .QN(n1224) );
  DFFRX1 \D_cache/cache_reg[5][74]  ( .D(\D_cache/n1199 ), .CK(clk), .RN(n5893), .Q(\D_cache/cache[5][74] ), .QN(n2761) );
  DFFRX1 \D_cache/cache_reg[6][74]  ( .D(\D_cache/n1198 ), .CK(clk), .RN(n5893), .Q(\D_cache/cache[6][74] ), .QN(n1230) );
  DFFRX1 \D_cache/cache_reg[7][74]  ( .D(\D_cache/n1197 ), .CK(clk), .RN(n5893), .Q(\D_cache/cache[7][74] ), .QN(n2768) );
  DFFRX1 \D_cache/cache_reg[0][75]  ( .D(\D_cache/n1196 ), .CK(clk), .RN(n5893), .Q(\D_cache/cache[0][75] ), .QN(n1118) );
  DFFRX1 \D_cache/cache_reg[1][75]  ( .D(\D_cache/n1195 ), .CK(clk), .RN(n5893), .Q(\D_cache/cache[1][75] ), .QN(n2667) );
  DFFRX1 \D_cache/cache_reg[2][75]  ( .D(\D_cache/n1194 ), .CK(clk), .RN(n5893), .Q(\D_cache/cache[2][75] ), .QN(n1078) );
  DFFRX1 \D_cache/cache_reg[3][75]  ( .D(\D_cache/n1193 ), .CK(clk), .RN(n5893), .Q(\D_cache/cache[3][75] ), .QN(n2656) );
  DFFRX1 \D_cache/cache_reg[4][75]  ( .D(\D_cache/n1192 ), .CK(clk), .RN(n5893), .Q(\D_cache/cache[4][75] ), .QN(n1132) );
  DFFRX1 \D_cache/cache_reg[5][75]  ( .D(\D_cache/n1191 ), .CK(clk), .RN(n5893), .Q(\D_cache/cache[5][75] ), .QN(n2668) );
  DFFRX1 \D_cache/cache_reg[6][75]  ( .D(\D_cache/n1190 ), .CK(clk), .RN(n5893), .Q(\D_cache/cache[6][75] ), .QN(n1131) );
  DFFRX1 \D_cache/cache_reg[7][75]  ( .D(\D_cache/n1189 ), .CK(clk), .RN(n5893), .Q(\D_cache/cache[7][75] ), .QN(n2666) );
  DFFRX1 \D_cache/cache_reg[0][76]  ( .D(\D_cache/n1188 ), .CK(clk), .RN(n5892), .Q(\D_cache/cache[0][76] ), .QN(n659) );
  DFFRX1 \D_cache/cache_reg[1][76]  ( .D(\D_cache/n1187 ), .CK(clk), .RN(n5892), .Q(\D_cache/cache[1][76] ), .QN(n2245) );
  DFFRX1 \D_cache/cache_reg[2][76]  ( .D(\D_cache/n1186 ), .CK(clk), .RN(n5892), .Q(\D_cache/cache[2][76] ), .QN(n807) );
  DFFRX1 \D_cache/cache_reg[3][76]  ( .D(\D_cache/n1185 ), .CK(clk), .RN(n5892), .Q(\D_cache/cache[3][76] ), .QN(n2370) );
  DFFRX1 \D_cache/cache_reg[4][76]  ( .D(\D_cache/n1184 ), .CK(clk), .RN(n5892), .Q(\D_cache/cache[4][76] ), .QN(n2290) );
  DFFRX1 \D_cache/cache_reg[5][76]  ( .D(\D_cache/n1183 ), .CK(clk), .RN(n5892), .Q(\D_cache/cache[5][76] ), .QN(n721) );
  DFFRX1 \D_cache/cache_reg[6][76]  ( .D(\D_cache/n1182 ), .CK(clk), .RN(n5892), .Q(\D_cache/cache[6][76] ), .QN(n806) );
  DFFRX1 \D_cache/cache_reg[7][76]  ( .D(\D_cache/n1181 ), .CK(clk), .RN(n5892), .Q(\D_cache/cache[7][76] ), .QN(n2369) );
  DFFRX1 \D_cache/cache_reg[0][77]  ( .D(\D_cache/n1180 ), .CK(clk), .RN(n5892), .Q(\D_cache/cache[0][77] ), .QN(n660) );
  DFFRX1 \D_cache/cache_reg[1][77]  ( .D(\D_cache/n1179 ), .CK(clk), .RN(n5892), .Q(\D_cache/cache[1][77] ), .QN(n2248) );
  DFFRX1 \D_cache/cache_reg[2][77]  ( .D(\D_cache/n1178 ), .CK(clk), .RN(n5892), .Q(\D_cache/cache[2][77] ), .QN(n1261) );
  DFFRX1 \D_cache/cache_reg[3][77]  ( .D(\D_cache/n1177 ), .CK(clk), .RN(n5892), .Q(\D_cache/cache[3][77] ), .QN(n2803) );
  DFFRX1 \D_cache/cache_reg[4][77]  ( .D(\D_cache/n1176 ), .CK(clk), .RN(n5891), .Q(\D_cache/cache[4][77] ), .QN(n2771) );
  DFFRX1 \D_cache/cache_reg[5][77]  ( .D(\D_cache/n1175 ), .CK(clk), .RN(n5891), .Q(\D_cache/cache[5][77] ), .QN(n1137) );
  DFFRX1 \D_cache/cache_reg[6][77]  ( .D(\D_cache/n1174 ), .CK(clk), .RN(n5891), .Q(\D_cache/cache[6][77] ), .QN(n844) );
  DFFRX1 \D_cache/cache_reg[7][77]  ( .D(\D_cache/n1173 ), .CK(clk), .RN(n5891), .Q(\D_cache/cache[7][77] ), .QN(n2407) );
  DFFRX1 \D_cache/cache_reg[0][78]  ( .D(\D_cache/n1172 ), .CK(clk), .RN(n5891), .Q(\D_cache/cache[0][78] ), .QN(n657) );
  DFFRX1 \D_cache/cache_reg[1][78]  ( .D(\D_cache/n1171 ), .CK(clk), .RN(n5891), .Q(\D_cache/cache[1][78] ), .QN(n2240) );
  DFFRX1 \D_cache/cache_reg[2][78]  ( .D(\D_cache/n1170 ), .CK(clk), .RN(n5891), .Q(\D_cache/cache[2][78] ), .QN(n803) );
  DFFRX1 \D_cache/cache_reg[3][78]  ( .D(\D_cache/n1169 ), .CK(clk), .RN(n5891), .Q(\D_cache/cache[3][78] ), .QN(n2366) );
  DFFRX1 \D_cache/cache_reg[4][78]  ( .D(\D_cache/n1168 ), .CK(clk), .RN(n5891), .Q(\D_cache/cache[4][78] ), .QN(n2105) );
  DFFRX1 \D_cache/cache_reg[5][78]  ( .D(\D_cache/n1167 ), .CK(clk), .RN(n5891), .Q(\D_cache/cache[5][78] ), .QN(n482) );
  DFFRX1 \D_cache/cache_reg[6][78]  ( .D(\D_cache/n1166 ), .CK(clk), .RN(n5891), .Q(\D_cache/cache[6][78] ), .QN(n802) );
  DFFRX1 \D_cache/cache_reg[7][78]  ( .D(\D_cache/n1165 ), .CK(clk), .RN(n5890), .Q(\D_cache/cache[7][78] ), .QN(n2365) );
  DFFRX1 \D_cache/cache_reg[0][79]  ( .D(\D_cache/n1164 ), .CK(clk), .RN(n5890), .Q(\D_cache/cache[0][79] ), .QN(n656) );
  DFFRX1 \D_cache/cache_reg[1][79]  ( .D(\D_cache/n1163 ), .CK(clk), .RN(n5890), .Q(\D_cache/cache[1][79] ), .QN(n2237) );
  DFFRX1 \D_cache/cache_reg[2][79]  ( .D(\D_cache/n1162 ), .CK(clk), .RN(n5890), .Q(\D_cache/cache[2][79] ), .QN(n2074) );
  DFFRX1 \D_cache/cache_reg[3][79]  ( .D(\D_cache/n1161 ), .CK(clk), .RN(n5890), .Q(\D_cache/cache[3][79] ), .QN(n484) );
  DFFRX1 \D_cache/cache_reg[4][79]  ( .D(\D_cache/n1160 ), .CK(clk), .RN(n5890), .Q(\D_cache/cache[4][79] ), .QN(n2075) );
  DFFRX1 \D_cache/cache_reg[5][79]  ( .D(\D_cache/n1159 ), .CK(clk), .RN(n5890), .Q(\D_cache/cache[5][79] ), .QN(n487) );
  DFFRX1 \D_cache/cache_reg[6][79]  ( .D(\D_cache/n1158 ), .CK(clk), .RN(n5890), .Q(\D_cache/cache[6][79] ), .QN(n666) );
  DFFRX1 \D_cache/cache_reg[7][79]  ( .D(\D_cache/n1157 ), .CK(clk), .RN(n5890), .Q(\D_cache/cache[7][79] ), .QN(n2236) );
  DFFRX1 \D_cache/cache_reg[0][80]  ( .D(\D_cache/n1156 ), .CK(clk), .RN(n5890), .Q(\D_cache/cache[0][80] ), .QN(n801) );
  DFFRX1 \D_cache/cache_reg[1][80]  ( .D(\D_cache/n1155 ), .CK(clk), .RN(n5890), .Q(\D_cache/cache[1][80] ), .QN(n2364) );
  DFFRX1 \D_cache/cache_reg[2][80]  ( .D(\D_cache/n1154 ), .CK(clk), .RN(n5890), .Q(\D_cache/cache[2][80] ), .QN(n800) );
  DFFRX1 \D_cache/cache_reg[3][80]  ( .D(\D_cache/n1153 ), .CK(clk), .RN(n5889), .Q(\D_cache/cache[3][80] ), .QN(n2363) );
  DFFRX1 \D_cache/cache_reg[4][80]  ( .D(\D_cache/n1152 ), .CK(clk), .RN(n5889), .Q(\D_cache/cache[4][80] ), .QN(n1296) );
  DFFRX1 \D_cache/cache_reg[5][80]  ( .D(\D_cache/n1151 ), .CK(clk), .RN(n5889), .Q(\D_cache/cache[5][80] ), .QN(n2827) );
  DFFRX1 \D_cache/cache_reg[6][80]  ( .D(\D_cache/n1150 ), .CK(clk), .RN(n5889), .Q(\D_cache/cache[6][80] ), .QN(n799) );
  DFFRX1 \D_cache/cache_reg[7][80]  ( .D(\D_cache/n1149 ), .CK(clk), .RN(n5889), .Q(\D_cache/cache[7][80] ), .QN(n2362) );
  DFFRX1 \D_cache/cache_reg[0][81]  ( .D(\D_cache/n1148 ), .CK(clk), .RN(n5889), .Q(\D_cache/cache[0][81] ), .QN(n1115) );
  DFFRX1 \D_cache/cache_reg[1][81]  ( .D(\D_cache/n1147 ), .CK(clk), .RN(n5889), .Q(\D_cache/cache[1][81] ), .QN(n2662) );
  DFFRX1 \D_cache/cache_reg[2][81]  ( .D(\D_cache/n1146 ), .CK(clk), .RN(n5889), .Q(\D_cache/cache[2][81] ), .QN(n2073) );
  DFFRX1 \D_cache/cache_reg[3][81]  ( .D(\D_cache/n1145 ), .CK(clk), .RN(n5889), .Q(\D_cache/cache[3][81] ), .QN(n483) );
  DFFRX1 \D_cache/cache_reg[4][81]  ( .D(\D_cache/n1144 ), .CK(clk), .RN(n5889), .Q(\D_cache/cache[4][81] ), .QN(n663) );
  DFFRX1 \D_cache/cache_reg[5][81]  ( .D(\D_cache/n1143 ), .CK(clk), .RN(n5889), .Q(\D_cache/cache[5][81] ), .QN(n2233) );
  DFFRX1 \D_cache/cache_reg[6][81]  ( .D(\D_cache/n1142 ), .CK(clk), .RN(n5889), .Q(\D_cache/cache[6][81] ), .QN(n665) );
  DFFRX1 \D_cache/cache_reg[7][81]  ( .D(\D_cache/n1141 ), .CK(clk), .RN(n5888), .Q(\D_cache/cache[7][81] ), .QN(n2235) );
  DFFRX1 \D_cache/cache_reg[0][82]  ( .D(\D_cache/n1140 ), .CK(clk), .RN(n5888), .Q(\D_cache/cache[0][82] ), .QN(n2770) );
  DFFRX1 \D_cache/cache_reg[1][82]  ( .D(\D_cache/n1139 ), .CK(clk), .RN(n5888), .Q(\D_cache/cache[1][82] ), .QN(n1122) );
  DFFRX1 \D_cache/cache_reg[2][82]  ( .D(\D_cache/n1138 ), .CK(clk), .RN(n5888), .Q(\D_cache/cache[2][82] ), .QN(n662) );
  DFFRX1 \D_cache/cache_reg[3][82]  ( .D(\D_cache/n1137 ), .CK(clk), .RN(n5888), .Q(\D_cache/cache[3][82] ), .QN(n2231) );
  DFFRX1 \D_cache/cache_reg[4][82]  ( .D(\D_cache/n1136 ), .CK(clk), .RN(n5888), .Q(\D_cache/cache[4][82] ), .QN(n2071) );
  DFFRX1 \D_cache/cache_reg[5][82]  ( .D(\D_cache/n1135 ), .CK(clk), .RN(n5888), .Q(\D_cache/cache[5][82] ), .QN(n486) );
  DFFRX1 \D_cache/cache_reg[6][82]  ( .D(\D_cache/n1134 ), .CK(clk), .RN(n5888), .Q(\D_cache/cache[6][82] ), .QN(n661) );
  DFFRX1 \D_cache/cache_reg[7][82]  ( .D(\D_cache/n1133 ), .CK(clk), .RN(n5888), .Q(\D_cache/cache[7][82] ), .QN(n2250) );
  DFFRX1 \D_cache/cache_reg[1][83]  ( .D(\D_cache/n1131 ), .CK(clk), .RN(n5888), .Q(\D_cache/cache[1][83] ), .QN(n677) );
  DFFRX1 \D_cache/cache_reg[3][83]  ( .D(\D_cache/n1129 ), .CK(clk), .RN(n5887), .Q(\D_cache/cache[3][83] ), .QN(n1422) );
  DFFRX1 \D_cache/cache_reg[4][83]  ( .D(\D_cache/n1128 ), .CK(clk), .RN(n5887), .Q(\D_cache/cache[4][83] ), .QN(n652) );
  DFFRX1 \D_cache/cache_reg[5][83]  ( .D(\D_cache/n1127 ), .CK(clk), .RN(n5887), .Q(\D_cache/cache[5][83] ), .QN(n2228) );
  DFFRX1 \D_cache/cache_reg[6][83]  ( .D(\D_cache/n1126 ), .CK(clk), .RN(n5887), .Q(\D_cache/cache[6][83] ), .QN(n2131) );
  DFFRX1 \D_cache/cache_reg[7][83]  ( .D(\D_cache/n1125 ), .CK(clk), .RN(n5887), .Q(\D_cache/cache[7][83] ), .QN(n545) );
  DFFRX1 \D_cache/cache_reg[0][84]  ( .D(\D_cache/n1124 ), .CK(clk), .RN(n5887), .Q(\D_cache/cache[0][84] ), .QN(n1051) );
  DFFRX1 \D_cache/cache_reg[1][84]  ( .D(\D_cache/n1123 ), .CK(clk), .RN(n5887), .Q(\D_cache/cache[1][84] ), .QN(n2646) );
  DFFRX1 \D_cache/cache_reg[2][84]  ( .D(\D_cache/n1122 ), .CK(clk), .RN(n5887), .Q(\D_cache/cache[2][84] ), .QN(n669) );
  DFFRX1 \D_cache/cache_reg[3][84]  ( .D(\D_cache/n1121 ), .CK(clk), .RN(n5887), .Q(\D_cache/cache[3][84] ), .QN(n2241) );
  DFFRX1 \D_cache/cache_reg[4][84]  ( .D(\D_cache/n1120 ), .CK(clk), .RN(n5887), .Q(\D_cache/cache[4][84] ), .QN(n655) );
  DFFRX1 \D_cache/cache_reg[5][84]  ( .D(\D_cache/n1119 ), .CK(clk), .RN(n5887), .Q(\D_cache/cache[5][84] ), .QN(n2232) );
  DFFRX1 \D_cache/cache_reg[6][84]  ( .D(\D_cache/n1118 ), .CK(clk), .RN(n5887), .Q(\D_cache/cache[6][84] ), .QN(n705) );
  DFFRX1 \D_cache/cache_reg[7][84]  ( .D(\D_cache/n1117 ), .CK(clk), .RN(n5886), .Q(\D_cache/cache[7][84] ), .QN(n2273) );
  DFFRX1 \D_cache/cache_reg[0][85]  ( .D(\D_cache/n1116 ), .CK(clk), .RN(n5886), .Q(\D_cache/cache[0][85] ), .QN(n2767) );
  DFFRX1 \D_cache/cache_reg[1][85]  ( .D(\D_cache/n1115 ), .CK(clk), .RN(n5886), .Q(\D_cache/cache[1][85] ), .QN(n1121) );
  DFFRX1 \D_cache/cache_reg[2][85]  ( .D(\D_cache/n1114 ), .CK(clk), .RN(n5886), .Q(\D_cache/cache[2][85] ), .QN(n1128) );
  DFFRX1 \D_cache/cache_reg[3][85]  ( .D(\D_cache/n1113 ), .CK(clk), .RN(n5886), .Q(\D_cache/cache[3][85] ), .QN(n2661) );
  DFFRX1 \D_cache/cache_reg[4][85]  ( .D(\D_cache/n1112 ), .CK(clk), .RN(n5886), .Q(\D_cache/cache[4][85] ), .QN(n653) );
  DFFRX1 \D_cache/cache_reg[5][85]  ( .D(\D_cache/n1111 ), .CK(clk), .RN(n5886), .Q(\D_cache/cache[5][85] ), .QN(n2230) );
  DFFRX1 \D_cache/cache_reg[6][85]  ( .D(\D_cache/n1110 ), .CK(clk), .RN(n5891), .Q(\D_cache/cache[6][85] ), .QN(n1082) );
  DFFRX1 \D_cache/cache_reg[7][85]  ( .D(\D_cache/n1109 ), .CK(clk), .RN(n5906), .Q(\D_cache/cache[7][85] ), .QN(n2675) );
  DFFRX1 \D_cache/cache_reg[0][86]  ( .D(\D_cache/n1108 ), .CK(clk), .RN(n5906), .Q(\D_cache/cache[0][86] ), .QN(n1052) );
  DFFRX1 \D_cache/cache_reg[1][86]  ( .D(\D_cache/n1107 ), .CK(clk), .RN(n5906), .Q(\D_cache/cache[1][86] ), .QN(n2650) );
  DFFRX1 \D_cache/cache_reg[2][86]  ( .D(\D_cache/n1106 ), .CK(clk), .RN(n5906), .Q(\D_cache/cache[2][86] ), .QN(n819) );
  DFFRX1 \D_cache/cache_reg[3][86]  ( .D(\D_cache/n1105 ), .CK(clk), .RN(n5905), .Q(\D_cache/cache[3][86] ), .QN(n2382) );
  DFFRX1 \D_cache/cache_reg[4][86]  ( .D(\D_cache/n1104 ), .CK(clk), .RN(n5905), .Q(\D_cache/cache[4][86] ), .QN(n1716) );
  DFFRX1 \D_cache/cache_reg[5][86]  ( .D(\D_cache/n1103 ), .CK(clk), .RN(n5905), .Q(\D_cache/cache[5][86] ), .QN(n3314) );
  DFFRX1 \D_cache/cache_reg[6][86]  ( .D(\D_cache/n1102 ), .CK(clk), .RN(n5905), .Q(\D_cache/cache[6][86] ), .QN(n818) );
  DFFRX1 \D_cache/cache_reg[7][86]  ( .D(\D_cache/n1101 ), .CK(clk), .RN(n5905), .Q(\D_cache/cache[7][86] ), .QN(n2381) );
  DFFRX1 \D_cache/cache_reg[1][87]  ( .D(\D_cache/n1099 ), .CK(clk), .RN(n5905), .Q(\D_cache/cache[1][87] ), .QN(n1144) );
  DFFRX1 \D_cache/cache_reg[2][87]  ( .D(\D_cache/n1098 ), .CK(clk), .RN(n5905), .Q(\D_cache/cache[2][87] ), .QN(n1084) );
  DFFRX1 \D_cache/cache_reg[3][87]  ( .D(\D_cache/n1097 ), .CK(clk), .RN(n5905), .Q(\D_cache/cache[3][87] ), .QN(n2678) );
  DFFRX1 \D_cache/cache_reg[4][87]  ( .D(\D_cache/n1096 ), .CK(clk), .RN(n5905), .Q(\D_cache/cache[4][87] ), .QN(n2088) );
  DFFRX1 \D_cache/cache_reg[5][87]  ( .D(\D_cache/n1095 ), .CK(clk), .RN(n5905), .Q(\D_cache/cache[5][87] ), .QN(n501) );
  DFFRX1 \D_cache/cache_reg[6][87]  ( .D(\D_cache/n1094 ), .CK(clk), .RN(n5905), .Q(\D_cache/cache[6][87] ), .QN(n1081) );
  DFFRX1 \D_cache/cache_reg[7][87]  ( .D(\D_cache/n1093 ), .CK(clk), .RN(n5904), .Q(\D_cache/cache[7][87] ), .QN(n2674) );
  DFFRX1 \D_cache/cache_reg[0][88]  ( .D(\D_cache/n1092 ), .CK(clk), .RN(n5904), .Q(\D_cache/cache[0][88] ), .QN(n658) );
  DFFRX1 \D_cache/cache_reg[1][88]  ( .D(\D_cache/n1091 ), .CK(clk), .RN(n5904), .Q(\D_cache/cache[1][88] ), .QN(n2244) );
  DFFRX1 \D_cache/cache_reg[2][88]  ( .D(\D_cache/n1090 ), .CK(clk), .RN(n5904), .Q(\D_cache/cache[2][88] ), .QN(n671) );
  DFFRX1 \D_cache/cache_reg[3][88]  ( .D(\D_cache/n1089 ), .CK(clk), .RN(n5904), .Q(\D_cache/cache[3][88] ), .QN(n2243) );
  DFFRX1 \D_cache/cache_reg[4][88]  ( .D(\D_cache/n1088 ), .CK(clk), .RN(n5904), .Q(\D_cache/cache[4][88] ), .QN(n1133) );
  DFFRX1 \D_cache/cache_reg[5][88]  ( .D(\D_cache/n1087 ), .CK(clk), .RN(n5904), .Q(\D_cache/cache[5][88] ), .QN(n2669) );
  DFFRX1 \D_cache/cache_reg[6][88]  ( .D(\D_cache/n1086 ), .CK(clk), .RN(n5904), .Q(\D_cache/cache[6][88] ), .QN(n670) );
  DFFRX1 \D_cache/cache_reg[7][88]  ( .D(\D_cache/n1085 ), .CK(clk), .RN(n5904), .Q(\D_cache/cache[7][88] ), .QN(n2242) );
  DFFRX1 \D_cache/cache_reg[0][89]  ( .D(\D_cache/n1084 ), .CK(clk), .RN(n5904), .Q(\D_cache/cache[0][89] ), .QN(n2293) );
  DFFRX1 \D_cache/cache_reg[1][89]  ( .D(\D_cache/n1083 ), .CK(clk), .RN(n5904), .Q(\D_cache/cache[1][89] ), .QN(n676) );
  DFFRX1 \D_cache/cache_reg[2][89]  ( .D(\D_cache/n1082 ), .CK(clk), .RN(n5904), .Q(\D_cache/cache[2][89] ), .QN(n672) );
  DFFRX1 \D_cache/cache_reg[3][89]  ( .D(\D_cache/n1081 ), .CK(clk), .RN(n5903), .Q(\D_cache/cache[3][89] ), .QN(n2246) );
  DFFRX1 \D_cache/cache_reg[4][89]  ( .D(\D_cache/n1080 ), .CK(clk), .RN(n5903), .Q(\D_cache/cache[4][89] ), .QN(n1114) );
  DFFRX1 \D_cache/cache_reg[5][89]  ( .D(\D_cache/n1079 ), .CK(clk), .RN(n5903), .Q(\D_cache/cache[5][89] ), .QN(n2660) );
  DFFRX1 \D_cache/cache_reg[6][89]  ( .D(\D_cache/n1078 ), .CK(clk), .RN(n5903), .Q(\D_cache/cache[6][89] ), .QN(n664) );
  DFFRX1 \D_cache/cache_reg[7][89]  ( .D(\D_cache/n1077 ), .CK(clk), .RN(n5903), .Q(\D_cache/cache[7][89] ), .QN(n2234) );
  DFFRX1 \D_cache/cache_reg[0][90]  ( .D(\D_cache/n1076 ), .CK(clk), .RN(n5903), .Q(\D_cache/cache[0][90] ), .QN(n1330) );
  DFFRX1 \D_cache/cache_reg[1][90]  ( .D(\D_cache/n1075 ), .CK(clk), .RN(n5903), .Q(\D_cache/cache[1][90] ), .QN(n2859) );
  DFFRX1 \D_cache/cache_reg[2][90]  ( .D(\D_cache/n1074 ), .CK(clk), .RN(n5903), .Q(\D_cache/cache[2][90] ), .QN(n2144) );
  DFFRX1 \D_cache/cache_reg[3][90]  ( .D(\D_cache/n1073 ), .CK(clk), .RN(n5903), .Q(\D_cache/cache[3][90] ), .QN(n564) );
  DFFRX1 \D_cache/cache_reg[4][90]  ( .D(\D_cache/n1072 ), .CK(clk), .RN(n5903), .Q(\D_cache/cache[4][90] ), .QN(n2145) );
  DFFRX1 \D_cache/cache_reg[5][90]  ( .D(\D_cache/n1071 ), .CK(clk), .RN(n5903), .Q(\D_cache/cache[5][90] ), .QN(n565) );
  DFFRX1 \D_cache/cache_reg[6][90]  ( .D(\D_cache/n1070 ), .CK(clk), .RN(n5903), .Q(\D_cache/cache[6][90] ), .QN(n2152) );
  DFFRX1 \D_cache/cache_reg[7][90]  ( .D(\D_cache/n1069 ), .CK(clk), .RN(n5902), .Q(\D_cache/cache[7][90] ), .QN(n573) );
  DFFRX1 \D_cache/cache_reg[0][91]  ( .D(\D_cache/n1068 ), .CK(clk), .RN(n5902), .Q(\D_cache/cache[0][91] ), .QN(n798) );
  DFFRX1 \D_cache/cache_reg[1][91]  ( .D(\D_cache/n1067 ), .CK(clk), .RN(n5902), .Q(\D_cache/cache[1][91] ), .QN(n2361) );
  DFFRX1 \D_cache/cache_reg[2][91]  ( .D(\D_cache/n1066 ), .CK(clk), .RN(n5902), .Q(\D_cache/cache[2][91] ), .QN(n797) );
  DFFRX1 \D_cache/cache_reg[3][91]  ( .D(\D_cache/n1065 ), .CK(clk), .RN(n5902), .Q(\D_cache/cache[3][91] ), .QN(n2360) );
  DFFRX1 \D_cache/cache_reg[4][91]  ( .D(\D_cache/n1064 ), .CK(clk), .RN(n5902), .Q(\D_cache/cache[4][91] ), .QN(n1214) );
  DFFRX1 \D_cache/cache_reg[5][91]  ( .D(\D_cache/n1063 ), .CK(clk), .RN(n5902), .Q(\D_cache/cache[5][91] ), .QN(n2751) );
  DFFRX1 \D_cache/cache_reg[6][91]  ( .D(\D_cache/n1062 ), .CK(clk), .RN(n5902), .Q(\D_cache/cache[6][91] ), .QN(n2123) );
  DFFRX1 \D_cache/cache_reg[7][91]  ( .D(\D_cache/n1061 ), .CK(clk), .RN(n5902), .Q(\D_cache/cache[7][91] ), .QN(n536) );
  DFFRX1 \D_cache/cache_reg[0][92]  ( .D(\D_cache/n1060 ), .CK(clk), .RN(n5902), .Q(\D_cache/cache[0][92] ), .QN(n2161) );
  DFFRX1 \D_cache/cache_reg[1][92]  ( .D(\D_cache/n1059 ), .CK(clk), .RN(n5902), .Q(\D_cache/cache[1][92] ), .QN(n585) );
  DFFRX1 \D_cache/cache_reg[2][92]  ( .D(\D_cache/n1058 ), .CK(clk), .RN(n5902), .Q(\D_cache/cache[2][92] ), .QN(n1339) );
  DFFRX1 \D_cache/cache_reg[3][92]  ( .D(\D_cache/n1057 ), .CK(clk), .RN(n5901), .Q(\D_cache/cache[3][92] ), .QN(n2868) );
  DFFRX1 \D_cache/cache_reg[4][92]  ( .D(\D_cache/n1056 ), .CK(clk), .RN(n5901), .Q(\D_cache/cache[4][92] ), .QN(n1366) );
  DFFRX1 \D_cache/cache_reg[5][92]  ( .D(\D_cache/n1055 ), .CK(clk), .RN(n5901), .Q(\D_cache/cache[5][92] ), .QN(n2896) );
  DFFRX1 \D_cache/cache_reg[6][92]  ( .D(\D_cache/n1054 ), .CK(clk), .RN(n5901), .Q(\D_cache/cache[6][92] ), .QN(n2130) );
  DFFRX1 \D_cache/cache_reg[7][92]  ( .D(\D_cache/n1053 ), .CK(clk), .RN(n5901), .Q(\D_cache/cache[7][92] ), .QN(n544) );
  DFFRX1 \D_cache/cache_reg[0][93]  ( .D(\D_cache/n1052 ), .CK(clk), .RN(n5901), .Q(\D_cache/cache[0][93] ), .QN(n1117) );
  DFFRX1 \D_cache/cache_reg[1][93]  ( .D(\D_cache/n1051 ), .CK(clk), .RN(n5901), .Q(\D_cache/cache[1][93] ), .QN(n2665) );
  DFFRX1 \D_cache/cache_reg[2][93]  ( .D(\D_cache/n1050 ), .CK(clk), .RN(n5901), .Q(\D_cache/cache[2][93] ), .QN(n1130) );
  DFFRX1 \D_cache/cache_reg[3][93]  ( .D(\D_cache/n1049 ), .CK(clk), .RN(n5901), .Q(\D_cache/cache[3][93] ), .QN(n2664) );
  DFFRX1 \D_cache/cache_reg[4][93]  ( .D(\D_cache/n1048 ), .CK(clk), .RN(n5901), .Q(\D_cache/cache[4][93] ), .QN(n1134) );
  DFFRX1 \D_cache/cache_reg[5][93]  ( .D(\D_cache/n1047 ), .CK(clk), .RN(n5901), .Q(\D_cache/cache[5][93] ), .QN(n2670) );
  DFFRX1 \D_cache/cache_reg[6][93]  ( .D(\D_cache/n1046 ), .CK(clk), .RN(n5900), .Q(\D_cache/cache[6][93] ), .QN(n1129) );
  DFFRX1 \D_cache/cache_reg[7][93]  ( .D(\D_cache/n1045 ), .CK(clk), .RN(n5900), .Q(\D_cache/cache[7][93] ), .QN(n2663) );
  DFFRX1 \D_cache/cache_reg[0][94]  ( .D(\D_cache/n1044 ), .CK(clk), .RN(n5900), .Q(\D_cache/cache[0][94] ), .QN(n2785) );
  DFFRX1 \D_cache/cache_reg[1][94]  ( .D(\D_cache/n1043 ), .CK(clk), .RN(n5900), .Q(\D_cache/cache[1][94] ), .QN(n1126) );
  DFFRX1 \D_cache/cache_reg[2][94]  ( .D(\D_cache/n1042 ), .CK(clk), .RN(n5900), .Q(\D_cache/cache[2][94] ), .QN(n1176) );
  DFFRX1 \D_cache/cache_reg[3][94]  ( .D(\D_cache/n1041 ), .CK(clk), .RN(n5900), .Q(\D_cache/cache[3][94] ), .QN(n2726) );
  DFFRX1 \D_cache/cache_reg[4][94]  ( .D(\D_cache/n1040 ), .CK(clk), .RN(n5900), .Q(\D_cache/cache[4][94] ), .QN(n1456) );
  DFFRX1 \D_cache/cache_reg[5][94]  ( .D(\D_cache/n1039 ), .CK(clk), .RN(n5900), .Q(\D_cache/cache[5][94] ), .QN(n3026) );
  DFFRX1 \D_cache/cache_reg[6][94]  ( .D(\D_cache/n1038 ), .CK(clk), .RN(n5900), .Q(\D_cache/cache[6][94] ), .QN(n1142) );
  DFFRX1 \D_cache/cache_reg[7][94]  ( .D(\D_cache/n1037 ), .CK(clk), .RN(n5900), .Q(\D_cache/cache[7][94] ), .QN(n2704) );
  DFFRX1 \D_cache/cache_reg[0][95]  ( .D(\D_cache/n1036 ), .CK(clk), .RN(n5900), .Q(\D_cache/cache[0][95] ), .QN(n2737) );
  DFFRX1 \D_cache/cache_reg[1][95]  ( .D(\D_cache/n1035 ), .CK(clk), .RN(n5900), .Q(\D_cache/cache[1][95] ), .QN(n1138) );
  DFFRX1 \D_cache/cache_reg[2][95]  ( .D(\D_cache/n1034 ), .CK(clk), .RN(n5899), .Q(\D_cache/cache[2][95] ), .QN(n673) );
  DFFRX1 \D_cache/cache_reg[3][95]  ( .D(\D_cache/n1033 ), .CK(clk), .RN(n5899), .Q(\D_cache/cache[3][95] ), .QN(n2247) );
  DFFRX1 \D_cache/cache_reg[4][95]  ( .D(\D_cache/n1032 ), .CK(clk), .RN(n5899), .Q(\D_cache/cache[4][95] ), .QN(n1457) );
  DFFRX1 \D_cache/cache_reg[5][95]  ( .D(\D_cache/n1031 ), .CK(clk), .RN(n5899), .Q(\D_cache/cache[5][95] ), .QN(n3027) );
  DFFRX1 \D_cache/cache_reg[6][95]  ( .D(\D_cache/n1030 ), .CK(clk), .RN(n5899), .Q(\D_cache/cache[6][95] ), .QN(n1127) );
  DFFRX1 \D_cache/cache_reg[7][95]  ( .D(\D_cache/n1029 ), .CK(clk), .RN(n5899), .Q(\D_cache/cache[7][95] ), .QN(n2658) );
  DFFRX1 \D_cache/cache_reg[0][96]  ( .D(\D_cache/n1028 ), .CK(clk), .RN(n5899), .Q(\D_cache/cache[0][96] ), .QN(n1336) );
  DFFRX1 \D_cache/cache_reg[1][96]  ( .D(\D_cache/n1027 ), .CK(clk), .RN(n5899), .Q(\D_cache/cache[1][96] ), .QN(n2865) );
  DFFRX1 \D_cache/cache_reg[2][96]  ( .D(\D_cache/n1026 ), .CK(clk), .RN(n5899), .Q(\D_cache/cache[2][96] ), .QN(n1335) );
  DFFRX1 \D_cache/cache_reg[3][96]  ( .D(\D_cache/n1025 ), .CK(clk), .RN(n5899), .Q(\D_cache/cache[3][96] ), .QN(n2864) );
  DFFRX1 \D_cache/cache_reg[4][96]  ( .D(\D_cache/n1024 ), .CK(clk), .RN(n5899), .Q(\D_cache/cache[4][96] ), .QN(n1362) );
  DFFRX1 \D_cache/cache_reg[5][96]  ( .D(\D_cache/n1023 ), .CK(clk), .RN(n5899), .Q(\D_cache/cache[5][96] ), .QN(n2892) );
  DFFRX1 \D_cache/cache_reg[6][96]  ( .D(\D_cache/n1022 ), .CK(clk), .RN(n5898), .Q(\D_cache/cache[6][96] ), .QN(n741) );
  DFFRX1 \D_cache/cache_reg[7][96]  ( .D(\D_cache/n1021 ), .CK(clk), .RN(n5898), .Q(\D_cache/cache[7][96] ), .QN(n2302) );
  DFFRX1 \D_cache/cache_reg[0][97]  ( .D(\D_cache/n1020 ), .CK(clk), .RN(n5898), .Q(\D_cache/cache[0][97] ), .QN(n1332) );
  DFFRX1 \D_cache/cache_reg[1][97]  ( .D(\D_cache/n1019 ), .CK(clk), .RN(n5898), .Q(\D_cache/cache[1][97] ), .QN(n2861) );
  DFFRX1 \D_cache/cache_reg[2][97]  ( .D(\D_cache/n1018 ), .CK(clk), .RN(n5898), .Q(\D_cache/cache[2][97] ), .QN(n2117) );
  DFFRX1 \D_cache/cache_reg[3][97]  ( .D(\D_cache/n1017 ), .CK(clk), .RN(n5898), .Q(\D_cache/cache[3][97] ), .QN(n530) );
  DFFRX1 \D_cache/cache_reg[4][97]  ( .D(\D_cache/n1016 ), .CK(clk), .RN(n5898), .Q(\D_cache/cache[4][97] ), .QN(n758) );
  DFFRX1 \D_cache/cache_reg[5][97]  ( .D(\D_cache/n1015 ), .CK(clk), .RN(n5898), .Q(\D_cache/cache[5][97] ), .QN(n2319) );
  DFFRX1 \D_cache/cache_reg[6][97]  ( .D(\D_cache/n1014 ), .CK(clk), .RN(n5898), .Q(\D_cache/cache[6][97] ), .QN(n2129) );
  DFFRX1 \D_cache/cache_reg[7][97]  ( .D(\D_cache/n1013 ), .CK(clk), .RN(n5898), .Q(\D_cache/cache[7][97] ), .QN(n543) );
  DFFRX1 \D_cache/cache_reg[0][98]  ( .D(\D_cache/n1012 ), .CK(clk), .RN(n5898), .Q(\D_cache/cache[0][98] ), .QN(n1348) );
  DFFRX1 \D_cache/cache_reg[1][98]  ( .D(\D_cache/n1011 ), .CK(clk), .RN(n5898), .Q(\D_cache/cache[1][98] ), .QN(n2877) );
  DFFRX1 \D_cache/cache_reg[2][98]  ( .D(\D_cache/n1010 ), .CK(clk), .RN(n5897), .Q(\D_cache/cache[2][98] ), .QN(n1347) );
  DFFRX1 \D_cache/cache_reg[3][98]  ( .D(\D_cache/n1009 ), .CK(clk), .RN(n5897), .Q(\D_cache/cache[3][98] ), .QN(n2876) );
  DFFRX1 \D_cache/cache_reg[4][98]  ( .D(\D_cache/n1008 ), .CK(clk), .RN(n5897), .Q(\D_cache/cache[4][98] ), .QN(n1360) );
  DFFRX1 \D_cache/cache_reg[5][98]  ( .D(\D_cache/n1007 ), .CK(clk), .RN(n5897), .Q(\D_cache/cache[5][98] ), .QN(n2890) );
  DFFRX1 \D_cache/cache_reg[6][98]  ( .D(\D_cache/n1006 ), .CK(clk), .RN(n5897), .Q(\D_cache/cache[6][98] ), .QN(n1346) );
  DFFRX1 \D_cache/cache_reg[7][98]  ( .D(\D_cache/n1005 ), .CK(clk), .RN(n5897), .Q(\D_cache/cache[7][98] ), .QN(n2875) );
  DFFRX1 \D_cache/cache_reg[0][99]  ( .D(\D_cache/n1004 ), .CK(clk), .RN(n5897), .Q(\D_cache/cache[0][99] ), .QN(n763) );
  DFFRX1 \D_cache/cache_reg[1][99]  ( .D(\D_cache/n1003 ), .CK(clk), .RN(n5897), .Q(\D_cache/cache[1][99] ), .QN(n2325) );
  DFFRX1 \D_cache/cache_reg[2][99]  ( .D(\D_cache/n1002 ), .CK(clk), .RN(n5897), .Q(\D_cache/cache[2][99] ), .QN(n1221) );
  DFFRX1 \D_cache/cache_reg[3][99]  ( .D(\D_cache/n1001 ), .CK(clk), .RN(n5897), .Q(\D_cache/cache[3][99] ), .QN(n2758) );
  DFFRX1 \D_cache/cache_reg[4][99]  ( .D(\D_cache/n1000 ), .CK(clk), .RN(n5897), .Q(\D_cache/cache[4][99] ), .QN(n753) );
  DFFRX1 \D_cache/cache_reg[5][99]  ( .D(\D_cache/n999 ), .CK(clk), .RN(n5897), 
        .Q(\D_cache/cache[5][99] ), .QN(n2314) );
  DFFRX1 \D_cache/cache_reg[6][99]  ( .D(\D_cache/n998 ), .CK(clk), .RN(n5896), 
        .Q(\D_cache/cache[6][99] ), .QN(n762) );
  DFFRX1 \D_cache/cache_reg[7][99]  ( .D(\D_cache/n997 ), .CK(clk), .RN(n5896), 
        .Q(\D_cache/cache[7][99] ), .QN(n2324) );
  DFFRX1 \D_cache/cache_reg[0][100]  ( .D(\D_cache/n996 ), .CK(clk), .RN(n5896), .Q(\D_cache/cache[0][100] ), .QN(n822) );
  DFFRX1 \D_cache/cache_reg[1][100]  ( .D(\D_cache/n995 ), .CK(clk), .RN(n5896), .Q(\D_cache/cache[1][100] ), .QN(n2385) );
  DFFRX1 \D_cache/cache_reg[2][100]  ( .D(\D_cache/n994 ), .CK(clk), .RN(n5896), .Q(\D_cache/cache[2][100] ), .QN(n1245) );
  DFFRX1 \D_cache/cache_reg[3][100]  ( .D(\D_cache/n993 ), .CK(clk), .RN(n5896), .Q(\D_cache/cache[3][100] ), .QN(n2787) );
  DFFRX1 \D_cache/cache_reg[4][100]  ( .D(\D_cache/n992 ), .CK(clk), .RN(n5896), .Q(\D_cache/cache[4][100] ), .QN(n1357) );
  DFFRX1 \D_cache/cache_reg[5][100]  ( .D(\D_cache/n991 ), .CK(clk), .RN(n5901), .Q(\D_cache/cache[5][100] ), .QN(n2887) );
  DFFRX1 \D_cache/cache_reg[6][100]  ( .D(\D_cache/n990 ), .CK(clk), .RN(n5876), .Q(\D_cache/cache[6][100] ), .QN(n821) );
  DFFRX1 \D_cache/cache_reg[7][100]  ( .D(\D_cache/n989 ), .CK(clk), .RN(n5876), .Q(\D_cache/cache[7][100] ), .QN(n2384) );
  DFFRX1 \D_cache/cache_reg[0][101]  ( .D(\D_cache/n988 ), .CK(clk), .RN(n5876), .Q(\D_cache/cache[0][101] ), .QN(n1178) );
  DFFRX1 \D_cache/cache_reg[1][101]  ( .D(\D_cache/n987 ), .CK(clk), .RN(n5876), .Q(\D_cache/cache[1][101] ), .QN(n2925) );
  DFFRX1 \D_cache/cache_reg[2][101]  ( .D(\D_cache/n986 ), .CK(clk), .RN(n5876), .Q(\D_cache/cache[2][101] ), .QN(n1249) );
  DFFRX1 \D_cache/cache_reg[3][101]  ( .D(\D_cache/n985 ), .CK(clk), .RN(n5875), .Q(\D_cache/cache[3][101] ), .QN(n2791) );
  DFFRX1 \D_cache/cache_reg[4][101]  ( .D(\D_cache/n984 ), .CK(clk), .RN(n5875), .Q(\D_cache/cache[4][101] ), .QN(n1717) );
  DFFRX1 \D_cache/cache_reg[5][101]  ( .D(\D_cache/n983 ), .CK(clk), .RN(n5875), .Q(\D_cache/cache[5][101] ), .QN(n3315) );
  DFFRX1 \D_cache/cache_reg[6][101]  ( .D(\D_cache/n982 ), .CK(clk), .RN(n5875), .Q(\D_cache/cache[6][101] ), .QN(n2294) );
  DFFRX1 \D_cache/cache_reg[7][101]  ( .D(\D_cache/n981 ), .CK(clk), .RN(n5875), .Q(\D_cache/cache[7][101] ), .QN(n732) );
  DFFRX1 \D_cache/cache_reg[1][102]  ( .D(\D_cache/n979 ), .CK(clk), .RN(n5875), .Q(\D_cache/cache[1][102] ), .QN(n1194) );
  DFFRX1 \D_cache/cache_reg[2][102]  ( .D(\D_cache/n978 ), .CK(clk), .RN(n5875), .Q(\D_cache/cache[2][102] ), .QN(n1156) );
  DFFRX1 \D_cache/cache_reg[3][102]  ( .D(\D_cache/n977 ), .CK(clk), .RN(n5875), .Q(\D_cache/cache[3][102] ), .QN(n2713) );
  DFFRX1 \D_cache/cache_reg[4][102]  ( .D(\D_cache/n976 ), .CK(clk), .RN(n5875), .Q(\D_cache/cache[4][102] ), .QN(n1162) );
  DFFRX1 \D_cache/cache_reg[5][102]  ( .D(\D_cache/n975 ), .CK(clk), .RN(n5875), .Q(\D_cache/cache[5][102] ), .QN(n2718) );
  DFFRX1 \D_cache/cache_reg[6][102]  ( .D(\D_cache/n974 ), .CK(clk), .RN(n5875), .Q(\D_cache/cache[6][102] ), .QN(n1155) );
  DFFRX1 \D_cache/cache_reg[7][102]  ( .D(\D_cache/n973 ), .CK(clk), .RN(n5874), .Q(\D_cache/cache[7][102] ), .QN(n2712) );
  DFFRX1 \D_cache/cache_reg[0][103]  ( .D(\D_cache/n972 ), .CK(clk), .RN(n5874), .Q(\D_cache/cache[0][103] ), .QN(n1338) );
  DFFRX1 \D_cache/cache_reg[1][103]  ( .D(\D_cache/n971 ), .CK(clk), .RN(n5874), .Q(\D_cache/cache[1][103] ), .QN(n2867) );
  DFFRX1 \D_cache/cache_reg[2][103]  ( .D(\D_cache/n970 ), .CK(clk), .RN(n5874), .Q(\D_cache/cache[2][103] ), .QN(n1213) );
  DFFRX1 \D_cache/cache_reg[3][103]  ( .D(\D_cache/n969 ), .CK(clk), .RN(n5874), .Q(\D_cache/cache[3][103] ), .QN(n2750) );
  DFFRX1 \D_cache/cache_reg[4][103]  ( .D(\D_cache/n968 ), .CK(clk), .RN(n5874), .Q(\D_cache/cache[4][103] ), .QN(n1375) );
  DFFRX1 \D_cache/cache_reg[5][103]  ( .D(\D_cache/n967 ), .CK(clk), .RN(n5874), .Q(\D_cache/cache[5][103] ), .QN(n2905) );
  DFFRX1 \D_cache/cache_reg[6][103]  ( .D(\D_cache/n966 ), .CK(clk), .RN(n5874), .Q(\D_cache/cache[6][103] ), .QN(n1337) );
  DFFRX1 \D_cache/cache_reg[7][103]  ( .D(\D_cache/n965 ), .CK(clk), .RN(n5874), .Q(\D_cache/cache[7][103] ), .QN(n2866) );
  DFFRX1 \D_cache/cache_reg[0][104]  ( .D(\D_cache/n964 ), .CK(clk), .RN(n5874), .Q(\D_cache/cache[0][104] ), .QN(n1318) );
  DFFRX1 \D_cache/cache_reg[1][104]  ( .D(\D_cache/n963 ), .CK(clk), .RN(n5874), .Q(\D_cache/cache[1][104] ), .QN(n2847) );
  DFFRX1 \D_cache/cache_reg[2][104]  ( .D(\D_cache/n962 ), .CK(clk), .RN(n5874), .Q(\D_cache/cache[2][104] ), .QN(n1317) );
  DFFRX1 \D_cache/cache_reg[3][104]  ( .D(\D_cache/n961 ), .CK(clk), .RN(n5873), .Q(\D_cache/cache[3][104] ), .QN(n2846) );
  DFFRX1 \D_cache/cache_reg[4][104]  ( .D(\D_cache/n960 ), .CK(clk), .RN(n5873), .Q(\D_cache/cache[4][104] ), .QN(n1361) );
  DFFRX1 \D_cache/cache_reg[5][104]  ( .D(\D_cache/n959 ), .CK(clk), .RN(n5873), .Q(\D_cache/cache[5][104] ), .QN(n2891) );
  DFFRX1 \D_cache/cache_reg[6][104]  ( .D(\D_cache/n958 ), .CK(clk), .RN(n5873), .Q(\D_cache/cache[6][104] ), .QN(n1226) );
  DFFRX1 \D_cache/cache_reg[7][104]  ( .D(\D_cache/n957 ), .CK(clk), .RN(n5873), .Q(\D_cache/cache[7][104] ), .QN(n2763) );
  DFFRX1 \D_cache/cache_reg[1][105]  ( .D(\D_cache/n955 ), .CK(clk), .RN(n5873), .Q(\D_cache/cache[1][105] ), .QN(n847) );
  DFFRX1 \D_cache/cache_reg[2][105]  ( .D(\D_cache/n954 ), .CK(clk), .RN(n5873), .Q(\D_cache/cache[2][105] ), .QN(n1331) );
  DFFRX1 \D_cache/cache_reg[3][105]  ( .D(\D_cache/n953 ), .CK(clk), .RN(n5873), .Q(\D_cache/cache[3][105] ), .QN(n2860) );
  DFFRX1 \D_cache/cache_reg[4][105]  ( .D(\D_cache/n952 ), .CK(clk), .RN(n5873), .Q(\D_cache/cache[4][105] ), .QN(n1119) );
  DFFRX1 \D_cache/cache_reg[5][105]  ( .D(\D_cache/n951 ), .CK(clk), .RN(n5873), .Q(\D_cache/cache[5][105] ), .QN(n2655) );
  DFFRX1 \D_cache/cache_reg[6][105]  ( .D(\D_cache/n950 ), .CK(clk), .RN(n5873), .Q(\D_cache/cache[6][105] ), .QN(n1116) );
  DFFRX1 \D_cache/cache_reg[7][105]  ( .D(\D_cache/n949 ), .CK(clk), .RN(n5872), .Q(\D_cache/cache[7][105] ), .QN(n2654) );
  DFFRX1 \D_cache/cache_reg[0][106]  ( .D(\D_cache/n948 ), .CK(clk), .RN(n5872), .Q(\D_cache/cache[0][106] ), .QN(n1208) );
  DFFRX1 \D_cache/cache_reg[1][106]  ( .D(\D_cache/n947 ), .CK(clk), .RN(n5872), .Q(\D_cache/cache[1][106] ), .QN(n2745) );
  DFFRX1 \D_cache/cache_reg[2][106]  ( .D(\D_cache/n946 ), .CK(clk), .RN(n5872), .Q(\D_cache/cache[2][106] ), .QN(n1324) );
  DFFRX1 \D_cache/cache_reg[3][106]  ( .D(\D_cache/n945 ), .CK(clk), .RN(n5872), .Q(\D_cache/cache[3][106] ), .QN(n2853) );
  DFFRX1 \D_cache/cache_reg[4][106]  ( .D(\D_cache/n944 ), .CK(clk), .RN(n5872), .Q(\D_cache/cache[4][106] ), .QN(n1223) );
  DFFRX1 \D_cache/cache_reg[5][106]  ( .D(\D_cache/n943 ), .CK(clk), .RN(n5872), .Q(\D_cache/cache[5][106] ), .QN(n2760) );
  DFFRX1 \D_cache/cache_reg[6][106]  ( .D(\D_cache/n942 ), .CK(clk), .RN(n5872), .Q(\D_cache/cache[6][106] ), .QN(n1323) );
  DFFRX1 \D_cache/cache_reg[7][106]  ( .D(\D_cache/n941 ), .CK(clk), .RN(n5872), .Q(\D_cache/cache[7][106] ), .QN(n2852) );
  DFFRX1 \D_cache/cache_reg[1][107]  ( .D(\D_cache/n939 ), .CK(clk), .RN(n5872), .Q(\D_cache/cache[1][107] ), .QN(n1192) );
  DFFRX1 \D_cache/cache_reg[2][107]  ( .D(\D_cache/n938 ), .CK(clk), .RN(n5872), .Q(\D_cache/cache[2][107] ), .QN(n1153) );
  DFFRX1 \D_cache/cache_reg[3][107]  ( .D(\D_cache/n937 ), .CK(clk), .RN(n5871), .Q(\D_cache/cache[3][107] ), .QN(n2710) );
  DFFRX1 \D_cache/cache_reg[4][107]  ( .D(\D_cache/n936 ), .CK(clk), .RN(n5871), .Q(\D_cache/cache[4][107] ), .QN(n2681) );
  DFFRX1 \D_cache/cache_reg[5][107]  ( .D(\D_cache/n935 ), .CK(clk), .RN(n5871), .Q(\D_cache/cache[5][107] ), .QN(n1125) );
  DFFRX1 \D_cache/cache_reg[6][107]  ( .D(\D_cache/n934 ), .CK(clk), .RN(n5871), .Q(\D_cache/cache[6][107] ), .QN(n1152) );
  DFFRX1 \D_cache/cache_reg[7][107]  ( .D(\D_cache/n933 ), .CK(clk), .RN(n5871), .Q(\D_cache/cache[7][107] ), .QN(n2709) );
  DFFRX1 \D_cache/cache_reg[1][108]  ( .D(\D_cache/n931 ), .CK(clk), .RN(n5871), .Q(\D_cache/cache[1][108] ), .QN(n513) );
  DFFRX1 \D_cache/cache_reg[2][108]  ( .D(\D_cache/n930 ), .CK(clk), .RN(n5871), .Q(\D_cache/cache[2][108] ), .QN(n736) );
  DFFRX1 \D_cache/cache_reg[3][108]  ( .D(\D_cache/n929 ), .CK(clk), .RN(n5871), .Q(\D_cache/cache[3][108] ), .QN(n2295) );
  DFFRX1 \D_cache/cache_reg[4][108]  ( .D(\D_cache/n928 ), .CK(clk), .RN(n5871), .Q(\D_cache/cache[4][108] ), .QN(n739) );
  DFFRX1 \D_cache/cache_reg[5][108]  ( .D(\D_cache/n927 ), .CK(clk), .RN(n5871), .Q(\D_cache/cache[5][108] ), .QN(n2300) );
  DFFRX1 \D_cache/cache_reg[6][108]  ( .D(\D_cache/n926 ), .CK(clk), .RN(n5870), .Q(\D_cache/cache[6][108] ), .QN(n738) );
  DFFRX1 \D_cache/cache_reg[7][108]  ( .D(\D_cache/n925 ), .CK(clk), .RN(n5870), .Q(\D_cache/cache[7][108] ), .QN(n2297) );
  DFFRX1 \D_cache/cache_reg[0][109]  ( .D(\D_cache/n924 ), .CK(clk), .RN(n5870), .Q(\D_cache/cache[0][109] ), .QN(n1298) );
  DFFRX1 \D_cache/cache_reg[1][109]  ( .D(\D_cache/n923 ), .CK(clk), .RN(n5870), .Q(\D_cache/cache[1][109] ), .QN(n2829) );
  DFFRX1 \D_cache/cache_reg[2][109]  ( .D(\D_cache/n922 ), .CK(clk), .RN(n5870), .Q(\D_cache/cache[2][109] ), .QN(n1343) );
  DFFRX1 \D_cache/cache_reg[3][109]  ( .D(\D_cache/n921 ), .CK(clk), .RN(n5870), .Q(\D_cache/cache[3][109] ), .QN(n2872) );
  DFFRX1 \D_cache/cache_reg[4][109]  ( .D(\D_cache/n920 ), .CK(clk), .RN(n5870), .Q(\D_cache/cache[4][109] ), .QN(n2108) );
  DFFRX1 \D_cache/cache_reg[5][109]  ( .D(\D_cache/n919 ), .CK(clk), .RN(n5870), .Q(\D_cache/cache[5][109] ), .QN(n521) );
  DFFRX1 \D_cache/cache_reg[6][109]  ( .D(\D_cache/n918 ), .CK(clk), .RN(n5870), .Q(\D_cache/cache[6][109] ), .QN(n1299) );
  DFFRX1 \D_cache/cache_reg[7][109]  ( .D(\D_cache/n917 ), .CK(clk), .RN(n5870), .Q(\D_cache/cache[7][109] ), .QN(n2830) );
  DFFRX1 \D_cache/cache_reg[0][110]  ( .D(\D_cache/n916 ), .CK(clk), .RN(n5870), .Q(\D_cache/cache[0][110] ), .QN(n1344) );
  DFFRX1 \D_cache/cache_reg[1][110]  ( .D(\D_cache/n915 ), .CK(clk), .RN(n5870), .Q(\D_cache/cache[1][110] ), .QN(n2873) );
  DFFRX1 \D_cache/cache_reg[3][110]  ( .D(\D_cache/n913 ), .CK(clk), .RN(n5869), .Q(\D_cache/cache[3][110] ), .QN(n1290) );
  DFFRX1 \D_cache/cache_reg[4][110]  ( .D(\D_cache/n912 ), .CK(clk), .RN(n5869), .Q(\D_cache/cache[4][110] ), .QN(n2107) );
  DFFRX1 \D_cache/cache_reg[5][110]  ( .D(\D_cache/n911 ), .CK(clk), .RN(n5869), .Q(\D_cache/cache[5][110] ), .QN(n520) );
  DFFRX1 \D_cache/cache_reg[6][110]  ( .D(\D_cache/n910 ), .CK(clk), .RN(n5869), .Q(\D_cache/cache[6][110] ), .QN(n743) );
  DFFRX1 \D_cache/cache_reg[7][110]  ( .D(\D_cache/n909 ), .CK(clk), .RN(n5869), .Q(\D_cache/cache[7][110] ), .QN(n2304) );
  DFFRX1 \D_cache/cache_reg[0][111]  ( .D(\D_cache/n908 ), .CK(clk), .RN(n5869), .Q(\D_cache/cache[0][111] ), .QN(n1222) );
  DFFRX1 \D_cache/cache_reg[1][111]  ( .D(\D_cache/n907 ), .CK(clk), .RN(n5869), .Q(\D_cache/cache[1][111] ), .QN(n2759) );
  DFFRX1 \D_cache/cache_reg[2][111]  ( .D(\D_cache/n906 ), .CK(clk), .RN(n5869), .Q(\D_cache/cache[2][111] ), .QN(n1329) );
  DFFRX1 \D_cache/cache_reg[3][111]  ( .D(\D_cache/n905 ), .CK(clk), .RN(n5869), .Q(\D_cache/cache[3][111] ), .QN(n2858) );
  DFFRX1 \D_cache/cache_reg[4][111]  ( .D(\D_cache/n904 ), .CK(clk), .RN(n5869), .Q(\D_cache/cache[4][111] ), .QN(n764) );
  DFFRX1 \D_cache/cache_reg[5][111]  ( .D(\D_cache/n903 ), .CK(clk), .RN(n5869), .Q(\D_cache/cache[5][111] ), .QN(n2326) );
  DFFRX1 \D_cache/cache_reg[6][111]  ( .D(\D_cache/n902 ), .CK(clk), .RN(n5868), .Q(\D_cache/cache[6][111] ), .QN(n1328) );
  DFFRX1 \D_cache/cache_reg[7][111]  ( .D(\D_cache/n901 ), .CK(clk), .RN(n5868), .Q(\D_cache/cache[7][111] ), .QN(n2857) );
  DFFRX1 \D_cache/cache_reg[1][112]  ( .D(\D_cache/n899 ), .CK(clk), .RN(n5868), .Q(\D_cache/cache[1][112] ), .QN(n1195) );
  DFFRX1 \D_cache/cache_reg[2][112]  ( .D(\D_cache/n898 ), .CK(clk), .RN(n5868), .Q(\D_cache/cache[2][112] ), .QN(n684) );
  DFFRX1 \D_cache/cache_reg[3][112]  ( .D(\D_cache/n897 ), .CK(clk), .RN(n5868), .Q(\D_cache/cache[3][112] ), .QN(n2256) );
  DFFRX1 \D_cache/cache_reg[4][112]  ( .D(\D_cache/n896 ), .CK(clk), .RN(n5868), .Q(\D_cache/cache[4][112] ), .QN(n1164) );
  DFFRX1 \D_cache/cache_reg[5][112]  ( .D(\D_cache/n895 ), .CK(clk), .RN(n5868), .Q(\D_cache/cache[5][112] ), .QN(n2720) );
  DFFRX1 \D_cache/cache_reg[6][112]  ( .D(\D_cache/n894 ), .CK(clk), .RN(n5868), .Q(\D_cache/cache[6][112] ), .QN(n694) );
  DFFRX1 \D_cache/cache_reg[7][112]  ( .D(\D_cache/n893 ), .CK(clk), .RN(n5868), .Q(\D_cache/cache[7][112] ), .QN(n2263) );
  DFFRX1 \D_cache/cache_reg[0][113]  ( .D(\D_cache/n892 ), .CK(clk), .RN(n5868), .Q(\D_cache/cache[0][113] ), .QN(n827) );
  DFFRX1 \D_cache/cache_reg[1][113]  ( .D(\D_cache/n891 ), .CK(clk), .RN(n5868), .Q(\D_cache/cache[1][113] ), .QN(n2390) );
  DFFRX1 \D_cache/cache_reg[2][113]  ( .D(\D_cache/n890 ), .CK(clk), .RN(n5867), .Q(\D_cache/cache[2][113] ), .QN(n749) );
  DFFRX1 \D_cache/cache_reg[3][113]  ( .D(\D_cache/n889 ), .CK(clk), .RN(n5867), .Q(\D_cache/cache[3][113] ), .QN(n2310) );
  DFFRX1 \D_cache/cache_reg[4][113]  ( .D(\D_cache/n888 ), .CK(clk), .RN(n5867), .Q(\D_cache/cache[4][113] ), .QN(n755) );
  DFFRX1 \D_cache/cache_reg[5][113]  ( .D(\D_cache/n887 ), .CK(clk), .RN(n5867), .Q(\D_cache/cache[5][113] ), .QN(n2316) );
  DFFRX1 \D_cache/cache_reg[6][113]  ( .D(\D_cache/n886 ), .CK(clk), .RN(n5867), .Q(\D_cache/cache[6][113] ), .QN(n826) );
  DFFRX1 \D_cache/cache_reg[7][113]  ( .D(\D_cache/n885 ), .CK(clk), .RN(n5867), .Q(\D_cache/cache[7][113] ), .QN(n2389) );
  DFFRX1 \D_cache/cache_reg[1][114]  ( .D(\D_cache/n883 ), .CK(clk), .RN(n5867), .Q(\D_cache/cache[1][114] ), .QN(n1139) );
  DFFRX1 \D_cache/cache_reg[2][114]  ( .D(\D_cache/n882 ), .CK(clk), .RN(n5867), .Q(\D_cache/cache[2][114] ), .QN(n1154) );
  DFFRX1 \D_cache/cache_reg[3][114]  ( .D(\D_cache/n881 ), .CK(clk), .RN(n5867), .Q(\D_cache/cache[3][114] ), .QN(n2711) );
  DFFRX1 \D_cache/cache_reg[4][114]  ( .D(\D_cache/n880 ), .CK(clk), .RN(n5867), .Q(\D_cache/cache[4][114] ), .QN(n683) );
  DFFRX1 \D_cache/cache_reg[5][114]  ( .D(\D_cache/n879 ), .CK(clk), .RN(n5867), .Q(\D_cache/cache[5][114] ), .QN(n2255) );
  DFFRX1 \D_cache/cache_reg[6][114]  ( .D(\D_cache/n878 ), .CK(clk), .RN(n5866), .Q(\D_cache/cache[6][114] ), .QN(n679) );
  DFFRX1 \D_cache/cache_reg[7][114]  ( .D(\D_cache/n877 ), .CK(clk), .RN(n5866), .Q(\D_cache/cache[7][114] ), .QN(n2251) );
  DFFRX1 \D_cache/cache_reg[0][115]  ( .D(\D_cache/n876 ), .CK(clk), .RN(n5866), .Q(\D_cache/cache[0][115] ), .QN(n820) );
  DFFRX1 \D_cache/cache_reg[1][115]  ( .D(\D_cache/n875 ), .CK(clk), .RN(n5866), .Q(\D_cache/cache[1][115] ), .QN(n2383) );
  DFFRX1 \D_cache/cache_reg[2][115]  ( .D(\D_cache/n874 ), .CK(clk), .RN(n5866), .Q(\D_cache/cache[2][115] ), .QN(n1244) );
  DFFRX1 \D_cache/cache_reg[3][115]  ( .D(\D_cache/n873 ), .CK(clk), .RN(n5866), .Q(\D_cache/cache[3][115] ), .QN(n2786) );
  DFFRX1 \D_cache/cache_reg[4][115]  ( .D(\D_cache/n872 ), .CK(clk), .RN(n5871), .Q(\D_cache/cache[4][115] ), .QN(n1211) );
  DFFRX1 \D_cache/cache_reg[5][115]  ( .D(\D_cache/n871 ), .CK(clk), .RN(n5886), .Q(\D_cache/cache[5][115] ), .QN(n2748) );
  DFFRX1 \D_cache/cache_reg[6][115]  ( .D(\D_cache/n870 ), .CK(clk), .RN(n5886), .Q(\D_cache/cache[6][115] ), .QN(n2132) );
  DFFRX1 \D_cache/cache_reg[7][115]  ( .D(\D_cache/n869 ), .CK(clk), .RN(n5886), .Q(\D_cache/cache[7][115] ), .QN(n546) );
  DFFRX1 \D_cache/cache_reg[1][116]  ( .D(\D_cache/n867 ), .CK(clk), .RN(n5885), .Q(\D_cache/cache[1][116] ), .QN(n728) );
  DFFRX1 \D_cache/cache_reg[2][116]  ( .D(\D_cache/n866 ), .CK(clk), .RN(n5885), .Q(\D_cache/cache[2][116] ), .QN(n707) );
  DFFRX1 \D_cache/cache_reg[3][116]  ( .D(\D_cache/n865 ), .CK(clk), .RN(n5885), .Q(\D_cache/cache[3][116] ), .QN(n2275) );
  DFFRX1 \D_cache/cache_reg[4][116]  ( .D(\D_cache/n864 ), .CK(clk), .RN(n5885), .Q(\D_cache/cache[4][116] ), .QN(n1165) );
  DFFRX1 \D_cache/cache_reg[5][116]  ( .D(\D_cache/n863 ), .CK(clk), .RN(n5885), .Q(\D_cache/cache[5][116] ), .QN(n2721) );
  DFFRX1 \D_cache/cache_reg[6][116]  ( .D(\D_cache/n862 ), .CK(clk), .RN(n5885), .Q(\D_cache/cache[6][116] ), .QN(n706) );
  DFFRX1 \D_cache/cache_reg[7][116]  ( .D(\D_cache/n861 ), .CK(clk), .RN(n5885), .Q(\D_cache/cache[7][116] ), .QN(n2274) );
  DFFRX1 \D_cache/cache_reg[1][117]  ( .D(\D_cache/n859 ), .CK(clk), .RN(n5885), .Q(\D_cache/cache[1][117] ), .QN(n1423) );
  DFFRX1 \D_cache/cache_reg[2][117]  ( .D(\D_cache/n858 ), .CK(clk), .RN(n5885), .Q(\D_cache/cache[2][117] ), .QN(n1309) );
  DFFRX1 \D_cache/cache_reg[3][117]  ( .D(\D_cache/n857 ), .CK(clk), .RN(n5885), .Q(\D_cache/cache[3][117] ), .QN(n2838) );
  DFFRX1 \D_cache/cache_reg[4][117]  ( .D(\D_cache/n856 ), .CK(clk), .RN(n5885), .Q(\D_cache/cache[4][117] ), .QN(n1715) );
  DFFRX1 \D_cache/cache_reg[5][117]  ( .D(\D_cache/n855 ), .CK(clk), .RN(n5884), .Q(\D_cache/cache[5][117] ), .QN(n3313) );
  DFFRX1 \D_cache/cache_reg[6][117]  ( .D(\D_cache/n854 ), .CK(clk), .RN(n5884), .Q(\D_cache/cache[6][117] ), .QN(n2729) );
  DFFRX1 \D_cache/cache_reg[7][117]  ( .D(\D_cache/n853 ), .CK(clk), .RN(n5884), .Q(\D_cache/cache[7][117] ), .QN(n1188) );
  DFFRX1 \D_cache/cache_reg[1][118]  ( .D(\D_cache/n851 ), .CK(clk), .RN(n5884), .Q(\D_cache/cache[1][118] ), .QN(n1074) );
  DFFRX1 \D_cache/cache_reg[2][118]  ( .D(\D_cache/n850 ), .CK(clk), .RN(n5884), .Q(\D_cache/cache[2][118] ), .QN(n1111) );
  DFFRX1 \D_cache/cache_reg[3][118]  ( .D(\D_cache/n849 ), .CK(clk), .RN(n5884), .Q(\D_cache/cache[3][118] ), .QN(n2700) );
  DFFRX1 \D_cache/cache_reg[4][118]  ( .D(\D_cache/n848 ), .CK(clk), .RN(n5884), .Q(\D_cache/cache[4][118] ), .QN(n1629) );
  DFFRX1 \D_cache/cache_reg[5][118]  ( .D(\D_cache/n847 ), .CK(clk), .RN(n5884), .Q(\D_cache/cache[5][118] ), .QN(n3205) );
  DFFRX1 \D_cache/cache_reg[6][118]  ( .D(\D_cache/n846 ), .CK(clk), .RN(n5884), .Q(\D_cache/cache[6][118] ), .QN(n714) );
  DFFRX1 \D_cache/cache_reg[7][118]  ( .D(\D_cache/n845 ), .CK(clk), .RN(n5884), .Q(\D_cache/cache[7][118] ), .QN(n2282) );
  DFFRX1 \D_cache/cache_reg[1][119]  ( .D(\D_cache/n843 ), .CK(clk), .RN(n5883), .Q(\D_cache/cache[1][119] ), .QN(n1123) );
  DFFRX1 \D_cache/cache_reg[3][119]  ( .D(\D_cache/n841 ), .CK(clk), .RN(n5883), .Q(\D_cache/cache[3][119] ), .QN(n674) );
  DFFRX1 \D_cache/cache_reg[4][119]  ( .D(\D_cache/n840 ), .CK(clk), .RN(n5883), .Q(\D_cache/cache[4][119] ), .QN(n2089) );
  DFFRX1 \D_cache/cache_reg[5][119]  ( .D(\D_cache/n839 ), .CK(clk), .RN(n5883), .Q(\D_cache/cache[5][119] ), .QN(n502) );
  DFFRX1 \D_cache/cache_reg[6][119]  ( .D(\D_cache/n838 ), .CK(clk), .RN(n5883), .Q(\D_cache/cache[6][119] ), .QN(n2078) );
  DFFRX1 \D_cache/cache_reg[7][119]  ( .D(\D_cache/n837 ), .CK(clk), .RN(n5883), .Q(\D_cache/cache[7][119] ), .QN(n490) );
  DFFRX1 \D_cache/cache_reg[0][120]  ( .D(\D_cache/n836 ), .CK(clk), .RN(n5883), .Q(\D_cache/cache[0][120] ), .QN(n1316) );
  DFFRX1 \D_cache/cache_reg[1][120]  ( .D(\D_cache/n835 ), .CK(clk), .RN(n5883), .Q(\D_cache/cache[1][120] ), .QN(n2845) );
  DFFRX1 \D_cache/cache_reg[2][120]  ( .D(\D_cache/n834 ), .CK(clk), .RN(n5883), .Q(\D_cache/cache[2][120] ), .QN(n1315) );
  DFFRX1 \D_cache/cache_reg[3][120]  ( .D(\D_cache/n833 ), .CK(clk), .RN(n5883), .Q(\D_cache/cache[3][120] ), .QN(n2844) );
  DFFRX1 \D_cache/cache_reg[4][120]  ( .D(\D_cache/n832 ), .CK(clk), .RN(n5883), .Q(\D_cache/cache[4][120] ), .QN(n1371) );
  DFFRX1 \D_cache/cache_reg[5][120]  ( .D(\D_cache/n831 ), .CK(clk), .RN(n5882), .Q(\D_cache/cache[5][120] ), .QN(n2901) );
  DFFRX1 \D_cache/cache_reg[6][120]  ( .D(\D_cache/n830 ), .CK(clk), .RN(n5882), .Q(\D_cache/cache[6][120] ), .QN(n1314) );
  DFFRX1 \D_cache/cache_reg[7][120]  ( .D(\D_cache/n829 ), .CK(clk), .RN(n5882), .Q(\D_cache/cache[7][120] ), .QN(n2843) );
  DFFRX1 \D_cache/cache_reg[1][121]  ( .D(\D_cache/n827 ), .CK(clk), .RN(n5882), .Q(\D_cache/cache[1][121] ), .QN(n1189) );
  DFFRX1 \D_cache/cache_reg[2][121]  ( .D(\D_cache/n826 ), .CK(clk), .RN(n5882), .Q(\D_cache/cache[2][121] ), .QN(n1140) );
  DFFRX1 \D_cache/cache_reg[3][121]  ( .D(\D_cache/n825 ), .CK(clk), .RN(n5882), .Q(\D_cache/cache[3][121] ), .QN(n2702) );
  DFFRX1 \D_cache/cache_reg[4][121]  ( .D(\D_cache/n824 ), .CK(clk), .RN(n5882), .Q(\D_cache/cache[4][121] ), .QN(n2076) );
  DFFRX1 \D_cache/cache_reg[5][121]  ( .D(\D_cache/n823 ), .CK(clk), .RN(n5882), .Q(\D_cache/cache[5][121] ), .QN(n488) );
  DFFRX1 \D_cache/cache_reg[6][121]  ( .D(\D_cache/n822 ), .CK(clk), .RN(n5882), .Q(\D_cache/cache[6][121] ), .QN(n685) );
  DFFRX1 \D_cache/cache_reg[7][121]  ( .D(\D_cache/n821 ), .CK(clk), .RN(n5882), .Q(\D_cache/cache[7][121] ), .QN(n2257) );
  DFFRX1 \D_cache/cache_reg[1][122]  ( .D(\D_cache/n819 ), .CK(clk), .RN(n5881), .Q(\D_cache/cache[1][122] ), .QN(n730) );
  DFFRX1 \D_cache/cache_reg[2][122]  ( .D(\D_cache/n818 ), .CK(clk), .RN(n5881), .Q(\D_cache/cache[2][122] ), .QN(n1109) );
  DFFRX1 \D_cache/cache_reg[3][122]  ( .D(\D_cache/n817 ), .CK(clk), .RN(n5881), .Q(\D_cache/cache[3][122] ), .QN(n2698) );
  DFFRX1 \D_cache/cache_reg[4][122]  ( .D(\D_cache/n816 ), .CK(clk), .RN(n5881), .Q(\D_cache/cache[4][122] ), .QN(n1163) );
  DFFRX1 \D_cache/cache_reg[5][122]  ( .D(\D_cache/n815 ), .CK(clk), .RN(n5881), .Q(\D_cache/cache[5][122] ), .QN(n2719) );
  DFFRX1 \D_cache/cache_reg[6][122]  ( .D(\D_cache/n814 ), .CK(clk), .RN(n5881), .Q(\D_cache/cache[6][122] ), .QN(n712) );
  DFFRX1 \D_cache/cache_reg[7][122]  ( .D(\D_cache/n813 ), .CK(clk), .RN(n5881), .Q(\D_cache/cache[7][122] ), .QN(n2280) );
  DFFRX1 \D_cache/cache_reg[1][123]  ( .D(\D_cache/n811 ), .CK(clk), .RN(n5881), .Q(\D_cache/cache[1][123] ), .QN(n727) );
  DFFRX1 \D_cache/cache_reg[2][123]  ( .D(\D_cache/n810 ), .CK(clk), .RN(n5881), .Q(\D_cache/cache[2][123] ), .QN(n704) );
  DFFRX1 \D_cache/cache_reg[3][123]  ( .D(\D_cache/n809 ), .CK(clk), .RN(n5881), .Q(\D_cache/cache[3][123] ), .QN(n2272) );
  DFFRX1 \D_cache/cache_reg[4][123]  ( .D(\D_cache/n808 ), .CK(clk), .RN(n5880), .Q(\D_cache/cache[4][123] ), .QN(n1149) );
  DFFRX1 \D_cache/cache_reg[5][123]  ( .D(\D_cache/n807 ), .CK(clk), .RN(n5880), .Q(\D_cache/cache[5][123] ), .QN(n2707) );
  DFFRX1 \D_cache/cache_reg[6][123]  ( .D(\D_cache/n806 ), .CK(clk), .RN(n5880), .Q(\D_cache/cache[6][123] ), .QN(n703) );
  DFFRX1 \D_cache/cache_reg[7][123]  ( .D(\D_cache/n805 ), .CK(clk), .RN(n5880), .Q(\D_cache/cache[7][123] ), .QN(n2271) );
  DFFRX1 \D_cache/cache_reg[1][124]  ( .D(\D_cache/n803 ), .CK(clk), .RN(n5880), .Q(\D_cache/cache[1][124] ), .QN(n587) );
  DFFRX1 \D_cache/cache_reg[2][124]  ( .D(\D_cache/n802 ), .CK(clk), .RN(n5880), .Q(\D_cache/cache[2][124] ), .QN(n1345) );
  DFFRX1 \D_cache/cache_reg[3][124]  ( .D(\D_cache/n801 ), .CK(clk), .RN(n5880), .Q(\D_cache/cache[3][124] ), .QN(n2874) );
  DFFRX1 \D_cache/cache_reg[4][124]  ( .D(\D_cache/n800 ), .CK(clk), .RN(n5880), .Q(\D_cache/cache[4][124] ), .QN(n1368) );
  DFFRX1 \D_cache/cache_reg[5][124]  ( .D(\D_cache/n799 ), .CK(clk), .RN(n5880), .Q(\D_cache/cache[5][124] ), .QN(n2898) );
  DFFRX1 \D_cache/cache_reg[6][124]  ( .D(\D_cache/n798 ), .CK(clk), .RN(n5880), .Q(\D_cache/cache[6][124] ), .QN(n2086) );
  DFFRX1 \D_cache/cache_reg[7][124]  ( .D(\D_cache/n797 ), .CK(clk), .RN(n5880), .Q(\D_cache/cache[7][124] ), .QN(n498) );
  DFFRX1 \D_cache/cache_reg[0][125]  ( .D(\D_cache/n796 ), .CK(clk), .RN(n5879), .Q(\D_cache/cache[0][125] ), .QN(n825) );
  DFFRX1 \D_cache/cache_reg[1][125]  ( .D(\D_cache/n795 ), .CK(clk), .RN(n5879), .Q(\D_cache/cache[1][125] ), .QN(n2388) );
  DFFRX1 \D_cache/cache_reg[2][125]  ( .D(\D_cache/n794 ), .CK(clk), .RN(n5879), .Q(\D_cache/cache[2][125] ), .QN(n1247) );
  DFFRX1 \D_cache/cache_reg[3][125]  ( .D(\D_cache/n793 ), .CK(clk), .RN(n5879), .Q(\D_cache/cache[3][125] ), .QN(n2789) );
  DFFRX1 \D_cache/cache_reg[4][125]  ( .D(\D_cache/n792 ), .CK(clk), .RN(n5879), .Q(\D_cache/cache[4][125] ), .QN(n1378) );
  DFFRX1 \D_cache/cache_reg[5][125]  ( .D(\D_cache/n791 ), .CK(clk), .RN(n5879), .Q(\D_cache/cache[5][125] ), .QN(n2908) );
  DFFRX1 \D_cache/cache_reg[6][125]  ( .D(\D_cache/n790 ), .CK(clk), .RN(n5879), .Q(\D_cache/cache[6][125] ), .QN(n824) );
  DFFRX1 \D_cache/cache_reg[7][125]  ( .D(\D_cache/n789 ), .CK(clk), .RN(n5879), .Q(\D_cache/cache[7][125] ), .QN(n2387) );
  DFFRX1 \D_cache/cache_reg[1][126]  ( .D(\D_cache/n787 ), .CK(clk), .RN(n5879), .Q(\D_cache/cache[1][126] ), .QN(n1204) );
  DFFRX1 \D_cache/cache_reg[2][126]  ( .D(\D_cache/n786 ), .CK(clk), .RN(n5879), .Q(\D_cache/cache[2][126] ), .QN(n1177) );
  DFFRX1 \D_cache/cache_reg[3][126]  ( .D(\D_cache/n785 ), .CK(clk), .RN(n5879), .Q(\D_cache/cache[3][126] ), .QN(n2727) );
  DFFRX1 \D_cache/cache_reg[4][126]  ( .D(\D_cache/n784 ), .CK(clk), .RN(n5878), .Q(\D_cache/cache[4][126] ), .QN(n1632) );
  DFFRX1 \D_cache/cache_reg[5][126]  ( .D(\D_cache/n783 ), .CK(clk), .RN(n5878), .Q(\D_cache/cache[5][126] ), .QN(n3208) );
  DFFRX1 \D_cache/cache_reg[6][126]  ( .D(\D_cache/n782 ), .CK(clk), .RN(n5878), .Q(\D_cache/cache[6][126] ), .QN(n1141) );
  DFFRX1 \D_cache/cache_reg[7][126]  ( .D(\D_cache/n781 ), .CK(clk), .RN(n5878), .Q(\D_cache/cache[7][126] ), .QN(n2703) );
  DFFRX1 \D_cache/cache_reg[0][127]  ( .D(\D_cache/n780 ), .CK(clk), .RN(n5878), .Q(\D_cache/cache[0][127] ), .QN(n1393) );
  DFFRX1 \D_cache/cache_reg[1][127]  ( .D(\D_cache/n779 ), .CK(clk), .RN(n5878), .Q(\D_cache/cache[1][127] ), .QN(n2923) );
  DFFRX1 \D_cache/cache_reg[2][127]  ( .D(\D_cache/n778 ), .CK(clk), .RN(n5878), .Q(\D_cache/cache[2][127] ), .QN(n1246) );
  DFFRX1 \D_cache/cache_reg[3][127]  ( .D(\D_cache/n777 ), .CK(clk), .RN(n5878), .Q(\D_cache/cache[3][127] ), .QN(n2788) );
  DFFRX1 \D_cache/cache_reg[4][127]  ( .D(\D_cache/n776 ), .CK(clk), .RN(n5878), .Q(\D_cache/cache[4][127] ), .QN(n1720) );
  DFFRX1 \D_cache/cache_reg[5][127]  ( .D(\D_cache/n775 ), .CK(clk), .RN(n5878), .Q(\D_cache/cache[5][127] ), .QN(n3318) );
  DFFRX1 \D_cache/cache_reg[6][127]  ( .D(\D_cache/n774 ), .CK(clk), .RN(n5878), .Q(\D_cache/cache[6][127] ), .QN(n823) );
  DFFRX1 \D_cache/cache_reg[7][127]  ( .D(\D_cache/n773 ), .CK(clk), .RN(n5878), .Q(\D_cache/cache[7][127] ), .QN(n2386) );
  DFFRX1 \D_cache/cache_reg[0][128]  ( .D(\D_cache/n772 ), .CK(clk), .RN(n5877), .Q(\D_cache/cache[0][128] ), .QN(n3029) );
  DFFRX1 \D_cache/cache_reg[1][128]  ( .D(\D_cache/n771 ), .CK(clk), .RN(n5877), .Q(\D_cache/cache[1][128] ), .QN(n848) );
  DFFRX1 \D_cache/cache_reg[2][128]  ( .D(\D_cache/n770 ), .CK(clk), .RN(n5877), .Q(\D_cache/cache[2][128] ), .QN(n3215) );
  DFFRX1 \D_cache/cache_reg[3][128]  ( .D(\D_cache/n769 ), .CK(clk), .RN(n5877), .Q(\D_cache/cache[3][128] ), .QN(n1291) );
  DFFRX1 \D_cache/cache_reg[4][128]  ( .D(\D_cache/n768 ), .CK(clk), .RN(n5877), .Q(\D_cache/cache[4][128] ), .QN(n1460) );
  DFFRX1 \D_cache/cache_reg[5][128]  ( .D(\D_cache/n767 ), .CK(clk), .RN(n5877), .Q(\D_cache/cache[5][128] ), .QN(n3034) );
  DFFRX1 \D_cache/cache_reg[6][128]  ( .D(\D_cache/n766 ), .CK(clk), .RN(n5877), .Q(\D_cache/cache[6][128] ), .QN(n751) );
  DFFRX1 \D_cache/cache_reg[0][130]  ( .D(\D_cache/n756 ), .CK(clk), .RN(n5876), .Q(\D_cache/cache[0][130] ), .QN(n2208) );
  DFFRX1 \D_cache/cache_reg[1][130]  ( .D(\D_cache/n755 ), .CK(clk), .RN(n5876), .Q(\D_cache/cache[1][130] ), .QN(n2018) );
  DFFRX1 \D_cache/cache_reg[2][130]  ( .D(\D_cache/n754 ), .CK(clk), .RN(n5876), .Q(\D_cache/cache[2][130] ), .QN(n511) );
  DFFRX1 \D_cache/cache_reg[3][130]  ( .D(\D_cache/n753 ), .CK(clk), .RN(n5876), .Q(\D_cache/cache[3][130] ), .QN(n2098) );
  DFFRX1 \D_cache/cache_reg[4][130]  ( .D(\D_cache/n752 ), .CK(clk), .RN(n5881), .Q(\D_cache/cache[4][130] ), .QN(n2165) );
  DFFRX1 \D_cache/cache_reg[5][130]  ( .D(\D_cache/n751 ), .CK(clk), .RN(n5886), .Q(\D_cache/cache[5][130] ), .QN(n591) );
  DFFRX1 \D_cache/cache_reg[6][130]  ( .D(\D_cache/n750 ), .CK(clk), .RN(n5936), .Q(\D_cache/cache[6][130] ), .QN(n2124) );
  DFFRX1 \D_cache/cache_reg[0][131]  ( .D(\D_cache/n748 ), .CK(clk), .RN(n5936), .Q(\D_cache/cache[0][131] ), .QN(n2112) );
  DFFRX1 \D_cache/cache_reg[1][131]  ( .D(\D_cache/n747 ), .CK(clk), .RN(n5936), .Q(\D_cache/cache[1][131] ), .QN(n525) );
  DFFRX1 \D_cache/cache_reg[2][131]  ( .D(\D_cache/n746 ), .CK(clk), .RN(n5936), .Q(\D_cache/cache[2][131] ), .QN(n2113) );
  DFFRX1 \D_cache/cache_reg[3][131]  ( .D(\D_cache/n745 ), .CK(clk), .RN(n5935), .Q(\D_cache/cache[3][131] ), .QN(n526) );
  DFFRX1 \D_cache/cache_reg[4][131]  ( .D(\D_cache/n744 ), .CK(clk), .RN(n5935), .Q(\D_cache/cache[4][131] ), .QN(n2146) );
  DFFRX1 \D_cache/cache_reg[6][131]  ( .D(\D_cache/n742 ), .CK(clk), .RN(n5935), .Q(\D_cache/cache[6][131] ), .QN(n2125) );
  DFFRX1 \D_cache/cache_reg[0][133]  ( .D(\D_cache/n732 ), .CK(clk), .RN(n5934), .Q(\D_cache/cache[0][133] ), .QN(n631) );
  DFFRX1 \D_cache/cache_reg[2][133]  ( .D(\D_cache/n730 ), .CK(clk), .RN(n5934), .Q(\D_cache/cache[2][133] ), .QN(n632) );
  DFFRX1 \D_cache/cache_reg[0][134]  ( .D(\D_cache/n724 ), .CK(clk), .RN(n5934), .Q(\D_cache/cache[0][134] ), .QN(n633) );
  DFFRX1 \D_cache/cache_reg[0][136]  ( .D(\D_cache/n708 ), .CK(clk), .RN(n5932), .Q(\D_cache/cache[0][136] ), .QN(n3005) );
  DFFRX1 \D_cache/cache_reg[1][136]  ( .D(\D_cache/n707 ), .CK(clk), .RN(n5932), .Q(\D_cache/cache[1][136] ), .QN(n577) );
  DFFRX1 \D_cache/cache_reg[2][136]  ( .D(\D_cache/n706 ), .CK(clk), .RN(n5932), .Q(\D_cache/cache[2][136] ), .QN(n3008) );
  DFFRX1 \D_cache/cache_reg[3][136]  ( .D(\D_cache/n705 ), .CK(clk), .RN(n5932), .Q(\D_cache/cache[3][136] ), .QN(n584) );
  DFFRX1 \D_cache/cache_reg[4][136]  ( .D(\D_cache/n704 ), .CK(clk), .RN(n5932), .Q(\D_cache/cache[4][136] ), .QN(n2999) );
  DFFRX1 \D_cache/cache_reg[5][136]  ( .D(\D_cache/n703 ), .CK(clk), .RN(n5932), .Q(\D_cache/cache[5][136] ), .QN(n557) );
  DFFRX1 \D_cache/cache_reg[6][136]  ( .D(\D_cache/n702 ), .CK(clk), .RN(n5932), .Q(\D_cache/cache[6][136] ), .QN(n756) );
  DFFRX1 \D_cache/cache_reg[7][136]  ( .D(\D_cache/n701 ), .CK(clk), .RN(n5932), .Q(\D_cache/cache[7][136] ), .QN(n2317) );
  DFFRX1 \D_cache/cache_reg[0][138]  ( .D(\D_cache/n692 ), .CK(clk), .RN(n5931), .Q(\D_cache/cache[0][138] ), .QN(n634) );
  DFFRX1 \D_cache/cache_reg[0][140]  ( .D(\D_cache/n676 ), .CK(clk), .RN(n5930), .Q(\D_cache/cache[0][140] ) );
  DFFRX1 \D_cache/cache_reg[4][140]  ( .D(\D_cache/n672 ), .CK(clk), .RN(n5929), .Q(\D_cache/cache[4][140] ), .QN(n3014) );
  DFFRX1 \D_cache/cache_reg[5][140]  ( .D(\D_cache/n671 ), .CK(clk), .RN(n5929), .Q(\D_cache/cache[5][140] ), .QN(n2222) );
  DFFRX1 \D_cache/cache_reg[0][141]  ( .D(\D_cache/n668 ), .CK(clk), .RN(n5929), .Q(\D_cache/cache[0][141] ), .QN(n2987) );
  DFFRX1 \D_cache/cache_reg[1][141]  ( .D(\D_cache/n667 ), .CK(clk), .RN(n5929), .Q(\D_cache/cache[1][141] ), .QN(n540) );
  DFFRX1 \D_cache/cache_reg[2][141]  ( .D(\D_cache/n666 ), .CK(clk), .RN(n5929), .Q(\D_cache/cache[2][141] ), .QN(n2652) );
  DFFRX1 \D_cache/cache_reg[3][141]  ( .D(\D_cache/n665 ), .CK(clk), .RN(n5929), .Q(\D_cache/cache[3][141] ), .QN(n590) );
  DFFRX1 \D_cache/cache_reg[4][141]  ( .D(\D_cache/n664 ), .CK(clk), .RN(n5929), .Q(\D_cache/cache[4][141] ), .QN(n1771) );
  DFFRX1 \D_cache/cache_reg[5][141]  ( .D(\D_cache/n663 ), .CK(clk), .RN(n5929), .Q(\D_cache/cache[5][141] ), .QN(n3401) );
  DFFRX1 \D_cache/cache_reg[6][141]  ( .D(\D_cache/n662 ), .CK(clk), .RN(n5928), .Q(\D_cache/cache[6][141] ), .QN(n635) );
  DFFRX1 \D_cache/cache_reg[0][143]  ( .D(\D_cache/n652 ), .CK(clk), .RN(n5928), .Q(\D_cache/cache[0][143] ), .QN(n3028) );
  DFFRX1 \D_cache/cache_reg[1][143]  ( .D(\D_cache/n651 ), .CK(clk), .RN(n5928), .Q(\D_cache/cache[1][143] ), .QN(n846) );
  DFFRX1 \D_cache/cache_reg[2][143]  ( .D(\D_cache/n650 ), .CK(clk), .RN(n5927), .Q(\D_cache/cache[2][143] ), .QN(n2996) );
  DFFRX1 \D_cache/cache_reg[3][143]  ( .D(\D_cache/n649 ), .CK(clk), .RN(n5927), .Q(\D_cache/cache[3][143] ), .QN(n554) );
  DFFRX1 \D_cache/cache_reg[4][143]  ( .D(\D_cache/n648 ), .CK(clk), .RN(n5927), .Q(\D_cache/cache[4][143] ), .QN(n1772) );
  DFFRX1 \D_cache/cache_reg[6][143]  ( .D(\D_cache/n646 ), .CK(clk), .RN(n5927), .Q(\D_cache/cache[6][143] ), .QN(n636) );
  DFFRX1 \D_cache/cache_reg[0][145]  ( .D(\D_cache/n636 ), .CK(clk), .RN(n5926), .Q(\D_cache/cache[0][145] ), .QN(n2019) );
  DFFRX1 \D_cache/cache_reg[2][145]  ( .D(\D_cache/n634 ), .CK(clk), .RN(n5926), .Q(\D_cache/cache[2][145] ), .QN(n2164) );
  DFFRX1 \D_cache/cache_reg[0][146]  ( .D(\D_cache/n628 ), .CK(clk), .RN(n5954), .Q(\D_cache/cache[0][146] ), .QN(n2155) );
  DFFRX1 \D_cache/cache_reg[2][146]  ( .D(\D_cache/n626 ), .CK(clk), .RN(n5945), .Q(\D_cache/cache[2][146] ), .QN(n768) );
  DFFRX1 \D_cache/cache_reg[0][147]  ( .D(\D_cache/n620 ), .CK(clk), .RN(n5945), .Q(\D_cache/cache[0][147] ), .QN(n3003) );
  DFFRX1 \D_cache/cache_reg[1][147]  ( .D(\D_cache/n619 ), .CK(clk), .RN(n5945), .Q(\D_cache/cache[1][147] ), .QN(n570) );
  DFFRX1 \D_cache/cache_reg[2][147]  ( .D(\D_cache/n618 ), .CK(clk), .RN(n5944), .Q(\D_cache/cache[2][147] ), .QN(n2998) );
  DFFRX1 \D_cache/cache_reg[3][147]  ( .D(\D_cache/n617 ), .CK(clk), .RN(n5945), .Q(\D_cache/cache[3][147] ), .QN(n556) );
  DFFRX1 \D_cache/cache_reg[4][147]  ( .D(\D_cache/n616 ), .CK(clk), .RN(n5945), .Q(\D_cache/cache[4][147] ), .QN(n3320) );
  DFFRX1 \D_cache/cache_reg[5][147]  ( .D(\D_cache/n615 ), .CK(clk), .RN(n5945), .Q(\D_cache/cache[5][147] ) );
  DFFRX1 \D_cache/cache_reg[6][147]  ( .D(\D_cache/n614 ), .CK(clk), .RN(n5944), .Q(\D_cache/cache[6][147] ), .QN(n1392) );
  DFFRX1 \D_cache/cache_reg[7][147]  ( .D(\D_cache/n613 ), .CK(clk), .RN(n5944), .Q(\D_cache/cache[7][147] ), .QN(n2922) );
  DFFRX1 \D_cache/cache_reg[0][149]  ( .D(\D_cache/n604 ), .CK(clk), .RN(n5944), .Q(\D_cache/cache[0][149] ), .QN(n3265) );
  DFFRX1 \D_cache/cache_reg[1][149]  ( .D(\D_cache/n603 ), .CK(clk), .RN(n5943), .Q(\D_cache/cache[1][149] ), .QN(n1425) );
  DFFRX1 \D_cache/cache_reg[2][149]  ( .D(\D_cache/n602 ), .CK(clk), .RN(n5943), .Q(\D_cache/cache[2][149] ), .QN(n2997) );
  DFFRX1 \D_cache/cache_reg[3][149]  ( .D(\D_cache/n601 ), .CK(clk), .RN(n5943), .Q(\D_cache/cache[3][149] ), .QN(n555) );
  DFFRX1 \D_cache/cache_reg[4][149]  ( .D(\D_cache/n600 ), .CK(clk), .RN(n5943), .Q(\D_cache/cache[4][149] ), .QN(n1773) );
  DFFRX1 \D_cache/cache_reg[5][149]  ( .D(\D_cache/n599 ), .CK(clk), .RN(n5943), .Q(\D_cache/cache[5][149] ), .QN(n3404) );
  DFFRX1 \D_cache/cache_reg[6][149]  ( .D(\D_cache/n598 ), .CK(clk), .RN(n5943), .Q(\D_cache/cache[6][149] ), .QN(n1391) );
  DFFRX1 \D_cache/cache_reg[7][149]  ( .D(\D_cache/n597 ), .CK(clk), .RN(n5943), .Q(\D_cache/cache[7][149] ), .QN(n2921) );
  DFFRX1 \D_cache/cache_reg[0][150]  ( .D(\D_cache/n596 ), .CK(clk), .RN(n5943), .Q(\D_cache/cache[0][150] ), .QN(n2127) );
  DFFRX1 \D_cache/cache_reg[1][150]  ( .D(\D_cache/n595 ), .CK(clk), .RN(n5943), .Q(\D_cache/cache[1][150] ), .QN(n541) );
  DFFRX1 \D_cache/cache_reg[2][150]  ( .D(\D_cache/n594 ), .CK(clk), .RN(n5943), .Q(\D_cache/cache[2][150] ), .QN(n2138) );
  DFFRX1 \D_cache/cache_reg[3][150]  ( .D(\D_cache/n593 ), .CK(clk), .RN(n5942), .Q(\D_cache/cache[3][150] ), .QN(n553) );
  DFFRX1 \D_cache/cache_reg[4][150]  ( .D(\D_cache/n592 ), .CK(clk), .RN(n5943), .Q(\D_cache/cache[4][150] ), .QN(n1469) );
  DFFRX1 \D_cache/cache_reg[6][150]  ( .D(\D_cache/n590 ), .CK(clk), .RN(n5942), .Q(\D_cache/cache[6][150] ), .QN(n2951) );
  DFFRX1 \D_cache/cache_reg[0][151]  ( .D(\D_cache/n588 ), .CK(clk), .RN(n5942), .Q(\D_cache/cache[0][151] ), .QN(n3004) );
  DFFRX1 \D_cache/cache_reg[1][151]  ( .D(\D_cache/n587 ), .CK(clk), .RN(n5942), .Q(\D_cache/cache[1][151] ), .QN(n576) );
  DFFRX1 \D_cache/cache_reg[2][151]  ( .D(\D_cache/n586 ), .CK(clk), .RN(n5942), .Q(\D_cache/cache[2][151] ), .QN(n3007) );
  DFFRX1 \D_cache/cache_reg[3][151]  ( .D(\D_cache/n585 ), .CK(clk), .RN(n5942), .Q(\D_cache/cache[3][151] ), .QN(n583) );
  DFFRX1 \D_cache/cache_reg[4][151]  ( .D(\D_cache/n584 ), .CK(clk), .RN(n5942), .Q(\D_cache/cache[4][151] ), .QN(n3000) );
  DFFRX1 \D_cache/cache_reg[5][151]  ( .D(\D_cache/n583 ), .CK(clk), .RN(n5942), .Q(\D_cache/cache[5][151] ), .QN(n558) );
  DFFRX1 \D_cache/cache_reg[6][151]  ( .D(\D_cache/n582 ), .CK(clk), .RN(n5942), .Q(\D_cache/cache[6][151] ), .QN(n628) );
  DFFRX1 \D_cache/cache_reg[0][152]  ( .D(\D_cache/n580 ), .CK(clk), .RN(n5942), .Q(\D_cache/cache[0][152] ), .QN(n3346) );
  DFFRX1 \D_cache/cache_reg[0][153]  ( .D(\D_cache/n572 ), .CK(clk), .RN(n5941), .Q(\D_cache/cache[0][153] ), .QN(n1485) );
  DFFRX1 \D_cache/cache_reg[1][153]  ( .D(\D_cache/n571 ), .CK(clk), .RN(n5941), .Q(\D_cache/cache[1][153] ), .QN(n3068) );
  DFFRX1 \D_cache/cache_reg[2][153]  ( .D(\D_cache/n570 ), .CK(clk), .RN(n5941), .Q(\D_cache/cache[2][153] ), .QN(n1594) );
  DFFRX1 \D_cache/cache_reg[3][153]  ( .D(\D_cache/n569 ), .CK(clk), .RN(n5941), .Q(\D_cache/cache[3][153] ), .QN(n3171) );
  DFFRX1 \D_cache/cache_reg[4][153]  ( .D(\D_cache/n568 ), .CK(clk), .RN(n5940), .Q(\D_cache/cache[4][153] ), .QN(n3328) );
  DFFRX1 \D_cache/cache_reg[5][153]  ( .D(\D_cache/n567 ), .CK(clk), .RN(n5940), .Q(\D_cache/cache[5][153] ), .QN(n1726) );
  DFFRX1 \D_cache/cache_reg[6][153]  ( .D(\D_cache/n566 ), .CK(clk), .RN(n5940), .Q(\D_cache/cache[6][153] ), .QN(n2744) );
  DFFRX1 \D_cache/cache_reg[7][153]  ( .D(\D_cache/n565 ), .CK(clk), .RN(n5940), .Q(\D_cache/cache[7][153] ), .QN(n1284) );
  DFFRX1 \D_cache/cache_reg[7][128]  ( .D(\D_cache/n765 ), .CK(clk), .RN(n5940), .Q(\D_cache/cache[7][128] ), .QN(n2312) );
  DFFRX1 \I_cache/cache_reg[0][0]  ( .D(n12786), .CK(clk), .RN(n5939), .Q(
        \I_cache/cache[0][0] ), .QN(n1677) );
  DFFRX1 \I_cache/cache_reg[1][0]  ( .D(n12785), .CK(clk), .RN(n5939), .Q(
        \I_cache/cache[1][0] ), .QN(n3267) );
  DFFRX1 \I_cache/cache_reg[2][0]  ( .D(n12784), .CK(clk), .RN(n5939), .Q(
        \I_cache/cache[2][0] ), .QN(n1679) );
  DFFRX1 \I_cache/cache_reg[3][0]  ( .D(n12783), .CK(clk), .RN(n5939), .Q(
        \I_cache/cache[3][0] ), .QN(n3269) );
  DFFRX1 \I_cache/cache_reg[4][0]  ( .D(n12782), .CK(clk), .RN(n5939), .Q(
        \I_cache/cache[4][0] ), .QN(n1678) );
  DFFRX1 \I_cache/cache_reg[5][0]  ( .D(n12781), .CK(clk), .RN(n5939), .Q(
        \I_cache/cache[5][0] ), .QN(n3268) );
  DFFRX1 \I_cache/cache_reg[6][0]  ( .D(n12780), .CK(clk), .RN(n5939), .Q(
        \I_cache/cache[6][0] ), .QN(n3002) );
  DFFRX1 \I_cache/cache_reg[7][0]  ( .D(n12787), .CK(clk), .RN(n5939), .Q(
        \I_cache/cache[7][0] ), .QN(n1439) );
  DFFRX1 \I_cache/cache_reg[0][1]  ( .D(n12779), .CK(clk), .RN(n5939), .Q(
        \I_cache/cache[0][1] ), .QN(n1709) );
  DFFRX1 \I_cache/cache_reg[1][1]  ( .D(n12778), .CK(clk), .RN(n5939), .Q(
        \I_cache/cache[1][1] ), .QN(n3306) );
  DFFRX1 \I_cache/cache_reg[2][1]  ( .D(n12777), .CK(clk), .RN(n5939), .Q(
        \I_cache/cache[2][1] ), .QN(n1680) );
  DFFRX1 \I_cache/cache_reg[3][1]  ( .D(n12776), .CK(clk), .RN(n5938), .Q(
        \I_cache/cache[3][1] ), .QN(n3271) );
  DFFRX1 \I_cache/cache_reg[4][1]  ( .D(n12775), .CK(clk), .RN(n5938), .Q(
        \I_cache/cache[4][1] ), .QN(n2994) );
  DFFRX1 \I_cache/cache_reg[5][1]  ( .D(n12774), .CK(clk), .RN(n5938), .Q(
        \I_cache/cache[5][1] ), .QN(n1436) );
  DFFRX1 \I_cache/cache_reg[6][1]  ( .D(n12773), .CK(clk), .RN(n5938), .Q(
        \I_cache/cache[6][1] ), .QN(n1713) );
  DFFRX1 \I_cache/cache_reg[7][1]  ( .D(n12772), .CK(clk), .RN(n5938), .Q(
        \I_cache/cache[7][1] ), .QN(n3310) );
  DFFRX1 \I_cache/cache_reg[0][2]  ( .D(n12771), .CK(clk), .RN(n5938), .Q(
        \I_cache/cache[0][2] ), .QN(n1617) );
  DFFRX1 \I_cache/cache_reg[1][2]  ( .D(n12770), .CK(clk), .RN(n5938), .Q(
        \I_cache/cache[1][2] ), .QN(n3194) );
  DFFRX1 \I_cache/cache_reg[2][2]  ( .D(n12769), .CK(clk), .RN(n5938), .Q(
        \I_cache/cache[2][2] ), .QN(n1577) );
  DFFRX1 \I_cache/cache_reg[3][2]  ( .D(n12768), .CK(clk), .RN(n5938), .Q(
        \I_cache/cache[3][2] ), .QN(n3159) );
  DFFRX1 \I_cache/cache_reg[4][2]  ( .D(n12767), .CK(clk), .RN(n5938), .Q(
        \I_cache/cache[4][2] ), .QN(n1286) );
  DFFRX1 \I_cache/cache_reg[5][2]  ( .D(n12766), .CK(clk), .RN(n5938), .Q(
        \I_cache/cache[5][2] ), .QN(n2982) );
  DFFRX1 \I_cache/cache_reg[6][2]  ( .D(n12765), .CK(clk), .RN(n5938), .Q(
        \I_cache/cache[6][2] ), .QN(n1625) );
  DFFRX1 \I_cache/cache_reg[7][2]  ( .D(n12764), .CK(clk), .RN(n5937), .Q(
        \I_cache/cache[7][2] ), .QN(n3311) );
  DFFRX1 \I_cache/cache_reg[0][3]  ( .D(n12763), .CK(clk), .RN(n5937), .Q(
        \I_cache/cache[0][3] ), .QN(n1683) );
  DFFRX1 \I_cache/cache_reg[1][3]  ( .D(n12762), .CK(clk), .RN(n5937), .Q(
        \I_cache/cache[1][3] ), .QN(n3274) );
  DFFRX1 \I_cache/cache_reg[2][3]  ( .D(n12761), .CK(clk), .RN(n5937), .Q(
        \I_cache/cache[2][3] ), .QN(n1669) );
  DFFRX1 \I_cache/cache_reg[3][3]  ( .D(n12760), .CK(clk), .RN(n5937), .Q(
        \I_cache/cache[3][3] ), .QN(n3253) );
  DFFRX1 \I_cache/cache_reg[4][3]  ( .D(n12759), .CK(clk), .RN(n5937), .Q(
        \I_cache/cache[4][3] ), .QN(n1668) );
  DFFRX1 \I_cache/cache_reg[5][3]  ( .D(n12758), .CK(clk), .RN(n5937), .Q(
        \I_cache/cache[5][3] ), .QN(n3252) );
  DFFRX1 \I_cache/cache_reg[6][3]  ( .D(n12757), .CK(clk), .RN(n5937), .Q(
        \I_cache/cache[6][3] ), .QN(n769) );
  DFFRX1 \I_cache/cache_reg[7][3]  ( .D(n12756), .CK(clk), .RN(n5937), .Q(
        \I_cache/cache[7][3] ), .QN(n2331) );
  DFFRX1 \I_cache/cache_reg[0][4]  ( .D(n12755), .CK(clk), .RN(n5937), .Q(
        \I_cache/cache[0][4] ), .QN(n1710) );
  DFFRX1 \I_cache/cache_reg[1][4]  ( .D(n12754), .CK(clk), .RN(n5937), .Q(
        \I_cache/cache[1][4] ), .QN(n3307) );
  DFFRX1 \I_cache/cache_reg[2][4]  ( .D(n12753), .CK(clk), .RN(n5937), .Q(
        \I_cache/cache[2][4] ), .QN(n1681) );
  DFFRX1 \I_cache/cache_reg[3][4]  ( .D(n12752), .CK(clk), .RN(n5936), .Q(
        \I_cache/cache[3][4] ), .QN(n3272) );
  DFFRX1 \I_cache/cache_reg[4][4]  ( .D(n12751), .CK(clk), .RN(n5936), .Q(
        \I_cache/cache[4][4] ), .QN(n2995) );
  DFFRX1 \I_cache/cache_reg[5][4]  ( .D(n12750), .CK(clk), .RN(n5936), .Q(
        \I_cache/cache[5][4] ), .QN(n1437) );
  DFFRX1 \I_cache/cache_reg[6][4]  ( .D(n12749), .CK(clk), .RN(n5936), .Q(
        \I_cache/cache[6][4] ), .QN(n1714) );
  DFFRX1 \I_cache/cache_reg[7][4]  ( .D(n12748), .CK(clk), .RN(n5936), .Q(
        \I_cache/cache[7][4] ), .QN(n3312) );
  DFFRX1 \I_cache/cache_reg[0][5]  ( .D(n12747), .CK(clk), .RN(n5936), .Q(
        \I_cache/cache[0][5] ), .QN(n2742) );
  DFFRX1 \I_cache/cache_reg[1][5]  ( .D(n12746), .CK(clk), .RN(n5936), .Q(
        \I_cache/cache[1][5] ), .QN(n1282) );
  DFFRX1 \I_cache/cache_reg[2][5]  ( .D(n12745), .CK(clk), .RN(n5941), .Q(
        \I_cache/cache[2][5] ), .QN(n1508) );
  DFFRX1 \I_cache/cache_reg[3][5]  ( .D(n12744), .CK(clk), .RN(n5916), .Q(
        \I_cache/cache[3][5] ), .QN(n3088) );
  DFFRX1 \I_cache/cache_reg[4][5]  ( .D(n12743), .CK(clk), .RN(n5916), .Q(
        \I_cache/cache[4][5] ), .QN(n1507) );
  DFFRX1 \I_cache/cache_reg[5][5]  ( .D(n12742), .CK(clk), .RN(n5916), .Q(
        \I_cache/cache[5][5] ), .QN(n3087) );
  DFFRX1 \I_cache/cache_reg[6][5]  ( .D(n12741), .CK(clk), .RN(n5916), .Q(
        \I_cache/cache[6][5] ), .QN(n1488) );
  DFFRX1 \I_cache/cache_reg[7][5]  ( .D(n12740), .CK(clk), .RN(n5916), .Q(
        \I_cache/cache[7][5] ), .QN(n3072) );
  DFFRX1 \I_cache/cache_reg[0][6]  ( .D(n12739), .CK(clk), .RN(n5915), .Q(
        \I_cache/cache[0][6] ), .QN(n1651) );
  DFFRX1 \I_cache/cache_reg[1][6]  ( .D(n12738), .CK(clk), .RN(n5915), .Q(
        \I_cache/cache[1][6] ), .QN(n3233) );
  DFFRX1 \I_cache/cache_reg[2][6]  ( .D(n12737), .CK(clk), .RN(n5915), .Q(
        \I_cache/cache[2][6] ), .QN(n1652) );
  DFFRX1 \I_cache/cache_reg[3][6]  ( .D(n12736), .CK(clk), .RN(n5915), .Q(
        \I_cache/cache[3][6] ), .QN(n3234) );
  DFFRX1 \I_cache/cache_reg[4][6]  ( .D(n12735), .CK(clk), .RN(n5915), .Q(
        \I_cache/cache[4][6] ), .QN(n3216) );
  DFFRX1 \I_cache/cache_reg[5][6]  ( .D(n12734), .CK(clk), .RN(n5915), .Q(
        \I_cache/cache[5][6] ), .QN(n1419) );
  DFFRX1 \I_cache/cache_reg[6][6]  ( .D(n12733), .CK(clk), .RN(n5915), .Q(
        \I_cache/cache[6][6] ), .QN(n1689) );
  DFFRX1 \I_cache/cache_reg[7][6]  ( .D(n12732), .CK(clk), .RN(n5915), .Q(
        \I_cache/cache[7][6] ), .QN(n3284) );
  DFFRX1 \I_cache/cache_reg[0][7]  ( .D(n12731), .CK(clk), .RN(n5915), .Q(
        \I_cache/cache[0][7] ), .QN(n1478) );
  DFFRX1 \I_cache/cache_reg[1][7]  ( .D(n12730), .CK(clk), .RN(n5915), .Q(
        \I_cache/cache[1][7] ), .QN(n3052) );
  DFFRX1 \I_cache/cache_reg[2][7]  ( .D(n12729), .CK(clk), .RN(n5915), .Q(
        \I_cache/cache[2][7] ), .QN(n3009) );
  DFFRX1 \I_cache/cache_reg[3][7]  ( .D(n12728), .CK(clk), .RN(n5915), .Q(
        \I_cache/cache[3][7] ), .QN(n1441) );
  DFFRX1 \I_cache/cache_reg[4][7]  ( .D(n12727), .CK(clk), .RN(n5914), .Q(
        \I_cache/cache[4][7] ), .QN(n3030) );
  DFFRX1 \I_cache/cache_reg[5][7]  ( .D(n12726), .CK(clk), .RN(n5914), .Q(
        \I_cache/cache[5][7] ), .QN(n850) );
  DFFRX1 \I_cache/cache_reg[6][7]  ( .D(n12725), .CK(clk), .RN(n5914), .Q(
        \I_cache/cache[6][7] ), .QN(n1479) );
  DFFRX1 \I_cache/cache_reg[7][7]  ( .D(n12724), .CK(clk), .RN(n5914), .Q(
        \I_cache/cache[7][7] ), .QN(n3053) );
  DFFRX1 \I_cache/cache_reg[0][8]  ( .D(n12723), .CK(clk), .RN(n5914), .Q(
        \I_cache/cache[0][8] ), .QN(n1593) );
  DFFRX1 \I_cache/cache_reg[1][8]  ( .D(n12722), .CK(clk), .RN(n5914), .Q(
        \I_cache/cache[1][8] ), .QN(n3303) );
  DFFRX1 \I_cache/cache_reg[2][8]  ( .D(n12721), .CK(clk), .RN(n5914), .Q(
        \I_cache/cache[2][8] ), .QN(n1648) );
  DFFRX1 \I_cache/cache_reg[3][8]  ( .D(n12720), .CK(clk), .RN(n5914), .Q(
        \I_cache/cache[3][8] ), .QN(n3230) );
  DFFRX1 \I_cache/cache_reg[4][8]  ( .D(n12719), .CK(clk), .RN(n5914), .Q(
        \I_cache/cache[4][8] ), .QN(n3217) );
  DFFRX1 \I_cache/cache_reg[5][8]  ( .D(n12718), .CK(clk), .RN(n5914), .Q(
        \I_cache/cache[5][8] ), .QN(n1420) );
  DFFRX1 \I_cache/cache_reg[6][8]  ( .D(n12717), .CK(clk), .RN(n5914), .Q(
        \I_cache/cache[6][8] ), .QN(n1707) );
  DFFRX1 \I_cache/cache_reg[7][8]  ( .D(n12716), .CK(clk), .RN(n5914), .Q(
        \I_cache/cache[7][8] ), .QN(n3304) );
  DFFRX1 \I_cache/cache_reg[0][9]  ( .D(n12715), .CK(clk), .RN(n5913), .Q(
        \I_cache/cache[0][9] ), .QN(n1705) );
  DFFRX1 \I_cache/cache_reg[1][9]  ( .D(n12714), .CK(clk), .RN(n5913), .Q(
        \I_cache/cache[1][9] ), .QN(n3301) );
  DFFRX1 \I_cache/cache_reg[2][9]  ( .D(n12713), .CK(clk), .RN(n5913), .Q(
        \I_cache/cache[2][9] ), .QN(n1704) );
  DFFRX1 \I_cache/cache_reg[3][9]  ( .D(n12712), .CK(clk), .RN(n5913), .Q(
        \I_cache/cache[3][9] ), .QN(n3300) );
  DFFRX1 \I_cache/cache_reg[4][9]  ( .D(n12711), .CK(clk), .RN(n5913), .Q(
        \I_cache/cache[4][9] ), .QN(n1288) );
  DFFRX1 \I_cache/cache_reg[5][9]  ( .D(n12710), .CK(clk), .RN(n5913), .Q(
        \I_cache/cache[5][9] ), .QN(n2821) );
  DFFRX1 \I_cache/cache_reg[6][9]  ( .D(n12709), .CK(clk), .RN(n5913), .Q(
        \I_cache/cache[6][9] ), .QN(n1706) );
  DFFRX1 \I_cache/cache_reg[7][9]  ( .D(n12708), .CK(clk), .RN(n5913), .Q(
        \I_cache/cache[7][9] ), .QN(n3302) );
  DFFRX1 \I_cache/cache_reg[0][10]  ( .D(n12707), .CK(clk), .RN(n5913), .Q(
        \I_cache/cache[0][10] ), .QN(n1495) );
  DFFRX1 \I_cache/cache_reg[1][10]  ( .D(n12706), .CK(clk), .RN(n5913), .Q(
        \I_cache/cache[1][10] ), .QN(n3255) );
  DFFRX1 \I_cache/cache_reg[2][10]  ( .D(n12705), .CK(clk), .RN(n5913), .Q(
        \I_cache/cache[2][10] ), .QN(n1670) );
  DFFRX1 \I_cache/cache_reg[3][10]  ( .D(n12704), .CK(clk), .RN(n5913), .Q(
        \I_cache/cache[3][10] ), .QN(n3254) );
  DFFRX1 \I_cache/cache_reg[4][10]  ( .D(n12703), .CK(clk), .RN(n5912), .Q(
        \I_cache/cache[4][10] ), .QN(n1475) );
  DFFRX1 \I_cache/cache_reg[5][10]  ( .D(n12702), .CK(clk), .RN(n5912), .Q(
        \I_cache/cache[5][10] ), .QN(n3049) );
  DFFRX1 \I_cache/cache_reg[6][10]  ( .D(n12701), .CK(clk), .RN(n5912), .Q(
        \I_cache/cache[6][10] ), .QN(n1671) );
  DFFRX1 \I_cache/cache_reg[7][10]  ( .D(n12700), .CK(clk), .RN(n5912), .Q(
        \I_cache/cache[7][10] ), .QN(n3256) );
  DFFRX1 \I_cache/cache_reg[0][11]  ( .D(n12699), .CK(clk), .RN(n5912), .Q(
        \I_cache/cache[0][11] ), .QN(n646) );
  DFFRX1 \I_cache/cache_reg[1][11]  ( .D(n12698), .CK(clk), .RN(n5912), .Q(
        \I_cache/cache[1][11] ), .QN(n2224) );
  DFFRX1 \I_cache/cache_reg[2][11]  ( .D(n12697), .CK(clk), .RN(n5912), .Q(
        \I_cache/cache[2][11] ), .QN(n1143) );
  DFFRX1 \I_cache/cache_reg[3][11]  ( .D(n12696), .CK(clk), .RN(n5912), .Q(
        \I_cache/cache[3][11] ), .QN(n2738) );
  DFFRX1 \I_cache/cache_reg[4][11]  ( .D(n12695), .CK(clk), .RN(n5912), .Q(
        \I_cache/cache[4][11] ), .QN(n1567) );
  DFFRX1 \I_cache/cache_reg[5][11]  ( .D(n12694), .CK(clk), .RN(n5912), .Q(
        \I_cache/cache[5][11] ), .QN(n3213) );
  DFFRX1 \I_cache/cache_reg[6][11]  ( .D(n12693), .CK(clk), .RN(n5912), .Q(
        \I_cache/cache[6][11] ), .QN(n1096) );
  DFFRX1 \I_cache/cache_reg[7][11]  ( .D(n12692), .CK(clk), .RN(n5912), .Q(
        \I_cache/cache[7][11] ), .QN(n2735) );
  DFFRX1 \I_cache/cache_reg[0][12]  ( .D(n12691), .CK(clk), .RN(n5911), .Q(
        \I_cache/cache[0][12] ), .QN(n647) );
  DFFRX1 \I_cache/cache_reg[1][12]  ( .D(n12690), .CK(clk), .RN(n5911), .Q(
        \I_cache/cache[1][12] ), .QN(n2223) );
  DFFRX1 \I_cache/cache_reg[2][12]  ( .D(n12689), .CK(clk), .RN(n5911), .Q(
        \I_cache/cache[2][12] ), .QN(n3017) );
  DFFRX1 \I_cache/cache_reg[3][12]  ( .D(n12688), .CK(clk), .RN(n5911), .Q(
        \I_cache/cache[3][12] ), .QN(n723) );
  DFFRX1 \I_cache/cache_reg[4][12]  ( .D(n12687), .CK(clk), .RN(n5911), .Q(
        \I_cache/cache[4][12] ), .QN(n1569) );
  DFFRX1 \I_cache/cache_reg[5][12]  ( .D(n12686), .CK(clk), .RN(n5911), .Q(
        \I_cache/cache[5][12] ), .QN(n3151) );
  DFFRX1 \I_cache/cache_reg[6][12]  ( .D(n12685), .CK(clk), .RN(n5911), .Q(
        \I_cache/cache[6][12] ), .QN(n3067) );
  DFFRX1 \I_cache/cache_reg[7][12]  ( .D(n12684), .CK(clk), .RN(n5911), .Q(
        \I_cache/cache[7][12] ), .QN(n1175) );
  DFFRX1 \I_cache/cache_reg[0][13]  ( .D(n12683), .CK(clk), .RN(n5911), .Q(
        \I_cache/cache[0][13] ), .QN(n1585) );
  DFFRX1 \I_cache/cache_reg[1][13]  ( .D(n12682), .CK(clk), .RN(n5911), .Q(
        \I_cache/cache[1][13] ), .QN(n3165) );
  DFFRX1 \I_cache/cache_reg[2][13]  ( .D(n12681), .CK(clk), .RN(n5911), .Q(
        \I_cache/cache[2][13] ), .QN(n1584) );
  DFFRX1 \I_cache/cache_reg[3][13]  ( .D(n12680), .CK(clk), .RN(n5910), .Q(
        \I_cache/cache[3][13] ), .QN(n3164) );
  DFFRX1 \I_cache/cache_reg[4][13]  ( .D(n12679), .CK(clk), .RN(n5910), .Q(
        \I_cache/cache[4][13] ), .QN(n760) );
  DFFRX1 \I_cache/cache_reg[5][13]  ( .D(n12678), .CK(clk), .RN(n5910), .Q(
        \I_cache/cache[5][13] ), .QN(n2321) );
  DFFRX1 \I_cache/cache_reg[6][13]  ( .D(n12677), .CK(clk), .RN(n5910), .Q(
        \I_cache/cache[6][13] ), .QN(n3075) );
  DFFRX1 \I_cache/cache_reg[7][13]  ( .D(n12676), .CK(clk), .RN(n5910), .Q(
        \I_cache/cache[7][13] ), .QN(n1421) );
  DFFRX1 \I_cache/cache_reg[0][14]  ( .D(n12675), .CK(clk), .RN(n5910), .Q(
        \I_cache/cache[0][14] ), .QN(n1446) );
  DFFRX1 \I_cache/cache_reg[1][14]  ( .D(n12674), .CK(clk), .RN(n5910), .Q(
        \I_cache/cache[1][14] ), .QN(n3015) );
  DFFRX1 \I_cache/cache_reg[2][14]  ( .D(n12673), .CK(clk), .RN(n5910), .Q(
        \I_cache/cache[2][14] ), .QN(n1504) );
  DFFRX1 \I_cache/cache_reg[3][14]  ( .D(n12672), .CK(clk), .RN(n5910), .Q(
        \I_cache/cache[3][14] ), .QN(n3084) );
  DFFRX1 \I_cache/cache_reg[4][14]  ( .D(n12671), .CK(clk), .RN(n5910), .Q(
        \I_cache/cache[4][14] ), .QN(n1568) );
  DFFRX1 \I_cache/cache_reg[5][14]  ( .D(n12670), .CK(clk), .RN(n5910), .Q(
        \I_cache/cache[5][14] ), .QN(n3150) );
  DFFRX1 \I_cache/cache_reg[6][14]  ( .D(n12669), .CK(clk), .RN(n5910), .Q(
        \I_cache/cache[6][14] ), .QN(n1505) );
  DFFRX1 \I_cache/cache_reg[7][14]  ( .D(n12668), .CK(clk), .RN(n5909), .Q(
        \I_cache/cache[7][14] ), .QN(n3085) );
  DFFRX1 \I_cache/cache_reg[0][28]  ( .D(n12563), .CK(clk), .RN(n5921), .Q(
        \I_cache/cache[0][28] ), .QN(n1618) );
  DFFRX1 \I_cache/cache_reg[1][28]  ( .D(n12562), .CK(clk), .RN(n5921), .Q(
        \I_cache/cache[1][28] ), .QN(n3195) );
  DFFRX1 \I_cache/cache_reg[2][28]  ( .D(n12561), .CK(clk), .RN(n5920), .Q(
        \I_cache/cache[2][28] ), .QN(n1620) );
  DFFRX1 \I_cache/cache_reg[3][28]  ( .D(n12560), .CK(clk), .RN(n5920), .Q(
        \I_cache/cache[3][28] ), .QN(n3197) );
  DFFRX1 \I_cache/cache_reg[4][28]  ( .D(n12559), .CK(clk), .RN(n5920), .Q(
        \I_cache/cache[4][28] ), .QN(n1619) );
  DFFRX1 \I_cache/cache_reg[5][28]  ( .D(n12558), .CK(clk), .RN(n5920), .Q(
        \I_cache/cache[5][28] ), .QN(n3196) );
  DFFRX1 \I_cache/cache_reg[6][28]  ( .D(n12557), .CK(clk), .RN(n5920), .Q(
        \I_cache/cache[6][28] ), .QN(n1626) );
  DFFRX1 \I_cache/cache_reg[7][28]  ( .D(n12556), .CK(clk), .RN(n5920), .Q(
        \I_cache/cache[7][28] ), .QN(n3202) );
  DFFRX1 \I_cache/cache_reg[1][29]  ( .D(n12554), .CK(clk), .RN(n5920), .Q(
        \I_cache/cache[1][29] ), .QN(n3095) );
  DFFRX1 \I_cache/cache_reg[2][29]  ( .D(n12553), .CK(clk), .RN(n5920), .Q(
        \I_cache/cache[2][29] ), .QN(n1514) );
  DFFRX1 \I_cache/cache_reg[3][29]  ( .D(n12552), .CK(clk), .RN(n5920), .Q(
        \I_cache/cache[3][29] ), .QN(n3094) );
  DFFRX1 \I_cache/cache_reg[4][29]  ( .D(n12551), .CK(clk), .RN(n5920), .Q(
        \I_cache/cache[4][29] ), .QN(n3059) );
  DFFRX1 \I_cache/cache_reg[5][29]  ( .D(n12550), .CK(clk), .RN(n5920), .Q(
        \I_cache/cache[5][29] ), .QN(n1145) );
  DFFRX1 \I_cache/cache_reg[6][29]  ( .D(n12549), .CK(clk), .RN(n5919), .Q(
        \I_cache/cache[6][29] ), .QN(n1516) );
  DFFRX1 \I_cache/cache_reg[7][29]  ( .D(n12548), .CK(clk), .RN(n5919), .Q(
        \I_cache/cache[7][29] ), .QN(n3096) );
  DFFRX1 \I_cache/cache_reg[0][30]  ( .D(n12547), .CK(clk), .RN(n5919), .Q(
        \I_cache/cache[0][30] ), .QN(n1526) );
  DFFRX1 \I_cache/cache_reg[1][30]  ( .D(n12546), .CK(clk), .RN(n5919), .Q(
        \I_cache/cache[1][30] ), .QN(n3106) );
  DFFRX1 \I_cache/cache_reg[2][30]  ( .D(n12545), .CK(clk), .RN(n5919), .Q(
        \I_cache/cache[2][30] ), .QN(n1578) );
  DFFRX1 \I_cache/cache_reg[3][30]  ( .D(n12544), .CK(clk), .RN(n5919), .Q(
        \I_cache/cache[3][30] ), .QN(n3160) );
  DFFRX1 \I_cache/cache_reg[4][30]  ( .D(n12543), .CK(clk), .RN(n5919), .Q(
        \I_cache/cache[4][30] ), .QN(n1600) );
  DFFRX1 \I_cache/cache_reg[5][30]  ( .D(n12542), .CK(clk), .RN(n5919), .Q(
        \I_cache/cache[5][30] ), .QN(n3177) );
  DFFRX1 \I_cache/cache_reg[6][30]  ( .D(n12541), .CK(clk), .RN(n5919), .Q(
        \I_cache/cache[6][30] ), .QN(n1527) );
  DFFRX1 \I_cache/cache_reg[7][30]  ( .D(n12540), .CK(clk), .RN(n5919), .Q(
        \I_cache/cache[7][30] ), .QN(n3107) );
  DFFRX1 \I_cache/cache_reg[5][31]  ( .D(n12534), .CK(clk), .RN(n5918), .Q(
        \I_cache/cache[5][31] ), .QN(n3182) );
  DFFRX1 \I_cache/cache_reg[7][31]  ( .D(n12532), .CK(clk), .RN(n5918), .Q(
        \I_cache/cache[7][31] ), .QN(n3131) );
  DFFRX1 \I_cache/cache_reg[0][32]  ( .D(n12531), .CK(clk), .RN(n5918), .Q(
        \I_cache/cache[0][32] ), .QN(n1658) );
  DFFRX1 \I_cache/cache_reg[1][32]  ( .D(n12530), .CK(clk), .RN(n5918), .Q(
        \I_cache/cache[1][32] ), .QN(n3242) );
  DFFRX1 \I_cache/cache_reg[2][32]  ( .D(n12529), .CK(clk), .RN(n5918), .Q(
        \I_cache/cache[2][32] ), .QN(n1659) );
  DFFRX1 \I_cache/cache_reg[3][32]  ( .D(n12528), .CK(clk), .RN(n5918), .Q(
        \I_cache/cache[3][32] ), .QN(n3243) );
  DFFRX1 \I_cache/cache_reg[4][32]  ( .D(n12527), .CK(clk), .RN(n5918), .Q(
        \I_cache/cache[4][32] ), .QN(n1645) );
  DFFRX1 \I_cache/cache_reg[5][32]  ( .D(n12526), .CK(clk), .RN(n5918), .Q(
        \I_cache/cache[5][32] ), .QN(n3227) );
  DFFRX1 \I_cache/cache_reg[6][32]  ( .D(n12525), .CK(clk), .RN(n5917), .Q(
        \I_cache/cache[6][32] ), .QN(n1646) );
  DFFRX1 \I_cache/cache_reg[7][32]  ( .D(n12524), .CK(clk), .RN(n5917), .Q(
        \I_cache/cache[7][32] ), .QN(n3228) );
  DFFRX1 \I_cache/cache_reg[0][33]  ( .D(n12523), .CK(clk), .RN(n5917), .Q(
        \I_cache/cache[0][33] ), .QN(n1474) );
  DFFRX1 \I_cache/cache_reg[1][33]  ( .D(n12522), .CK(clk), .RN(n5917), .Q(
        \I_cache/cache[1][33] ), .QN(n3048) );
  DFFRX1 \I_cache/cache_reg[2][33]  ( .D(n12521), .CK(clk), .RN(n5917), .Q(
        \I_cache/cache[2][33] ), .QN(n2988) );
  DFFRX1 \I_cache/cache_reg[3][33]  ( .D(n12520), .CK(clk), .RN(n5917), .Q(
        \I_cache/cache[3][33] ), .QN(n1431) );
  DFFRX1 \I_cache/cache_reg[4][33]  ( .D(n12519), .CK(clk), .RN(n5917), .Q(
        \I_cache/cache[4][33] ), .QN(n1467) );
  DFFRX1 \I_cache/cache_reg[5][33]  ( .D(n12518), .CK(clk), .RN(n5917), .Q(
        \I_cache/cache[5][33] ), .QN(n3041) );
  DFFRX1 \I_cache/cache_reg[6][33]  ( .D(n12517), .CK(clk), .RN(n5917), .Q(
        \I_cache/cache[6][33] ), .QN(n1650) );
  DFFRX1 \I_cache/cache_reg[7][33]  ( .D(n12516), .CK(clk), .RN(n5917), .Q(
        \I_cache/cache[7][33] ), .QN(n3232) );
  DFFRX1 \I_cache/cache_reg[0][34]  ( .D(n12515), .CK(clk), .RN(n5917), .Q(
        \I_cache/cache[0][34] ), .QN(n1614) );
  DFFRX1 \I_cache/cache_reg[1][34]  ( .D(n12514), .CK(clk), .RN(n5917), .Q(
        \I_cache/cache[1][34] ), .QN(n3191) );
  DFFRX1 \I_cache/cache_reg[2][34]  ( .D(n12513), .CK(clk), .RN(n5916), .Q(
        \I_cache/cache[2][34] ), .QN(n1616) );
  DFFRX1 \I_cache/cache_reg[3][34]  ( .D(n12512), .CK(clk), .RN(n5916), .Q(
        \I_cache/cache[3][34] ), .QN(n3193) );
  DFFRX1 \I_cache/cache_reg[4][34]  ( .D(n12511), .CK(clk), .RN(n5916), .Q(
        \I_cache/cache[4][34] ), .QN(n1615) );
  DFFRX1 \I_cache/cache_reg[5][34]  ( .D(n12510), .CK(clk), .RN(n5916), .Q(
        \I_cache/cache[5][34] ), .QN(n3192) );
  DFFRX1 \I_cache/cache_reg[6][34]  ( .D(n12509), .CK(clk), .RN(n5916), .Q(
        \I_cache/cache[6][34] ), .QN(n1624) );
  DFFRX1 \I_cache/cache_reg[7][34]  ( .D(n12508), .CK(clk), .RN(n5916), .Q(
        \I_cache/cache[7][34] ), .QN(n3201) );
  DFFRX1 \I_cache/cache_reg[0][35]  ( .D(n12507), .CK(clk), .RN(n5916), .Q(
        \I_cache/cache[0][35] ), .QN(n1682) );
  DFFRX1 \I_cache/cache_reg[1][35]  ( .D(n12506), .CK(clk), .RN(n5921), .Q(
        \I_cache/cache[1][35] ), .QN(n3273) );
  DFFRX1 \I_cache/cache_reg[2][35]  ( .D(n12505), .CK(clk), .RN(n5926), .Q(
        \I_cache/cache[2][35] ), .QN(n1667) );
  DFFRX1 \I_cache/cache_reg[3][35]  ( .D(n12504), .CK(clk), .RN(n5826), .Q(
        \I_cache/cache[3][35] ), .QN(n3251) );
  DFFRX1 \I_cache/cache_reg[4][35]  ( .D(n12503), .CK(clk), .RN(n5816), .Q(
        \I_cache/cache[4][35] ), .QN(n1666) );
  DFFRX1 \I_cache/cache_reg[5][35]  ( .D(n12502), .CK(clk), .RN(n5816), .Q(
        \I_cache/cache[5][35] ), .QN(n3250) );
  DFFRX1 \I_cache/cache_reg[6][35]  ( .D(n12501), .CK(clk), .RN(n5816), .Q(
        \I_cache/cache[6][35] ), .QN(n1225) );
  DFFRX1 \I_cache/cache_reg[7][35]  ( .D(n12500), .CK(clk), .RN(n5816), .Q(
        \I_cache/cache[7][35] ), .QN(n2762) );
  DFFRX1 \I_cache/cache_reg[0][36]  ( .D(n12499), .CK(clk), .RN(n5816), .Q(
        \I_cache/cache[0][36] ), .QN(n2990) );
  DFFRX1 \I_cache/cache_reg[1][36]  ( .D(n12498), .CK(clk), .RN(n5816), .Q(
        \I_cache/cache[1][36] ), .QN(n1432) );
  DFFRX1 \I_cache/cache_reg[2][36]  ( .D(n12497), .CK(clk), .RN(n5816), .Q(
        \I_cache/cache[2][36] ), .QN(n1675) );
  DFFRX1 \I_cache/cache_reg[3][36]  ( .D(n12496), .CK(clk), .RN(n5815), .Q(
        \I_cache/cache[3][36] ), .QN(n3263) );
  DFFRX1 \I_cache/cache_reg[4][36]  ( .D(n12495), .CK(clk), .RN(n5815), .Q(
        \I_cache/cache[4][36] ), .QN(n1674) );
  DFFRX1 \I_cache/cache_reg[5][36]  ( .D(n12494), .CK(clk), .RN(n5815), .Q(
        \I_cache/cache[5][36] ), .QN(n3262) );
  DFFRX1 \I_cache/cache_reg[6][36]  ( .D(n12493), .CK(clk), .RN(n5815), .Q(
        \I_cache/cache[6][36] ), .QN(n1708) );
  DFFRX1 \I_cache/cache_reg[7][36]  ( .D(n12492), .CK(clk), .RN(n5815), .Q(
        \I_cache/cache[7][36] ), .QN(n3305) );
  DFFRX1 \I_cache/cache_reg[0][37]  ( .D(n12491), .CK(clk), .RN(n5815), .Q(
        \I_cache/cache[0][37] ), .QN(n2741) );
  DFFRX1 \I_cache/cache_reg[1][37]  ( .D(n12490), .CK(clk), .RN(n5815), .Q(
        \I_cache/cache[1][37] ), .QN(n1281) );
  DFFRX1 \I_cache/cache_reg[2][37]  ( .D(n12489), .CK(clk), .RN(n5815), .Q(
        \I_cache/cache[2][37] ), .QN(n1506) );
  DFFRX1 \I_cache/cache_reg[3][37]  ( .D(n12488), .CK(clk), .RN(n5815), .Q(
        \I_cache/cache[3][37] ), .QN(n3086) );
  DFFRX1 \I_cache/cache_reg[4][37]  ( .D(n12487), .CK(clk), .RN(n5815), .Q(
        \I_cache/cache[4][37] ), .QN(n1579) );
  DFFRX1 \I_cache/cache_reg[5][37]  ( .D(n12486), .CK(clk), .RN(n5815), .Q(
        \I_cache/cache[5][37] ), .QN(n3161) );
  DFFRX1 \I_cache/cache_reg[6][37]  ( .D(n12485), .CK(clk), .RN(n5815), .Q(
        \I_cache/cache[6][37] ), .QN(n1596) );
  DFFRX1 \I_cache/cache_reg[7][37]  ( .D(n12484), .CK(clk), .RN(n5814), .Q(
        \I_cache/cache[7][37] ), .QN(n3173) );
  DFFRX1 \I_cache/cache_reg[0][38]  ( .D(n12483), .CK(clk), .RN(n5814), .Q(
        \I_cache/cache[0][38] ), .QN(n1702) );
  DFFRX1 \I_cache/cache_reg[1][38]  ( .D(n12482), .CK(clk), .RN(n5814), .Q(
        \I_cache/cache[1][38] ), .QN(n3298) );
  DFFRX1 \I_cache/cache_reg[2][38]  ( .D(n12481), .CK(clk), .RN(n5814), .Q(
        \I_cache/cache[2][38] ), .QN(n1701) );
  DFFRX1 \I_cache/cache_reg[3][38]  ( .D(n12480), .CK(clk), .RN(n5814), .Q(
        \I_cache/cache[3][38] ), .QN(n3297) );
  DFFRX1 \I_cache/cache_reg[4][38]  ( .D(n12479), .CK(clk), .RN(n5814), .Q(
        \I_cache/cache[4][38] ), .QN(n1383) );
  DFFRX1 \I_cache/cache_reg[5][38]  ( .D(n12478), .CK(clk), .RN(n5814), .Q(
        \I_cache/cache[5][38] ), .QN(n2913) );
  DFFRX1 \I_cache/cache_reg[6][38]  ( .D(n12477), .CK(clk), .RN(n5814), .Q(
        \I_cache/cache[6][38] ), .QN(n1703) );
  DFFRX1 \I_cache/cache_reg[7][38]  ( .D(n12476), .CK(clk), .RN(n5814), .Q(
        \I_cache/cache[7][38] ), .QN(n3299) );
  DFFRX1 \I_cache/cache_reg[0][39]  ( .D(n12475), .CK(clk), .RN(n5814), .Q(
        \I_cache/cache[0][39] ), .QN(n1649) );
  DFFRX1 \I_cache/cache_reg[1][39]  ( .D(n12474), .CK(clk), .RN(n5814), .Q(
        \I_cache/cache[1][39] ), .QN(n3231) );
  DFFRX1 \I_cache/cache_reg[2][39]  ( .D(n12473), .CK(clk), .RN(n5814), .Q(
        \I_cache/cache[2][39] ), .QN(n1696) );
  DFFRX1 \I_cache/cache_reg[3][39]  ( .D(n12472), .CK(clk), .RN(n5813), .Q(
        \I_cache/cache[3][39] ), .QN(n3292) );
  DFFRX1 \I_cache/cache_reg[4][39]  ( .D(n12471), .CK(clk), .RN(n5813), .Q(
        \I_cache/cache[4][39] ), .QN(n1220) );
  DFFRX1 \I_cache/cache_reg[5][39]  ( .D(n12470), .CK(clk), .RN(n5813), .Q(
        \I_cache/cache[5][39] ), .QN(n2757) );
  DFFRX1 \I_cache/cache_reg[6][39]  ( .D(n12469), .CK(clk), .RN(n5813), .Q(
        \I_cache/cache[6][39] ), .QN(n1461) );
  DFFRX1 \I_cache/cache_reg[7][39]  ( .D(n12468), .CK(clk), .RN(n5813), .Q(
        \I_cache/cache[7][39] ), .QN(n3035) );
  DFFRX1 \I_cache/cache_reg[0][40]  ( .D(n12467), .CK(clk), .RN(n5813), .Q(
        \I_cache/cache[0][40] ), .QN(n1684) );
  DFFRX1 \I_cache/cache_reg[1][40]  ( .D(n12466), .CK(clk), .RN(n5813), .Q(
        \I_cache/cache[1][40] ), .QN(n3277) );
  DFFRX1 \I_cache/cache_reg[2][40]  ( .D(n12465), .CK(clk), .RN(n5813), .Q(
        \I_cache/cache[2][40] ), .QN(n1643) );
  DFFRX1 \I_cache/cache_reg[3][40]  ( .D(n12464), .CK(clk), .RN(n5813), .Q(
        \I_cache/cache[3][40] ), .QN(n3225) );
  DFFRX1 \I_cache/cache_reg[4][40]  ( .D(n12463), .CK(clk), .RN(n5813), .Q(
        \I_cache/cache[4][40] ), .QN(n1287) );
  DFFRX1 \I_cache/cache_reg[5][40]  ( .D(n12462), .CK(clk), .RN(n5813), .Q(
        \I_cache/cache[5][40] ), .QN(n2820) );
  DFFRX1 \I_cache/cache_reg[6][40]  ( .D(n12461), .CK(clk), .RN(n5813), .Q(
        \I_cache/cache[6][40] ), .QN(n1642) );
  DFFRX1 \I_cache/cache_reg[7][40]  ( .D(n12460), .CK(clk), .RN(n5812), .Q(
        \I_cache/cache[7][40] ), .QN(n3224) );
  DFFRX1 \I_cache/cache_reg[0][41]  ( .D(n12459), .CK(clk), .RN(n5812), .Q(
        \I_cache/cache[0][41] ), .QN(n1692) );
  DFFRX1 \I_cache/cache_reg[1][41]  ( .D(n12458), .CK(clk), .RN(n5812), .Q(
        \I_cache/cache[1][41] ), .QN(n3288) );
  DFFRX1 \I_cache/cache_reg[2][41]  ( .D(n12457), .CK(clk), .RN(n5812), .Q(
        \I_cache/cache[2][41] ), .QN(n1473) );
  DFFRX1 \I_cache/cache_reg[3][41]  ( .D(n12456), .CK(clk), .RN(n5812), .Q(
        \I_cache/cache[3][41] ), .QN(n3047) );
  DFFRX1 \I_cache/cache_reg[4][41]  ( .D(n12455), .CK(clk), .RN(n5812), .Q(
        \I_cache/cache[4][41] ), .QN(n765) );
  DFFRX1 \I_cache/cache_reg[5][41]  ( .D(n12454), .CK(clk), .RN(n5812), .Q(
        \I_cache/cache[5][41] ), .QN(n2327) );
  DFFRX1 \I_cache/cache_reg[6][41]  ( .D(n12453), .CK(clk), .RN(n5812), .Q(
        \I_cache/cache[6][41] ), .QN(n1638) );
  DFFRX1 \I_cache/cache_reg[7][41]  ( .D(n12452), .CK(clk), .RN(n5812), .Q(
        \I_cache/cache[7][41] ), .QN(n3220) );
  DFFRX1 \I_cache/cache_reg[0][42]  ( .D(n12451), .CK(clk), .RN(n5812), .Q(
        \I_cache/cache[0][42] ), .QN(n1493) );
  DFFRX1 \I_cache/cache_reg[1][42]  ( .D(n12450), .CK(clk), .RN(n5812), .Q(
        \I_cache/cache[1][42] ), .QN(n3211) );
  DFFRX1 \I_cache/cache_reg[2][42]  ( .D(n12449), .CK(clk), .RN(n5812), .Q(
        \I_cache/cache[2][42] ), .QN(n1492) );
  DFFRX1 \I_cache/cache_reg[3][42]  ( .D(n12448), .CK(clk), .RN(n5811), .Q(
        \I_cache/cache[3][42] ), .QN(n3210) );
  DFFRX1 \I_cache/cache_reg[4][42]  ( .D(n12447), .CK(clk), .RN(n5811), .Q(
        \I_cache/cache[4][42] ), .QN(n1451) );
  DFFRX1 \I_cache/cache_reg[5][42]  ( .D(n12446), .CK(clk), .RN(n5811), .Q(
        \I_cache/cache[5][42] ), .QN(n3024) );
  DFFRX1 \I_cache/cache_reg[6][42]  ( .D(n12445), .CK(clk), .RN(n5811), .Q(
        \I_cache/cache[6][42] ), .QN(n1494) );
  DFFRX1 \I_cache/cache_reg[7][42]  ( .D(n12444), .CK(clk), .RN(n5811), .Q(
        \I_cache/cache[7][42] ), .QN(n3212) );
  DFFRX1 \I_cache/cache_reg[0][43]  ( .D(n12443), .CK(clk), .RN(n5811), .Q(
        \I_cache/cache[0][43] ), .QN(n1092) );
  DFFRX1 \I_cache/cache_reg[1][43]  ( .D(n12442), .CK(clk), .RN(n5811), .Q(
        \I_cache/cache[1][43] ), .QN(n2684) );
  DFFRX1 \I_cache/cache_reg[2][43]  ( .D(n12441), .CK(clk), .RN(n5811), .Q(
        \I_cache/cache[2][43] ), .QN(n1091) );
  DFFRX1 \I_cache/cache_reg[3][43]  ( .D(n12440), .CK(clk), .RN(n5811), .Q(
        \I_cache/cache[3][43] ), .QN(n2683) );
  DFFRX1 \I_cache/cache_reg[4][43]  ( .D(n12439), .CK(clk), .RN(n5811), .Q(
        \I_cache/cache[4][43] ), .QN(n687) );
  DFFRX1 \I_cache/cache_reg[5][43]  ( .D(n12438), .CK(clk), .RN(n5811), .Q(
        \I_cache/cache[5][43] ), .QN(n2298) );
  DFFRX1 \I_cache/cache_reg[6][43]  ( .D(n12437), .CK(clk), .RN(n5810), .Q(
        \I_cache/cache[6][43] ), .QN(n1093) );
  DFFRX1 \I_cache/cache_reg[7][43]  ( .D(n12436), .CK(clk), .RN(n5810), .Q(
        \I_cache/cache[7][43] ), .QN(n2734) );
  DFFRX1 \I_cache/cache_reg[0][44]  ( .D(n12435), .CK(clk), .RN(n5810), .Q(
        \I_cache/cache[0][44] ), .QN(n1102) );
  DFFRX1 \I_cache/cache_reg[1][44]  ( .D(n12434), .CK(clk), .RN(n5810), .Q(
        \I_cache/cache[1][44] ), .QN(n2691) );
  DFFRX1 \I_cache/cache_reg[2][44]  ( .D(n12433), .CK(clk), .RN(n5810), .Q(
        \I_cache/cache[2][44] ), .QN(n1101) );
  DFFRX1 \I_cache/cache_reg[3][44]  ( .D(n12432), .CK(clk), .RN(n5810), .Q(
        \I_cache/cache[3][44] ), .QN(n2690) );
  DFFRX1 \I_cache/cache_reg[4][44]  ( .D(n12431), .CK(clk), .RN(n5810), .Q(
        \I_cache/cache[4][44] ), .QN(n1169) );
  DFFRX1 \I_cache/cache_reg[5][44]  ( .D(n12430), .CK(clk), .RN(n5810), .Q(
        \I_cache/cache[5][44] ), .QN(n2725) );
  DFFRX1 \I_cache/cache_reg[6][44]  ( .D(n12429), .CK(clk), .RN(n5810), .Q(
        \I_cache/cache[6][44] ), .QN(n1103) );
  DFFRX1 \I_cache/cache_reg[7][44]  ( .D(n12428), .CK(clk), .RN(n5810), .Q(
        \I_cache/cache[7][44] ), .QN(n2692) );
  DFFRX1 \I_cache/cache_reg[0][45]  ( .D(n12427), .CK(clk), .RN(n5810), .Q(
        \I_cache/cache[0][45] ), .QN(n1491) );
  DFFRX1 \I_cache/cache_reg[1][45]  ( .D(n12426), .CK(clk), .RN(n5810), .Q(
        \I_cache/cache[1][45] ), .QN(n3236) );
  DFFRX1 \I_cache/cache_reg[2][45]  ( .D(n12425), .CK(clk), .RN(n5809), .Q(
        \I_cache/cache[2][45] ), .QN(n1490) );
  DFFRX1 \I_cache/cache_reg[3][45]  ( .D(n12424), .CK(clk), .RN(n5809), .Q(
        \I_cache/cache[3][45] ), .QN(n3235) );
  DFFRX1 \I_cache/cache_reg[4][45]  ( .D(n12423), .CK(clk), .RN(n5809), .Q(
        \I_cache/cache[4][45] ), .QN(n2989) );
  DFFRX1 \I_cache/cache_reg[5][45]  ( .D(n12422), .CK(clk), .RN(n5809), .Q(
        \I_cache/cache[5][45] ), .QN(n548) );
  DFFRX1 \I_cache/cache_reg[6][45]  ( .D(n12421), .CK(clk), .RN(n5809), .Q(
        \I_cache/cache[6][45] ), .QN(n1653) );
  DFFRX1 \I_cache/cache_reg[7][45]  ( .D(n12420), .CK(clk), .RN(n5809), .Q(
        \I_cache/cache[7][45] ), .QN(n3237) );
  DFFRX1 \I_cache/cache_reg[0][46]  ( .D(n12419), .CK(clk), .RN(n5809), .Q(
        \I_cache/cache[0][46] ), .QN(n1499) );
  DFFRX1 \I_cache/cache_reg[1][46]  ( .D(n12418), .CK(clk), .RN(n5809), .Q(
        \I_cache/cache[1][46] ), .QN(n3079) );
  DFFRX1 \I_cache/cache_reg[2][46]  ( .D(n12417), .CK(clk), .RN(n5809), .Q(
        \I_cache/cache[2][46] ), .QN(n3064) );
  DFFRX1 \I_cache/cache_reg[3][46]  ( .D(n12416), .CK(clk), .RN(n5809), .Q(
        \I_cache/cache[3][46] ), .QN(n1173) );
  DFFRX1 \I_cache/cache_reg[4][46]  ( .D(n12415), .CK(clk), .RN(n5809), .Q(
        \I_cache/cache[4][46] ), .QN(n1080) );
  DFFRX1 \I_cache/cache_reg[5][46]  ( .D(n12414), .CK(clk), .RN(n5809), .Q(
        \I_cache/cache[5][46] ), .QN(n2673) );
  DFFRX1 \I_cache/cache_reg[6][46]  ( .D(n12413), .CK(clk), .RN(n5808), .Q(
        \I_cache/cache[6][46] ), .QN(n3071) );
  DFFRX1 \I_cache/cache_reg[7][46]  ( .D(n12412), .CK(clk), .RN(n5808), .Q(
        \I_cache/cache[7][46] ), .QN(n1183) );
  DFFRX1 \I_cache/cache_reg[0][60]  ( .D(n12307), .CK(clk), .RN(n5819), .Q(
        \I_cache/cache[0][60] ), .QN(n1621) );
  DFFRX1 \I_cache/cache_reg[1][60]  ( .D(n12306), .CK(clk), .RN(n5819), .Q(
        \I_cache/cache[1][60] ), .QN(n3198) );
  DFFRX1 \I_cache/cache_reg[2][60]  ( .D(n12305), .CK(clk), .RN(n5819), .Q(
        \I_cache/cache[2][60] ), .QN(n3113) );
  DFFRX1 \I_cache/cache_reg[3][60]  ( .D(n12304), .CK(clk), .RN(n5819), .Q(
        \I_cache/cache[3][60] ), .QN(n1203) );
  DFFRX1 \I_cache/cache_reg[4][60]  ( .D(n12303), .CK(clk), .RN(n5819), .Q(
        \I_cache/cache[4][60] ), .QN(n3112) );
  DFFRX1 \I_cache/cache_reg[5][60]  ( .D(n12302), .CK(clk), .RN(n5819), .Q(
        \I_cache/cache[5][60] ), .QN(n1202) );
  DFFRX1 \I_cache/cache_reg[6][60]  ( .D(n12301), .CK(clk), .RN(n5819), .Q(
        \I_cache/cache[6][60] ), .QN(n1627) );
  DFFRX1 \I_cache/cache_reg[7][60]  ( .D(n12300), .CK(clk), .RN(n5819), .Q(
        \I_cache/cache[7][60] ), .QN(n3203) );
  DFFRX1 \I_cache/cache_reg[0][61]  ( .D(n12299), .CK(clk), .RN(n5819), .Q(
        \I_cache/cache[0][61] ), .QN(n1521) );
  DFFRX1 \I_cache/cache_reg[1][61]  ( .D(n12298), .CK(clk), .RN(n5819), .Q(
        \I_cache/cache[1][61] ), .QN(n3101) );
  DFFRX1 \I_cache/cache_reg[2][61]  ( .D(n12297), .CK(clk), .RN(n5819), .Q(
        \I_cache/cache[2][61] ), .QN(n1520) );
  DFFRX1 \I_cache/cache_reg[3][61]  ( .D(n12296), .CK(clk), .RN(n5819), .Q(
        \I_cache/cache[3][61] ), .QN(n3100) );
  DFFRX1 \I_cache/cache_reg[4][61]  ( .D(n12295), .CK(clk), .RN(n5818), .Q(
        \I_cache/cache[4][61] ), .QN(n1599) );
  DFFRX1 \I_cache/cache_reg[5][61]  ( .D(n12294), .CK(clk), .RN(n5818), .Q(
        \I_cache/cache[5][61] ), .QN(n3176) );
  DFFRX1 \I_cache/cache_reg[6][61]  ( .D(n12293), .CK(clk), .RN(n5818), .Q(
        \I_cache/cache[6][61] ), .QN(n1522) );
  DFFRX1 \I_cache/cache_reg[7][61]  ( .D(n12292), .CK(clk), .RN(n5818), .Q(
        \I_cache/cache[7][61] ), .QN(n3102) );
  DFFRX1 \I_cache/cache_reg[0][62]  ( .D(n12291), .CK(clk), .RN(n5818), .Q(
        \I_cache/cache[0][62] ), .QN(n1530) );
  DFFRX1 \I_cache/cache_reg[1][62]  ( .D(n12290), .CK(clk), .RN(n5818), .Q(
        \I_cache/cache[1][62] ), .QN(n3110) );
  DFFRX1 \I_cache/cache_reg[2][62]  ( .D(n12289), .CK(clk), .RN(n5818), .Q(
        \I_cache/cache[2][62] ), .QN(n1529) );
  DFFRX1 \I_cache/cache_reg[3][62]  ( .D(n12288), .CK(clk), .RN(n5818), .Q(
        \I_cache/cache[3][62] ), .QN(n3109) );
  DFFRX1 \I_cache/cache_reg[4][62]  ( .D(n12287), .CK(clk), .RN(n5818), .Q(
        \I_cache/cache[4][62] ), .QN(n1598) );
  DFFRX1 \I_cache/cache_reg[5][62]  ( .D(n12286), .CK(clk), .RN(n5818), .Q(
        \I_cache/cache[5][62] ), .QN(n3175) );
  DFFRX1 \I_cache/cache_reg[6][62]  ( .D(n12285), .CK(clk), .RN(n5818), .Q(
        \I_cache/cache[6][62] ), .QN(n1531) );
  DFFRX1 \I_cache/cache_reg[7][62]  ( .D(n12284), .CK(clk), .RN(n5818), .Q(
        \I_cache/cache[7][62] ), .QN(n3111) );
  DFFRX1 \I_cache/cache_reg[3][63]  ( .D(n12280), .CK(clk), .RN(n5817), .Q(
        \I_cache/cache[3][63] ), .QN(n3135) );
  DFFRX1 \I_cache/cache_reg[5][63]  ( .D(n12278), .CK(clk), .RN(n5817), .Q(
        \I_cache/cache[5][63] ), .QN(n3180) );
  DFFRX1 \I_cache/cache_reg[7][63]  ( .D(n12276), .CK(clk), .RN(n5817), .Q(
        \I_cache/cache[7][63] ), .QN(n3137) );
  DFFRX1 \I_cache/cache_reg[0][64]  ( .D(n12275), .CK(clk), .RN(n5817), .Q(
        \I_cache/cache[0][64] ), .QN(n1459) );
  DFFRX1 \I_cache/cache_reg[1][64]  ( .D(n12274), .CK(clk), .RN(n5817), .Q(
        \I_cache/cache[1][64] ), .QN(n3033) );
  DFFRX1 \I_cache/cache_reg[2][64]  ( .D(n12273), .CK(clk), .RN(n5817), .Q(
        \I_cache/cache[2][64] ), .QN(n1657) );
  DFFRX1 \I_cache/cache_reg[3][64]  ( .D(n12272), .CK(clk), .RN(n5817), .Q(
        \I_cache/cache[3][64] ), .QN(n3241) );
  DFFRX1 \I_cache/cache_reg[4][64]  ( .D(n12271), .CK(clk), .RN(n5816), .Q(
        \I_cache/cache[4][64] ), .QN(n1656) );
  DFFRX1 \I_cache/cache_reg[5][64]  ( .D(n12270), .CK(clk), .RN(n5816), .Q(
        \I_cache/cache[5][64] ), .QN(n3240) );
  DFFRX1 \I_cache/cache_reg[6][64]  ( .D(n12269), .CK(clk), .RN(n5816), .Q(
        \I_cache/cache[6][64] ), .QN(n3001) );
  DFFRX1 \I_cache/cache_reg[7][64]  ( .D(n12268), .CK(clk), .RN(n5816), .Q(
        \I_cache/cache[7][64] ), .QN(n1438) );
  DFFRX1 \I_cache/cache_reg[0][65]  ( .D(n12267), .CK(clk), .RN(n5816), .Q(
        \I_cache/cache[0][65] ), .QN(n1655) );
  DFFRX1 \I_cache/cache_reg[1][65]  ( .D(n12266), .CK(clk), .RN(n5821), .Q(
        \I_cache/cache[1][65] ), .QN(n3239) );
  DFFRX1 \I_cache/cache_reg[2][65]  ( .D(n12265), .CK(clk), .RN(n5796), .Q(
        \I_cache/cache[2][65] ), .QN(n1464) );
  DFFRX1 \I_cache/cache_reg[3][65]  ( .D(n12264), .CK(clk), .RN(n5796), .Q(
        \I_cache/cache[3][65] ), .QN(n3038) );
  DFFRX1 \I_cache/cache_reg[4][65]  ( .D(n12263), .CK(clk), .RN(n5796), .Q(
        \I_cache/cache[4][65] ), .QN(n1636) );
  DFFRX1 \I_cache/cache_reg[5][65]  ( .D(n12262), .CK(clk), .RN(n5796), .Q(
        \I_cache/cache[5][65] ), .QN(n3218) );
  DFFRX1 \I_cache/cache_reg[6][65]  ( .D(n12261), .CK(clk), .RN(n5796), .Q(
        \I_cache/cache[6][65] ), .QN(n1462) );
  DFFRX1 \I_cache/cache_reg[7][65]  ( .D(n12260), .CK(clk), .RN(n5796), .Q(
        \I_cache/cache[7][65] ), .QN(n3036) );
  DFFRX1 \I_cache/cache_reg[0][66]  ( .D(n12259), .CK(clk), .RN(n5796), .Q(
        \I_cache/cache[0][66] ), .QN(n1611) );
  DFFRX1 \I_cache/cache_reg[1][66]  ( .D(n12258), .CK(clk), .RN(n5796), .Q(
        \I_cache/cache[1][66] ), .QN(n3188) );
  DFFRX1 \I_cache/cache_reg[2][66]  ( .D(n12257), .CK(clk), .RN(n5795), .Q(
        \I_cache/cache[2][66] ), .QN(n1613) );
  DFFRX1 \I_cache/cache_reg[3][66]  ( .D(n12256), .CK(clk), .RN(n5795), .Q(
        \I_cache/cache[3][66] ), .QN(n3190) );
  DFFRX1 \I_cache/cache_reg[4][66]  ( .D(n12255), .CK(clk), .RN(n5795), .Q(
        \I_cache/cache[4][66] ), .QN(n1612) );
  DFFRX1 \I_cache/cache_reg[5][66]  ( .D(n12254), .CK(clk), .RN(n5795), .Q(
        \I_cache/cache[5][66] ), .QN(n3189) );
  DFFRX1 \I_cache/cache_reg[6][66]  ( .D(n12253), .CK(clk), .RN(n5795), .Q(
        \I_cache/cache[6][66] ), .QN(n1589) );
  DFFRX1 \I_cache/cache_reg[7][66]  ( .D(n12252), .CK(clk), .RN(n5795), .Q(
        \I_cache/cache[7][66] ), .QN(n3167) );
  DFFRX1 \I_cache/cache_reg[0][67]  ( .D(n12251), .CK(clk), .RN(n5795), .Q(
        \I_cache/cache[0][67] ), .QN(n1639) );
  DFFRX1 \I_cache/cache_reg[1][67]  ( .D(n12250), .CK(clk), .RN(n5795), .Q(
        \I_cache/cache[1][67] ), .QN(n3221) );
  DFFRX1 \I_cache/cache_reg[2][67]  ( .D(n12249), .CK(clk), .RN(n5795), .Q(
        \I_cache/cache[2][67] ), .QN(n1665) );
  DFFRX1 \I_cache/cache_reg[3][67]  ( .D(n12248), .CK(clk), .RN(n5795), .Q(
        \I_cache/cache[3][67] ), .QN(n3249) );
  DFFRX1 \I_cache/cache_reg[4][67]  ( .D(n12247), .CK(clk), .RN(n5795), .Q(
        \I_cache/cache[4][67] ), .QN(n1664) );
  DFFRX1 \I_cache/cache_reg[5][67]  ( .D(n12246), .CK(clk), .RN(n5795), .Q(
        \I_cache/cache[5][67] ), .QN(n3248) );
  DFFRX1 \I_cache/cache_reg[6][67]  ( .D(n12245), .CK(clk), .RN(n5794), .Q(
        \I_cache/cache[6][67] ), .QN(n2986) );
  DFFRX1 \I_cache/cache_reg[7][67]  ( .D(n12244), .CK(clk), .RN(n5794), .Q(
        \I_cache/cache[7][67] ), .QN(n1430) );
  DFFRX1 \I_cache/cache_reg[0][68]  ( .D(n12243), .CK(clk), .RN(n5794), .Q(
        \I_cache/cache[0][68] ), .QN(n2991) );
  DFFRX1 \I_cache/cache_reg[1][68]  ( .D(n12242), .CK(clk), .RN(n5794), .Q(
        \I_cache/cache[1][68] ), .QN(n1433) );
  DFFRX1 \I_cache/cache_reg[2][68]  ( .D(n12241), .CK(clk), .RN(n5794), .Q(
        \I_cache/cache[2][68] ), .QN(n1673) );
  DFFRX1 \I_cache/cache_reg[3][68]  ( .D(n12240), .CK(clk), .RN(n5794), .Q(
        \I_cache/cache[3][68] ), .QN(n3261) );
  DFFRX1 \I_cache/cache_reg[4][68]  ( .D(n12239), .CK(clk), .RN(n5794), .Q(
        \I_cache/cache[4][68] ), .QN(n1672) );
  DFFRX1 \I_cache/cache_reg[5][68]  ( .D(n12238), .CK(clk), .RN(n5794), .Q(
        \I_cache/cache[5][68] ), .QN(n3260) );
  DFFRX1 \I_cache/cache_reg[6][68]  ( .D(n12237), .CK(clk), .RN(n5794), .Q(
        \I_cache/cache[6][68] ), .QN(n1641) );
  DFFRX1 \I_cache/cache_reg[7][68]  ( .D(n12236), .CK(clk), .RN(n5794), .Q(
        \I_cache/cache[7][68] ), .QN(n3223) );
  DFFRX1 \I_cache/cache_reg[0][69]  ( .D(n12235), .CK(clk), .RN(n5794), .Q(
        \I_cache/cache[0][69] ), .QN(n1500) );
  DFFRX1 \I_cache/cache_reg[1][69]  ( .D(n12234), .CK(clk), .RN(n5794), .Q(
        \I_cache/cache[1][69] ), .QN(n3080) );
  DFFRX1 \I_cache/cache_reg[2][69]  ( .D(n12233), .CK(clk), .RN(n5793), .Q(
        \I_cache/cache[2][69] ), .QN(n1610) );
  DFFRX1 \I_cache/cache_reg[3][69]  ( .D(n12232), .CK(clk), .RN(n5793), .Q(
        \I_cache/cache[3][69] ), .QN(n3187) );
  DFFRX1 \I_cache/cache_reg[4][69]  ( .D(n12231), .CK(clk), .RN(n5793), .Q(
        \I_cache/cache[4][69] ), .QN(n1609) );
  DFFRX1 \I_cache/cache_reg[5][69]  ( .D(n12230), .CK(clk), .RN(n5793), .Q(
        \I_cache/cache[5][69] ), .QN(n3186) );
  DFFRX1 \I_cache/cache_reg[6][69]  ( .D(n12229), .CK(clk), .RN(n5793), .Q(
        \I_cache/cache[6][69] ), .QN(n1623) );
  DFFRX1 \I_cache/cache_reg[7][69]  ( .D(n12228), .CK(clk), .RN(n5793), .Q(
        \I_cache/cache[7][69] ), .QN(n3200) );
  DFFRX1 \I_cache/cache_reg[0][70]  ( .D(n12227), .CK(clk), .RN(n5793), .Q(
        \I_cache/cache[0][70] ), .QN(n1470) );
  DFFRX1 \I_cache/cache_reg[1][70]  ( .D(n12226), .CK(clk), .RN(n5793), .Q(
        \I_cache/cache[1][70] ), .QN(n3044) );
  DFFRX1 \I_cache/cache_reg[2][70]  ( .D(n12225), .CK(clk), .RN(n5793), .Q(
        \I_cache/cache[2][70] ), .QN(n1686) );
  DFFRX1 \I_cache/cache_reg[3][70]  ( .D(n12224), .CK(clk), .RN(n5793), .Q(
        \I_cache/cache[3][70] ), .QN(n3279) );
  DFFRX1 \I_cache/cache_reg[4][70]  ( .D(n12223), .CK(clk), .RN(n5793), .Q(
        \I_cache/cache[4][70] ), .QN(n1382) );
  DFFRX1 \I_cache/cache_reg[5][70]  ( .D(n12222), .CK(clk), .RN(n5793), .Q(
        \I_cache/cache[5][70] ), .QN(n2912) );
  DFFRX1 \I_cache/cache_reg[6][70]  ( .D(n12221), .CK(clk), .RN(n5792), .Q(
        \I_cache/cache[6][70] ), .QN(n1687) );
  DFFRX1 \I_cache/cache_reg[7][70]  ( .D(n12220), .CK(clk), .RN(n5792), .Q(
        \I_cache/cache[7][70] ), .QN(n3280) );
  DFFRX1 \I_cache/cache_reg[0][71]  ( .D(n12219), .CK(clk), .RN(n5792), .Q(
        \I_cache/cache[0][71] ), .QN(n1644) );
  DFFRX1 \I_cache/cache_reg[1][71]  ( .D(n12218), .CK(clk), .RN(n5792), .Q(
        \I_cache/cache[1][71] ), .QN(n3226) );
  DFFRX1 \I_cache/cache_reg[2][71]  ( .D(n12217), .CK(clk), .RN(n5792), .Q(
        \I_cache/cache[2][71] ), .QN(n1685) );
  DFFRX1 \I_cache/cache_reg[3][71]  ( .D(n12216), .CK(clk), .RN(n5792), .Q(
        \I_cache/cache[3][71] ), .QN(n3278) );
  DFFRX1 \I_cache/cache_reg[4][71]  ( .D(n12215), .CK(clk), .RN(n5792), .Q(
        \I_cache/cache[4][71] ), .QN(n1303) );
  DFFRX1 \I_cache/cache_reg[5][71]  ( .D(n12214), .CK(clk), .RN(n5792), .Q(
        \I_cache/cache[5][71] ), .QN(n3285) );
  DFFRX1 \I_cache/cache_reg[6][71]  ( .D(n12213), .CK(clk), .RN(n5792), .Q(
        \I_cache/cache[6][71] ), .QN(n3006) );
  DFFRX1 \I_cache/cache_reg[7][71]  ( .D(n12212), .CK(clk), .RN(n5792), .Q(
        \I_cache/cache[7][71] ), .QN(n1440) );
  DFFRX1 \I_cache/cache_reg[0][72]  ( .D(n12211), .CK(clk), .RN(n5792), .Q(
        \I_cache/cache[0][72] ), .QN(n1690) );
  DFFRX1 \I_cache/cache_reg[1][72]  ( .D(n12210), .CK(clk), .RN(n5792), .Q(
        \I_cache/cache[1][72] ), .QN(n3286) );
  DFFRX1 \I_cache/cache_reg[2][72]  ( .D(n12209), .CK(clk), .RN(n5791), .Q(
        \I_cache/cache[2][72] ), .QN(n1640) );
  DFFRX1 \I_cache/cache_reg[3][72]  ( .D(n12208), .CK(clk), .RN(n5791), .Q(
        \I_cache/cache[3][72] ), .QN(n3222) );
  DFFRX1 \I_cache/cache_reg[4][72]  ( .D(n12207), .CK(clk), .RN(n5791), .Q(
        \I_cache/cache[4][72] ), .QN(n1381) );
  DFFRX1 \I_cache/cache_reg[5][72]  ( .D(n12206), .CK(clk), .RN(n5791), .Q(
        \I_cache/cache[5][72] ), .QN(n2911) );
  DFFRX1 \I_cache/cache_reg[6][72]  ( .D(n12205), .CK(clk), .RN(n5791), .Q(
        \I_cache/cache[6][72] ), .QN(n1691) );
  DFFRX1 \I_cache/cache_reg[7][72]  ( .D(n12204), .CK(clk), .RN(n5791), .Q(
        \I_cache/cache[7][72] ), .QN(n3287) );
  DFFRX1 \I_cache/cache_reg[0][73]  ( .D(n12203), .CK(clk), .RN(n5791), .Q(
        \I_cache/cache[0][73] ), .QN(n480) );
  DFFRX1 \I_cache/cache_reg[1][73]  ( .D(n12202), .CK(clk), .RN(n5791), .Q(
        \I_cache/cache[1][73] ), .QN(n2070) );
  DFFRX1 \I_cache/cache_reg[2][73]  ( .D(n12201), .CK(clk), .RN(n5791), .Q(
        \I_cache/cache[2][73] ), .QN(n1482) );
  DFFRX1 \I_cache/cache_reg[3][73]  ( .D(n12200), .CK(clk), .RN(n5791), .Q(
        \I_cache/cache[3][73] ), .QN(n3056) );
  DFFRX1 \I_cache/cache_reg[4][73]  ( .D(n12199), .CK(clk), .RN(n5791), .Q(
        \I_cache/cache[4][73] ), .QN(n630) );
  DFFRX1 \I_cache/cache_reg[5][73]  ( .D(n12198), .CK(clk), .RN(n5790), .Q(
        \I_cache/cache[5][73] ), .QN(n2983) );
  DFFRX1 \I_cache/cache_reg[6][73]  ( .D(n12197), .CK(clk), .RN(n5790), .Q(
        \I_cache/cache[6][73] ), .QN(n1483) );
  DFFRX1 \I_cache/cache_reg[7][73]  ( .D(n12196), .CK(clk), .RN(n5790), .Q(
        \I_cache/cache[7][73] ), .QN(n3057) );
  DFFRX1 \I_cache/cache_reg[0][74]  ( .D(n12195), .CK(clk), .RN(n5790), .Q(
        \I_cache/cache[0][74] ), .QN(n1591) );
  DFFRX1 \I_cache/cache_reg[1][74]  ( .D(n12194), .CK(clk), .RN(n5790), .Q(
        \I_cache/cache[1][74] ), .QN(n3169) );
  DFFRX1 \I_cache/cache_reg[2][74]  ( .D(n12193), .CK(clk), .RN(n5790), .Q(
        \I_cache/cache[2][74] ), .QN(n1590) );
  DFFRX1 \I_cache/cache_reg[3][74]  ( .D(n12192), .CK(clk), .RN(n5790), .Q(
        \I_cache/cache[3][74] ), .QN(n3168) );
  DFFRX1 \I_cache/cache_reg[4][74]  ( .D(n12191), .CK(clk), .RN(n5790), .Q(
        \I_cache/cache[4][74] ), .QN(n1633) );
  DFFRX1 \I_cache/cache_reg[5][74]  ( .D(n12190), .CK(clk), .RN(n5790), .Q(
        \I_cache/cache[5][74] ), .QN(n3319) );
  DFFRX1 \I_cache/cache_reg[6][74]  ( .D(n12189), .CK(clk), .RN(n5790), .Q(
        \I_cache/cache[6][74] ), .QN(n1592) );
  DFFRX1 \I_cache/cache_reg[7][74]  ( .D(n12188), .CK(clk), .RN(n5790), .Q(
        \I_cache/cache[7][74] ), .QN(n3170) );
  DFFRX1 \I_cache/cache_reg[0][75]  ( .D(n12187), .CK(clk), .RN(n5790), .Q(
        \I_cache/cache[0][75] ), .QN(n1089) );
  DFFRX1 \I_cache/cache_reg[1][75]  ( .D(n12186), .CK(clk), .RN(n5789), .Q(
        \I_cache/cache[1][75] ), .QN(n2732) );
  DFFRX1 \I_cache/cache_reg[2][75]  ( .D(n12185), .CK(clk), .RN(n5789), .Q(
        \I_cache/cache[2][75] ), .QN(n1088) );
  DFFRX1 \I_cache/cache_reg[3][75]  ( .D(n12184), .CK(clk), .RN(n5789), .Q(
        \I_cache/cache[3][75] ), .QN(n2731) );
  DFFRX1 \I_cache/cache_reg[4][75]  ( .D(n12183), .CK(clk), .RN(n5789), .Q(
        \I_cache/cache[4][75] ), .QN(n688) );
  DFFRX1 \I_cache/cache_reg[5][75]  ( .D(n12182), .CK(clk), .RN(n5789), .Q(
        \I_cache/cache[5][75] ), .QN(n2299) );
  DFFRX1 \I_cache/cache_reg[6][75]  ( .D(n12181), .CK(clk), .RN(n5789), .Q(
        \I_cache/cache[6][75] ), .QN(n1090) );
  DFFRX1 \I_cache/cache_reg[7][75]  ( .D(n12180), .CK(clk), .RN(n5789), .Q(
        \I_cache/cache[7][75] ), .QN(n2733) );
  DFFRX1 \I_cache/cache_reg[0][76]  ( .D(n12179), .CK(clk), .RN(n5789), .Q(
        \I_cache/cache[0][76] ), .QN(n698) );
  DFFRX1 \I_cache/cache_reg[1][76]  ( .D(n12178), .CK(clk), .RN(n5789), .Q(
        \I_cache/cache[1][76] ), .QN(n2267) );
  DFFRX1 \I_cache/cache_reg[2][76]  ( .D(n12177), .CK(clk), .RN(n5789), .Q(
        \I_cache/cache[2][76] ), .QN(n1094) );
  DFFRX1 \I_cache/cache_reg[3][76]  ( .D(n12176), .CK(clk), .RN(n5789), .Q(
        \I_cache/cache[3][76] ), .QN(n2685) );
  DFFRX1 \I_cache/cache_reg[4][76]  ( .D(n12175), .CK(clk), .RN(n5789), .Q(
        \I_cache/cache[4][76] ), .QN(n1166) );
  DFFRX1 \I_cache/cache_reg[5][76]  ( .D(n12174), .CK(clk), .RN(n5788), .Q(
        \I_cache/cache[5][76] ), .QN(n2722) );
  DFFRX1 \I_cache/cache_reg[6][76]  ( .D(n12173), .CK(clk), .RN(n5788), .Q(
        \I_cache/cache[6][76] ), .QN(n1095) );
  DFFRX1 \I_cache/cache_reg[7][76]  ( .D(n12172), .CK(clk), .RN(n5788), .Q(
        \I_cache/cache[7][76] ), .QN(n2686) );
  DFFRX1 \I_cache/cache_reg[0][77]  ( .D(n12171), .CK(clk), .RN(n5788), .Q(
        \I_cache/cache[0][77] ), .QN(n1588) );
  DFFRX1 \I_cache/cache_reg[1][77]  ( .D(n12170), .CK(clk), .RN(n5788), .Q(
        \I_cache/cache[1][77] ), .QN(n3282) );
  DFFRX1 \I_cache/cache_reg[2][77]  ( .D(n12169), .CK(clk), .RN(n5788), .Q(
        \I_cache/cache[2][77] ), .QN(n1587) );
  DFFRX1 \I_cache/cache_reg[3][77]  ( .D(n12168), .CK(clk), .RN(n5788), .Q(
        \I_cache/cache[3][77] ), .QN(n3281) );
  DFFRX1 \I_cache/cache_reg[4][77]  ( .D(n12167), .CK(clk), .RN(n5788), .Q(
        \I_cache/cache[4][77] ), .QN(n629) );
  DFFRX1 \I_cache/cache_reg[5][77]  ( .D(n12166), .CK(clk), .RN(n5788), .Q(
        \I_cache/cache[5][77] ), .QN(n2981) );
  DFFRX1 \I_cache/cache_reg[6][77]  ( .D(n12165), .CK(clk), .RN(n5788), .Q(
        \I_cache/cache[6][77] ), .QN(n1688) );
  DFFRX1 \I_cache/cache_reg[7][77]  ( .D(n12164), .CK(clk), .RN(n5788), .Q(
        \I_cache/cache[7][77] ), .QN(n3283) );
  DFFRX1 \I_cache/cache_reg[0][78]  ( .D(n12163), .CK(clk), .RN(n5788), .Q(
        \I_cache/cache[0][78] ), .QN(n3062) );
  DFFRX1 \I_cache/cache_reg[1][78]  ( .D(n12162), .CK(clk), .RN(n5787), .Q(
        \I_cache/cache[1][78] ), .QN(n1171) );
  DFFRX1 \I_cache/cache_reg[2][78]  ( .D(n12161), .CK(clk), .RN(n5787), .Q(
        \I_cache/cache[2][78] ), .QN(n3061) );
  DFFRX1 \I_cache/cache_reg[3][78]  ( .D(n12160), .CK(clk), .RN(n5787), .Q(
        \I_cache/cache[3][78] ), .QN(n1170) );
  DFFRX1 \I_cache/cache_reg[4][78]  ( .D(n12159), .CK(clk), .RN(n5787), .Q(
        \I_cache/cache[4][78] ), .QN(n1167) );
  DFFRX1 \I_cache/cache_reg[5][78]  ( .D(n12158), .CK(clk), .RN(n5787), .Q(
        \I_cache/cache[5][78] ), .QN(n2723) );
  DFFRX1 \I_cache/cache_reg[6][78]  ( .D(n12157), .CK(clk), .RN(n5787), .Q(
        \I_cache/cache[6][78] ), .QN(n3063) );
  DFFRX1 \I_cache/cache_reg[7][78]  ( .D(n12156), .CK(clk), .RN(n5787), .Q(
        \I_cache/cache[7][78] ), .QN(n1172) );
  DFFRX1 \I_cache/cache_reg[7][91]  ( .D(n12052), .CK(clk), .RN(n5798), .Q(
        \I_cache/cache[7][91] ), .QN(n3122) );
  DFFRX1 \I_cache/cache_reg[0][92]  ( .D(n12051), .CK(clk), .RN(n5798), .Q(
        \I_cache/cache[0][92] ), .QN(n1106) );
  DFFRX1 \I_cache/cache_reg[2][92]  ( .D(n12049), .CK(clk), .RN(n5798), .Q(
        \I_cache/cache[2][92] ), .QN(n1108) );
  DFFRX1 \I_cache/cache_reg[3][92]  ( .D(n12048), .CK(clk), .RN(n5798), .Q(
        \I_cache/cache[3][92] ), .QN(n2697) );
  DFFRX1 \I_cache/cache_reg[4][92]  ( .D(n12047), .CK(clk), .RN(n5798), .Q(
        \I_cache/cache[4][92] ), .QN(n1107) );
  DFFRX1 \I_cache/cache_reg[5][92]  ( .D(n12046), .CK(clk), .RN(n5798), .Q(
        \I_cache/cache[5][92] ), .QN(n2696) );
  DFFRX1 \I_cache/cache_reg[6][92]  ( .D(n12045), .CK(clk), .RN(n5798), .Q(
        \I_cache/cache[6][92] ), .QN(n3077) );
  DFFRX1 \I_cache/cache_reg[7][92]  ( .D(n12044), .CK(clk), .RN(n5797), .Q(
        \I_cache/cache[7][92] ), .QN(n1187) );
  DFFRX1 \I_cache/cache_reg[0][93]  ( .D(n12043), .CK(clk), .RN(n5797), .Q(
        \I_cache/cache[0][93] ), .QN(n1518) );
  DFFRX1 \I_cache/cache_reg[1][93]  ( .D(n12042), .CK(clk), .RN(n5797), .Q(
        \I_cache/cache[1][93] ), .QN(n3098) );
  DFFRX1 \I_cache/cache_reg[2][93]  ( .D(n12041), .CK(clk), .RN(n5797), .Q(
        \I_cache/cache[2][93] ), .QN(n1517) );
  DFFRX1 \I_cache/cache_reg[3][93]  ( .D(n12040), .CK(clk), .RN(n5797), .Q(
        \I_cache/cache[3][93] ), .QN(n3097) );
  DFFRX1 \I_cache/cache_reg[4][93]  ( .D(n12039), .CK(clk), .RN(n5797), .Q(
        \I_cache/cache[4][93] ), .QN(n3076) );
  DFFRX1 \I_cache/cache_reg[5][93]  ( .D(n12038), .CK(clk), .RN(n5797), .Q(
        \I_cache/cache[5][93] ), .QN(n1186) );
  DFFRX1 \I_cache/cache_reg[6][93]  ( .D(n12037), .CK(clk), .RN(n5797), .Q(
        \I_cache/cache[6][93] ), .QN(n1519) );
  DFFRX1 \I_cache/cache_reg[7][93]  ( .D(n12036), .CK(clk), .RN(n5797), .Q(
        \I_cache/cache[7][93] ), .QN(n3099) );
  DFFRX1 \I_cache/cache_reg[2][94]  ( .D(n12033), .CK(clk), .RN(n5797), .Q(
        \I_cache/cache[2][94] ), .QN(n1576) );
  DFFRX1 \I_cache/cache_reg[3][94]  ( .D(n12032), .CK(clk), .RN(n5796), .Q(
        \I_cache/cache[3][94] ), .QN(n3158) );
  DFFRX1 \I_cache/cache_reg[4][94]  ( .D(n12031), .CK(clk), .RN(n5796), .Q(
        \I_cache/cache[4][94] ), .QN(n1597) );
  DFFRX1 \I_cache/cache_reg[5][94]  ( .D(n12030), .CK(clk), .RN(n5796), .Q(
        \I_cache/cache[5][94] ), .QN(n3174) );
  DFFRX1 \I_cache/cache_reg[6][94]  ( .D(n12029), .CK(clk), .RN(n5796), .Q(
        \I_cache/cache[6][94] ), .QN(n1575) );
  DFFRX1 \I_cache/cache_reg[7][94]  ( .D(n12028), .CK(clk), .RN(n5801), .Q(
        \I_cache/cache[7][94] ), .QN(n3157) );
  DFFRX1 \I_cache/cache_reg[1][95]  ( .D(n12026), .CK(clk), .RN(n5856), .Q(
        \I_cache/cache[1][95] ), .QN(n3133) );
  DFFRX1 \I_cache/cache_reg[3][95]  ( .D(n12024), .CK(clk), .RN(n5856), .Q(
        \I_cache/cache[3][95] ), .QN(n3132) );
  DFFRX1 \I_cache/cache_reg[4][95]  ( .D(n12023), .CK(clk), .RN(n5856), .Q(
        \I_cache/cache[4][95] ), .QN(n1601) );
  DFFRX1 \I_cache/cache_reg[5][95]  ( .D(n12022), .CK(clk), .RN(n5866), .Q(
        \I_cache/cache[5][95] ), .QN(n3178) );
  DFFRX1 \I_cache/cache_reg[6][95]  ( .D(n12021), .CK(clk), .RN(n5856), .Q(
        \I_cache/cache[6][95] ), .QN(n1552) );
  DFFRX1 \I_cache/cache_reg[7][95]  ( .D(n12020), .CK(clk), .RN(n5856), .Q(
        \I_cache/cache[7][95] ), .QN(n3134) );
  DFFRX1 \I_cache/cache_reg[0][96]  ( .D(n12019), .CK(clk), .RN(n5855), .Q(
        \I_cache/cache[0][96] ), .QN(n1660) );
  DFFRX1 \I_cache/cache_reg[1][96]  ( .D(n12018), .CK(clk), .RN(n5855), .Q(
        \I_cache/cache[1][96] ), .QN(n3244) );
  DFFRX1 \I_cache/cache_reg[2][96]  ( .D(n12017), .CK(clk), .RN(n5855), .Q(
        \I_cache/cache[2][96] ), .QN(n1662) );
  DFFRX1 \I_cache/cache_reg[3][96]  ( .D(n12016), .CK(clk), .RN(n5855), .Q(
        \I_cache/cache[3][96] ), .QN(n3246) );
  DFFRX1 \I_cache/cache_reg[4][96]  ( .D(n12015), .CK(clk), .RN(n5855), .Q(
        \I_cache/cache[4][96] ), .QN(n1661) );
  DFFRX1 \I_cache/cache_reg[5][96]  ( .D(n12014), .CK(clk), .RN(n5855), .Q(
        \I_cache/cache[5][96] ), .QN(n3245) );
  DFFRX1 \I_cache/cache_reg[6][96]  ( .D(n12013), .CK(clk), .RN(n5855), .Q(
        \I_cache/cache[6][96] ), .QN(n1458) );
  DFFRX1 \I_cache/cache_reg[7][96]  ( .D(n12012), .CK(clk), .RN(n5855), .Q(
        \I_cache/cache[7][96] ), .QN(n3032) );
  DFFRX1 \I_cache/cache_reg[0][97]  ( .D(n12011), .CK(clk), .RN(n5855), .Q(
        \I_cache/cache[0][97] ), .QN(n1663) );
  DFFRX1 \I_cache/cache_reg[1][97]  ( .D(n12010), .CK(clk), .RN(n5855), .Q(
        \I_cache/cache[1][97] ), .QN(n3247) );
  DFFRX1 \I_cache/cache_reg[2][97]  ( .D(n12009), .CK(clk), .RN(n5855), .Q(
        \I_cache/cache[2][97] ), .QN(n1471) );
  DFFRX1 \I_cache/cache_reg[3][97]  ( .D(n12008), .CK(clk), .RN(n5855), .Q(
        \I_cache/cache[3][97] ), .QN(n3045) );
  DFFRX1 \I_cache/cache_reg[4][97]  ( .D(n12007), .CK(clk), .RN(n5854), .Q(
        \I_cache/cache[4][97] ), .QN(n1472) );
  DFFRX1 \I_cache/cache_reg[5][97]  ( .D(n12006), .CK(clk), .RN(n5854), .Q(
        \I_cache/cache[5][97] ), .QN(n3046) );
  DFFRX1 \I_cache/cache_reg[6][97]  ( .D(n12005), .CK(clk), .RN(n5854), .Q(
        \I_cache/cache[6][97] ), .QN(n1477) );
  DFFRX1 \I_cache/cache_reg[7][97]  ( .D(n12004), .CK(clk), .RN(n5854), .Q(
        \I_cache/cache[7][97] ), .QN(n3051) );
  DFFRX1 \I_cache/cache_reg[0][98]  ( .D(n12003), .CK(clk), .RN(n5854), .Q(
        \I_cache/cache[0][98] ), .QN(n1489) );
  DFFRX1 \I_cache/cache_reg[1][98]  ( .D(n12002), .CK(clk), .RN(n5854), .Q(
        \I_cache/cache[1][98] ), .QN(n3073) );
  DFFRX1 \I_cache/cache_reg[2][98]  ( .D(n12001), .CK(clk), .RN(n5854), .Q(
        \I_cache/cache[2][98] ), .QN(n2740) );
  DFFRX1 \I_cache/cache_reg[3][98]  ( .D(n12000), .CK(clk), .RN(n5854), .Q(
        \I_cache/cache[3][98] ), .QN(n1280) );
  DFFRX1 \I_cache/cache_reg[4][98]  ( .D(n11999), .CK(clk), .RN(n5854), .Q(
        \I_cache/cache[4][98] ), .QN(n1486) );
  DFFRX1 \I_cache/cache_reg[5][98]  ( .D(n11998), .CK(clk), .RN(n5854), .Q(
        \I_cache/cache[5][98] ), .QN(n3069) );
  DFFRX1 \I_cache/cache_reg[6][98]  ( .D(n11997), .CK(clk), .RN(n5854), .Q(
        \I_cache/cache[6][98] ), .QN(n1487) );
  DFFRX1 \I_cache/cache_reg[7][98]  ( .D(n11996), .CK(clk), .RN(n5854), .Q(
        \I_cache/cache[7][98] ), .QN(n3070) );
  DFFRX1 \I_cache/cache_reg[2][99]  ( .D(n11993), .CK(clk), .RN(n5853), .Q(
        \I_cache/cache[2][99] ), .QN(n1448) );
  DFFRX1 \I_cache/cache_reg[3][99]  ( .D(n11992), .CK(clk), .RN(n5853), .Q(
        \I_cache/cache[3][99] ), .QN(n3019) );
  DFFRX1 \I_cache/cache_reg[4][99]  ( .D(n11991), .CK(clk), .RN(n5853), .Q(
        \I_cache/cache[4][99] ), .QN(n1580) );
  DFFRX1 \I_cache/cache_reg[5][99]  ( .D(n11990), .CK(clk), .RN(n5853), .Q(
        \I_cache/cache[5][99] ), .QN(n3162) );
  DFFRX1 \I_cache/cache_reg[6][99]  ( .D(n11989), .CK(clk), .RN(n5853), .Q(
        \I_cache/cache[6][99] ), .QN(n1450) );
  DFFRX1 \I_cache/cache_reg[7][99]  ( .D(n11988), .CK(clk), .RN(n5853), .Q(
        \I_cache/cache[7][99] ), .QN(n3021) );
  DFFRX1 \I_cache/cache_reg[0][100]  ( .D(n11987), .CK(clk), .RN(n5853), .Q(
        \I_cache/cache[0][100] ), .QN(n2992) );
  DFFRX1 \I_cache/cache_reg[1][100]  ( .D(n11986), .CK(clk), .RN(n5853), .Q(
        \I_cache/cache[1][100] ), .QN(n1434) );
  DFFRX1 \I_cache/cache_reg[2][100]  ( .D(n11985), .CK(clk), .RN(n5853), .Q(
        \I_cache/cache[2][100] ), .QN(n1468) );
  DFFRX1 \I_cache/cache_reg[3][100]  ( .D(n11984), .CK(clk), .RN(n5853), .Q(
        \I_cache/cache[3][100] ), .QN(n3042) );
  DFFRX1 \I_cache/cache_reg[4][100]  ( .D(n11983), .CK(clk), .RN(n5852), .Q(
        \I_cache/cache[4][100] ), .QN(n1676) );
  DFFRX1 \I_cache/cache_reg[5][100]  ( .D(n11982), .CK(clk), .RN(n5852), .Q(
        \I_cache/cache[5][100] ), .QN(n3264) );
  DFFRX1 \I_cache/cache_reg[6][100]  ( .D(n11981), .CK(clk), .RN(n5852), .Q(
        \I_cache/cache[6][100] ), .QN(n1654) );
  DFFRX1 \I_cache/cache_reg[7][100]  ( .D(n11980), .CK(clk), .RN(n5852), .Q(
        \I_cache/cache[7][100] ), .QN(n3238) );
  DFFRX1 \I_cache/cache_reg[0][101]  ( .D(n11979), .CK(clk), .RN(n5852), .Q(
        \I_cache/cache[0][101] ), .QN(n2743) );
  DFFRX1 \I_cache/cache_reg[1][101]  ( .D(n11978), .CK(clk), .RN(n5852), .Q(
        \I_cache/cache[1][101] ), .QN(n1283) );
  DFFRX1 \I_cache/cache_reg[2][101]  ( .D(n11977), .CK(clk), .RN(n5852), .Q(
        \I_cache/cache[2][101] ), .QN(n1510) );
  DFFRX1 \I_cache/cache_reg[3][101]  ( .D(n11976), .CK(clk), .RN(n5852), .Q(
        \I_cache/cache[3][101] ), .QN(n3090) );
  DFFRX1 \I_cache/cache_reg[4][101]  ( .D(n11975), .CK(clk), .RN(n5852), .Q(
        \I_cache/cache[4][101] ), .QN(n1509) );
  DFFRX1 \I_cache/cache_reg[5][101]  ( .D(n11974), .CK(clk), .RN(n5852), .Q(
        \I_cache/cache[5][101] ), .QN(n3089) );
  DFFRX1 \I_cache/cache_reg[6][101]  ( .D(n11973), .CK(clk), .RN(n5852), .Q(
        \I_cache/cache[6][101] ), .QN(n1595) );
  DFFRX1 \I_cache/cache_reg[7][101]  ( .D(n11972), .CK(clk), .RN(n5852), .Q(
        \I_cache/cache[7][101] ), .QN(n3172) );
  DFFRX1 \I_cache/cache_reg[0][102]  ( .D(n11971), .CK(clk), .RN(n5851), .Q(
        \I_cache/cache[0][102] ), .QN(n1699) );
  DFFRX1 \I_cache/cache_reg[1][102]  ( .D(n11970), .CK(clk), .RN(n5851), .Q(
        \I_cache/cache[1][102] ), .QN(n3295) );
  DFFRX1 \I_cache/cache_reg[2][102]  ( .D(n11969), .CK(clk), .RN(n5851), .Q(
        \I_cache/cache[2][102] ), .QN(n1698) );
  DFFRX1 \I_cache/cache_reg[3][102]  ( .D(n11968), .CK(clk), .RN(n5851), .Q(
        \I_cache/cache[3][102] ), .QN(n3294) );
  DFFRX1 \I_cache/cache_reg[4][102]  ( .D(n11967), .CK(clk), .RN(n5851), .Q(
        \I_cache/cache[4][102] ), .QN(n750) );
  DFFRX1 \I_cache/cache_reg[5][102]  ( .D(n11966), .CK(clk), .RN(n5851), .Q(
        \I_cache/cache[5][102] ), .QN(n2311) );
  DFFRX1 \I_cache/cache_reg[6][102]  ( .D(n11965), .CK(clk), .RN(n5851), .Q(
        \I_cache/cache[6][102] ), .QN(n1700) );
  DFFRX1 \I_cache/cache_reg[7][102]  ( .D(n11964), .CK(clk), .RN(n5851), .Q(
        \I_cache/cache[7][102] ), .QN(n3296) );
  DFFRX1 \I_cache/cache_reg[0][103]  ( .D(n11963), .CK(clk), .RN(n5851), .Q(
        \I_cache/cache[0][103] ), .QN(n1647) );
  DFFRX1 \I_cache/cache_reg[1][103]  ( .D(n11962), .CK(clk), .RN(n5851), .Q(
        \I_cache/cache[1][103] ), .QN(n3229) );
  DFFRX1 \I_cache/cache_reg[2][103]  ( .D(n11961), .CK(clk), .RN(n5851), .Q(
        \I_cache/cache[2][103] ), .QN(n1463) );
  DFFRX1 \I_cache/cache_reg[3][103]  ( .D(n11960), .CK(clk), .RN(n5850), .Q(
        \I_cache/cache[3][103] ), .QN(n3037) );
  DFFRX1 \I_cache/cache_reg[4][103]  ( .D(n11959), .CK(clk), .RN(n5850), .Q(
        \I_cache/cache[4][103] ), .QN(n1218) );
  DFFRX1 \I_cache/cache_reg[5][103]  ( .D(n11958), .CK(clk), .RN(n5850), .Q(
        \I_cache/cache[5][103] ), .QN(n2755) );
  DFFRX1 \I_cache/cache_reg[6][103]  ( .D(n11957), .CK(clk), .RN(n5850), .Q(
        \I_cache/cache[6][103] ), .QN(n1466) );
  DFFRX1 \I_cache/cache_reg[7][103]  ( .D(n11956), .CK(clk), .RN(n5850), .Q(
        \I_cache/cache[7][103] ), .QN(n3040) );
  DFFRX1 \I_cache/cache_reg[0][104]  ( .D(n11955), .CK(clk), .RN(n5850), .Q(
        \I_cache/cache[0][104] ), .QN(n1697) );
  DFFRX1 \I_cache/cache_reg[1][104]  ( .D(n11954), .CK(clk), .RN(n5850), .Q(
        \I_cache/cache[1][104] ), .QN(n3293) );
  DFFRX1 \I_cache/cache_reg[2][104]  ( .D(n11953), .CK(clk), .RN(n5850), .Q(
        \I_cache/cache[2][104] ), .QN(n1465) );
  DFFRX1 \I_cache/cache_reg[3][104]  ( .D(n11952), .CK(clk), .RN(n5850), .Q(
        \I_cache/cache[3][104] ), .QN(n3039) );
  DFFRX1 \I_cache/cache_reg[4][104]  ( .D(n11951), .CK(clk), .RN(n5850), .Q(
        \I_cache/cache[4][104] ), .QN(n1209) );
  DFFRX1 \I_cache/cache_reg[5][104]  ( .D(n11950), .CK(clk), .RN(n5850), .Q(
        \I_cache/cache[5][104] ), .QN(n2746) );
  DFFRX1 \I_cache/cache_reg[6][104]  ( .D(n11949), .CK(clk), .RN(n5850), .Q(
        \I_cache/cache[6][104] ), .QN(n1637) );
  DFFRX1 \I_cache/cache_reg[7][104]  ( .D(n11948), .CK(clk), .RN(n5849), .Q(
        \I_cache/cache[7][104] ), .QN(n3219) );
  DFFRX1 \I_cache/cache_reg[0][105]  ( .D(n11947), .CK(clk), .RN(n5849), .Q(
        \I_cache/cache[0][105] ), .QN(n1694) );
  DFFRX1 \I_cache/cache_reg[1][105]  ( .D(n11946), .CK(clk), .RN(n5849), .Q(
        \I_cache/cache[1][105] ), .QN(n3290) );
  DFFRX1 \I_cache/cache_reg[2][105]  ( .D(n11945), .CK(clk), .RN(n5849), .Q(
        \I_cache/cache[2][105] ), .QN(n1693) );
  DFFRX1 \I_cache/cache_reg[3][105]  ( .D(n11944), .CK(clk), .RN(n5849), .Q(
        \I_cache/cache[3][105] ), .QN(n3289) );
  DFFRX1 \I_cache/cache_reg[4][105]  ( .D(n11943), .CK(clk), .RN(n5849), .Q(
        \I_cache/cache[4][105] ), .QN(n1384) );
  DFFRX1 \I_cache/cache_reg[5][105]  ( .D(n11942), .CK(clk), .RN(n5849), .Q(
        \I_cache/cache[5][105] ), .QN(n2914) );
  DFFRX1 \I_cache/cache_reg[6][105]  ( .D(n11941), .CK(clk), .RN(n5849), .Q(
        \I_cache/cache[6][105] ), .QN(n1695) );
  DFFRX1 \I_cache/cache_reg[7][105]  ( .D(n11940), .CK(clk), .RN(n5849), .Q(
        \I_cache/cache[7][105] ), .QN(n3291) );
  DFFRX1 \I_cache/cache_reg[0][106]  ( .D(n11939), .CK(clk), .RN(n5849), .Q(
        \I_cache/cache[0][106] ), .QN(n1497) );
  DFFRX1 \I_cache/cache_reg[1][106]  ( .D(n11938), .CK(clk), .RN(n5849), .Q(
        \I_cache/cache[1][106] ), .QN(n3258) );
  DFFRX1 \I_cache/cache_reg[2][106]  ( .D(n11937), .CK(clk), .RN(n5849), .Q(
        \I_cache/cache[2][106] ), .QN(n1496) );
  DFFRX1 \I_cache/cache_reg[3][106]  ( .D(n11936), .CK(clk), .RN(n5848), .Q(
        \I_cache/cache[3][106] ), .QN(n3257) );
  DFFRX1 \I_cache/cache_reg[4][106]  ( .D(n11935), .CK(clk), .RN(n5848), .Q(
        \I_cache/cache[4][106] ), .QN(n1476) );
  DFFRX1 \I_cache/cache_reg[5][106]  ( .D(n11934), .CK(clk), .RN(n5848), .Q(
        \I_cache/cache[5][106] ), .QN(n3050) );
  DFFRX1 \I_cache/cache_reg[6][106]  ( .D(n11933), .CK(clk), .RN(n5848), .Q(
        \I_cache/cache[6][106] ), .QN(n1498) );
  DFFRX1 \I_cache/cache_reg[7][106]  ( .D(n11932), .CK(clk), .RN(n5848), .Q(
        \I_cache/cache[7][106] ), .QN(n3259) );
  DFFRX1 \I_cache/cache_reg[0][107]  ( .D(n11931), .CK(clk), .RN(n5848), .Q(
        \I_cache/cache[0][107] ), .QN(n3066) );
  DFFRX1 \I_cache/cache_reg[1][107]  ( .D(n11930), .CK(clk), .RN(n5848), .Q(
        \I_cache/cache[1][107] ), .QN(n1174) );
  DFFRX1 \I_cache/cache_reg[2][107]  ( .D(n11929), .CK(clk), .RN(n5848), .Q(
        \I_cache/cache[2][107] ), .QN(n3065) );
  DFFRX1 \I_cache/cache_reg[3][107]  ( .D(n11928), .CK(clk), .RN(n5848), .Q(
        \I_cache/cache[3][107] ), .QN(n1277) );
  DFFRX1 \I_cache/cache_reg[4][107]  ( .D(n11927), .CK(clk), .RN(n5848), .Q(
        \I_cache/cache[4][107] ), .QN(n3018) );
  DFFRX1 \I_cache/cache_reg[5][107]  ( .D(n11926), .CK(clk), .RN(n5848), .Q(
        \I_cache/cache[5][107] ), .QN(n845) );
  DFFRX1 \I_cache/cache_reg[6][107]  ( .D(n11925), .CK(clk), .RN(n5848), .Q(
        \I_cache/cache[6][107] ), .QN(n1097) );
  DFFRX1 \I_cache/cache_reg[7][107]  ( .D(n11924), .CK(clk), .RN(n5847), .Q(
        \I_cache/cache[7][107] ), .QN(n2736) );
  DFFRX1 \I_cache/cache_reg[0][108]  ( .D(n11923), .CK(clk), .RN(n5847), .Q(
        \I_cache/cache[0][108] ), .QN(n1099) );
  DFFRX1 \I_cache/cache_reg[1][108]  ( .D(n11922), .CK(clk), .RN(n5847), .Q(
        \I_cache/cache[1][108] ), .QN(n2688) );
  DFFRX1 \I_cache/cache_reg[2][108]  ( .D(n11921), .CK(clk), .RN(n5847), .Q(
        \I_cache/cache[2][108] ), .QN(n1098) );
  DFFRX1 \I_cache/cache_reg[3][108]  ( .D(n11920), .CK(clk), .RN(n5847), .Q(
        \I_cache/cache[3][108] ), .QN(n2687) );
  DFFRX1 \I_cache/cache_reg[4][108]  ( .D(n11919), .CK(clk), .RN(n5847), .Q(
        \I_cache/cache[4][108] ), .QN(n1168) );
  DFFRX1 \I_cache/cache_reg[5][108]  ( .D(n11918), .CK(clk), .RN(n5847), .Q(
        \I_cache/cache[5][108] ), .QN(n2724) );
  DFFRX1 \I_cache/cache_reg[6][108]  ( .D(n11917), .CK(clk), .RN(n5847), .Q(
        \I_cache/cache[6][108] ), .QN(n1100) );
  DFFRX1 \I_cache/cache_reg[7][108]  ( .D(n11916), .CK(clk), .RN(n5847), .Q(
        \I_cache/cache[7][108] ), .QN(n2689) );
  DFFRX1 \I_cache/cache_reg[0][109]  ( .D(n11915), .CK(clk), .RN(n5847), .Q(
        \I_cache/cache[0][109] ), .QN(n1583) );
  DFFRX1 \I_cache/cache_reg[1][109]  ( .D(n11914), .CK(clk), .RN(n5847), .Q(
        \I_cache/cache[1][109] ), .QN(n3163) );
  DFFRX1 \I_cache/cache_reg[2][109]  ( .D(n11913), .CK(clk), .RN(n5847), .Q(
        \I_cache/cache[2][109] ), .QN(n1582) );
  DFFRX1 \I_cache/cache_reg[3][109]  ( .D(n11912), .CK(clk), .RN(n5846), .Q(
        \I_cache/cache[3][109] ), .QN(n3276) );
  DFFRX1 \I_cache/cache_reg[4][109]  ( .D(n11911), .CK(clk), .RN(n5846), .Q(
        \I_cache/cache[4][109] ), .QN(n2134) );
  DFFRX1 \I_cache/cache_reg[5][109]  ( .D(n11910), .CK(clk), .RN(n5846), .Q(
        \I_cache/cache[5][109] ), .QN(n549) );
  DFFRX1 \I_cache/cache_reg[6][109]  ( .D(n11909), .CK(clk), .RN(n5846), .Q(
        \I_cache/cache[6][109] ), .QN(n1581) );
  DFFRX1 \I_cache/cache_reg[7][109]  ( .D(n11908), .CK(clk), .RN(n5846), .Q(
        \I_cache/cache[7][109] ), .QN(n3275) );
  DFFRX1 \I_cache/cache_reg[0][110]  ( .D(n11907), .CK(clk), .RN(n5846), .Q(
        \I_cache/cache[0][110] ), .QN(n1502) );
  DFFRX1 \I_cache/cache_reg[1][110]  ( .D(n11906), .CK(clk), .RN(n5851), .Q(
        \I_cache/cache[1][110] ), .QN(n3082) );
  DFFRX1 \I_cache/cache_reg[2][110]  ( .D(n11905), .CK(clk), .RN(n5866), .Q(
        \I_cache/cache[2][110] ), .QN(n1501) );
  DFFRX1 \I_cache/cache_reg[3][110]  ( .D(n11904), .CK(clk), .RN(n5866), .Q(
        \I_cache/cache[3][110] ), .QN(n3081) );
  DFFRX1 \I_cache/cache_reg[4][110]  ( .D(n11903), .CK(clk), .RN(n5866), .Q(
        \I_cache/cache[4][110] ), .QN(n1586) );
  DFFRX1 \I_cache/cache_reg[5][110]  ( .D(n11902), .CK(clk), .RN(n5866), .Q(
        \I_cache/cache[5][110] ), .QN(n3166) );
  DFFRX1 \I_cache/cache_reg[6][110]  ( .D(n11901), .CK(clk), .RN(n5866), .Q(
        \I_cache/cache[6][110] ), .QN(n1503) );
  DFFRX1 \I_cache/cache_reg[7][110]  ( .D(n11900), .CK(clk), .RN(n5865), .Q(
        \I_cache/cache[7][110] ), .QN(n3083) );
  DFFRX1 \I_cache/cache_reg[0][124]  ( .D(n11795), .CK(clk), .RN(n5857), .Q(
        \I_cache/cache[0][124] ), .QN(n3016) );
  DFFRX1 \I_cache/cache_reg[1][124]  ( .D(n11794), .CK(clk), .RN(n5857), .Q(
        \I_cache/cache[1][124] ), .QN(n722) );
  DFFRX1 \I_cache/cache_reg[2][124]  ( .D(n11793), .CK(clk), .RN(n5856), .Q(
        \I_cache/cache[2][124] ), .QN(n1105) );
  DFFRX1 \I_cache/cache_reg[3][124]  ( .D(n11792), .CK(clk), .RN(n5856), .Q(
        \I_cache/cache[3][124] ), .QN(n2694) );
  DFFRX1 \I_cache/cache_reg[4][124]  ( .D(n11791), .CK(clk), .RN(n5856), .Q(
        \I_cache/cache[4][124] ), .QN(n1104) );
  DFFRX1 \I_cache/cache_reg[5][124]  ( .D(n11790), .CK(clk), .RN(n5856), .Q(
        \I_cache/cache[5][124] ), .QN(n2693) );
  DFFRX1 \I_cache/cache_reg[6][124]  ( .D(n11789), .CK(clk), .RN(n5856), .Q(
        \I_cache/cache[6][124] ), .QN(n1086) );
  DFFRX1 \I_cache/cache_reg[7][124]  ( .D(n11788), .CK(clk), .RN(n5856), .Q(
        \I_cache/cache[7][124] ), .QN(n2680) );
  DFFRX1 \I_cache/cache_reg[0][125]  ( .D(n11787), .CK(clk), .RN(n5861), .Q(
        \I_cache/cache[0][125] ), .QN(n1512) );
  DFFRX1 \I_cache/cache_reg[1][125]  ( .D(n11786), .CK(clk), .RN(n5836), .Q(
        \I_cache/cache[1][125] ), .QN(n3092) );
  DFFRX1 \I_cache/cache_reg[2][125]  ( .D(n11785), .CK(clk), .RN(n5836), .Q(
        \I_cache/cache[2][125] ), .QN(n1511) );
  DFFRX1 \I_cache/cache_reg[3][125]  ( .D(n11784), .CK(clk), .RN(n5836), .Q(
        \I_cache/cache[3][125] ), .QN(n3091) );
  DFFRX1 \I_cache/cache_reg[4][125]  ( .D(n11783), .CK(clk), .RN(n5836), .Q(
        \I_cache/cache[4][125] ), .QN(n3060) );
  DFFRX1 \I_cache/cache_reg[5][125]  ( .D(n11782), .CK(clk), .RN(n5836), .Q(
        \I_cache/cache[5][125] ), .QN(n1150) );
  DFFRX1 \I_cache/cache_reg[6][125]  ( .D(n11781), .CK(clk), .RN(n5836), .Q(
        \I_cache/cache[6][125] ), .QN(n1513) );
  DFFRX1 \I_cache/cache_reg[7][125]  ( .D(n11780), .CK(clk), .RN(n5835), .Q(
        \I_cache/cache[7][125] ), .QN(n3093) );
  DFFRX1 \I_cache/cache_reg[1][126]  ( .D(n11778), .CK(clk), .RN(n5835), .Q(
        \I_cache/cache[1][126] ), .QN(n3104) );
  DFFRX1 \I_cache/cache_reg[2][126]  ( .D(n11777), .CK(clk), .RN(n5835), .Q(
        \I_cache/cache[2][126] ), .QN(n1523) );
  DFFRX1 \I_cache/cache_reg[3][126]  ( .D(n11776), .CK(clk), .RN(n5835), .Q(
        \I_cache/cache[3][126] ), .QN(n3103) );
  DFFRX1 \I_cache/cache_reg[4][126]  ( .D(n11775), .CK(clk), .RN(n5835), .Q(
        \I_cache/cache[4][126] ), .QN(n3074) );
  DFFRX1 \I_cache/cache_reg[5][126]  ( .D(n11774), .CK(clk), .RN(n5835), .Q(
        \I_cache/cache[5][126] ), .QN(n1184) );
  DFFRX1 \I_cache/cache_reg[6][126]  ( .D(n11773), .CK(clk), .RN(n5835), .Q(
        \I_cache/cache[6][126] ), .QN(n1525) );
  DFFRX1 \I_cache/cache_reg[1][127]  ( .D(n11770), .CK(clk), .RN(n5835), .Q(
        \I_cache/cache[1][127] ), .QN(n3127) );
  DFFRX1 \I_cache/cache_reg[3][127]  ( .D(n11768), .CK(clk), .RN(n5834), .Q(
        \I_cache/cache[3][127] ), .QN(n3126) );
  DFFRX1 \I_cache/cache_reg[5][127]  ( .D(n11766), .CK(clk), .RN(n5834), .Q(
        \I_cache/cache[5][127] ), .QN(n3179) );
  DFFRX1 \I_cache/cache_reg[6][127]  ( .D(n11765), .CK(clk), .RN(n5834), .Q(
        \I_cache/cache[6][127] ), .QN(n1546) );
  DFFRX1 \I_cache/cache_reg[7][127]  ( .D(n11764), .CK(clk), .RN(n5834), .Q(
        \I_cache/cache[7][127] ), .QN(n3128) );
  DFFRX1 \I_cache/cache_reg[0][130]  ( .D(n11747), .CK(clk), .RN(n5833), .Q(
        \I_cache/cache[0][130] ), .QN(n740) );
  DFFRX1 \I_cache/cache_reg[0][145]  ( .D(n11627), .CK(clk), .RN(n5843), .Q(
        \I_cache/cache[0][145] ), .QN(n1251) );
  DFFRX1 \I_cache/cache_reg[0][143]  ( .D(n11643), .CK(clk), .RN(n5844), .Q(
        \I_cache/cache[0][143] ), .QN(n2173) );
  DFFRX1 \I_cache/cache_reg[4][141]  ( .D(n11655), .CK(clk), .RN(n5845), .Q(
        \I_cache/cache[4][141] ), .QN(n2181) );
  DFFRX1 \I_cache/cache_reg[2][142]  ( .D(n11649), .CK(clk), .RN(n5844), .Q(
        \I_cache/cache[2][142] ), .QN(n2177) );
  DFFRX1 \I_cache/cache_reg[0][129]  ( .D(n11755), .CK(clk), .RN(n5833), .Q(
        \I_cache/cache[0][129] ), .QN(n2182) );
  DFFRX1 \I_cache/cache_reg[2][146]  ( .D(n11617), .CK(clk), .RN(n5842), .Q(
        \I_cache/cache[2][146] ), .QN(n2186) );
  DFFRX1 \I_cache/cache_reg[1][141]  ( .D(n11658), .CK(clk), .RN(n5845), .Q(
        \I_cache/cache[1][141] ), .QN(n605) );
  DFFRX1 \I_cache/cache_reg[6][141]  ( .D(n11653), .CK(clk), .RN(n5845), .Q(
        \I_cache/cache[6][141] ), .QN(n794) );
  DFFRX1 \I_cache/cache_reg[0][131]  ( .D(n11739), .CK(clk), .RN(n5832), .Q(
        \I_cache/cache[0][131] ), .QN(n1234) );
  DFFRX1 \I_cache/cache_reg[0][150]  ( .D(n11587), .CK(clk), .RN(n5839), .Q(
        \I_cache/cache[0][150] ), .QN(n1400) );
  DFFRX1 \I_cache/cache_reg[2][130]  ( .D(n11745), .CK(clk), .RN(n5833), .Q(
        \I_cache/cache[2][130] ), .QN(n1236) );
  DFFRX1 \I_cache/cache_reg[2][143]  ( .D(n11641), .CK(clk), .RN(n5844), .Q(
        \I_cache/cache[2][143] ), .QN(n2174) );
  DFFRX1 \I_cache/cache_reg[4][142]  ( .D(n11647), .CK(clk), .RN(n5844), .Q(
        \I_cache/cache[4][142] ), .QN(n2178) );
  DFFRX1 \I_cache/cache_reg[4][146]  ( .D(n11615), .CK(clk), .RN(n5842), .Q(
        \I_cache/cache[4][146] ), .QN(n2187) );
  DFFRX1 \I_cache/cache_reg[0][147]  ( .D(n11611), .CK(clk), .RN(n5841), .Q(
        \I_cache/cache[0][147] ), .QN(n1397) );
  DFFRX1 \I_cache/cache_reg[2][145]  ( .D(n11625), .CK(clk), .RN(n5842), .Q(
        \I_cache/cache[2][145] ), .QN(n1252) );
  DFFRX1 \I_cache/cache_reg[2][129]  ( .D(n11753), .CK(clk), .RN(n5833), .Q(
        \I_cache/cache[2][129] ), .QN(n2183) );
  DFFRX1 \I_cache/cache_reg[1][146]  ( .D(n11618), .CK(clk), .RN(n5842), .Q(
        \I_cache/cache[1][146] ), .QN(n611) );
  DFFRX1 \I_cache/cache_reg[1][142]  ( .D(n11650), .CK(clk), .RN(n5845), .Q(
        \I_cache/cache[1][142] ), .QN(n602) );
  DFFRX1 \I_cache/cache_reg[6][142]  ( .D(n11645), .CK(clk), .RN(n5844), .Q(
        \I_cache/cache[6][142] ), .QN(n793) );
  DFFRX1 \I_cache/cache_reg[3][141]  ( .D(n11656), .CK(clk), .RN(n5845), .Q(
        \I_cache/cache[3][141] ), .QN(n606) );
  DFFRX1 \I_cache/cache_reg[6][146]  ( .D(n11613), .CK(clk), .RN(n5841), .Q(
        \I_cache/cache[6][146] ), .QN(n2151) );
  DFFRX1 \I_cache/cache_reg[2][131]  ( .D(n11737), .CK(clk), .RN(n5832), .Q(
        \I_cache/cache[2][131] ), .QN(n1235) );
  DFFRX1 \I_cache/cache_reg[4][130]  ( .D(n11743), .CK(clk), .RN(n5832), .Q(
        \I_cache/cache[4][130] ), .QN(n1237) );
  DFFRX1 \I_cache/cache_reg[4][143]  ( .D(n11639), .CK(clk), .RN(n5844), .Q(
        \I_cache/cache[4][143] ), .QN(n2175) );
  DFFRX1 \I_cache/cache_reg[4][129]  ( .D(n11751), .CK(clk), .RN(n5833), .Q(
        \I_cache/cache[4][129] ), .QN(n2184) );
  DFFRX1 \I_cache/cache_reg[1][130]  ( .D(n11746), .CK(clk), .RN(n5833), .Q(
        \I_cache/cache[1][130] ), .QN(n2301) );
  DFFRX1 \I_cache/cache_reg[6][130]  ( .D(n11741), .CK(clk), .RN(n5832), .Q(
        \I_cache/cache[6][130] ), .QN(n788) );
  DFFRX1 \I_cache/cache_reg[6][145]  ( .D(n11621), .CK(clk), .RN(n5842), .Q(
        \I_cache/cache[6][145] ), .QN(n785) );
  DFFRX1 \I_cache/cache_reg[2][150]  ( .D(n11585), .CK(clk), .RN(n5839), .Q(
        \I_cache/cache[2][150] ), .QN(n1401) );
  DFFRX1 \I_cache/cache_reg[0][149]  ( .D(n11595), .CK(clk), .RN(n5840), .Q(
        \I_cache/cache[0][149] ), .QN(n1228) );
  DFFRX1 \I_cache/cache_reg[1][143]  ( .D(n11642), .CK(clk), .RN(n5844), .Q(
        \I_cache/cache[1][143] ), .QN(n599) );
  DFFRX1 \I_cache/cache_reg[0][134]  ( .D(n11715), .CK(clk), .RN(n5830), .Q(
        \I_cache/cache[0][134] ), .QN(n2170) );
  DFFRX1 \I_cache/cache_reg[6][143]  ( .D(n11637), .CK(clk), .RN(n5843), .Q(
        \I_cache/cache[6][143] ), .QN(n792) );
  DFFRX1 \I_cache/cache_reg[4][145]  ( .D(n11623), .CK(clk), .RN(n5842), .Q(
        \I_cache/cache[4][145] ), .QN(n742) );
  DFFRX1 \I_cache/cache_reg[1][129]  ( .D(n11754), .CK(clk), .RN(n5833), .Q(
        \I_cache/cache[1][129] ), .QN(n608) );
  DFFRX1 \I_cache/cache_reg[4][131]  ( .D(n11735), .CK(clk), .RN(n5832), .Q(
        \I_cache/cache[4][131] ), .QN(n770) );
  DFFRX1 \I_cache/cache_reg[0][151]  ( .D(n11579), .CK(clk), .RN(n5839), .Q(
        \I_cache/cache[0][151] ), .QN(n1417) );
  DFFRX1 \I_cache/cache_reg[2][147]  ( .D(n11609), .CK(clk), .RN(n5841), .Q(
        \I_cache/cache[2][147] ), .QN(n1398) );
  DFFRX1 \I_cache/cache_reg[6][129]  ( .D(n11749), .CK(clk), .RN(n5833), .Q(
        \I_cache/cache[6][129] ), .QN(n786) );
  DFFRX1 \I_cache/cache_reg[3][146]  ( .D(n11616), .CK(clk), .RN(n5842), .Q(
        \I_cache/cache[3][146] ), .QN(n612) );
  DFFRX1 \I_cache/cache_reg[3][142]  ( .D(n11648), .CK(clk), .RN(n5844), .Q(
        \I_cache/cache[3][142] ), .QN(n603) );
  DFFRX1 \I_cache/cache_reg[5][141]  ( .D(n11654), .CK(clk), .RN(n5845), .Q(
        \I_cache/cache[5][141] ), .QN(n607) );
  DFFRX1 \I_cache/cache_reg[1][145]  ( .D(n11626), .CK(clk), .RN(n5843), .Q(
        \I_cache/cache[1][145] ), .QN(n2793) );
  DFFRX1 \I_cache/cache_reg[1][131]  ( .D(n11738), .CK(clk), .RN(n5832), .Q(
        \I_cache/cache[1][131] ), .QN(n2775) );
  DFFRX1 \I_cache/cache_reg[6][150]  ( .D(n11581), .CK(clk), .RN(n5839), .Q(
        \I_cache/cache[6][150] ), .QN(n1389) );
  DFFRX1 \I_cache/cache_reg[6][131]  ( .D(n11733), .CK(clk), .RN(n5832), .Q(
        \I_cache/cache[6][131] ), .QN(n787) );
  DFFRX1 \I_cache/cache_reg[0][144]  ( .D(n11635), .CK(clk), .RN(n5843), .Q(
        \I_cache/cache[0][144] ), .QN(n1415) );
  DFFRX1 \I_cache/cache_reg[0][128]  ( .D(n11763), .CK(clk), .RN(n5834), .Q(
        \I_cache/cache[0][128] ), .QN(n649) );
  DFFRX1 \I_cache/cache_reg[0][137]  ( .D(n11691), .CK(clk), .RN(n5828), .Q(
        \I_cache/cache[0][137] ), .QN(n1409) );
  DFFRX1 \I_cache/cache_reg[6][147]  ( .D(n11605), .CK(clk), .RN(n5841), .Q(
        \I_cache/cache[6][147] ), .QN(n1388) );
  DFFRX1 \I_cache/cache_reg[2][134]  ( .D(n11713), .CK(clk), .RN(n5830), .Q(
        \I_cache/cache[2][134] ), .QN(n2171) );
  DFFRX1 \I_cache/cache_reg[0][135]  ( .D(n11707), .CK(clk), .RN(n5829), .Q(
        \I_cache/cache[0][135] ), .QN(n1238) );
  DFFRX1 \I_cache/cache_reg[4][150]  ( .D(n11583), .CK(clk), .RN(n5839), .Q(
        \I_cache/cache[4][150] ), .QN(n1402) );
  DFFRX1 \I_cache/cache_reg[3][130]  ( .D(n11744), .CK(clk), .RN(n5833), .Q(
        \I_cache/cache[3][130] ), .QN(n2777) );
  DFFRX1 \I_cache/cache_reg[3][143]  ( .D(n11640), .CK(clk), .RN(n5844), .Q(
        \I_cache/cache[3][143] ), .QN(n600) );
  DFFRX1 \I_cache/cache_reg[0][133]  ( .D(n11723), .CK(clk), .RN(n5831), .Q(
        \I_cache/cache[0][133] ), .QN(n1240) );
  DFFRX1 \I_cache/cache_reg[2][151]  ( .D(n11577), .CK(clk), .RN(n5838), .Q(
        \I_cache/cache[2][151] ), .QN(n1289) );
  DFFRX1 \I_cache/cache_reg[2][149]  ( .D(n11593), .CK(clk), .RN(n5840), .Q(
        \I_cache/cache[2][149] ), .QN(n1395) );
  DFFRX1 \I_cache/cache_reg[4][147]  ( .D(n11607), .CK(clk), .RN(n5841), .Q(
        \I_cache/cache[4][147] ), .QN(n1399) );
  DFFRX1 \I_cache/cache_reg[3][129]  ( .D(n11752), .CK(clk), .RN(n5833), .Q(
        \I_cache/cache[3][129] ), .QN(n609) );
  DFFRX1 \I_cache/cache_reg[5][146]  ( .D(n11614), .CK(clk), .RN(n5842), .Q(
        \I_cache/cache[5][146] ), .QN(n613) );
  DFFRX1 \I_cache/cache_reg[5][142]  ( .D(n11646), .CK(clk), .RN(n5844), .Q(
        \I_cache/cache[5][142] ), .QN(n604) );
  DFFRX1 \I_cache/cache_reg[7][141]  ( .D(n11652), .CK(clk), .RN(n5845), .Q(
        \I_cache/cache[7][141] ), .QN(n2356) );
  DFFRX1 \I_cache/cache_reg[1][150]  ( .D(n11586), .CK(clk), .RN(n5839), .Q(
        \I_cache/cache[1][150] ), .QN(n2931) );
  DFFRX1 \I_cache/cache_reg[6][149]  ( .D(n11589), .CK(clk), .RN(n5839), .Q(
        \I_cache/cache[6][149] ), .QN(n1390) );
  DFFRX1 \I_cache/cache_reg[2][144]  ( .D(n11633), .CK(clk), .RN(n5843), .Q(
        \I_cache/cache[2][144] ), .QN(n1416) );
  DFFRX1 \I_cache/cache_reg[4][134]  ( .D(n11711), .CK(clk), .RN(n5830), .Q(
        \I_cache/cache[4][134] ), .QN(n2172) );
  DFFRX1 \I_cache/cache_reg[2][128]  ( .D(n11761), .CK(clk), .RN(n5834), .Q(
        \I_cache/cache[2][128] ), .QN(n1243) );
  DFFRX1 \I_cache/cache_reg[3][131]  ( .D(n11736), .CK(clk), .RN(n5832), .Q(
        \I_cache/cache[3][131] ), .QN(n2776) );
  DFFRX1 \I_cache/cache_reg[0][138]  ( .D(n11683), .CK(clk), .RN(n5827), .Q(
        \I_cache/cache[0][138] ), .QN(n1253) );
  DFFRX1 \I_cache/cache_reg[1][147]  ( .D(n11610), .CK(clk), .RN(n5841), .Q(
        \I_cache/cache[1][147] ), .QN(n2928) );
  DFFRX1 \I_cache/cache_reg[0][139]  ( .D(n11675), .CK(clk), .RN(n5827), .Q(
        \I_cache/cache[0][139] ), .QN(n1413) );
  DFFRX1 \I_cache/cache_reg[2][137]  ( .D(n11689), .CK(clk), .RN(n5828), .Q(
        \I_cache/cache[2][137] ), .QN(n1410) );
  DFFRX1 \I_cache/cache_reg[0][136]  ( .D(n11699), .CK(clk), .RN(n5829), .Q(
        \I_cache/cache[0][136] ), .QN(n1406) );
  DFFRX1 \I_cache/cache_reg[2][135]  ( .D(n11705), .CK(clk), .RN(n5829), .Q(
        \I_cache/cache[2][135] ), .QN(n1239) );
  DFFRX1 \I_cache/cache_reg[4][151]  ( .D(n11575), .CK(clk), .RN(n5838), .Q(
        \I_cache/cache[4][151] ), .QN(n2137) );
  DFFRX1 \I_cache/cache_reg[1][134]  ( .D(n11714), .CK(clk), .RN(n5830), .Q(
        \I_cache/cache[1][134] ), .QN(n596) );
  DFFRX1 \I_cache/cache_reg[2][133]  ( .D(n11721), .CK(clk), .RN(n5831), .Q(
        \I_cache/cache[2][133] ), .QN(n1241) );
  DFFRX1 \I_cache/cache_reg[0][132]  ( .D(n11731), .CK(clk), .RN(n5831), .Q(
        \I_cache/cache[0][132] ), .QN(n776) );
  DFFRX1 \I_cache/cache_reg[3][145]  ( .D(n11624), .CK(clk), .RN(n5842), .Q(
        \I_cache/cache[3][145] ), .QN(n2794) );
  DFFRX1 \I_cache/cache_reg[5][143]  ( .D(n11638), .CK(clk), .RN(n5844), .Q(
        \I_cache/cache[5][143] ), .QN(n601) );
  DFFRX1 \I_cache/cache_reg[5][130]  ( .D(n11742), .CK(clk), .RN(n5832), .Q(
        \I_cache/cache[5][130] ), .QN(n2778) );
  DFFRX1 \I_cache/cache_reg[6][134]  ( .D(n11709), .CK(clk), .RN(n5830), .Q(
        \I_cache/cache[6][134] ), .QN(n791) );
  DFFRX1 \I_cache/cache_reg[4][149]  ( .D(n11591), .CK(clk), .RN(n5840), .Q(
        \I_cache/cache[4][149] ), .QN(n1396) );
  DFFRX1 \I_cache/cache_reg[1][151]  ( .D(n11578), .CK(clk), .RN(n5838), .Q(
        \I_cache/cache[1][151] ), .QN(n2948) );
  DFFRX1 \I_cache/cache_reg[5][129]  ( .D(n11750), .CK(clk), .RN(n5833), .Q(
        \I_cache/cache[5][129] ), .QN(n610) );
  DFFRX1 \I_cache/cache_reg[4][144]  ( .D(n11631), .CK(clk), .RN(n5843), .Q(
        \I_cache/cache[4][144] ), .QN(n2159) );
  DFFRX1 \I_cache/cache_reg[7][146]  ( .D(n11612), .CK(clk), .RN(n5841), .Q(
        \I_cache/cache[7][146] ), .QN(n572) );
  DFFRX1 \I_cache/cache_reg[7][142]  ( .D(n11644), .CK(clk), .RN(n5844), .Q(
        \I_cache/cache[7][142] ), .QN(n2355) );
  DFFRX1 \I_cache/cache_reg[4][128]  ( .D(n11759), .CK(clk), .RN(n5834), .Q(
        \I_cache/cache[4][128] ), .QN(n2158) );
  DFFRX1 \I_cache/cache_reg[6][151]  ( .D(n11573), .CK(clk), .RN(n5838), .Q(
        \I_cache/cache[6][151] ), .QN(n1385) );
  DFFRX1 \I_cache/cache_reg[4][137]  ( .D(n11687), .CK(clk), .RN(n5828), .Q(
        \I_cache/cache[4][137] ), .QN(n1411) );
  DFFRX1 \I_cache/cache_reg[4][135]  ( .D(n11703), .CK(clk), .RN(n5829), .Q(
        \I_cache/cache[4][135] ), .QN(n777) );
  DFFRX1 \I_cache/cache_reg[2][138]  ( .D(n11681), .CK(clk), .RN(n5827), .Q(
        \I_cache/cache[2][138] ), .QN(n1254) );
  DFFRX1 \I_cache/cache_reg[1][149]  ( .D(n11594), .CK(clk), .RN(n5840), .Q(
        \I_cache/cache[1][149] ), .QN(n2765) );
  DFFRX1 \I_cache/cache_reg[2][139]  ( .D(n11673), .CK(clk), .RN(n5827), .Q(
        \I_cache/cache[2][139] ), .QN(n1414) );
  DFFRX1 \I_cache/cache_reg[0][148]  ( .D(n11603), .CK(clk), .RN(n5841), .Q(
        \I_cache/cache[0][148] ), .QN(n1403) );
  DFFRX1 \I_cache/cache_reg[1][144]  ( .D(n11634), .CK(clk), .RN(n5843), .Q(
        \I_cache/cache[1][144] ), .QN(n2946) );
  DFFRX1 \I_cache/cache_reg[0][140]  ( .D(n11667), .CK(clk), .RN(n5831), .Q(
        \I_cache/cache[0][140] ), .QN(n1210) );
  DFFRX1 \I_cache/cache_reg[1][128]  ( .D(n11762), .CK(clk), .RN(n5834), .Q(
        \I_cache/cache[1][128] ), .QN(n2226) );
  DFFRX1 \I_cache/cache_reg[2][136]  ( .D(n11697), .CK(clk), .RN(n5829), .Q(
        \I_cache/cache[2][136] ), .QN(n1407) );
  DFFRX1 \I_cache/cache_reg[4][133]  ( .D(n11719), .CK(clk), .RN(n5830), .Q(
        \I_cache/cache[4][133] ), .QN(n2168) );
  DFFRX1 \I_cache/cache_reg[7][130]  ( .D(n11740), .CK(clk), .RN(n5832), .Q(
        \I_cache/cache[7][130] ), .QN(n2350) );
  DFFRX1 \I_cache/cache_reg[5][131]  ( .D(n11734), .CK(clk), .RN(n5832), .Q(
        \I_cache/cache[5][131] ), .QN(n2332) );
  DFFRX1 \I_cache/cache_reg[3][150]  ( .D(n11584), .CK(clk), .RN(n5839), .Q(
        \I_cache/cache[3][150] ), .QN(n2932) );
  DFFRX1 \I_cache/cache_reg[6][144]  ( .D(n11629), .CK(clk), .RN(n5843), .Q(
        \I_cache/cache[6][144] ), .QN(n1276) );
  DFFRX1 \I_cache/cache_reg[7][145]  ( .D(n11620), .CK(clk), .RN(n5842), .Q(
        \I_cache/cache[7][145] ), .QN(n2347) );
  DFFRX1 \I_cache/cache_reg[1][137]  ( .D(n11690), .CK(clk), .RN(n5828), .Q(
        \I_cache/cache[1][137] ), .QN(n2940) );
  DFFRX1 \I_cache/cache_reg[6][128]  ( .D(n11757), .CK(clk), .RN(n5834), .Q(
        \I_cache/cache[6][128] ), .QN(n1305) );
  DFFRX1 \I_cache/cache_reg[1][135]  ( .D(n11706), .CK(clk), .RN(n5829), .Q(
        \I_cache/cache[1][135] ), .QN(n2779) );
  DFFRX1 \I_cache/cache_reg[2][132]  ( .D(n11729), .CK(clk), .RN(n5831), .Q(
        \I_cache/cache[2][132] ), .QN(n1242) );
  DFFRX1 \I_cache/cache_reg[3][134]  ( .D(n11712), .CK(clk), .RN(n5830), .Q(
        \I_cache/cache[3][134] ), .QN(n597) );
  DFFRX1 \I_cache/cache_reg[6][137]  ( .D(n11685), .CK(clk), .RN(n5828), .Q(
        \I_cache/cache[6][137] ), .QN(n1227) );
  DFFRX1 \I_cache/cache_reg[7][143]  ( .D(n11636), .CK(clk), .RN(n5843), .Q(
        \I_cache/cache[7][143] ), .QN(n2354) );
  DFFRX1 \I_cache/cache_reg[1][133]  ( .D(n11722), .CK(clk), .RN(n5831), .Q(
        \I_cache/cache[1][133] ), .QN(n2781) );
  DFFRX1 \I_cache/cache_reg[6][135]  ( .D(n11701), .CK(clk), .RN(n5829), .Q(
        \I_cache/cache[6][135] ), .QN(n1275) );
  DFFRX1 \I_cache/cache_reg[3][147]  ( .D(n11608), .CK(clk), .RN(n5841), .Q(
        \I_cache/cache[3][147] ), .QN(n2929) );
  DFFRX1 \I_cache/cache_reg[6][133]  ( .D(n11717), .CK(clk), .RN(n5830), .Q(
        \I_cache/cache[6][133] ), .QN(n790) );
  DFFRX1 \I_cache/cache_reg[7][129]  ( .D(n11748), .CK(clk), .RN(n5833), .Q(
        \I_cache/cache[7][129] ), .QN(n2348) );
  DFFRX1 \I_cache/cache_reg[3][151]  ( .D(n11576), .CK(clk), .RN(n5838), .Q(
        \I_cache/cache[3][151] ), .QN(n2822) );
  DFFRX1 \I_cache/cache_reg[4][138]  ( .D(n11679), .CK(clk), .RN(n5827), .Q(
        \I_cache/cache[4][138] ), .QN(n1255) );
  DFFRX1 \I_cache/cache_reg[4][139]  ( .D(n11671), .CK(clk), .RN(n5826), .Q(
        \I_cache/cache[4][139] ), .QN(n2157) );
  DFFRX1 \I_cache/cache_reg[4][136]  ( .D(n11695), .CK(clk), .RN(n5828), .Q(
        \I_cache/cache[4][136] ), .QN(n1408) );
  DFFRX1 \I_cache/cache_reg[5][145]  ( .D(n11622), .CK(clk), .RN(n5842), .Q(
        \I_cache/cache[5][145] ), .QN(n2303) );
  DFFRX1 \I_cache/cache_reg[7][131]  ( .D(n11732), .CK(clk), .RN(n5832), .Q(
        \I_cache/cache[7][131] ), .QN(n2349) );
  DFFRX1 \I_cache/cache_reg[7][150]  ( .D(n11580), .CK(clk), .RN(n5839), .Q(
        \I_cache/cache[7][150] ), .QN(n2919) );
  DFFRX1 \I_cache/cache_reg[0][152]  ( .D(n11571), .CK(clk), .RN(n5838), .Q(
        \I_cache/cache[0][152] ), .QN(n1135) );
  DFFRX1 \I_cache/cache_reg[2][148]  ( .D(n11601), .CK(clk), .RN(n5840), .Q(
        \I_cache/cache[2][148] ), .QN(n1404) );
  DFFRX1 \I_cache/cache_reg[2][140]  ( .D(n11665), .CK(clk), .RN(n5846), .Q(
        \I_cache/cache[2][140] ), .QN(n1412) );
  DFFRX1 \I_cache/cache_reg[4][132]  ( .D(n11727), .CK(clk), .RN(n5831), .Q(
        \I_cache/cache[4][132] ), .QN(n2169) );
  DFFRX1 \I_cache/cache_reg[3][144]  ( .D(n11632), .CK(clk), .RN(n5843), .Q(
        \I_cache/cache[3][144] ), .QN(n2947) );
  DFFRX1 \I_cache/cache_reg[3][128]  ( .D(n11760), .CK(clk), .RN(n5834), .Q(
        \I_cache/cache[3][128] ), .QN(n2784) );
  DFFRX1 \I_cache/cache_reg[1][138]  ( .D(n11682), .CK(clk), .RN(n5827), .Q(
        \I_cache/cache[1][138] ), .QN(n2795) );
  DFFRX1 \I_cache/cache_reg[1][139]  ( .D(n11674), .CK(clk), .RN(n5827), .Q(
        \I_cache/cache[1][139] ), .QN(n2944) );
  DFFRX1 \I_cache/cache_reg[7][147]  ( .D(n11604), .CK(clk), .RN(n5841), .Q(
        \I_cache/cache[7][147] ), .QN(n2918) );
  DFFRX1 \I_cache/cache_reg[1][136]  ( .D(n11698), .CK(clk), .RN(n5829), .Q(
        \I_cache/cache[1][136] ), .QN(n2937) );
  DFFRX1 \I_cache/cache_reg[6][138]  ( .D(n11677), .CK(clk), .RN(n5827), .Q(
        \I_cache/cache[6][138] ), .QN(n789) );
  DFFRX1 \I_cache/cache_reg[3][137]  ( .D(n11688), .CK(clk), .RN(n5828), .Q(
        \I_cache/cache[3][137] ), .QN(n2941) );
  DFFRX1 \I_cache/cache_reg[6][139]  ( .D(n11669), .CK(clk), .RN(n5826), .Q(
        \I_cache/cache[6][139] ), .QN(n1274) );
  DFFRX1 \I_cache/cache_reg[3][135]  ( .D(n11704), .CK(clk), .RN(n5829), .Q(
        \I_cache/cache[3][135] ), .QN(n2780) );
  DFFRX1 \I_cache/cache_reg[6][136]  ( .D(n11693), .CK(clk), .RN(n5828), .Q(
        \I_cache/cache[6][136] ), .QN(n1386) );
  DFFRX1 \I_cache/cache_reg[1][132]  ( .D(n11730), .CK(clk), .RN(n5831), .Q(
        \I_cache/cache[1][132] ), .QN(n2338) );
  DFFRX1 \I_cache/cache_reg[5][134]  ( .D(n11710), .CK(clk), .RN(n5830), .Q(
        \I_cache/cache[5][134] ), .QN(n598) );
  DFFRX1 \I_cache/cache_reg[3][149]  ( .D(n11592), .CK(clk), .RN(n5840), .Q(
        \I_cache/cache[3][149] ), .QN(n2926) );
  DFFRX1 \I_cache/cache_reg[3][133]  ( .D(n11720), .CK(clk), .RN(n5830), .Q(
        \I_cache/cache[3][133] ), .QN(n2782) );
  DFFRX1 \I_cache/cache_reg[6][132]  ( .D(n11725), .CK(clk), .RN(n5831), .Q(
        \I_cache/cache[6][132] ), .QN(n2101) );
  DFFRX1 \I_cache/cache_reg[5][150]  ( .D(n11582), .CK(clk), .RN(n5839), .Q(
        \I_cache/cache[5][150] ), .QN(n2933) );
  DFFRX1 \I_cache/cache_reg[4][148]  ( .D(n11599), .CK(clk), .RN(n5840), .Q(
        \I_cache/cache[4][148] ), .QN(n1405) );
  DFFRX1 \I_cache/cache_reg[4][140]  ( .D(n11663), .CK(clk), .RN(n5846), .Q(
        \I_cache/cache[4][140] ), .QN(n2156) );
  DFFRX1 \I_cache/cache_reg[5][151]  ( .D(n11574), .CK(clk), .RN(n5838), .Q(
        \I_cache/cache[5][151] ), .QN(n552) );
  DFFRX1 \I_cache/cache_reg[7][149]  ( .D(n11588), .CK(clk), .RN(n5839), .Q(
        \I_cache/cache[7][149] ), .QN(n2920) );
  DFFRX1 \I_cache/cache_reg[2][152]  ( .D(n11569), .CK(clk), .RN(n5838), .Q(
        \I_cache/cache[2][152] ), .QN(n1136) );
  DFFRX1 \I_cache/cache_reg[5][147]  ( .D(n11606), .CK(clk), .RN(n5841), .Q(
        \I_cache/cache[5][147] ), .QN(n2930) );
  DFFRX1 \I_cache/cache_reg[1][148]  ( .D(n11602), .CK(clk), .RN(n5840), .Q(
        \I_cache/cache[1][148] ), .QN(n2934) );
  DFFRX1 \I_cache/cache_reg[1][140]  ( .D(n11666), .CK(clk), .RN(n5846), .Q(
        \I_cache/cache[1][140] ), .QN(n2747) );
  DFFRX1 \I_cache/cache_reg[5][144]  ( .D(n11630), .CK(clk), .RN(n5843), .Q(
        \I_cache/cache[5][144] ), .QN(n582) );
  DFFRX1 \I_cache/cache_reg[5][128]  ( .D(n11758), .CK(clk), .RN(n5834), .Q(
        \I_cache/cache[5][128] ), .QN(n581) );
  DFFRX1 \I_cache/cache_reg[3][138]  ( .D(n11680), .CK(clk), .RN(n5827), .Q(
        \I_cache/cache[3][138] ), .QN(n2796) );
  DFFRX1 \I_cache/cache_reg[3][139]  ( .D(n11672), .CK(clk), .RN(n5826), .Q(
        \I_cache/cache[3][139] ), .QN(n2945) );
  DFFRX1 \I_cache/cache_reg[6][148]  ( .D(n11597), .CK(clk), .RN(n5840), .Q(
        \I_cache/cache[6][148] ), .QN(n1387) );
  DFFRX1 \I_cache/cache_reg[3][136]  ( .D(n11696), .CK(clk), .RN(n5828), .Q(
        \I_cache/cache[3][136] ), .QN(n2938) );
  DFFRX1 \I_cache/cache_reg[6][140]  ( .D(n11661), .CK(clk), .RN(n5845), .Q(
        \I_cache/cache[6][140] ), .QN(n1273) );
  DFFRX1 \I_cache/cache_reg[5][137]  ( .D(n11686), .CK(clk), .RN(n5828), .Q(
        \I_cache/cache[5][137] ), .QN(n2942) );
  DFFRX1 \I_cache/cache_reg[5][135]  ( .D(n11702), .CK(clk), .RN(n5829), .Q(
        \I_cache/cache[5][135] ), .QN(n2339) );
  DFFRX1 \I_cache/cache_reg[3][132]  ( .D(n11728), .CK(clk), .RN(n5831), .Q(
        \I_cache/cache[3][132] ), .QN(n2783) );
  DFFRX1 \I_cache/cache_reg[7][134]  ( .D(n11708), .CK(clk), .RN(n5829), .Q(
        \I_cache/cache[7][134] ), .QN(n2353) );
  DFFRX1 \I_cache/cache_reg[5][133]  ( .D(n11718), .CK(clk), .RN(n5830), .Q(
        \I_cache/cache[5][133] ), .QN(n594) );
  DFFRX1 \I_cache/cache_reg[7][151]  ( .D(n11572), .CK(clk), .RN(n5838), .Q(
        \I_cache/cache[7][151] ), .QN(n2915) );
  DFFRX1 \I_cache/cache_reg[5][149]  ( .D(n11590), .CK(clk), .RN(n5839), .Q(
        \I_cache/cache[5][149] ), .QN(n2927) );
  DFFRX1 \I_cache/cache_reg[1][152]  ( .D(n11570), .CK(clk), .RN(n5838), .Q(
        \I_cache/cache[1][152] ), .QN(n2671) );
  DFFRX1 \I_cache/cache_reg[3][148]  ( .D(n11600), .CK(clk), .RN(n5840), .Q(
        \I_cache/cache[3][148] ), .QN(n2935) );
  DFFRX1 \I_cache/cache_reg[6][152]  ( .D(n11565), .CK(clk), .RN(n5837), .Q(
        \I_cache/cache[6][152] ), .QN(n1079) );
  DFFRX1 \I_cache/cache_reg[3][140]  ( .D(n11664), .CK(clk), .RN(n5846), .Q(
        \I_cache/cache[3][140] ), .QN(n2943) );
  DFFRX1 \I_cache/cache_reg[7][144]  ( .D(n11628), .CK(clk), .RN(n5843), .Q(
        \I_cache/cache[7][144] ), .QN(n2819) );
  DFFRX1 \I_cache/cache_reg[7][128]  ( .D(n11756), .CK(clk), .RN(n5837), .Q(
        \I_cache/cache[7][128] ), .QN(n2834) );
  DFFRX1 \I_cache/cache_reg[5][138]  ( .D(n11678), .CK(clk), .RN(n5827), .Q(
        \I_cache/cache[5][138] ), .QN(n2797) );
  DFFRX1 \I_cache/cache_reg[5][139]  ( .D(n11670), .CK(clk), .RN(n5826), .Q(
        \I_cache/cache[5][139] ), .QN(n580) );
  DFFRX1 \I_cache/cache_reg[5][136]  ( .D(n11694), .CK(clk), .RN(n5828), .Q(
        \I_cache/cache[5][136] ), .QN(n2939) );
  DFFRX1 \I_cache/cache_reg[7][137]  ( .D(n11684), .CK(clk), .RN(n5827), .Q(
        \I_cache/cache[7][137] ), .QN(n2764) );
  DFFRX1 \I_cache/cache_reg[7][135]  ( .D(n11700), .CK(clk), .RN(n5829), .Q(
        \I_cache/cache[7][135] ), .QN(n2818) );
  DFFRX1 \I_cache/cache_reg[5][132]  ( .D(n11726), .CK(clk), .RN(n5831), .Q(
        \I_cache/cache[5][132] ), .QN(n595) );
  DFFRX1 \I_cache/cache_reg[7][133]  ( .D(n11716), .CK(clk), .RN(n5830), .Q(
        \I_cache/cache[7][133] ), .QN(n2352) );
  DFFRX1 \I_cache/cache_reg[3][152]  ( .D(n11568), .CK(clk), .RN(n5838), .Q(
        \I_cache/cache[3][152] ), .QN(n2672) );
  DFFRX1 \I_cache/cache_reg[5][148]  ( .D(n11598), .CK(clk), .RN(n5840), .Q(
        \I_cache/cache[5][148] ), .QN(n2936) );
  DFFRX1 \I_cache/cache_reg[5][140]  ( .D(n11662), .CK(clk), .RN(n5846), .Q(
        \I_cache/cache[5][140] ), .QN(n579) );
  DFFRX1 \I_cache/cache_reg[7][138]  ( .D(n11676), .CK(clk), .RN(n5827), .Q(
        \I_cache/cache[7][138] ), .QN(n2351) );
  DFFRX1 \I_cache/cache_reg[7][139]  ( .D(n11668), .CK(clk), .RN(n5826), .Q(
        \I_cache/cache[7][139] ), .QN(n2817) );
  DFFRX1 \I_cache/cache_reg[7][136]  ( .D(n11692), .CK(clk), .RN(n5828), .Q(
        \I_cache/cache[7][136] ), .QN(n2916) );
  DFFRX1 \I_cache/cache_reg[7][132]  ( .D(n11724), .CK(clk), .RN(n5831), .Q(
        \I_cache/cache[7][132] ), .QN(n516) );
  DFFRX1 \I_cache/cache_reg[5][152]  ( .D(n11566), .CK(clk), .RN(n5837), .Q(
        \I_cache/cache[5][152] ), .QN(n485) );
  DFFRX1 \I_cache/cache_reg[7][148]  ( .D(n11596), .CK(clk), .RN(n5840), .Q(
        \I_cache/cache[7][148] ), .QN(n2917) );
  DFFRX1 \I_cache/cache_reg[7][140]  ( .D(n11660), .CK(clk), .RN(n5845), .Q(
        \I_cache/cache[7][140] ), .QN(n2816) );
  DFFRX1 \I_cache/cache_reg[7][152]  ( .D(n11564), .CK(clk), .RN(n5837), .Q(
        \I_cache/cache[7][152] ), .QN(n2657) );
  DFFRX1 \I_cache/cache_reg[6][15]  ( .D(n12661), .CK(clk), .RN(n5909), .Q(
        \I_cache/cache[6][15] ), .QN(n1481) );
  DFFRX1 \I_cache/cache_reg[7][15]  ( .D(n12660), .CK(clk), .RN(n5909), .Q(
        \I_cache/cache[7][15] ), .QN(n3055) );
  DFFRX1 \I_cache/cache_reg[0][47]  ( .D(n12411), .CK(clk), .RN(n5808), .Q(
        \I_cache/cache[0][47] ), .QN(n2984) );
  DFFRX1 \I_cache/cache_reg[1][47]  ( .D(n12410), .CK(clk), .RN(n5808), .Q(
        \I_cache/cache[1][47] ), .QN(n1428) );
  DFFRX1 \I_cache/cache_reg[2][47]  ( .D(n12409), .CK(clk), .RN(n5808), .Q(
        \I_cache/cache[2][47] ), .QN(n2985) );
  DFFRX1 \I_cache/cache_reg[3][47]  ( .D(n12408), .CK(clk), .RN(n5808), .Q(
        \I_cache/cache[3][47] ), .QN(n1429) );
  DFFRX1 \I_cache/cache_reg[4][47]  ( .D(n12407), .CK(clk), .RN(n5808), .Q(
        \I_cache/cache[4][47] ), .QN(n2993) );
  DFFRX1 \I_cache/cache_reg[5][47]  ( .D(n12406), .CK(clk), .RN(n5808), .Q(
        \I_cache/cache[5][47] ), .QN(n1435) );
  DFFRX1 \I_cache/cache_reg[6][47]  ( .D(n12405), .CK(clk), .RN(n5808), .Q(
        \I_cache/cache[6][47] ), .QN(n2163) );
  DFFRX1 \I_cache/cache_reg[7][47]  ( .D(n12404), .CK(clk), .RN(n5808), .Q(
        \I_cache/cache[7][47] ), .QN(n588) );
  DFFRX1 \I_cache/cache_reg[2][79]  ( .D(n12153), .CK(clk), .RN(n5787), .Q(
        \I_cache/cache[2][79] ), .QN(n2739) );
  DFFRX1 \I_cache/cache_reg[3][79]  ( .D(n12152), .CK(clk), .RN(n5787), .Q(
        \I_cache/cache[3][79] ), .QN(n1279) );
  DFFRX1 \I_cache/cache_reg[4][79]  ( .D(n12151), .CK(clk), .RN(n5787), .Q(
        \I_cache/cache[4][79] ), .QN(n1449) );
  DFFRX1 \I_cache/cache_reg[5][79]  ( .D(n12150), .CK(clk), .RN(n5786), .Q(
        \I_cache/cache[5][79] ), .QN(n3020) );
  DFFRX1 \I_cache/cache_reg[6][79]  ( .D(n12149), .CK(clk), .RN(n5786), .Q(
        \I_cache/cache[6][79] ), .QN(n701) );
  DFFRX1 \I_cache/cache_reg[7][79]  ( .D(n12148), .CK(clk), .RN(n5786), .Q(
        \I_cache/cache[7][79] ), .QN(n2270) );
  DFFRX1 \I_cache/cache_reg[4][111]  ( .D(n11895), .CK(clk), .RN(n5865), .Q(
        \I_cache/cache[4][111] ), .QN(n1480) );
  DFFRX1 \I_cache/cache_reg[5][111]  ( .D(n11894), .CK(clk), .RN(n5865), .Q(
        \I_cache/cache[5][111] ), .QN(n3054) );
  DFFRX1 \I_cache/cache_reg[0][141]  ( .D(n11659), .CK(clk), .RN(n5845), .Q(
        \I_cache/cache[0][141] ), .QN(n2179) );
  DFFRX1 \I_cache/cache_reg[2][141]  ( .D(n11657), .CK(clk), .RN(n5845), .Q(
        \I_cache/cache[2][141] ), .QN(n2180) );
  DFFRX1 \I_cache/cache_reg[0][142]  ( .D(n11651), .CK(clk), .RN(n5845), .Q(
        \I_cache/cache[0][142] ), .QN(n2176) );
  DFFRX1 \I_cache/cache_reg[0][146]  ( .D(n11619), .CK(clk), .RN(n5842), .Q(
        \I_cache/cache[0][146] ), .QN(n2185) );
  DFFRX1 \I_cache/cache_reg[6][153]  ( .D(n11557), .CK(clk), .RN(n5837), .Q(
        \I_cache/cache[6][153] ), .QN(n1634) );
  DFFRX1 \I_cache/cache_reg[7][153]  ( .D(n11556), .CK(clk), .RN(n5837), .Q(
        \I_cache/cache[7][153] ), .QN(n3214) );
  DFFRX1 \I_cache/cache_reg[0][15]  ( .D(n12667), .CK(clk), .RN(n5909), .Q(
        \I_cache/cache[0][15] ), .QN(n1484) );
  DFFRX1 \I_cache/cache_reg[1][15]  ( .D(n12666), .CK(clk), .RN(n5909), .Q(
        \I_cache/cache[1][15] ), .QN(n3058) );
  DFFRX1 \I_cache/cache_reg[2][15]  ( .D(n12665), .CK(clk), .RN(n5909), .Q(
        \I_cache/cache[2][15] ), .QN(n3031) );
  DFFRX1 \I_cache/cache_reg[3][15]  ( .D(n12664), .CK(clk), .RN(n5909), .Q(
        \I_cache/cache[3][15] ), .QN(n1447) );
  DFFRX1 \I_cache/cache_reg[4][15]  ( .D(n12663), .CK(clk), .RN(n5909), .Q(
        \I_cache/cache[4][15] ), .QN(n3010) );
  DFFRX1 \I_cache/cache_reg[5][15]  ( .D(n12662), .CK(clk), .RN(n5909), .Q(
        \I_cache/cache[5][15] ), .QN(n1442) );
  DFFRX1 \I_cache/cache_reg[0][111]  ( .D(n11899), .CK(clk), .RN(n5865), .Q(
        \I_cache/cache[0][111] ), .QN(n3011) );
  DFFRX1 \I_cache/cache_reg[1][111]  ( .D(n11898), .CK(clk), .RN(n5865), .Q(
        \I_cache/cache[1][111] ), .QN(n1443) );
  DFFRX1 \I_cache/cache_reg[2][111]  ( .D(n11897), .CK(clk), .RN(n5865), .Q(
        \I_cache/cache[2][111] ), .QN(n3012) );
  DFFRX1 \I_cache/cache_reg[3][111]  ( .D(n11896), .CK(clk), .RN(n5865), .Q(
        \I_cache/cache[3][111] ), .QN(n1444) );
  DFFRX1 \I_cache/cache_reg[6][111]  ( .D(n11893), .CK(clk), .RN(n5865), .Q(
        \I_cache/cache[6][111] ), .QN(n3013) );
  DFFRX1 \I_cache/cache_reg[7][111]  ( .D(n11892), .CK(clk), .RN(n5865), .Q(
        \I_cache/cache[7][111] ), .QN(n1445) );
  DFFRX1 \D_cache/cache_reg[4][142]  ( .D(\D_cache/n656 ), .CK(clk), .RN(n5928), .Q(\D_cache/cache[4][142] ), .QN(n2189) );
  DFFRX1 \D_cache/cache_reg[5][142]  ( .D(\D_cache/n655 ), .CK(clk), .RN(n5928), .Q(\D_cache/cache[5][142] ), .QN(n615) );
  DFFRX1 \D_cache/cache_reg[4][129]  ( .D(\D_cache/n760 ), .CK(clk), .RN(n5877), .Q(\D_cache/cache[4][129] ), .QN(n2188) );
  DFFRX1 \D_cache/cache_reg[5][129]  ( .D(\D_cache/n759 ), .CK(clk), .RN(n5876), .Q(\D_cache/cache[5][129] ), .QN(n614) );
  DFFRX1 \D_cache/cache_reg[5][131]  ( .D(\D_cache/n743 ), .CK(clk), .RN(n5935), .Q(\D_cache/cache[5][131] ), .QN(n566) );
  DFFRX1 \I_cache/cache_reg[0][153]  ( .D(n11563), .CK(clk), .RN(n5837), .Q(
        \I_cache/cache[0][153] ), .QN(n1729) );
  DFFRX1 \I_cache/cache_reg[1][153]  ( .D(n11562), .CK(clk), .RN(n5837), .Q(
        \I_cache/cache[1][153] ), .QN(n3336) );
  DFFRX1 \I_cache/cache_reg[2][153]  ( .D(n11561), .CK(clk), .RN(n5837), .Q(
        \I_cache/cache[2][153] ), .QN(n1728) );
  DFFRX1 \I_cache/cache_reg[3][153]  ( .D(n11560), .CK(clk), .RN(n5837), .Q(
        \I_cache/cache[3][153] ), .QN(n3335) );
  DFFRX1 \I_cache/cache_reg[4][153]  ( .D(n11559), .CK(clk), .RN(n5837), .Q(
        \I_cache/cache[4][153] ), .QN(n3325) );
  DFFRX1 \I_cache/cache_reg[5][153]  ( .D(n11558), .CK(clk), .RN(n5837), .Q(
        \I_cache/cache[5][153] ), .QN(n1723) );
  DFFRX1 \D_cache/cache_reg[0][142]  ( .D(\D_cache/n660 ), .CK(clk), .RN(n5928), .Q(\D_cache/cache[0][142] ), .QN(n2103) );
  DFFRX1 \D_cache/cache_reg[1][142]  ( .D(\D_cache/n659 ), .CK(clk), .RN(n5928), .Q(\D_cache/cache[1][142] ), .QN(n518) );
  DFFRX1 \D_cache/cache_reg[2][142]  ( .D(\D_cache/n658 ), .CK(clk), .RN(n5928), .Q(\D_cache/cache[2][142] ), .QN(n2109) );
  DFFRX1 \D_cache/cache_reg[3][142]  ( .D(\D_cache/n657 ), .CK(clk), .RN(n5928), .Q(\D_cache/cache[3][142] ), .QN(n522) );
  DFFRX1 \D_cache/cache_reg[6][142]  ( .D(\D_cache/n654 ), .CK(clk), .RN(n5928), .Q(\D_cache/cache[6][142] ), .QN(n2206) );
  DFFRX1 \D_cache/cache_reg[7][142]  ( .D(\D_cache/n653 ), .CK(clk), .RN(n5928), .Q(\D_cache/cache[7][142] ), .QN(n2207) );
  DFFRX1 \D_cache/cache_reg[0][129]  ( .D(\D_cache/n764 ), .CK(clk), .RN(n5877), .Q(\D_cache/cache[0][129] ), .QN(n2150) );
  DFFRX1 \D_cache/cache_reg[1][129]  ( .D(\D_cache/n763 ), .CK(clk), .RN(n5877), .Q(\D_cache/cache[1][129] ), .QN(n571) );
  DFFRX1 \D_cache/cache_reg[2][129]  ( .D(\D_cache/n762 ), .CK(clk), .RN(n5877), .Q(\D_cache/cache[2][129] ), .QN(n2121) );
  DFFRX1 \D_cache/cache_reg[3][129]  ( .D(\D_cache/n761 ), .CK(clk), .RN(n5877), .Q(\D_cache/cache[3][129] ), .QN(n534) );
  DFFRX1 \D_cache/cache_reg[6][129]  ( .D(\D_cache/n758 ), .CK(clk), .RN(n5876), .Q(\D_cache/cache[6][129] ), .QN(n2122) );
  DFFRX1 \D_cache/cache_reg[7][129]  ( .D(\D_cache/n757 ), .CK(clk), .RN(n5876), .Q(\D_cache/cache[7][129] ), .QN(n535) );
  DFFRX1 \D_cache/cache_reg[4][145]  ( .D(\D_cache/n632 ), .CK(clk), .RN(n5926), .Q(\D_cache/cache[4][145] ), .QN(n3367) );
  DFFRX1 \D_cache/cache_reg[5][145]  ( .D(\D_cache/n631 ), .CK(clk), .RN(n5931), .Q(\D_cache/cache[5][145] ), .QN(n1738) );
  DFFRX1 \D_cache/cache_reg[7][130]  ( .D(\D_cache/n749 ), .CK(clk), .RN(n5936), .Q(\D_cache/cache[7][130] ), .QN(n537) );
  DFFRX1 \D_cache/cache_reg[7][131]  ( .D(\D_cache/n741 ), .CK(clk), .RN(n5935), .Q(\D_cache/cache[7][131] ), .QN(n538) );
  DFFRX1 \D_cache/cache_reg[4][138]  ( .D(\D_cache/n688 ), .CK(clk), .RN(n5931), .Q(\D_cache/cache[4][138] ), .QN(n3393) );
  DFFRX1 \D_cache/cache_reg[5][138]  ( .D(\D_cache/n687 ), .CK(clk), .RN(n5931), .Q(\D_cache/cache[5][138] ), .QN(n1764) );
  DFFRX1 \D_cache/cache_reg[4][134]  ( .D(\D_cache/n720 ), .CK(clk), .RN(n5933), .Q(\D_cache/cache[4][134] ), .QN(n3390) );
  DFFRX1 \D_cache/cache_reg[5][134]  ( .D(\D_cache/n719 ), .CK(clk), .RN(n5933), .Q(\D_cache/cache[5][134] ), .QN(n1761) );
  DFFRX1 \D_cache/cache_reg[4][146]  ( .D(\D_cache/n624 ), .CK(clk), .RN(n5945), .Q(\D_cache/cache[4][146] ), .QN(n3392) );
  DFFRX1 \D_cache/cache_reg[5][146]  ( .D(\D_cache/n623 ), .CK(clk), .RN(n5945), .Q(\D_cache/cache[5][146] ), .QN(n1763) );
  DFFRX1 \D_cache/cache_reg[4][133]  ( .D(\D_cache/n728 ), .CK(clk), .RN(n5934), .Q(\D_cache/cache[4][133] ), .QN(n3387) );
  DFFRX1 \D_cache/cache_reg[5][133]  ( .D(\D_cache/n727 ), .CK(clk), .RN(n5934), .Q(\D_cache/cache[5][133] ), .QN(n1758) );
  DFFRX1 \D_cache/cache_reg[5][143]  ( .D(\D_cache/n647 ), .CK(clk), .RN(n5927), .Q(\D_cache/cache[5][143] ), .QN(n3402) );
  DFFRX1 \D_cache/cache_reg[5][150]  ( .D(\D_cache/n591 ), .CK(clk), .RN(n5943), .Q(\D_cache/cache[5][150] ), .QN(n3043) );
  DFFRX1 \D_cache/cache_reg[4][148]  ( .D(\D_cache/n608 ), .CK(clk), .RN(n5944), .Q(\D_cache/cache[4][148] ), .QN(n3376) );
  DFFRX1 \D_cache/cache_reg[5][148]  ( .D(\D_cache/n607 ), .CK(clk), .RN(n5944), .Q(\D_cache/cache[5][148] ), .QN(n1747) );
  DFFRX1 \D_cache/cache_reg[4][135]  ( .D(\D_cache/n712 ), .CK(clk), .RN(n5933), .Q(\D_cache/cache[4][135] ), .QN(n3382) );
  DFFRX1 \D_cache/cache_reg[5][135]  ( .D(\D_cache/n711 ), .CK(clk), .RN(n5933), .Q(\D_cache/cache[5][135] ), .QN(n1753) );
  DFFRX1 \D_cache/cache_reg[4][132]  ( .D(\D_cache/n736 ), .CK(clk), .RN(n5935), .Q(\D_cache/cache[4][132] ), .QN(n3379) );
  DFFRX1 \D_cache/cache_reg[5][132]  ( .D(\D_cache/n735 ), .CK(clk), .RN(n5935), .Q(\D_cache/cache[5][132] ), .QN(n1750) );
  DFFRX1 \D_cache/cache_reg[4][137]  ( .D(\D_cache/n696 ), .CK(clk), .RN(n5931), .Q(\D_cache/cache[4][137] ), .QN(n3385) );
  DFFRX1 \D_cache/cache_reg[5][137]  ( .D(\D_cache/n695 ), .CK(clk), .RN(n5931), .Q(\D_cache/cache[5][137] ), .QN(n1756) );
  DFFRX1 \D_cache/cache_reg[6][152]  ( .D(\D_cache/n574 ), .CK(clk), .RN(n5941), .Q(\D_cache/cache[6][152] ), .QN(n3373) );
  DFFRX1 \D_cache/cache_reg[7][152]  ( .D(\D_cache/n573 ), .CK(clk), .RN(n5941), .Q(\D_cache/cache[7][152] ), .QN(n1744) );
  DFFRX1 \D_cache/cache_reg[3][145]  ( .D(\D_cache/n633 ), .CK(clk), .RN(n5926), .Q(\D_cache/cache[3][145] ), .QN(n589) );
  DFFRX1 \D_cache/cache_reg[6][145]  ( .D(\D_cache/n630 ), .CK(clk), .RN(n5945), .Q(\D_cache/cache[6][145] ), .QN(n2102) );
  DFFRX1 \D_cache/cache_reg[7][145]  ( .D(\D_cache/n629 ), .CK(clk), .RN(n5955), .Q(\D_cache/cache[7][145] ), .QN(n517) );
  DFFRX1 \D_cache/cache_reg[2][152]  ( .D(\D_cache/n578 ), .CK(clk), .RN(n5941), .Q(\D_cache/cache[2][152] ), .QN(n3372) );
  DFFRX1 \D_cache/cache_reg[3][152]  ( .D(\D_cache/n577 ), .CK(clk), .RN(n5941), .Q(\D_cache/cache[3][152] ), .QN(n1743) );
  DFFRX1 \D_cache/cache_reg[6][139]  ( .D(\D_cache/n678 ), .CK(clk), .RN(n5930), .Q(\D_cache/cache[6][139] ) );
  DFFRX1 \D_cache/cache_reg[7][139]  ( .D(\D_cache/n677 ), .CK(clk), .RN(n5930), .Q(\D_cache/cache[7][139] ), .QN(n3345) );
  DFFRX1 \D_cache/cache_reg[2][139]  ( .D(\D_cache/n682 ), .CK(clk), .RN(n5930), .Q(\D_cache/cache[2][139] ), .QN(n3354) );
  DFFRX1 \D_cache/cache_reg[3][139]  ( .D(\D_cache/n681 ), .CK(clk), .RN(n5930), .Q(\D_cache/cache[3][139] ), .QN(n1734) );
  DFFRX1 \D_cache/cache_reg[6][144]  ( .D(\D_cache/n638 ), .CK(clk), .RN(n5926), .Q(\D_cache/cache[6][144] ), .QN(n3374) );
  DFFRX1 \D_cache/cache_reg[7][144]  ( .D(\D_cache/n637 ), .CK(clk), .RN(n5926), .Q(\D_cache/cache[7][144] ), .QN(n1745) );
  DFFRX1 \D_cache/cache_reg[2][144]  ( .D(\D_cache/n642 ), .CK(clk), .RN(n5927), .Q(\D_cache/cache[2][144] ), .QN(n3369) );
  DFFRX1 \D_cache/cache_reg[3][144]  ( .D(\D_cache/n641 ), .CK(clk), .RN(n5927), .Q(\D_cache/cache[3][144] ), .QN(n1740) );
  DFFRX1 \D_cache/cache_reg[2][140]  ( .D(\D_cache/n674 ), .CK(clk), .RN(n5929), .Q(\D_cache/cache[2][140] ), .QN(n2160) );
  DFFRX1 \D_cache/cache_reg[3][140]  ( .D(\D_cache/n673 ), .CK(clk), .RN(n5929), .Q(\D_cache/cache[3][140] ), .QN(n438) );
  DFFRX1 \D_cache/cache_reg[1][138]  ( .D(\D_cache/n691 ), .CK(clk), .RN(n5931), .Q(\D_cache/cache[1][138] ), .QN(n3364) );
  DFFRX1 \D_cache/cache_reg[2][138]  ( .D(\D_cache/n690 ), .CK(clk), .RN(n5931), .Q(\D_cache/cache[2][138] ), .QN(n2154) );
  DFFRX1 \D_cache/cache_reg[3][138]  ( .D(\D_cache/n689 ), .CK(clk), .RN(n5931), .Q(\D_cache/cache[3][138] ), .QN(n575) );
  DFFRX1 \D_cache/cache_reg[6][138]  ( .D(\D_cache/n686 ), .CK(clk), .RN(n5930), .Q(\D_cache/cache[6][138] ), .QN(n2139) );
  DFFRX1 \D_cache/cache_reg[7][138]  ( .D(\D_cache/n685 ), .CK(clk), .RN(n5930), .Q(\D_cache/cache[7][138] ), .QN(n559) );
  DFFRX1 \D_cache/cache_reg[1][134]  ( .D(\D_cache/n723 ), .CK(clk), .RN(n5934), .Q(\D_cache/cache[1][134] ), .QN(n3363) );
  DFFRX1 \D_cache/cache_reg[2][134]  ( .D(\D_cache/n722 ), .CK(clk), .RN(n5934), .Q(\D_cache/cache[2][134] ), .QN(n3389) );
  DFFRX1 \D_cache/cache_reg[3][134]  ( .D(\D_cache/n721 ), .CK(clk), .RN(n5933), .Q(\D_cache/cache[3][134] ), .QN(n1760) );
  DFFRX1 \D_cache/cache_reg[6][134]  ( .D(\D_cache/n718 ), .CK(clk), .RN(n5933), .Q(\D_cache/cache[6][134] ), .QN(n3391) );
  DFFRX1 \D_cache/cache_reg[7][134]  ( .D(\D_cache/n717 ), .CK(clk), .RN(n5933), .Q(\D_cache/cache[7][134] ), .QN(n1762) );
  DFFRX1 \D_cache/cache_reg[6][140]  ( .D(\D_cache/n670 ), .CK(clk), .RN(n5929), .Q(\D_cache/cache[6][140] ), .QN(n2111) );
  DFFRX1 \D_cache/cache_reg[7][140]  ( .D(\D_cache/n669 ), .CK(clk), .RN(n5929), .Q(\D_cache/cache[7][140] ), .QN(n524) );
  DFFRX1 \D_cache/cache_reg[1][146]  ( .D(\D_cache/n627 ), .CK(clk), .RN(n5971), .Q(\D_cache/cache[1][146] ), .QN(n578) );
  DFFRX1 \D_cache/cache_reg[3][146]  ( .D(\D_cache/n625 ), .CK(clk), .RN(n5945), .Q(\D_cache/cache[3][146] ), .QN(n2330) );
  DFFRX1 \D_cache/cache_reg[6][146]  ( .D(\D_cache/n622 ), .CK(clk), .RN(n5945), .Q(\D_cache/cache[6][146] ), .QN(n2104) );
  DFFRX1 \D_cache/cache_reg[7][146]  ( .D(\D_cache/n621 ), .CK(clk), .RN(n5945), .Q(\D_cache/cache[7][146] ), .QN(n519) );
  DFFRX1 \D_cache/cache_reg[1][133]  ( .D(\D_cache/n731 ), .CK(clk), .RN(n5934), .Q(\D_cache/cache[1][133] ), .QN(n3361) );
  DFFRX1 \D_cache/cache_reg[3][133]  ( .D(\D_cache/n729 ), .CK(clk), .RN(n5934), .Q(\D_cache/cache[3][133] ), .QN(n3362) );
  DFFRX1 \D_cache/cache_reg[6][133]  ( .D(\D_cache/n726 ), .CK(clk), .RN(n5934), .Q(\D_cache/cache[6][133] ), .QN(n3388) );
  DFFRX1 \D_cache/cache_reg[7][133]  ( .D(\D_cache/n725 ), .CK(clk), .RN(n5934), .Q(\D_cache/cache[7][133] ), .QN(n1759) );
  DFFRX1 \D_cache/cache_reg[7][141]  ( .D(\D_cache/n661 ), .CK(clk), .RN(n5928), .Q(\D_cache/cache[7][141] ), .QN(n3353) );
  DFFRX1 \D_cache/cache_reg[7][143]  ( .D(\D_cache/n645 ), .CK(clk), .RN(n5927), .Q(\D_cache/cache[7][143] ), .QN(n3365) );
  DFFRX1 \D_cache/cache_reg[7][150]  ( .D(\D_cache/n589 ), .CK(clk), .RN(n5942), .Q(\D_cache/cache[7][150] ), .QN(n3209) );
  DFFRX1 \D_cache/cache_reg[4][152]  ( .D(\D_cache/n576 ), .CK(clk), .RN(n5941), .Q(\D_cache/cache[4][152] ), .QN(n2221) );
  DFFRX1 \D_cache/cache_reg[5][152]  ( .D(\D_cache/n575 ), .CK(clk), .RN(n5941), .Q(\D_cache/cache[5][152] ), .QN(n2436) );
  DFFRX1 \D_cache/cache_reg[0][148]  ( .D(\D_cache/n612 ), .CK(clk), .RN(n5944), .Q(\D_cache/cache[0][148] ), .QN(n3366) );
  DFFRX1 \D_cache/cache_reg[1][148]  ( .D(\D_cache/n611 ), .CK(clk), .RN(n5944), .Q(\D_cache/cache[1][148] ), .QN(n1737) );
  DFFRX1 \D_cache/cache_reg[2][148]  ( .D(\D_cache/n610 ), .CK(clk), .RN(n5944), .Q(\D_cache/cache[2][148] ), .QN(n3375) );
  DFFRX1 \D_cache/cache_reg[3][148]  ( .D(\D_cache/n609 ), .CK(clk), .RN(n5944), .Q(\D_cache/cache[3][148] ), .QN(n1746) );
  DFFRX1 \D_cache/cache_reg[6][148]  ( .D(\D_cache/n606 ), .CK(clk), .RN(n5944), .Q(\D_cache/cache[6][148] ), .QN(n3377) );
  DFFRX1 \D_cache/cache_reg[7][148]  ( .D(\D_cache/n605 ), .CK(clk), .RN(n5944), .Q(\D_cache/cache[7][148] ), .QN(n1748) );
  DFFRX1 \D_cache/cache_reg[0][135]  ( .D(\D_cache/n716 ), .CK(clk), .RN(n5933), .Q(\D_cache/cache[0][135] ), .QN(n3371) );
  DFFRX1 \D_cache/cache_reg[1][135]  ( .D(\D_cache/n715 ), .CK(clk), .RN(n5933), .Q(\D_cache/cache[1][135] ), .QN(n1742) );
  DFFRX1 \D_cache/cache_reg[2][135]  ( .D(\D_cache/n714 ), .CK(clk), .RN(n5933), .Q(\D_cache/cache[2][135] ), .QN(n3381) );
  DFFRX1 \D_cache/cache_reg[3][135]  ( .D(\D_cache/n713 ), .CK(clk), .RN(n5933), .Q(\D_cache/cache[3][135] ), .QN(n1752) );
  DFFRX1 \D_cache/cache_reg[6][135]  ( .D(\D_cache/n710 ), .CK(clk), .RN(n5933), .Q(\D_cache/cache[6][135] ), .QN(n3383) );
  DFFRX1 \D_cache/cache_reg[7][135]  ( .D(\D_cache/n709 ), .CK(clk), .RN(n5932), .Q(\D_cache/cache[7][135] ), .QN(n1754) );
  DFFRX1 \D_cache/cache_reg[0][132]  ( .D(\D_cache/n740 ), .CK(clk), .RN(n5935), .Q(\D_cache/cache[0][132] ), .QN(n3370) );
  DFFRX1 \D_cache/cache_reg[1][132]  ( .D(\D_cache/n739 ), .CK(clk), .RN(n5935), .Q(\D_cache/cache[1][132] ), .QN(n1741) );
  DFFRX1 \D_cache/cache_reg[2][132]  ( .D(\D_cache/n738 ), .CK(clk), .RN(n5935), .Q(\D_cache/cache[2][132] ), .QN(n3378) );
  DFFRX1 \D_cache/cache_reg[3][132]  ( .D(\D_cache/n737 ), .CK(clk), .RN(n5935), .Q(\D_cache/cache[3][132] ), .QN(n1749) );
  DFFRX1 \D_cache/cache_reg[6][132]  ( .D(\D_cache/n734 ), .CK(clk), .RN(n5935), .Q(\D_cache/cache[6][132] ), .QN(n3380) );
  DFFRX1 \D_cache/cache_reg[7][132]  ( .D(\D_cache/n733 ), .CK(clk), .RN(n5934), .Q(\D_cache/cache[7][132] ), .QN(n1751) );
  DFFRX1 \D_cache/cache_reg[0][137]  ( .D(\D_cache/n700 ), .CK(clk), .RN(n5932), .Q(\D_cache/cache[0][137] ), .QN(n3368) );
  DFFRX1 \D_cache/cache_reg[1][137]  ( .D(\D_cache/n699 ), .CK(clk), .RN(n5932), .Q(\D_cache/cache[1][137] ), .QN(n1739) );
  DFFRX1 \D_cache/cache_reg[2][137]  ( .D(\D_cache/n698 ), .CK(clk), .RN(n5932), .Q(\D_cache/cache[2][137] ), .QN(n3384) );
  DFFRX1 \D_cache/cache_reg[3][137]  ( .D(\D_cache/n697 ), .CK(clk), .RN(n5931), .Q(\D_cache/cache[3][137] ), .QN(n1755) );
  DFFRX1 \D_cache/cache_reg[6][137]  ( .D(\D_cache/n694 ), .CK(clk), .RN(n5931), .Q(\D_cache/cache[6][137] ), .QN(n3386) );
  DFFRX1 \D_cache/cache_reg[7][137]  ( .D(\D_cache/n693 ), .CK(clk), .RN(n5931), .Q(\D_cache/cache[7][137] ), .QN(n1757) );
  DFFRX1 \i_MIPS/ID_EX_reg[98]  ( .D(\i_MIPS/n487 ), .CK(clk), .RN(n5742), .Q(
        \i_MIPS/ID_EX[98] ) );
  DFFRX1 \i_MIPS/ID_EX_reg[103]  ( .D(\i_MIPS/n482 ), .CK(clk), .RN(n5742), 
        .Q(\i_MIPS/ID_EX[103] ), .QN(n4492) );
  DFFRX1 \i_MIPS/ID_EX_reg[93]  ( .D(\i_MIPS/n492 ), .CK(clk), .RN(n5741), .Q(
        \i_MIPS/ID_EX[93] ), .QN(n4497) );
  DFFRX1 \i_MIPS/ID_EX_reg[90]  ( .D(\i_MIPS/n495 ), .CK(clk), .RN(n5741), .Q(
        \i_MIPS/ID_EX[90] ), .QN(n4495) );
  DFFRX1 \i_MIPS/ID_EX_reg[91]  ( .D(\i_MIPS/n494 ), .CK(clk), .RN(n5741), .Q(
        \i_MIPS/ID_EX[91] ), .QN(n4494) );
  DFFRX1 \i_MIPS/ID_EX_reg[92]  ( .D(\i_MIPS/n493 ), .CK(clk), .RN(n5741), .Q(
        \i_MIPS/ID_EX[92] ), .QN(n4496) );
  DFFRX1 \D_cache/cache_reg[0][154]  ( .D(\D_cache/n564 ), .CK(clk), .RN(n5940), .Q(\D_cache/cache[0][154] ) );
  DFFRX1 \D_cache/cache_reg[1][154]  ( .D(\D_cache/n563 ), .CK(clk), .RN(n5940), .Q(\D_cache/cache[1][154] ) );
  DFFRX1 \D_cache/cache_reg[2][154]  ( .D(\D_cache/n562 ), .CK(clk), .RN(n5940), .Q(\D_cache/cache[2][154] ) );
  DFFRX1 \D_cache/cache_reg[3][154]  ( .D(\D_cache/n561 ), .CK(clk), .RN(n5940), .Q(\D_cache/cache[3][154] ) );
  DFFRX1 \D_cache/cache_reg[4][154]  ( .D(\D_cache/n560 ), .CK(clk), .RN(n5940), .Q(\D_cache/cache[4][154] ) );
  DFFRX1 \D_cache/cache_reg[5][154]  ( .D(\D_cache/n559 ), .CK(clk), .RN(n5940), .Q(\D_cache/cache[5][154] ) );
  DFFRX1 \D_cache/cache_reg[6][154]  ( .D(\D_cache/n558 ), .CK(clk), .RN(n5940), .Q(\D_cache/cache[6][154] ) );
  DFFRX1 \D_cache/cache_reg[7][154]  ( .D(\D_cache/n557 ), .CK(clk), .RN(n5939), .Q(\D_cache/cache[7][154] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][0]  ( .D(\i_MIPS/Register/n148 ), 
        .CK(clk), .RN(n5706), .Q(\i_MIPS/Register/register[30][0] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][1]  ( .D(\i_MIPS/Register/n149 ), 
        .CK(clk), .RN(n5711), .Q(\i_MIPS/Register/register[30][1] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][2]  ( .D(\i_MIPS/Register/n150 ), 
        .CK(clk), .RN(n5726), .Q(\i_MIPS/Register/register[30][2] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][3]  ( .D(\i_MIPS/Register/n151 ), 
        .CK(clk), .RN(n5726), .Q(\i_MIPS/Register/register[30][3] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][4]  ( .D(\i_MIPS/Register/n152 ), 
        .CK(clk), .RN(n5726), .Q(\i_MIPS/Register/register[30][4] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][5]  ( .D(\i_MIPS/Register/n153 ), 
        .CK(clk), .RN(n5726), .Q(\i_MIPS/Register/register[30][5] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][6]  ( .D(\i_MIPS/Register/n154 ), 
        .CK(clk), .RN(n5726), .Q(\i_MIPS/Register/register[30][6] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][7]  ( .D(\i_MIPS/Register/n155 ), 
        .CK(clk), .RN(n5726), .Q(\i_MIPS/Register/register[30][7] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][8]  ( .D(\i_MIPS/Register/n156 ), 
        .CK(clk), .RN(n5726), .Q(\i_MIPS/Register/register[30][8] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][9]  ( .D(\i_MIPS/Register/n157 ), 
        .CK(clk), .RN(n5726), .Q(\i_MIPS/Register/register[30][9] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][10]  ( .D(\i_MIPS/Register/n158 ), 
        .CK(clk), .RN(n5726), .Q(\i_MIPS/Register/register[30][10] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][11]  ( .D(\i_MIPS/Register/n159 ), 
        .CK(clk), .RN(n5725), .Q(\i_MIPS/Register/register[30][11] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][12]  ( .D(\i_MIPS/Register/n160 ), 
        .CK(clk), .RN(n5725), .Q(\i_MIPS/Register/register[30][12] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][13]  ( .D(\i_MIPS/Register/n161 ), 
        .CK(clk), .RN(n5725), .Q(\i_MIPS/Register/register[30][13] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][14]  ( .D(\i_MIPS/Register/n162 ), 
        .CK(clk), .RN(n5725), .Q(\i_MIPS/Register/register[30][14] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][15]  ( .D(\i_MIPS/Register/n163 ), 
        .CK(clk), .RN(n5725), .Q(\i_MIPS/Register/register[30][15] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][16]  ( .D(\i_MIPS/Register/n164 ), 
        .CK(clk), .RN(n5725), .Q(\i_MIPS/Register/register[30][16] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][17]  ( .D(\i_MIPS/Register/n165 ), 
        .CK(clk), .RN(n5725), .Q(\i_MIPS/Register/register[30][17] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][18]  ( .D(\i_MIPS/Register/n166 ), 
        .CK(clk), .RN(n5725), .Q(\i_MIPS/Register/register[30][18] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][20]  ( .D(\i_MIPS/Register/n168 ), 
        .CK(clk), .RN(n5725), .Q(\i_MIPS/Register/register[30][20] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][21]  ( .D(\i_MIPS/Register/n169 ), 
        .CK(clk), .RN(n5725), .Q(\i_MIPS/Register/register[30][21] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][22]  ( .D(\i_MIPS/Register/n170 ), 
        .CK(clk), .RN(n5725), .Q(\i_MIPS/Register/register[30][22] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][23]  ( .D(\i_MIPS/Register/n171 ), 
        .CK(clk), .RN(n5724), .Q(\i_MIPS/Register/register[30][23] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][24]  ( .D(\i_MIPS/Register/n172 ), 
        .CK(clk), .RN(n5724), .Q(\i_MIPS/Register/register[30][24] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][25]  ( .D(\i_MIPS/Register/n173 ), 
        .CK(clk), .RN(n5724), .Q(\i_MIPS/Register/register[30][25] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][26]  ( .D(\i_MIPS/Register/n174 ), 
        .CK(clk), .RN(n5724), .Q(\i_MIPS/Register/register[30][26] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][27]  ( .D(\i_MIPS/Register/n175 ), 
        .CK(clk), .RN(n5724), .Q(\i_MIPS/Register/register[30][27] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][28]  ( .D(\i_MIPS/Register/n176 ), 
        .CK(clk), .RN(n5724), .Q(\i_MIPS/Register/register[30][28] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][29]  ( .D(\i_MIPS/Register/n177 ), 
        .CK(clk), .RN(n5724), .Q(\i_MIPS/Register/register[30][29] ) );
  DFFRX1 \i_MIPS/Register/register_reg[29][27]  ( .D(\i_MIPS/Register/n207 ), 
        .CK(clk), .RN(n5721), .Q(\i_MIPS/Register/register[29][27] ) );
  DFFRX1 \i_MIPS/Register/register_reg[27][27]  ( .D(\i_MIPS/Register/n271 ), 
        .CK(clk), .RN(n5776), .Q(\i_MIPS/Register/register[27][27] ) );
  DFFRX1 \i_MIPS/Register/register_reg[25][27]  ( .D(\i_MIPS/Register/n335 ), 
        .CK(clk), .RN(n5771), .Q(\i_MIPS/Register/register[25][27] ) );
  DFFRX1 \i_MIPS/Register/register_reg[15][27]  ( .D(\i_MIPS/Register/n655 ), 
        .CK(clk), .RN(n5764), .Q(\i_MIPS/Register/register[15][27] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][0]  ( .D(\i_MIPS/Register/n660 ), 
        .CK(clk), .RN(n5763), .Q(\i_MIPS/Register/register[14][0] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][1]  ( .D(\i_MIPS/Register/n661 ), 
        .CK(clk), .RN(n5763), .Q(\i_MIPS/Register/register[14][1] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][2]  ( .D(\i_MIPS/Register/n662 ), 
        .CK(clk), .RN(n5763), .Q(\i_MIPS/Register/register[14][2] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][3]  ( .D(\i_MIPS/Register/n663 ), 
        .CK(clk), .RN(n5763), .Q(\i_MIPS/Register/register[14][3] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][4]  ( .D(\i_MIPS/Register/n664 ), 
        .CK(clk), .RN(n5763), .Q(\i_MIPS/Register/register[14][4] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][5]  ( .D(\i_MIPS/Register/n665 ), 
        .CK(clk), .RN(n5763), .Q(\i_MIPS/Register/register[14][5] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][6]  ( .D(\i_MIPS/Register/n666 ), 
        .CK(clk), .RN(n5763), .Q(\i_MIPS/Register/register[14][6] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][7]  ( .D(\i_MIPS/Register/n667 ), 
        .CK(clk), .RN(n5763), .Q(\i_MIPS/Register/register[14][7] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][8]  ( .D(\i_MIPS/Register/n668 ), 
        .CK(clk), .RN(n5763), .Q(\i_MIPS/Register/register[14][8] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][9]  ( .D(\i_MIPS/Register/n669 ), 
        .CK(clk), .RN(n5763), .Q(\i_MIPS/Register/register[14][9] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][10]  ( .D(\i_MIPS/Register/n670 ), 
        .CK(clk), .RN(n5763), .Q(\i_MIPS/Register/register[14][10] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][11]  ( .D(\i_MIPS/Register/n671 ), 
        .CK(clk), .RN(n5763), .Q(\i_MIPS/Register/register[14][11] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][12]  ( .D(\i_MIPS/Register/n672 ), 
        .CK(clk), .RN(n5762), .Q(\i_MIPS/Register/register[14][12] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][13]  ( .D(\i_MIPS/Register/n673 ), 
        .CK(clk), .RN(n5762), .Q(\i_MIPS/Register/register[14][13] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][14]  ( .D(\i_MIPS/Register/n674 ), 
        .CK(clk), .RN(n5762), .Q(\i_MIPS/Register/register[14][14] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][15]  ( .D(\i_MIPS/Register/n675 ), 
        .CK(clk), .RN(n5762), .Q(\i_MIPS/Register/register[14][15] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][16]  ( .D(\i_MIPS/Register/n676 ), 
        .CK(clk), .RN(n5762), .Q(\i_MIPS/Register/register[14][16] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][17]  ( .D(\i_MIPS/Register/n677 ), 
        .CK(clk), .RN(n5762), .Q(\i_MIPS/Register/register[14][17] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][18]  ( .D(\i_MIPS/Register/n678 ), 
        .CK(clk), .RN(n5762), .Q(\i_MIPS/Register/register[14][18] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][20]  ( .D(\i_MIPS/Register/n680 ), 
        .CK(clk), .RN(n5762), .Q(\i_MIPS/Register/register[14][20] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][21]  ( .D(\i_MIPS/Register/n681 ), 
        .CK(clk), .RN(n5762), .Q(\i_MIPS/Register/register[14][21] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][22]  ( .D(\i_MIPS/Register/n682 ), 
        .CK(clk), .RN(n5762), .Q(\i_MIPS/Register/register[14][22] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][23]  ( .D(\i_MIPS/Register/n683 ), 
        .CK(clk), .RN(n5762), .Q(\i_MIPS/Register/register[14][23] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][24]  ( .D(\i_MIPS/Register/n684 ), 
        .CK(clk), .RN(n5761), .Q(\i_MIPS/Register/register[14][24] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][25]  ( .D(\i_MIPS/Register/n685 ), 
        .CK(clk), .RN(n5761), .Q(\i_MIPS/Register/register[14][25] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][26]  ( .D(\i_MIPS/Register/n686 ), 
        .CK(clk), .RN(n5761), .Q(\i_MIPS/Register/register[14][26] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][27]  ( .D(\i_MIPS/Register/n687 ), 
        .CK(clk), .RN(n5761), .Q(\i_MIPS/Register/register[14][27] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][28]  ( .D(\i_MIPS/Register/n688 ), 
        .CK(clk), .RN(n5761), .Q(\i_MIPS/Register/register[14][28] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][29]  ( .D(\i_MIPS/Register/n689 ), 
        .CK(clk), .RN(n5761), .Q(\i_MIPS/Register/register[14][29] ) );
  DFFRX1 \i_MIPS/Register/register_reg[13][27]  ( .D(\i_MIPS/Register/n719 ), 
        .CK(clk), .RN(n5758), .Q(\i_MIPS/Register/register[13][27] ) );
  DFFRX1 \i_MIPS/Register/register_reg[11][27]  ( .D(\i_MIPS/Register/n783 ), 
        .CK(clk), .RN(n5654), .Q(\i_MIPS/Register/register[11][27] ) );
  DFFRX1 \i_MIPS/Register/register_reg[9][27]  ( .D(\i_MIPS/Register/n847 ), 
        .CK(clk), .RN(n5648), .Q(\i_MIPS/Register/register[9][27] ) );
  DFFRX1 \i_MIPS/Register/register_reg[23][27]  ( .D(\i_MIPS/Register/n399 ), 
        .CK(clk), .RN(n5785), .Q(\i_MIPS/Register/register[23][27] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][0]  ( .D(\i_MIPS/Register/n404 ), 
        .CK(clk), .RN(n5785), .Q(\i_MIPS/Register/register[22][0] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][1]  ( .D(\i_MIPS/Register/n405 ), 
        .CK(clk), .RN(n5785), .Q(\i_MIPS/Register/register[22][1] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][2]  ( .D(\i_MIPS/Register/n406 ), 
        .CK(clk), .RN(n5785), .Q(\i_MIPS/Register/register[22][2] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][3]  ( .D(\i_MIPS/Register/n407 ), 
        .CK(clk), .RN(n5785), .Q(\i_MIPS/Register/register[22][3] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][4]  ( .D(\i_MIPS/Register/n408 ), 
        .CK(clk), .RN(n5785), .Q(\i_MIPS/Register/register[22][4] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][5]  ( .D(\i_MIPS/Register/n409 ), 
        .CK(clk), .RN(n5785), .Q(\i_MIPS/Register/register[22][5] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][6]  ( .D(\i_MIPS/Register/n410 ), 
        .CK(clk), .RN(n5784), .Q(\i_MIPS/Register/register[22][6] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][7]  ( .D(\i_MIPS/Register/n411 ), 
        .CK(clk), .RN(n5784), .Q(\i_MIPS/Register/register[22][7] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][8]  ( .D(\i_MIPS/Register/n412 ), 
        .CK(clk), .RN(n5784), .Q(\i_MIPS/Register/register[22][8] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][9]  ( .D(\i_MIPS/Register/n413 ), 
        .CK(clk), .RN(n5784), .Q(\i_MIPS/Register/register[22][9] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][10]  ( .D(\i_MIPS/Register/n414 ), 
        .CK(clk), .RN(n5784), .Q(\i_MIPS/Register/register[22][10] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][11]  ( .D(\i_MIPS/Register/n415 ), 
        .CK(clk), .RN(n5784), .Q(\i_MIPS/Register/register[22][11] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][12]  ( .D(\i_MIPS/Register/n416 ), 
        .CK(clk), .RN(n5784), .Q(\i_MIPS/Register/register[22][12] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][13]  ( .D(\i_MIPS/Register/n417 ), 
        .CK(clk), .RN(n5784), .Q(\i_MIPS/Register/register[22][13] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][14]  ( .D(\i_MIPS/Register/n418 ), 
        .CK(clk), .RN(n5784), .Q(\i_MIPS/Register/register[22][14] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][15]  ( .D(\i_MIPS/Register/n419 ), 
        .CK(clk), .RN(n5784), .Q(\i_MIPS/Register/register[22][15] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][16]  ( .D(\i_MIPS/Register/n420 ), 
        .CK(clk), .RN(n5784), .Q(\i_MIPS/Register/register[22][16] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][17]  ( .D(\i_MIPS/Register/n421 ), 
        .CK(clk), .RN(n5784), .Q(\i_MIPS/Register/register[22][17] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][18]  ( .D(\i_MIPS/Register/n422 ), 
        .CK(clk), .RN(n5783), .Q(\i_MIPS/Register/register[22][18] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][20]  ( .D(\i_MIPS/Register/n424 ), 
        .CK(clk), .RN(n5783), .Q(\i_MIPS/Register/register[22][20] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][21]  ( .D(\i_MIPS/Register/n425 ), 
        .CK(clk), .RN(n5783), .Q(\i_MIPS/Register/register[22][21] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][23]  ( .D(\i_MIPS/Register/n427 ), 
        .CK(clk), .RN(n5783), .Q(\i_MIPS/Register/register[22][23] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][24]  ( .D(\i_MIPS/Register/n428 ), 
        .CK(clk), .RN(n5783), .Q(\i_MIPS/Register/register[22][24] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][25]  ( .D(\i_MIPS/Register/n429 ), 
        .CK(clk), .RN(n5783), .Q(\i_MIPS/Register/register[22][25] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][26]  ( .D(\i_MIPS/Register/n430 ), 
        .CK(clk), .RN(n5783), .Q(\i_MIPS/Register/register[22][26] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][27]  ( .D(\i_MIPS/Register/n431 ), 
        .CK(clk), .RN(n5783), .Q(\i_MIPS/Register/register[22][27] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][28]  ( .D(\i_MIPS/Register/n432 ), 
        .CK(clk), .RN(n5783), .Q(\i_MIPS/Register/register[22][28] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][29]  ( .D(\i_MIPS/Register/n433 ), 
        .CK(clk), .RN(n5783), .Q(\i_MIPS/Register/register[22][29] ) );
  DFFRX1 \i_MIPS/Register/register_reg[21][27]  ( .D(\i_MIPS/Register/n463 ), 
        .CK(clk), .RN(n5780), .Q(\i_MIPS/Register/register[21][27] ) );
  DFFRX1 \i_MIPS/Register/register_reg[19][27]  ( .D(\i_MIPS/Register/n527 ), 
        .CK(clk), .RN(n5755), .Q(\i_MIPS/Register/register[19][27] ) );
  DFFRX1 \i_MIPS/Register/register_reg[17][27]  ( .D(\i_MIPS/Register/n591 ), 
        .CK(clk), .RN(n5749), .Q(\i_MIPS/Register/register[17][27] ) );
  DFFRX1 \i_MIPS/Register/register_reg[7][27]  ( .D(\i_MIPS/Register/n911 ), 
        .CK(clk), .RN(n5663), .Q(\i_MIPS/Register/register[7][27] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][0]  ( .D(\i_MIPS/Register/n916 ), 
        .CK(clk), .RN(n5662), .Q(\i_MIPS/Register/register[6][0] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][1]  ( .D(\i_MIPS/Register/n917 ), 
        .CK(clk), .RN(n5662), .Q(\i_MIPS/Register/register[6][1] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][2]  ( .D(\i_MIPS/Register/n918 ), 
        .CK(clk), .RN(n5662), .Q(\i_MIPS/Register/register[6][2] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][3]  ( .D(\i_MIPS/Register/n919 ), 
        .CK(clk), .RN(n5662), .Q(\i_MIPS/Register/register[6][3] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][4]  ( .D(\i_MIPS/Register/n920 ), 
        .CK(clk), .RN(n5662), .Q(\i_MIPS/Register/register[6][4] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][5]  ( .D(\i_MIPS/Register/n921 ), 
        .CK(clk), .RN(n5662), .Q(\i_MIPS/Register/register[6][5] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][6]  ( .D(\i_MIPS/Register/n922 ), 
        .CK(clk), .RN(n5662), .Q(\i_MIPS/Register/register[6][6] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][7]  ( .D(\i_MIPS/Register/n923 ), 
        .CK(clk), .RN(n5662), .Q(\i_MIPS/Register/register[6][7] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][8]  ( .D(\i_MIPS/Register/n924 ), 
        .CK(clk), .RN(n5662), .Q(\i_MIPS/Register/register[6][8] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][9]  ( .D(\i_MIPS/Register/n925 ), 
        .CK(clk), .RN(n5662), .Q(\i_MIPS/Register/register[6][9] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][10]  ( .D(\i_MIPS/Register/n926 ), 
        .CK(clk), .RN(n5662), .Q(\i_MIPS/Register/register[6][10] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][11]  ( .D(\i_MIPS/Register/n927 ), 
        .CK(clk), .RN(n5662), .Q(\i_MIPS/Register/register[6][11] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][13]  ( .D(\i_MIPS/Register/n929 ), 
        .CK(clk), .RN(n5661), .Q(\i_MIPS/Register/register[6][13] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][14]  ( .D(\i_MIPS/Register/n930 ), 
        .CK(clk), .RN(n5661), .Q(\i_MIPS/Register/register[6][14] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][15]  ( .D(\i_MIPS/Register/n931 ), 
        .CK(clk), .RN(n5661), .Q(\i_MIPS/Register/register[6][15] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][16]  ( .D(\i_MIPS/Register/n932 ), 
        .CK(clk), .RN(n5661), .Q(\i_MIPS/Register/register[6][16] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][18]  ( .D(\i_MIPS/Register/n934 ), 
        .CK(clk), .RN(n5661), .Q(\i_MIPS/Register/register[6][18] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][20]  ( .D(\i_MIPS/Register/n936 ), 
        .CK(clk), .RN(n5661), .Q(\i_MIPS/Register/register[6][20] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][21]  ( .D(\i_MIPS/Register/n937 ), 
        .CK(clk), .RN(n5661), .Q(\i_MIPS/Register/register[6][21] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][23]  ( .D(\i_MIPS/Register/n939 ), 
        .CK(clk), .RN(n5660), .Q(\i_MIPS/Register/register[6][23] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][24]  ( .D(\i_MIPS/Register/n940 ), 
        .CK(clk), .RN(n5660), .Q(\i_MIPS/Register/register[6][24] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][25]  ( .D(\i_MIPS/Register/n941 ), 
        .CK(clk), .RN(n5660), .Q(\i_MIPS/Register/register[6][25] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][26]  ( .D(\i_MIPS/Register/n942 ), 
        .CK(clk), .RN(n5660), .Q(\i_MIPS/Register/register[6][26] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][27]  ( .D(\i_MIPS/Register/n943 ), 
        .CK(clk), .RN(n5660), .Q(\i_MIPS/Register/register[6][27] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][28]  ( .D(\i_MIPS/Register/n944 ), 
        .CK(clk), .RN(n5660), .Q(\i_MIPS/Register/register[6][28] ) );
  DFFRX1 \i_MIPS/Register/register_reg[5][27]  ( .D(\i_MIPS/Register/n975 ), 
        .CK(clk), .RN(n5657), .Q(\i_MIPS/Register/register[5][27] ) );
  DFFRX1 \i_MIPS/Register/register_reg[3][27]  ( .D(\i_MIPS/Register/n1039 ), 
        .CK(clk), .RN(n5632), .Q(\i_MIPS/Register/register[3][27] ) );
  DFFRX1 \i_MIPS/Register/register_reg[1][27]  ( .D(\i_MIPS/Register/n1103 ), 
        .CK(clk), .RN(n5627), .Q(\i_MIPS/Register/register[1][27] ) );
  DFFRX1 \i_MIPS/Register/register_reg[29][0]  ( .D(\i_MIPS/Register/n180 ), 
        .CK(clk), .RN(n5724), .Q(\i_MIPS/Register/register[29][0] ), .QN(n290)
         );
  DFFRX1 \i_MIPS/Register/register_reg[29][1]  ( .D(\i_MIPS/Register/n181 ), 
        .CK(clk), .RN(n5724), .Q(\i_MIPS/Register/register[29][1] ), .QN(n996)
         );
  DFFRX1 \i_MIPS/Register/register_reg[29][2]  ( .D(\i_MIPS/Register/n182 ), 
        .CK(clk), .RN(n5724), .Q(\i_MIPS/Register/register[29][2] ), .QN(n948)
         );
  DFFRX1 \i_MIPS/Register/register_reg[29][3]  ( .D(\i_MIPS/Register/n183 ), 
        .CK(clk), .RN(n5723), .Q(\i_MIPS/Register/register[29][3] ), .QN(n473)
         );
  DFFRX1 \i_MIPS/Register/register_reg[29][4]  ( .D(\i_MIPS/Register/n184 ), 
        .CK(clk), .RN(n5723), .Q(\i_MIPS/Register/register[29][4] ), .QN(n868)
         );
  DFFRX1 \i_MIPS/Register/register_reg[29][5]  ( .D(\i_MIPS/Register/n185 ), 
        .CK(clk), .RN(n5723), .Q(\i_MIPS/Register/register[29][5] ), .QN(n893)
         );
  DFFRX1 \i_MIPS/Register/register_reg[29][6]  ( .D(\i_MIPS/Register/n186 ), 
        .CK(clk), .RN(n5723), .Q(\i_MIPS/Register/register[29][6] ), .QN(n951)
         );
  DFFRX1 \i_MIPS/Register/register_reg[29][7]  ( .D(\i_MIPS/Register/n187 ), 
        .CK(clk), .RN(n5723), .Q(\i_MIPS/Register/register[29][7] ), .QN(n474)
         );
  DFFRX1 \i_MIPS/Register/register_reg[29][8]  ( .D(\i_MIPS/Register/n188 ), 
        .CK(clk), .RN(n5723), .Q(\i_MIPS/Register/register[29][8] ), .QN(n892)
         );
  DFFRX1 \i_MIPS/Register/register_reg[29][9]  ( .D(\i_MIPS/Register/n189 ), 
        .CK(clk), .RN(n5723), .Q(\i_MIPS/Register/register[29][9] ), .QN(n454)
         );
  DFFRX1 \i_MIPS/Register/register_reg[29][10]  ( .D(\i_MIPS/Register/n190 ), 
        .CK(clk), .RN(n5723), .Q(\i_MIPS/Register/register[29][10] ), .QN(n298) );
  DFFRX1 \i_MIPS/Register/register_reg[29][11]  ( .D(\i_MIPS/Register/n191 ), 
        .CK(clk), .RN(n5723), .Q(\i_MIPS/Register/register[29][11] ), .QN(n296) );
  DFFRX1 \i_MIPS/Register/register_reg[29][12]  ( .D(\i_MIPS/Register/n192 ), 
        .CK(clk), .RN(n5723), .Q(\i_MIPS/Register/register[29][12] ), .QN(n291) );
  DFFRX1 \i_MIPS/Register/register_reg[29][13]  ( .D(\i_MIPS/Register/n193 ), 
        .CK(clk), .RN(n5723), .Q(\i_MIPS/Register/register[29][13] ), .QN(n439) );
  DFFRX1 \i_MIPS/Register/register_reg[29][14]  ( .D(\i_MIPS/Register/n194 ), 
        .CK(clk), .RN(n5723), .Q(\i_MIPS/Register/register[29][14] ), .QN(n287) );
  DFFRX1 \i_MIPS/Register/register_reg[29][15]  ( .D(\i_MIPS/Register/n195 ), 
        .CK(clk), .RN(n5722), .Q(\i_MIPS/Register/register[29][15] ), .QN(n294) );
  DFFRX1 \i_MIPS/Register/register_reg[29][16]  ( .D(\i_MIPS/Register/n196 ), 
        .CK(clk), .RN(n5722), .Q(\i_MIPS/Register/register[29][16] ), .QN(n458) );
  DFFRX1 \i_MIPS/Register/register_reg[29][17]  ( .D(\i_MIPS/Register/n197 ), 
        .CK(clk), .RN(n5722), .Q(\i_MIPS/Register/register[29][17] ), .QN(n642) );
  DFFRX1 \i_MIPS/Register/register_reg[29][18]  ( .D(\i_MIPS/Register/n198 ), 
        .CK(clk), .RN(n5722), .Q(\i_MIPS/Register/register[29][18] ), .QN(n450) );
  DFFRX1 \i_MIPS/Register/register_reg[29][20]  ( .D(\i_MIPS/Register/n200 ), 
        .CK(clk), .RN(n5722), .Q(\i_MIPS/Register/register[29][20] ), .QN(n468) );
  DFFRX1 \i_MIPS/Register/register_reg[29][21]  ( .D(\i_MIPS/Register/n201 ), 
        .CK(clk), .RN(n5722), .Q(\i_MIPS/Register/register[29][21] ), .QN(n986) );
  DFFRX1 \i_MIPS/Register/register_reg[29][22]  ( .D(\i_MIPS/Register/n202 ), 
        .CK(clk), .RN(n5722), .Q(\i_MIPS/Register/register[29][22] ), .QN(n472) );
  DFFRX1 \i_MIPS/Register/register_reg[29][23]  ( .D(\i_MIPS/Register/n203 ), 
        .CK(clk), .RN(n5722), .Q(\i_MIPS/Register/register[29][23] ), .QN(n881) );
  DFFRX1 \i_MIPS/Register/register_reg[29][24]  ( .D(\i_MIPS/Register/n204 ), 
        .CK(clk), .RN(n5722), .Q(\i_MIPS/Register/register[29][24] ), .QN(n639) );
  DFFRX1 \i_MIPS/Register/register_reg[29][25]  ( .D(\i_MIPS/Register/n205 ), 
        .CK(clk), .RN(n5722), .Q(\i_MIPS/Register/register[29][25] ), .QN(n447) );
  DFFRX1 \i_MIPS/Register/register_reg[29][26]  ( .D(\i_MIPS/Register/n206 ), 
        .CK(clk), .RN(n5722), .Q(\i_MIPS/Register/register[29][26] ), .QN(n470) );
  DFFRX1 \i_MIPS/Register/register_reg[29][28]  ( .D(\i_MIPS/Register/n208 ), 
        .CK(clk), .RN(n5721), .Q(\i_MIPS/Register/register[29][28] ), .QN(n643) );
  DFFRX1 \i_MIPS/Register/register_reg[29][29]  ( .D(\i_MIPS/Register/n209 ), 
        .CK(clk), .RN(n5721), .Q(\i_MIPS/Register/register[29][29] ), .QN(n475) );
  DFFRX1 \i_MIPS/Register/register_reg[28][0]  ( .D(\i_MIPS/Register/n212 ), 
        .CK(clk), .RN(n5721), .Q(\i_MIPS/Register/register[28][0] ), .QN(n396)
         );
  DFFRX1 \i_MIPS/Register/register_reg[28][1]  ( .D(\i_MIPS/Register/n213 ), 
        .CK(clk), .RN(n5721), .Q(\i_MIPS/Register/register[28][1] ), .QN(n1009) );
  DFFRX1 \i_MIPS/Register/register_reg[28][2]  ( .D(\i_MIPS/Register/n214 ), 
        .CK(clk), .RN(n5721), .Q(\i_MIPS/Register/register[28][2] ), .QN(n939)
         );
  DFFRX1 \i_MIPS/Register/register_reg[28][3]  ( .D(\i_MIPS/Register/n215 ), 
        .CK(clk), .RN(n5721), .Q(\i_MIPS/Register/register[28][3] ), .QN(n1012) );
  DFFRX1 \i_MIPS/Register/register_reg[28][4]  ( .D(\i_MIPS/Register/n216 ), 
        .CK(clk), .RN(n5721), .Q(\i_MIPS/Register/register[28][4] ), .QN(n1015) );
  DFFRX1 \i_MIPS/Register/register_reg[28][6]  ( .D(\i_MIPS/Register/n218 ), 
        .CK(clk), .RN(n5720), .Q(\i_MIPS/Register/register[28][6] ), .QN(n940)
         );
  DFFRX1 \i_MIPS/Register/register_reg[28][7]  ( .D(\i_MIPS/Register/n219 ), 
        .CK(clk), .RN(n5720), .Q(\i_MIPS/Register/register[28][7] ), .QN(n889)
         );
  DFFRX1 \i_MIPS/Register/register_reg[28][9]  ( .D(\i_MIPS/Register/n221 ), 
        .CK(clk), .RN(n5720), .Q(\i_MIPS/Register/register[28][9] ), .QN(n1013) );
  DFFRX1 \i_MIPS/Register/register_reg[28][10]  ( .D(\i_MIPS/Register/n222 ), 
        .CK(clk), .RN(n5720), .Q(\i_MIPS/Register/register[28][10] ), .QN(n394) );
  DFFRX1 \i_MIPS/Register/register_reg[28][13]  ( .D(\i_MIPS/Register/n225 ), 
        .CK(clk), .RN(n5720), .Q(\i_MIPS/Register/register[28][13] ), .QN(n890) );
  DFFRX1 \i_MIPS/Register/register_reg[28][14]  ( .D(\i_MIPS/Register/n226 ), 
        .CK(clk), .RN(n5720), .Q(\i_MIPS/Register/register[28][14] ), .QN(n395) );
  DFFRX1 \i_MIPS/Register/register_reg[28][15]  ( .D(\i_MIPS/Register/n227 ), 
        .CK(clk), .RN(n5720), .Q(\i_MIPS/Register/register[28][15] ), .QN(n397) );
  DFFRX1 \i_MIPS/Register/register_reg[28][16]  ( .D(\i_MIPS/Register/n228 ), 
        .CK(clk), .RN(n5720), .Q(\i_MIPS/Register/register[28][16] ), .QN(n891) );
  DFFRX1 \i_MIPS/Register/register_reg[28][18]  ( .D(\i_MIPS/Register/n230 ), 
        .CK(clk), .RN(n5719), .Q(\i_MIPS/Register/register[28][18] ), .QN(
        n1008) );
  DFFRX1 \i_MIPS/Register/register_reg[28][20]  ( .D(\i_MIPS/Register/n232 ), 
        .CK(clk), .RN(n5719), .Q(\i_MIPS/Register/register[28][20] ), .QN(n958) );
  DFFRX1 \i_MIPS/Register/register_reg[28][21]  ( .D(\i_MIPS/Register/n233 ), 
        .CK(clk), .RN(n5719), .Q(\i_MIPS/Register/register[28][21] ), .QN(
        n1010) );
  DFFRX1 \i_MIPS/Register/register_reg[28][23]  ( .D(\i_MIPS/Register/n235 ), 
        .CK(clk), .RN(n5719), .Q(\i_MIPS/Register/register[28][23] ), .QN(
        n1011) );
  DFFRX1 \i_MIPS/Register/register_reg[28][25]  ( .D(\i_MIPS/Register/n237 ), 
        .CK(clk), .RN(n5719), .Q(\i_MIPS/Register/register[28][25] ), .QN(
        n1014) );
  DFFRX1 \i_MIPS/Register/register_reg[28][26]  ( .D(\i_MIPS/Register/n238 ), 
        .CK(clk), .RN(n5719), .Q(\i_MIPS/Register/register[28][26] ), .QN(n960) );
  DFFRX1 \i_MIPS/Register/register_reg[28][28]  ( .D(\i_MIPS/Register/n240 ), 
        .CK(clk), .RN(n5719), .Q(\i_MIPS/Register/register[28][28] ), .QN(n959) );
  DFFRX1 \i_MIPS/Register/register_reg[27][0]  ( .D(\i_MIPS/Register/n244 ), 
        .CK(clk), .RN(n5718), .Q(\i_MIPS/Register/register[27][0] ), .QN(n390)
         );
  DFFRX1 \i_MIPS/Register/register_reg[27][1]  ( .D(\i_MIPS/Register/n245 ), 
        .CK(clk), .RN(n5718), .Q(\i_MIPS/Register/register[27][1] ), .QN(n995)
         );
  DFFRX1 \i_MIPS/Register/register_reg[27][2]  ( .D(\i_MIPS/Register/n246 ), 
        .CK(clk), .RN(n5718), .Q(\i_MIPS/Register/register[27][2] ), .QN(n1005) );
  DFFRX1 \i_MIPS/Register/register_reg[27][3]  ( .D(\i_MIPS/Register/n247 ), 
        .CK(clk), .RN(n5718), .Q(\i_MIPS/Register/register[27][3] ), .QN(n352)
         );
  DFFRX1 \i_MIPS/Register/register_reg[27][4]  ( .D(\i_MIPS/Register/n248 ), 
        .CK(clk), .RN(n5718), .Q(\i_MIPS/Register/register[27][4] ), .QN(n917)
         );
  DFFRX1 \i_MIPS/Register/register_reg[27][5]  ( .D(\i_MIPS/Register/n249 ), 
        .CK(clk), .RN(n5718), .Q(\i_MIPS/Register/register[27][5] ), .QN(n919)
         );
  DFFRX1 \i_MIPS/Register/register_reg[27][6]  ( .D(\i_MIPS/Register/n250 ), 
        .CK(clk), .RN(n5718), .Q(\i_MIPS/Register/register[27][6] ), .QN(n950)
         );
  DFFRX1 \i_MIPS/Register/register_reg[27][7]  ( .D(\i_MIPS/Register/n251 ), 
        .CK(clk), .RN(n5718), .Q(\i_MIPS/Register/register[27][7] ), .QN(n901)
         );
  DFFRX1 \i_MIPS/Register/register_reg[27][8]  ( .D(\i_MIPS/Register/n252 ), 
        .CK(clk), .RN(n5718), .Q(\i_MIPS/Register/register[27][8] ), .QN(n983)
         );
  DFFRX1 \i_MIPS/Register/register_reg[27][9]  ( .D(\i_MIPS/Register/n253 ), 
        .CK(clk), .RN(n5718), .Q(\i_MIPS/Register/register[27][9] ), .QN(n382)
         );
  DFFRX1 \i_MIPS/Register/register_reg[27][10]  ( .D(\i_MIPS/Register/n254 ), 
        .CK(clk), .RN(n5717), .Q(\i_MIPS/Register/register[27][10] ), .QN(n370) );
  DFFRX1 \i_MIPS/Register/register_reg[27][11]  ( .D(\i_MIPS/Register/n255 ), 
        .CK(clk), .RN(n5717), .Q(\i_MIPS/Register/register[27][11] ), .QN(n327) );
  DFFRX1 \i_MIPS/Register/register_reg[27][12]  ( .D(\i_MIPS/Register/n256 ), 
        .CK(clk), .RN(n5717), .Q(\i_MIPS/Register/register[27][12] ), .QN(n365) );
  DFFRX1 \i_MIPS/Register/register_reg[27][13]  ( .D(\i_MIPS/Register/n257 ), 
        .CK(clk), .RN(n5717), .Q(\i_MIPS/Register/register[27][13] ), .QN(
        n1002) );
  DFFRX1 \i_MIPS/Register/register_reg[27][14]  ( .D(\i_MIPS/Register/n258 ), 
        .CK(clk), .RN(n5717), .Q(\i_MIPS/Register/register[27][14] ), .QN(n393) );
  DFFRX1 \i_MIPS/Register/register_reg[27][15]  ( .D(\i_MIPS/Register/n259 ), 
        .CK(clk), .RN(n5717), .Q(\i_MIPS/Register/register[27][15] ), .QN(n388) );
  DFFRX1 \i_MIPS/Register/register_reg[27][16]  ( .D(\i_MIPS/Register/n260 ), 
        .CK(clk), .RN(n5717), .Q(\i_MIPS/Register/register[27][16] ), .QN(n998) );
  DFFRX1 \i_MIPS/Register/register_reg[27][17]  ( .D(\i_MIPS/Register/n261 ), 
        .CK(clk), .RN(n5717), .Q(\i_MIPS/Register/register[27][17] ), .QN(n906) );
  DFFRX1 \i_MIPS/Register/register_reg[27][18]  ( .D(\i_MIPS/Register/n262 ), 
        .CK(clk), .RN(n5717), .Q(\i_MIPS/Register/register[27][18] ), .QN(n337) );
  DFFRX1 \i_MIPS/Register/register_reg[27][20]  ( .D(\i_MIPS/Register/n264 ), 
        .CK(clk), .RN(n5717), .Q(\i_MIPS/Register/register[27][20] ), .QN(n994) );
  DFFRX1 \i_MIPS/Register/register_reg[27][21]  ( .D(\i_MIPS/Register/n265 ), 
        .CK(clk), .RN(n5717), .Q(\i_MIPS/Register/register[27][21] ), .QN(n455) );
  DFFRX1 \i_MIPS/Register/register_reg[27][22]  ( .D(\i_MIPS/Register/n266 ), 
        .CK(clk), .RN(n5716), .Q(\i_MIPS/Register/register[27][22] ), .QN(n903) );
  DFFRX1 \i_MIPS/Register/register_reg[27][23]  ( .D(\i_MIPS/Register/n267 ), 
        .CK(clk), .RN(n5716), .Q(\i_MIPS/Register/register[27][23] ), .QN(n477) );
  DFFRX1 \i_MIPS/Register/register_reg[27][24]  ( .D(\i_MIPS/Register/n268 ), 
        .CK(clk), .RN(n5721), .Q(\i_MIPS/Register/register[27][24] ), .QN(n322) );
  DFFRX1 \i_MIPS/Register/register_reg[27][25]  ( .D(\i_MIPS/Register/n269 ), 
        .CK(clk), .RN(n5726), .Q(\i_MIPS/Register/register[27][25] ), .QN(n988) );
  DFFRX1 \i_MIPS/Register/register_reg[27][26]  ( .D(\i_MIPS/Register/n270 ), 
        .CK(clk), .RN(n5776), .Q(\i_MIPS/Register/register[27][26] ), .QN(n912) );
  DFFRX1 \i_MIPS/Register/register_reg[27][28]  ( .D(\i_MIPS/Register/n272 ), 
        .CK(clk), .RN(n5776), .Q(\i_MIPS/Register/register[27][28] ), .QN(n353) );
  DFFRX1 \i_MIPS/Register/register_reg[27][29]  ( .D(\i_MIPS/Register/n273 ), 
        .CK(clk), .RN(n5776), .Q(\i_MIPS/Register/register[27][29] ), .QN(n909) );
  DFFRX1 \i_MIPS/Register/register_reg[25][0]  ( .D(\i_MIPS/Register/n308 ), 
        .CK(clk), .RN(n5773), .Q(\i_MIPS/Register/register[25][0] ), .QN(n385)
         );
  DFFRX1 \i_MIPS/Register/register_reg[25][1]  ( .D(\i_MIPS/Register/n309 ), 
        .CK(clk), .RN(n5773), .Q(\i_MIPS/Register/register[25][1] ), .QN(n985)
         );
  DFFRX1 \i_MIPS/Register/register_reg[25][2]  ( .D(\i_MIPS/Register/n310 ), 
        .CK(clk), .RN(n5773), .Q(\i_MIPS/Register/register[25][2] ), .QN(n963)
         );
  DFFRX1 \i_MIPS/Register/register_reg[25][3]  ( .D(\i_MIPS/Register/n311 ), 
        .CK(clk), .RN(n5773), .Q(\i_MIPS/Register/register[25][3] ), .QN(n384)
         );
  DFFRX1 \i_MIPS/Register/register_reg[25][4]  ( .D(\i_MIPS/Register/n312 ), 
        .CK(clk), .RN(n5773), .Q(\i_MIPS/Register/register[25][4] ), .QN(n878)
         );
  DFFRX1 \i_MIPS/Register/register_reg[25][5]  ( .D(\i_MIPS/Register/n313 ), 
        .CK(clk), .RN(n5773), .Q(\i_MIPS/Register/register[25][5] ), .QN(n926)
         );
  DFFRX1 \i_MIPS/Register/register_reg[25][6]  ( .D(\i_MIPS/Register/n314 ), 
        .CK(clk), .RN(n5773), .Q(\i_MIPS/Register/register[25][6] ), .QN(n964)
         );
  DFFRX1 \i_MIPS/Register/register_reg[25][7]  ( .D(\i_MIPS/Register/n315 ), 
        .CK(clk), .RN(n5772), .Q(\i_MIPS/Register/register[25][7] ), .QN(n934)
         );
  DFFRX1 \i_MIPS/Register/register_reg[25][8]  ( .D(\i_MIPS/Register/n316 ), 
        .CK(clk), .RN(n5772), .Q(\i_MIPS/Register/register[25][8] ), .QN(n924)
         );
  DFFRX1 \i_MIPS/Register/register_reg[25][9]  ( .D(\i_MIPS/Register/n317 ), 
        .CK(clk), .RN(n5772), .Q(\i_MIPS/Register/register[25][9] ), .QN(n342)
         );
  DFFRX1 \i_MIPS/Register/register_reg[25][10]  ( .D(\i_MIPS/Register/n318 ), 
        .CK(clk), .RN(n5772), .Q(\i_MIPS/Register/register[25][10] ), .QN(n330) );
  DFFRX1 \i_MIPS/Register/register_reg[25][11]  ( .D(\i_MIPS/Register/n319 ), 
        .CK(clk), .RN(n5772), .Q(\i_MIPS/Register/register[25][11] ), .QN(n349) );
  DFFRX1 \i_MIPS/Register/register_reg[25][12]  ( .D(\i_MIPS/Register/n320 ), 
        .CK(clk), .RN(n5772), .Q(\i_MIPS/Register/register[25][12] ), .QN(n333) );
  DFFRX1 \i_MIPS/Register/register_reg[25][13]  ( .D(\i_MIPS/Register/n321 ), 
        .CK(clk), .RN(n5772), .Q(\i_MIPS/Register/register[25][13] ), .QN(n962) );
  DFFRX1 \i_MIPS/Register/register_reg[25][14]  ( .D(\i_MIPS/Register/n322 ), 
        .CK(clk), .RN(n5772), .Q(\i_MIPS/Register/register[25][14] ), .QN(n377) );
  DFFRX1 \i_MIPS/Register/register_reg[25][15]  ( .D(\i_MIPS/Register/n323 ), 
        .CK(clk), .RN(n5772), .Q(\i_MIPS/Register/register[25][15] ), .QN(n332) );
  DFFRX1 \i_MIPS/Register/register_reg[25][16]  ( .D(\i_MIPS/Register/n324 ), 
        .CK(clk), .RN(n5772), .Q(\i_MIPS/Register/register[25][16] ), .QN(n854) );
  DFFRX1 \i_MIPS/Register/register_reg[25][17]  ( .D(\i_MIPS/Register/n325 ), 
        .CK(clk), .RN(n5772), .Q(\i_MIPS/Register/register[25][17] ), .QN(n921) );
  DFFRX1 \i_MIPS/Register/register_reg[25][18]  ( .D(\i_MIPS/Register/n326 ), 
        .CK(clk), .RN(n5772), .Q(\i_MIPS/Register/register[25][18] ), .QN(n372) );
  DFFRX1 \i_MIPS/Register/register_reg[25][20]  ( .D(\i_MIPS/Register/n328 ), 
        .CK(clk), .RN(n5771), .Q(\i_MIPS/Register/register[25][20] ), .QN(n375) );
  DFFRX1 \i_MIPS/Register/register_reg[25][21]  ( .D(\i_MIPS/Register/n329 ), 
        .CK(clk), .RN(n5771), .Q(\i_MIPS/Register/register[25][21] ), .QN(n300) );
  DFFRX1 \i_MIPS/Register/register_reg[25][22]  ( .D(\i_MIPS/Register/n330 ), 
        .CK(clk), .RN(n5771), .Q(\i_MIPS/Register/register[25][22] ), .QN(n361) );
  DFFRX1 \i_MIPS/Register/register_reg[25][23]  ( .D(\i_MIPS/Register/n331 ), 
        .CK(clk), .RN(n5771), .Q(\i_MIPS/Register/register[25][23] ), .QN(n369) );
  DFFRX1 \i_MIPS/Register/register_reg[25][24]  ( .D(\i_MIPS/Register/n332 ), 
        .CK(clk), .RN(n5771), .Q(\i_MIPS/Register/register[25][24] ), .QN(n345) );
  DFFRX1 \i_MIPS/Register/register_reg[25][25]  ( .D(\i_MIPS/Register/n333 ), 
        .CK(clk), .RN(n5771), .Q(\i_MIPS/Register/register[25][25] ), .QN(n347) );
  DFFRX1 \i_MIPS/Register/register_reg[25][26]  ( .D(\i_MIPS/Register/n334 ), 
        .CK(clk), .RN(n5771), .Q(\i_MIPS/Register/register[25][26] ), .QN(n363) );
  DFFRX1 \i_MIPS/Register/register_reg[25][28]  ( .D(\i_MIPS/Register/n336 ), 
        .CK(clk), .RN(n5771), .Q(\i_MIPS/Register/register[25][28] ), .QN(n360) );
  DFFRX1 \i_MIPS/Register/register_reg[25][29]  ( .D(\i_MIPS/Register/n337 ), 
        .CK(clk), .RN(n5771), .Q(\i_MIPS/Register/register[25][29] ), .QN(n923) );
  DFFRX1 \i_MIPS/Register/register_reg[24][0]  ( .D(\i_MIPS/Register/n340 ), 
        .CK(clk), .RN(n5770), .Q(\i_MIPS/Register/register[24][0] ), .QN(n900)
         );
  DFFRX1 \i_MIPS/Register/register_reg[24][1]  ( .D(\i_MIPS/Register/n341 ), 
        .CK(clk), .RN(n5770), .Q(\i_MIPS/Register/register[24][1] ), .QN(n392)
         );
  DFFRX1 \i_MIPS/Register/register_reg[24][2]  ( .D(\i_MIPS/Register/n342 ), 
        .CK(clk), .RN(n5770), .Q(\i_MIPS/Register/register[24][2] ), .QN(n640)
         );
  DFFRX1 \i_MIPS/Register/register_reg[24][3]  ( .D(\i_MIPS/Register/n343 ), 
        .CK(clk), .RN(n5770), .Q(\i_MIPS/Register/register[24][3] ), .QN(n931)
         );
  DFFRX1 \i_MIPS/Register/register_reg[24][4]  ( .D(\i_MIPS/Register/n344 ), 
        .CK(clk), .RN(n5770), .Q(\i_MIPS/Register/register[24][4] ), .QN(n465)
         );
  DFFRX1 \i_MIPS/Register/register_reg[24][6]  ( .D(\i_MIPS/Register/n346 ), 
        .CK(clk), .RN(n5770), .Q(\i_MIPS/Register/register[24][6] ), .QN(n446)
         );
  DFFRX1 \i_MIPS/Register/register_reg[24][7]  ( .D(\i_MIPS/Register/n347 ), 
        .CK(clk), .RN(n5770), .Q(\i_MIPS/Register/register[24][7] ), .QN(n358)
         );
  DFFRX1 \i_MIPS/Register/register_reg[24][8]  ( .D(\i_MIPS/Register/n348 ), 
        .CK(clk), .RN(n5770), .Q(\i_MIPS/Register/register[24][8] ), .QN(n467)
         );
  DFFRX1 \i_MIPS/Register/register_reg[24][9]  ( .D(\i_MIPS/Register/n349 ), 
        .CK(clk), .RN(n5770), .Q(\i_MIPS/Register/register[24][9] ), .QN(n930)
         );
  DFFRX1 \i_MIPS/Register/register_reg[24][10]  ( .D(\i_MIPS/Register/n350 ), 
        .CK(clk), .RN(n5769), .Q(\i_MIPS/Register/register[24][10] ), .QN(n853) );
  DFFRX1 \i_MIPS/Register/register_reg[24][11]  ( .D(\i_MIPS/Register/n351 ), 
        .CK(clk), .RN(n5769), .Q(\i_MIPS/Register/register[24][11] ), .QN(n896) );
  DFFRX1 \i_MIPS/Register/register_reg[24][13]  ( .D(\i_MIPS/Register/n353 ), 
        .CK(clk), .RN(n5769), .Q(\i_MIPS/Register/register[24][13] ), .QN(n356) );
  DFFRX1 \i_MIPS/Register/register_reg[24][14]  ( .D(\i_MIPS/Register/n354 ), 
        .CK(clk), .RN(n5769), .Q(\i_MIPS/Register/register[24][14] ), .QN(n894) );
  DFFRX1 \i_MIPS/Register/register_reg[24][15]  ( .D(\i_MIPS/Register/n355 ), 
        .CK(clk), .RN(n5769), .Q(\i_MIPS/Register/register[24][15] ), .QN(n898) );
  DFFRX1 \i_MIPS/Register/register_reg[24][16]  ( .D(\i_MIPS/Register/n356 ), 
        .CK(clk), .RN(n5769), .Q(\i_MIPS/Register/register[24][16] ), .QN(n340) );
  DFFRX1 \i_MIPS/Register/register_reg[24][18]  ( .D(\i_MIPS/Register/n358 ), 
        .CK(clk), .RN(n5769), .Q(\i_MIPS/Register/register[24][18] ), .QN(n857) );
  DFFRX1 \i_MIPS/Register/register_reg[24][20]  ( .D(\i_MIPS/Register/n360 ), 
        .CK(clk), .RN(n5769), .Q(\i_MIPS/Register/register[24][20] ), .QN(n441) );
  DFFRX1 \i_MIPS/Register/register_reg[24][21]  ( .D(\i_MIPS/Register/n361 ), 
        .CK(clk), .RN(n5769), .Q(\i_MIPS/Register/register[24][21] ), .QN(n461) );
  DFFRX1 \i_MIPS/Register/register_reg[24][23]  ( .D(\i_MIPS/Register/n363 ), 
        .CK(clk), .RN(n5768), .Q(\i_MIPS/Register/register[24][23] ), .QN(n929) );
  DFFRX1 \i_MIPS/Register/register_reg[24][24]  ( .D(\i_MIPS/Register/n364 ), 
        .CK(clk), .RN(n5768), .Q(\i_MIPS/Register/register[24][24] ), .QN(n932) );
  DFFRX1 \i_MIPS/Register/register_reg[24][25]  ( .D(\i_MIPS/Register/n365 ), 
        .CK(clk), .RN(n5768), .Q(\i_MIPS/Register/register[24][25] ), .QN(n463) );
  DFFRX1 \i_MIPS/Register/register_reg[24][26]  ( .D(\i_MIPS/Register/n366 ), 
        .CK(clk), .RN(n5768), .Q(\i_MIPS/Register/register[24][26] ), .QN(n442) );
  DFFRX1 \i_MIPS/Register/register_reg[24][28]  ( .D(\i_MIPS/Register/n368 ), 
        .CK(clk), .RN(n5768), .Q(\i_MIPS/Register/register[24][28] ), .QN(n886) );
  DFFRX1 \i_MIPS/Register/register_reg[15][0]  ( .D(\i_MIPS/Register/n628 ), 
        .CK(clk), .RN(n5766), .Q(\i_MIPS/Register/register[15][0] ), .QN(n943)
         );
  DFFRX1 \i_MIPS/Register/register_reg[15][1]  ( .D(\i_MIPS/Register/n629 ), 
        .CK(clk), .RN(n5766), .Q(\i_MIPS/Register/register[15][1] ), .QN(n999)
         );
  DFFRX1 \i_MIPS/Register/register_reg[15][2]  ( .D(\i_MIPS/Register/n630 ), 
        .CK(clk), .RN(n5766), .Q(\i_MIPS/Register/register[15][2] ), .QN(n952)
         );
  DFFRX1 \i_MIPS/Register/register_reg[15][3]  ( .D(\i_MIPS/Register/n631 ), 
        .CK(clk), .RN(n5766), .Q(\i_MIPS/Register/register[15][3] ), .QN(n874)
         );
  DFFRX1 \i_MIPS/Register/register_reg[15][4]  ( .D(\i_MIPS/Register/n632 ), 
        .CK(clk), .RN(n5766), .Q(\i_MIPS/Register/register[15][4] ), .QN(n876)
         );
  DFFRX1 \i_MIPS/Register/register_reg[15][5]  ( .D(\i_MIPS/Register/n633 ), 
        .CK(clk), .RN(n5766), .Q(\i_MIPS/Register/register[15][5] ), .QN(n877)
         );
  DFFRX1 \i_MIPS/Register/register_reg[15][6]  ( .D(\i_MIPS/Register/n634 ), 
        .CK(clk), .RN(n5766), .Q(\i_MIPS/Register/register[15][6] ), .QN(n954)
         );
  DFFRX1 \i_MIPS/Register/register_reg[15][7]  ( .D(\i_MIPS/Register/n635 ), 
        .CK(clk), .RN(n5766), .Q(\i_MIPS/Register/register[15][7] ), .QN(n982)
         );
  DFFRX1 \i_MIPS/Register/register_reg[15][8]  ( .D(\i_MIPS/Register/n636 ), 
        .CK(clk), .RN(n5765), .Q(\i_MIPS/Register/register[15][8] ), .QN(n916)
         );
  DFFRX1 \i_MIPS/Register/register_reg[15][9]  ( .D(\i_MIPS/Register/n637 ), 
        .CK(clk), .RN(n5765), .Q(\i_MIPS/Register/register[15][9] ), .QN(n872)
         );
  DFFRX1 \i_MIPS/Register/register_reg[15][10]  ( .D(\i_MIPS/Register/n638 ), 
        .CK(clk), .RN(n5765), .Q(\i_MIPS/Register/register[15][10] ), .QN(n942) );
  DFFRX1 \i_MIPS/Register/register_reg[15][11]  ( .D(\i_MIPS/Register/n639 ), 
        .CK(clk), .RN(n5765), .Q(\i_MIPS/Register/register[15][11] ), .QN(n941) );
  DFFRX1 \i_MIPS/Register/register_reg[15][12]  ( .D(\i_MIPS/Register/n640 ), 
        .CK(clk), .RN(n5765), .Q(\i_MIPS/Register/register[15][12] ), .QN(n990) );
  DFFRX1 \i_MIPS/Register/register_reg[15][13]  ( .D(\i_MIPS/Register/n641 ), 
        .CK(clk), .RN(n5765), .Q(\i_MIPS/Register/register[15][13] ), .QN(n949) );
  DFFRX1 \i_MIPS/Register/register_reg[15][14]  ( .D(\i_MIPS/Register/n642 ), 
        .CK(clk), .RN(n5765), .Q(\i_MIPS/Register/register[15][14] ), .QN(n436) );
  DFFRX1 \i_MIPS/Register/register_reg[15][15]  ( .D(\i_MIPS/Register/n643 ), 
        .CK(clk), .RN(n5765), .Q(\i_MIPS/Register/register[15][15] ), .QN(n991) );
  DFFRX1 \i_MIPS/Register/register_reg[15][16]  ( .D(\i_MIPS/Register/n644 ), 
        .CK(clk), .RN(n5765), .Q(\i_MIPS/Register/register[15][16] ), .QN(
        n1003) );
  DFFRX1 \i_MIPS/Register/register_reg[15][17]  ( .D(\i_MIPS/Register/n645 ), 
        .CK(clk), .RN(n5765), .Q(\i_MIPS/Register/register[15][17] ), .QN(n908) );
  DFFRX1 \i_MIPS/Register/register_reg[15][18]  ( .D(\i_MIPS/Register/n646 ), 
        .CK(clk), .RN(n5765), .Q(\i_MIPS/Register/register[15][18] ), .QN(n871) );
  DFFRX1 \i_MIPS/Register/register_reg[15][20]  ( .D(\i_MIPS/Register/n648 ), 
        .CK(clk), .RN(n5764), .Q(\i_MIPS/Register/register[15][20] ), .QN(n947) );
  DFFRX1 \i_MIPS/Register/register_reg[15][21]  ( .D(\i_MIPS/Register/n649 ), 
        .CK(clk), .RN(n5764), .Q(\i_MIPS/Register/register[15][21] ), .QN(n937) );
  DFFRX1 \i_MIPS/Register/register_reg[15][22]  ( .D(\i_MIPS/Register/n650 ), 
        .CK(clk), .RN(n5764), .Q(\i_MIPS/Register/register[15][22] ), .QN(n905) );
  DFFRX1 \i_MIPS/Register/register_reg[15][23]  ( .D(\i_MIPS/Register/n651 ), 
        .CK(clk), .RN(n5764), .Q(\i_MIPS/Register/register[15][23] ), .QN(n873) );
  DFFRX1 \i_MIPS/Register/register_reg[15][24]  ( .D(\i_MIPS/Register/n652 ), 
        .CK(clk), .RN(n5764), .Q(\i_MIPS/Register/register[15][24] ), .QN(n432) );
  DFFRX1 \i_MIPS/Register/register_reg[15][25]  ( .D(\i_MIPS/Register/n653 ), 
        .CK(clk), .RN(n5764), .Q(\i_MIPS/Register/register[15][25] ), .QN(
        n2443) );
  DFFRX1 \i_MIPS/Register/register_reg[15][26]  ( .D(\i_MIPS/Register/n654 ), 
        .CK(clk), .RN(n5764), .Q(\i_MIPS/Register/register[15][26] ), .QN(n914) );
  DFFRX1 \i_MIPS/Register/register_reg[15][28]  ( .D(\i_MIPS/Register/n656 ), 
        .CK(clk), .RN(n5764), .Q(\i_MIPS/Register/register[15][28] ), .QN(n875) );
  DFFRX1 \i_MIPS/Register/register_reg[15][29]  ( .D(\i_MIPS/Register/n657 ), 
        .CK(clk), .RN(n5764), .Q(\i_MIPS/Register/register[15][29] ), .QN(n911) );
  DFFRX1 \i_MIPS/Register/register_reg[13][0]  ( .D(\i_MIPS/Register/n692 ), 
        .CK(clk), .RN(n5761), .Q(\i_MIPS/Register/register[13][0] ), .QN(n299)
         );
  DFFRX1 \i_MIPS/Register/register_reg[13][1]  ( .D(\i_MIPS/Register/n693 ), 
        .CK(clk), .RN(n5761), .Q(\i_MIPS/Register/register[13][1] ), .QN(n1001) );
  DFFRX1 \i_MIPS/Register/register_reg[13][2]  ( .D(\i_MIPS/Register/n694 ), 
        .CK(clk), .RN(n5761), .Q(\i_MIPS/Register/register[13][2] ), .QN(n953)
         );
  DFFRX1 \i_MIPS/Register/register_reg[13][3]  ( .D(\i_MIPS/Register/n695 ), 
        .CK(clk), .RN(n5760), .Q(\i_MIPS/Register/register[13][3] ), .QN(n452)
         );
  DFFRX1 \i_MIPS/Register/register_reg[13][4]  ( .D(\i_MIPS/Register/n696 ), 
        .CK(clk), .RN(n5760), .Q(\i_MIPS/Register/register[13][4] ), .QN(n869)
         );
  DFFRX1 \i_MIPS/Register/register_reg[13][5]  ( .D(\i_MIPS/Register/n697 ), 
        .CK(clk), .RN(n5760), .Q(\i_MIPS/Register/register[13][5] ), .QN(n870)
         );
  DFFRX1 \i_MIPS/Register/register_reg[13][6]  ( .D(\i_MIPS/Register/n698 ), 
        .CK(clk), .RN(n5760), .Q(\i_MIPS/Register/register[13][6] ), .QN(n956)
         );
  DFFRX1 \i_MIPS/Register/register_reg[13][7]  ( .D(\i_MIPS/Register/n699 ), 
        .CK(clk), .RN(n5760), .Q(\i_MIPS/Register/register[13][7] ), .QN(n456)
         );
  DFFRX1 \i_MIPS/Register/register_reg[13][8]  ( .D(\i_MIPS/Register/n700 ), 
        .CK(clk), .RN(n5760), .Q(\i_MIPS/Register/register[13][8] ), .QN(n867)
         );
  DFFRX1 \i_MIPS/Register/register_reg[13][9]  ( .D(\i_MIPS/Register/n701 ), 
        .CK(clk), .RN(n5760), .Q(\i_MIPS/Register/register[13][9] ), .QN(n638)
         );
  DFFRX1 \i_MIPS/Register/register_reg[13][10]  ( .D(\i_MIPS/Register/n702 ), 
        .CK(clk), .RN(n5760), .Q(\i_MIPS/Register/register[13][10] ), .QN(n289) );
  DFFRX1 \i_MIPS/Register/register_reg[13][11]  ( .D(\i_MIPS/Register/n703 ), 
        .CK(clk), .RN(n5760), .Q(\i_MIPS/Register/register[13][11] ), .QN(n297) );
  DFFRX1 \i_MIPS/Register/register_reg[13][12]  ( .D(\i_MIPS/Register/n704 ), 
        .CK(clk), .RN(n5760), .Q(\i_MIPS/Register/register[13][12] ), .QN(n292) );
  DFFRX1 \i_MIPS/Register/register_reg[13][13]  ( .D(\i_MIPS/Register/n705 ), 
        .CK(clk), .RN(n5760), .Q(\i_MIPS/Register/register[13][13] ), .QN(n440) );
  DFFRX1 \i_MIPS/Register/register_reg[13][14]  ( .D(\i_MIPS/Register/n706 ), 
        .CK(clk), .RN(n5760), .Q(\i_MIPS/Register/register[13][14] ), .QN(n288) );
  DFFRX1 \i_MIPS/Register/register_reg[13][15]  ( .D(\i_MIPS/Register/n707 ), 
        .CK(clk), .RN(n5759), .Q(\i_MIPS/Register/register[13][15] ), .QN(n293) );
  DFFRX1 \i_MIPS/Register/register_reg[13][16]  ( .D(\i_MIPS/Register/n708 ), 
        .CK(clk), .RN(n5759), .Q(\i_MIPS/Register/register[13][16] ), .QN(n459) );
  DFFRX1 \i_MIPS/Register/register_reg[13][17]  ( .D(\i_MIPS/Register/n709 ), 
        .CK(clk), .RN(n5759), .Q(\i_MIPS/Register/register[13][17] ), .QN(n457) );
  DFFRX1 \i_MIPS/Register/register_reg[13][18]  ( .D(\i_MIPS/Register/n710 ), 
        .CK(clk), .RN(n5759), .Q(\i_MIPS/Register/register[13][18] ), .QN(n451) );
  DFFRX1 \i_MIPS/Register/register_reg[13][20]  ( .D(\i_MIPS/Register/n712 ), 
        .CK(clk), .RN(n5759), .Q(\i_MIPS/Register/register[13][20] ), .QN(n469) );
  DFFRX1 \i_MIPS/Register/register_reg[13][21]  ( .D(\i_MIPS/Register/n713 ), 
        .CK(clk), .RN(n5759), .Q(\i_MIPS/Register/register[13][21] ), .QN(n987) );
  DFFRX1 \i_MIPS/Register/register_reg[13][22]  ( .D(\i_MIPS/Register/n714 ), 
        .CK(clk), .RN(n5759), .Q(\i_MIPS/Register/register[13][22] ), .QN(n981) );
  DFFRX1 \i_MIPS/Register/register_reg[13][23]  ( .D(\i_MIPS/Register/n715 ), 
        .CK(clk), .RN(n5759), .Q(\i_MIPS/Register/register[13][23] ), .QN(n882) );
  DFFRX1 \i_MIPS/Register/register_reg[13][24]  ( .D(\i_MIPS/Register/n716 ), 
        .CK(clk), .RN(n5759), .Q(\i_MIPS/Register/register[13][24] ), .QN(n453) );
  DFFRX1 \i_MIPS/Register/register_reg[13][25]  ( .D(\i_MIPS/Register/n717 ), 
        .CK(clk), .RN(n5759), .Q(\i_MIPS/Register/register[13][25] ), .QN(n448) );
  DFFRX1 \i_MIPS/Register/register_reg[13][26]  ( .D(\i_MIPS/Register/n718 ), 
        .CK(clk), .RN(n5759), .Q(\i_MIPS/Register/register[13][26] ), .QN(n471) );
  DFFRX1 \i_MIPS/Register/register_reg[13][28]  ( .D(\i_MIPS/Register/n720 ), 
        .CK(clk), .RN(n5758), .Q(\i_MIPS/Register/register[13][28] ), .QN(n449) );
  DFFRX1 \i_MIPS/Register/register_reg[13][29]  ( .D(\i_MIPS/Register/n721 ), 
        .CK(clk), .RN(n5758), .Q(\i_MIPS/Register/register[13][29] ), .QN(n476) );
  DFFRX1 \i_MIPS/Register/register_reg[12][0]  ( .D(\i_MIPS/Register/n724 ), 
        .CK(clk), .RN(n5758), .Q(\i_MIPS/Register/register[12][0] ), .QN(n335)
         );
  DFFRX1 \i_MIPS/Register/register_reg[12][1]  ( .D(\i_MIPS/Register/n725 ), 
        .CK(clk), .RN(n5758), .Q(\i_MIPS/Register/register[12][1] ), .QN(n969)
         );
  DFFRX1 \i_MIPS/Register/register_reg[12][2]  ( .D(\i_MIPS/Register/n726 ), 
        .CK(clk), .RN(n5758), .Q(\i_MIPS/Register/register[12][2] ), .QN(n938)
         );
  DFFRX1 \i_MIPS/Register/register_reg[12][3]  ( .D(\i_MIPS/Register/n727 ), 
        .CK(clk), .RN(n5758), .Q(\i_MIPS/Register/register[12][3] ), .QN(n975)
         );
  DFFRX1 \i_MIPS/Register/register_reg[12][4]  ( .D(\i_MIPS/Register/n728 ), 
        .CK(clk), .RN(n5758), .Q(\i_MIPS/Register/register[12][4] ), .QN(n865)
         );
  DFFRX1 \i_MIPS/Register/register_reg[12][6]  ( .D(\i_MIPS/Register/n730 ), 
        .CK(clk), .RN(n5758), .Q(\i_MIPS/Register/register[12][6] ), .QN(n972)
         );
  DFFRX1 \i_MIPS/Register/register_reg[12][7]  ( .D(\i_MIPS/Register/n731 ), 
        .CK(clk), .RN(n5757), .Q(\i_MIPS/Register/register[12][7] ), .QN(n863)
         );
  DFFRX1 \i_MIPS/Register/register_reg[12][9]  ( .D(\i_MIPS/Register/n733 ), 
        .CK(clk), .RN(n5757), .Q(\i_MIPS/Register/register[12][9] ), .QN(n862)
         );
  DFFRX1 \i_MIPS/Register/register_reg[12][10]  ( .D(\i_MIPS/Register/n734 ), 
        .CK(clk), .RN(n5757), .Q(\i_MIPS/Register/register[12][10] ), .QN(n334) );
  DFFRX1 \i_MIPS/Register/register_reg[12][13]  ( .D(\i_MIPS/Register/n737 ), 
        .CK(clk), .RN(n5757), .Q(\i_MIPS/Register/register[12][13] ), .QN(n970) );
  DFFRX1 \i_MIPS/Register/register_reg[12][14]  ( .D(\i_MIPS/Register/n738 ), 
        .CK(clk), .RN(n5757), .Q(\i_MIPS/Register/register[12][14] ), .QN(n381) );
  DFFRX1 \i_MIPS/Register/register_reg[12][15]  ( .D(\i_MIPS/Register/n739 ), 
        .CK(clk), .RN(n5757), .Q(\i_MIPS/Register/register[12][15] ), .QN(n401) );
  DFFRX1 \i_MIPS/Register/register_reg[12][16]  ( .D(\i_MIPS/Register/n740 ), 
        .CK(clk), .RN(n5757), .Q(\i_MIPS/Register/register[12][16] ), .QN(n973) );
  DFFRX1 \i_MIPS/Register/register_reg[12][18]  ( .D(\i_MIPS/Register/n742 ), 
        .CK(clk), .RN(n5757), .Q(\i_MIPS/Register/register[12][18] ), .QN(n860) );
  DFFRX1 \i_MIPS/Register/register_reg[12][20]  ( .D(\i_MIPS/Register/n744 ), 
        .CK(clk), .RN(n5756), .Q(\i_MIPS/Register/register[12][20] ), .QN(n971) );
  DFFRX1 \i_MIPS/Register/register_reg[12][21]  ( .D(\i_MIPS/Register/n745 ), 
        .CK(clk), .RN(n5756), .Q(\i_MIPS/Register/register[12][21] ), .QN(
        n1020) );
  DFFRX1 \i_MIPS/Register/register_reg[12][23]  ( .D(\i_MIPS/Register/n747 ), 
        .CK(clk), .RN(n5766), .Q(\i_MIPS/Register/register[12][23] ), .QN(n861) );
  DFFRX1 \i_MIPS/Register/register_reg[12][25]  ( .D(\i_MIPS/Register/n749 ), 
        .CK(clk), .RN(n5656), .Q(\i_MIPS/Register/register[12][25] ), .QN(n864) );
  DFFRX1 \i_MIPS/Register/register_reg[12][26]  ( .D(\i_MIPS/Register/n750 ), 
        .CK(clk), .RN(n5656), .Q(\i_MIPS/Register/register[12][26] ), .QN(n976) );
  DFFRX1 \i_MIPS/Register/register_reg[12][28]  ( .D(\i_MIPS/Register/n752 ), 
        .CK(clk), .RN(n5656), .Q(\i_MIPS/Register/register[12][28] ), .QN(n974) );
  DFFRX1 \i_MIPS/Register/register_reg[11][0]  ( .D(\i_MIPS/Register/n756 ), 
        .CK(clk), .RN(n5656), .Q(\i_MIPS/Register/register[11][0] ), .QN(n391)
         );
  DFFRX1 \i_MIPS/Register/register_reg[11][1]  ( .D(\i_MIPS/Register/n757 ), 
        .CK(clk), .RN(n5656), .Q(\i_MIPS/Register/register[11][1] ), .QN(n1000) );
  DFFRX1 \i_MIPS/Register/register_reg[11][2]  ( .D(\i_MIPS/Register/n758 ), 
        .CK(clk), .RN(n5656), .Q(\i_MIPS/Register/register[11][2] ), .QN(n1007) );
  DFFRX1 \i_MIPS/Register/register_reg[11][3]  ( .D(\i_MIPS/Register/n759 ), 
        .CK(clk), .RN(n5656), .Q(\i_MIPS/Register/register[11][3] ), .QN(n354)
         );
  DFFRX1 \i_MIPS/Register/register_reg[11][4]  ( .D(\i_MIPS/Register/n760 ), 
        .CK(clk), .RN(n5656), .Q(\i_MIPS/Register/register[11][4] ), .QN(n918)
         );
  DFFRX1 \i_MIPS/Register/register_reg[11][5]  ( .D(\i_MIPS/Register/n761 ), 
        .CK(clk), .RN(n5655), .Q(\i_MIPS/Register/register[11][5] ), .QN(n920)
         );
  DFFRX1 \i_MIPS/Register/register_reg[11][6]  ( .D(\i_MIPS/Register/n762 ), 
        .CK(clk), .RN(n5655), .Q(\i_MIPS/Register/register[11][6] ), .QN(n955)
         );
  DFFRX1 \i_MIPS/Register/register_reg[11][7]  ( .D(\i_MIPS/Register/n763 ), 
        .CK(clk), .RN(n5655), .Q(\i_MIPS/Register/register[11][7] ), .QN(n902)
         );
  DFFRX1 \i_MIPS/Register/register_reg[11][8]  ( .D(\i_MIPS/Register/n764 ), 
        .CK(clk), .RN(n5655), .Q(\i_MIPS/Register/register[11][8] ), .QN(n915)
         );
  DFFRX1 \i_MIPS/Register/register_reg[11][9]  ( .D(\i_MIPS/Register/n765 ), 
        .CK(clk), .RN(n5655), .Q(\i_MIPS/Register/register[11][9] ), .QN(n355)
         );
  DFFRX1 \i_MIPS/Register/register_reg[11][10]  ( .D(\i_MIPS/Register/n766 ), 
        .CK(clk), .RN(n5655), .Q(\i_MIPS/Register/register[11][10] ), .QN(n371) );
  DFFRX1 \i_MIPS/Register/register_reg[11][11]  ( .D(\i_MIPS/Register/n767 ), 
        .CK(clk), .RN(n5655), .Q(\i_MIPS/Register/register[11][11] ), .QN(n387) );
  DFFRX1 \i_MIPS/Register/register_reg[11][12]  ( .D(\i_MIPS/Register/n768 ), 
        .CK(clk), .RN(n5655), .Q(\i_MIPS/Register/register[11][12] ), .QN(n386) );
  DFFRX1 \i_MIPS/Register/register_reg[11][13]  ( .D(\i_MIPS/Register/n769 ), 
        .CK(clk), .RN(n5655), .Q(\i_MIPS/Register/register[11][13] ), .QN(
        n1006) );
  DFFRX1 \i_MIPS/Register/register_reg[11][14]  ( .D(\i_MIPS/Register/n770 ), 
        .CK(clk), .RN(n5655), .Q(\i_MIPS/Register/register[11][14] ), .QN(n326) );
  DFFRX1 \i_MIPS/Register/register_reg[11][15]  ( .D(\i_MIPS/Register/n771 ), 
        .CK(clk), .RN(n5655), .Q(\i_MIPS/Register/register[11][15] ), .QN(n389) );
  DFFRX1 \i_MIPS/Register/register_reg[11][16]  ( .D(\i_MIPS/Register/n772 ), 
        .CK(clk), .RN(n5655), .Q(\i_MIPS/Register/register[11][16] ), .QN(
        n1004) );
  DFFRX1 \i_MIPS/Register/register_reg[11][17]  ( .D(\i_MIPS/Register/n773 ), 
        .CK(clk), .RN(n5654), .Q(\i_MIPS/Register/register[11][17] ), .QN(n907) );
  DFFRX1 \i_MIPS/Register/register_reg[11][18]  ( .D(\i_MIPS/Register/n774 ), 
        .CK(clk), .RN(n5654), .Q(\i_MIPS/Register/register[11][18] ), .QN(n367) );
  DFFRX1 \i_MIPS/Register/register_reg[11][20]  ( .D(\i_MIPS/Register/n776 ), 
        .CK(clk), .RN(n5654), .Q(\i_MIPS/Register/register[11][20] ), .QN(n997) );
  DFFRX1 \i_MIPS/Register/register_reg[11][21]  ( .D(\i_MIPS/Register/n777 ), 
        .CK(clk), .RN(n5654), .Q(\i_MIPS/Register/register[11][21] ), .QN(n645) );
  DFFRX1 \i_MIPS/Register/register_reg[11][22]  ( .D(\i_MIPS/Register/n778 ), 
        .CK(clk), .RN(n5654), .Q(\i_MIPS/Register/register[11][22] ), .QN(n904) );
  DFFRX1 \i_MIPS/Register/register_reg[11][23]  ( .D(\i_MIPS/Register/n779 ), 
        .CK(clk), .RN(n5654), .Q(\i_MIPS/Register/register[11][23] ), .QN(n644) );
  DFFRX1 \i_MIPS/Register/register_reg[11][24]  ( .D(\i_MIPS/Register/n780 ), 
        .CK(clk), .RN(n5654), .Q(\i_MIPS/Register/register[11][24] ), .QN(n323) );
  DFFRX1 \i_MIPS/Register/register_reg[11][25]  ( .D(\i_MIPS/Register/n781 ), 
        .CK(clk), .RN(n5654), .Q(\i_MIPS/Register/register[11][25] ), .QN(n989) );
  DFFRX1 \i_MIPS/Register/register_reg[11][26]  ( .D(\i_MIPS/Register/n782 ), 
        .CK(clk), .RN(n5654), .Q(\i_MIPS/Register/register[11][26] ), .QN(n913) );
  DFFRX1 \i_MIPS/Register/register_reg[11][28]  ( .D(\i_MIPS/Register/n784 ), 
        .CK(clk), .RN(n5654), .Q(\i_MIPS/Register/register[11][28] ), .QN(n383) );
  DFFRX1 \i_MIPS/Register/register_reg[11][29]  ( .D(\i_MIPS/Register/n785 ), 
        .CK(clk), .RN(n5653), .Q(\i_MIPS/Register/register[11][29] ), .QN(n910) );
  DFFRX1 \i_MIPS/Register/register_reg[9][0]  ( .D(\i_MIPS/Register/n820 ), 
        .CK(clk), .RN(n5650), .Q(\i_MIPS/Register/register[9][0] ), .QN(n351)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][1]  ( .D(\i_MIPS/Register/n821 ), 
        .CK(clk), .RN(n5650), .Q(\i_MIPS/Register/register[9][1] ), .QN(n927)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][2]  ( .D(\i_MIPS/Register/n822 ), 
        .CK(clk), .RN(n5650), .Q(\i_MIPS/Register/register[9][2] ), .QN(n965)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][3]  ( .D(\i_MIPS/Register/n823 ), 
        .CK(clk), .RN(n5650), .Q(\i_MIPS/Register/register[9][3] ), .QN(n368)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][4]  ( .D(\i_MIPS/Register/n824 ), 
        .CK(clk), .RN(n5650), .Q(\i_MIPS/Register/register[9][4] ), .QN(n879)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][5]  ( .D(\i_MIPS/Register/n825 ), 
        .CK(clk), .RN(n5650), .Q(\i_MIPS/Register/register[9][5] ), .QN(n880)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][6]  ( .D(\i_MIPS/Register/n826 ), 
        .CK(clk), .RN(n5650), .Q(\i_MIPS/Register/register[9][6] ), .QN(n966)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][7]  ( .D(\i_MIPS/Register/n827 ), 
        .CK(clk), .RN(n5650), .Q(\i_MIPS/Register/register[9][7] ), .QN(n935)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][8]  ( .D(\i_MIPS/Register/n828 ), 
        .CK(clk), .RN(n5650), .Q(\i_MIPS/Register/register[9][8] ), .QN(n925)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][9]  ( .D(\i_MIPS/Register/n829 ), 
        .CK(clk), .RN(n5650), .Q(\i_MIPS/Register/register[9][9] ), .QN(n343)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][10]  ( .D(\i_MIPS/Register/n830 ), 
        .CK(clk), .RN(n5650), .Q(\i_MIPS/Register/register[9][10] ), .QN(n331)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][11]  ( .D(\i_MIPS/Register/n831 ), 
        .CK(clk), .RN(n5650), .Q(\i_MIPS/Register/register[9][11] ), .QN(n350)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][12]  ( .D(\i_MIPS/Register/n832 ), 
        .CK(clk), .RN(n5649), .Q(\i_MIPS/Register/register[9][12] ), .QN(n329)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][13]  ( .D(\i_MIPS/Register/n833 ), 
        .CK(clk), .RN(n5649), .Q(\i_MIPS/Register/register[9][13] ), .QN(n852)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][14]  ( .D(\i_MIPS/Register/n834 ), 
        .CK(clk), .RN(n5649), .Q(\i_MIPS/Register/register[9][14] ), .QN(n378)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][15]  ( .D(\i_MIPS/Register/n835 ), 
        .CK(clk), .RN(n5649), .Q(\i_MIPS/Register/register[9][15] ), .QN(n366)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][16]  ( .D(\i_MIPS/Register/n836 ), 
        .CK(clk), .RN(n5649), .Q(\i_MIPS/Register/register[9][16] ), .QN(n855)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][17]  ( .D(\i_MIPS/Register/n837 ), 
        .CK(clk), .RN(n5649), .Q(\i_MIPS/Register/register[9][17] ), .QN(n922)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][18]  ( .D(\i_MIPS/Register/n838 ), 
        .CK(clk), .RN(n5649), .Q(\i_MIPS/Register/register[9][18] ), .QN(n373)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][20]  ( .D(\i_MIPS/Register/n840 ), 
        .CK(clk), .RN(n5649), .Q(\i_MIPS/Register/register[9][20] ), .QN(n376)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][21]  ( .D(\i_MIPS/Register/n841 ), 
        .CK(clk), .RN(n5649), .Q(\i_MIPS/Register/register[9][21] ), .QN(n374)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][22]  ( .D(\i_MIPS/Register/n842 ), 
        .CK(clk), .RN(n5649), .Q(\i_MIPS/Register/register[9][22] ), .QN(n362)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][23]  ( .D(\i_MIPS/Register/n843 ), 
        .CK(clk), .RN(n5649), .Q(\i_MIPS/Register/register[9][23] ), .QN(n295)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][24]  ( .D(\i_MIPS/Register/n844 ), 
        .CK(clk), .RN(n5648), .Q(\i_MIPS/Register/register[9][24] ), .QN(n346)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][25]  ( .D(\i_MIPS/Register/n845 ), 
        .CK(clk), .RN(n5648), .Q(\i_MIPS/Register/register[9][25] ), .QN(n348)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][26]  ( .D(\i_MIPS/Register/n846 ), 
        .CK(clk), .RN(n5648), .Q(\i_MIPS/Register/register[9][26] ), .QN(n364)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][28]  ( .D(\i_MIPS/Register/n848 ), 
        .CK(clk), .RN(n5648), .Q(\i_MIPS/Register/register[9][28] ), .QN(n344)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][29]  ( .D(\i_MIPS/Register/n849 ), 
        .CK(clk), .RN(n5648), .Q(\i_MIPS/Register/register[9][29] ), .QN(n984)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][0]  ( .D(\i_MIPS/Register/n852 ), 
        .CK(clk), .RN(n5648), .Q(\i_MIPS/Register/register[8][0] ), .QN(n899)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][1]  ( .D(\i_MIPS/Register/n853 ), 
        .CK(clk), .RN(n5648), .Q(\i_MIPS/Register/register[8][1] ), .QN(n338)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][2]  ( .D(\i_MIPS/Register/n854 ), 
        .CK(clk), .RN(n5648), .Q(\i_MIPS/Register/register[8][2] ), .QN(n443)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][3]  ( .D(\i_MIPS/Register/n855 ), 
        .CK(clk), .RN(n5648), .Q(\i_MIPS/Register/register[8][3] ), .QN(n885)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][4]  ( .D(\i_MIPS/Register/n856 ), 
        .CK(clk), .RN(n5647), .Q(\i_MIPS/Register/register[8][4] ), .QN(n464)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][6]  ( .D(\i_MIPS/Register/n858 ), 
        .CK(clk), .RN(n5647), .Q(\i_MIPS/Register/register[8][6] ), .QN(n444)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][7]  ( .D(\i_MIPS/Register/n859 ), 
        .CK(clk), .RN(n5647), .Q(\i_MIPS/Register/register[8][7] ), .QN(n357)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][8]  ( .D(\i_MIPS/Register/n860 ), 
        .CK(clk), .RN(n5647), .Q(\i_MIPS/Register/register[8][8] ), .QN(n933)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][9]  ( .D(\i_MIPS/Register/n861 ), 
        .CK(clk), .RN(n5647), .Q(\i_MIPS/Register/register[8][9] ), .QN(n884)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][10]  ( .D(\i_MIPS/Register/n862 ), 
        .CK(clk), .RN(n5647), .Q(\i_MIPS/Register/register[8][10] ), .QN(n856)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][13]  ( .D(\i_MIPS/Register/n865 ), 
        .CK(clk), .RN(n5647), .Q(\i_MIPS/Register/register[8][13] ), .QN(n341)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][14]  ( .D(\i_MIPS/Register/n866 ), 
        .CK(clk), .RN(n5647), .Q(\i_MIPS/Register/register[8][14] ), .QN(n641)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][15]  ( .D(\i_MIPS/Register/n867 ), 
        .CK(clk), .RN(n5647), .Q(\i_MIPS/Register/register[8][15] ), .QN(n897)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][16]  ( .D(\i_MIPS/Register/n868 ), 
        .CK(clk), .RN(n5651), .Q(\i_MIPS/Register/register[8][16] ), .QN(n339)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][18]  ( .D(\i_MIPS/Register/n870 ), 
        .CK(clk), .RN(n5666), .Q(\i_MIPS/Register/register[8][18] ), .QN(n858)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][20]  ( .D(\i_MIPS/Register/n872 ), 
        .CK(clk), .RN(n5666), .Q(\i_MIPS/Register/register[8][20] ), .QN(n967)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][21]  ( .D(\i_MIPS/Register/n873 ), 
        .CK(clk), .RN(n5666), .Q(\i_MIPS/Register/register[8][21] ), .QN(n460)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][23]  ( .D(\i_MIPS/Register/n875 ), 
        .CK(clk), .RN(n5666), .Q(\i_MIPS/Register/register[8][23] ), .QN(n928)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][24]  ( .D(\i_MIPS/Register/n876 ), 
        .CK(clk), .RN(n5666), .Q(\i_MIPS/Register/register[8][24] ), .QN(n887)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][25]  ( .D(\i_MIPS/Register/n877 ), 
        .CK(clk), .RN(n5666), .Q(\i_MIPS/Register/register[8][25] ), .QN(n462)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][26]  ( .D(\i_MIPS/Register/n878 ), 
        .CK(clk), .RN(n5666), .Q(\i_MIPS/Register/register[8][26] ), .QN(n946)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][28]  ( .D(\i_MIPS/Register/n880 ), 
        .CK(clk), .RN(n5665), .Q(\i_MIPS/Register/register[8][28] ), .QN(n883)
         );
  DFFRX1 \i_MIPS/Register/register_reg[23][0]  ( .D(\i_MIPS/Register/n372 ), 
        .CK(clk), .RN(n5768), .Q(\i_MIPS/Register/register[23][0] ), .QN(n2515) );
  DFFRX1 \i_MIPS/Register/register_reg[23][1]  ( .D(\i_MIPS/Register/n373 ), 
        .CK(clk), .RN(n5768), .Q(\i_MIPS/Register/register[23][1] ), .QN(n2519) );
  DFFRX1 \i_MIPS/Register/register_reg[23][2]  ( .D(\i_MIPS/Register/n374 ), 
        .CK(clk), .RN(n5767), .Q(\i_MIPS/Register/register[23][2] ), .QN(n2462) );
  DFFRX1 \i_MIPS/Register/register_reg[23][3]  ( .D(\i_MIPS/Register/n375 ), 
        .CK(clk), .RN(n5767), .Q(\i_MIPS/Register/register[23][3] ), .QN(n2616) );
  DFFRX1 \i_MIPS/Register/register_reg[23][4]  ( .D(\i_MIPS/Register/n376 ), 
        .CK(clk), .RN(n5767), .Q(\i_MIPS/Register/register[23][4] ), .QN(n2622) );
  DFFRX1 \i_MIPS/Register/register_reg[23][5]  ( .D(\i_MIPS/Register/n377 ), 
        .CK(clk), .RN(n5767), .Q(\i_MIPS/Register/register[23][5] ), .QN(n2625) );
  DFFRX1 \i_MIPS/Register/register_reg[23][6]  ( .D(\i_MIPS/Register/n378 ), 
        .CK(clk), .RN(n5767), .Q(\i_MIPS/Register/register[23][6] ), .QN(n2465) );
  DFFRX1 \i_MIPS/Register/register_reg[23][7]  ( .D(\i_MIPS/Register/n379 ), 
        .CK(clk), .RN(n5767), .Q(\i_MIPS/Register/register[23][7] ), .QN(n2497) );
  DFFRX1 \i_MIPS/Register/register_reg[23][8]  ( .D(\i_MIPS/Register/n380 ), 
        .CK(clk), .RN(n5767), .Q(\i_MIPS/Register/register[23][8] ), .QN(n2617) );
  DFFRX1 \i_MIPS/Register/register_reg[23][9]  ( .D(\i_MIPS/Register/n381 ), 
        .CK(clk), .RN(n5767), .Q(\i_MIPS/Register/register[23][9] ), .QN(n2601) );
  DFFRX1 \i_MIPS/Register/register_reg[23][10]  ( .D(\i_MIPS/Register/n382 ), 
        .CK(clk), .RN(n5767), .Q(\i_MIPS/Register/register[23][10] ), .QN(
        n2452) );
  DFFRX1 \i_MIPS/Register/register_reg[23][11]  ( .D(\i_MIPS/Register/n383 ), 
        .CK(clk), .RN(n5767), .Q(\i_MIPS/Register/register[23][11] ), .QN(
        n2512) );
  DFFRX1 \i_MIPS/Register/register_reg[23][12]  ( .D(\i_MIPS/Register/n384 ), 
        .CK(clk), .RN(n5767), .Q(\i_MIPS/Register/register[23][12] ), .QN(
        n2633) );
  DFFRX1 \i_MIPS/Register/register_reg[23][13]  ( .D(\i_MIPS/Register/n385 ), 
        .CK(clk), .RN(n5767), .Q(\i_MIPS/Register/register[23][13] ), .QN(
        n2460) );
  DFFRX1 \i_MIPS/Register/register_reg[23][14]  ( .D(\i_MIPS/Register/n386 ), 
        .CK(clk), .RN(n5766), .Q(\i_MIPS/Register/register[23][14] ), .QN(
        n2046) );
  DFFRX1 \i_MIPS/Register/register_reg[23][15]  ( .D(\i_MIPS/Register/n387 ), 
        .CK(clk), .RN(n5766), .Q(\i_MIPS/Register/register[23][15] ), .QN(
        n2513) );
  DFFRX1 \i_MIPS/Register/register_reg[23][16]  ( .D(\i_MIPS/Register/n388 ), 
        .CK(clk), .RN(n5766), .Q(\i_MIPS/Register/register[23][16] ), .QN(
        n2523) );
  DFFRX1 \i_MIPS/Register/register_reg[23][17]  ( .D(\i_MIPS/Register/n389 ), 
        .CK(clk), .RN(n5771), .Q(\i_MIPS/Register/register[23][17] ), .QN(
        n2500) );
  DFFRX1 \i_MIPS/Register/register_reg[23][18]  ( .D(\i_MIPS/Register/n390 ), 
        .CK(clk), .RN(n5786), .Q(\i_MIPS/Register/register[23][18] ), .QN(
        n2567) );
  DFFRX1 \i_MIPS/Register/register_reg[23][20]  ( .D(\i_MIPS/Register/n392 ), 
        .CK(clk), .RN(n5786), .Q(\i_MIPS/Register/register[23][20] ), .QN(
        n2022) );
  DFFRX1 \i_MIPS/Register/register_reg[23][21]  ( .D(\i_MIPS/Register/n393 ), 
        .CK(clk), .RN(n5786), .Q(\i_MIPS/Register/register[23][21] ), .QN(
        n2455) );
  DFFRX1 \i_MIPS/Register/register_reg[23][22]  ( .D(\i_MIPS/Register/n394 ), 
        .CK(clk), .RN(n5786), .Q(\i_MIPS/Register/register[23][22] ), .QN(
        n2603) );
  DFFRX1 \i_MIPS/Register/register_reg[23][23]  ( .D(\i_MIPS/Register/n395 ), 
        .CK(clk), .RN(n5786), .Q(\i_MIPS/Register/register[23][23] ), .QN(
        n2568) );
  DFFRX1 \i_MIPS/Register/register_reg[23][24]  ( .D(\i_MIPS/Register/n396 ), 
        .CK(clk), .RN(n5786), .Q(\i_MIPS/Register/register[23][24] ), .QN(
        n2560) );
  DFFRX1 \i_MIPS/Register/register_reg[23][25]  ( .D(\i_MIPS/Register/n397 ), 
        .CK(clk), .RN(n5786), .Q(\i_MIPS/Register/register[23][25] ), .QN(
        n2021) );
  DFFRX1 \i_MIPS/Register/register_reg[23][26]  ( .D(\i_MIPS/Register/n398 ), 
        .CK(clk), .RN(n5785), .Q(\i_MIPS/Register/register[23][26] ), .QN(
        n2613) );
  DFFRX1 \i_MIPS/Register/register_reg[23][28]  ( .D(\i_MIPS/Register/n400 ), 
        .CK(clk), .RN(n5785), .Q(\i_MIPS/Register/register[23][28] ), .QN(
        n2620) );
  DFFRX1 \i_MIPS/Register/register_reg[23][29]  ( .D(\i_MIPS/Register/n401 ), 
        .CK(clk), .RN(n5785), .Q(\i_MIPS/Register/register[23][29] ), .QN(
        n2502) );
  DFFRX1 \i_MIPS/Register/register_reg[21][0]  ( .D(\i_MIPS/Register/n436 ), 
        .CK(clk), .RN(n5782), .Q(\i_MIPS/Register/register[21][0] ), .QN(n2060) );
  DFFRX1 \i_MIPS/Register/register_reg[21][1]  ( .D(\i_MIPS/Register/n437 ), 
        .CK(clk), .RN(n5782), .Q(\i_MIPS/Register/register[21][1] ), .QN(n2521) );
  DFFRX1 \i_MIPS/Register/register_reg[21][2]  ( .D(\i_MIPS/Register/n438 ), 
        .CK(clk), .RN(n5782), .Q(\i_MIPS/Register/register[21][2] ), .QN(n2463) );
  DFFRX1 \i_MIPS/Register/register_reg[21][3]  ( .D(\i_MIPS/Register/n439 ), 
        .CK(clk), .RN(n5782), .Q(\i_MIPS/Register/register[21][3] ), .QN(n2065) );
  DFFRX1 \i_MIPS/Register/register_reg[21][4]  ( .D(\i_MIPS/Register/n440 ), 
        .CK(clk), .RN(n5782), .Q(\i_MIPS/Register/register[21][4] ), .QN(n2552) );
  DFFRX1 \i_MIPS/Register/register_reg[21][5]  ( .D(\i_MIPS/Register/n441 ), 
        .CK(clk), .RN(n5782), .Q(\i_MIPS/Register/register[21][5] ), .QN(n2591) );
  DFFRX1 \i_MIPS/Register/register_reg[21][6]  ( .D(\i_MIPS/Register/n442 ), 
        .CK(clk), .RN(n5782), .Q(\i_MIPS/Register/register[21][6] ), .QN(n2467) );
  DFFRX1 \i_MIPS/Register/register_reg[21][7]  ( .D(\i_MIPS/Register/n443 ), 
        .CK(clk), .RN(n5782), .Q(\i_MIPS/Register/register[21][7] ), .QN(n2066) );
  DFFRX1 \i_MIPS/Register/register_reg[21][8]  ( .D(\i_MIPS/Register/n444 ), 
        .CK(clk), .RN(n5782), .Q(\i_MIPS/Register/register[21][8] ), .QN(n2590) );
  DFFRX1 \i_MIPS/Register/register_reg[21][9]  ( .D(\i_MIPS/Register/n445 ), 
        .CK(clk), .RN(n5782), .Q(\i_MIPS/Register/register[21][9] ), .QN(n2040) );
  DFFRX1 \i_MIPS/Register/register_reg[21][10]  ( .D(\i_MIPS/Register/n446 ), 
        .CK(clk), .RN(n5781), .Q(\i_MIPS/Register/register[21][10] ), .QN(
        n2572) );
  DFFRX1 \i_MIPS/Register/register_reg[21][11]  ( .D(\i_MIPS/Register/n447 ), 
        .CK(clk), .RN(n5781), .Q(\i_MIPS/Register/register[21][11] ), .QN(
        n2570) );
  DFFRX1 \i_MIPS/Register/register_reg[21][12]  ( .D(\i_MIPS/Register/n448 ), 
        .CK(clk), .RN(n5781), .Q(\i_MIPS/Register/register[21][12] ), .QN(
        n2061) );
  DFFRX1 \i_MIPS/Register/register_reg[21][13]  ( .D(\i_MIPS/Register/n449 ), 
        .CK(clk), .RN(n5781), .Q(\i_MIPS/Register/register[21][13] ), .QN(
        n2020) );
  DFFRX1 \i_MIPS/Register/register_reg[21][14]  ( .D(\i_MIPS/Register/n450 ), 
        .CK(clk), .RN(n5781), .Q(\i_MIPS/Register/register[21][14] ), .QN(
        n2032) );
  DFFRX1 \i_MIPS/Register/register_reg[21][15]  ( .D(\i_MIPS/Register/n451 ), 
        .CK(clk), .RN(n5781), .Q(\i_MIPS/Register/register[21][15] ), .QN(
        n2064) );
  DFFRX1 \i_MIPS/Register/register_reg[21][16]  ( .D(\i_MIPS/Register/n452 ), 
        .CK(clk), .RN(n5781), .Q(\i_MIPS/Register/register[21][16] ), .QN(
        n2044) );
  DFFRX1 \i_MIPS/Register/register_reg[21][17]  ( .D(\i_MIPS/Register/n453 ), 
        .CK(clk), .RN(n5781), .Q(\i_MIPS/Register/register[21][17] ), .QN(
        n2217) );
  DFFRX1 \i_MIPS/Register/register_reg[21][18]  ( .D(\i_MIPS/Register/n454 ), 
        .CK(clk), .RN(n5781), .Q(\i_MIPS/Register/register[21][18] ), .QN(
        n2036) );
  DFFRX1 \i_MIPS/Register/register_reg[21][20]  ( .D(\i_MIPS/Register/n456 ), 
        .CK(clk), .RN(n5781), .Q(\i_MIPS/Register/register[21][20] ), .QN(
        n2055) );
  DFFRX1 \i_MIPS/Register/register_reg[21][21]  ( .D(\i_MIPS/Register/n457 ), 
        .CK(clk), .RN(n5780), .Q(\i_MIPS/Register/register[21][21] ), .QN(
        n2506) );
  DFFRX1 \i_MIPS/Register/register_reg[21][22]  ( .D(\i_MIPS/Register/n458 ), 
        .CK(clk), .RN(n5780), .Q(\i_MIPS/Register/register[21][22] ), .QN(
        n2059) );
  DFFRX1 \i_MIPS/Register/register_reg[21][23]  ( .D(\i_MIPS/Register/n459 ), 
        .CK(clk), .RN(n5780), .Q(\i_MIPS/Register/register[21][23] ), .QN(
        n2569) );
  DFFRX1 \i_MIPS/Register/register_reg[21][24]  ( .D(\i_MIPS/Register/n460 ), 
        .CK(clk), .RN(n5780), .Q(\i_MIPS/Register/register[21][24] ), .QN(
        n2214) );
  DFFRX1 \i_MIPS/Register/register_reg[21][25]  ( .D(\i_MIPS/Register/n461 ), 
        .CK(clk), .RN(n5780), .Q(\i_MIPS/Register/register[21][25] ), .QN(
        n2030) );
  DFFRX1 \i_MIPS/Register/register_reg[21][26]  ( .D(\i_MIPS/Register/n462 ), 
        .CK(clk), .RN(n5780), .Q(\i_MIPS/Register/register[21][26] ), .QN(
        n2057) );
  DFFRX1 \i_MIPS/Register/register_reg[21][28]  ( .D(\i_MIPS/Register/n464 ), 
        .CK(clk), .RN(n5780), .Q(\i_MIPS/Register/register[21][28] ), .QN(
        n2218) );
  DFFRX1 \i_MIPS/Register/register_reg[21][29]  ( .D(\i_MIPS/Register/n465 ), 
        .CK(clk), .RN(n5780), .Q(\i_MIPS/Register/register[21][29] ), .QN(
        n2067) );
  DFFRX1 \i_MIPS/Register/register_reg[20][0]  ( .D(\i_MIPS/Register/n468 ), 
        .CK(clk), .RN(n5780), .Q(\i_MIPS/Register/register[20][0] ), .QN(n1045) );
  DFFRX1 \i_MIPS/Register/register_reg[20][1]  ( .D(\i_MIPS/Register/n469 ), 
        .CK(clk), .RN(n5779), .Q(\i_MIPS/Register/register[20][1] ), .QN(n2535) );
  DFFRX1 \i_MIPS/Register/register_reg[20][2]  ( .D(\i_MIPS/Register/n470 ), 
        .CK(clk), .RN(n5779), .Q(\i_MIPS/Register/register[20][2] ), .QN(n2449) );
  DFFRX1 \i_MIPS/Register/register_reg[20][3]  ( .D(\i_MIPS/Register/n471 ), 
        .CK(clk), .RN(n5779), .Q(\i_MIPS/Register/register[20][3] ), .QN(n2538) );
  DFFRX1 \i_MIPS/Register/register_reg[20][4]  ( .D(\i_MIPS/Register/n472 ), 
        .CK(clk), .RN(n5779), .Q(\i_MIPS/Register/register[20][4] ), .QN(n2541) );
  DFFRX1 \i_MIPS/Register/register_reg[20][5]  ( .D(\i_MIPS/Register/n473 ), 
        .CK(clk), .RN(n5779), .Q(\i_MIPS/Register/register[20][5] ), .QN(n2543) );
  DFFRX1 \i_MIPS/Register/register_reg[20][6]  ( .D(\i_MIPS/Register/n474 ), 
        .CK(clk), .RN(n5779), .Q(\i_MIPS/Register/register[20][6] ), .QN(n2450) );
  DFFRX1 \i_MIPS/Register/register_reg[20][7]  ( .D(\i_MIPS/Register/n475 ), 
        .CK(clk), .RN(n5779), .Q(\i_MIPS/Register/register[20][7] ), .QN(n2583) );
  DFFRX1 \i_MIPS/Register/register_reg[20][8]  ( .D(\i_MIPS/Register/n476 ), 
        .CK(clk), .RN(n5779), .Q(\i_MIPS/Register/register[20][8] ), .QN(n2477) );
  DFFRX1 \i_MIPS/Register/register_reg[20][9]  ( .D(\i_MIPS/Register/n477 ), 
        .CK(clk), .RN(n5779), .Q(\i_MIPS/Register/register[20][9] ), .QN(n2539) );
  DFFRX1 \i_MIPS/Register/register_reg[20][10]  ( .D(\i_MIPS/Register/n478 ), 
        .CK(clk), .RN(n5779), .Q(\i_MIPS/Register/register[20][10] ), .QN(
        n1043) );
  DFFRX1 \i_MIPS/Register/register_reg[20][11]  ( .D(\i_MIPS/Register/n479 ), 
        .CK(clk), .RN(n5779), .Q(\i_MIPS/Register/register[20][11] ), .QN(
        n1047) );
  DFFRX1 \i_MIPS/Register/register_reg[20][12]  ( .D(\i_MIPS/Register/n480 ), 
        .CK(clk), .RN(n5779), .Q(\i_MIPS/Register/register[20][12] ), .QN(
        n1048) );
  DFFRX1 \i_MIPS/Register/register_reg[20][13]  ( .D(\i_MIPS/Register/n481 ), 
        .CK(clk), .RN(n5778), .Q(\i_MIPS/Register/register[20][13] ), .QN(
        n2584) );
  DFFRX1 \i_MIPS/Register/register_reg[20][14]  ( .D(\i_MIPS/Register/n482 ), 
        .CK(clk), .RN(n5778), .Q(\i_MIPS/Register/register[20][14] ), .QN(
        n1044) );
  DFFRX1 \i_MIPS/Register/register_reg[20][15]  ( .D(\i_MIPS/Register/n483 ), 
        .CK(clk), .RN(n5778), .Q(\i_MIPS/Register/register[20][15] ), .QN(
        n1046) );
  DFFRX1 \i_MIPS/Register/register_reg[20][16]  ( .D(\i_MIPS/Register/n484 ), 
        .CK(clk), .RN(n5778), .Q(\i_MIPS/Register/register[20][16] ), .QN(
        n2585) );
  DFFRX1 \i_MIPS/Register/register_reg[20][17]  ( .D(\i_MIPS/Register/n485 ), 
        .CK(clk), .RN(n5778), .Q(\i_MIPS/Register/register[20][17] ), .QN(
        n2544) );
  DFFRX1 \i_MIPS/Register/register_reg[20][18]  ( .D(\i_MIPS/Register/n486 ), 
        .CK(clk), .RN(n5778), .Q(\i_MIPS/Register/register[20][18] ), .QN(
        n2534) );
  DFFRX1 \i_MIPS/Register/register_reg[20][20]  ( .D(\i_MIPS/Register/n488 ), 
        .CK(clk), .RN(n5778), .Q(\i_MIPS/Register/register[20][20] ), .QN(
        n2474) );
  DFFRX1 \i_MIPS/Register/register_reg[20][21]  ( .D(\i_MIPS/Register/n489 ), 
        .CK(clk), .RN(n5778), .Q(\i_MIPS/Register/register[20][21] ), .QN(
        n2536) );
  DFFRX1 \i_MIPS/Register/register_reg[20][23]  ( .D(\i_MIPS/Register/n491 ), 
        .CK(clk), .RN(n5778), .Q(\i_MIPS/Register/register[20][23] ), .QN(
        n2537) );
  DFFRX1 \i_MIPS/Register/register_reg[20][24]  ( .D(\i_MIPS/Register/n492 ), 
        .CK(clk), .RN(n5778), .Q(\i_MIPS/Register/register[20][24] ), .QN(
        n2542) );
  DFFRX1 \i_MIPS/Register/register_reg[20][25]  ( .D(\i_MIPS/Register/n493 ), 
        .CK(clk), .RN(n5777), .Q(\i_MIPS/Register/register[20][25] ), .QN(
        n2540) );
  DFFRX1 \i_MIPS/Register/register_reg[20][26]  ( .D(\i_MIPS/Register/n494 ), 
        .CK(clk), .RN(n5777), .Q(\i_MIPS/Register/register[20][26] ), .QN(
        n2476) );
  DFFRX1 \i_MIPS/Register/register_reg[20][28]  ( .D(\i_MIPS/Register/n496 ), 
        .CK(clk), .RN(n5777), .Q(\i_MIPS/Register/register[20][28] ), .QN(
        n2475) );
  DFFRX1 \i_MIPS/Register/register_reg[20][29]  ( .D(\i_MIPS/Register/n497 ), 
        .CK(clk), .RN(n5777), .Q(\i_MIPS/Register/register[20][29] ), .QN(
        n2582) );
  DFFRX1 \i_MIPS/Register/register_reg[19][0]  ( .D(\i_MIPS/Register/n500 ), 
        .CK(clk), .RN(n5777), .Q(\i_MIPS/Register/register[19][0] ), .QN(n1039) );
  DFFRX1 \i_MIPS/Register/register_reg[19][1]  ( .D(\i_MIPS/Register/n501 ), 
        .CK(clk), .RN(n5777), .Q(\i_MIPS/Register/register[19][1] ), .QN(n2520) );
  DFFRX1 \i_MIPS/Register/register_reg[19][2]  ( .D(\i_MIPS/Register/n502 ), 
        .CK(clk), .RN(n5777), .Q(\i_MIPS/Register/register[19][2] ), .QN(n2531) );
  DFFRX1 \i_MIPS/Register/register_reg[19][3]  ( .D(\i_MIPS/Register/n503 ), 
        .CK(clk), .RN(n5777), .Q(\i_MIPS/Register/register[19][3] ), .QN(n2586) );
  DFFRX1 \i_MIPS/Register/register_reg[19][4]  ( .D(\i_MIPS/Register/n504 ), 
        .CK(clk), .RN(n5777), .Q(\i_MIPS/Register/register[19][4] ), .QN(n2621) );
  DFFRX1 \i_MIPS/Register/register_reg[19][5]  ( .D(\i_MIPS/Register/n505 ), 
        .CK(clk), .RN(n5776), .Q(\i_MIPS/Register/register[19][5] ), .QN(n2624) );
  DFFRX1 \i_MIPS/Register/register_reg[19][6]  ( .D(\i_MIPS/Register/n506 ), 
        .CK(clk), .RN(n5776), .Q(\i_MIPS/Register/register[19][6] ), .QN(n2466) );
  DFFRX1 \i_MIPS/Register/register_reg[19][7]  ( .D(\i_MIPS/Register/n507 ), 
        .CK(clk), .RN(n5776), .Q(\i_MIPS/Register/register[19][7] ), .QN(n2599) );
  DFFRX1 \i_MIPS/Register/register_reg[19][8]  ( .D(\i_MIPS/Register/n508 ), 
        .CK(clk), .RN(n5781), .Q(\i_MIPS/Register/register[19][8] ), .QN(n2499) );
  DFFRX1 \i_MIPS/Register/register_reg[19][9]  ( .D(\i_MIPS/Register/n509 ), 
        .CK(clk), .RN(n5756), .Q(\i_MIPS/Register/register[19][9] ), .QN(n2503) );
  DFFRX1 \i_MIPS/Register/register_reg[19][10]  ( .D(\i_MIPS/Register/n510 ), 
        .CK(clk), .RN(n5756), .Q(\i_MIPS/Register/register[19][10] ), .QN(
        n1024) );
  DFFRX1 \i_MIPS/Register/register_reg[19][11]  ( .D(\i_MIPS/Register/n511 ), 
        .CK(clk), .RN(n5756), .Q(\i_MIPS/Register/register[19][11] ), .QN(n479) );
  DFFRX1 \i_MIPS/Register/register_reg[19][12]  ( .D(\i_MIPS/Register/n512 ), 
        .CK(clk), .RN(n5756), .Q(\i_MIPS/Register/register[19][12] ), .QN(
        n1073) );
  DFFRX1 \i_MIPS/Register/register_reg[19][13]  ( .D(\i_MIPS/Register/n513 ), 
        .CK(clk), .RN(n5756), .Q(\i_MIPS/Register/register[19][13] ), .QN(
        n2528) );
  DFFRX1 \i_MIPS/Register/register_reg[19][14]  ( .D(\i_MIPS/Register/n514 ), 
        .CK(clk), .RN(n5756), .Q(\i_MIPS/Register/register[19][14] ), .QN(
        n1042) );
  DFFRX1 \i_MIPS/Register/register_reg[19][15]  ( .D(\i_MIPS/Register/n515 ), 
        .CK(clk), .RN(n5756), .Q(\i_MIPS/Register/register[19][15] ), .QN(
        n1037) );
  DFFRX1 \i_MIPS/Register/register_reg[19][16]  ( .D(\i_MIPS/Register/n516 ), 
        .CK(clk), .RN(n5756), .Q(\i_MIPS/Register/register[19][16] ), .QN(
        n2524) );
  DFFRX1 \i_MIPS/Register/register_reg[19][17]  ( .D(\i_MIPS/Register/n517 ), 
        .CK(clk), .RN(n5756), .Q(\i_MIPS/Register/register[19][17] ), .QN(
        n2606) );
  DFFRX1 \i_MIPS/Register/register_reg[19][18]  ( .D(\i_MIPS/Register/n518 ), 
        .CK(clk), .RN(n5755), .Q(\i_MIPS/Register/register[19][18] ), .QN(
        n2550) );
  DFFRX1 \i_MIPS/Register/register_reg[19][20]  ( .D(\i_MIPS/Register/n520 ), 
        .CK(clk), .RN(n5755), .Q(\i_MIPS/Register/register[19][20] ), .QN(
        n2518) );
  DFFRX1 \i_MIPS/Register/register_reg[19][21]  ( .D(\i_MIPS/Register/n521 ), 
        .CK(clk), .RN(n5755), .Q(\i_MIPS/Register/register[19][21] ), .QN(
        n2041) );
  DFFRX1 \i_MIPS/Register/register_reg[19][22]  ( .D(\i_MIPS/Register/n522 ), 
        .CK(clk), .RN(n5755), .Q(\i_MIPS/Register/register[19][22] ), .QN(
        n2602) );
  DFFRX1 \i_MIPS/Register/register_reg[19][23]  ( .D(\i_MIPS/Register/n523 ), 
        .CK(clk), .RN(n5755), .Q(\i_MIPS/Register/register[19][23] ), .QN(
        n2069) );
  DFFRX1 \i_MIPS/Register/register_reg[19][24]  ( .D(\i_MIPS/Register/n524 ), 
        .CK(clk), .RN(n5755), .Q(\i_MIPS/Register/register[19][24] ), .QN(
        n2549) );
  DFFRX1 \i_MIPS/Register/register_reg[19][25]  ( .D(\i_MIPS/Register/n525 ), 
        .CK(clk), .RN(n5755), .Q(\i_MIPS/Register/register[19][25] ), .QN(
        n2509) );
  DFFRX1 \i_MIPS/Register/register_reg[19][26]  ( .D(\i_MIPS/Register/n526 ), 
        .CK(clk), .RN(n5755), .Q(\i_MIPS/Register/register[19][26] ), .QN(
        n2612) );
  DFFRX1 \i_MIPS/Register/register_reg[19][28]  ( .D(\i_MIPS/Register/n528 ), 
        .CK(clk), .RN(n5755), .Q(\i_MIPS/Register/register[19][28] ), .QN(
        n2587) );
  DFFRX1 \i_MIPS/Register/register_reg[19][29]  ( .D(\i_MIPS/Register/n529 ), 
        .CK(clk), .RN(n5755), .Q(\i_MIPS/Register/register[19][29] ), .QN(
        n2609) );
  DFFRX1 \i_MIPS/Register/register_reg[17][0]  ( .D(\i_MIPS/Register/n564 ), 
        .CK(clk), .RN(n5752), .Q(\i_MIPS/Register/register[17][0] ), .QN(n2508) );
  DFFRX1 \i_MIPS/Register/register_reg[17][1]  ( .D(\i_MIPS/Register/n565 ), 
        .CK(clk), .RN(n5752), .Q(\i_MIPS/Register/register[17][1] ), .QN(n2505) );
  DFFRX1 \i_MIPS/Register/register_reg[17][2]  ( .D(\i_MIPS/Register/n566 ), 
        .CK(clk), .RN(n5751), .Q(\i_MIPS/Register/register[17][2] ), .QN(n2481) );
  DFFRX1 \i_MIPS/Register/register_reg[17][3]  ( .D(\i_MIPS/Register/n567 ), 
        .CK(clk), .RN(n5751), .Q(\i_MIPS/Register/register[17][3] ), .QN(n1034) );
  DFFRX1 \i_MIPS/Register/register_reg[17][4]  ( .D(\i_MIPS/Register/n568 ), 
        .CK(clk), .RN(n5751), .Q(\i_MIPS/Register/register[17][4] ), .QN(n2564) );
  DFFRX1 \i_MIPS/Register/register_reg[17][5]  ( .D(\i_MIPS/Register/n569 ), 
        .CK(clk), .RN(n5751), .Q(\i_MIPS/Register/register[17][5] ), .QN(n2632) );
  DFFRX1 \i_MIPS/Register/register_reg[17][6]  ( .D(\i_MIPS/Register/n570 ), 
        .CK(clk), .RN(n5751), .Q(\i_MIPS/Register/register[17][6] ), .QN(n2482) );
  DFFRX1 \i_MIPS/Register/register_reg[17][7]  ( .D(\i_MIPS/Register/n571 ), 
        .CK(clk), .RN(n5751), .Q(\i_MIPS/Register/register[17][7] ), .QN(n2641) );
  DFFRX1 \i_MIPS/Register/register_reg[17][8]  ( .D(\i_MIPS/Register/n572 ), 
        .CK(clk), .RN(n5751), .Q(\i_MIPS/Register/register[17][8] ), .QN(n2630) );
  DFFRX1 \i_MIPS/Register/register_reg[17][9]  ( .D(\i_MIPS/Register/n573 ), 
        .CK(clk), .RN(n5751), .Q(\i_MIPS/Register/register[17][9] ), .QN(n1057) );
  DFFRX1 \i_MIPS/Register/register_reg[17][10]  ( .D(\i_MIPS/Register/n574 ), 
        .CK(clk), .RN(n5751), .Q(\i_MIPS/Register/register[17][10] ), .QN(
        n2439) );
  DFFRX1 \i_MIPS/Register/register_reg[17][11]  ( .D(\i_MIPS/Register/n575 ), 
        .CK(clk), .RN(n5751), .Q(\i_MIPS/Register/register[17][11] ), .QN(
        n2579) );
  DFFRX1 \i_MIPS/Register/register_reg[17][12]  ( .D(\i_MIPS/Register/n576 ), 
        .CK(clk), .RN(n5751), .Q(\i_MIPS/Register/register[17][12] ), .QN(
        n2435) );
  DFFRX1 \i_MIPS/Register/register_reg[17][13]  ( .D(\i_MIPS/Register/n577 ), 
        .CK(clk), .RN(n5750), .Q(\i_MIPS/Register/register[17][13] ), .QN(
        n2479) );
  DFFRX1 \i_MIPS/Register/register_reg[17][14]  ( .D(\i_MIPS/Register/n578 ), 
        .CK(clk), .RN(n5750), .Q(\i_MIPS/Register/register[17][14] ), .QN(
        n2478) );
  DFFRX1 \i_MIPS/Register/register_reg[17][15]  ( .D(\i_MIPS/Register/n579 ), 
        .CK(clk), .RN(n5750), .Q(\i_MIPS/Register/register[17][15] ), .QN(
        n2441) );
  DFFRX1 \i_MIPS/Register/register_reg[17][16]  ( .D(\i_MIPS/Register/n580 ), 
        .CK(clk), .RN(n5750), .Q(\i_MIPS/Register/register[17][16] ), .QN(
        n2422) );
  DFFRX1 \i_MIPS/Register/register_reg[17][17]  ( .D(\i_MIPS/Register/n581 ), 
        .CK(clk), .RN(n5750), .Q(\i_MIPS/Register/register[17][17] ), .QN(
        n2627) );
  DFFRX1 \i_MIPS/Register/register_reg[17][18]  ( .D(\i_MIPS/Register/n582 ), 
        .CK(clk), .RN(n5750), .Q(\i_MIPS/Register/register[17][18] ), .QN(
        n1026) );
  DFFRX1 \i_MIPS/Register/register_reg[17][20]  ( .D(\i_MIPS/Register/n584 ), 
        .CK(clk), .RN(n5750), .Q(\i_MIPS/Register/register[17][20] ), .QN(
        n1029) );
  DFFRX1 \i_MIPS/Register/register_reg[17][21]  ( .D(\i_MIPS/Register/n585 ), 
        .CK(clk), .RN(n5750), .Q(\i_MIPS/Register/register[17][21] ), .QN(n403) );
  DFFRX1 \i_MIPS/Register/register_reg[17][22]  ( .D(\i_MIPS/Register/n586 ), 
        .CK(clk), .RN(n5750), .Q(\i_MIPS/Register/register[17][22] ), .QN(
        n1069) );
  DFFRX1 \i_MIPS/Register/register_reg[17][23]  ( .D(\i_MIPS/Register/n587 ), 
        .CK(clk), .RN(n5750), .Q(\i_MIPS/Register/register[17][23] ), .QN(
        n1023) );
  DFFRX1 \i_MIPS/Register/register_reg[17][24]  ( .D(\i_MIPS/Register/n588 ), 
        .CK(clk), .RN(n5750), .Q(\i_MIPS/Register/register[17][24] ), .QN(
        n1060) );
  DFFRX1 \i_MIPS/Register/register_reg[17][25]  ( .D(\i_MIPS/Register/n589 ), 
        .CK(clk), .RN(n5749), .Q(\i_MIPS/Register/register[17][25] ), .QN(
        n1062) );
  DFFRX1 \i_MIPS/Register/register_reg[17][26]  ( .D(\i_MIPS/Register/n590 ), 
        .CK(clk), .RN(n5749), .Q(\i_MIPS/Register/register[17][26] ), .QN(
        n1071) );
  DFFRX1 \i_MIPS/Register/register_reg[17][28]  ( .D(\i_MIPS/Register/n592 ), 
        .CK(clk), .RN(n5749), .Q(\i_MIPS/Register/register[17][28] ), .QN(
        n1068) );
  DFFRX1 \i_MIPS/Register/register_reg[17][29]  ( .D(\i_MIPS/Register/n593 ), 
        .CK(clk), .RN(n5749), .Q(\i_MIPS/Register/register[17][29] ), .QN(
        n2629) );
  DFFRX1 \i_MIPS/Register/register_reg[16][0]  ( .D(\i_MIPS/Register/n596 ), 
        .CK(clk), .RN(n5749), .Q(\i_MIPS/Register/register[16][0] ), .QN(n2598) );
  DFFRX1 \i_MIPS/Register/register_reg[16][1]  ( .D(\i_MIPS/Register/n597 ), 
        .CK(clk), .RN(n5749), .Q(\i_MIPS/Register/register[16][1] ), .QN(n1041) );
  DFFRX1 \i_MIPS/Register/register_reg[16][2]  ( .D(\i_MIPS/Register/n598 ), 
        .CK(clk), .RN(n5749), .Q(\i_MIPS/Register/register[16][2] ), .QN(n2215) );
  DFFRX1 \i_MIPS/Register/register_reg[16][3]  ( .D(\i_MIPS/Register/n599 ), 
        .CK(clk), .RN(n5749), .Q(\i_MIPS/Register/register[16][3] ), .QN(n2638) );
  DFFRX1 \i_MIPS/Register/register_reg[16][4]  ( .D(\i_MIPS/Register/n600 ), 
        .CK(clk), .RN(n5749), .Q(\i_MIPS/Register/register[16][4] ), .QN(n2052) );
  DFFRX1 \i_MIPS/Register/register_reg[16][5]  ( .D(\i_MIPS/Register/n601 ), 
        .CK(clk), .RN(n5748), .Q(\i_MIPS/Register/register[16][5] ), .QN(n2053) );
  DFFRX1 \i_MIPS/Register/register_reg[16][6]  ( .D(\i_MIPS/Register/n602 ), 
        .CK(clk), .RN(n5748), .Q(\i_MIPS/Register/register[16][6] ), .QN(n2029) );
  DFFRX1 \i_MIPS/Register/register_reg[16][7]  ( .D(\i_MIPS/Register/n603 ), 
        .CK(clk), .RN(n5748), .Q(\i_MIPS/Register/register[16][7] ), .QN(n1066) );
  DFFRX1 \i_MIPS/Register/register_reg[16][8]  ( .D(\i_MIPS/Register/n604 ), 
        .CK(clk), .RN(n5748), .Q(\i_MIPS/Register/register[16][8] ), .QN(n2054) );
  DFFRX1 \i_MIPS/Register/register_reg[16][9]  ( .D(\i_MIPS/Register/n605 ), 
        .CK(clk), .RN(n5748), .Q(\i_MIPS/Register/register[16][9] ), .QN(n2637) );
  DFFRX1 \i_MIPS/Register/register_reg[16][10]  ( .D(\i_MIPS/Register/n606 ), 
        .CK(clk), .RN(n5748), .Q(\i_MIPS/Register/register[16][10] ), .QN(
        n2434) );
  DFFRX1 \i_MIPS/Register/register_reg[16][11]  ( .D(\i_MIPS/Register/n607 ), 
        .CK(clk), .RN(n5748), .Q(\i_MIPS/Register/register[16][11] ), .QN(
        n2594) );
  DFFRX1 \i_MIPS/Register/register_reg[16][12]  ( .D(\i_MIPS/Register/n608 ), 
        .CK(clk), .RN(n5748), .Q(\i_MIPS/Register/register[16][12] ), .QN(
        n2516) );
  DFFRX1 \i_MIPS/Register/register_reg[16][13]  ( .D(\i_MIPS/Register/n609 ), 
        .CK(clk), .RN(n5748), .Q(\i_MIPS/Register/register[16][13] ), .QN(
        n1064) );
  DFFRX1 \i_MIPS/Register/register_reg[16][14]  ( .D(\i_MIPS/Register/n610 ), 
        .CK(clk), .RN(n5748), .Q(\i_MIPS/Register/register[16][14] ), .QN(
        n2592) );
  DFFRX1 \i_MIPS/Register/register_reg[16][15]  ( .D(\i_MIPS/Register/n611 ), 
        .CK(clk), .RN(n5748), .Q(\i_MIPS/Register/register[16][15] ), .QN(
        n2596) );
  DFFRX1 \i_MIPS/Register/register_reg[16][16]  ( .D(\i_MIPS/Register/n612 ), 
        .CK(clk), .RN(n5748), .Q(\i_MIPS/Register/register[16][16] ), .QN(
        n1055) );
  DFFRX1 \i_MIPS/Register/register_reg[16][17]  ( .D(\i_MIPS/Register/n613 ), 
        .CK(clk), .RN(n5747), .Q(\i_MIPS/Register/register[16][17] ), .QN(
        n1067) );
  DFFRX1 \i_MIPS/Register/register_reg[16][18]  ( .D(\i_MIPS/Register/n614 ), 
        .CK(clk), .RN(n5747), .Q(\i_MIPS/Register/register[16][18] ), .QN(
        n2425) );
  DFFRX1 \i_MIPS/Register/register_reg[16][20]  ( .D(\i_MIPS/Register/n616 ), 
        .CK(clk), .RN(n5747), .Q(\i_MIPS/Register/register[16][20] ), .QN(
        n2024) );
  DFFRX1 \i_MIPS/Register/register_reg[16][21]  ( .D(\i_MIPS/Register/n617 ), 
        .CK(clk), .RN(n5747), .Q(\i_MIPS/Register/register[16][21] ), .QN(
        n2048) );
  DFFRX1 \i_MIPS/Register/register_reg[16][23]  ( .D(\i_MIPS/Register/n619 ), 
        .CK(clk), .RN(n5747), .Q(\i_MIPS/Register/register[16][23] ), .QN(
        n2636) );
  DFFRX1 \i_MIPS/Register/register_reg[16][24]  ( .D(\i_MIPS/Register/n620 ), 
        .CK(clk), .RN(n5747), .Q(\i_MIPS/Register/register[16][24] ), .QN(
        n2639) );
  DFFRX1 \i_MIPS/Register/register_reg[16][25]  ( .D(\i_MIPS/Register/n621 ), 
        .CK(clk), .RN(n5747), .Q(\i_MIPS/Register/register[16][25] ), .QN(
        n2050) );
  DFFRX1 \i_MIPS/Register/register_reg[16][26]  ( .D(\i_MIPS/Register/n622 ), 
        .CK(clk), .RN(n5747), .Q(\i_MIPS/Register/register[16][26] ), .QN(
        n2025) );
  DFFRX1 \i_MIPS/Register/register_reg[16][28]  ( .D(\i_MIPS/Register/n624 ), 
        .CK(clk), .RN(n5747), .Q(\i_MIPS/Register/register[16][28] ), .QN(
        n2577) );
  DFFRX1 \i_MIPS/Register/register_reg[16][29]  ( .D(\i_MIPS/Register/n625 ), 
        .CK(clk), .RN(n5746), .Q(\i_MIPS/Register/register[16][29] ), .QN(
        n1049) );
  DFFRX1 \i_MIPS/Register/register_reg[7][0]  ( .D(\i_MIPS/Register/n884 ), 
        .CK(clk), .RN(n5665), .Q(\i_MIPS/Register/register[7][0] ), .QN(n2454)
         );
  DFFRX1 \i_MIPS/Register/register_reg[7][1]  ( .D(\i_MIPS/Register/n885 ), 
        .CK(clk), .RN(n5665), .Q(\i_MIPS/Register/register[7][1] ), .QN(n2525)
         );
  DFFRX1 \i_MIPS/Register/register_reg[7][2]  ( .D(\i_MIPS/Register/n886 ), 
        .CK(clk), .RN(n5665), .Q(\i_MIPS/Register/register[7][2] ), .QN(n2468)
         );
  DFFRX1 \i_MIPS/Register/register_reg[7][3]  ( .D(\i_MIPS/Register/n887 ), 
        .CK(clk), .RN(n5665), .Q(\i_MIPS/Register/register[7][3] ), .QN(n2558)
         );
  DFFRX1 \i_MIPS/Register/register_reg[7][4]  ( .D(\i_MIPS/Register/n888 ), 
        .CK(clk), .RN(n5665), .Q(\i_MIPS/Register/register[7][4] ), .QN(n2562)
         );
  DFFRX1 \i_MIPS/Register/register_reg[7][5]  ( .D(\i_MIPS/Register/n889 ), 
        .CK(clk), .RN(n5665), .Q(\i_MIPS/Register/register[7][5] ), .QN(n2563)
         );
  DFFRX1 \i_MIPS/Register/register_reg[7][6]  ( .D(\i_MIPS/Register/n890 ), 
        .CK(clk), .RN(n5665), .Q(\i_MIPS/Register/register[7][6] ), .QN(n2470)
         );
  DFFRX1 \i_MIPS/Register/register_reg[7][7]  ( .D(\i_MIPS/Register/n891 ), 
        .CK(clk), .RN(n5665), .Q(\i_MIPS/Register/register[7][7] ), .QN(n2498)
         );
  DFFRX1 \i_MIPS/Register/register_reg[7][8]  ( .D(\i_MIPS/Register/n892 ), 
        .CK(clk), .RN(n5664), .Q(\i_MIPS/Register/register[7][8] ), .QN(n2619)
         );
  DFFRX1 \i_MIPS/Register/register_reg[7][9]  ( .D(\i_MIPS/Register/n893 ), 
        .CK(clk), .RN(n5664), .Q(\i_MIPS/Register/register[7][9] ), .QN(n2556)
         );
  DFFRX1 \i_MIPS/Register/register_reg[7][10]  ( .D(\i_MIPS/Register/n894 ), 
        .CK(clk), .RN(n5664), .Q(\i_MIPS/Register/register[7][10] ), .QN(n2453) );
  DFFRX1 \i_MIPS/Register/register_reg[7][11]  ( .D(\i_MIPS/Register/n895 ), 
        .CK(clk), .RN(n5664), .Q(\i_MIPS/Register/register[7][11] ), .QN(n2451) );
  DFFRX1 \i_MIPS/Register/register_reg[7][12]  ( .D(\i_MIPS/Register/n896 ), 
        .CK(clk), .RN(n5664), .Q(\i_MIPS/Register/register[7][12] ), .QN(n2511) );
  DFFRX1 \i_MIPS/Register/register_reg[7][13]  ( .D(\i_MIPS/Register/n897 ), 
        .CK(clk), .RN(n5664), .Q(\i_MIPS/Register/register[7][13] ), .QN(n2464) );
  DFFRX1 \i_MIPS/Register/register_reg[7][14]  ( .D(\i_MIPS/Register/n898 ), 
        .CK(clk), .RN(n5664), .Q(\i_MIPS/Register/register[7][14] ), .QN(n2461) );
  DFFRX1 \i_MIPS/Register/register_reg[7][15]  ( .D(\i_MIPS/Register/n899 ), 
        .CK(clk), .RN(n5664), .Q(\i_MIPS/Register/register[7][15] ), .QN(n2514) );
  DFFRX1 \i_MIPS/Register/register_reg[7][16]  ( .D(\i_MIPS/Register/n900 ), 
        .CK(clk), .RN(n5664), .Q(\i_MIPS/Register/register[7][16] ), .QN(n2529) );
  DFFRX1 \i_MIPS/Register/register_reg[7][17]  ( .D(\i_MIPS/Register/n901 ), 
        .CK(clk), .RN(n5664), .Q(\i_MIPS/Register/register[7][17] ), .QN(n2608) );
  DFFRX1 \i_MIPS/Register/register_reg[7][18]  ( .D(\i_MIPS/Register/n902 ), 
        .CK(clk), .RN(n5664), .Q(\i_MIPS/Register/register[7][18] ), .QN(n2555) );
  DFFRX1 \i_MIPS/Register/register_reg[7][20]  ( .D(\i_MIPS/Register/n904 ), 
        .CK(clk), .RN(n5663), .Q(\i_MIPS/Register/register[7][20] ), .QN(n2459) );
  DFFRX1 \i_MIPS/Register/register_reg[7][21]  ( .D(\i_MIPS/Register/n905 ), 
        .CK(clk), .RN(n5663), .Q(\i_MIPS/Register/register[7][21] ), .QN(n2444) );
  DFFRX1 \i_MIPS/Register/register_reg[7][22]  ( .D(\i_MIPS/Register/n906 ), 
        .CK(clk), .RN(n5663), .Q(\i_MIPS/Register/register[7][22] ), .QN(n2605) );
  DFFRX1 \i_MIPS/Register/register_reg[7][23]  ( .D(\i_MIPS/Register/n907 ), 
        .CK(clk), .RN(n5663), .Q(\i_MIPS/Register/register[7][23] ), .QN(n2557) );
  DFFRX1 \i_MIPS/Register/register_reg[7][24]  ( .D(\i_MIPS/Register/n908 ), 
        .CK(clk), .RN(n5663), .Q(\i_MIPS/Register/register[7][24] ), .QN(n2561) );
  DFFRX1 \i_MIPS/Register/register_reg[7][25]  ( .D(\i_MIPS/Register/n909 ), 
        .CK(clk), .RN(n5663), .Q(\i_MIPS/Register/register[7][25] ) );
  DFFRX1 \i_MIPS/Register/register_reg[7][26]  ( .D(\i_MIPS/Register/n910 ), 
        .CK(clk), .RN(n5663), .Q(\i_MIPS/Register/register[7][26] ), .QN(n2615) );
  DFFRX1 \i_MIPS/Register/register_reg[7][28]  ( .D(\i_MIPS/Register/n912 ), 
        .CK(clk), .RN(n5663), .Q(\i_MIPS/Register/register[7][28] ), .QN(n2559) );
  DFFRX1 \i_MIPS/Register/register_reg[7][29]  ( .D(\i_MIPS/Register/n913 ), 
        .CK(clk), .RN(n5663), .Q(\i_MIPS/Register/register[7][29] ), .QN(n2611) );
  DFFRX1 \i_MIPS/Register/register_reg[5][0]  ( .D(\i_MIPS/Register/n948 ), 
        .CK(clk), .RN(n5660), .Q(\i_MIPS/Register/register[5][0] ), .QN(n2447)
         );
  DFFRX1 \i_MIPS/Register/register_reg[5][1]  ( .D(\i_MIPS/Register/n949 ), 
        .CK(clk), .RN(n5660), .Q(\i_MIPS/Register/register[5][1] ), .QN(n2527)
         );
  DFFRX1 \i_MIPS/Register/register_reg[5][2]  ( .D(\i_MIPS/Register/n950 ), 
        .CK(clk), .RN(n5660), .Q(\i_MIPS/Register/register[5][2] ), .QN(n2469)
         );
  DFFRX1 \i_MIPS/Register/register_reg[5][3]  ( .D(\i_MIPS/Register/n951 ), 
        .CK(clk), .RN(n5659), .Q(\i_MIPS/Register/register[5][3] ), .QN(n2038)
         );
  DFFRX1 \i_MIPS/Register/register_reg[5][4]  ( .D(\i_MIPS/Register/n952 ), 
        .CK(clk), .RN(n5659), .Q(\i_MIPS/Register/register[5][4] ), .QN(n2553)
         );
  DFFRX1 \i_MIPS/Register/register_reg[5][5]  ( .D(\i_MIPS/Register/n953 ), 
        .CK(clk), .RN(n5659), .Q(\i_MIPS/Register/register[5][5] ), .QN(n2554)
         );
  DFFRX1 \i_MIPS/Register/register_reg[5][6]  ( .D(\i_MIPS/Register/n954 ), 
        .CK(clk), .RN(n5659), .Q(\i_MIPS/Register/register[5][6] ), .QN(n2472)
         );
  DFFRX1 \i_MIPS/Register/register_reg[5][7]  ( .D(\i_MIPS/Register/n955 ), 
        .CK(clk), .RN(n5659), .Q(\i_MIPS/Register/register[5][7] ), .QN(n2042)
         );
  DFFRX1 \i_MIPS/Register/register_reg[5][8]  ( .D(\i_MIPS/Register/n956 ), 
        .CK(clk), .RN(n5659), .Q(\i_MIPS/Register/register[5][8] ), .QN(n2551)
         );
  DFFRX1 \i_MIPS/Register/register_reg[5][9]  ( .D(\i_MIPS/Register/n957 ), 
        .CK(clk), .RN(n5659), .Q(\i_MIPS/Register/register[5][9] ), .QN(n2213)
         );
  DFFRX1 \i_MIPS/Register/register_reg[5][10]  ( .D(\i_MIPS/Register/n958 ), 
        .CK(clk), .RN(n5659), .Q(\i_MIPS/Register/register[5][10] ), .QN(n2034) );
  DFFRX1 \i_MIPS/Register/register_reg[5][11]  ( .D(\i_MIPS/Register/n959 ), 
        .CK(clk), .RN(n5659), .Q(\i_MIPS/Register/register[5][11] ), .QN(n2571) );
  DFFRX1 \i_MIPS/Register/register_reg[5][12]  ( .D(\i_MIPS/Register/n960 ), 
        .CK(clk), .RN(n5659), .Q(\i_MIPS/Register/register[5][12] ), .QN(n2062) );
  DFFRX1 \i_MIPS/Register/register_reg[5][13]  ( .D(\i_MIPS/Register/n961 ), 
        .CK(clk), .RN(n5659), .Q(\i_MIPS/Register/register[5][13] ), .QN(n2023) );
  DFFRX1 \i_MIPS/Register/register_reg[5][14]  ( .D(\i_MIPS/Register/n962 ), 
        .CK(clk), .RN(n5659), .Q(\i_MIPS/Register/register[5][14] ), .QN(n2033) );
  DFFRX1 \i_MIPS/Register/register_reg[5][15]  ( .D(\i_MIPS/Register/n963 ), 
        .CK(clk), .RN(n5658), .Q(\i_MIPS/Register/register[5][15] ), .QN(n2063) );
  DFFRX1 \i_MIPS/Register/register_reg[5][16]  ( .D(\i_MIPS/Register/n964 ), 
        .CK(clk), .RN(n5658), .Q(\i_MIPS/Register/register[5][16] ), .QN(n2045) );
  DFFRX1 \i_MIPS/Register/register_reg[5][17]  ( .D(\i_MIPS/Register/n965 ), 
        .CK(clk), .RN(n5658), .Q(\i_MIPS/Register/register[5][17] ), .QN(n2043) );
  DFFRX1 \i_MIPS/Register/register_reg[5][18]  ( .D(\i_MIPS/Register/n966 ), 
        .CK(clk), .RN(n5658), .Q(\i_MIPS/Register/register[5][18] ), .QN(n2037) );
  DFFRX1 \i_MIPS/Register/register_reg[5][20]  ( .D(\i_MIPS/Register/n968 ), 
        .CK(clk), .RN(n5658), .Q(\i_MIPS/Register/register[5][20] ), .QN(n2056) );
  DFFRX1 \i_MIPS/Register/register_reg[5][21]  ( .D(\i_MIPS/Register/n969 ), 
        .CK(clk), .RN(n5658), .Q(\i_MIPS/Register/register[5][21] ), .QN(n2507) );
  DFFRX1 \i_MIPS/Register/register_reg[5][22]  ( .D(\i_MIPS/Register/n970 ), 
        .CK(clk), .RN(n5658), .Q(\i_MIPS/Register/register[5][22] ), .QN(n2496) );
  DFFRX1 \i_MIPS/Register/register_reg[5][23]  ( .D(\i_MIPS/Register/n971 ), 
        .CK(clk), .RN(n5658), .Q(\i_MIPS/Register/register[5][23] ), .QN(n2573) );
  DFFRX1 \i_MIPS/Register/register_reg[5][24]  ( .D(\i_MIPS/Register/n972 ), 
        .CK(clk), .RN(n5658), .Q(\i_MIPS/Register/register[5][24] ), .QN(n2039) );
  DFFRX1 \i_MIPS/Register/register_reg[5][25]  ( .D(\i_MIPS/Register/n973 ), 
        .CK(clk), .RN(n5658), .Q(\i_MIPS/Register/register[5][25] ), .QN(n2031) );
  DFFRX1 \i_MIPS/Register/register_reg[5][26]  ( .D(\i_MIPS/Register/n974 ), 
        .CK(clk), .RN(n5658), .Q(\i_MIPS/Register/register[5][26] ), .QN(n2058) );
  DFFRX1 \i_MIPS/Register/register_reg[5][28]  ( .D(\i_MIPS/Register/n976 ), 
        .CK(clk), .RN(n5657), .Q(\i_MIPS/Register/register[5][28] ), .QN(n2035) );
  DFFRX1 \i_MIPS/Register/register_reg[5][29]  ( .D(\i_MIPS/Register/n977 ), 
        .CK(clk), .RN(n5657), .Q(\i_MIPS/Register/register[5][29] ), .QN(n2068) );
  DFFRX1 \i_MIPS/Register/register_reg[4][0]  ( .D(\i_MIPS/Register/n980 ), 
        .CK(clk), .RN(n5657), .Q(\i_MIPS/Register/register[4][0] ), .QN(n979)
         );
  DFFRX1 \i_MIPS/Register/register_reg[4][1]  ( .D(\i_MIPS/Register/n981 ), 
        .CK(clk), .RN(n5657), .Q(\i_MIPS/Register/register[4][1] ), .QN(n2487)
         );
  DFFRX1 \i_MIPS/Register/register_reg[4][2]  ( .D(\i_MIPS/Register/n982 ), 
        .CK(clk), .RN(n5657), .Q(\i_MIPS/Register/register[4][2] ), .QN(n2448)
         );
  DFFRX1 \i_MIPS/Register/register_reg[4][3]  ( .D(\i_MIPS/Register/n983 ), 
        .CK(clk), .RN(n5657), .Q(\i_MIPS/Register/register[4][3] ), .QN(n2493)
         );
  DFFRX1 \i_MIPS/Register/register_reg[4][4]  ( .D(\i_MIPS/Register/n984 ), 
        .CK(clk), .RN(n5657), .Q(\i_MIPS/Register/register[4][4] ), .QN(n2433)
         );
  DFFRX1 \i_MIPS/Register/register_reg[4][5]  ( .D(\i_MIPS/Register/n985 ), 
        .CK(clk), .RN(n5657), .Q(\i_MIPS/Register/register[4][5] ), .QN(n2486)
         );
  DFFRX1 \i_MIPS/Register/register_reg[4][6]  ( .D(\i_MIPS/Register/n986 ), 
        .CK(clk), .RN(n5657), .Q(\i_MIPS/Register/register[4][6] ), .QN(n2490)
         );
  DFFRX1 \i_MIPS/Register/register_reg[4][7]  ( .D(\i_MIPS/Register/n987 ), 
        .CK(clk), .RN(n5661), .Q(\i_MIPS/Register/register[4][7] ), .QN(n2431)
         );
  DFFRX1 \i_MIPS/Register/register_reg[4][8]  ( .D(\i_MIPS/Register/n988 ), 
        .CK(clk), .RN(n5636), .Q(\i_MIPS/Register/register[4][8] ), .QN(n2547)
         );
  DFFRX1 \i_MIPS/Register/register_reg[4][9]  ( .D(\i_MIPS/Register/n989 ), 
        .CK(clk), .RN(n5636), .Q(\i_MIPS/Register/register[4][9] ), .QN(n2430)
         );
  DFFRX1 \i_MIPS/Register/register_reg[4][10]  ( .D(\i_MIPS/Register/n990 ), 
        .CK(clk), .RN(n5636), .Q(\i_MIPS/Register/register[4][10] ), .QN(n978)
         );
  DFFRX1 \i_MIPS/Register/register_reg[4][11]  ( .D(\i_MIPS/Register/n991 ), 
        .CK(clk), .RN(n5636), .Q(\i_MIPS/Register/register[4][11] ), .QN(n980)
         );
  DFFRX1 \i_MIPS/Register/register_reg[4][12]  ( .D(\i_MIPS/Register/n992 ), 
        .CK(clk), .RN(n5636), .Q(\i_MIPS/Register/register[4][12] ), .QN(n1032) );
  DFFRX1 \i_MIPS/Register/register_reg[4][13]  ( .D(\i_MIPS/Register/n993 ), 
        .CK(clk), .RN(n5636), .Q(\i_MIPS/Register/register[4][13] ), .QN(n2488) );
  DFFRX1 \i_MIPS/Register/register_reg[4][14]  ( .D(\i_MIPS/Register/n994 ), 
        .CK(clk), .RN(n5636), .Q(\i_MIPS/Register/register[4][14] ), .QN(n1033) );
  DFFRX1 \i_MIPS/Register/register_reg[4][15]  ( .D(\i_MIPS/Register/n995 ), 
        .CK(clk), .RN(n5636), .Q(\i_MIPS/Register/register[4][15] ), .QN(n1050) );
  DFFRX1 \i_MIPS/Register/register_reg[4][16]  ( .D(\i_MIPS/Register/n996 ), 
        .CK(clk), .RN(n5636), .Q(\i_MIPS/Register/register[4][16] ), .QN(n2491) );
  DFFRX1 \i_MIPS/Register/register_reg[4][17]  ( .D(\i_MIPS/Register/n997 ), 
        .CK(clk), .RN(n5636), .Q(\i_MIPS/Register/register[4][17] ), .QN(n2427) );
  DFFRX1 \i_MIPS/Register/register_reg[4][18]  ( .D(\i_MIPS/Register/n998 ), 
        .CK(clk), .RN(n5636), .Q(\i_MIPS/Register/register[4][18] ), .QN(n2428) );
  DFFRX1 \i_MIPS/Register/register_reg[4][20]  ( .D(\i_MIPS/Register/n1000 ), 
        .CK(clk), .RN(n5635), .Q(\i_MIPS/Register/register[4][20] ), .QN(n2489) );
  DFFRX1 \i_MIPS/Register/register_reg[4][21]  ( .D(\i_MIPS/Register/n1001 ), 
        .CK(clk), .RN(n5635), .Q(\i_MIPS/Register/register[4][21] ), .QN(n2546) );
  DFFRX1 \i_MIPS/Register/register_reg[4][23]  ( .D(\i_MIPS/Register/n1003 ), 
        .CK(clk), .RN(n5635), .Q(\i_MIPS/Register/register[4][23] ), .QN(n2429) );
  DFFRX1 \i_MIPS/Register/register_reg[4][24]  ( .D(\i_MIPS/Register/n1004 ), 
        .CK(clk), .RN(n5635), .Q(\i_MIPS/Register/register[4][24] ), .QN(n2495) );
  DFFRX1 \i_MIPS/Register/register_reg[4][25]  ( .D(\i_MIPS/Register/n1005 ), 
        .CK(clk), .RN(n5635), .Q(\i_MIPS/Register/register[4][25] ), .QN(n2432) );
  DFFRX1 \i_MIPS/Register/register_reg[4][26]  ( .D(\i_MIPS/Register/n1006 ), 
        .CK(clk), .RN(n5635), .Q(\i_MIPS/Register/register[4][26] ), .QN(n2494) );
  DFFRX1 \i_MIPS/Register/register_reg[4][28]  ( .D(\i_MIPS/Register/n1008 ), 
        .CK(clk), .RN(n5635), .Q(\i_MIPS/Register/register[4][28] ), .QN(n2492) );
  DFFRX1 \i_MIPS/Register/register_reg[4][29]  ( .D(\i_MIPS/Register/n1009 ), 
        .CK(clk), .RN(n5635), .Q(\i_MIPS/Register/register[4][29] ), .QN(n2548) );
  DFFRX1 \i_MIPS/Register/register_reg[3][0]  ( .D(\i_MIPS/Register/n1012 ), 
        .CK(clk), .RN(n5634), .Q(\i_MIPS/Register/register[3][0] ), .QN(n1040)
         );
  DFFRX1 \i_MIPS/Register/register_reg[3][1]  ( .D(\i_MIPS/Register/n1013 ), 
        .CK(clk), .RN(n5634), .Q(\i_MIPS/Register/register[3][1] ), .QN(n2526)
         );
  DFFRX1 \i_MIPS/Register/register_reg[3][2]  ( .D(\i_MIPS/Register/n1014 ), 
        .CK(clk), .RN(n5634), .Q(\i_MIPS/Register/register[3][2] ), .QN(n2533)
         );
  DFFRX1 \i_MIPS/Register/register_reg[3][3]  ( .D(\i_MIPS/Register/n1015 ), 
        .CK(clk), .RN(n5634), .Q(\i_MIPS/Register/register[3][3] ), .QN(n2588)
         );
  DFFRX1 \i_MIPS/Register/register_reg[3][4]  ( .D(\i_MIPS/Register/n1016 ), 
        .CK(clk), .RN(n5634), .Q(\i_MIPS/Register/register[3][4] ), .QN(n2623)
         );
  DFFRX1 \i_MIPS/Register/register_reg[3][5]  ( .D(\i_MIPS/Register/n1017 ), 
        .CK(clk), .RN(n5634), .Q(\i_MIPS/Register/register[3][5] ), .QN(n2626)
         );
  DFFRX1 \i_MIPS/Register/register_reg[3][6]  ( .D(\i_MIPS/Register/n1018 ), 
        .CK(clk), .RN(n5634), .Q(\i_MIPS/Register/register[3][6] ), .QN(n2471)
         );
  DFFRX1 \i_MIPS/Register/register_reg[3][7]  ( .D(\i_MIPS/Register/n1019 ), 
        .CK(clk), .RN(n5634), .Q(\i_MIPS/Register/register[3][7] ), .QN(n2600)
         );
  DFFRX1 \i_MIPS/Register/register_reg[3][8]  ( .D(\i_MIPS/Register/n1020 ), 
        .CK(clk), .RN(n5634), .Q(\i_MIPS/Register/register[3][8] ), .QN(n2618)
         );
  DFFRX1 \i_MIPS/Register/register_reg[3][9]  ( .D(\i_MIPS/Register/n1021 ), 
        .CK(clk), .RN(n5634), .Q(\i_MIPS/Register/register[3][9] ), .QN(n2589)
         );
  DFFRX1 \i_MIPS/Register/register_reg[3][10]  ( .D(\i_MIPS/Register/n1022 ), 
        .CK(clk), .RN(n5634), .Q(\i_MIPS/Register/register[3][10] ), .QN(n1025) );
  DFFRX1 \i_MIPS/Register/register_reg[3][11]  ( .D(\i_MIPS/Register/n1023 ), 
        .CK(clk), .RN(n5634), .Q(\i_MIPS/Register/register[3][11] ), .QN(n1036) );
  DFFRX1 \i_MIPS/Register/register_reg[3][12]  ( .D(\i_MIPS/Register/n1024 ), 
        .CK(clk), .RN(n5633), .Q(\i_MIPS/Register/register[3][12] ), .QN(n1035) );
  DFFRX1 \i_MIPS/Register/register_reg[3][13]  ( .D(\i_MIPS/Register/n1025 ), 
        .CK(clk), .RN(n5633), .Q(\i_MIPS/Register/register[3][13] ), .QN(n2532) );
  DFFRX1 \i_MIPS/Register/register_reg[3][14]  ( .D(\i_MIPS/Register/n1026 ), 
        .CK(clk), .RN(n5633), .Q(\i_MIPS/Register/register[3][14] ), .QN(n478)
         );
  DFFRX1 \i_MIPS/Register/register_reg[3][15]  ( .D(\i_MIPS/Register/n1027 ), 
        .CK(clk), .RN(n5633), .Q(\i_MIPS/Register/register[3][15] ), .QN(n1038) );
  DFFRX1 \i_MIPS/Register/register_reg[3][16]  ( .D(\i_MIPS/Register/n1028 ), 
        .CK(clk), .RN(n5633), .Q(\i_MIPS/Register/register[3][16] ), .QN(n2530) );
  DFFRX1 \i_MIPS/Register/register_reg[3][17]  ( .D(\i_MIPS/Register/n1029 ), 
        .CK(clk), .RN(n5633), .Q(\i_MIPS/Register/register[3][17] ), .QN(n2607) );
  DFFRX1 \i_MIPS/Register/register_reg[3][18]  ( .D(\i_MIPS/Register/n1030 ), 
        .CK(clk), .RN(n5633), .Q(\i_MIPS/Register/register[3][18] ), .QN(n2446) );
  DFFRX1 \i_MIPS/Register/register_reg[3][20]  ( .D(\i_MIPS/Register/n1032 ), 
        .CK(clk), .RN(n5633), .Q(\i_MIPS/Register/register[3][20] ), .QN(n2522) );
  DFFRX1 \i_MIPS/Register/register_reg[3][21]  ( .D(\i_MIPS/Register/n1033 ), 
        .CK(clk), .RN(n5633), .Q(\i_MIPS/Register/register[3][21] ), .QN(n2220) );
  DFFRX1 \i_MIPS/Register/register_reg[3][22]  ( .D(\i_MIPS/Register/n1034 ), 
        .CK(clk), .RN(n5633), .Q(\i_MIPS/Register/register[3][22] ), .QN(n2604) );
  DFFRX1 \i_MIPS/Register/register_reg[3][23]  ( .D(\i_MIPS/Register/n1035 ), 
        .CK(clk), .RN(n5633), .Q(\i_MIPS/Register/register[3][23] ), .QN(n2219) );
  DFFRX1 \i_MIPS/Register/register_reg[3][24]  ( .D(\i_MIPS/Register/n1036 ), 
        .CK(clk), .RN(n5632), .Q(\i_MIPS/Register/register[3][24] ), .QN(n2445) );
  DFFRX1 \i_MIPS/Register/register_reg[3][25]  ( .D(\i_MIPS/Register/n1037 ), 
        .CK(clk), .RN(n5632), .Q(\i_MIPS/Register/register[3][25] ), .QN(n2510) );
  DFFRX1 \i_MIPS/Register/register_reg[3][26]  ( .D(\i_MIPS/Register/n1038 ), 
        .CK(clk), .RN(n5632), .Q(\i_MIPS/Register/register[3][26] ), .QN(n2614) );
  DFFRX1 \i_MIPS/Register/register_reg[3][28]  ( .D(\i_MIPS/Register/n1040 ), 
        .CK(clk), .RN(n5632), .Q(\i_MIPS/Register/register[3][28] ), .QN(n2504) );
  DFFRX1 \i_MIPS/Register/register_reg[3][29]  ( .D(\i_MIPS/Register/n1041 ), 
        .CK(clk), .RN(n5632), .Q(\i_MIPS/Register/register[3][29] ), .QN(n2610) );
  DFFRX1 \i_MIPS/Register/register_reg[1][0]  ( .D(\i_MIPS/Register/n1076 ), 
        .CK(clk), .RN(n5629), .Q(\i_MIPS/Register/register[1][0] ), .QN(n2581)
         );
  DFFRX1 \i_MIPS/Register/register_reg[1][1]  ( .D(\i_MIPS/Register/n1077 ), 
        .CK(clk), .RN(n5629), .Q(\i_MIPS/Register/register[1][1] ), .QN(n2634)
         );
  DFFRX1 \i_MIPS/Register/register_reg[1][2]  ( .D(\i_MIPS/Register/n1078 ), 
        .CK(clk), .RN(n5629), .Q(\i_MIPS/Register/register[1][2] ), .QN(n2483)
         );
  DFFRX1 \i_MIPS/Register/register_reg[1][3]  ( .D(\i_MIPS/Register/n1079 ), 
        .CK(clk), .RN(n5629), .Q(\i_MIPS/Register/register[1][3] ), .QN(n1022)
         );
  DFFRX1 \i_MIPS/Register/register_reg[1][4]  ( .D(\i_MIPS/Register/n1080 ), 
        .CK(clk), .RN(n5629), .Q(\i_MIPS/Register/register[1][4] ), .QN(n2565)
         );
  DFFRX1 \i_MIPS/Register/register_reg[1][5]  ( .D(\i_MIPS/Register/n1081 ), 
        .CK(clk), .RN(n5629), .Q(\i_MIPS/Register/register[1][5] ), .QN(n2566)
         );
  DFFRX1 \i_MIPS/Register/register_reg[1][6]  ( .D(\i_MIPS/Register/n1082 ), 
        .CK(clk), .RN(n5629), .Q(\i_MIPS/Register/register[1][6] ), .QN(n2484)
         );
  DFFRX1 \i_MIPS/Register/register_reg[1][7]  ( .D(\i_MIPS/Register/n1083 ), 
        .CK(clk), .RN(n5628), .Q(\i_MIPS/Register/register[1][7] ), .QN(n2642)
         );
  DFFRX1 \i_MIPS/Register/register_reg[1][8]  ( .D(\i_MIPS/Register/n1084 ), 
        .CK(clk), .RN(n5628), .Q(\i_MIPS/Register/register[1][8] ), .QN(n2631)
         );
  DFFRX1 \i_MIPS/Register/register_reg[1][9]  ( .D(\i_MIPS/Register/n1085 ), 
        .CK(clk), .RN(n5628), .Q(\i_MIPS/Register/register[1][9] ), .QN(n1058)
         );
  DFFRX1 \i_MIPS/Register/register_reg[1][10]  ( .D(\i_MIPS/Register/n1086 ), 
        .CK(clk), .RN(n5628), .Q(\i_MIPS/Register/register[1][10] ), .QN(n2440) );
  DFFRX1 \i_MIPS/Register/register_reg[1][11]  ( .D(\i_MIPS/Register/n1087 ), 
        .CK(clk), .RN(n5628), .Q(\i_MIPS/Register/register[1][11] ), .QN(n2580) );
  DFFRX1 \i_MIPS/Register/register_reg[1][12]  ( .D(\i_MIPS/Register/n1088 ), 
        .CK(clk), .RN(n5628), .Q(\i_MIPS/Register/register[1][12] ), .QN(n2438) );
  DFFRX1 \i_MIPS/Register/register_reg[1][13]  ( .D(\i_MIPS/Register/n1089 ), 
        .CK(clk), .RN(n5628), .Q(\i_MIPS/Register/register[1][13] ), .QN(n2437) );
  DFFRX1 \i_MIPS/Register/register_reg[1][14]  ( .D(\i_MIPS/Register/n1090 ), 
        .CK(clk), .RN(n5628), .Q(\i_MIPS/Register/register[1][14] ), .QN(n2480) );
  DFFRX1 \i_MIPS/Register/register_reg[1][15]  ( .D(\i_MIPS/Register/n1091 ), 
        .CK(clk), .RN(n5628), .Q(\i_MIPS/Register/register[1][15] ), .QN(n2643) );
  DFFRX1 \i_MIPS/Register/register_reg[1][16]  ( .D(\i_MIPS/Register/n1092 ), 
        .CK(clk), .RN(n5628), .Q(\i_MIPS/Register/register[1][16] ), .QN(n2423) );
  DFFRX1 \i_MIPS/Register/register_reg[1][17]  ( .D(\i_MIPS/Register/n1093 ), 
        .CK(clk), .RN(n5628), .Q(\i_MIPS/Register/register[1][17] ), .QN(n2628) );
  DFFRX1 \i_MIPS/Register/register_reg[1][18]  ( .D(\i_MIPS/Register/n1094 ), 
        .CK(clk), .RN(n5628), .Q(\i_MIPS/Register/register[1][18] ), .QN(n1027) );
  DFFRX1 \i_MIPS/Register/register_reg[1][20]  ( .D(\i_MIPS/Register/n1096 ), 
        .CK(clk), .RN(n5627), .Q(\i_MIPS/Register/register[1][20] ), .QN(n1030) );
  DFFRX1 \i_MIPS/Register/register_reg[1][21]  ( .D(\i_MIPS/Register/n1097 ), 
        .CK(clk), .RN(n5627), .Q(\i_MIPS/Register/register[1][21] ), .QN(n1028) );
  DFFRX1 \i_MIPS/Register/register_reg[1][22]  ( .D(\i_MIPS/Register/n1098 ), 
        .CK(clk), .RN(n5627), .Q(\i_MIPS/Register/register[1][22] ), .QN(n1070) );
  DFFRX1 \i_MIPS/Register/register_reg[1][23]  ( .D(\i_MIPS/Register/n1099 ), 
        .CK(clk), .RN(n5627), .Q(\i_MIPS/Register/register[1][23] ), .QN(n404)
         );
  DFFRX1 \i_MIPS/Register/register_reg[1][24]  ( .D(\i_MIPS/Register/n1100 ), 
        .CK(clk), .RN(n5627), .Q(\i_MIPS/Register/register[1][24] ), .QN(n1061) );
  DFFRX1 \i_MIPS/Register/register_reg[1][25]  ( .D(\i_MIPS/Register/n1101 ), 
        .CK(clk), .RN(n5627), .Q(\i_MIPS/Register/register[1][25] ), .QN(n1063) );
  DFFRX1 \i_MIPS/Register/register_reg[1][26]  ( .D(\i_MIPS/Register/n1102 ), 
        .CK(clk), .RN(n5627), .Q(\i_MIPS/Register/register[1][26] ), .QN(n1072) );
  DFFRX1 \i_MIPS/Register/register_reg[1][28]  ( .D(\i_MIPS/Register/n1104 ), 
        .CK(clk), .RN(n5627), .Q(\i_MIPS/Register/register[1][28] ), .QN(n1059) );
  DFFRX1 \i_MIPS/Register/register_reg[1][29]  ( .D(\i_MIPS/Register/n1105 ), 
        .CK(clk), .RN(n5627), .Q(\i_MIPS/Register/register[1][29] ), .QN(n2501) );
  DFFRX1 \i_MIPS/Register/register_reg[0][0]  ( .D(\i_MIPS/Register/n1108 ), 
        .CK(clk), .RN(n5646), .Q(\i_MIPS/Register/register[0][0] ), .QN(n2597)
         );
  DFFRX1 \i_MIPS/Register/register_reg[0][1]  ( .D(\i_MIPS/Register/n1109 ), 
        .CK(clk), .RN(n5646), .Q(\i_MIPS/Register/register[0][1] ), .QN(n1053)
         );
  DFFRX1 \i_MIPS/Register/register_reg[0][2]  ( .D(\i_MIPS/Register/n1110 ), 
        .CK(clk), .RN(n5646), .Q(\i_MIPS/Register/register[0][2] ), .QN(n2026)
         );
  DFFRX1 \i_MIPS/Register/register_reg[0][3]  ( .D(\i_MIPS/Register/n1111 ), 
        .CK(clk), .RN(n5646), .Q(\i_MIPS/Register/register[0][3] ), .QN(n2576)
         );
  DFFRX1 \i_MIPS/Register/register_reg[0][4]  ( .D(\i_MIPS/Register/n1112 ), 
        .CK(clk), .RN(n5646), .Q(\i_MIPS/Register/register[0][4] ), .QN(n2051)
         );
  DFFRX1 \i_MIPS/Register/register_reg[0][5]  ( .D(\i_MIPS/Register/n1113 ), 
        .CK(clk), .RN(n5646), .Q(\i_MIPS/Register/register[0][5] ), .QN(n2028)
         );
  DFFRX1 \i_MIPS/Register/register_reg[0][6]  ( .D(\i_MIPS/Register/n1114 ), 
        .CK(clk), .RN(n5646), .Q(\i_MIPS/Register/register[0][6] ), .QN(n2027)
         );
  DFFRX1 \i_MIPS/Register/register_reg[0][7]  ( .D(\i_MIPS/Register/n1115 ), 
        .CK(clk), .RN(n5646), .Q(\i_MIPS/Register/register[0][7] ), .QN(n1065)
         );
  DFFRX1 \i_MIPS/Register/register_reg[0][8]  ( .D(\i_MIPS/Register/n1116 ), 
        .CK(clk), .RN(n5646), .Q(\i_MIPS/Register/register[0][8] ), .QN(n2640)
         );
  DFFRX1 \i_MIPS/Register/register_reg[0][9]  ( .D(\i_MIPS/Register/n1117 ), 
        .CK(clk), .RN(n5646), .Q(\i_MIPS/Register/register[0][9] ), .QN(n2575)
         );
  DFFRX1 \i_MIPS/Register/register_reg[0][10]  ( .D(\i_MIPS/Register/n1118 ), 
        .CK(clk), .RN(n5645), .Q(\i_MIPS/Register/register[0][10] ), .QN(n2424) );
  DFFRX1 \i_MIPS/Register/register_reg[0][11]  ( .D(\i_MIPS/Register/n1119 ), 
        .CK(clk), .RN(n5645), .Q(\i_MIPS/Register/register[0][11] ), .QN(n2593) );
  DFFRX1 \i_MIPS/Register/register_reg[0][12]  ( .D(\i_MIPS/Register/n1120 ), 
        .CK(clk), .RN(n5645), .Q(\i_MIPS/Register/register[0][12] ), .QN(n2456) );
  DFFRX1 \i_MIPS/Register/register_reg[0][13]  ( .D(\i_MIPS/Register/n1121 ), 
        .CK(clk), .RN(n5645), .Q(\i_MIPS/Register/register[0][13] ), .QN(n1056) );
  DFFRX1 \i_MIPS/Register/register_reg[0][14]  ( .D(\i_MIPS/Register/n1122 ), 
        .CK(clk), .RN(n5645), .Q(\i_MIPS/Register/register[0][14] ), .QN(n2216) );
  DFFRX1 \i_MIPS/Register/register_reg[0][15]  ( .D(\i_MIPS/Register/n1123 ), 
        .CK(clk), .RN(n5645), .Q(\i_MIPS/Register/register[0][15] ), .QN(n2595) );
  DFFRX1 \i_MIPS/Register/register_reg[0][16]  ( .D(\i_MIPS/Register/n1124 ), 
        .CK(clk), .RN(n5645), .Q(\i_MIPS/Register/register[0][16] ), .QN(n1054) );
  DFFRX1 \i_MIPS/Register/register_reg[0][17]  ( .D(\i_MIPS/Register/n1125 ), 
        .CK(clk), .RN(n5645), .Q(\i_MIPS/Register/register[0][17] ), .QN(n651)
         );
  DFFRX1 \i_MIPS/Register/register_reg[0][18]  ( .D(\i_MIPS/Register/n1126 ), 
        .CK(clk), .RN(n5645), .Q(\i_MIPS/Register/register[0][18] ), .QN(n2426) );
  DFFRX1 \i_MIPS/Register/register_reg[0][20]  ( .D(\i_MIPS/Register/n1128 ), 
        .CK(clk), .RN(n5645), .Q(\i_MIPS/Register/register[0][20] ), .QN(n2485) );
  DFFRX1 \i_MIPS/Register/register_reg[0][21]  ( .D(\i_MIPS/Register/n1129 ), 
        .CK(clk), .RN(n5645), .Q(\i_MIPS/Register/register[0][21] ), .QN(n2047) );
  DFFRX1 \i_MIPS/Register/register_reg[0][23]  ( .D(\i_MIPS/Register/n1131 ), 
        .CK(clk), .RN(n5644), .Q(\i_MIPS/Register/register[0][23] ), .QN(n2635) );
  DFFRX1 \i_MIPS/Register/register_reg[0][24]  ( .D(\i_MIPS/Register/n1132 ), 
        .CK(clk), .RN(n5644), .Q(\i_MIPS/Register/register[0][24] ), .QN(n2578) );
  DFFRX1 \i_MIPS/Register/register_reg[0][25]  ( .D(\i_MIPS/Register/n1133 ), 
        .CK(clk), .RN(n5644), .Q(\i_MIPS/Register/register[0][25] ), .QN(n2049) );
  DFFRX1 \i_MIPS/Register/register_reg[0][26]  ( .D(\i_MIPS/Register/n1134 ), 
        .CK(clk), .RN(n5644), .Q(\i_MIPS/Register/register[0][26] ), .QN(n2458) );
  DFFRX1 \i_MIPS/Register/register_reg[0][28]  ( .D(\i_MIPS/Register/n1136 ), 
        .CK(clk), .RN(n5644), .Q(\i_MIPS/Register/register[0][28] ), .QN(n2574) );
  DFFRX1 \i_MIPS/Register/register_reg[0][29]  ( .D(\i_MIPS/Register/n1137 ), 
        .CK(clk), .RN(n5644), .Q(\i_MIPS/Register/register[0][29] ), .QN(n1031) );
  DFFRX1 \i_MIPS/Register/register_reg[31][27]  ( .D(n11518), .CK(clk), .RN(
        n5707), .Q(\i_MIPS/Register/register[31][27] ), .QN(n1938) );
  DFFRX1 \i_MIPS/ID_EX_reg[114]  ( .D(\i_MIPS/n516 ), .CK(clk), .RN(n5738), 
        .Q(\i_MIPS/ID_EX[114] ), .QN(\i_MIPS/n319 ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][1]  ( .D(\i_MIPS/Register/n533 ), 
        .CK(clk), .RN(n5754), .Q(\i_MIPS/Register/register[18][1] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][10]  ( .D(\i_MIPS/Register/n542 ), 
        .CK(clk), .RN(n5753), .Q(\i_MIPS/Register/register[18][10] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][13]  ( .D(\i_MIPS/Register/n545 ), 
        .CK(clk), .RN(n5753), .Q(\i_MIPS/Register/register[18][13] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][18]  ( .D(\i_MIPS/Register/n550 ), 
        .CK(clk), .RN(n5753), .Q(\i_MIPS/Register/register[18][18] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][24]  ( .D(\i_MIPS/Register/n556 ), 
        .CK(clk), .RN(n5752), .Q(\i_MIPS/Register/register[18][24] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][1]  ( .D(\i_MIPS/Register/n1045 ), 
        .CK(clk), .RN(n5632), .Q(\i_MIPS/Register/register[2][1] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][10]  ( .D(\i_MIPS/Register/n1054 ), 
        .CK(clk), .RN(n5631), .Q(\i_MIPS/Register/register[2][10] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][13]  ( .D(\i_MIPS/Register/n1057 ), 
        .CK(clk), .RN(n5631), .Q(\i_MIPS/Register/register[2][13] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][18]  ( .D(\i_MIPS/Register/n1062 ), 
        .CK(clk), .RN(n5630), .Q(\i_MIPS/Register/register[2][18] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][24]  ( .D(\i_MIPS/Register/n1068 ), 
        .CK(clk), .RN(n5630), .Q(\i_MIPS/Register/register[2][24] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][0]  ( .D(\i_MIPS/Register/n276 ), 
        .CK(clk), .RN(n5776), .Q(\i_MIPS/Register/register[26][0] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][1]  ( .D(\i_MIPS/Register/n277 ), 
        .CK(clk), .RN(n5776), .Q(\i_MIPS/Register/register[26][1] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][2]  ( .D(\i_MIPS/Register/n278 ), 
        .CK(clk), .RN(n5776), .Q(\i_MIPS/Register/register[26][2] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][6]  ( .D(\i_MIPS/Register/n282 ), 
        .CK(clk), .RN(n5775), .Q(\i_MIPS/Register/register[26][6] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][7]  ( .D(\i_MIPS/Register/n283 ), 
        .CK(clk), .RN(n5775), .Q(\i_MIPS/Register/register[26][7] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][9]  ( .D(\i_MIPS/Register/n285 ), 
        .CK(clk), .RN(n5775), .Q(\i_MIPS/Register/register[26][9] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][10]  ( .D(\i_MIPS/Register/n286 ), 
        .CK(clk), .RN(n5775), .Q(\i_MIPS/Register/register[26][10] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][13]  ( .D(\i_MIPS/Register/n289 ), 
        .CK(clk), .RN(n5775), .Q(\i_MIPS/Register/register[26][13] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][14]  ( .D(\i_MIPS/Register/n290 ), 
        .CK(clk), .RN(n5775), .Q(\i_MIPS/Register/register[26][14] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][16]  ( .D(\i_MIPS/Register/n292 ), 
        .CK(clk), .RN(n5774), .Q(\i_MIPS/Register/register[26][16] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][18]  ( .D(\i_MIPS/Register/n294 ), 
        .CK(clk), .RN(n5774), .Q(\i_MIPS/Register/register[26][18] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][20]  ( .D(\i_MIPS/Register/n296 ), 
        .CK(clk), .RN(n5774), .Q(\i_MIPS/Register/register[26][20] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][21]  ( .D(\i_MIPS/Register/n297 ), 
        .CK(clk), .RN(n5774), .Q(\i_MIPS/Register/register[26][21] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][23]  ( .D(\i_MIPS/Register/n299 ), 
        .CK(clk), .RN(n5774), .Q(\i_MIPS/Register/register[26][23] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][24]  ( .D(\i_MIPS/Register/n300 ), 
        .CK(clk), .RN(n5774), .Q(\i_MIPS/Register/register[26][24] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][28]  ( .D(\i_MIPS/Register/n304 ), 
        .CK(clk), .RN(n5773), .Q(\i_MIPS/Register/register[26][28] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][1]  ( .D(\i_MIPS/Register/n789 ), 
        .CK(clk), .RN(n5653), .Q(\i_MIPS/Register/register[10][1] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][2]  ( .D(\i_MIPS/Register/n790 ), 
        .CK(clk), .RN(n5653), .Q(\i_MIPS/Register/register[10][2] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][6]  ( .D(\i_MIPS/Register/n794 ), 
        .CK(clk), .RN(n5653), .Q(\i_MIPS/Register/register[10][6] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][9]  ( .D(\i_MIPS/Register/n797 ), 
        .CK(clk), .RN(n5652), .Q(\i_MIPS/Register/register[10][9] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][10]  ( .D(\i_MIPS/Register/n798 ), 
        .CK(clk), .RN(n5652), .Q(\i_MIPS/Register/register[10][10] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][13]  ( .D(\i_MIPS/Register/n801 ), 
        .CK(clk), .RN(n5652), .Q(\i_MIPS/Register/register[10][13] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][14]  ( .D(\i_MIPS/Register/n802 ), 
        .CK(clk), .RN(n5652), .Q(\i_MIPS/Register/register[10][14] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][16]  ( .D(\i_MIPS/Register/n804 ), 
        .CK(clk), .RN(n5652), .Q(\i_MIPS/Register/register[10][16] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][18]  ( .D(\i_MIPS/Register/n806 ), 
        .CK(clk), .RN(n5652), .Q(\i_MIPS/Register/register[10][18] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][20]  ( .D(\i_MIPS/Register/n808 ), 
        .CK(clk), .RN(n5652), .Q(\i_MIPS/Register/register[10][20] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][21]  ( .D(\i_MIPS/Register/n809 ), 
        .CK(clk), .RN(n5651), .Q(\i_MIPS/Register/register[10][21] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][23]  ( .D(\i_MIPS/Register/n811 ), 
        .CK(clk), .RN(n5651), .Q(\i_MIPS/Register/register[10][23] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][24]  ( .D(\i_MIPS/Register/n812 ), 
        .CK(clk), .RN(n5651), .Q(\i_MIPS/Register/register[10][24] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][28]  ( .D(\i_MIPS/Register/n816 ), 
        .CK(clk), .RN(n5651), .Q(\i_MIPS/Register/register[10][28] ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[0]  ( .D(\i_MIPS/n563 ), .CK(clk), .RN(n5713), .Q(
        \i_MIPS/EX_MEM_0 ), .QN(\i_MIPS/n373 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[16]  ( .D(\i_MIPS/n458 ), .CK(clk), .RN(n5744), 
        .Q(n12948) );
  DFFRX1 \i_MIPS/EX_MEM_reg[30]  ( .D(\i_MIPS/n444 ), .CK(clk), .RN(n5745), 
        .Q(n12934) );
  DFFRX1 \i_MIPS/EX_MEM_reg[19]  ( .D(\i_MIPS/n455 ), .CK(clk), .RN(n5744), 
        .Q(n12945), .QN(n3409) );
  DFFRX1 \i_MIPS/EX_MEM_reg[27]  ( .D(\i_MIPS/n447 ), .CK(clk), .RN(n5745), 
        .Q(n12937), .QN(n3716) );
  DFFRX1 \i_MIPS/EX_MEM_reg[20]  ( .D(\i_MIPS/n454 ), .CK(clk), .RN(n5744), 
        .Q(n12944) );
  DFFRX1 \i_MIPS/EX_MEM_reg[32]  ( .D(\i_MIPS/n442 ), .CK(clk), .RN(n5745), 
        .Q(n12932) );
  DFFRXL \i_MIPS/EX_MEM_reg[35]  ( .D(\i_MIPS/n439 ), .CK(clk), .RN(n5746), 
        .Q(n12929), .QN(n3411) );
  DFFRX1 \i_MIPS/EX_MEM_reg[34]  ( .D(\i_MIPS/n440 ), .CK(clk), .RN(n5746), 
        .Q(n12930), .QN(n4626) );
  DFFRX1 \i_MIPS/EX_MEM_reg[13]  ( .D(\i_MIPS/n461 ), .CK(clk), .RN(n5744), 
        .Q(n12951), .QN(n1776) );
  DFFRX2 \i_MIPS/ID_EX_reg[34]  ( .D(\i_MIPS/n537 ), .CK(clk), .RN(n5715), .Q(
        \i_MIPS/ALUin1[25] ), .QN(\i_MIPS/n346 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[33]  ( .D(\i_MIPS/n538 ), .CK(clk), .RN(n5715), .Q(
        \i_MIPS/ALUin1[24] ), .QN(\i_MIPS/n347 ) );
  DFFRX2 \i_MIPS/EX_MEM_reg[3]  ( .D(\i_MIPS/n524 ), .CK(clk), .RN(n5716), .Q(
        DCACHE_ren), .QN(\i_MIPS/n334 ) );
  DFFRX2 \i_MIPS/EX_MEM_reg[72]  ( .D(\i_MIPS/n474 ), .CK(clk), .RN(n5743), 
        .Q(\i_MIPS/Reg_W[3] ), .QN(n4543) );
  DFFRX2 \i_MIPS/EX_MEM_reg[69]  ( .D(\i_MIPS/n477 ), .CK(clk), .RN(n5743), 
        .Q(\i_MIPS/Reg_W[0] ), .QN(n415) );
  DFFRX2 \i_MIPS/EX_MEM_reg[70]  ( .D(\i_MIPS/n476 ), .CK(clk), .RN(n5743), 
        .Q(\i_MIPS/Reg_W[1] ), .QN(n303) );
  DFFRX2 \i_MIPS/EX_MEM_reg[73]  ( .D(\i_MIPS/n473 ), .CK(clk), .RN(n5743), 
        .Q(\i_MIPS/Reg_W[4] ), .QN(n4542) );
  DFFRX2 \i_MIPS/EX_MEM_reg[71]  ( .D(\i_MIPS/n475 ), .CK(clk), .RN(n5743), 
        .Q(\i_MIPS/Reg_W[2] ), .QN(n4534) );
  DFFRX1 \i_MIPS/EX_MEM_reg[24]  ( .D(\i_MIPS/n450 ), .CK(clk), .RN(n5745), 
        .Q(n12940), .QN(n4633) );
  DFFRX1 \i_MIPS/EX_MEM_reg[22]  ( .D(\i_MIPS/n452 ), .CK(clk), .RN(n5745), 
        .Q(n12942), .QN(n4598) );
  DFFRX1 \i_MIPS/EX_MEM_reg[18]  ( .D(\i_MIPS/n456 ), .CK(clk), .RN(n5744), 
        .Q(n12946), .QN(n4596) );
  DFFRX1 \i_MIPS/EX_MEM_reg[17]  ( .D(\i_MIPS/n457 ), .CK(clk), .RN(n5744), 
        .Q(n12947), .QN(n4594) );
  DFFRX1 \i_MIPS/EX_MEM_reg[23]  ( .D(\i_MIPS/n451 ), .CK(clk), .RN(n5745), 
        .Q(n12941), .QN(n4629) );
  DFFRX1 \D_cache/cache_reg[0][139]  ( .D(\D_cache/n684 ), .CK(clk), .RN(n5930), .Q(\D_cache/cache[0][139] ), .QN(n3347) );
  DFFRX1 \D_cache/cache_reg[1][139]  ( .D(\D_cache/n683 ), .CK(clk), .RN(n5930), .Q(\D_cache/cache[1][139] ), .QN(n405) );
  DFFRX1 \D_cache/cache_reg[4][139]  ( .D(\D_cache/n680 ), .CK(clk), .RN(n5930), .Q(\D_cache/cache[4][139] ), .QN(n3344) );
  DFFRX1 \D_cache/cache_reg[5][139]  ( .D(\D_cache/n679 ), .CK(clk), .RN(n5930), .Q(\D_cache/cache[5][139] ), .QN(n1730) );
  DFFRX1 \D_cache/cache_reg[0][144]  ( .D(\D_cache/n644 ), .CK(clk), .RN(n5927), .Q(\D_cache/cache[0][144] ), .QN(n3348) );
  DFFRX1 \D_cache/cache_reg[1][144]  ( .D(\D_cache/n643 ), .CK(clk), .RN(n5927), .Q(\D_cache/cache[1][144] ), .QN(n1732) );
  DFFRX1 \D_cache/cache_reg[4][144]  ( .D(\D_cache/n640 ), .CK(clk), .RN(n5927), .Q(\D_cache/cache[4][144] ), .QN(n3349) );
  DFFRX1 \D_cache/cache_reg[5][144]  ( .D(\D_cache/n639 ), .CK(clk), .RN(n5927), .Q(\D_cache/cache[5][144] ), .QN(n1733) );
  DFFRHQX8 \i_MIPS/ID_EX_reg[8]  ( .D(\i_MIPS/n470 ), .CK(clk), .RN(n5743), 
        .Q(n4323) );
  DFFRX1 \D_cache/cache_reg[7][151]  ( .D(\D_cache/n581 ), .CK(clk), .RN(n5942), .Q(\D_cache/cache[7][151] ), .QN(n3360) );
  DFFRX1 \D_cache/cache_reg[1][152]  ( .D(\D_cache/n579 ), .CK(clk), .RN(n5941), .Q(\D_cache/cache[1][152] ), .QN(n1731) );
  DFFRX1 \D_cache/cache_reg[1][140]  ( .D(\D_cache/n675 ), .CK(clk), .RN(n5930), .Q(\D_cache/cache[1][140] ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[7]  ( .D(\i_MIPS/n467 ), .CK(clk), .RN(n5743), .Q(
        n12955), .QN(n2651) );
  DFFRX4 \i_MIPS/ID_EX_reg[9]  ( .D(\i_MIPS/n562 ), .CK(clk), .RN(n5713), .Q(
        \i_MIPS/ALUin1[0] ), .QN(\i_MIPS/n371 ) );
  DFFRX4 \i_MIPS/PC/PC_o_reg[12]  ( .D(\i_MIPS/PC/n46 ), .CK(clk), .RN(n5711), 
        .Q(ICACHE_addr[10]), .QN(\i_MIPS/PC/n14 ) );
  DFFRX4 \i_MIPS/ID_EX_reg[88]  ( .D(\i_MIPS/n497 ), .CK(clk), .RN(n5741), .Q(
        \i_MIPS/ID_EX[88] ) );
  DFFRX4 \i_MIPS/PC/PC_o_reg[7]  ( .D(\i_MIPS/PC/n41 ), .CK(clk), .RN(n5711), 
        .Q(ICACHE_addr[5]), .QN(\i_MIPS/PC/n9 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[44]  ( .D(\i_MIPS/n431 ), .CK(clk), .RN(n5726), 
        .QN(\i_MIPS/n303 ) );
  DFFRHQX8 \i_MIPS/EX_MEM_reg[10]  ( .D(\i_MIPS/n464 ), .CK(clk), .RN(n5744), 
        .Q(n4382) );
  DFFRX4 \i_MIPS/ID_EX_reg[106]  ( .D(\i_MIPS/n519 ), .CK(clk), .RN(n5737), 
        .Q(\i_MIPS/ID_EX[106] ), .QN(\i_MIPS/n325 ) );
  DFFRX4 \i_MIPS/PC/PC_o_reg[10]  ( .D(\i_MIPS/PC/n44 ), .CK(clk), .RN(n5711), 
        .Q(ICACHE_addr[8]), .QN(\i_MIPS/PC/n12 ) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[26]  ( .D(\i_MIPS/PC/n60 ), .CK(clk), .RN(n5710), 
        .Q(ICACHE_addr[24]), .QN(\i_MIPS/PC/n28 ) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[1]  ( .D(\i_MIPS/PC/n35 ), .CK(clk), .RN(n5712), 
        .Q(\i_MIPS/PC_o[1] ), .QN(\i_MIPS/PC/n3 ) );
  DFFRX4 \D_cache/cache_reg[0][21]  ( .D(\D_cache/n1628 ), .CK(clk), .RN(n5690), .Q(\D_cache/cache[0][21] ), .QN(n2648) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[0]  ( .D(\i_MIPS/PC/n34 ), .CK(clk), .RN(n5712), 
        .Q(\i_MIPS/BranchAddr[0] ), .QN(\i_MIPS/PC/n2 ) );
  DFFRX4 \D_cache/cache_reg[0][48]  ( .D(\D_cache/n1412 ), .CK(clk), .RN(n5672), .Q(\D_cache/cache[0][48] ), .QN(n2967) );
  DFFRX4 \D_cache/cache_reg[0][8]  ( .D(\D_cache/n1732 ), .CK(clk), .RN(n5638), 
        .Q(\D_cache/cache[0][8] ), .QN(n2419) );
  DFFRX4 \D_cache/cache_reg[0][0]  ( .D(\D_cache/n1795 ), .CK(clk), .RN(n5644), 
        .Q(\D_cache/cache[0][0] ), .QN(n3333) );
  DFFRX4 \i_MIPS/PC/PC_o_reg[29]  ( .D(\i_MIPS/PC/n63 ), .CK(clk), .RN(n5709), 
        .Q(ICACHE_addr[27]), .QN(\i_MIPS/PC/n31 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[96]  ( .D(\i_MIPS/N122 ), .CK(clk), .RN(n5627), .Q(
        \i_MIPS/IF_ID[96] ), .QN(\i_MIPS/n182 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[73]  ( .D(\i_MIPS/N99 ), .CK(clk), .RN(n5735), .Q(
        \i_MIPS/IF_ID[73] ), .QN(\i_MIPS/n245 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[85]  ( .D(\i_MIPS/N111 ), .CK(clk), .RN(n5736), .Q(
        \i_MIPS/IF_ID[85] ), .QN(\i_MIPS/n171 ) );
  DFFRX4 \i_MIPS/ID_EX_reg[107]  ( .D(\i_MIPS/n520 ), .CK(clk), .RN(n5736), 
        .Q(\i_MIPS/ID_EX[107] ), .QN(\i_MIPS/n327 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[40]  ( .D(\i_MIPS/N66 ), .CK(clk), .RN(n5739), .Q(
        \i_MIPS/Sign_Extend_ID[8] ), .QN(\i_MIPS/n223 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[88]  ( .D(\i_MIPS/N114 ), .CK(clk), .RN(n5736), .Q(
        \i_MIPS/IF_ID[88] ), .QN(\i_MIPS/n174 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[82]  ( .D(\i_MIPS/N108 ), .CK(clk), .RN(n5735), .Q(
        \i_MIPS/IF_ID[82] ), .QN(\i_MIPS/n168 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[80]  ( .D(\i_MIPS/N106 ), .CK(clk), .RN(n5735), .Q(
        \i_MIPS/IF_ID[80] ), .QN(\i_MIPS/n166 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[3]  ( .D(\i_MIPS/N29 ), .CK(clk), .RN(n5732), .QN(
        \i_MIPS/n186 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[2]  ( .D(\i_MIPS/N28 ), .CK(clk), .RN(n5732), .QN(
        \i_MIPS/n185 ) );
  DFFRX4 \i_MIPS/IF_ID_reg[57]  ( .D(\i_MIPS/N83 ), .CK(clk), .RN(n5737), .Q(
        \i_MIPS/IR_ID[25] ), .QN(\i_MIPS/n235 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[79]  ( .D(\i_MIPS/N105 ), .CK(clk), .RN(n5735), .Q(
        \i_MIPS/IF_ID[79] ), .QN(\i_MIPS/n165 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[33]  ( .D(\i_MIPS/N59 ), .CK(clk), .RN(n5739), .Q(
        \i_MIPS/Sign_Extend_ID[1] ), .QN(\i_MIPS/n216 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[37]  ( .D(\i_MIPS/N63 ), .CK(clk), .RN(n5739), .Q(
        \i_MIPS/Sign_Extend_ID[5] ), .QN(\i_MIPS/n220 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[75]  ( .D(\i_MIPS/N101 ), .CK(clk), .RN(n5735), .Q(
        \i_MIPS/IF_ID[75] ), .QN(\i_MIPS/n161 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[92]  ( .D(\i_MIPS/N118 ), .CK(clk), .RN(n5736), .Q(
        \i_MIPS/IF_ID[92] ), .QN(\i_MIPS/n178 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[71]  ( .D(\i_MIPS/N97 ), .CK(clk), .RN(n5734), .Q(
        \i_MIPS/IF_ID[71] ), .QN(\i_MIPS/n243 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[91]  ( .D(\i_MIPS/N117 ), .CK(clk), .RN(n5736), .Q(
        \i_MIPS/IF_ID[91] ), .QN(\i_MIPS/n177 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[74]  ( .D(\i_MIPS/N100 ), .CK(clk), .RN(n5731), .Q(
        \i_MIPS/IF_ID[74] ), .QN(\i_MIPS/n160 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[35]  ( .D(\i_MIPS/N61 ), .CK(clk), .RN(n5739), .Q(
        \i_MIPS/Sign_Extend_ID[3] ), .QN(\i_MIPS/n218 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[77]  ( .D(\i_MIPS/N103 ), .CK(clk), .RN(n5735), .Q(
        \i_MIPS/IF_ID[77] ), .QN(\i_MIPS/n163 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[90]  ( .D(\i_MIPS/N116 ), .CK(clk), .RN(n5736), .Q(
        \i_MIPS/IF_ID[90] ), .QN(\i_MIPS/n176 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[38]  ( .D(\i_MIPS/N64 ), .CK(clk), .RN(n5739), .Q(
        \i_MIPS/Sign_Extend_ID[6] ), .QN(\i_MIPS/n221 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[39]  ( .D(\i_MIPS/N65 ), .CK(clk), .RN(n5739), .QN(
        \i_MIPS/n222 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[36]  ( .D(\i_MIPS/N62 ), .CK(clk), .RN(n5739), .Q(
        \i_MIPS/Sign_Extend_ID[4] ), .QN(\i_MIPS/n219 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[41]  ( .D(\i_MIPS/N67 ), .CK(clk), .RN(n5739), .QN(
        \i_MIPS/n224 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[42]  ( .D(\i_MIPS/N68 ), .CK(clk), .RN(n5739), .QN(
        \i_MIPS/n225 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[32]  ( .D(\i_MIPS/N58 ), .CK(clk), .RN(n5715), .Q(
        \i_MIPS/Sign_Extend_ID[0] ), .QN(\i_MIPS/n215 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[34]  ( .D(\i_MIPS/N60 ), .CK(clk), .RN(n5739), .Q(
        \i_MIPS/Sign_Extend_ID[2] ), .QN(\i_MIPS/n217 ) );
  DFFRX4 \i_MIPS/PC/PC_o_reg[31]  ( .D(\i_MIPS/PC/n65 ), .CK(clk), .RN(n5709), 
        .Q(ICACHE_addr[29]), .QN(\i_MIPS/PC/n33 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[86]  ( .D(\i_MIPS/N112 ), .CK(clk), .RN(n5736), .Q(
        \i_MIPS/IF_ID[86] ), .QN(\i_MIPS/n172 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[69]  ( .D(\i_MIPS/N95 ), .CK(clk), .RN(n5734), .Q(
        \i_MIPS/IF_ID[69] ), .QN(\i_MIPS/n241 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[70]  ( .D(\i_MIPS/N96 ), .CK(clk), .RN(n5734), .Q(
        \i_MIPS/IF_ID[70] ), .QN(\i_MIPS/n242 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[68]  ( .D(\i_MIPS/N94 ), .CK(clk), .RN(n5734), .Q(
        \i_MIPS/IF_ID[68] ), .QN(\i_MIPS/n240 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[81]  ( .D(\i_MIPS/N107 ), .CK(clk), .RN(n5735), .Q(
        \i_MIPS/IF_ID[81] ), .QN(\i_MIPS/n167 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[72]  ( .D(\i_MIPS/N98 ), .CK(clk), .RN(n5735), .Q(
        \i_MIPS/IF_ID[72] ), .QN(\i_MIPS/n244 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[84]  ( .D(\i_MIPS/N110 ), .CK(clk), .RN(n5735), .Q(
        \i_MIPS/IF_ID[84] ), .QN(\i_MIPS/n170 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[76]  ( .D(\i_MIPS/N102 ), .CK(clk), .RN(n5735), .Q(
        \i_MIPS/IF_ID[76] ), .QN(\i_MIPS/n162 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[87]  ( .D(\i_MIPS/N113 ), .CK(clk), .RN(n5736), .Q(
        \i_MIPS/IF_ID[87] ), .QN(\i_MIPS/n173 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[78]  ( .D(\i_MIPS/N104 ), .CK(clk), .RN(n5735), .Q(
        \i_MIPS/IF_ID[78] ), .QN(\i_MIPS/n164 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[94]  ( .D(\i_MIPS/N120 ), .CK(clk), .RN(n5736), .Q(
        \i_MIPS/IF_ID[94] ), .QN(\i_MIPS/n180 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[44]  ( .D(\i_MIPS/N70 ), .CK(clk), .RN(n5738), .QN(
        \i_MIPS/n227 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[45]  ( .D(\i_MIPS/N71 ), .CK(clk), .RN(n5738), .QN(
        \i_MIPS/n228 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[46]  ( .D(\i_MIPS/N72 ), .CK(clk), .RN(n5738), .QN(
        \i_MIPS/n229 ) );
  DFFRX4 \i_MIPS/PC/PC_o_reg[30]  ( .D(\i_MIPS/PC/n64 ), .CK(clk), .RN(n5709), 
        .Q(ICACHE_addr[28]), .QN(\i_MIPS/PC/n32 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[43]  ( .D(\i_MIPS/N69 ), .CK(clk), .RN(n5738), .QN(
        \i_MIPS/n226 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[47]  ( .D(\i_MIPS/N73 ), .CK(clk), .RN(n5738), .Q(
        \i_MIPS/Sign_Extend_ID[31] ), .QN(\i_MIPS/n230 ) );
  DFFRX4 \i_MIPS/ID_EX_reg[108]  ( .D(\i_MIPS/n521 ), .CK(clk), .RN(n5741), 
        .Q(net133414), .QN(\i_MIPS/n329 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[20]  ( .D(\i_MIPS/N46 ), .CK(clk), .RN(n5733), .QN(
        \i_MIPS/n203 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[16]  ( .D(\i_MIPS/N42 ), .CK(clk), .RN(n5733), .QN(
        \i_MIPS/n199 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[12]  ( .D(\i_MIPS/N38 ), .CK(clk), .RN(n5732), .QN(
        \i_MIPS/n195 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[11]  ( .D(\i_MIPS/N37 ), .CK(clk), .RN(n5732), .QN(
        \i_MIPS/n194 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[15]  ( .D(\i_MIPS/N41 ), .CK(clk), .RN(n5733), .QN(
        \i_MIPS/n198 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[14]  ( .D(\i_MIPS/N40 ), .CK(clk), .RN(n5733), .QN(
        \i_MIPS/n197 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[28]  ( .D(\i_MIPS/N54 ), .CK(clk), .RN(n5734), .Q(
        \i_MIPS/IF_ID_28 ), .QN(\i_MIPS/n211 ) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[21]  ( .D(\i_MIPS/PC/n55 ), .CK(clk), .RN(n5710), 
        .Q(ICACHE_addr[19]), .QN(\i_MIPS/PC/n23 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[27]  ( .D(\i_MIPS/N53 ), .CK(clk), .RN(n5734), .QN(
        \i_MIPS/n210 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[9]  ( .D(\i_MIPS/N35 ), .CK(clk), .RN(n5732), .QN(
        \i_MIPS/n192 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[7]  ( .D(\i_MIPS/N33 ), .CK(clk), .RN(n5732), .QN(
        \i_MIPS/n190 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[23]  ( .D(\i_MIPS/N49 ), .CK(clk), .RN(n5733), .QN(
        \i_MIPS/n206 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[6]  ( .D(\i_MIPS/N32 ), .CK(clk), .RN(n5732), .QN(
        \i_MIPS/n189 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[67]  ( .D(\i_MIPS/N93 ), .CK(clk), .RN(n5734), .Q(
        \i_MIPS/IF_ID[67] ), .QN(\i_MIPS/n239 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[10]  ( .D(\i_MIPS/N36 ), .CK(clk), .RN(n5732), .QN(
        \i_MIPS/n193 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[5]  ( .D(\i_MIPS/N31 ), .CK(clk), .RN(n5732), .QN(
        \i_MIPS/n188 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[26]  ( .D(\i_MIPS/N52 ), .CK(clk), .RN(n5734), .QN(
        \i_MIPS/n209 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[8]  ( .D(\i_MIPS/N34 ), .CK(clk), .RN(n5732), .QN(
        \i_MIPS/n191 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[18]  ( .D(\i_MIPS/N44 ), .CK(clk), .RN(n5733), .QN(
        \i_MIPS/n201 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[24]  ( .D(\i_MIPS/N50 ), .CK(clk), .RN(n5733), .QN(
        \i_MIPS/n207 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[25]  ( .D(\i_MIPS/N51 ), .CK(clk), .RN(n5733), .QN(
        \i_MIPS/n208 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[31]  ( .D(\i_MIPS/N57 ), .CK(clk), .RN(n5786), .Q(
        \i_MIPS/IF_ID_31 ), .QN(\i_MIPS/n214 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[29]  ( .D(\i_MIPS/N55 ), .CK(clk), .RN(n5734), .Q(
        \i_MIPS/IF_ID_29 ), .QN(\i_MIPS/n212 ) );
  DFFRX4 \i_MIPS/PC/PC_o_reg[28]  ( .D(\i_MIPS/PC/n62 ), .CK(clk), .RN(n5709), 
        .Q(ICACHE_addr[26]), .QN(\i_MIPS/PC/n30 ) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[19]  ( .D(\i_MIPS/PC/n53 ), .CK(clk), .RN(n5710), 
        .Q(ICACHE_addr[17]), .QN(\i_MIPS/PC/n21 ) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[16]  ( .D(\i_MIPS/PC/n50 ), .CK(clk), .RN(n5710), 
        .Q(ICACHE_addr[14]), .QN(\i_MIPS/PC/n18 ) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[15]  ( .D(\i_MIPS/PC/n49 ), .CK(clk), .RN(n5711), 
        .Q(ICACHE_addr[13]), .QN(\i_MIPS/PC/n17 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[87]  ( .D(\i_MIPS/n498 ), .CK(clk), .RN(n5741), 
        .QN(n4540) );
  DFFRX2 \i_MIPS/EX_MEM_reg[1]  ( .D(\i_MIPS/n526 ), .CK(clk), .RN(n5716), .Q(
        \i_MIPS/EX_MEM_1 ), .QN(\i_MIPS/n336 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[93]  ( .D(\i_MIPS/N119 ), .CK(clk), .RN(n5736), .Q(
        \i_MIPS/IF_ID[93] ), .QN(\i_MIPS/n179 ) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[24]  ( .D(\i_MIPS/PC/n58 ), .CK(clk), .RN(n5710), 
        .Q(ICACHE_addr[22]), .QN(\i_MIPS/PC/n26 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[111]  ( .D(\i_MIPS/n513 ), .CK(clk), .RN(n5738), 
        .QN(\i_MIPS/n313 ) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[23]  ( .D(\i_MIPS/PC/n57 ), .CK(clk), .RN(n5710), 
        .Q(ICACHE_addr[21]), .QN(\i_MIPS/PC/n25 ) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[14]  ( .D(\i_MIPS/PC/n48 ), .CK(clk), .RN(n5711), 
        .Q(ICACHE_addr[12]), .QN(\i_MIPS/PC/n16 ) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[13]  ( .D(\i_MIPS/PC/n47 ), .CK(clk), .RN(n5711), 
        .Q(ICACHE_addr[11]), .QN(\i_MIPS/PC/n15 ) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[17]  ( .D(\i_MIPS/PC/n51 ), .CK(clk), .RN(n5710), 
        .Q(ICACHE_addr[15]), .QN(\i_MIPS/PC/n19 ) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[20]  ( .D(\i_MIPS/PC/n54 ), .CK(clk), .RN(n5710), 
        .Q(ICACHE_addr[18]), .QN(\i_MIPS/PC/n22 ) );
  DFFRX4 \D_cache/cache_reg[0][50]  ( .D(\D_cache/n1396 ), .CK(clk), .RN(n5670), .Q(\D_cache/cache[0][50] ), .QN(n2963) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[18]  ( .D(\i_MIPS/PC/n52 ), .CK(clk), .RN(n5710), 
        .Q(ICACHE_addr[16]), .QN(\i_MIPS/PC/n20 ) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[27]  ( .D(\i_MIPS/PC/n61 ), .CK(clk), .RN(n5710), 
        .Q(ICACHE_addr[25]), .QN(\i_MIPS/PC/n29 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[102]  ( .D(\i_MIPS/n483 ), .CK(clk), .RN(n5742), 
        .Q(\i_MIPS/ID_EX[102] ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[15]  ( .D(\i_MIPS/n459 ), .CK(clk), .RN(n5744), 
        .Q(n12949) );
  DFFRHQX8 \i_MIPS/PC/PC_o_reg[4]  ( .D(\i_MIPS/PC/n38 ), .CK(clk), .RN(n5712), 
        .Q(n3783) );
  DFFRX2 \i_MIPS/IF_ID_reg[58]  ( .D(\i_MIPS/N84 ), .CK(clk), .RN(n5737), .Q(
        \i_MIPS/IR_ID[26] ), .QN(\i_MIPS/n322 ) );
  DFFRX4 \i_MIPS/ID_EX_reg[19]  ( .D(\i_MIPS/n552 ), .CK(clk), .RN(n5713), .Q(
        \i_MIPS/ALUin1[10] ), .QN(\i_MIPS/n361 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[42]  ( .D(\i_MIPS/n435 ), .CK(clk), .RN(n5746), .Q(
        \i_MIPS/ID_EX[42] ), .QN(\i_MIPS/n307 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[28]  ( .D(\i_MIPS/n446 ), .CK(clk), .RN(n5745), 
        .Q(n12936), .QN(n4631) );
  DFFRX4 \i_MIPS/ID_EX_reg[52]  ( .D(\i_MIPS/n415 ), .CK(clk), .RN(n5728), .Q(
        n3699), .QN(\i_MIPS/n287 ) );
  DFFRX4 \i_MIPS/ID_EX_reg[51]  ( .D(\i_MIPS/n417 ), .CK(clk), .RN(n5728), .Q(
        n3695), .QN(\i_MIPS/n289 ) );
  DFFRX4 \i_MIPS/ID_EX_reg[109]  ( .D(\i_MIPS/n522 ), .CK(clk), .RN(n5716), 
        .QN(\i_MIPS/n331 ) );
  DFFRX4 \i_MIPS/ID_EX_reg[50]  ( .D(\i_MIPS/n419 ), .CK(clk), .RN(n5727), .Q(
        \i_MIPS/ID_EX[50] ), .QN(\i_MIPS/n291 ) );
  DFFRX4 \i_MIPS/ID_EX_reg[110]  ( .D(\i_MIPS/n523 ), .CK(clk), .RN(n5716), 
        .QN(\i_MIPS/n333 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[112]  ( .D(\i_MIPS/n514 ), .CK(clk), .RN(n5738), 
        .Q(\i_MIPS/ID_EX[112] ), .QN(\i_MIPS/n315 ) );
  DFFRHQX4 \i_MIPS/EX_MEM_reg[11]  ( .D(\i_MIPS/n463 ), .CK(clk), .RN(n5744), 
        .Q(n4296) );
  DFFRX1 \i_MIPS/EX_MEM_reg[29]  ( .D(\i_MIPS/n445 ), .CK(clk), .RN(n5745), 
        .Q(n12935), .QN(n3763) );
  DFFRX1 \i_MIPS/EX_MEM_reg[36]  ( .D(\i_MIPS/n438 ), .CK(clk), .RN(n5746), 
        .Q(n12928), .QN(n3928) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[22]  ( .D(\i_MIPS/PC/n56 ), .CK(clk), .RN(n5710), 
        .Q(ICACHE_addr[20]), .QN(\i_MIPS/PC/n24 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[60]  ( .D(\i_MIPS/N86 ), .CK(clk), .RN(n5736), .Q(
        \i_MIPS/IR_ID[28] ), .QN(\i_MIPS/n326 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[59]  ( .D(\i_MIPS/N85 ), .CK(clk), .RN(n5737), .Q(
        \i_MIPS/IR_ID[27] ), .QN(\i_MIPS/n324 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[65]  ( .D(\i_MIPS/n389 ), .CK(clk), .RN(n5730), .Q(
        n3613), .QN(\i_MIPS/n261 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[64]  ( .D(\i_MIPS/n391 ), .CK(clk), .RN(n5730), .Q(
        \i_MIPS/ID_EX[64] ), .QN(\i_MIPS/n263 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[63]  ( .D(\i_MIPS/n393 ), .CK(clk), .RN(n5730), .Q(
        n3611), .QN(\i_MIPS/n265 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[72]  ( .D(\i_MIPS/n375 ), .CK(clk), .RN(n5731), .Q(
        n3610), .QN(\i_MIPS/n247 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[63]  ( .D(\i_MIPS/N89 ), .CK(clk), .RN(n5716), .Q(
        \i_MIPS/IR_ID[31] ), .QN(\i_MIPS/n332 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[52]  ( .D(\i_MIPS/N78 ), .CK(clk), .RN(n5737), .Q(
        \i_MIPS/IR_ID[20] ), .QN(\i_MIPS/n320 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[4]  ( .D(\i_MIPS/N30 ), .CK(clk), .RN(n5732), .QN(
        \i_MIPS/n187 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[17]  ( .D(\i_MIPS/N43 ), .CK(clk), .RN(n5733), .QN(
        \i_MIPS/n200 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[21]  ( .D(\i_MIPS/N47 ), .CK(clk), .RN(n5733), .QN(
        \i_MIPS/n204 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[19]  ( .D(\i_MIPS/N45 ), .CK(clk), .RN(n5733), .QN(
        \i_MIPS/n202 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[22]  ( .D(\i_MIPS/N48 ), .CK(clk), .RN(n5733), .QN(
        \i_MIPS/n205 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[60]  ( .D(\i_MIPS/n399 ), .CK(clk), .RN(n5729), .Q(
        n3604), .QN(\i_MIPS/n271 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[53]  ( .D(\i_MIPS/n413 ), .CK(clk), .RN(n5728), .Q(
        n3601), .QN(\i_MIPS/n285 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[48]  ( .D(\i_MIPS/n423 ), .CK(clk), .RN(n5727), .Q(
        n3596), .QN(\i_MIPS/n295 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[45]  ( .D(\i_MIPS/n429 ), .CK(clk), .RN(n5727), .Q(
        n3593), .QN(\i_MIPS/n301 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[25]  ( .D(\i_MIPS/n449 ), .CK(clk), .RN(n5745), 
        .Q(n12939), .QN(n4593) );
  DFFRX1 \I_cache/cache_reg[3][22]  ( .D(n12608), .CK(clk), .RN(n5924), .Q(
        \I_cache/cache[3][22] ), .QN(n3592) );
  DFFRX1 \I_cache/cache_reg[5][22]  ( .D(n12606), .CK(clk), .RN(n5924), .Q(
        \I_cache/cache[5][22] ), .QN(n3591) );
  DFFRX1 \I_cache/cache_reg[6][22]  ( .D(n12605), .CK(clk), .RN(n5924), .Q(
        \I_cache/cache[6][22] ), .QN(n3590) );
  DFFRX2 \I_cache/cache_reg[2][118]  ( .D(n11841), .CK(clk), .RN(n5860), .Q(
        \I_cache/cache[2][118] ), .QN(n3589) );
  DFFRX1 \I_cache/cache_reg[1][22]  ( .D(n12610), .CK(clk), .RN(n5925), .Q(
        \I_cache/cache[1][22] ), .QN(n3588) );
  DFFRX2 \i_MIPS/IF_ID_reg[97]  ( .D(\i_MIPS/N123 ), .CK(clk), .RN(n5742), .Q(
        \i_MIPS/IF_ID[97] ), .QN(\i_MIPS/n567 ) );
  DFFRX1 \I_cache/cache_reg[6][154]  ( .D(n11549), .CK(clk), .RN(n5841), .Q(
        \I_cache/cache[6][154] ), .QN(n3408) );
  DFFRX1 \I_cache/cache_reg[3][154]  ( .D(n11552), .CK(clk), .RN(n5836), .Q(
        \I_cache/cache[3][154] ), .QN(n3407) );
  DFFRX1 \I_cache/cache_reg[1][154]  ( .D(n11554), .CK(clk), .RN(n5836), .Q(
        \I_cache/cache[1][154] ), .QN(n3406) );
  DFFRX2 \i_MIPS/IF_ID_reg[56]  ( .D(\i_MIPS/N82 ), .CK(clk), .RN(n5737), .Q(
        \i_MIPS/IR_ID[24] ), .QN(\i_MIPS/n234 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[38]  ( .D(\i_MIPS/n533 ), .CK(clk), .RN(n5715), .Q(
        \i_MIPS/ALUin1[29] ), .QN(n3358) );
  DFFRX1 \i_MIPS/EX_MEM_reg[26]  ( .D(\i_MIPS/n448 ), .CK(clk), .RN(n5745), 
        .Q(n12938), .QN(n3713) );
  DFFRX2 \i_MIPS/ID_EX_reg[13]  ( .D(\i_MIPS/n558 ), .CK(clk), .RN(n5713), .Q(
        \i_MIPS/ALUin1[4] ), .QN(\i_MIPS/n367 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[31]  ( .D(\i_MIPS/n540 ), .CK(clk), .RN(n5714), .Q(
        \i_MIPS/ALUin1[22] ), .QN(\i_MIPS/n349 ) );
  DFFRX1 \I_cache/cache_reg[0][79]  ( .D(n12155), .CK(clk), .RN(n5787), .Q(
        \I_cache/cache[0][79] ), .QN(n3323) );
  DFFRX2 \i_MIPS/ID_EX_reg[40]  ( .D(\i_MIPS/n531 ), .CK(clk), .RN(n5715), .Q(
        \i_MIPS/ALU/N303 ), .QN(\i_MIPS/n340 ) );
  DFFRX1 \I_cache/cache_reg[1][99]  ( .D(n11994), .CK(clk), .RN(n5853), .Q(
        \I_cache/cache[1][99] ), .QN(n3322) );
  DFFRX2 \i_MIPS/ID_EX_reg[105]  ( .D(\i_MIPS/n518 ), .CK(clk), .RN(n5737), 
        .Q(\i_MIPS/ID_EX[105] ), .QN(\i_MIPS/n323 ) );
  DFFRX1 \D_cache/cache_reg[5][41]  ( .D(\D_cache/n1463 ), .CK(clk), .RN(n5676), .Q(\D_cache/cache[5][41] ), .QN(n2980) );
  DFFRX2 \D_cache/cache_reg[0][31]  ( .D(\D_cache/n1548 ), .CK(clk), .RN(n5703), .Q(\D_cache/cache[0][31] ), .QN(n2979) );
  DFFRX1 \D_cache/cache_reg[0][62]  ( .D(\D_cache/n1300 ), .CK(clk), .RN(n5682), .Q(\D_cache/cache[0][62] ), .QN(n2978) );
  DFFRX2 \D_cache/cache_reg[0][63]  ( .D(\D_cache/n1292 ), .CK(clk), .RN(n5681), .Q(\D_cache/cache[0][63] ), .QN(n2977) );
  DFFRX2 \D_cache/cache_reg[0][126]  ( .D(\D_cache/n788 ), .CK(clk), .RN(n5879), .Q(\D_cache/cache[0][126] ), .QN(n2976) );
  DFFRX1 \D_cache/cache_reg[0][55]  ( .D(\D_cache/n1356 ), .CK(clk), .RN(n5667), .Q(\D_cache/cache[0][55] ), .QN(n2975) );
  DFFRX2 \D_cache/cache_reg[0][46]  ( .D(\D_cache/n1428 ), .CK(clk), .RN(n5673), .Q(\D_cache/cache[0][46] ), .QN(n2974) );
  DFFRX1 \D_cache/cache_reg[0][49]  ( .D(\D_cache/n1404 ), .CK(clk), .RN(n5671), .Q(\D_cache/cache[0][49] ), .QN(n2973) );
  DFFRX1 \D_cache/cache_reg[0][23]  ( .D(\D_cache/n1612 ), .CK(clk), .RN(n5688), .Q(\D_cache/cache[0][23] ), .QN(n2971) );
  DFFRX1 \D_cache/cache_reg[0][20]  ( .D(\D_cache/n1636 ), .CK(clk), .RN(n5690), .Q(\D_cache/cache[0][20] ), .QN(n2970) );
  DFFRX2 \D_cache/cache_reg[0][112]  ( .D(\D_cache/n900 ), .CK(clk), .RN(n5868), .Q(\D_cache/cache[0][112] ), .QN(n2969) );
  DFFRX1 \D_cache/cache_reg[0][102]  ( .D(\D_cache/n980 ), .CK(clk), .RN(n5875), .Q(\D_cache/cache[0][102] ), .QN(n2968) );
  DFFRX2 \D_cache/cache_reg[0][119]  ( .D(\D_cache/n844 ), .CK(clk), .RN(n5884), .Q(\D_cache/cache[0][119] ), .QN(n2966) );
  DFFRX1 \D_cache/cache_reg[0][107]  ( .D(\D_cache/n940 ), .CK(clk), .RN(n5872), .Q(\D_cache/cache[0][107] ), .QN(n2965) );
  DFFRX1 \D_cache/cache_reg[0][121]  ( .D(\D_cache/n828 ), .CK(clk), .RN(n5882), .Q(\D_cache/cache[0][121] ), .QN(n2962) );
  DFFRX1 \D_cache/cache_reg[0][117]  ( .D(\D_cache/n860 ), .CK(clk), .RN(n5885), .Q(\D_cache/cache[0][117] ), .QN(n2961) );
  DFFRX1 \D_cache/cache_reg[2][83]  ( .D(\D_cache/n1130 ), .CK(clk), .RN(n5888), .Q(\D_cache/cache[2][83] ), .QN(n2960) );
  DFFRX2 \D_cache/cache_reg[0][44]  ( .D(\D_cache/n1444 ), .CK(clk), .RN(n5674), .Q(\D_cache/cache[0][44] ), .QN(n2959) );
  DFFRX1 \D_cache/cache_reg[0][14]  ( .D(\D_cache/n1684 ), .CK(clk), .RN(n5694), .Q(\D_cache/cache[0][14] ), .QN(n2958) );
  DFFRX1 \D_cache/cache_reg[0][13]  ( .D(\D_cache/n1692 ), .CK(clk), .RN(n5695), .Q(\D_cache/cache[0][13] ), .QN(n2957) );
  DFFRX1 \D_cache/cache_reg[0][30]  ( .D(\D_cache/n1556 ), .CK(clk), .RN(n5704), .Q(\D_cache/cache[0][30] ), .QN(n2956) );
  DFFRX1 \D_cache/cache_reg[0][45]  ( .D(\D_cache/n1436 ), .CK(clk), .RN(n5674), .Q(\D_cache/cache[0][45] ), .QN(n2955) );
  DFFRX1 \D_cache/cache_reg[2][110]  ( .D(\D_cache/n914 ), .CK(clk), .RN(n5869), .Q(\D_cache/cache[2][110] ), .QN(n2953) );
  DFFRX2 \i_MIPS/ID_EX_reg[36]  ( .D(\i_MIPS/n535 ), .CK(clk), .RN(n5715), .Q(
        \i_MIPS/ALUin1[27] ), .QN(\i_MIPS/n344 ) );
  DFFRX1 \D_cache/cache_reg[1][51]  ( .D(\D_cache/n1387 ), .CK(clk), .RN(n5669), .Q(\D_cache/cache[1][51] ), .QN(n2421) );
  DFFRX1 \D_cache/cache_reg[0][4]  ( .D(\D_cache/n1764 ), .CK(clk), .RN(n5641), 
        .Q(\D_cache/cache[0][4] ), .QN(n2420) );
  DFFRX1 \D_cache/cache_reg[0][69]  ( .D(\D_cache/n1244 ), .CK(clk), .RN(n5677), .Q(\D_cache/cache[0][69] ), .QN(n2417) );
  DFFRX1 \D_cache/cache_reg[0][122]  ( .D(\D_cache/n820 ), .CK(clk), .RN(n5882), .Q(\D_cache/cache[0][122] ), .QN(n2416) );
  DFFRX1 \D_cache/cache_reg[0][57]  ( .D(\D_cache/n1340 ), .CK(clk), .RN(n5685), .Q(\D_cache/cache[0][57] ), .QN(n2415) );
  DFFRX1 \D_cache/cache_reg[0][116]  ( .D(\D_cache/n868 ), .CK(clk), .RN(n5886), .Q(\D_cache/cache[0][116] ), .QN(n2414) );
  DFFRX1 \D_cache/cache_reg[0][83]  ( .D(\D_cache/n1132 ), .CK(clk), .RN(n5888), .Q(\D_cache/cache[0][83] ), .QN(n2413) );
  DFFRX1 \D_cache/cache_reg[0][123]  ( .D(\D_cache/n812 ), .CK(clk), .RN(n5881), .Q(\D_cache/cache[0][123] ), .QN(n2412) );
  DFFRX1 \D_cache/cache_reg[0][19]  ( .D(\D_cache/n1644 ), .CK(clk), .RN(n5691), .Q(\D_cache/cache[0][19] ), .QN(n2411) );
  DFFRX1 \D_cache/cache_reg[0][64]  ( .D(\D_cache/n1284 ), .CK(clk), .RN(n5681), .Q(\D_cache/cache[0][64] ), .QN(n2410) );
  DFFRX1 \D_cache/cache_reg[0][105]  ( .D(\D_cache/n956 ), .CK(clk), .RN(n5873), .Q(\D_cache/cache[0][105] ), .QN(n2409) );
  DFFRX1 \D_cache/cache_reg[2][119]  ( .D(\D_cache/n842 ), .CK(clk), .RN(n5883), .Q(\D_cache/cache[2][119] ), .QN(n2408) );
  DFFRX1 \D_cache/cache_reg[0][28]  ( .D(\D_cache/n1572 ), .CK(clk), .RN(n5705), .Q(\D_cache/cache[0][28] ), .QN(n2205) );
  DFFRX1 \D_cache/cache_reg[0][124]  ( .D(\D_cache/n804 ), .CK(clk), .RN(n5880), .Q(\D_cache/cache[0][124] ), .QN(n2204) );
  DFFRX2 \D_cache/cache_reg[0][108]  ( .D(\D_cache/n932 ), .CK(clk), .RN(n5871), .Q(\D_cache/cache[0][108] ), .QN(n2203) );
  DFFRX1 \I_cache/cache_reg[4][152]  ( .D(n11567), .CK(clk), .RN(n5838), .Q(
        \I_cache/cache[4][152] ), .QN(n2202) );
  DFFRX2 \i_MIPS/ID_EX_reg[11]  ( .D(\i_MIPS/n560 ), .CK(clk), .RN(n5713), .Q(
        \i_MIPS/ALUin1[2] ), .QN(\i_MIPS/n369 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[14]  ( .D(\i_MIPS/n460 ), .CK(clk), .RN(n5744), 
        .Q(n12950), .QN(n3901) );
  DFFRX2 \i_MIPS/ID_EX_reg[23]  ( .D(\i_MIPS/n548 ), .CK(clk), .RN(n5714), .Q(
        \i_MIPS/ALUin1[14] ), .QN(\i_MIPS/n357 ) );
  DFFRX1 \I_cache/cache_reg[2][22]  ( .D(n12609), .CK(clk), .RN(n5925), .Q(
        \I_cache/cache[2][22] ), .QN(n1936) );
  DFFRX1 \I_cache/cache_reg[4][22]  ( .D(n12607), .CK(clk), .RN(n5924), .Q(
        \I_cache/cache[4][22] ), .QN(n1935) );
  DFFRX1 \I_cache/cache_reg[0][22]  ( .D(n12611), .CK(clk), .RN(n5925), .Q(
        \I_cache/cache[0][22] ), .QN(n1934) );
  DFFRX1 \I_cache/cache_reg[7][154]  ( .D(n11548), .CK(clk), .RN(n5846), .Q(
        \I_cache/cache[7][154] ), .QN(n1775) );
  DFFRX2 \i_MIPS/ID_EX_reg[26]  ( .D(\i_MIPS/n545 ), .CK(clk), .RN(n5714), .Q(
        \i_MIPS/ALUin1[17] ), .QN(\i_MIPS/n354 ) );
  DFFRX2 \I_cache/cache_reg[1][79]  ( .D(n12154), .CK(clk), .RN(n5787), .Q(
        \I_cache/cache[1][79] ), .QN(n1722) );
  DFFRX2 \i_MIPS/ID_EX_reg[32]  ( .D(\i_MIPS/n539 ), .CK(clk), .RN(n5715), .Q(
        \i_MIPS/ALUin1[23] ), .QN(\i_MIPS/n348 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[30]  ( .D(\i_MIPS/n541 ), .CK(clk), .RN(n5714), .Q(
        \i_MIPS/ALUin1[21] ), .QN(\i_MIPS/n350 ) );
  DFFRX1 \D_cache/cache_reg[0][51]  ( .D(\D_cache/n1388 ), .CK(clk), .RN(n5669), .Q(\D_cache/cache[0][51] ), .QN(n851) );
  DFFRX2 \i_MIPS/ID_EX_reg[39]  ( .D(\i_MIPS/n532 ), .CK(clk), .RN(n5715), .Q(
        \i_MIPS/ALUin1[30] ), .QN(\i_MIPS/n341 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[35]  ( .D(\i_MIPS/n536 ), .CK(clk), .RN(n5715), .Q(
        \i_MIPS/ALUin1[26] ), .QN(\i_MIPS/n345 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[8]  ( .D(\i_MIPS/n466 ), .CK(clk), .RN(n5743), .Q(
        n12954), .QN(n437) );
  DFFRX4 \i_MIPS/IF_ID_reg[49]  ( .D(\i_MIPS/N75 ), .CK(clk), .RN(n5738), .Q(
        \i_MIPS/IR_ID[17] ), .QN(\i_MIPS/n314 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[21]  ( .D(\i_MIPS/n453 ), .CK(clk), .RN(n5745), 
        .Q(n12943), .QN(n4628) );
  DFFRX2 \i_MIPS/ID_EX_reg[24]  ( .D(\i_MIPS/n547 ), .CK(clk), .RN(n5714), .Q(
        \i_MIPS/ALUin1[15] ), .QN(\i_MIPS/n356 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[21]  ( .D(\i_MIPS/n550 ), .CK(clk), .RN(n5714), .Q(
        \i_MIPS/ALUin1[12] ), .QN(\i_MIPS/n359 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[14]  ( .D(\i_MIPS/n557 ), .CK(clk), .RN(n5713), .Q(
        \i_MIPS/ALUin1[5] ), .QN(\i_MIPS/n366 ) );
  DFFRHQX4 \i_MIPS/PC/PC_o_reg[2]  ( .D(\i_MIPS/PC/n36 ), .CK(clk), .RN(n5712), 
        .Q(n4301) );
  DFFRX2 \i_MIPS/ID_EX_reg[27]  ( .D(\i_MIPS/n544 ), .CK(clk), .RN(n5714), .Q(
        \i_MIPS/ALUin1[18] ), .QN(\i_MIPS/n353 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[31]  ( .D(\i_MIPS/n443 ), .CK(clk), .RN(n5745), 
        .Q(n12933), .QN(n4293) );
  DFFRX1 \i_MIPS/EX_MEM_reg[33]  ( .D(\i_MIPS/n441 ), .CK(clk), .RN(n5746), 
        .Q(n12931), .QN(n4291) );
  DFFRX1 \i_MIPS/EX_MEM_reg[12]  ( .D(\i_MIPS/n462 ), .CK(clk), .RN(n5744), 
        .Q(n12952), .QN(n4289) );
  DFFRX1 \i_MIPS/EX_MEM_reg[56]  ( .D(\i_MIPS/n398 ), .CK(clk), .RN(n5729), 
        .Q(n12968), .QN(\i_MIPS/n270 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[39]  ( .D(\i_MIPS/n432 ), .CK(clk), .RN(n5731), 
        .Q(n12985), .QN(\i_MIPS/n304 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[63]  ( .D(\i_MIPS/n384 ), .CK(clk), .RN(n5730), 
        .Q(n12961), .QN(\i_MIPS/n256 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[65]  ( .D(\i_MIPS/n380 ), .CK(clk), .RN(n5731), 
        .Q(n12959), .QN(\i_MIPS/n252 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[37]  ( .D(\i_MIPS/n436 ), .CK(clk), .RN(n5746), 
        .Q(n12987), .QN(\i_MIPS/n308 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[38]  ( .D(\i_MIPS/n434 ), .CK(clk), .RN(n5746), 
        .Q(n12986), .QN(\i_MIPS/n306 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[40]  ( .D(\i_MIPS/n430 ), .CK(clk), .RN(n5726), 
        .Q(n12984), .QN(\i_MIPS/n302 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[41]  ( .D(\i_MIPS/n428 ), .CK(clk), .RN(n5727), 
        .Q(n12983), .QN(\i_MIPS/n300 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[42]  ( .D(\i_MIPS/n426 ), .CK(clk), .RN(n5727), 
        .Q(n12982), .QN(\i_MIPS/n298 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[43]  ( .D(\i_MIPS/n424 ), .CK(clk), .RN(n5727), 
        .Q(n12981), .QN(\i_MIPS/n296 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[44]  ( .D(\i_MIPS/n422 ), .CK(clk), .RN(n5727), 
        .Q(n12980), .QN(\i_MIPS/n294 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[45]  ( .D(\i_MIPS/n420 ), .CK(clk), .RN(n5727), 
        .Q(n12979), .QN(\i_MIPS/n292 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[46]  ( .D(\i_MIPS/n418 ), .CK(clk), .RN(n5727), 
        .Q(n12978), .QN(\i_MIPS/n290 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[47]  ( .D(\i_MIPS/n416 ), .CK(clk), .RN(n5728), 
        .Q(n12977), .QN(\i_MIPS/n288 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[48]  ( .D(\i_MIPS/n414 ), .CK(clk), .RN(n5728), 
        .Q(n12976), .QN(\i_MIPS/n286 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[49]  ( .D(\i_MIPS/n412 ), .CK(clk), .RN(n5728), 
        .Q(n12975), .QN(\i_MIPS/n284 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[50]  ( .D(\i_MIPS/n410 ), .CK(clk), .RN(n5728), 
        .Q(n12974), .QN(\i_MIPS/n282 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[51]  ( .D(\i_MIPS/n408 ), .CK(clk), .RN(n5728), 
        .Q(n12973), .QN(\i_MIPS/n280 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[52]  ( .D(\i_MIPS/n406 ), .CK(clk), .RN(n5728), 
        .Q(n12972), .QN(\i_MIPS/n278 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[53]  ( .D(\i_MIPS/n404 ), .CK(clk), .RN(n5729), 
        .Q(n12971), .QN(\i_MIPS/n276 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[54]  ( .D(\i_MIPS/n402 ), .CK(clk), .RN(n5729), 
        .Q(n12970), .QN(\i_MIPS/n274 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[55]  ( .D(\i_MIPS/n400 ), .CK(clk), .RN(n5729), 
        .Q(n12969), .QN(\i_MIPS/n272 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[57]  ( .D(\i_MIPS/n396 ), .CK(clk), .RN(n5729), 
        .Q(n12967), .QN(\i_MIPS/n268 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[58]  ( .D(\i_MIPS/n394 ), .CK(clk), .RN(n5729), 
        .Q(n12966), .QN(\i_MIPS/n266 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[59]  ( .D(\i_MIPS/n392 ), .CK(clk), .RN(n5730), 
        .Q(n12965), .QN(\i_MIPS/n264 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[60]  ( .D(\i_MIPS/n390 ), .CK(clk), .RN(n5730), 
        .Q(n12964), .QN(\i_MIPS/n262 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[61]  ( .D(\i_MIPS/n388 ), .CK(clk), .RN(n5730), 
        .Q(n12963), .QN(\i_MIPS/n260 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[62]  ( .D(\i_MIPS/n386 ), .CK(clk), .RN(n5730), 
        .Q(n12962), .QN(\i_MIPS/n258 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[64]  ( .D(\i_MIPS/n382 ), .CK(clk), .RN(n5730), 
        .Q(n12960), .QN(\i_MIPS/n254 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[66]  ( .D(\i_MIPS/n378 ), .CK(clk), .RN(n5731), 
        .Q(n12958), .QN(\i_MIPS/n250 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[67]  ( .D(\i_MIPS/n376 ), .CK(clk), .RN(n5731), 
        .Q(n12957), .QN(\i_MIPS/n248 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[68]  ( .D(\i_MIPS/n374 ), .CK(clk), .RN(n5731), 
        .Q(n12956), .QN(\i_MIPS/n246 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[4]  ( .D(\i_MIPS/n479 ), .CK(clk), .RN(n5742), .Q(
        n12988), .QN(\i_MIPS/n310 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[22]  ( .D(\i_MIPS/n549 ), .CK(clk), .RN(n5714), .Q(
        \i_MIPS/ALUin1[13] ), .QN(\i_MIPS/n358 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[10]  ( .D(\i_MIPS/n561 ), .CK(clk), .RN(n5713), .Q(
        \i_MIPS/ALUin1[1] ), .QN(\i_MIPS/n370 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[12]  ( .D(\i_MIPS/n559 ), .CK(clk), .RN(n5713), .Q(
        \i_MIPS/ALUin1[3] ), .QN(\i_MIPS/n368 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[85]  ( .D(\i_MIPS/n500 ), .CK(clk), .RN(n5740), .Q(
        \i_MIPS/ID_EX[85] ), .QN(n4539) );
  DFFRX2 \i_MIPS/ID_EX_reg[29]  ( .D(\i_MIPS/n542 ), .CK(clk), .RN(n5714), .Q(
        \i_MIPS/ALUin1[20] ), .QN(\i_MIPS/n351 ) );
  DFFRX2 \D_cache/cache_reg[0][114]  ( .D(\D_cache/n884 ), .CK(clk), .RN(n5867), .Q(\D_cache/cache[0][114] ), .QN(n2952) );
  DFFRX2 \D_cache/cache_reg[0][118]  ( .D(\D_cache/n852 ), .CK(clk), .RN(n5884), .Q(\D_cache/cache[0][118] ), .QN(n2647) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[11]  ( .D(\i_MIPS/PC/n45 ), .CK(clk), .RN(n5711), 
        .Q(ICACHE_addr[9]), .QN(\i_MIPS/PC/n13 ) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[25]  ( .D(\i_MIPS/PC/n59 ), .CK(clk), .RN(n5710), 
        .Q(ICACHE_addr[23]), .QN(\i_MIPS/PC/n27 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[100]  ( .D(\i_MIPS/n485 ), .CK(clk), .RN(n5742), 
        .Q(\i_MIPS/ID_EX[100] ) );
  DFFRX1 \I_cache/cache_reg[0][99]  ( .D(n11995), .CK(clk), .RN(n5853), .Q(
        \I_cache/cache[0][99] ), .QN(n1721) );
  DFFRX1 \i_MIPS/ID_EX_reg[96]  ( .D(\i_MIPS/n489 ), .CK(clk), .RN(n5741), .Q(
        \i_MIPS/ID_EX[96] ) );
  DFFRX2 \i_MIPS/ID_EX_reg[49]  ( .D(\i_MIPS/n421 ), .CK(clk), .RN(n5727), .Q(
        \i_MIPS/ID_EX[49] ), .QN(\i_MIPS/n293 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[83]  ( .D(\i_MIPS/N109 ), .CK(clk), .RN(n5735), .Q(
        \i_MIPS/IF_ID[83] ), .QN(\i_MIPS/n169 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[95]  ( .D(\i_MIPS/N121 ), .CK(clk), .RN(n5746), .Q(
        \i_MIPS/IF_ID[95] ), .QN(\i_MIPS/n181 ) );
  DFFRX2 \D_cache/cache_reg[0][32]  ( .D(\D_cache/n1540 ), .CK(clk), .RN(n5702), .Q(\D_cache/cache[0][32] ), .QN(n2964) );
  DFFRX2 \i_MIPS/IF_ID_reg[89]  ( .D(\i_MIPS/N115 ), .CK(clk), .RN(n5736), .Q(
        \i_MIPS/IF_ID[89] ), .QN(\i_MIPS/n175 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[66]  ( .D(\i_MIPS/N92 ), .CK(clk), .RN(n5734), .Q(
        \i_MIPS/IF_ID[66] ), .QN(\i_MIPS/n238 ) );
  DFFRX1 \D_cache/cache_reg[3][0]  ( .D(\D_cache/n1792 ), .CK(clk), .RN(n5643), 
        .Q(\D_cache/cache[3][0] ), .QN(n1427) );
  DFFRHQX4 \i_MIPS/ID_EX_reg[74]  ( .D(\i_MIPS/n511 ), .CK(clk), .RN(n5739), 
        .Q(n3812) );
  DFFRX1 \D_cache/cache_reg[1][145]  ( .D(\D_cache/n635 ), .CK(clk), .RN(n5926), .Q(\D_cache/cache[1][145] ) );
  DFFRX1 \i_MIPS/IF_ID_reg[61]  ( .D(\i_MIPS/N87 ), .CK(clk), .RN(n5716), .Q(
        \i_MIPS/IR_ID[29] ), .QN(\i_MIPS/n328 ) );
  DFFRHQX4 \i_MIPS/ID_EX_reg[6]  ( .D(\i_MIPS/n472 ), .CK(clk), .RN(n5743), 
        .Q(n3704) );
  DFFRX2 \i_MIPS/ID_EX_reg[84]  ( .D(\i_MIPS/n501 ), .CK(clk), .RN(n5740), .Q(
        \i_MIPS/ID_EX[84] ), .QN(n4537) );
  DFFRHQX4 \i_MIPS/ID_EX_reg[76]  ( .D(\i_MIPS/n509 ), .CK(clk), .RN(n5740), 
        .Q(n3696) );
  DFFRX1 \i_MIPS/ID_EX_reg[99]  ( .D(\i_MIPS/n486 ), .CK(clk), .RN(n5742), .Q(
        \i_MIPS/ID_EX[99] ) );
  DFFRX1 \i_MIPS/ID_EX_reg[101]  ( .D(\i_MIPS/n484 ), .CK(clk), .RN(n5742), 
        .Q(\i_MIPS/ID_EX[101] ) );
  DFFRX1 \i_MIPS/IF_ID_reg[64]  ( .D(\i_MIPS/N90 ), .CK(clk), .RN(n5742), .Q(
        \i_MIPS/IF_ID[64] ), .QN(\i_MIPS/n236 ) );
  DFFRX1 \D_cache/cache_reg[0][58]  ( .D(\D_cache/n1332 ), .CK(clk), .RN(n5685), .Q(\D_cache/cache[0][58] ), .QN(n2972) );
  DFFRX1 \D_cache/cache_reg[0][87]  ( .D(\D_cache/n1100 ), .CK(clk), .RN(n5905), .Q(\D_cache/cache[0][87] ), .QN(n2954) );
  DFFRX1 \D_cache/cache_reg[0][59]  ( .D(\D_cache/n1324 ), .CK(clk), .RN(n5684), .Q(\D_cache/cache[0][59] ), .QN(n2418) );
  DFFRX1 \i_MIPS/ID_EX_reg[59]  ( .D(\i_MIPS/n401 ), .CK(clk), .RN(n5729), .Q(
        n3595), .QN(\i_MIPS/n273 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[56]  ( .D(\i_MIPS/n407 ), .CK(clk), .RN(n5728), .Q(
        n4378), .QN(\i_MIPS/n279 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[58]  ( .D(\i_MIPS/n403 ), .CK(clk), .RN(n5729), .Q(
        n3594), .QN(\i_MIPS/n275 ) );
  DFFRX4 \i_MIPS/PC/PC_o_reg[9]  ( .D(\i_MIPS/PC/n43 ), .CK(clk), .RN(n5711), 
        .Q(ICACHE_addr[7]), .QN(\i_MIPS/PC/n11 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[55]  ( .D(\i_MIPS/n409 ), .CK(clk), .RN(n5728), .Q(
        n3599), .QN(\i_MIPS/n281 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[86]  ( .D(\i_MIPS/n499 ), .CK(clk), .RN(n5740), .Q(
        \i_MIPS/ID_EX[86] ), .QN(n4538) );
  DFFRX2 \i_MIPS/ID_EX_reg[54]  ( .D(\i_MIPS/n411 ), .CK(clk), .RN(n5728), .Q(
        n3607), .QN(\i_MIPS/n283 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[46]  ( .D(\i_MIPS/n427 ), .CK(clk), .RN(n5727), .Q(
        n3603), .QN(\i_MIPS/n299 ) );
  DFFRHQX4 \i_MIPS/PC/PC_o_reg[8]  ( .D(\i_MIPS/PC/n42 ), .CK(clk), .RN(n5711), 
        .Q(n3781) );
  DFFRX4 \i_MIPS/ID_EX_reg[47]  ( .D(\i_MIPS/n425 ), .CK(clk), .RN(n5727), .Q(
        n3612), .QN(\i_MIPS/n297 ) );
  DFFRX4 \i_MIPS/ID_EX_reg[89]  ( .D(\i_MIPS/n496 ), .CK(clk), .RN(n5741), .Q(
        \i_MIPS/ID_EX[89] ), .QN(n4493) );
  DFFRX4 \i_MIPS/ID_EX_reg[57]  ( .D(\i_MIPS/n405 ), .CK(clk), .RN(n5729), .Q(
        n3600), .QN(\i_MIPS/n277 ) );
  DFFRX4 \i_MIPS/ID_EX_reg[41]  ( .D(\i_MIPS/n437 ), .CK(clk), .RN(n5746), 
        .QN(\i_MIPS/n309 ) );
  DFFRX2 \D_cache/cache_reg[1][21]  ( .D(\D_cache/n1627 ), .CK(clk), .RN(n5689), .Q(\D_cache/cache[1][21] ), .QN(n1075) );
  DFFRX2 \i_MIPS/ID_EX_reg[115]  ( .D(\i_MIPS/n517 ), .CK(clk), .RN(n5737), 
        .Q(\i_MIPS/ID_EX[115] ), .QN(\i_MIPS/n321 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[113]  ( .D(\i_MIPS/n515 ), .CK(clk), .RN(n5738), 
        .QN(\i_MIPS/n317 ) );
  DFFRHQX8 \i_MIPS/PC/PC_o_reg[6]  ( .D(\i_MIPS/PC/n40 ), .CK(clk), .RN(n5711), 
        .Q(n3785) );
  DFFRX4 \I_cache/cache_reg[1][92]  ( .D(n12050), .CK(clk), .RN(n5798), .Q(
        \I_cache/cache[1][92] ), .QN(n2695) );
  DFFRX2 \I_cache/cache_reg[0][94]  ( .D(n12035), .CK(clk), .RN(n5797), .Q(
        \I_cache/cache[0][94] ), .QN(n1528) );
  DFFRX2 \I_cache/cache_reg[0][126]  ( .D(n11779), .CK(clk), .RN(n5835), .Q(
        \I_cache/cache[0][126] ), .QN(n1524) );
  DFFRX4 \I_cache/cache_reg[0][29]  ( .D(n12555), .CK(clk), .RN(n5920), .Q(
        \I_cache/cache[0][29] ), .QN(n1515) );
  DFFRX4 \I_cache/cache_reg[1][94]  ( .D(n12034), .CK(clk), .RN(n5797), .Q(
        \I_cache/cache[1][94] ), .QN(n3108) );
  DFFRX4 \I_cache/cache_reg[7][126]  ( .D(n11772), .CK(clk), .RN(n5835), .Q(
        \I_cache/cache[7][126] ), .QN(n3105) );
  DFFRX2 \i_MIPS/PHT_2/current_state_1_reg[0]  ( .D(n11508), .CK(clk), .RN(
        n5712), .Q(n3606), .QN(\i_MIPS/PHT_2/n8 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[37]  ( .D(\i_MIPS/n534 ), .CK(clk), .RN(n5715), .Q(
        \i_MIPS/ALUin1[28] ), .QN(\i_MIPS/n343 ) );
  DFFRX4 \i_MIPS/ID_EX_reg[43]  ( .D(\i_MIPS/n433 ), .CK(clk), .RN(n5746), .Q(
        \i_MIPS/ID_EX[43] ), .QN(\i_MIPS/n305 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[61]  ( .D(\i_MIPS/n397 ), .CK(clk), .RN(n5729), .Q(
        n3602), .QN(\i_MIPS/n269 ) );
  NAND3X8 U2 ( .A(n7219), .B(n7891), .C(n7218), .Y(n7220) );
  INVX6 U3 ( .A(n11173), .Y(n11163) );
  OAI221XL U4 ( .A0(net103954), .A1(net111624), .B0(net103955), .B1(net111636), 
        .C0(net103956), .Y(n2) );
  CLKMX2X2 U5 ( .A(n7462), .B(n7461), .S0(net107812), .Y(net103954) );
  INVX12 U6 ( .A(net112676), .Y(net97445) );
  INVX3 U7 ( .A(net98063), .Y(net103955) );
  AND2X6 U8 ( .A(n3425), .B(net98755), .Y(n3693) );
  NAND2X6 U9 ( .A(net100400), .B(n324), .Y(n4146) );
  NAND3BX4 U10 ( .AN(n8757), .B(n8758), .C(net112294), .Y(n8762) );
  INVX1 U11 ( .A(n8758), .Y(n8759) );
  NAND4X4 U12 ( .A(n8735), .B(n8734), .C(n4658), .D(n8733), .Y(n8743) );
  OA22X1 U13 ( .A0(n4969), .A1(n714), .B0(n5019), .B1(n2282), .Y(n9507) );
  OA22X1 U14 ( .A0(n4969), .A1(n2152), .B0(n5014), .B1(n573), .Y(n8991) );
  OA22X1 U15 ( .A0(n4969), .A1(n708), .B0(n5014), .B1(n2276), .Y(n9080) );
  OA22X1 U16 ( .A0(n4969), .A1(n2097), .B0(n5014), .B1(n510), .Y(n8983) );
  BUFX2 U17 ( .A(n4994), .Y(n4969) );
  INVX3 U18 ( .A(net103070), .Y(n3) );
  INVX3 U19 ( .A(n3), .Y(n4) );
  AO21XL U20 ( .A0(net102429), .A1(net102430), .B0(net102431), .Y(n8340) );
  NAND2X6 U21 ( .A(net102430), .B(n8360), .Y(n6756) );
  NAND2X2 U22 ( .A(\i_MIPS/ALUin1[2] ), .B(net105677), .Y(net105034) );
  CLKMX2X2 U23 ( .A(n8956), .B(n6492), .S0(net107798), .Y(n9460) );
  NAND2X1 U24 ( .A(n9328), .B(n6493), .Y(n6499) );
  CLKBUFX8 U25 ( .A(n5533), .Y(n5530) );
  BUFX16 U26 ( .A(n9986), .Y(n4838) );
  INVX3 U27 ( .A(n3899), .Y(n9355) );
  NAND4X2 U28 ( .A(n6035), .B(n6034), .C(n6033), .D(n6032), .Y(n11337) );
  OA22X2 U29 ( .A0(n5101), .A1(n1251), .B0(n5061), .B1(n2793), .Y(n6035) );
  AND4X8 U30 ( .A(n9359), .B(n9360), .C(n9358), .D(n9357), .Y(n3412) );
  NOR3X6 U31 ( .A(n4309), .B(n4310), .C(net100583), .Y(n7241) );
  BUFX6 U32 ( .A(net97815), .Y(n5) );
  MX2X4 U33 ( .A(n7981), .B(net100585), .S0(n6538), .Y(n7970) );
  CLKINVX6 U34 ( .A(n6538), .Y(n7969) );
  NAND4X2 U35 ( .A(n6291), .B(n6290), .C(n6289), .D(n6288), .Y(n9566) );
  NAND2BX2 U36 ( .AN(n5429), .B(n11247), .Y(n6288) );
  INVX16 U37 ( .A(net102393), .Y(net101906) );
  BUFX20 U38 ( .A(n4891), .Y(n4928) );
  AND2X1 U39 ( .A(n7683), .B(n7409), .Y(n3667) );
  AOI2BB2X1 U40 ( .B0(net111960), .B1(n8978), .A0N(n3773), .A1N(n3721), .Y(n6)
         );
  INVXL U41 ( .A(n7981), .Y(n7983) );
  OA22XL U42 ( .A0(n4920), .A1(n778), .B0(n4949), .B1(n2340), .Y(n7426) );
  OA22XL U43 ( .A0(n4920), .A1(n2290), .B0(n4949), .B1(n721), .Y(n7438) );
  OA22XL U44 ( .A0(n4920), .A1(n1223), .B0(n4949), .B1(n2760), .Y(n7353) );
  OA22XL U45 ( .A0(n4920), .A1(n1224), .B0(n4949), .B1(n2761), .Y(n7357) );
  OA22X1 U46 ( .A0(n4920), .A1(n2677), .B0(n4949), .B1(n1120), .Y(n7430) );
  BUFX4 U47 ( .A(n9987), .Y(n4890) );
  OA22X1 U48 ( .A0(n5398), .A1(n1714), .B0(n5331), .B1(n3312), .Y(n6127) );
  INVX6 U49 ( .A(net97817), .Y(net104583) );
  BUFX8 U50 ( .A(net98080), .Y(net112999) );
  AND4X6 U51 ( .A(n8566), .B(n8565), .C(n8564), .D(n8563), .Y(n3405) );
  NAND4X2 U52 ( .A(n8963), .B(n8962), .C(n4658), .D(n8961), .Y(n8973) );
  CLKMX2X2 U53 ( .A(net112438), .B(net100573), .S0(n8955), .Y(n8963) );
  INVX6 U54 ( .A(net133688), .Y(net101402) );
  CLKBUFX3 U55 ( .A(n3820), .Y(n7) );
  OR2X8 U56 ( .A(n6312), .B(n6311), .Y(n8) );
  OR2X8 U57 ( .A(n6312), .B(n6311), .Y(n9) );
  INVX16 U58 ( .A(n2017), .Y(n4246) );
  OAI221X2 U59 ( .A0(net103954), .A1(net111624), .B0(net103955), .B1(net111636), .C0(net103956), .Y(net98061) );
  NAND2BX1 U60 ( .AN(n5429), .B(n11246), .Y(n6292) );
  AO22X4 U61 ( .A0(mem_rdata_I[60]), .A1(n5542), .B0(n249), .B1(n11246), .Y(
        n6176) );
  NAND4X2 U62 ( .A(n6175), .B(n6174), .C(n6173), .D(n6172), .Y(n11246) );
  INVX1 U63 ( .A(n8), .Y(n9980) );
  AOI22X1 U64 ( .A0(n7686), .A1(net112292), .B0(net111996), .B1(n3730), .Y(
        n7716) );
  INVX3 U65 ( .A(n7691), .Y(n3730) );
  OR2X8 U66 ( .A(net103417), .B(net111636), .Y(n3651) );
  OR2X4 U67 ( .A(net103416), .B(net111624), .Y(n3650) );
  OAI221X1 U68 ( .A0(net112368), .A1(\i_MIPS/n364 ), .B0(net112350), .B1(
        \i_MIPS/n363 ), .C0(n6486), .Y(n10) );
  CLKXOR2X2 U69 ( .A(n10175), .B(n3781), .Y(n10373) );
  NAND2X6 U70 ( .A(n10370), .B(n10368), .Y(n10228) );
  AOI222X1 U71 ( .A0(n5510), .A1(n11407), .B0(mem_rdata_D[57]), .B1(n234), 
        .C0(n12962), .C1(n5506), .Y(n10501) );
  CLKAND2X3 U72 ( .A(n4199), .B(n4200), .Y(n3337) );
  NAND2X2 U73 ( .A(n10664), .B(n4201), .Y(n4202) );
  NAND2X2 U74 ( .A(n10518), .B(n4237), .Y(n4238) );
  CLKAND2X3 U75 ( .A(n7703), .B(net100585), .Y(n4149) );
  XOR2X1 U76 ( .A(n6605), .B(\i_MIPS/IR_ID[21] ), .Y(n6448) );
  NAND2X2 U77 ( .A(net100682), .B(n6453), .Y(n6455) );
  NAND4X6 U78 ( .A(n6452), .B(n6451), .C(n6608), .D(n6450), .Y(net100682) );
  BUFX6 U79 ( .A(n5268), .Y(n5264) );
  BUFX4 U80 ( .A(n4885), .Y(n4869) );
  OA22X1 U81 ( .A0(n4823), .A1(n2117), .B0(n4869), .B1(n530), .Y(n8019) );
  OA22X1 U82 ( .A0(n4823), .A1(n2118), .B0(n4869), .B1(n531), .Y(n8015) );
  OA22XL U83 ( .A0(n4823), .A1(n2119), .B0(n4869), .B1(n532), .Y(n7945) );
  OA22X1 U84 ( .A0(n4823), .A1(n2120), .B0(n4869), .B1(n533), .Y(n8023) );
  OA22X1 U85 ( .A0(n4823), .A1(n2116), .B0(n4869), .B1(n529), .Y(n8011) );
  OA22X1 U86 ( .A0(n4824), .A1(n749), .B0(n4869), .B1(n2310), .Y(n7847) );
  OA22X1 U87 ( .A0(n4824), .A1(n737), .B0(n4869), .B1(n2296), .Y(n7843) );
  INVX8 U88 ( .A(n5622), .Y(n4163) );
  INVX6 U89 ( .A(n6756), .Y(n6501) );
  OA22X1 U90 ( .A0(n4827), .A1(n736), .B0(n4872), .B1(n2295), .Y(n7435) );
  OA22X1 U91 ( .A0(n4827), .A1(n748), .B0(n4872), .B1(n2309), .Y(n7427) );
  OA22X1 U92 ( .A0(n4827), .A1(n690), .B0(n4872), .B1(n2259), .Y(n7579) );
  OA22X1 U93 ( .A0(n4827), .A1(n807), .B0(n4872), .B1(n2370), .Y(n7439) );
  BUFX4 U94 ( .A(n4883), .Y(n4872) );
  INVX4 U95 ( .A(net97736), .Y(net103719) );
  MX2X6 U96 ( .A(n7813), .B(n7812), .S0(net107798), .Y(n8655) );
  NAND4X8 U97 ( .A(n7832), .B(n7834), .C(n7833), .D(n7835), .Y(net97995) );
  MX2X8 U98 ( .A(\i_MIPS/n301 ), .B(net127933), .S0(n5623), .Y(n6542) );
  NAND2X6 U99 ( .A(n3683), .B(n4417), .Y(n7159) );
  XNOR2X4 U100 ( .A(ICACHE_addr[14]), .B(n11329), .Y(n6062) );
  NAND4X2 U101 ( .A(n6063), .B(n6062), .C(n6061), .D(n6060), .Y(n6075) );
  CLKINVX1 U102 ( .A(net98495), .Y(net98501) );
  NAND4X2 U103 ( .A(net129200), .B(net100415), .C(net100416), .D(net100417), 
        .Y(n11) );
  AND4X8 U104 ( .A(n3956), .B(n3957), .C(n3955), .D(n3958), .Y(net100415) );
  INVX4 U105 ( .A(n9488), .Y(n9148) );
  OAI211X4 U106 ( .A0(n9143), .A1(n9142), .B0(n9262), .C0(n9141), .Y(n9488) );
  OR2X6 U107 ( .A(n3901), .B(n11485), .Y(n4185) );
  AO22XL U108 ( .A0(n5528), .A1(DCACHE_addr[7]), .B0(n5527), .B1(n11485), .Y(
        n11036) );
  NAND4X8 U109 ( .A(n3799), .B(n3800), .C(n6397), .D(n6398), .Y(n11485) );
  NOR4X6 U110 ( .A(n6404), .B(n6403), .C(n6401), .D(n6402), .Y(n6427) );
  INVXL U111 ( .A(n7825), .Y(n12) );
  CLKINVX1 U112 ( .A(n9158), .Y(n7825) );
  INVX3 U113 ( .A(n8163), .Y(n7701) );
  CLKINVX1 U114 ( .A(n10645), .Y(n10635) );
  BUFX2 U115 ( .A(n4768), .Y(n4755) );
  BUFX8 U116 ( .A(n4767), .Y(n4768) );
  INVX6 U117 ( .A(n10502), .Y(n8825) );
  NAND2X4 U118 ( .A(n3419), .B(n10519), .Y(n8827) );
  BUFX4 U119 ( .A(n5395), .Y(n5388) );
  NAND2BX2 U120 ( .AN(n4247), .B(n11284), .Y(n9949) );
  NAND4X4 U121 ( .A(n6126), .B(n6125), .C(n6124), .D(n6123), .Y(n11284) );
  OAI221X2 U122 ( .A0(net112366), .A1(\i_MIPS/n350 ), .B0(net112348), .B1(
        \i_MIPS/n351 ), .C0(n6921), .Y(n6976) );
  OA22X1 U123 ( .A0(n5382), .A1(n1706), .B0(n5345), .B1(n3302), .Y(n10017) );
  NAND2BX2 U124 ( .AN(n4247), .B(n11291), .Y(n10039) );
  AO21X2 U125 ( .A0(n6704), .A1(n6705), .B0(net112306), .Y(n6716) );
  NAND2X6 U126 ( .A(n4216), .B(n8165), .Y(n6704) );
  NOR2X8 U127 ( .A(n9550), .B(n9551), .Y(net100417) );
  BUFX12 U128 ( .A(n10994), .Y(n5499) );
  OA22X2 U129 ( .A0(n3713), .A1(n3804), .B0(n4649), .B1(n3769), .Y(n3712) );
  INVX16 U130 ( .A(n3715), .Y(mem_addr_D[22]) );
  INVX16 U131 ( .A(n3732), .Y(mem_addr_D[23]) );
  INVX6 U132 ( .A(n7686), .Y(n7690) );
  AND4X8 U133 ( .A(n3946), .B(n3945), .C(n3948), .D(n3947), .Y(net102783) );
  BUFX20 U134 ( .A(n5508), .Y(n5511) );
  AND2X4 U135 ( .A(n4205), .B(n4206), .Y(n3331) );
  NAND2X1 U136 ( .A(\i_MIPS/ALUin1[24] ), .B(n6567), .Y(n8236) );
  CLKINVX1 U137 ( .A(n6567), .Y(n6564) );
  NAND2X1 U138 ( .A(n6567), .B(\i_MIPS/n347 ), .Y(n8253) );
  CLKMX2X8 U139 ( .A(\i_MIPS/n261 ), .B(n4489), .S0(n4323), .Y(n6567) );
  AND2X4 U140 ( .A(n4233), .B(n4234), .Y(n3327) );
  AND2X4 U141 ( .A(n4242), .B(n4243), .Y(n3332) );
  INVX4 U142 ( .A(net103076), .Y(net103079) );
  BUFX4 U143 ( .A(n5353), .Y(n5332) );
  NAND2X1 U144 ( .A(n9330), .B(n9329), .Y(n9354) );
  OAI211X1 U145 ( .A0(n3638), .A1(n7800), .B0(n9268), .C0(n9266), .Y(n7537) );
  INVX4 U146 ( .A(n6525), .Y(n3644) );
  INVXL U147 ( .A(net103955), .Y(n13) );
  AND4X8 U148 ( .A(n3749), .B(n3748), .C(n3750), .D(n3751), .Y(net100416) );
  BUFX2 U149 ( .A(n9986), .Y(n4844) );
  OA22X4 U150 ( .A0(n5284), .A1(n2168), .B0(n5239), .B1(n594), .Y(n6017) );
  BUFX8 U151 ( .A(n10651), .Y(n14) );
  CLKBUFX6 U152 ( .A(n5176), .Y(n5155) );
  NAND4X6 U153 ( .A(n6295), .B(n6294), .C(n6293), .D(n6292), .Y(n10347) );
  NAND2BX1 U154 ( .AN(n5428), .B(n11214), .Y(n6293) );
  OA22X2 U155 ( .A0(n5285), .A1(n742), .B0(n5238), .B1(n2303), .Y(n6033) );
  OA22X1 U156 ( .A0(n5210), .A1(n1616), .B0(n5167), .B1(n3193), .Y(n9936) );
  OAI222X1 U157 ( .A0(n3782), .A1(net108688), .B0(n3637), .B1(n10373), .C0(
        n4431), .C1(net108704), .Y(n10381) );
  BUFX12 U158 ( .A(n4384), .Y(n5502) );
  NAND4X2 U159 ( .A(n6195), .B(n6194), .C(n6193), .D(n6192), .Y(n11249) );
  NAND2BX2 U160 ( .AN(n5428), .B(n11217), .Y(n6281) );
  BUFX2 U161 ( .A(n5308), .Y(n5286) );
  MX2X1 U162 ( .A(\I_cache/cache[7][126] ), .B(n6211), .S0(n5317), .Y(n11772)
         );
  CLKMX2X3 U163 ( .A(\I_cache/cache[2][126] ), .B(n6211), .S0(n5184), .Y(
        n11777) );
  MX2X1 U164 ( .A(\I_cache/cache[1][94] ), .B(n6216), .S0(n5051), .Y(n12034)
         );
  CLKMX2X3 U165 ( .A(\I_cache/cache[6][94] ), .B(n6216), .S0(n5362), .Y(n12029) );
  MX2X1 U166 ( .A(\I_cache/cache[0][29] ), .B(n6221), .S0(n5094), .Y(n12555)
         );
  CLKMX2X3 U167 ( .A(\I_cache/cache[7][29] ), .B(n6221), .S0(n5317), .Y(n12548) );
  MX2X1 U168 ( .A(\I_cache/cache[1][92] ), .B(n6176), .S0(n5053), .Y(n12050)
         );
  CLKMX2X3 U169 ( .A(\I_cache/cache[6][92] ), .B(n6176), .S0(n5364), .Y(n12045) );
  AND3X8 U170 ( .A(\i_MIPS/IF_ID[64] ), .B(net97574), .C(net97444), .Y(n15) );
  OAI221XL U171 ( .A0(n9461), .A1(n8261), .B0(n9336), .B1(n8260), .C0(n4658), 
        .Y(n8090) );
  AND2X1 U172 ( .A(n4656), .B(n11308), .Y(n12824) );
  OAI2BB2X1 U173 ( .B0(net108192), .B1(\i_MIPS/n322 ), .A0N(n5545), .A1N(n9565), .Y(\i_MIPS/N84 ) );
  NAND4X2 U174 ( .A(n6279), .B(n6278), .C(n6277), .D(n6276), .Y(n9565) );
  CLKINVX4 U175 ( .A(n10416), .Y(n10417) );
  NAND2X4 U176 ( .A(n3418), .B(net98550), .Y(n4095) );
  NAND4X8 U177 ( .A(n10135), .B(n10134), .C(n10133), .D(n10132), .Y(n10236) );
  NAND2BX4 U178 ( .AN(n5427), .B(n11193), .Y(n10133) );
  NAND2X6 U179 ( .A(n10464), .B(n10463), .Y(n10822) );
  NAND2X8 U180 ( .A(n3357), .B(n10570), .Y(n10464) );
  OAI2BB2X4 U181 ( .B0(\i_MIPS/n182 ), .B1(net108192), .A0N(n5545), .A1N(n4326), .Y(\i_MIPS/N122 ) );
  NAND2BX1 U182 ( .AN(n4247), .B(n11309), .Y(n6259) );
  NAND4X4 U183 ( .A(n6259), .B(n6258), .C(n6257), .D(n6256), .Y(n10348) );
  INVX3 U184 ( .A(n11353), .Y(n10920) );
  NAND2BX1 U185 ( .AN(n4247), .B(n11310), .Y(n6295) );
  NOR2X1 U186 ( .A(n10347), .B(n10346), .Y(n10351) );
  CLKAND2X12 U187 ( .A(net97686), .B(net97687), .Y(n3835) );
  NAND3X6 U188 ( .A(n6504), .B(n7400), .C(n3413), .Y(n6514) );
  NAND3X4 U189 ( .A(n3642), .B(n3643), .C(net104409), .Y(n4136) );
  BUFX12 U190 ( .A(net100791), .Y(net112420) );
  CLKAND2X4 U191 ( .A(n3785), .B(n4661), .Y(n4525) );
  NAND2BX4 U192 ( .AN(n4247), .B(n11282), .Y(n9953) );
  CLKAND2X12 U193 ( .A(\i_MIPS/ID_EX[80] ), .B(\i_MIPS/ID_EX[79] ), .Y(
        net127709) );
  NAND2BX4 U194 ( .AN(n5428), .B(n11199), .Y(n9711) );
  OR2X6 U195 ( .A(n10336), .B(n10337), .Y(n10539) );
  NAND4XL U196 ( .A(\i_MIPS/PHT_2/current_state_2[1] ), .B(n270), .C(n11064), 
        .D(net97592), .Y(n11056) );
  CLKAND2X3 U197 ( .A(n4194), .B(n4195), .Y(n3342) );
  CLKAND2X3 U198 ( .A(n4235), .B(n4236), .Y(n3341) );
  OAI221X4 U199 ( .A0(\i_MIPS/Register/register[18][28] ), .A1(n4691), .B0(
        \i_MIPS/Register/register[26][28] ), .B1(n4687), .C0(n8514), .Y(n8522)
         );
  INVX4 U200 ( .A(n6611), .Y(n6612) );
  CLKAND2X3 U201 ( .A(\i_MIPS/n316 ), .B(\i_MIPS/n318 ), .Y(n4445) );
  AO21X4 U202 ( .A0(net98371), .A1(net98372), .B0(net111904), .Y(net98572) );
  NAND2X4 U203 ( .A(net98571), .B(net98572), .Y(n4096) );
  INVX4 U204 ( .A(n10665), .Y(n9219) );
  OA22X2 U205 ( .A0(n10139), .A1(n4675), .B0(n10142), .B1(n4250), .Y(n6439) );
  CLKBUFX8 U206 ( .A(n5041), .Y(n5036) );
  NAND2X6 U207 ( .A(net98363), .B(net98364), .Y(n3898) );
  OA21X2 U208 ( .A0(n7498), .A1(n7515), .B0(n7528), .Y(n7499) );
  NAND2X2 U209 ( .A(n6550), .B(\i_MIPS/n359 ), .Y(n7684) );
  OA22X2 U210 ( .A0(net133471), .A1(n7154), .B0(n7147), .B1(n7901), .Y(n7180)
         );
  NAND2X8 U211 ( .A(net128301), .B(\i_MIPS/ID_EX[83] ), .Y(n9455) );
  INVX6 U212 ( .A(n10206), .Y(n10247) );
  BUFX8 U213 ( .A(n5313), .Y(n5305) );
  NAND4X4 U214 ( .A(n9957), .B(n9956), .C(n9955), .D(n9954), .Y(n11251) );
  NAND3BX4 U215 ( .AN(n9275), .B(n2210), .C(n9274), .Y(n9277) );
  NAND2X8 U216 ( .A(n7969), .B(\i_MIPS/n370 ), .Y(n7975) );
  BUFX8 U217 ( .A(n10666), .Y(n225) );
  CLKINVX3 U218 ( .A(n5623), .Y(n54) );
  CLKINVX3 U219 ( .A(n5623), .Y(n50) );
  NAND3X2 U220 ( .A(n8537), .B(n8544), .C(net112294), .Y(n8565) );
  INVX4 U221 ( .A(n9068), .Y(n9070) );
  NAND2X6 U222 ( .A(n3666), .B(\i_MIPS/n356 ), .Y(n7805) );
  CLKAND2X12 U223 ( .A(n4164), .B(n4165), .Y(n3666) );
  INVX8 U224 ( .A(n8537), .Y(n8545) );
  INVX8 U225 ( .A(n3430), .Y(n3802) );
  INVX6 U226 ( .A(n3714), .Y(n3830) );
  AND4X6 U227 ( .A(\i_MIPS/n323 ), .B(\i_MIPS/ALUOp[1] ), .C(
        \i_MIPS/ALU_Control/n11 ), .D(\i_MIPS/ID_EX[106] ), .Y(
        \i_MIPS/ALU_Control/n10 ) );
  INVX6 U228 ( .A(n9463), .Y(n9327) );
  MX2X4 U229 ( .A(net103092), .B(net103093), .S0(net107812), .Y(net103089) );
  NAND4BX2 U230 ( .AN(n7966), .B(n7965), .C(n7964), .D(n7963), .Y(net103093)
         );
  CLKBUFX4 U231 ( .A(n5308), .Y(n5288) );
  OAI2BB1X4 U232 ( .A0N(n6941), .A1N(n6940), .B0(n3720), .Y(net99003) );
  OAI222X2 U233 ( .A0(n7984), .A1(net103076), .B0(n9162), .B1(n7901), .C0(
        net101914), .C1(n9151), .Y(n6774) );
  INVX3 U234 ( .A(net98029), .Y(net103582) );
  AOI22X2 U235 ( .A0(net111966), .A1(net98029), .B0(net111962), .B1(n7645), 
        .Y(n3418) );
  AOI2BB1X2 U236 ( .A0N(net137891), .A1N(n7620), .B0(n7619), .Y(n7621) );
  INVXL U237 ( .A(n8336), .Y(n16) );
  XNOR2X4 U238 ( .A(n17), .B(n10775), .Y(n8530) );
  NAND2X2 U239 ( .A(n3423), .B(n10455), .Y(n17) );
  NOR3X6 U240 ( .A(n8271), .B(n8272), .C(n8273), .Y(n18) );
  NOR2X8 U241 ( .A(n8274), .B(n19), .Y(n8275) );
  INVX6 U242 ( .A(n18), .Y(n19) );
  INVX8 U243 ( .A(n10774), .Y(n8336) );
  OAI33X4 U244 ( .A0(n8859), .A1(n8865), .A2(n8266), .B0(n8247), .B1(net101257), .B2(n8259), .Y(n8274) );
  NAND2X4 U245 ( .A(n3821), .B(n8256), .Y(n8273) );
  NAND4X4 U246 ( .A(n8270), .B(n8269), .C(n8268), .D(n8267), .Y(n8271) );
  NAND2X8 U247 ( .A(n8275), .B(net138213), .Y(n10774) );
  INVX6 U248 ( .A(n8850), .Y(n8859) );
  NOR3X6 U249 ( .A(n4149), .B(n4148), .C(n4150), .Y(n7705) );
  CLKAND2X8 U250 ( .A(n7704), .B(net103548), .Y(n4148) );
  INVX16 U251 ( .A(n9461), .Y(n9170) );
  AND4X8 U252 ( .A(n3755), .B(n6368), .C(n6367), .D(n6366), .Y(n3656) );
  AND4X4 U253 ( .A(n3852), .B(n3851), .C(n3850), .D(n3853), .Y(n3755) );
  NAND4X4 U254 ( .A(n6350), .B(n6349), .C(n6348), .D(n6347), .Y(n11506) );
  AOI222X4 U255 ( .A0(n5512), .A1(n11387), .B0(mem_rdata_D[37]), .B1(n235), 
        .C0(n12982), .C1(n5507), .Y(n10988) );
  INVX4 U256 ( .A(n11387), .Y(n10987) );
  NAND2X6 U257 ( .A(n3768), .B(n10285), .Y(n9019) );
  INVX6 U258 ( .A(n5547), .Y(n3729) );
  BUFX20 U259 ( .A(n5549), .Y(n5547) );
  NAND2X6 U260 ( .A(n4185), .B(n4186), .Y(n6402) );
  NAND2X2 U261 ( .A(n4157), .B(n4158), .Y(n6404) );
  CLKAND2X8 U262 ( .A(n4130), .B(n4131), .Y(n3935) );
  INVX6 U263 ( .A(net98012), .Y(net104408) );
  OAI31X2 U264 ( .A0(n9481), .A1(n8542), .A2(n8726), .B0(n8541), .Y(n8561) );
  NAND2X6 U265 ( .A(n3416), .B(n10580), .Y(n4325) );
  XNOR2XL U266 ( .A(n9885), .B(\i_MIPS/IR_ID[18] ), .Y(n4531) );
  MX2X6 U267 ( .A(\i_MIPS/n317 ), .B(n6444), .S0(\i_MIPS/ID_EX_5 ), .Y(n9885)
         );
  INVX4 U268 ( .A(n10578), .Y(n3753) );
  NAND2X4 U269 ( .A(n10463), .B(n10823), .Y(n10572) );
  NAND2X2 U270 ( .A(n9163), .B(net101908), .Y(n3429) );
  NAND3BX4 U271 ( .AN(n6580), .B(n4450), .C(n9144), .Y(n6581) );
  NAND2X8 U272 ( .A(n6556), .B(\i_MIPS/n356 ), .Y(n7527) );
  INVX6 U273 ( .A(n3666), .Y(n6556) );
  MXI2X8 U274 ( .A(n3699), .B(\i_MIPS/ID_EX[84] ), .S0(n5623), .Y(n6549) );
  INVX16 U275 ( .A(n6549), .Y(n6545) );
  INVX4 U276 ( .A(net97753), .Y(net101465) );
  OAI2BB2X2 U277 ( .B0(n3787), .B1(n3655), .A0N(net111968), .A1N(net97753), 
        .Y(net101552) );
  OR2X4 U278 ( .A(net101465), .B(net111634), .Y(n4177) );
  CLKAND2X12 U279 ( .A(net97574), .B(n4141), .Y(n4140) );
  INVX6 U280 ( .A(n6680), .Y(n6706) );
  AND4X4 U281 ( .A(n3908), .B(n6499), .C(n6498), .D(n6497), .Y(n3907) );
  NAND2X4 U282 ( .A(n6587), .B(\i_MIPS/n345 ), .Y(n8949) );
  NAND3X4 U283 ( .A(n25), .B(n26), .C(net104741), .Y(net99151) );
  AOI32X4 U284 ( .A0(n8863), .A1(n8862), .A2(n4443), .B0(n8861), .B1(net100585), .Y(n8870) );
  AOI33X4 U285 ( .A0(n8863), .A1(n4662), .A2(net101910), .B0(net137952), .B1(
        n7889), .B2(n7888), .Y(n7908) );
  NAND2X1 U286 ( .A(n4519), .B(net107804), .Y(n7887) );
  OA22X1 U287 ( .A0(n5121), .A1(n1692), .B0(n5063), .B1(n3288), .Y(n10025) );
  CLKBUFX6 U288 ( .A(n5125), .Y(n5121) );
  OAI2BB2X1 U289 ( .B0(\i_MIPS/n173 ), .B1(net108192), .A0N(n4315), .A1N(
        n10547), .Y(\i_MIPS/N113 ) );
  CLKINVX2 U290 ( .A(n10551), .Y(n10547) );
  INVX6 U291 ( .A(n10787), .Y(n6640) );
  INVX6 U292 ( .A(\i_MIPS/ALUin1[9] ), .Y(net103561) );
  NAND2X6 U293 ( .A(net103561), .B(n6529), .Y(n8641) );
  NAND2X8 U294 ( .A(\i_MIPS/ALUin1[9] ), .B(n6543), .Y(n8642) );
  NAND2X4 U295 ( .A(n6543), .B(net103561), .Y(n8631) );
  INVX16 U296 ( .A(n9350), .Y(n9044) );
  AND3X4 U297 ( .A(n6296), .B(n10349), .C(n10347), .Y(n6297) );
  BUFX16 U298 ( .A(n5268), .Y(n5265) );
  OA22XL U299 ( .A0(n5198), .A1(n1529), .B0(n5155), .B1(n3109), .Y(n6204) );
  AND2X4 U300 ( .A(n4208), .B(n4209), .Y(n3330) );
  XNOR2X2 U301 ( .A(n3411), .B(n11506), .Y(n6351) );
  NAND2BX1 U302 ( .AN(n5428), .B(n11215), .Y(n6289) );
  AND2XL U303 ( .A(n5557), .B(n11215), .Y(n12905) );
  OR2X6 U304 ( .A(net102791), .B(net111634), .Y(n3703) );
  INVX12 U305 ( .A(n8946), .Y(n4320) );
  BUFX20 U306 ( .A(n9989), .Y(n4955) );
  INVX16 U307 ( .A(n4330), .Y(n9989) );
  AO21X4 U308 ( .A0(net99164), .A1(net99165), .B0(net111904), .Y(net99161) );
  XOR2X4 U309 ( .A(n3916), .B(n4633), .Y(n3851) );
  INVX6 U310 ( .A(n3704), .Y(n3705) );
  INVX8 U311 ( .A(n3696), .Y(net105783) );
  INVX3 U312 ( .A(net97770), .Y(net105046) );
  OAI222X2 U313 ( .A0(net101914), .A1(n9246), .B0(net103076), .B1(n7488), .C0(
        n3762), .C1(n7420), .Y(n6855) );
  INVX1 U314 ( .A(n11433), .Y(n10995) );
  NAND3X6 U315 ( .A(n71), .B(n72), .C(n8603), .Y(n8627) );
  OR2X2 U316 ( .A(n10995), .B(n4250), .Y(n72) );
  OA22X1 U317 ( .A0(n4912), .A1(n1161), .B0(n4249), .B1(n2717), .Y(n8592) );
  OR2X8 U318 ( .A(n3714), .B(net111634), .Y(n3692) );
  NAND3BX2 U319 ( .AN(n264), .B(n8175), .C(net111994), .Y(n8185) );
  NAND3BX2 U320 ( .AN(n8453), .B(n8175), .C(net112294), .Y(n8152) );
  INVX4 U321 ( .A(n6594), .Y(n6585) );
  NAND3X8 U322 ( .A(n7170), .B(n7169), .C(n7168), .Y(n9145) );
  NAND3X6 U323 ( .A(n6540), .B(net102427), .C(n8338), .Y(n7050) );
  NAND3X8 U324 ( .A(n6917), .B(net103889), .C(n6916), .Y(n6540) );
  NAND3X6 U325 ( .A(n7161), .B(n7162), .C(n7160), .Y(n7169) );
  CLKAND2X2 U326 ( .A(n10567), .B(n10566), .Y(n1987) );
  AOI222X4 U327 ( .A0(n5505), .A1(n11374), .B0(mem_rdata_D[24]), .B1(n235), 
        .C0(n12963), .C1(n5502), .Y(n10783) );
  INVX6 U328 ( .A(n11374), .Y(n10782) );
  NAND4X4 U329 ( .A(n8308), .B(n8307), .C(n8306), .D(n8305), .Y(n11374) );
  NAND3X6 U330 ( .A(n255), .B(n9065), .C(n9066), .Y(n8952) );
  NAND2X4 U331 ( .A(n6538), .B(\i_MIPS/n370 ), .Y(n7982) );
  AO22X4 U332 ( .A0(mem_rdata_I[27]), .A1(n5535), .B0(n252), .B1(n11213), .Y(
        n11159) );
  NAND4X2 U333 ( .A(n6251), .B(n6250), .C(n6249), .D(n6248), .Y(n11213) );
  OR2X6 U334 ( .A(n9115), .B(net111634), .Y(n3775) );
  CLKAND2X12 U335 ( .A(n6966), .B(n7876), .Y(n4618) );
  MX2X1 U336 ( .A(DCACHE_addr[23]), .B(n10487), .S0(n204), .Y(\i_MIPS/n444 )
         );
  OA22XL U337 ( .A0(n4760), .A1(n2417), .B0(n4796), .B1(n731), .Y(n6814) );
  OA22XL U338 ( .A0(n4760), .A1(n1394), .B0(n4795), .B1(n2924), .Y(n6806) );
  OA22XL U339 ( .A0(n4760), .A1(n2420), .B0(n4796), .B1(n735), .Y(n6883) );
  CLKBUFX3 U340 ( .A(n4767), .Y(n4760) );
  INVX8 U341 ( .A(net112999), .Y(net104252) );
  OA22X1 U342 ( .A0(n5367), .A1(n1689), .B0(n5348), .B1(n3284), .Y(n10088) );
  OAI2BB2X1 U343 ( .B0(\i_MIPS/n178 ), .B1(net108190), .A0N(n4073), .A1N(
        n10837), .Y(\i_MIPS/N118 ) );
  NAND4X4 U344 ( .A(n6399), .B(n3806), .C(n6400), .D(n3805), .Y(n11486) );
  XOR2X2 U345 ( .A(n12949), .B(n11486), .Y(n6401) );
  MXI2X4 U346 ( .A(n10957), .B(n10956), .S0(n5522), .Y(n10958) );
  NAND3BX4 U347 ( .AN(n11058), .B(n11064), .C(n11060), .Y(n11059) );
  CLKMX2X6 U348 ( .A(n11057), .B(n3605), .S0(net112691), .Y(n11058) );
  CLKINVX16 U349 ( .A(n5625), .Y(n5623) );
  INVX4 U350 ( .A(net100402), .Y(net98620) );
  NAND2X6 U351 ( .A(n9164), .B(net107804), .Y(n8457) );
  CLKINVX12 U352 ( .A(n9467), .Y(n9164) );
  INVX12 U353 ( .A(net98630), .Y(net97452) );
  INVX16 U354 ( .A(n11347), .Y(n5549) );
  AOI222X4 U355 ( .A0(n5498), .A1(n11432), .B0(mem_rdata_D[82]), .B1(n234), 
        .C0(n12969), .C1(n4385), .Y(n10512) );
  NAND2X8 U356 ( .A(n3819), .B(n6749), .Y(n10867) );
  NAND4BX2 U357 ( .AN(n6699), .B(n6698), .C(n6697), .D(n6696), .Y(n6700) );
  OAI221X4 U358 ( .A0(n9342), .A1(n9335), .B0(n6692), .B1(net133688), .C0(
        n6691), .Y(n6701) );
  CLKBUFX4 U359 ( .A(n5305), .Y(n5300) );
  OAI2BB2X1 U360 ( .B0(\i_MIPS/n172 ), .B1(net108190), .A0N(n4315), .A1N(
        n11122), .Y(\i_MIPS/N112 ) );
  XOR3X1 U361 ( .A(net112400), .B(n11121), .C(n11120), .Y(n11125) );
  NOR2X4 U362 ( .A(n6011), .B(n6010), .Y(n6110) );
  NAND3X2 U363 ( .A(n5999), .B(n5998), .C(n5997), .Y(n6011) );
  CLKBUFX16 U364 ( .A(n12868), .Y(mem_wdata_I[74]) );
  CLKAND2X12 U365 ( .A(n4468), .B(n8535), .Y(n2210) );
  OAI222X1 U366 ( .A0(\i_MIPS/PC/n11 ), .A1(net97444), .B0(net97445), .B1(
        n10585), .C0(n4404), .C1(net108704), .Y(n10590) );
  INVX8 U367 ( .A(n7617), .Y(n7806) );
  NAND3X6 U368 ( .A(\i_MIPS/PC/n5 ), .B(n10176), .C(n9569), .Y(n3428) );
  XNOR2X4 U369 ( .A(n10453), .B(net112404), .Y(n10458) );
  BUFX20 U370 ( .A(net100398), .Y(n3917) );
  AO22X2 U371 ( .A0(net111992), .A1(n6706), .B0(net112296), .B1(n6704), .Y(
        n6600) );
  CLKINVX6 U372 ( .A(n8486), .Y(n10356) );
  AOI2BB1X4 U373 ( .A0N(n9044), .A1N(n8449), .B0(net101257), .Y(n8461) );
  INVX12 U374 ( .A(n8072), .Y(n7800) );
  NAND2X8 U375 ( .A(n6552), .B(\i_MIPS/n353 ), .Y(n8737) );
  INVX8 U376 ( .A(n6574), .Y(n6552) );
  MXI2X4 U377 ( .A(n10292), .B(n10291), .S0(n5515), .Y(n10293) );
  OA22XL U378 ( .A0(n4761), .A1(n3003), .B0(n4795), .B1(n570), .Y(n6431) );
  INVX4 U379 ( .A(n4761), .Y(n4507) );
  NAND2X6 U380 ( .A(n10851), .B(n10850), .Y(n10792) );
  NAND2X6 U381 ( .A(n3754), .B(n3753), .Y(n4231) );
  NAND3X4 U382 ( .A(n10571), .B(n10570), .C(n3357), .Y(n3754) );
  INVX20 U383 ( .A(n4142), .Y(net97444) );
  NAND2X8 U384 ( .A(net98620), .B(n4146), .Y(n4142) );
  CLKBUFX20 U385 ( .A(n10638), .Y(n4247) );
  CLKBUFX12 U386 ( .A(n3428), .Y(n5427) );
  NAND2BX4 U387 ( .AN(n10252), .B(n10325), .Y(n10634) );
  INVX16 U388 ( .A(net112676), .Y(n3637) );
  NAND3X8 U389 ( .A(n3924), .B(n3925), .C(n3923), .Y(n3922) );
  INVX6 U390 ( .A(n80), .Y(n81) );
  NAND4X6 U391 ( .A(n4350), .B(n4351), .C(n9973), .D(n9972), .Y(n11349) );
  BUFX2 U392 ( .A(n4924), .Y(n4918) );
  AND2X4 U393 ( .A(n4214), .B(n4215), .Y(n3338) );
  NAND3X6 U394 ( .A(n107), .B(n108), .C(net103720), .Y(n4133) );
  OR2X8 U395 ( .A(net103719), .B(net111636), .Y(n108) );
  OA22X2 U396 ( .A0(n10959), .A1(n4245), .B0(n10962), .B1(n4246), .Y(n7589) );
  INVX3 U397 ( .A(n11382), .Y(n10962) );
  AND4X8 U398 ( .A(n4460), .B(\i_MIPS/EX_MEM_1 ), .C(DCACHE_ren), .D(n11345), 
        .Y(n2017) );
  NAND2X4 U399 ( .A(n8240), .B(n7497), .Y(n7689) );
  INVX1 U400 ( .A(n7497), .Y(n7493) );
  CLKAND2X4 U401 ( .A(n7497), .B(n7523), .Y(n4451) );
  NAND2X4 U402 ( .A(n7497), .B(n7496), .Y(n7515) );
  INVXL U403 ( .A(n9547), .Y(n20) );
  OR2X2 U404 ( .A(n9548), .B(net111622), .Y(n21) );
  OR2X4 U405 ( .A(n9547), .B(net111634), .Y(n22) );
  NAND3X6 U406 ( .A(n21), .B(n22), .C(n9546), .Y(n3896) );
  CLKINVX8 U407 ( .A(n10557), .Y(n9547) );
  NAND4X4 U408 ( .A(n9498), .B(n9495), .C(n9496), .D(n9497), .Y(n10557) );
  AOI2BB2X4 U409 ( .B0(net111630), .B1(n9429), .A0N(net111644), .A1N(n10313), 
        .Y(n9432) );
  NAND2X2 U410 ( .A(n4505), .B(n4500), .Y(n9413) );
  CLKAND2X12 U411 ( .A(\i_MIPS/IR_ID[16] ), .B(\i_MIPS/n314 ), .Y(n4505) );
  INVX12 U412 ( .A(n6550), .Y(n6561) );
  NAND3BX4 U413 ( .AN(n11062), .B(n11064), .C(n11065), .Y(n11063) );
  CLKAND2X12 U414 ( .A(n8946), .B(n8748), .Y(n8756) );
  NAND3X8 U415 ( .A(ICACHE_addr[10]), .B(ICACHE_addr[9]), .C(n10233), .Y(
        n10235) );
  CLKINVX8 U416 ( .A(n10232), .Y(n10233) );
  NAND3X8 U417 ( .A(n4230), .B(n4231), .C(n10577), .Y(n10851) );
  INVX4 U418 ( .A(n10572), .Y(n10576) );
  NAND2X2 U419 ( .A(n10836), .B(net112404), .Y(n10573) );
  BUFX12 U420 ( .A(n3786), .Y(n224) );
  CLKINVX3 U421 ( .A(n10468), .Y(n10465) );
  OAI222X1 U422 ( .A0(\i_MIPS/PC/n27 ), .A1(net108686), .B0(n3637), .B1(n10468), .C0(n4398), .C1(net108704), .Y(n10473) );
  NOR2X8 U423 ( .A(n4101), .B(n4102), .Y(n4129) );
  OA22X4 U424 ( .A0(n10928), .A1(n4675), .B0(n10931), .B1(n4250), .Y(n6941) );
  INVX8 U425 ( .A(n3905), .Y(n8180) );
  NAND2BX2 U426 ( .AN(n4950), .B(\D_cache/cache[5][154] ), .Y(n6305) );
  AOI2BB2X1 U427 ( .B0(n11360), .B1(n3400), .A0N(n10266), .A1N(n4246), .Y(
        n7360) );
  OA22X2 U428 ( .A0(n4836), .A1(n3354), .B0(n4882), .B1(n1734), .Y(n6328) );
  AND2X4 U429 ( .A(n4196), .B(n4197), .Y(n3329) );
  BUFX12 U430 ( .A(n4421), .Y(n5507) );
  NAND2X6 U431 ( .A(n4319), .B(n10417), .Y(n10431) );
  INVX8 U432 ( .A(n10383), .Y(n10420) );
  NAND4X6 U433 ( .A(n9965), .B(n9964), .C(n9963), .D(n9962), .Y(n11219) );
  OA22X4 U434 ( .A0(n5211), .A1(n1464), .B0(n5168), .B1(n3038), .Y(n9964) );
  OA22X2 U435 ( .A0(n5111), .A1(n1655), .B0(n5056), .B1(n3239), .Y(n9965) );
  CLKBUFX6 U436 ( .A(n5134), .Y(n5111) );
  CLKBUFX6 U437 ( .A(n5087), .Y(n5056) );
  NAND2X2 U438 ( .A(net111960), .B(n8091), .Y(n23) );
  NAND2X2 U439 ( .A(net111968), .B(net98728), .Y(n24) );
  NAND2X4 U440 ( .A(n23), .B(n24), .Y(net102878) );
  BUFX20 U441 ( .A(net100535), .Y(net111960) );
  CLKMX2X4 U442 ( .A(n8066), .B(n8065), .S0(net107816), .Y(n8091) );
  BUFX12 U443 ( .A(net100537), .Y(net111968) );
  INVX6 U444 ( .A(net102878), .Y(net98707) );
  OR2X4 U445 ( .A(net104739), .B(net111624), .Y(n25) );
  OR2X6 U446 ( .A(net104740), .B(net111636), .Y(n26) );
  CLKINVX4 U447 ( .A(net97684), .Y(net104740) );
  OAI2BB1X2 U448 ( .A0N(n10064), .A1N(net99157), .B0(net112782), .Y(net104741)
         );
  OR2X6 U449 ( .A(n6121), .B(n9568), .Y(n27) );
  NAND2X6 U450 ( .A(n27), .B(n4060), .Y(n6119) );
  NAND4X6 U451 ( .A(n6118), .B(n6117), .C(n6116), .D(n6115), .Y(n6121) );
  CLKINVX8 U452 ( .A(n6122), .Y(n9568) );
  INVX12 U453 ( .A(n4059), .Y(n4060) );
  AND2X8 U454 ( .A(n6119), .B(n4651), .Y(n11171) );
  OA21X4 U455 ( .A0(n7047), .A1(n6965), .B0(n6964), .Y(n28) );
  NAND2X6 U456 ( .A(n28), .B(n3685), .Y(n6967) );
  INVX6 U457 ( .A(n6962), .Y(n7047) );
  NAND2X8 U458 ( .A(n8341), .B(n6844), .Y(n6965) );
  BUFX4 U459 ( .A(n6963), .Y(n3685) );
  NAND2X6 U460 ( .A(n6967), .B(n6966), .Y(n7878) );
  NAND2X1 U461 ( .A(n10869), .B(n29), .Y(n30) );
  NAND2X1 U462 ( .A(n10868), .B(n5520), .Y(n31) );
  NAND2X2 U463 ( .A(n30), .B(n31), .Y(n32) );
  CLKINVX1 U464 ( .A(n5520), .Y(n29) );
  INVX3 U465 ( .A(n32), .Y(n10870) );
  CLKINVX1 U466 ( .A(n11477), .Y(n10868) );
  OR2X8 U467 ( .A(n10327), .B(n10337), .Y(n33) );
  OR2X2 U468 ( .A(n4300), .B(net112404), .Y(n34) );
  NAND3X8 U469 ( .A(n33), .B(n34), .C(n10326), .Y(n10538) );
  CLKINVX8 U470 ( .A(n10323), .Y(n10327) );
  NAND2X8 U471 ( .A(n10325), .B(n10324), .Y(n10337) );
  CLKBUFX20 U472 ( .A(net97874), .Y(net112404) );
  CLKINVX8 U473 ( .A(n10538), .Y(n10331) );
  OR2X4 U474 ( .A(net103581), .B(net111624), .Y(n35) );
  OR2X8 U475 ( .A(net103582), .B(net111636), .Y(n36) );
  NAND3X2 U476 ( .A(n35), .B(n36), .C(net103583), .Y(net98027) );
  NOR2X1 U477 ( .A(n4743), .B(n2648), .Y(n37) );
  NOR2X1 U478 ( .A(n4788), .B(n1075), .Y(n38) );
  OR2X1 U479 ( .A(n37), .B(n38), .Y(n4348) );
  CLKBUFX4 U480 ( .A(n4771), .Y(n4743) );
  NAND4BX2 U481 ( .AN(n4348), .B(n9183), .C(n9182), .D(n9181), .Y(n11467) );
  OR2XL U482 ( .A(\i_MIPS/ALUin1[10] ), .B(net112364), .Y(n39) );
  OR2XL U483 ( .A(\i_MIPS/ALUin1[9] ), .B(net112346), .Y(n40) );
  NAND3X1 U484 ( .A(n39), .B(n40), .C(n7897), .Y(n8359) );
  CLKINVX12 U485 ( .A(net112374), .Y(net112364) );
  INVX16 U486 ( .A(net112356), .Y(net112346) );
  OAI222X1 U487 ( .A0(n8359), .A1(net103076), .B0(n8876), .B1(n7901), .C0(
        n8875), .C1(net101914), .Y(n7904) );
  OA21X4 U488 ( .A0(n6717), .A1(n6716), .B0(n6715), .Y(n41) );
  NAND2X8 U489 ( .A(n41), .B(n6714), .Y(n10866) );
  NAND2X1 U490 ( .A(n6695), .B(n6707), .Y(n6717) );
  OAI32X4 U491 ( .A0(n6713), .A1(n6712), .A2(n6711), .B0(n4455), .B1(n4509), 
        .Y(n6714) );
  NAND2X6 U492 ( .A(net111966), .B(n10866), .Y(n10859) );
  OR2X2 U493 ( .A(n10301), .B(n4675), .Y(n42) );
  OR2X2 U494 ( .A(n10304), .B(n4250), .Y(n43) );
  NAND3X6 U495 ( .A(n42), .B(n43), .C(n9398), .Y(n10315) );
  INVX3 U496 ( .A(n11473), .Y(n10301) );
  OA22X2 U497 ( .A0(n10307), .A1(n4245), .B0(n10310), .B1(n4246), .Y(n9398) );
  CLKINVX8 U498 ( .A(n10315), .Y(n9430) );
  OR2X2 U499 ( .A(n4660), .B(n260), .Y(n44) );
  OR2X4 U500 ( .A(net103552), .B(n4587), .Y(n45) );
  NAND3X6 U501 ( .A(n44), .B(n45), .C(n7471), .Y(n8084) );
  CLKBUFX6 U502 ( .A(n8651), .Y(n4660) );
  BUFX8 U503 ( .A(n7473), .Y(n260) );
  NAND2X4 U504 ( .A(n4662), .B(net107798), .Y(net103552) );
  BUFX16 U505 ( .A(n7472), .Y(n4587) );
  OA22X4 U506 ( .A0(n8353), .A1(n7470), .B0(n7469), .B1(n4659), .Y(n7471) );
  OAI32X4 U507 ( .A0(n8085), .A1(\i_MIPS/ID_EX[83] ), .A2(n8084), .B0(
        net133471), .B1(n8753), .Y(n8086) );
  NAND2X4 U508 ( .A(n8095), .B(n8092), .Y(n46) );
  NAND3X4 U509 ( .A(n8093), .B(n8094), .C(n47), .Y(n11462) );
  CLKINVX1 U510 ( .A(n46), .Y(n47) );
  OA22X2 U511 ( .A0(n4750), .A1(n1159), .B0(n4791), .B1(n2879), .Y(n8095) );
  OA22X1 U512 ( .A0(n4823), .A1(n2115), .B0(n4869), .B1(n528), .Y(n8094) );
  OA22XL U513 ( .A0(n4915), .A1(n2126), .B0(n4947), .B1(n539), .Y(n8093) );
  AOI222X1 U514 ( .A0(n5495), .A1(n11462), .B0(mem_rdata_D[112]), .B1(n234), 
        .C0(n12971), .C1(n5494), .Y(n10289) );
  OR2X4 U515 ( .A(n5300), .B(n1676), .Y(n48) );
  OR2X1 U516 ( .A(n5255), .B(n3264), .Y(n49) );
  AND2X4 U517 ( .A(n48), .B(n49), .Y(n9899) );
  NAND2X6 U518 ( .A(\i_MIPS/n309 ), .B(n50), .Y(n51) );
  NAND2X2 U519 ( .A(net137684), .B(n5623), .Y(n52) );
  NAND2X8 U520 ( .A(n51), .B(n52), .Y(n7464) );
  INVX8 U521 ( .A(n7464), .Y(n7475) );
  OR3X8 U522 ( .A(n8234), .B(n8233), .C(n8232), .Y(n53) );
  NAND2X8 U523 ( .A(n53), .B(n8231), .Y(n8235) );
  INVX4 U524 ( .A(n9141), .Y(n8234) );
  NAND2X8 U525 ( .A(n9262), .B(n9152), .Y(n8232) );
  INVX16 U526 ( .A(n8945), .Y(n8231) );
  NAND2X8 U527 ( .A(n9475), .B(n8235), .Y(n8850) );
  NAND2X6 U528 ( .A(\i_MIPS/n277 ), .B(n54), .Y(n55) );
  NAND2X2 U529 ( .A(n4493), .B(n5623), .Y(n56) );
  NAND2X8 U530 ( .A(n55), .B(n56), .Y(n6575) );
  NAND2X4 U531 ( .A(n6575), .B(\i_MIPS/n355 ), .Y(n8749) );
  INVX8 U532 ( .A(n6575), .Y(n6551) );
  NAND2X4 U533 ( .A(\i_MIPS/ALUin1[16] ), .B(n6575), .Y(n8071) );
  NAND2X1 U534 ( .A(n10950), .B(n57), .Y(n58) );
  NAND2XL U535 ( .A(n10949), .B(n5522), .Y(n59) );
  NAND2X2 U536 ( .A(n58), .B(n59), .Y(n60) );
  CLKINVX1 U537 ( .A(n5522), .Y(n57) );
  INVX3 U538 ( .A(n60), .Y(n10951) );
  INVX4 U539 ( .A(n11405), .Y(n10949) );
  OR2X1 U540 ( .A(n9469), .B(n8260), .Y(n61) );
  OR2X4 U541 ( .A(net102405), .B(n8264), .Y(n62) );
  OR2X8 U542 ( .A(n7463), .B(net137891), .Y(n63) );
  NAND3X6 U543 ( .A(n61), .B(n62), .C(n63), .Y(n7064) );
  NAND2X8 U544 ( .A(net128301), .B(n4443), .Y(n9469) );
  NAND2X2 U545 ( .A(n4520), .B(net107802), .Y(n8260) );
  CLKMX2X8 U546 ( .A(n7062), .B(n7061), .S0(net107794), .Y(n7463) );
  AO21X2 U547 ( .A0(n3838), .A1(n8249), .B0(n7064), .Y(n4170) );
  NAND2X2 U548 ( .A(n10848), .B(n65), .Y(n66) );
  NAND2X4 U549 ( .A(n64), .B(ICACHE_addr[29]), .Y(n67) );
  NAND2X6 U550 ( .A(n66), .B(n67), .Y(n10857) );
  INVX3 U551 ( .A(n10848), .Y(n64) );
  INVXL U552 ( .A(ICACHE_addr[29]), .Y(n65) );
  INVX4 U553 ( .A(n10857), .Y(n10863) );
  NAND2X4 U554 ( .A(n3839), .B(n68), .Y(n69) );
  NAND2X2 U555 ( .A(\i_MIPS/n297 ), .B(n5625), .Y(n70) );
  NAND2X8 U556 ( .A(n69), .B(n70), .Y(n6534) );
  CLKINVX2 U557 ( .A(n5625), .Y(n68) );
  NAND2X8 U558 ( .A(\i_MIPS/ALUin1[6] ), .B(n6534), .Y(n7511) );
  NAND2X6 U559 ( .A(n6534), .B(n7696), .Y(n7877) );
  INVX6 U560 ( .A(n6534), .Y(n6536) );
  OR2X2 U561 ( .A(n10991), .B(n4675), .Y(n71) );
  BUFX20 U562 ( .A(n3424), .Y(n4675) );
  OA22X2 U563 ( .A0(n10999), .A1(n4245), .B0(n11004), .B1(n4246), .Y(n8603) );
  OR2X1 U564 ( .A(n9250), .B(n9249), .Y(n73) );
  OR2XL U565 ( .A(n9248), .B(n9467), .Y(n74) );
  NAND3X2 U566 ( .A(n73), .B(n74), .C(n4658), .Y(n9259) );
  CLKINVX6 U567 ( .A(n8069), .Y(n9250) );
  NAND2X4 U568 ( .A(n9328), .B(net107804), .Y(n9249) );
  CLKINVX3 U569 ( .A(n6850), .Y(n9248) );
  CLKAND2X2 U570 ( .A(n4422), .B(n9154), .Y(n75) );
  AND2X6 U571 ( .A(n6764), .B(n6763), .Y(n76) );
  CLKAND2X3 U572 ( .A(n6762), .B(n6761), .Y(n77) );
  NOR3X4 U573 ( .A(n75), .B(n76), .C(n77), .Y(n6776) );
  AND2X2 U574 ( .A(net101910), .B(n8958), .Y(n4422) );
  OR2X4 U575 ( .A(n9018), .B(net111622), .Y(n78) );
  OR2X4 U576 ( .A(n3893), .B(net111634), .Y(n79) );
  NAND3X6 U577 ( .A(n78), .B(n79), .C(n9017), .Y(n10300) );
  BUFX16 U578 ( .A(n10300), .Y(n4592) );
  NOR3X4 U579 ( .A(n7176), .B(n7177), .C(n7175), .Y(n80) );
  NOR2X6 U580 ( .A(n7174), .B(n81), .Y(n7178) );
  OAI32X4 U581 ( .A0(net101257), .A1(n4441), .A2(n413), .B0(n413), .B1(n7173), 
        .Y(n7174) );
  OAI32X2 U582 ( .A0(n7156), .A1(n7155), .A2(net112300), .B0(n7887), .B1(n7234), .Y(n7176) );
  AND3X6 U583 ( .A(n4441), .B(n7171), .C(net137952), .Y(n7175) );
  CLKMX2X8 U584 ( .A(net112415), .B(net101082), .S0(n7153), .Y(n7177) );
  NAND4X8 U585 ( .A(n7180), .B(n7178), .C(n7179), .D(n4658), .Y(net98012) );
  NAND2X2 U586 ( .A(n6803), .B(n6805), .Y(n82) );
  NAND3X6 U587 ( .A(n6806), .B(n6804), .C(n83), .Y(n11419) );
  INVX3 U588 ( .A(n82), .Y(n83) );
  OA22X2 U589 ( .A0(n4833), .A1(n1248), .B0(n4878), .B1(n2790), .Y(n6805) );
  OA22X2 U590 ( .A0(n4985), .A1(n828), .B0(n5031), .B1(n2391), .Y(n6803) );
  AOI222X4 U591 ( .A0(n5500), .A1(n11419), .B0(mem_rdata_D[69]), .B1(n234), 
        .C0(n12982), .C1(n4385), .Y(n10982) );
  INVX8 U592 ( .A(n11419), .Y(n10981) );
  NAND3X2 U593 ( .A(n8699), .B(n8697), .C(n8698), .Y(n84) );
  NAND2X8 U594 ( .A(n85), .B(n8696), .Y(n11391) );
  INVX4 U595 ( .A(n84), .Y(n85) );
  OA22X2 U596 ( .A0(n4746), .A1(n810), .B0(n4789), .B1(n2373), .Y(n8699) );
  OA22XL U597 ( .A0(n4915), .A1(n2166), .B0(n4947), .B1(n592), .Y(n8697) );
  INVX8 U598 ( .A(n11391), .Y(n10704) );
  NAND2X1 U599 ( .A(n11333), .B(n87), .Y(n88) );
  NAND2X4 U600 ( .A(n86), .B(ICACHE_addr[18]), .Y(n89) );
  NAND2X2 U601 ( .A(n88), .B(n89), .Y(n5982) );
  INVX3 U602 ( .A(n11333), .Y(n86) );
  INVXL U603 ( .A(ICACHE_addr[18]), .Y(n87) );
  NAND4X4 U604 ( .A(n5976), .B(n5975), .C(n5974), .D(n5973), .Y(n11333) );
  NOR2X6 U605 ( .A(n5982), .B(n5981), .Y(n5999) );
  NAND2X1 U606 ( .A(n10476), .B(n90), .Y(n91) );
  NAND2X1 U607 ( .A(n10475), .B(n5515), .Y(n92) );
  NAND2X2 U608 ( .A(n91), .B(n92), .Y(n93) );
  CLKINVX1 U609 ( .A(n5515), .Y(n90) );
  INVX4 U610 ( .A(n93), .Y(n10477) );
  NAND2X2 U611 ( .A(n4416), .B(n4570), .Y(n94) );
  CLKINVX1 U612 ( .A(n8751), .Y(n95) );
  NAND2X6 U613 ( .A(n95), .B(n94), .Y(n8076) );
  CLKAND2X2 U614 ( .A(n7803), .B(n7805), .Y(n4416) );
  NAND2X4 U615 ( .A(n8076), .B(n8749), .Y(n7807) );
  CLKINVX4 U616 ( .A(n8076), .Y(n8078) );
  OR2X1 U617 ( .A(n4978), .B(n747), .Y(n96) );
  OR2X2 U618 ( .A(n5023), .B(n2308), .Y(n97) );
  AND2X2 U619 ( .A(n96), .B(n97), .Y(n7739) );
  NAND4X2 U620 ( .A(n7742), .B(n7741), .C(n7740), .D(n7739), .Y(n11459) );
  NOR2X2 U621 ( .A(n8578), .B(n8580), .Y(n98) );
  NOR3X2 U622 ( .A(n8577), .B(n99), .C(n8579), .Y(n8581) );
  INVX1 U623 ( .A(n98), .Y(n99) );
  AO22X1 U624 ( .A0(net112178), .A1(n272), .B0(net112160), .B1(n2004), .Y(
        n8580) );
  AO22XL U625 ( .A0(n145), .A1(n320), .B0(n226), .B1(n428), .Y(n8577) );
  NAND4BX2 U626 ( .AN(n8584), .B(n8583), .C(n8582), .D(n8581), .Y(n8585) );
  CLKAND2X3 U627 ( .A(n7756), .B(n7755), .Y(n100) );
  OR2X8 U628 ( .A(n100), .B(n3665), .Y(net112736) );
  NAND2X1 U629 ( .A(n9940), .B(n9938), .Y(n101) );
  NAND3X4 U630 ( .A(n9939), .B(n9941), .C(n102), .Y(n11188) );
  CLKINVX1 U631 ( .A(n101), .Y(n102) );
  OA22XL U632 ( .A0(n5120), .A1(n1489), .B0(n5088), .B1(n3073), .Y(n9941) );
  OA22X2 U633 ( .A0(n5210), .A1(n2740), .B0(n5167), .B1(n1280), .Y(n9940) );
  AO22X4 U634 ( .A0(mem_rdata_I[2]), .A1(n5536), .B0(n249), .B1(n11188), .Y(
        n11104) );
  NAND2BX4 U635 ( .AN(n5427), .B(n11188), .Y(n9947) );
  NAND2X1 U636 ( .A(n10305), .B(n103), .Y(n104) );
  NAND2X1 U637 ( .A(n10304), .B(n5515), .Y(n105) );
  NAND2X2 U638 ( .A(n104), .B(n105), .Y(n106) );
  CLKINVX1 U639 ( .A(n5515), .Y(n103) );
  INVX3 U640 ( .A(n106), .Y(n10306) );
  OR2X2 U641 ( .A(net103718), .B(net111624), .Y(n107) );
  OAI2BB1X2 U642 ( .A0N(net98366), .A1N(net98367), .B0(net112782), .Y(
        net103720) );
  CLKAND2X4 U643 ( .A(net100581), .B(net103354), .Y(n109) );
  NOR2X2 U644 ( .A(n109), .B(net105012), .Y(net128963) );
  CLKINVX2 U645 ( .A(net103710), .Y(net100581) );
  INVX8 U646 ( .A(net103552), .Y(net103354) );
  NAND2X1 U647 ( .A(net101910), .B(net128963), .Y(net105006) );
  OR2X2 U648 ( .A(net102405), .B(n8968), .Y(n110) );
  OR2X1 U649 ( .A(net101914), .B(n8964), .Y(n111) );
  OR2X2 U650 ( .A(net104229), .B(net137891), .Y(n112) );
  NAND3X2 U651 ( .A(n110), .B(n111), .C(n112), .Y(n7319) );
  NAND2X6 U652 ( .A(n8862), .B(\i_MIPS/ID_EX[83] ), .Y(net102405) );
  NAND2X2 U653 ( .A(n7316), .B(n4536), .Y(n8968) );
  MX2X2 U654 ( .A(net104885), .B(net104868), .S0(net107794), .Y(net104229) );
  BUFX20 U655 ( .A(net102393), .Y(net137891) );
  NAND2X6 U656 ( .A(n9952), .B(n9950), .Y(n113) );
  NAND3X8 U657 ( .A(n9953), .B(n9951), .C(n114), .Y(n11067) );
  INVX8 U658 ( .A(n113), .Y(n114) );
  NAND2BX2 U659 ( .AN(n5425), .B(n11250), .Y(n9952) );
  OAI2BB2X2 U660 ( .B0(\i_MIPS/n215 ), .B1(net108198), .A0N(n5545), .A1N(
        n11067), .Y(\i_MIPS/N58 ) );
  NAND2X2 U661 ( .A(net98335), .B(net98336), .Y(n115) );
  CLKINVX1 U662 ( .A(net111904), .Y(n116) );
  NAND2X4 U663 ( .A(n115), .B(n116), .Y(net97937) );
  INVX4 U664 ( .A(net111910), .Y(net111904) );
  AND2XL U665 ( .A(net97936), .B(net97937), .Y(n4405) );
  NAND2X6 U666 ( .A(n9968), .B(n9966), .Y(n117) );
  NAND3X8 U667 ( .A(n9967), .B(n9969), .C(n118), .Y(n11076) );
  CLKINVX8 U668 ( .A(n117), .Y(n118) );
  NAND2BX4 U669 ( .AN(n5425), .B(n11251), .Y(n9968) );
  NAND2BX4 U670 ( .AN(n5429), .B(n11219), .Y(n9966) );
  OAI2BB2X2 U671 ( .B0(\i_MIPS/n216 ), .B1(net108198), .A0N(n4072), .A1N(
        n11076), .Y(\i_MIPS/N59 ) );
  INVX12 U672 ( .A(n11076), .Y(n11081) );
  AND2XL U673 ( .A(n5498), .B(n11440), .Y(n119) );
  AND2X2 U674 ( .A(mem_rdata_D[90]), .B(n234), .Y(n120) );
  AND2XL U675 ( .A(n12961), .B(n4385), .Y(n121) );
  NOR3X1 U676 ( .A(n119), .B(n120), .C(n121), .Y(n10273) );
  BUFX20 U677 ( .A(n10994), .Y(n5498) );
  MXI2X4 U678 ( .A(n10273), .B(n10272), .S0(n5515), .Y(n10274) );
  OR2X2 U679 ( .A(n8527), .B(net111622), .Y(n122) );
  OR2X8 U680 ( .A(n8526), .B(net111634), .Y(n123) );
  NAND3X6 U681 ( .A(n122), .B(n123), .C(n8525), .Y(n10474) );
  INVX3 U682 ( .A(n10320), .Y(n8526) );
  BUFX16 U683 ( .A(n10474), .Y(n262) );
  OA21X2 U684 ( .A0(n4412), .A1(n7051), .B0(n4417), .Y(n124) );
  NAND2X2 U685 ( .A(n124), .B(n7160), .Y(n7222) );
  CLKAND2X12 U686 ( .A(n7509), .B(n7502), .Y(n4412) );
  AND2X4 U687 ( .A(n7874), .B(n7881), .Y(n4417) );
  AOI21X2 U688 ( .A0(n7222), .A1(n3343), .B0(n7223), .Y(n7224) );
  NAND2X4 U689 ( .A(n7222), .B(n7880), .Y(n8637) );
  NAND2XL U690 ( .A(n8632), .B(net100585), .Y(n125) );
  NAND2X2 U691 ( .A(n7057), .B(n7056), .Y(n126) );
  NAND2X1 U692 ( .A(n7055), .B(n7054), .Y(n127) );
  AND3X4 U693 ( .A(n125), .B(n126), .C(n127), .Y(n7066) );
  AO22X1 U694 ( .A0(n7052), .A1(net137952), .B0(net112296), .B1(n8634), .Y(
        n7055) );
  NAND2X2 U695 ( .A(n11321), .B(n129), .Y(n130) );
  NAND2X6 U696 ( .A(n128), .B(n3781), .Y(n131) );
  NAND2X4 U697 ( .A(n130), .B(n131), .Y(n5992) );
  INVX4 U698 ( .A(n11321), .Y(n128) );
  INVX1 U699 ( .A(n3781), .Y(n129) );
  NOR2X2 U700 ( .A(n5992), .B(n5991), .Y(n5998) );
  NAND2X1 U701 ( .A(n10295), .B(n132), .Y(n133) );
  NAND2X1 U702 ( .A(n10294), .B(n5515), .Y(n134) );
  NAND2X2 U703 ( .A(n133), .B(n134), .Y(n135) );
  CLKINVX1 U704 ( .A(n5515), .Y(n132) );
  INVX3 U705 ( .A(n135), .Y(n10296) );
  INVX3 U706 ( .A(n11366), .Y(n10294) );
  CLKAND2X3 U707 ( .A(mem_rdata_I[25]), .B(n5540), .Y(n136) );
  AND2X2 U708 ( .A(n251), .B(n11211), .Y(n137) );
  OR2X6 U709 ( .A(n136), .B(n137), .Y(n9817) );
  AND2X1 U710 ( .A(mem_rdata_I[12]), .B(n5540), .Y(n138) );
  AND2X2 U711 ( .A(n249), .B(n11198), .Y(n139) );
  OR2X8 U712 ( .A(n138), .B(n139), .Y(n9774) );
  NAND4X2 U713 ( .A(n9773), .B(n9772), .C(n9771), .D(n9770), .Y(n11198) );
  CLKMX2X4 U714 ( .A(\I_cache/cache[0][108] ), .B(n9774), .S0(n5095), .Y(
        n11923) );
  CLKMX2X4 U715 ( .A(\I_cache/cache[1][108] ), .B(n9774), .S0(n5051), .Y(
        n11922) );
  CLKMX2X4 U716 ( .A(\I_cache/cache[2][108] ), .B(n9774), .S0(n5187), .Y(
        n11921) );
  CLKMX2X4 U717 ( .A(\I_cache/cache[3][108] ), .B(n9774), .S0(n5141), .Y(
        n11920) );
  CLKMX2X4 U718 ( .A(\I_cache/cache[4][108] ), .B(n9774), .S0(n5273), .Y(
        n11919) );
  CLKMX2X4 U719 ( .A(\I_cache/cache[5][108] ), .B(n9774), .S0(n5230), .Y(
        n11918) );
  CLKMX2X4 U720 ( .A(\I_cache/cache[6][108] ), .B(n9774), .S0(n5361), .Y(
        n11917) );
  CLKMX2X4 U721 ( .A(\I_cache/cache[7][108] ), .B(n9774), .S0(n5319), .Y(
        n11916) );
  BUFX12 U722 ( .A(n6201), .Y(n140) );
  AO22X1 U723 ( .A0(mem_rdata_I[126]), .A1(n5542), .B0(n253), .B1(n11312), .Y(
        n6201) );
  BUFX12 U724 ( .A(n9634), .Y(n141) );
  AO22X1 U725 ( .A0(mem_rdata_I[52]), .A1(n5540), .B0(n252), .B1(n11238), .Y(
        n9634) );
  INVX3 U726 ( .A(net112286), .Y(n142) );
  INVX3 U727 ( .A(net112286), .Y(n143) );
  INVX1 U728 ( .A(net128157), .Y(n144) );
  INVX1 U729 ( .A(n144), .Y(n145) );
  INVX16 U730 ( .A(n142), .Y(n146) );
  INVX20 U731 ( .A(n146), .Y(n147) );
  INVX20 U732 ( .A(n146), .Y(n148) );
  INVX12 U733 ( .A(n143), .Y(n149) );
  INVX20 U734 ( .A(n149), .Y(n150) );
  INVX16 U735 ( .A(n149), .Y(n151) );
  AND2X1 U736 ( .A(n402), .B(n4504), .Y(net128157) );
  BUFX6 U737 ( .A(net128157), .Y(net112286) );
  OA22X2 U738 ( .A0(n4993), .A1(n756), .B0(n5034), .B1(n2317), .Y(n6343) );
  BUFX16 U739 ( .A(n3840), .Y(n5034) );
  CLKAND2X12 U740 ( .A(net98707), .B(net98708), .Y(net128955) );
  INVX8 U741 ( .A(n6530), .Y(n6544) );
  AOI222X4 U742 ( .A0(n5512), .A1(n11386), .B0(mem_rdata_D[36]), .B1(n233), 
        .C0(n12983), .C1(n5507), .Y(n10976) );
  INVX4 U743 ( .A(n11386), .Y(n10975) );
  NAND4X4 U744 ( .A(n6895), .B(n6894), .C(n6893), .D(n6892), .Y(n11386) );
  NAND2X8 U745 ( .A(\i_MIPS/ALUin1[14] ), .B(n6555), .Y(n7617) );
  CLKINVX8 U746 ( .A(n6576), .Y(n6555) );
  OA22X2 U747 ( .A0(n5302), .A1(n1636), .B0(n5256), .B1(n3218), .Y(n9963) );
  CLKBUFX4 U748 ( .A(n5305), .Y(n5302) );
  INVX4 U749 ( .A(n3926), .Y(net97574) );
  CLKBUFX8 U750 ( .A(n5400), .Y(n5398) );
  CLKBUFX20 U751 ( .A(n5400), .Y(n5399) );
  CLKBUFX12 U752 ( .A(n5400), .Y(n5397) );
  BUFX4 U753 ( .A(n5398), .Y(n5377) );
  BUFX4 U754 ( .A(n5398), .Y(n5378) );
  CLKBUFX3 U755 ( .A(n5398), .Y(n5379) );
  CLKBUFX4 U756 ( .A(n5399), .Y(n237) );
  CLKBUFX4 U757 ( .A(n5399), .Y(n5373) );
  CLKBUFX2 U758 ( .A(n5399), .Y(n5375) );
  CLKBUFX2 U759 ( .A(n5399), .Y(n5372) );
  CLKBUFX2 U760 ( .A(n5397), .Y(n5382) );
  CLKBUFX4 U761 ( .A(n5399), .Y(n5374) );
  CLKBUFX6 U762 ( .A(n5397), .Y(n5381) );
  BUFX20 U763 ( .A(n5397), .Y(n5380) );
  CLKBUFX2 U764 ( .A(n5394), .Y(n5393) );
  BUFX20 U765 ( .A(n5401), .Y(n5395) );
  BUFX20 U766 ( .A(n5399), .Y(n5371) );
  BUFX12 U767 ( .A(n5401), .Y(n5396) );
  BUFX6 U768 ( .A(n5398), .Y(n5376) );
  BUFX4 U769 ( .A(n5392), .Y(n5370) );
  CLKBUFX8 U770 ( .A(n5392), .Y(n5368) );
  CLKBUFX4 U771 ( .A(n5395), .Y(n5387) );
  CLKBUFX4 U772 ( .A(n5395), .Y(n5389) );
  BUFX16 U773 ( .A(n5396), .Y(n5385) );
  CLKBUFX6 U774 ( .A(n5396), .Y(n5386) );
  CLKBUFX8 U775 ( .A(n5396), .Y(n5383) );
  NAND2X8 U776 ( .A(n9559), .B(\i_MIPS/IF_ID[97] ), .Y(net97592) );
  BUFX12 U777 ( .A(n6226), .Y(n152) );
  AO22X1 U778 ( .A0(mem_rdata_I[93]), .A1(n5542), .B0(n252), .B1(n11279), .Y(
        n6226) );
  BUFX12 U779 ( .A(n9678), .Y(n153) );
  AO22X1 U780 ( .A0(mem_rdata_I[18]), .A1(n5540), .B0(n251), .B1(n11204), .Y(
        n9678) );
  BUFX12 U781 ( .A(n6196), .Y(n154) );
  AO22X1 U782 ( .A0(mem_rdata_I[63]), .A1(n5542), .B0(n251), .B1(n11249), .Y(
        n6196) );
  BUFX12 U783 ( .A(n9673), .Y(n155) );
  AO22X1 U784 ( .A0(mem_rdata_I[82]), .A1(n5540), .B0(n253), .B1(n11268), .Y(
        n9673) );
  OAI2BB2X1 U785 ( .B0(net108192), .B1(\i_MIPS/n328 ), .A0N(n4073), .A1N(n9566), .Y(\i_MIPS/N87 ) );
  OAI2BB2X1 U786 ( .B0(\i_MIPS/n236 ), .B1(net108190), .A0N(n11041), .A1N(
        n4073), .Y(\i_MIPS/N90 ) );
  BUFX12 U787 ( .A(n9813), .Y(n156) );
  AO22X1 U788 ( .A0(mem_rdata_I[89]), .A1(n5540), .B0(n252), .B1(n11275), .Y(
        n9813) );
  BUFX12 U789 ( .A(n6171), .Y(n157) );
  AO22X1 U790 ( .A0(mem_rdata_I[28]), .A1(n5542), .B0(n250), .B1(n11214), .Y(
        n6171) );
  NAND2X8 U791 ( .A(n11081), .B(n11078), .Y(n10177) );
  BUFX12 U792 ( .A(n9629), .Y(n158) );
  AO22X1 U793 ( .A0(mem_rdata_I[20]), .A1(n5540), .B0(n251), .B1(n11206), .Y(
        n9629) );
  BUFX12 U794 ( .A(n6181), .Y(n159) );
  AO22X1 U795 ( .A0(mem_rdata_I[127]), .A1(n5542), .B0(n249), .B1(n11313), .Y(
        n6181) );
  BUFX12 U796 ( .A(n9788), .Y(n160) );
  AO22X1 U797 ( .A0(mem_rdata_I[120]), .A1(n5540), .B0(n253), .B1(n11306), .Y(
        n9788) );
  BUFX12 U798 ( .A(n6206), .Y(n161) );
  AO22X1 U799 ( .A0(mem_rdata_I[94]), .A1(n5542), .B0(n251), .B1(n11280), .Y(
        n6206) );
  AOI2BB2X2 U800 ( .B0(n2649), .B1(net108664), .A0N(n10470), .A1N(net133585), 
        .Y(n10471) );
  CLKINVX16 U801 ( .A(n3921), .Y(net133585) );
  BUFX12 U802 ( .A(n9683), .Y(n162) );
  AO22X1 U803 ( .A0(mem_rdata_I[50]), .A1(n5540), .B0(n250), .B1(n11236), .Y(
        n9683) );
  BUFX12 U804 ( .A(n9668), .Y(n163) );
  AO22X1 U805 ( .A0(mem_rdata_I[114]), .A1(n5540), .B0(n253), .B1(n11300), .Y(
        n9668) );
  BUFX12 U806 ( .A(n6191), .Y(n164) );
  AO22X1 U807 ( .A0(mem_rdata_I[31]), .A1(n5542), .B0(n251), .B1(n11217), .Y(
        n6191) );
  BUFX12 U808 ( .A(n6186), .Y(n165) );
  AO22X1 U809 ( .A0(mem_rdata_I[95]), .A1(n5542), .B0(n253), .B1(n11281), .Y(
        n6186) );
  BUFX4 U810 ( .A(n10147), .Y(n166) );
  MXI2X1 U811 ( .A(n10146), .B(n10145), .S0(n5513), .Y(n10147) );
  AOI22X4 U812 ( .A0(\i_MIPS/IF_ID[95] ), .A1(n3930), .B0(n10795), .B1(
        net108664), .Y(n3932) );
  AO22X4 U813 ( .A0(mem_rdata_I[17]), .A1(n5536), .B0(n249), .B1(n11203), .Y(
        n10167) );
  BUFX6 U814 ( .A(n5529), .Y(n5536) );
  INVX2 U815 ( .A(n10629), .Y(n10626) );
  XOR3X4 U816 ( .A(net112400), .B(n10627), .C(n10625), .Y(n10629) );
  OAI21X2 U817 ( .A0(\i_MIPS/n238 ), .A1(net108190), .B0(n10529), .Y(
        \i_MIPS/N92 ) );
  OAI2BB2X2 U818 ( .B0(\i_MIPS/n203 ), .B1(net108198), .A0N(n4300), .A1N(n4072), .Y(\i_MIPS/N46 ) );
  NAND2X1 U819 ( .A(n4300), .B(net97874), .Y(n10540) );
  XNOR2X4 U820 ( .A(n10225), .B(ICACHE_addr[18]), .Y(n4300) );
  BUFX12 U821 ( .A(n10191), .Y(n167) );
  NAND3BX2 U822 ( .AN(n4661), .B(n3783), .C(n224), .Y(n10191) );
  CLKBUFX12 U823 ( .A(n12789), .Y(mem_addr_D[29]) );
  CLKINVX1 U824 ( .A(n4624), .Y(n12789) );
  BUFX4 U825 ( .A(n10895), .Y(n169) );
  MXI2X1 U826 ( .A(n10894), .B(n10893), .S0(n5520), .Y(n10895) );
  CLKAND2X12 U827 ( .A(mem_write_I), .B(n11240), .Y(mem_wdata_I[54]) );
  BUFX20 U828 ( .A(n4002), .Y(mem_wdata_I[72]) );
  BUFX4 U829 ( .A(n12870), .Y(n4002) );
  BUFX20 U830 ( .A(n4009), .Y(mem_wdata_I[78]) );
  BUFX4 U831 ( .A(n12864), .Y(n4009) );
  BUFX20 U832 ( .A(n4015), .Y(mem_wdata_I[84]) );
  BUFX4 U833 ( .A(n12858), .Y(n4015) );
  BUFX20 U834 ( .A(n4018), .Y(mem_wdata_I[87]) );
  BUFX4 U835 ( .A(n12855), .Y(n4018) );
  BUFX20 U836 ( .A(n4027), .Y(mem_wdata_I[96]) );
  BUFX4 U837 ( .A(n12846), .Y(n4027) );
  BUFX20 U838 ( .A(n4033), .Y(mem_wdata_I[102]) );
  BUFX4 U839 ( .A(n12841), .Y(n4033) );
  BUFX20 U840 ( .A(n4036), .Y(mem_wdata_I[105]) );
  BUFX4 U841 ( .A(n12838), .Y(n4036) );
  BUFX20 U842 ( .A(n4042), .Y(mem_wdata_I[114]) );
  BUFX4 U843 ( .A(n12832), .Y(n4042) );
  BUFX20 U844 ( .A(n4045), .Y(mem_wdata_I[117]) );
  BUFX4 U845 ( .A(n12829), .Y(n4045) );
  BUFX20 U846 ( .A(n4048), .Y(mem_wdata_I[120]) );
  BUFX4 U847 ( .A(n12826), .Y(n4048) );
  BUFX12 U848 ( .A(n5531), .Y(n5537) );
  BUFX12 U849 ( .A(n9919), .Y(n180) );
  AO22X1 U850 ( .A0(mem_rdata_I[69]), .A1(n5537), .B0(n251), .B1(n11255), .Y(
        n9919) );
  INVX20 U851 ( .A(net108680), .Y(net108676) );
  OAI32X4 U852 ( .A0(n10858), .A1(n10790), .A2(net138000), .B0(\i_MIPS/PC/n31 ), .B1(net97444), .Y(n10583) );
  NAND3BX2 U853 ( .AN(n10358), .B(net97592), .C(n10372), .Y(n10858) );
  INVXL U854 ( .A(net97444), .Y(net138000) );
  NAND2X2 U855 ( .A(n10316), .B(ICACHE_addr[23]), .Y(n10284) );
  AOI2BB2X4 U856 ( .B0(\i_MIPS/IF_ID[73] ), .B1(n3930), .A0N(net108674), .A1N(
        \i_MIPS/n191 ), .Y(n10380) );
  AOI2BB2X4 U857 ( .B0(\i_MIPS/IF_ID[66] ), .B1(n3930), .A0N(net108674), .A1N(
        \i_MIPS/n184 ), .Y(n10528) );
  BUFX20 U858 ( .A(n4140), .Y(n3930) );
  OAI222X2 U859 ( .A0(\i_MIPS/PC/n12 ), .A1(net108688), .B0(n3637), .B1(n10816), .C0(n4430), .C1(net108702), .Y(n10821) );
  OAI222X1 U860 ( .A0(\i_MIPS/PC/n13 ), .A1(net108688), .B0(n3637), .B1(n10595), .C0(n4396), .C1(net108704), .Y(n10600) );
  OAI222X2 U861 ( .A0(\i_MIPS/PC/n23 ), .A1(net108690), .B0(n3637), .B1(n11123), .C0(n4427), .C1(net108702), .Y(n11129) );
  OAI222X1 U862 ( .A0(n10176), .A1(net108686), .B0(n3637), .B1(n4301), .C0(
        net129005), .C1(net108702), .Y(n11072) );
  NAND2BX4 U863 ( .AN(n3637), .B(n409), .Y(n4221) );
  BUFX3 U864 ( .A(n5084), .Y(n181) );
  BUFX16 U865 ( .A(n167), .Y(n5089) );
  BUFX20 U866 ( .A(n167), .Y(n5088) );
  BUFX20 U867 ( .A(n5089), .Y(n5081) );
  BUFX12 U868 ( .A(n5088), .Y(n5083) );
  BUFX20 U869 ( .A(n5089), .Y(n5080) );
  BUFX6 U870 ( .A(n5089), .Y(n5086) );
  BUFX20 U871 ( .A(n5088), .Y(n5084) );
  BUFX20 U872 ( .A(n5089), .Y(n5082) );
  CLKBUFX8 U873 ( .A(n5080), .Y(n5077) );
  BUFX20 U874 ( .A(n5080), .Y(n5079) );
  BUFX20 U875 ( .A(n5088), .Y(n5087) );
  BUFX20 U876 ( .A(n5075), .Y(n5054) );
  BUFX4 U877 ( .A(n5086), .Y(n5058) );
  BUFX6 U878 ( .A(n5081), .Y(n5076) );
  BUFX20 U879 ( .A(n5085), .Y(n5063) );
  BUFX6 U880 ( .A(n5083), .Y(n5070) );
  CLKBUFX6 U881 ( .A(n5081), .Y(n5074) );
  BUFX6 U882 ( .A(n5086), .Y(n5059) );
  BUFX8 U883 ( .A(n5083), .Y(n5069) );
  CLKBUFX6 U884 ( .A(n5080), .Y(n5078) );
  BUFX4 U885 ( .A(n5083), .Y(n5068) );
  BUFX20 U886 ( .A(n5084), .Y(n5066) );
  CLKBUFX4 U887 ( .A(n5084), .Y(n5064) );
  CLKBUFX4 U888 ( .A(n5084), .Y(n5067) );
  BUFX20 U889 ( .A(n5084), .Y(n5065) );
  BUFX20 U890 ( .A(n5087), .Y(n5057) );
  CLKBUFX4 U891 ( .A(n5087), .Y(n5055) );
  CLKBUFX6 U892 ( .A(n5081), .Y(n5073) );
  BUFX20 U893 ( .A(n5082), .Y(n5072) );
  BUFX20 U894 ( .A(n5082), .Y(n5071) );
  CLKINVX3 U895 ( .A(n5054), .Y(n5053) );
  CLKINVX3 U896 ( .A(n5056), .Y(n5051) );
  CLKINVX3 U897 ( .A(n5057), .Y(n5049) );
  CLKINVX3 U898 ( .A(n5071), .Y(n5046) );
  CLKINVX3 U899 ( .A(n5071), .Y(n5050) );
  BUFX4 U900 ( .A(n10955), .Y(n182) );
  MXI2X1 U901 ( .A(n10954), .B(n10953), .S0(n5522), .Y(n10955) );
  OA22XL U902 ( .A0(n5382), .A1(n1086), .B0(n5333), .B1(n2680), .Y(n6167) );
  OA22XL U903 ( .A0(n269), .A1(n1537), .B0(n5335), .B1(n3119), .Y(n6240) );
  OA22XL U904 ( .A0(n5399), .A1(n1488), .B0(n5350), .B1(n3072), .Y(n9910) );
  BUFX16 U905 ( .A(n269), .Y(n5400) );
  BUFX20 U906 ( .A(n269), .Y(n5401) );
  BUFX8 U907 ( .A(n5158), .Y(n183) );
  AO22X4 U908 ( .A0(mem_rdata_I[51]), .A1(n5535), .B0(n253), .B1(n11237), .Y(
        n11119) );
  BUFX6 U909 ( .A(n5529), .Y(n5535) );
  XOR2X4 U910 ( .A(n10452), .B(n10456), .Y(n10453) );
  NAND3BX4 U911 ( .AN(n11101), .B(n11100), .C(n11099), .Y(\i_MIPS/PC/n40 ) );
  OA22X2 U912 ( .A0(n11098), .A1(net133585), .B0(n11097), .B1(net108658), .Y(
        n11099) );
  CLKINVX4 U913 ( .A(n10533), .Y(n10256) );
  XNOR2X4 U914 ( .A(n10255), .B(net112404), .Y(n10533) );
  CLKINVX8 U915 ( .A(n5021), .Y(n184) );
  INVX12 U916 ( .A(n184), .Y(n185) );
  AO22X4 U917 ( .A0(n5543), .A1(ICACHE_addr[19]), .B0(n239), .B1(n11334), .Y(
        n11131) );
  NAND4X4 U918 ( .A(n5980), .B(n5979), .C(n5978), .D(n5977), .Y(n11334) );
  AO22X4 U919 ( .A0(mem_rdata_I[75]), .A1(n5539), .B0(n252), .B1(n11261), .Y(
        n9746) );
  BUFX16 U920 ( .A(n5530), .Y(n5539) );
  CLKMX2X6 U921 ( .A(\i_MIPS/n299 ), .B(net127930), .S0(n5624), .Y(n6535) );
  NAND2BX4 U922 ( .AN(n8266), .B(n8861), .Y(n8267) );
  NAND2X2 U923 ( .A(net112294), .B(n8238), .Y(n8266) );
  AOI22X2 U924 ( .A0(net111910), .A1(n6747), .B0(net111962), .B1(n6679), .Y(
        n4457) );
  NAND2X6 U925 ( .A(n10137), .B(n10136), .Y(n6747) );
  NAND2X4 U926 ( .A(n6562), .B(\i_MIPS/n358 ), .Y(n7693) );
  INVX8 U927 ( .A(n6547), .Y(n6562) );
  NAND2X4 U928 ( .A(n10569), .B(ICACHE_addr[25]), .Y(n10343) );
  INVX4 U929 ( .A(n10342), .Y(n10569) );
  AOI2BB2X2 U930 ( .B0(\i_MIPS/IF_ID[89] ), .B1(n3930), .A0N(net108674), .A1N(
        \i_MIPS/n207 ), .Y(n10461) );
  AOI2BB2X2 U931 ( .B0(\i_MIPS/IF_ID[88] ), .B1(n3930), .A0N(net108674), .A1N(
        \i_MIPS/n206 ), .Y(n4144) );
  AOI2BB2X2 U932 ( .B0(\i_MIPS/IF_ID[80] ), .B1(n3930), .A0N(net108674), .A1N(
        \i_MIPS/n198 ), .Y(n10429) );
  AOI2BB2X2 U933 ( .B0(\i_MIPS/IF_ID[86] ), .B1(n3930), .A0N(net108678), .A1N(
        \i_MIPS/n204 ), .Y(n11128) );
  AOI2BB2X2 U934 ( .B0(\i_MIPS/IF_ID[82] ), .B1(n3930), .A0N(net108674), .A1N(
        \i_MIPS/n200 ), .Y(n10442) );
  AOI2BB2X2 U935 ( .B0(\i_MIPS/IF_ID[92] ), .B1(n3930), .A0N(net108676), .A1N(
        \i_MIPS/n210 ), .Y(n10844) );
  AOI2BB2X2 U936 ( .B0(\i_MIPS/IF_ID[84] ), .B1(n3930), .A0N(net108676), .A1N(
        \i_MIPS/n202 ), .Y(n10648) );
  AOI2BB2X2 U937 ( .B0(\i_MIPS/IF_ID[91] ), .B1(n3930), .A0N(net108676), .A1N(
        \i_MIPS/n209 ), .Y(n10833) );
  AOI2BB2X2 U938 ( .B0(\i_MIPS/IF_ID[85] ), .B1(n3930), .A0N(net108674), .A1N(
        \i_MIPS/n203 ), .Y(n10536) );
  AOI2BB2X2 U939 ( .B0(\i_MIPS/IF_ID[79] ), .B1(n3930), .A0N(net108674), .A1N(
        \i_MIPS/n197 ), .Y(n10414) );
  OR2XL U940 ( .A(n4649), .B(n10744), .Y(n3719) );
  INVX3 U941 ( .A(n11428), .Y(n10744) );
  INVXL U942 ( .A(n9532), .Y(n186) );
  INVXL U943 ( .A(n4719), .Y(n187) );
  INVXL U944 ( .A(n4719), .Y(n188) );
  INVXL U945 ( .A(n4719), .Y(n189) );
  INVX8 U946 ( .A(n9413), .Y(n9532) );
  BUFX20 U947 ( .A(n9532), .Y(n4718) );
  BUFX20 U948 ( .A(n4718), .Y(n4719) );
  NAND2X6 U949 ( .A(n7688), .B(n7693), .Y(n7164) );
  NOR2X6 U950 ( .A(n7223), .B(n3343), .Y(n7166) );
  CLKAND2X12 U951 ( .A(n6546), .B(n3343), .Y(n4388) );
  AND2X6 U952 ( .A(n7880), .B(n8635), .Y(n3343) );
  NAND3BX2 U953 ( .AN(n7802), .B(n7801), .C(net111994), .Y(n7835) );
  BUFX8 U954 ( .A(n10913), .Y(n190) );
  INVX8 U955 ( .A(net112218), .Y(n191) );
  CLKINVX16 U956 ( .A(n191), .Y(n192) );
  CLKINVX4 U957 ( .A(net112232), .Y(net112218) );
  AOI21X2 U958 ( .A0(n8174), .A1(n9350), .B0(n8173), .Y(n4425) );
  CLKBUFX8 U959 ( .A(n4929), .Y(n4916) );
  INVX8 U960 ( .A(net112214), .Y(n193) );
  CLKINVX2 U961 ( .A(net128161), .Y(n194) );
  CLKINVX1 U962 ( .A(n194), .Y(n195) );
  CLKINVX16 U963 ( .A(n193), .Y(n196) );
  INVX20 U964 ( .A(n196), .Y(n197) );
  INVX16 U965 ( .A(n196), .Y(n198) );
  INVX12 U966 ( .A(n196), .Y(n199) );
  INVX16 U967 ( .A(n196), .Y(n200) );
  AND2X1 U968 ( .A(n4521), .B(n4504), .Y(net128161) );
  BUFX6 U969 ( .A(net128161), .Y(net112214) );
  BUFX6 U970 ( .A(n9280), .Y(n4251) );
  NAND2X2 U971 ( .A(\i_MIPS/ALUin1[26] ), .B(n261), .Y(n8948) );
  BUFX8 U972 ( .A(n6591), .Y(n261) );
  AND4X6 U973 ( .A(n9287), .B(n9285), .C(n9286), .D(n9284), .Y(n3913) );
  CLKMX2X4 U974 ( .A(\i_MIPS/n283 ), .B(n4538), .S0(n5622), .Y(n6547) );
  CLKMX2X4 U975 ( .A(n8438), .B(n9250), .S0(net107796), .Y(n8261) );
  NAND2X4 U976 ( .A(net105676), .B(\i_MIPS/n369 ), .Y(net102430) );
  OA22XL U977 ( .A0(n4750), .A1(n796), .B0(n4791), .B1(n2359), .Y(n8191) );
  OA22X1 U978 ( .A0(n4750), .A1(n2969), .B0(n4791), .B1(n1195), .Y(n8103) );
  OA22X1 U979 ( .A0(n4750), .A1(n805), .B0(n4791), .B1(n2368), .Y(n8024) );
  BUFX2 U980 ( .A(n4769), .Y(n4750) );
  BUFX16 U981 ( .A(n5305), .Y(n5304) );
  OA22X4 U982 ( .A0(n4979), .A1(n2094), .B0(n5024), .B1(n507), .Y(n7650) );
  CLKBUFX12 U983 ( .A(n4992), .Y(n4979) );
  BUFX2 U984 ( .A(n4837), .Y(n4823) );
  OA22X4 U985 ( .A0(n5384), .A1(n1713), .B0(n5331), .B1(n3310), .Y(n6132) );
  BUFX8 U986 ( .A(n5392), .Y(n5369) );
  OAI2BB2X1 U987 ( .B0(\i_MIPS/n167 ), .B1(net108192), .A0N(n4073), .A1N(
        n10614), .Y(\i_MIPS/N107 ) );
  CLKINVX4 U988 ( .A(n10616), .Y(n10614) );
  INVX8 U989 ( .A(n11435), .Y(n10670) );
  NAND4X4 U990 ( .A(n9187), .B(n9186), .C(n9185), .D(n9184), .Y(n11435) );
  AOI33X2 U991 ( .A0(n8859), .A1(n8871), .A2(net112292), .B0(n8858), .B1(n8857), .B2(net137952), .Y(net101555) );
  NAND4X2 U992 ( .A(n8502), .B(n8501), .C(n8500), .D(n8499), .Y(n11410) );
  OA22X2 U993 ( .A0(n4972), .A1(n2130), .B0(n5017), .B1(n544), .Y(n8499) );
  INVXL U994 ( .A(net97410), .Y(n201) );
  INVX4 U995 ( .A(n201), .Y(n202) );
  INVX16 U996 ( .A(net108118), .Y(n203) );
  CLKINVX16 U997 ( .A(n203), .Y(n204) );
  CLKINVX16 U998 ( .A(n203), .Y(n205) );
  INVX16 U999 ( .A(net108108), .Y(n206) );
  CLKINVX16 U1000 ( .A(n206), .Y(n207) );
  CLKINVX16 U1001 ( .A(n206), .Y(n208) );
  INVX8 U1002 ( .A(net108098), .Y(n209) );
  CLKINVX12 U1003 ( .A(n209), .Y(n210) );
  CLKINVX12 U1004 ( .A(n209), .Y(n211) );
  INVX12 U1005 ( .A(net108112), .Y(n212) );
  CLKINVX12 U1006 ( .A(n212), .Y(n213) );
  CLKINVX12 U1007 ( .A(n212), .Y(n214) );
  INVX16 U1008 ( .A(net108110), .Y(n215) );
  CLKINVX16 U1009 ( .A(n215), .Y(n216) );
  CLKINVX16 U1010 ( .A(n215), .Y(n217) );
  INVX20 U1011 ( .A(net108116), .Y(n218) );
  INVX12 U1012 ( .A(n218), .Y(n219) );
  INVX20 U1013 ( .A(n218), .Y(n220) );
  INVX16 U1014 ( .A(net108114), .Y(n221) );
  CLKINVX16 U1015 ( .A(n221), .Y(n222) );
  CLKINVX16 U1016 ( .A(n221), .Y(n223) );
  CLKINVX1 U1017 ( .A(net108156), .Y(net108118) );
  CLKINVX3 U1018 ( .A(net108154), .Y(net108108) );
  INVX1 U1019 ( .A(net108156), .Y(net108112) );
  CLKINVX1 U1020 ( .A(net108132), .Y(net108110) );
  CLKINVX1 U1021 ( .A(net108126), .Y(net108116) );
  CLKINVX1 U1022 ( .A(net108128), .Y(net108114) );
  NAND3BX2 U1023 ( .AN(n11009), .B(n4060), .C(n9568), .Y(net97410) );
  BUFX12 U1024 ( .A(net97410), .Y(net108160) );
  BUFX4 U1025 ( .A(net108160), .Y(net108154) );
  BUFX20 U1026 ( .A(net108160), .Y(net108156) );
  BUFX8 U1027 ( .A(net108154), .Y(net108132) );
  BUFX16 U1028 ( .A(net108156), .Y(net108126) );
  CLKINVX3 U1029 ( .A(n3785), .Y(n3786) );
  AOI2BB2X2 U1030 ( .B0(\i_MIPS/IF_ID[71] ), .B1(net108670), .A0N(net108678), 
        .A1N(\i_MIPS/n189 ), .Y(n11100) );
  NAND2X2 U1031 ( .A(n8237), .B(n8236), .Y(net102573) );
  NAND2X2 U1032 ( .A(n6564), .B(\i_MIPS/n347 ), .Y(n8237) );
  OA22X4 U1033 ( .A0(n5120), .A1(n1614), .B0(n5074), .B1(n3191), .Y(n9937) );
  BUFX12 U1034 ( .A(n5125), .Y(n5120) );
  NOR2X8 U1035 ( .A(n6351), .B(n6352), .Y(n6367) );
  OA22X1 U1036 ( .A0(n5124), .A1(n1682), .B0(n5070), .B1(n3273), .Y(n10186) );
  OA22X4 U1037 ( .A0(n5105), .A1(n1660), .B0(n5067), .B1(n3244), .Y(n6150) );
  OA22X4 U1038 ( .A0(n5105), .A1(n1677), .B0(n181), .B1(n3267), .Y(n6140) );
  OA22X4 U1039 ( .A0(n5105), .A1(n1658), .B0(n5067), .B1(n3242), .Y(n6145) );
  OA22X2 U1040 ( .A0(n5105), .A1(n1618), .B0(n5078), .B1(n3195), .Y(n6160) );
  OA22X4 U1041 ( .A0(n5105), .A1(n1459), .B0(n5073), .B1(n3033), .Y(n6155) );
  OA22X1 U1042 ( .A0(n5105), .A1(n1621), .B0(n5064), .B1(n3198), .Y(n6165) );
  OA22X4 U1043 ( .A0(n5124), .A1(n1683), .B0(n5069), .B1(n3274), .Y(n10182) );
  CLKBUFX6 U1044 ( .A(n5125), .Y(n5124) );
  BUFX6 U1045 ( .A(n5530), .Y(n5542) );
  OA22X4 U1046 ( .A0(n5120), .A1(n1611), .B0(n5061), .B1(n3188), .Y(n9945) );
  BUFX20 U1047 ( .A(n5081), .Y(n5075) );
  NAND2X8 U1048 ( .A(n7520), .B(n7527), .Y(n7797) );
  AND2X1 U1049 ( .A(n5557), .B(n11187), .Y(n12927) );
  NAND4X4 U1050 ( .A(n9961), .B(n9960), .C(n9959), .D(n9958), .Y(n11187) );
  INVX6 U1051 ( .A(n11319), .Y(n11512) );
  BUFX12 U1052 ( .A(n11512), .Y(mem_read_I) );
  NAND3BX4 U1053 ( .AN(n11316), .B(n11315), .C(n11314), .Y(n11319) );
  AOI2BB2X2 U1054 ( .B0(\i_MIPS/IF_ID[76] ), .B1(n3930), .A0N(net108676), 
        .A1N(\i_MIPS/n194 ), .Y(n10599) );
  NAND3BX4 U1055 ( .AN(n10473), .B(n10472), .C(n10471), .Y(\i_MIPS/PC/n59 ) );
  AOI2BB2X2 U1056 ( .B0(\i_MIPS/IF_ID[90] ), .B1(n3930), .A0N(net108674), 
        .A1N(\i_MIPS/n208 ), .Y(n10472) );
  INVX8 U1057 ( .A(n11422), .Y(n10896) );
  NAND4X6 U1058 ( .A(n7096), .B(n7095), .C(n7094), .D(n7093), .Y(n11422) );
  INVX1 U1059 ( .A(net112258), .Y(n226) );
  INVX8 U1060 ( .A(net112260), .Y(n227) );
  INVX2 U1061 ( .A(net112254), .Y(n228) );
  INVX1 U1062 ( .A(net112258), .Y(n229) );
  CLKINVX12 U1063 ( .A(net112268), .Y(net112254) );
  CLKINVX12 U1064 ( .A(net112264), .Y(net112260) );
  CLKINVX12 U1065 ( .A(net112266), .Y(net112258) );
  AND2X1 U1066 ( .A(n402), .B(n4446), .Y(net128156) );
  BUFX4 U1067 ( .A(net128156), .Y(net112264) );
  BUFX4 U1068 ( .A(net128156), .Y(net112268) );
  AOI222XL U1069 ( .A0(n5503), .A1(n11351), .B0(mem_rdata_D[1]), .B1(n233), 
        .C0(n12986), .C1(n5502), .Y(n10912) );
  INVX8 U1070 ( .A(n11351), .Y(n10911) );
  NAND4X4 U1071 ( .A(n8020), .B(n8019), .C(n8018), .D(n8017), .Y(n11351) );
  NAND2X2 U1072 ( .A(net108664), .B(n4424), .Y(n10582) );
  XNOR3X2 U1073 ( .A(net112400), .B(n10791), .C(n10792), .Y(n4424) );
  OAI2BB2X4 U1074 ( .B0(\i_MIPS/n171 ), .B1(net108198), .A0N(n4072), .A1N(
        n10256), .Y(\i_MIPS/N111 ) );
  OAI222X4 U1075 ( .A0(n224), .A1(net108688), .B0(net97445), .B1(n11096), .C0(
        n4406), .C1(net108702), .Y(n11101) );
  OAI2BB2X4 U1076 ( .B0(\i_MIPS/n175 ), .B1(net108194), .A0N(n4073), .A1N(
        n10454), .Y(\i_MIPS/N115 ) );
  CLKINVX3 U1077 ( .A(n10458), .Y(n10454) );
  OAI2BB2X4 U1078 ( .B0(\i_MIPS/n181 ), .B1(net108192), .A0N(n10795), .A1N(
        n4315), .Y(\i_MIPS/N121 ) );
  NAND3BX2 U1079 ( .AN(n10600), .B(n10598), .C(n10599), .Y(\i_MIPS/PC/n45 ) );
  NOR2X4 U1080 ( .A(n7158), .B(n7157), .Y(n7170) );
  CLKINVX3 U1081 ( .A(n10426), .Y(n10424) );
  OAI2BB2X2 U1082 ( .B0(\i_MIPS/n169 ), .B1(net108192), .A0N(n5545), .A1N(
        n10626), .Y(\i_MIPS/N109 ) );
  CLKAND2X12 U1083 ( .A(n6518), .B(n4468), .Y(n4436) );
  NAND2X6 U1084 ( .A(n6518), .B(n9140), .Y(n8229) );
  CLKINVX8 U1085 ( .A(n9139), .Y(n6518) );
  NAND3BX4 U1086 ( .AN(n11072), .B(n11071), .C(n11070), .Y(\i_MIPS/PC/n36 ) );
  OA22X2 U1087 ( .A0(n11069), .A1(net133585), .B0(net108658), .B1(n11068), .Y(
        n11070) );
  AOI2BB2X2 U1088 ( .B0(\i_MIPS/IF_ID[67] ), .B1(net108670), .A0N(net108676), 
        .A1N(\i_MIPS/n185 ), .Y(n11071) );
  AOI21X4 U1089 ( .A0(n6546), .A1(n7223), .B0(n7163), .Y(n4433) );
  INVX8 U1090 ( .A(n7167), .Y(n6546) );
  NAND2X8 U1091 ( .A(n8636), .B(n8631), .Y(n7223) );
  BUFX16 U1092 ( .A(n5294), .Y(n230) );
  BUFX3 U1093 ( .A(n5307), .Y(n5294) );
  OA22X2 U1094 ( .A0(n10597), .A1(net133585), .B0(n10596), .B1(net108660), .Y(
        n10598) );
  XOR3X2 U1095 ( .A(n10593), .B(n10592), .C(n10591), .Y(n10596) );
  INVX8 U1096 ( .A(n10790), .Y(n10791) );
  NAND2XL U1097 ( .A(net112400), .B(n10790), .Y(n10853) );
  XOR2X4 U1098 ( .A(n10793), .B(ICACHE_addr[27]), .Y(n10790) );
  CLKMX2X8 U1099 ( .A(\i_MIPS/n281 ), .B(n4540), .S0(n5622), .Y(n6576) );
  MXI2X1 U1100 ( .A(\i_MIPS/n280 ), .B(\i_MIPS/n281 ), .S0(n207), .Y(
        \i_MIPS/n408 ) );
  MXI2X2 U1101 ( .A(n10963), .B(n10962), .S0(n5522), .Y(n10964) );
  NAND2X2 U1102 ( .A(n8448), .B(n3899), .Y(n8463) );
  AND2X8 U1103 ( .A(n3910), .B(n8970), .Y(n3899) );
  NAND4X2 U1104 ( .A(n9397), .B(n9396), .C(n9395), .D(n9394), .Y(n11409) );
  OA22X4 U1105 ( .A0(n4997), .A1(n2123), .B0(n5016), .B1(n536), .Y(n9394) );
  OA22XL U1106 ( .A0(n4907), .A1(n1214), .B0(n4947), .B1(n2751), .Y(n9395) );
  XOR2X4 U1107 ( .A(DCACHE_addr[18]), .B(n11496), .Y(n6414) );
  NAND4X4 U1108 ( .A(n6408), .B(n6407), .C(n6406), .D(n6405), .Y(n11496) );
  AOI33X4 U1109 ( .A0(n9150), .A1(n9488), .A2(net112292), .B0(n9149), .B1(
        n9168), .B2(net137952), .Y(n9177) );
  XOR2X4 U1110 ( .A(n6337), .B(n4631), .Y(n3852) );
  NAND2X4 U1111 ( .A(n11011), .B(n11012), .Y(n6337) );
  OAI22X4 U1112 ( .A0(n4836), .A1(n2160), .B0(n4882), .B1(n438), .Y(n3403) );
  BUFX20 U1113 ( .A(n4838), .Y(n4836) );
  NOR4X4 U1114 ( .A(n8171), .B(n8170), .C(n8169), .D(n8168), .Y(n8186) );
  OAI211X2 U1115 ( .A0(n10576), .A1(n10575), .B0(n10574), .C0(n10573), .Y(
        n10578) );
  NAND4X2 U1116 ( .A(n4352), .B(n7652), .C(n7651), .D(n7650), .Y(n11428) );
  MXI2X2 U1117 ( .A(n10261), .B(n10260), .S0(n5514), .Y(n10262) );
  OR2XL U1118 ( .A(n4649), .B(n10260), .Y(n3717) );
  OA22X4 U1119 ( .A0(n10257), .A1(n4676), .B0(n10260), .B1(n4250), .Y(n7361)
         );
  INVX3 U1120 ( .A(n11424), .Y(n10260) );
  CLKINVX8 U1121 ( .A(n6570), .Y(n6559) );
  CLKINVX8 U1122 ( .A(n4082), .Y(n4079) );
  NAND2X8 U1123 ( .A(n3836), .B(net137684), .Y(n4082) );
  INVX8 U1124 ( .A(net103889), .Y(net102428) );
  NAND2X4 U1125 ( .A(net105676), .B(\i_MIPS/ALUin1[2] ), .Y(net103889) );
  INVX20 U1126 ( .A(net102050), .Y(net100603) );
  NAND2X2 U1127 ( .A(n4503), .B(n4447), .Y(net102050) );
  AOI2BB2X4 U1128 ( .B0(net111960), .B1(n8978), .A0N(n3773), .A1N(n3721), .Y(
        n3768) );
  BUFX16 U1129 ( .A(n3893), .Y(n3721) );
  BUFX16 U1130 ( .A(n5126), .Y(n5114) );
  NAND2X1 U1131 ( .A(n10329), .B(ICACHE_addr[19]), .Y(n10330) );
  CLKINVX8 U1132 ( .A(n10328), .Y(n10329) );
  NAND2X4 U1133 ( .A(net105677), .B(\i_MIPS/n369 ), .Y(net102427) );
  INVX4 U1134 ( .A(net105677), .Y(net105676) );
  OA22X4 U1135 ( .A0(n10730), .A1(n4676), .B0(n10733), .B1(n4250), .Y(n7756)
         );
  OR2XL U1136 ( .A(n4649), .B(n10730), .Y(n4609) );
  INVX4 U1137 ( .A(n11459), .Y(n10730) );
  OA22X4 U1138 ( .A0(n4919), .A1(n3355), .B0(n4948), .B1(n1735), .Y(n7651) );
  OA22X4 U1139 ( .A0(n4919), .A1(n2730), .B0(n4948), .B1(n1124), .Y(n7586) );
  OA22X4 U1140 ( .A0(n4919), .A1(n2772), .B0(n4948), .B1(n1201), .Y(n7647) );
  OA22X2 U1141 ( .A0(n4919), .A1(n1365), .B0(n4949), .B1(n2895), .Y(n7265) );
  OA22X2 U1142 ( .A0(n4919), .A1(n1362), .B0(n4948), .B1(n2892), .Y(n7582) );
  OA22X2 U1143 ( .A0(n4919), .A1(n2084), .B0(n4948), .B1(n496), .Y(n7578) );
  CLKBUFX4 U1144 ( .A(n4929), .Y(n4919) );
  XOR2X4 U1145 ( .A(n11334), .B(ICACHE_addr[19]), .Y(n5981) );
  XOR2X4 U1146 ( .A(n11491), .B(n12944), .Y(n6352) );
  NAND4X4 U1147 ( .A(n6346), .B(n6345), .C(n6344), .D(n6343), .Y(n11491) );
  CLKMX2X3 U1148 ( .A(\I_cache/cache[1][33] ), .B(n11073), .S0(n5049), .Y(
        n12522) );
  CLKMX2X3 U1149 ( .A(\I_cache/cache[5][33] ), .B(n11073), .S0(n5228), .Y(
        n12518) );
  CLKMX2X3 U1150 ( .A(\I_cache/cache[4][33] ), .B(n11073), .S0(n5277), .Y(
        n12519) );
  CLKMX2X3 U1151 ( .A(\I_cache/cache[6][33] ), .B(n11073), .S0(n5358), .Y(
        n12517) );
  CLKMX2X3 U1152 ( .A(\I_cache/cache[3][33] ), .B(n11073), .S0(n5139), .Y(
        n12520) );
  CLKMX2X3 U1153 ( .A(\I_cache/cache[0][33] ), .B(n11073), .S0(n5099), .Y(
        n12523) );
  AO22X4 U1154 ( .A0(mem_rdata_I[65]), .A1(n5536), .B0(n253), .B1(n11251), .Y(
        n11073) );
  INVX6 U1155 ( .A(n6329), .Y(n11015) );
  INVX8 U1156 ( .A(n11088), .Y(n10362) );
  INVX3 U1157 ( .A(n10360), .Y(n10204) );
  XOR2X4 U1158 ( .A(n10343), .B(ICACHE_addr[26]), .Y(n10357) );
  NAND2X4 U1159 ( .A(n11015), .B(n11014), .Y(n6332) );
  OAI31X4 U1160 ( .A0(n9483), .A1(n9482), .A2(n9481), .B0(n9480), .Y(n9491) );
  AOI2BB1X4 U1161 ( .A0N(n9482), .A1N(n9479), .B0(n9478), .Y(n9480) );
  INVX12 U1162 ( .A(n10816), .Y(n10814) );
  XOR2X4 U1163 ( .A(n10231), .B(ICACHE_addr[8]), .Y(n10816) );
  CLKINVX12 U1164 ( .A(n11008), .Y(n231) );
  CLKINVX12 U1165 ( .A(n231), .Y(n232) );
  INVX12 U1166 ( .A(n231), .Y(n233) );
  INVX12 U1167 ( .A(n231), .Y(n234) );
  INVX12 U1168 ( .A(n231), .Y(n235) );
  INVX8 U1169 ( .A(n231), .Y(n236) );
  AND2X6 U1170 ( .A(n9982), .B(mem_ready_D), .Y(n11008) );
  AO21X2 U1171 ( .A0(n7689), .A1(n7688), .B0(n7687), .Y(n7691) );
  NAND2X8 U1172 ( .A(n4525), .B(n3784), .Y(n269) );
  BUFX20 U1173 ( .A(n5401), .Y(n5394) );
  BUFX6 U1174 ( .A(n5399), .Y(n5367) );
  CLKBUFX4 U1175 ( .A(n5394), .Y(n5391) );
  CLKBUFX4 U1176 ( .A(n5394), .Y(n5390) );
  BUFX20 U1177 ( .A(n5394), .Y(n5392) );
  BUFX6 U1178 ( .A(n5396), .Y(n5384) );
  CLKINVX4 U1179 ( .A(n5367), .Y(n5366) );
  CLKINVX4 U1180 ( .A(n5371), .Y(n5358) );
  CLKINVX3 U1181 ( .A(n5371), .Y(n5359) );
  CLKINVX3 U1182 ( .A(n5368), .Y(n5363) );
  CLKINVX3 U1183 ( .A(n5369), .Y(n5361) );
  CLKINVX3 U1184 ( .A(n5385), .Y(n5360) );
  CLKINVX3 U1185 ( .A(n5385), .Y(n5364) );
  CLKINVX3 U1186 ( .A(n5386), .Y(n5365) );
  CLKINVX3 U1187 ( .A(n5386), .Y(n5362) );
  NAND2X2 U1188 ( .A(\i_MIPS/ALUin1[28] ), .B(n6593), .Y(n8433) );
  INVX3 U1189 ( .A(n6593), .Y(n6589) );
  MXI2X2 U1190 ( .A(\i_MIPS/ID_EX[69] ), .B(\i_MIPS/ID_EX[101] ), .S0(n5624), 
        .Y(n6593) );
  INVX12 U1191 ( .A(n11123), .Y(n11121) );
  XOR2X4 U1192 ( .A(n10328), .B(ICACHE_addr[19]), .Y(n11123) );
  NAND3X6 U1193 ( .A(n3659), .B(n3660), .C(n10382), .Y(n10399) );
  NAND2X4 U1194 ( .A(n10597), .B(n10595), .Y(n10382) );
  XOR2X4 U1195 ( .A(n10338), .B(ICACHE_addr[23]), .Y(n10468) );
  NAND3X4 U1196 ( .A(ICACHE_addr[22]), .B(ICACHE_addr[21]), .C(net98662), .Y(
        n10338) );
  XOR2X2 U1197 ( .A(n10229), .B(ICACHE_addr[7]), .Y(n10585) );
  NAND2XL U1198 ( .A(n10230), .B(ICACHE_addr[7]), .Y(n10231) );
  XNOR2X4 U1199 ( .A(ICACHE_addr[7]), .B(n11322), .Y(n6009) );
  NAND3BX2 U1200 ( .AN(n11316), .B(n11185), .C(n4651), .Y(n11170) );
  CLKINVX8 U1201 ( .A(n6120), .Y(n11316) );
  INVX12 U1202 ( .A(n6571), .Y(n6558) );
  MX2X8 U1203 ( .A(\i_MIPS/n267 ), .B(n4491), .S0(n4299), .Y(n6571) );
  NAND2X4 U1204 ( .A(net112400), .B(n11123), .Y(n10544) );
  AND2X1 U1205 ( .A(net112400), .B(n10468), .Y(n4467) );
  NAND2X4 U1206 ( .A(net112400), .B(net98497), .Y(n10451) );
  BUFX20 U1207 ( .A(net97496), .Y(net112400) );
  NAND3X2 U1208 ( .A(n4166), .B(n4167), .C(n7152), .Y(n7227) );
  OA22X4 U1209 ( .A0(n4669), .A1(\i_MIPS/n351 ), .B0(n3828), .B1(\i_MIPS/n352 ), .Y(n7152) );
  INVX2 U1210 ( .A(n8232), .Y(n6516) );
  CLKAND2X2 U1211 ( .A(n10431), .B(n10421), .Y(n4386) );
  NAND2X6 U1212 ( .A(n10421), .B(n10609), .Y(n10433) );
  NAND2X4 U1213 ( .A(n10408), .B(n10406), .Y(n10421) );
  AND3X8 U1214 ( .A(n8952), .B(n9040), .C(n8953), .Y(n8954) );
  BUFX20 U1215 ( .A(n12820), .Y(mem_addr_I[15]) );
  BUFX20 U1216 ( .A(n12819), .Y(mem_addr_I[16]) );
  BUFX20 U1217 ( .A(n12818), .Y(mem_addr_I[17]) );
  BUFX20 U1218 ( .A(n12817), .Y(mem_addr_I[18]) );
  BUFX20 U1219 ( .A(n12816), .Y(mem_addr_I[19]) );
  BUFX20 U1220 ( .A(n12815), .Y(mem_addr_I[20]) );
  BUFX20 U1221 ( .A(n12814), .Y(mem_addr_I[21]) );
  BUFX20 U1222 ( .A(n12813), .Y(mem_addr_I[22]) );
  BUFX20 U1223 ( .A(n12812), .Y(mem_addr_I[23]) );
  BUFX20 U1224 ( .A(n12811), .Y(mem_addr_I[24]) );
  BUFX20 U1225 ( .A(n12810), .Y(mem_addr_I[25]) );
  BUFX20 U1226 ( .A(n12809), .Y(mem_addr_I[26]) );
  BUFX20 U1227 ( .A(n12808), .Y(mem_addr_I[27]) );
  BUFX20 U1228 ( .A(n12807), .Y(mem_addr_I[28]) );
  BUFX20 U1229 ( .A(n12806), .Y(mem_addr_I[29]) );
  BUFX20 U1230 ( .A(n12805), .Y(mem_addr_I[30]) );
  BUFX20 U1231 ( .A(n12804), .Y(mem_addr_I[31]) );
  AO22X4 U1232 ( .A0(mem_rdata_I[97]), .A1(n5543), .B0(n251), .B1(n11283), .Y(
        n6136) );
  BUFX20 U1233 ( .A(n5531), .Y(n5543) );
  INVX8 U1234 ( .A(n11155), .Y(n238) );
  INVX20 U1235 ( .A(n238), .Y(n239) );
  CLKINVX12 U1236 ( .A(n238), .Y(n240) );
  NAND2BX4 U1237 ( .AN(n11130), .B(n11315), .Y(n11155) );
  INVX20 U1238 ( .A(n9414), .Y(n9531) );
  INVX8 U1239 ( .A(n6541), .Y(n6539) );
  CLKMX2X6 U1240 ( .A(\i_MIPS/n303 ), .B(net105783), .S0(n5623), .Y(n6541) );
  OAI221X2 U1241 ( .A0(net112366), .A1(net103561), .B0(net112348), .B1(
        \i_MIPS/n361 ), .C0(n7418), .Y(n8069) );
  OA22X2 U1242 ( .A0(n4669), .A1(\i_MIPS/n360 ), .B0(n3828), .B1(\i_MIPS/n359 ), .Y(n7418) );
  OA22X2 U1243 ( .A0(n8551), .A1(net101914), .B0(n9334), .B1(net133688), .Y(
        n8365) );
  BUFX8 U1244 ( .A(net98046), .Y(n241) );
  INVX4 U1245 ( .A(n241), .Y(net103417) );
  NAND2X8 U1246 ( .A(n4498), .B(n7975), .Y(net105038) );
  AND2X8 U1247 ( .A(\i_MIPS/ALUin1[0] ), .B(n7475), .Y(n4498) );
  OAI221X4 U1248 ( .A0(net112306), .A1(n8340), .B0(n4419), .B1(net101257), 
        .C0(net112420), .Y(n8344) );
  XOR2X4 U1249 ( .A(n6332), .B(n4629), .Y(n3853) );
  AO21X2 U1250 ( .A0(n10282), .A1(n10281), .B0(net111902), .Y(n10285) );
  AO21X4 U1251 ( .A0(n7806), .A1(n7805), .B0(n7804), .Y(n8751) );
  CLKINVX8 U1252 ( .A(n7154), .Y(n7804) );
  CLKAND2X12 U1253 ( .A(\i_MIPS/Sign_Extend_ID[31] ), .B(n217), .Y(n4380) );
  CLKINVX8 U1254 ( .A(n4062), .Y(n242) );
  INVX20 U1255 ( .A(n242), .Y(mem_addr_I[8]) );
  INVX3 U1256 ( .A(n410), .Y(n4062) );
  CLKINVX8 U1257 ( .A(n4066), .Y(n244) );
  INVX20 U1258 ( .A(n244), .Y(mem_addr_I[11]) );
  INVX3 U1259 ( .A(n411), .Y(n4066) );
  CLKINVX8 U1260 ( .A(n4069), .Y(n246) );
  INVX20 U1261 ( .A(n246), .Y(mem_addr_I[14]) );
  INVX3 U1262 ( .A(n412), .Y(n4069) );
  INVX20 U1263 ( .A(n11170), .Y(n248) );
  INVX20 U1264 ( .A(n248), .Y(n249) );
  INVX20 U1265 ( .A(n248), .Y(n250) );
  INVX20 U1266 ( .A(n248), .Y(n251) );
  INVX20 U1267 ( .A(n248), .Y(n252) );
  INVX16 U1268 ( .A(n248), .Y(n253) );
  BUFX20 U1269 ( .A(n4884), .Y(n4882) );
  NAND3X6 U1270 ( .A(ICACHE_addr[12]), .B(ICACHE_addr[11]), .C(n10242), .Y(
        n10241) );
  INVX8 U1271 ( .A(n10235), .Y(n10242) );
  NAND2X4 U1272 ( .A(net97496), .B(n10439), .Y(n3707) );
  CLKINVX20 U1273 ( .A(net112404), .Y(net97496) );
  NAND2X2 U1274 ( .A(n6559), .B(\i_MIPS/n351 ), .Y(n9242) );
  AOI2BB1X2 U1275 ( .A0N(n7153), .A1N(n7617), .B0(n7804), .Y(n6517) );
  NAND2X6 U1276 ( .A(n4444), .B(n7468), .Y(net102393) );
  INVX8 U1277 ( .A(net107804), .Y(net107794) );
  AND4X4 U1278 ( .A(n6388), .B(n6387), .C(n6386), .D(n6385), .Y(n3906) );
  NAND2X4 U1279 ( .A(n6458), .B(n4499), .Y(net133470) );
  NAND2X4 U1280 ( .A(n4470), .B(n4451), .Y(n8241) );
  OR2X6 U1281 ( .A(n7224), .B(n7521), .Y(n7305) );
  INVXL U1282 ( .A(n9043), .Y(n3776) );
  CLKBUFX8 U1283 ( .A(net112104), .Y(net112096) );
  BUFX12 U1284 ( .A(net112014), .Y(net112006) );
  BUFX6 U1285 ( .A(net100601), .Y(net112046) );
  NAND2X4 U1286 ( .A(n4469), .B(n224), .Y(n4334) );
  BUFX16 U1287 ( .A(n5356), .Y(n5353) );
  CLKINVX4 U1288 ( .A(n4664), .Y(n4331) );
  BUFX8 U1289 ( .A(n8653), .Y(n3844) );
  MXI2X2 U1290 ( .A(n7978), .B(n7977), .S0(net107796), .Y(n4459) );
  INVX3 U1291 ( .A(n10384), .Y(n10238) );
  NAND3X6 U1292 ( .A(n4313), .B(n4314), .C(n9661), .Y(net97874) );
  NOR2X2 U1293 ( .A(n7538), .B(n7536), .Y(n6579) );
  BUFX8 U1294 ( .A(n4934), .Y(n4930) );
  CLKINVX6 U1295 ( .A(n8354), .Y(n9331) );
  CLKINVX1 U1296 ( .A(n8958), .Y(n3849) );
  INVX2 U1297 ( .A(n8352), .Y(n7231) );
  INVX8 U1298 ( .A(net100478), .Y(net111910) );
  INVXL U1299 ( .A(\i_MIPS/forward_unit/n10 ), .Y(n6454) );
  BUFX6 U1300 ( .A(n5153), .Y(n5172) );
  BUFX16 U1301 ( .A(n5223), .Y(n5195) );
  BUFX12 U1302 ( .A(n4839), .Y(n4820) );
  BUFX12 U1303 ( .A(n4839), .Y(n4821) );
  BUFX12 U1304 ( .A(n4839), .Y(n4822) );
  INVX4 U1305 ( .A(net101908), .Y(n3762) );
  AND2X4 U1306 ( .A(n10587), .B(n10585), .Y(n4466) );
  NAND2X4 U1307 ( .A(n10227), .B(n10236), .Y(n10810) );
  NOR4X2 U1308 ( .A(n8447), .B(n8446), .C(n9453), .D(n8445), .Y(n3900) );
  NAND2X2 U1309 ( .A(n9974), .B(n9557), .Y(n11346) );
  INVX4 U1310 ( .A(n11466), .Y(n10654) );
  OA22X2 U1311 ( .A0(n5385), .A1(n3006), .B0(n5347), .B1(n1440), .Y(n10127) );
  OA22X1 U1312 ( .A0(n5213), .A1(n3009), .B0(n5170), .B1(n1441), .Y(n10114) );
  NAND2X4 U1313 ( .A(n10356), .B(n10355), .Y(n4324) );
  AND3X4 U1314 ( .A(n7528), .B(n7527), .C(n7526), .Y(n7529) );
  NAND2X4 U1315 ( .A(net98530), .B(net98531), .Y(n4099) );
  INVX1 U1316 ( .A(n4535), .Y(n3694) );
  NOR2X4 U1317 ( .A(n6544), .B(\i_MIPS/ALUin1[10] ), .Y(n3824) );
  OAI221XL U1318 ( .A0(\i_MIPS/Register/register[18][27] ), .A1(net112078), 
        .B0(\i_MIPS/Register/register[26][27] ), .B1(net112100), .C0(n9374), 
        .Y(n9377) );
  OA22XL U1319 ( .A0(\i_MIPS/Register/register[22][27] ), .A1(net112116), .B0(
        \i_MIPS/Register/register[30][27] ), .B1(net112142), .Y(n9374) );
  NAND2X1 U1320 ( .A(n8852), .B(n8851), .Y(n8871) );
  NAND2X4 U1321 ( .A(n10542), .B(n10540), .Y(n10335) );
  NAND2X4 U1322 ( .A(n3663), .B(n10530), .Y(n9326) );
  INVX3 U1323 ( .A(n10444), .Y(n10333) );
  BUFX12 U1324 ( .A(net112032), .Y(net112026) );
  INVX12 U1325 ( .A(\i_MIPS/ALUin1[6] ), .Y(n7696) );
  NAND2X2 U1326 ( .A(net112376), .B(\i_MIPS/n353 ), .Y(n8153) );
  INVX6 U1327 ( .A(n6590), .Y(n6586) );
  CLKINVX1 U1328 ( .A(n9046), .Y(n255) );
  AND2X2 U1329 ( .A(n437), .B(n2651), .Y(n4392) );
  CLKAND2X6 U1330 ( .A(\i_MIPS/ALUin1[2] ), .B(n4671), .Y(n4517) );
  NAND2X4 U1331 ( .A(n6538), .B(\i_MIPS/ALUin1[1] ), .Y(net103070) );
  NAND2X4 U1332 ( .A(n3772), .B(net98231), .Y(n4098) );
  NAND2X4 U1333 ( .A(n3421), .B(net99161), .Y(n4127) );
  CLKAND2X8 U1334 ( .A(n3321), .B(net98514), .Y(n257) );
  BUFX12 U1335 ( .A(net112014), .Y(net112000) );
  NAND2X4 U1336 ( .A(n6073), .B(n6072), .Y(n6074) );
  NOR2X4 U1337 ( .A(n6106), .B(n6105), .Y(n6107) );
  AND2X4 U1338 ( .A(n7610), .B(n7527), .Y(n4393) );
  INVX3 U1339 ( .A(n3884), .Y(n8650) );
  AND2X2 U1340 ( .A(n4536), .B(n7822), .Y(n4444) );
  NAND2X4 U1341 ( .A(n6558), .B(\i_MIPS/n350 ), .Y(n9138) );
  NAND2X1 U1342 ( .A(\i_MIPS/ALU/N303 ), .B(n6693), .Y(n11178) );
  AND2XL U1343 ( .A(n6693), .B(\i_MIPS/n340 ), .Y(n4455) );
  OA22X1 U1344 ( .A0(\i_MIPS/Register/register[22][1] ), .A1(n4682), .B0(
        \i_MIPS/Register/register[30][1] ), .B1(n4679), .Y(n8036) );
  OAI221XL U1345 ( .A0(\i_MIPS/Register/register[2][1] ), .A1(n4692), .B0(
        \i_MIPS/Register/register[10][1] ), .B1(n4687), .C0(n8027), .Y(n8035)
         );
  OA22XL U1346 ( .A0(\i_MIPS/Register/register[6][1] ), .A1(n4682), .B0(
        \i_MIPS/Register/register[14][1] ), .B1(n4679), .Y(n8027) );
  AO22X1 U1347 ( .A0(net112002), .A1(n641), .B0(net112020), .B1(n2216), .Y(
        n7630) );
  OAI221XL U1348 ( .A0(\i_MIPS/Register/register[18][14] ), .A1(net112072), 
        .B0(\i_MIPS/Register/register[26][14] ), .B1(net112090), .C0(n7638), 
        .Y(n7641) );
  OAI221X1 U1349 ( .A0(\i_MIPS/Register/register[18][28] ), .A1(net112078), 
        .B0(\i_MIPS/Register/register[26][28] ), .B1(net112096), .C0(n8478), 
        .Y(n8481) );
  NAND2X4 U1350 ( .A(n10556), .B(net112404), .Y(n10446) );
  OAI221XL U1351 ( .A0(\i_MIPS/Register/register[2][2] ), .A1(n4692), .B0(
        \i_MIPS/Register/register[10][2] ), .B1(n4688), .C0(n6942), .Y(n6950)
         );
  OAI221XL U1352 ( .A0(\i_MIPS/Register/register[18][20] ), .A1(net112078), 
        .B0(\i_MIPS/Register/register[26][20] ), .B1(net112098), .C0(n9235), 
        .Y(n9238) );
  AO22XL U1353 ( .A0(net112008), .A1(n442), .B0(net112026), .B1(n2025), .Y(
        n8933) );
  NAND3BX1 U1354 ( .AN(n4523), .B(n7698), .C(n6765), .Y(n7976) );
  NOR4X2 U1355 ( .A(n8419), .B(n8418), .C(n8417), .D(n8416), .Y(n8420) );
  OAI221XL U1356 ( .A0(\i_MIPS/Register/register[18][1] ), .A1(net112076), 
        .B0(\i_MIPS/Register/register[26][1] ), .B1(net112090), .C0(n8002), 
        .Y(n8005) );
  OAI221XL U1357 ( .A0(\i_MIPS/Register/register[2][1] ), .A1(net112076), .B0(
        \i_MIPS/Register/register[10][1] ), .B1(net112090), .C0(n7993), .Y(
        n7996) );
  OA22X1 U1358 ( .A0(\i_MIPS/Register/register[6][0] ), .A1(net112112), .B0(
        \i_MIPS/Register/register[14][0] ), .B1(net112142), .Y(n7556) );
  OAI221XL U1359 ( .A0(\i_MIPS/Register/register[18][0] ), .A1(net112072), 
        .B0(\i_MIPS/Register/register[26][0] ), .B1(net112098), .C0(n7565), 
        .Y(n7568) );
  OAI221XL U1360 ( .A0(\i_MIPS/Register/register[2][13] ), .A1(net112076), 
        .B0(\i_MIPS/Register/register[10][13] ), .B1(net112090), .C0(n7722), 
        .Y(n7725) );
  NAND2X2 U1361 ( .A(n8731), .B(n9059), .Y(n7817) );
  CLKINVX6 U1362 ( .A(n6572), .Y(n6554) );
  INVX8 U1363 ( .A(n8737), .Y(n8542) );
  BUFX4 U1364 ( .A(n8649), .Y(n4659) );
  NAND2X6 U1365 ( .A(n6560), .B(\i_MIPS/n349 ), .Y(n9456) );
  INVX6 U1366 ( .A(\i_MIPS/ID_EX[83] ), .Y(n7822) );
  NAND3X6 U1367 ( .A(n4320), .B(n8231), .C(n4321), .Y(n4322) );
  OA22X2 U1368 ( .A0(n4918), .A1(n2106), .B0(n4948), .B1(n512), .Y(n7740) );
  OA22XL U1369 ( .A0(\i_MIPS/Register/register[6][30] ), .A1(n4682), .B0(
        \i_MIPS/Register/register[14][30] ), .B1(n4678), .Y(n6613) );
  OAI221XL U1370 ( .A0(\i_MIPS/Register/register[18][30] ), .A1(n4691), .B0(
        \i_MIPS/Register/register[26][30] ), .B1(n4687), .C0(n6622), .Y(n6630)
         );
  CLKAND2X4 U1371 ( .A(n9043), .B(n8949), .Y(n4423) );
  OA22X2 U1372 ( .A0(\i_MIPS/ALUin1[22] ), .A1(n4670), .B0(\i_MIPS/ALUin1[23] ), .B1(n3828), .Y(n6682) );
  INVX4 U1373 ( .A(n9560), .Y(n10350) );
  OAI221XL U1374 ( .A0(\i_MIPS/Register/register[18][15] ), .A1(net112072), 
        .B0(\i_MIPS/Register/register[26][15] ), .B1(net112098), .C0(n7140), 
        .Y(n7143) );
  OA22XL U1375 ( .A0(\i_MIPS/Register/register[17][15] ), .A1(net112260), .B0(
        \i_MIPS/Register/register[25][15] ), .B1(n148), .Y(n7139) );
  OAI221XL U1376 ( .A0(\i_MIPS/Register/register[2][15] ), .A1(net112072), 
        .B0(\i_MIPS/Register/register[10][15] ), .B1(net112098), .C0(n7131), 
        .Y(n7134) );
  OAI221XL U1377 ( .A0(\i_MIPS/Register/register[18][16] ), .A1(net112076), 
        .B0(\i_MIPS/Register/register[26][16] ), .B1(net112090), .C0(n8060), 
        .Y(n8063) );
  CLKAND2X3 U1378 ( .A(n4672), .B(\i_MIPS/ALUin1[29] ), .Y(n4516) );
  OA22X2 U1379 ( .A0(n5283), .A1(n1286), .B0(n5240), .B1(n2982), .Y(n6124) );
  BUFX12 U1380 ( .A(n4839), .Y(n4819) );
  BUFX16 U1381 ( .A(n4873), .Y(n4865) );
  AND2X4 U1382 ( .A(n4183), .B(n4184), .Y(n6393) );
  INVX3 U1383 ( .A(n6336), .Y(n11011) );
  NOR4X2 U1384 ( .A(n7868), .B(n7867), .C(n7866), .D(n7865), .Y(n7869) );
  OAI221XL U1385 ( .A0(\i_MIPS/Register/register[18][17] ), .A1(n4692), .B0(
        \i_MIPS/Register/register[26][17] ), .B1(n4687), .C0(n7864), .Y(n7872)
         );
  NOR4X2 U1386 ( .A(n8817), .B(n8816), .C(n8815), .D(n8814), .Y(n8818) );
  OR2X4 U1387 ( .A(net112304), .B(n8639), .Y(n4168) );
  INVX3 U1388 ( .A(n9162), .Y(n9166) );
  OAI221XL U1389 ( .A0(\i_MIPS/Register/register[18][4] ), .A1(n4692), .B0(
        \i_MIPS/Register/register[26][4] ), .B1(n4688), .C0(n6907), .Y(n6915)
         );
  NAND4BX2 U1390 ( .AN(n9312), .B(n9311), .C(n9310), .D(n9309), .Y(n9323) );
  NAND3BX2 U1391 ( .AN(n9271), .B(net111994), .C(n9270), .Y(n9286) );
  INVX3 U1392 ( .A(net97703), .Y(net105195) );
  INVXL U1393 ( .A(net111636), .Y(n3891) );
  NOR4X2 U1394 ( .A(n7295), .B(n7294), .C(n7293), .D(n7292), .Y(n7296) );
  AO22XL U1395 ( .A0(n9531), .A1(n327), .B0(n4716), .B1(n479), .Y(n7294) );
  NAND3X6 U1396 ( .A(ICACHE_addr[20]), .B(ICACHE_addr[19]), .C(n10329), .Y(
        net98663) );
  CLKINVX4 U1397 ( .A(n11265), .Y(n9660) );
  MX2X1 U1398 ( .A(n7976), .B(n7813), .S0(net107794), .Y(n7712) );
  AOI2BB1X1 U1399 ( .A0N(net112304), .A1N(n7882), .B0(net100583), .Y(n7883) );
  CLKINVX1 U1400 ( .A(n8443), .Y(n3726) );
  NAND2XL U1401 ( .A(n8539), .B(n3770), .Y(n7820) );
  NAND2XL U1402 ( .A(n9457), .B(n9456), .Y(n9492) );
  AND2X2 U1403 ( .A(net137952), .B(n7225), .Y(n4309) );
  CLKAND2X4 U1404 ( .A(n7893), .B(n8354), .Y(n7236) );
  OA22X1 U1405 ( .A0(n4978), .A1(n2744), .B0(n5023), .B1(n1284), .Y(n9972) );
  OA22X1 U1406 ( .A0(n4918), .A1(n3328), .B0(n4948), .B1(n1726), .Y(n9973) );
  BUFX12 U1407 ( .A(n4486), .Y(n5528) );
  CLKINVX4 U1408 ( .A(n11381), .Y(n10874) );
  INVX6 U1409 ( .A(n11379), .Y(n10687) );
  INVX6 U1410 ( .A(n11378), .Y(n10481) );
  INVX4 U1411 ( .A(n11376), .Y(n10275) );
  INVX4 U1412 ( .A(n11370), .Y(n10660) );
  INVX3 U1413 ( .A(n11369), .Y(n10999) );
  NAND4X2 U1414 ( .A(n7193), .B(n7192), .C(n7191), .D(n7190), .Y(n11365) );
  OA22X2 U1415 ( .A0(n4918), .A1(n2108), .B0(n4948), .B1(n521), .Y(n7748) );
  INVX4 U1416 ( .A(n11356), .Y(n10079) );
  INVX4 U1417 ( .A(n11355), .Y(n10984) );
  NAND4X2 U1418 ( .A(n8994), .B(n8993), .C(n8992), .D(n8991), .Y(n11408) );
  INVX4 U1419 ( .A(n11406), .Y(n10785) );
  INVX1 U1420 ( .A(n11404), .Y(n10218) );
  OA22XL U1421 ( .A0(n4752), .A1(n660), .B0(n4792), .B1(n2248), .Y(n7754) );
  OA22XL U1422 ( .A0(n4830), .A1(n771), .B0(n4875), .B1(n2333), .Y(n7103) );
  OA22XL U1423 ( .A0(n4982), .A1(n775), .B0(n5028), .B1(n2337), .Y(n7101) );
  INVX4 U1424 ( .A(n11389), .Y(n10890) );
  NAND4X2 U1425 ( .A(n6648), .B(n6647), .C(n6646), .D(n6645), .Y(n11445) );
  OA22X2 U1426 ( .A0(n4822), .A1(n2198), .B0(n4868), .B1(n624), .Y(n8194) );
  OA22XL U1427 ( .A0(n4747), .A1(n2162), .B0(n4790), .B1(n586), .Y(n8494) );
  OA22X1 U1428 ( .A0(n4973), .A1(n2142), .B0(n5018), .B1(n562), .Y(n8491) );
  OA22X2 U1429 ( .A0(n4911), .A1(n2091), .B0(n4949), .B1(n504), .Y(n8791) );
  NAND4X2 U1430 ( .A(n7938), .B(n7937), .C(n7936), .D(n7935), .Y(n11421) );
  INVX6 U1431 ( .A(n11472), .Y(n10269) );
  INVX3 U1432 ( .A(n11465), .Y(n10991) );
  OA22X2 U1433 ( .A0(n4977), .A1(n2128), .B0(n5022), .B1(n542), .Y(n7931) );
  NAND4X2 U1434 ( .A(n6802), .B(n6801), .C(n6800), .D(n6799), .Y(n11451) );
  CLKBUFX3 U1435 ( .A(n5525), .Y(n5513) );
  OA22XL U1436 ( .A0(n4977), .A1(n2092), .B0(n5025), .B1(n505), .Y(n7573) );
  OA22XL U1437 ( .A0(n4919), .A1(n1453), .B0(n4949), .B1(n3023), .Y(n7574) );
  CLKBUFX3 U1438 ( .A(n5525), .Y(n5522) );
  OAI221XL U1439 ( .A0(\i_MIPS/Register/register[2][26] ), .A1(n4690), .B0(
        \i_MIPS/Register/register[10][26] ), .B1(n4686), .C0(n8997), .Y(n9005)
         );
  NOR4X1 U1440 ( .A(n9107), .B(n9106), .C(n9105), .D(n9104), .Y(n9108) );
  BUFX8 U1441 ( .A(net137952), .Y(net111996) );
  INVX1 U1442 ( .A(n3848), .Y(n9333) );
  INVX12 U1443 ( .A(net112300), .Y(net112294) );
  BUFX4 U1444 ( .A(\i_MIPS/IR_ID[20] ), .Y(net107810) );
  NOR4X2 U1445 ( .A(n8671), .B(n8670), .C(n8669), .D(n8668), .Y(n8682) );
  OA22X2 U1446 ( .A0(\i_MIPS/ALUin1[9] ), .A1(n4670), .B0(\i_MIPS/ALUin1[8] ), 
        .B1(n3828), .Y(n6839) );
  MX2X1 U1447 ( .A(net101082), .B(net112415), .S0(n3685), .Y(n6854) );
  OA22X2 U1448 ( .A0(n5119), .A1(n2992), .B0(n5056), .B1(n1434), .Y(n9901) );
  NAND4X2 U1449 ( .A(n10101), .B(n10100), .C(n10099), .D(n10098), .Y(n11192)
         );
  NAND4X2 U1450 ( .A(n10030), .B(n10029), .C(n10028), .D(n10027), .Y(n11195)
         );
  OA22X2 U1451 ( .A0(n5400), .A1(n3001), .B0(n5332), .B1(n1438), .Y(n6152) );
  OA22X2 U1452 ( .A0(n5377), .A1(n2986), .B0(n5348), .B1(n1430), .Y(n10196) );
  OA22X2 U1453 ( .A0(n5119), .A1(n2991), .B0(n5089), .B1(n1433), .Y(n9905) );
  NAND4X2 U1454 ( .A(n10106), .B(n10105), .C(n10104), .D(n10103), .Y(n11224)
         );
  NAND4X2 U1455 ( .A(n10011), .B(n10010), .C(n10009), .D(n10008), .Y(n11226)
         );
  NAND4X2 U1456 ( .A(n9937), .B(n9936), .C(n9935), .D(n9934), .Y(n11252) );
  NAND4X2 U1457 ( .A(n9897), .B(n9896), .C(n9895), .D(n9894), .Y(n11254) );
  OA22X2 U1458 ( .A0(n5119), .A1(n2990), .B0(n5073), .B1(n1432), .Y(n9897) );
  NAND4X2 U1459 ( .A(n9918), .B(n9917), .C(n9916), .D(n9915), .Y(n11255) );
  OA22X2 U1460 ( .A0(n5381), .A1(n3002), .B0(n5332), .B1(n1439), .Y(n6137) );
  OA22X2 U1461 ( .A0(n5300), .A1(n2994), .B0(n5240), .B1(n1436), .Y(n6133) );
  NAND4X2 U1462 ( .A(n10182), .B(n10181), .C(n10180), .D(n10179), .Y(n11285)
         );
  OA22X2 U1463 ( .A0(n5290), .A1(n2995), .B0(n5240), .B1(n1437), .Y(n6128) );
  NAND4X2 U1464 ( .A(n10091), .B(n10090), .C(n10089), .D(n10088), .Y(n11288)
         );
  NAND4X2 U1465 ( .A(n9996), .B(n9995), .C(n9994), .D(n9993), .Y(n11290) );
  NAND4X2 U1466 ( .A(n10020), .B(n10019), .C(n10018), .D(n10017), .Y(n11291)
         );
  NAND4X4 U1467 ( .A(n9642), .B(n9641), .C(n9640), .D(n9639), .Y(n11297) );
  OA22XL U1468 ( .A0(n4822), .A1(n684), .B0(n4868), .B1(n2256), .Y(n8102) );
  OA22X1 U1469 ( .A0(n4830), .A1(n668), .B0(n4875), .B1(n2239), .Y(n7018) );
  NAND4X4 U1470 ( .A(n7197), .B(n7196), .C(n7195), .D(n7194), .Y(n11397) );
  OA22XL U1471 ( .A0(n4829), .A1(n2074), .B0(n4874), .B1(n484), .Y(n7196) );
  OA22X2 U1472 ( .A0(n4824), .A1(n2073), .B0(n4869), .B1(n483), .Y(n7851) );
  OA22XL U1473 ( .A0(n4831), .A1(n815), .B0(n4876), .B1(n2378), .Y(n7010) );
  OA22XL U1474 ( .A0(n4818), .A1(n2143), .B0(n263), .B1(n563), .Y(n8690) );
  OA22X2 U1475 ( .A0(n4971), .A1(n2153), .B0(n5016), .B1(n574), .Y(n8688) );
  OA22XL U1476 ( .A0(n4829), .A1(n2196), .B0(n4874), .B1(n622), .Y(n7270) );
  OA22XL U1477 ( .A0(n4756), .A1(n2195), .B0(n4793), .B1(n621), .Y(n7271) );
  NAND4X4 U1478 ( .A(n7189), .B(n7188), .C(n7187), .D(n7186), .Y(n11429) );
  OA22X1 U1479 ( .A0(n4829), .A1(n2149), .B0(n4874), .B1(n569), .Y(n7188) );
  OA22X2 U1480 ( .A0(n4981), .A1(n2147), .B0(n5027), .B1(n567), .Y(n7186) );
  OA22XL U1481 ( .A0(n4822), .A1(n691), .B0(n4868), .B1(n2260), .Y(n8098) );
  OA22X2 U1482 ( .A0(n4975), .A1(n2087), .B0(n5020), .B1(n499), .Y(n8096) );
  OA22X1 U1483 ( .A0(n4909), .A1(n3399), .B0(n4947), .B1(n1770), .Y(n9293) );
  OA22X2 U1484 ( .A0(n4911), .A1(n3356), .B0(n4949), .B1(n1736), .Y(n8886) );
  NAND4X2 U1485 ( .A(n8304), .B(n8303), .C(n8302), .D(n8301), .Y(n11438) );
  INVXL U1486 ( .A(n11446), .Y(n10953) );
  OA22XL U1487 ( .A0(n4751), .A1(n834), .B0(n4791), .B1(n2397), .Y(n8012) );
  OA22XL U1488 ( .A0(n4830), .A1(n699), .B0(n4875), .B1(n2268), .Y(n7091) );
  OA22X1 U1489 ( .A0(n4982), .A1(n718), .B0(n5028), .B1(n2286), .Y(n7089) );
  NAND4X2 U1490 ( .A(n9291), .B(n9290), .C(n9289), .D(n9288), .Y(n11466) );
  NAND4X2 U1491 ( .A(n8884), .B(n8883), .C(n8882), .D(n8881), .Y(n11469) );
  NAND4X2 U1492 ( .A(n8490), .B(n8489), .C(n8488), .D(n8487), .Y(n11474) );
  OA22X1 U1493 ( .A0(n4748), .A1(n2205), .B0(n4790), .B1(n500), .Y(n8490) );
  OA22X2 U1494 ( .A0(n4913), .A1(n2077), .B0(n4249), .B1(n489), .Y(n8488) );
  NAND4X2 U1495 ( .A(n6302), .B(n6301), .C(n6300), .D(n6299), .Y(n11476) );
  NAND4X4 U1496 ( .A(n4328), .B(n6362), .C(n6361), .D(n6360), .Y(n11490) );
  NAND4X4 U1497 ( .A(n6422), .B(n6421), .C(n6420), .D(n6419), .Y(n11500) );
  NAND4X4 U1498 ( .A(n6380), .B(n6379), .C(n6378), .D(n6377), .Y(n11501) );
  NAND4X2 U1499 ( .A(n6431), .B(n6430), .C(n6429), .D(n6428), .Y(n11502) );
  OA22X2 U1500 ( .A0(n4834), .A1(n2998), .B0(n4879), .B1(n556), .Y(n6430) );
  AOI2BB1X2 U1501 ( .A0N(n8362), .A1N(net137891), .B0(n8361), .Y(n8363) );
  CLKINVX4 U1502 ( .A(n11092), .Y(n11098) );
  XOR2X1 U1503 ( .A(n10225), .B(ICACHE_addr[18]), .Y(n10531) );
  XOR2X2 U1504 ( .A(net98663), .B(ICACHE_addr[21]), .Y(net98497) );
  CLKINVX1 U1505 ( .A(n11162), .Y(n11161) );
  XOR3X2 U1506 ( .A(net112400), .B(n10836), .C(n10835), .Y(n10841) );
  INVX12 U1507 ( .A(net108662), .Y(net108660) );
  NAND4X4 U1508 ( .A(n10063), .B(n10062), .C(n10061), .D(n10060), .Y(n10394)
         );
  CLKINVX1 U1509 ( .A(n11047), .Y(n11060) );
  AND2X6 U1510 ( .A(n11064), .B(n270), .Y(n4461) );
  NOR2X4 U1511 ( .A(n6545), .B(\i_MIPS/ALUin1[11] ), .Y(n3771) );
  AND2X4 U1512 ( .A(n3785), .B(n3783), .Y(n4527) );
  AND2X2 U1513 ( .A(\i_MIPS/IR_ID[21] ), .B(\i_MIPS/n232 ), .Y(n402) );
  NAND2X2 U1514 ( .A(n3324), .B(n10926), .Y(n8430) );
  NAND2X1 U1515 ( .A(n10446), .B(n10449), .Y(n10334) );
  CLKMX2X4 U1516 ( .A(\i_MIPS/n269 ), .B(n4497), .S0(n5622), .Y(n6570) );
  NAND2X4 U1517 ( .A(n7492), .B(n7500), .Y(n7163) );
  NAND2X2 U1518 ( .A(n4381), .B(n7511), .Y(n7051) );
  NAND2X6 U1519 ( .A(n4228), .B(n4229), .Y(n6403) );
  INVX4 U1520 ( .A(n3816), .Y(n4228) );
  NAND2X2 U1521 ( .A(n1776), .B(n11484), .Y(n4158) );
  OR2X4 U1522 ( .A(n1776), .B(n11484), .Y(n4157) );
  NAND2X2 U1523 ( .A(n3901), .B(n11485), .Y(n4186) );
  XNOR2X1 U1524 ( .A(n11500), .B(n3763), .Y(n6423) );
  XOR2X1 U1525 ( .A(n4628), .B(n11492), .Y(n4641) );
  XOR2X1 U1526 ( .A(n11490), .B(n3409), .Y(n4640) );
  XNOR2X1 U1527 ( .A(DCACHE_addr[9]), .B(n11487), .Y(n4639) );
  OA21XL U1528 ( .A0(n7493), .A1(n7492), .B0(n7527), .Y(n7501) );
  NAND2BX1 U1529 ( .AN(n7515), .B(n8635), .Y(n7522) );
  CLKAND2X8 U1530 ( .A(\i_MIPS/IR_ID[23] ), .B(\i_MIPS/n234 ), .Y(n4503) );
  AND2X4 U1531 ( .A(\i_MIPS/n234 ), .B(\i_MIPS/n233 ), .Y(n4446) );
  CLKAND2X8 U1532 ( .A(\i_MIPS/IR_ID[24] ), .B(\i_MIPS/n233 ), .Y(n4504) );
  CLKAND2X3 U1533 ( .A(\i_MIPS/n231 ), .B(\i_MIPS/n232 ), .Y(n4447) );
  INVX3 U1534 ( .A(n3812), .Y(n3813) );
  CLKINVX3 U1535 ( .A(\i_MIPS/ALU_Control/n10 ), .Y(n4077) );
  NAND2X6 U1536 ( .A(n4420), .B(n7050), .Y(n7160) );
  NAND2X4 U1537 ( .A(n8630), .B(n7496), .Y(n7167) );
  NAND3BX2 U1538 ( .AN(n4661), .B(n3785), .C(n3784), .Y(n10195) );
  NAND2X1 U1539 ( .A(n9328), .B(net107794), .Y(n9255) );
  NAND2X2 U1540 ( .A(\i_MIPS/IR_ID[17] ), .B(\i_MIPS/n312 ), .Y(n6611) );
  AND2X2 U1541 ( .A(net112374), .B(\i_MIPS/n358 ), .Y(n4473) );
  NAND2X1 U1542 ( .A(\i_MIPS/ALUin1[18] ), .B(net112338), .Y(n6920) );
  OA22X1 U1543 ( .A0(\i_MIPS/Register/register[22][28] ), .A1(net112116), .B0(
        \i_MIPS/Register/register[30][28] ), .B1(net112134), .Y(n8478) );
  NAND2X2 U1544 ( .A(n4389), .B(n10399), .Y(n10418) );
  NAND2X4 U1545 ( .A(net98499), .B(net98500), .Y(n8918) );
  NAND2X2 U1546 ( .A(n3422), .B(n10584), .Y(n8725) );
  NAND2X2 U1547 ( .A(n3417), .B(n10548), .Y(n9549) );
  OA22X1 U1548 ( .A0(\i_MIPS/Register/register[22][0] ), .A1(net112112), .B0(
        \i_MIPS/Register/register[30][0] ), .B1(net112142), .Y(n7565) );
  INVX6 U1549 ( .A(n4616), .Y(n6531) );
  NAND2X1 U1550 ( .A(n8433), .B(n11181), .Y(n8454) );
  NAND2X2 U1551 ( .A(n6593), .B(n7149), .Y(n8444) );
  CLKINVX1 U1552 ( .A(n8454), .Y(n8436) );
  NAND2X1 U1553 ( .A(net112294), .B(n8451), .Y(n8435) );
  NAND3BX1 U1554 ( .AN(n4526), .B(n6920), .C(n6491), .Y(n8740) );
  OA22X2 U1555 ( .A0(net112368), .A1(\i_MIPS/n356 ), .B0(net112350), .B1(
        \i_MIPS/n355 ), .Y(n6491) );
  NAND2X1 U1556 ( .A(net112356), .B(\i_MIPS/n357 ), .Y(n8068) );
  OAI2BB1X2 U1557 ( .A0N(\i_MIPS/n364 ), .A1N(\i_MIPS/n363 ), .B0(n6505), .Y(
        n6508) );
  INVX3 U1558 ( .A(n7400), .Y(n7402) );
  NAND2X2 U1559 ( .A(n6547), .B(\i_MIPS/n358 ), .Y(n7708) );
  INVX6 U1560 ( .A(n6573), .Y(n6553) );
  AND2X4 U1561 ( .A(n8753), .B(n8752), .Y(n4468) );
  NAND2X4 U1562 ( .A(n8751), .B(n8749), .Y(n8535) );
  NOR2X6 U1563 ( .A(n6572), .B(\i_MIPS/ALUin1[19] ), .Y(n3662) );
  NAND2X1 U1564 ( .A(n4393), .B(n8072), .Y(n8538) );
  AND2X4 U1565 ( .A(\i_MIPS/ALUin1[17] ), .B(n4671), .Y(n4526) );
  CLKMX2X4 U1566 ( .A(\i_MIPS/n293 ), .B(n3837), .S0(n5624), .Y(n7053) );
  INVX3 U1567 ( .A(n7053), .Y(n7495) );
  CLKAND2X6 U1568 ( .A(\i_MIPS/ALUin1[14] ), .B(n4671), .Y(n4523) );
  NAND2X4 U1569 ( .A(n4378), .B(n4163), .Y(n4164) );
  NAND2X4 U1570 ( .A(n8738), .B(n8546), .Y(n9139) );
  NAND2X4 U1571 ( .A(\i_MIPS/ALUin1[20] ), .B(n6559), .Y(n9262) );
  INVX4 U1572 ( .A(n6548), .Y(n6560) );
  CLKINVX4 U1573 ( .A(n8944), .Y(n4321) );
  CLKINVX1 U1574 ( .A(n9268), .Y(n7538) );
  CLKINVX1 U1575 ( .A(n9482), .Y(n3826) );
  NAND2X6 U1576 ( .A(\i_MIPS/ALUin1[11] ), .B(n6545), .Y(n7409) );
  OR2X1 U1577 ( .A(net112348), .B(\i_MIPS/n350 ), .Y(n4167) );
  AND2X2 U1578 ( .A(mem_ready_D), .B(n11478), .Y(n4524) );
  BUFX12 U1579 ( .A(n9988), .Y(n4891) );
  OAI221X1 U1580 ( .A0(\i_MIPS/ALUin1[19] ), .A1(net112364), .B0(
        \i_MIPS/ALUin1[20] ), .B1(net112346), .C0(n6490), .Y(n8956) );
  OA22X2 U1581 ( .A0(\i_MIPS/ALUin1[21] ), .A1(n4670), .B0(\i_MIPS/ALUin1[22] ), .B1(n3828), .Y(n6490) );
  CLKINVX1 U1582 ( .A(n8950), .Y(n8967) );
  AO22X1 U1583 ( .A0(n4723), .A1(n643), .B0(n4719), .B1(n2218), .Y(n8516) );
  INVX3 U1584 ( .A(n6592), .Y(n6588) );
  XNOR2X1 U1585 ( .A(n12952), .B(n11483), .Y(n6368) );
  AND4X4 U1586 ( .A(n4639), .B(n4638), .C(n4641), .D(n4640), .Y(n6366) );
  AND2X4 U1587 ( .A(\i_MIPS/IR_ID[18] ), .B(\i_MIPS/n318 ), .Y(n4500) );
  NAND2X4 U1588 ( .A(n4522), .B(n4445), .Y(n9415) );
  AND2X4 U1589 ( .A(\i_MIPS/IR_ID[19] ), .B(\i_MIPS/n316 ), .Y(n4502) );
  NAND2BX2 U1590 ( .AN(n4989), .B(\D_cache/cache[6][154] ), .Y(n6304) );
  NAND2BX2 U1591 ( .AN(n4927), .B(\D_cache/cache[4][154] ), .Y(n6306) );
  NAND2BX2 U1592 ( .AN(n4837), .B(\D_cache/cache[2][154] ), .Y(n6308) );
  NAND2BX2 U1593 ( .AN(n4765), .B(\D_cache/cache[0][154] ), .Y(n6310) );
  NAND2BX2 U1594 ( .AN(n4796), .B(\D_cache/cache[1][154] ), .Y(n6309) );
  BUFX12 U1595 ( .A(n10195), .Y(n5313) );
  NAND3BX2 U1596 ( .AN(n7482), .B(n4454), .C(n8433), .Y(net103914) );
  INVX3 U1597 ( .A(net133411), .Y(net103907) );
  INVX3 U1598 ( .A(n8948), .Y(n7490) );
  OR2X6 U1599 ( .A(n7821), .B(n4171), .Y(n7968) );
  OA22X1 U1600 ( .A0(\i_MIPS/Register/register[17][12] ), .A1(net112258), .B0(
        \i_MIPS/Register/register[25][12] ), .B1(n147), .Y(n7392) );
  OAI221X1 U1601 ( .A0(\i_MIPS/Register/register[18][19] ), .A1(net112078), 
        .B0(\i_MIPS/Register/register[26][19] ), .B1(net112096), .C0(n8576), 
        .Y(n8584) );
  AND4X1 U1602 ( .A(n415), .B(n303), .C(\i_MIPS/forward_unit/n25 ), .D(n4534), 
        .Y(\i_MIPS/forward_unit/n10 ) );
  XNOR2X1 U1603 ( .A(ICACHE_addr[23]), .B(n11338), .Y(n5997) );
  CLKMX2X2 U1604 ( .A(\i_MIPS/ID_EX[75] ), .B(net127930), .S0(n3812), .Y(
        net127703) );
  INVX6 U1605 ( .A(net103923), .Y(net103913) );
  INVX3 U1606 ( .A(n6755), .Y(n6757) );
  NAND2X1 U1607 ( .A(n7798), .B(n7797), .Y(n8070) );
  BUFX4 U1608 ( .A(n5090), .Y(n5134) );
  BUFX2 U1609 ( .A(n4999), .Y(n5040) );
  NAND2X6 U1610 ( .A(\i_MIPS/ALUin1[3] ), .B(n6539), .Y(n8341) );
  AO22X2 U1611 ( .A0(n4722), .A1(n292), .B0(n4719), .B1(n2062), .Y(n7445) );
  OAI221XL U1612 ( .A0(\i_MIPS/Register/register[2][12] ), .A1(n4692), .B0(
        \i_MIPS/Register/register[10][12] ), .B1(n4687), .C0(n7443), .Y(n7451)
         );
  NOR4X1 U1613 ( .A(n7456), .B(n7455), .C(n7454), .D(n7453), .Y(n7457) );
  AO22X2 U1614 ( .A0(n4723), .A1(n291), .B0(n4719), .B1(n2061), .Y(n7454) );
  AO22X1 U1615 ( .A0(n4720), .A1(n468), .B0(n4719), .B1(n2055), .Y(n9315) );
  AO22X1 U1616 ( .A0(n4713), .A1(n305), .B0(n4710), .B1(n2022), .Y(n9317) );
  AO22X1 U1617 ( .A0(n4723), .A1(n469), .B0(n4719), .B1(n2056), .Y(n9306) );
  NAND2X1 U1618 ( .A(n9243), .B(n9242), .Y(n9281) );
  CLKINVX1 U1619 ( .A(n4251), .Y(n9270) );
  NOR4X1 U1620 ( .A(n8328), .B(n8327), .C(n8326), .D(n8325), .Y(n8329) );
  AO22X1 U1621 ( .A0(n4723), .A1(n639), .B0(n4719), .B1(n2214), .Y(n8326) );
  OA22X1 U1622 ( .A0(\i_MIPS/Register/register[22][24] ), .A1(n4682), .B0(
        \i_MIPS/Register/register[30][24] ), .B1(n4679), .Y(n8324) );
  OA22X1 U1623 ( .A0(\i_MIPS/Register/register[6][24] ), .A1(n4682), .B0(
        \i_MIPS/Register/register[14][24] ), .B1(n4679), .Y(n8315) );
  CLKINVX1 U1624 ( .A(n8261), .Y(n8262) );
  CLKINVX1 U1625 ( .A(n7875), .Y(n6971) );
  OAI221X1 U1626 ( .A0(\i_MIPS/ALUin1[11] ), .A1(n4668), .B0(
        \i_MIPS/ALUin1[10] ), .B1(n3828), .C0(n6922), .Y(net104885) );
  AOI2BB1X1 U1627 ( .A0N(\i_MIPS/ALUin1[12] ), .A1N(net112350), .B0(n4473), 
        .Y(n6922) );
  AO22X1 U1628 ( .A0(net112000), .A1(n465), .B0(net112018), .B1(n2052), .Y(
        n6873) );
  AO22X1 U1629 ( .A0(net112000), .A1(n464), .B0(net112018), .B1(n2051), .Y(
        n6864) );
  CLKMX2X2 U1630 ( .A(n9380), .B(n9379), .S0(net107816), .Y(n9381) );
  AO22X1 U1631 ( .A0(net112008), .A1(n275), .B0(net112026), .B1(n307), .Y(
        n9375) );
  OAI221XL U1632 ( .A0(\i_MIPS/Register/register[18][17] ), .A1(net112076), 
        .B0(\i_MIPS/Register/register[26][17] ), .B1(net112090), .C0(n7790), 
        .Y(n7793) );
  OAI221XL U1633 ( .A0(\i_MIPS/Register/register[2][17] ), .A1(net112076), 
        .B0(\i_MIPS/Register/register[10][17] ), .B1(net112090), .C0(n7781), 
        .Y(n7784) );
  AO22X1 U1634 ( .A0(net112004), .A1(n328), .B0(net112030), .B1(n651), .Y(
        n7782) );
  NAND2X1 U1635 ( .A(n8857), .B(n8850), .Y(net101554) );
  AO22X1 U1636 ( .A0(net112008), .A1(n461), .B0(net112026), .B1(n2048), .Y(
        n9131) );
  AO22X1 U1637 ( .A0(net112008), .A1(n460), .B0(net112026), .B1(n2047), .Y(
        n9122) );
  CLKINVX1 U1638 ( .A(n10226), .Y(n10283) );
  CLKINVX1 U1639 ( .A(n11297), .Y(n9663) );
  CLKINVX1 U1640 ( .A(n11201), .Y(n9662) );
  OR2X1 U1641 ( .A(n10556), .B(net112404), .Y(n3681) );
  NAND2X2 U1642 ( .A(n10613), .B(n10611), .Y(n10435) );
  CLKINVX1 U1643 ( .A(n10575), .Y(n10571) );
  AND2X2 U1644 ( .A(n3432), .B(net97452), .Y(n1774) );
  NAND2X1 U1645 ( .A(n10448), .B(net112404), .Y(n10463) );
  OAI221XL U1646 ( .A0(\i_MIPS/Register/register[18][10] ), .A1(net112072), 
        .B0(\i_MIPS/Register/register[26][10] ), .B1(net112098), .C0(n7336), 
        .Y(n7339) );
  OA22X1 U1647 ( .A0(\i_MIPS/Register/register[17][10] ), .A1(net112260), .B0(
        \i_MIPS/Register/register[25][10] ), .B1(n147), .Y(n7335) );
  OAI221XL U1648 ( .A0(\i_MIPS/Register/register[2][10] ), .A1(net112072), 
        .B0(\i_MIPS/Register/register[10][10] ), .B1(net112098), .C0(n7327), 
        .Y(n7330) );
  NAND4X1 U1649 ( .A(n7326), .B(n7325), .C(n7324), .D(n7323), .Y(n7331) );
  OA22X1 U1650 ( .A0(\i_MIPS/Register/register[1][10] ), .A1(net112254), .B0(
        \i_MIPS/Register/register[9][10] ), .B1(n151), .Y(n7326) );
  OA22X1 U1651 ( .A0(\i_MIPS/Register/register[22][3] ), .A1(n4682), .B0(
        \i_MIPS/Register/register[30][3] ), .B1(n4679), .Y(n8415) );
  OA22X1 U1652 ( .A0(\i_MIPS/Register/register[6][3] ), .A1(n4682), .B0(
        \i_MIPS/Register/register[14][3] ), .B1(n4679), .Y(n8406) );
  AO22X1 U1653 ( .A0(n4722), .A1(n458), .B0(n4719), .B1(n2044), .Y(n8121) );
  OA22X1 U1654 ( .A0(\i_MIPS/Register/register[22][16] ), .A1(n4682), .B0(
        \i_MIPS/Register/register[30][16] ), .B1(n4679), .Y(n8119) );
  AO22X1 U1655 ( .A0(n4722), .A1(n459), .B0(n4719), .B1(n2045), .Y(n8112) );
  OA22X1 U1656 ( .A0(\i_MIPS/Register/register[6][16] ), .A1(n4682), .B0(
        \i_MIPS/Register/register[14][16] ), .B1(n4679), .Y(n8110) );
  NAND2X2 U1657 ( .A(n11090), .B(n11089), .Y(n10361) );
  OA22X1 U1658 ( .A0(\i_MIPS/ALUin1[8] ), .A1(n4670), .B0(\i_MIPS/ALUin1[7] ), 
        .B1(n3828), .Y(n7897) );
  AO22X2 U1659 ( .A0(net100583), .A1(n8454), .B0(n8453), .B1(net100585), .Y(
        n8459) );
  AOI211X1 U1660 ( .A0(n8441), .A1(net102253), .B0(n4512), .C0(n4510), .Y(
        n8442) );
  CLKMX2X2 U1661 ( .A(net101082), .B(net112415), .S0(n8444), .Y(n8445) );
  OAI2BB2X1 U1662 ( .B0(n8435), .B1(n9347), .A0N(n9338), .A1N(n8448), .Y(n8447) );
  OAI221XL U1663 ( .A0(\i_MIPS/Register/register[18][18] ), .A1(net112078), 
        .B0(\i_MIPS/Register/register[26][18] ), .B1(net112098), .C0(n8778), 
        .Y(n8781) );
  CLKAND2X3 U1664 ( .A(\i_MIPS/ALUin1[5] ), .B(net112372), .Y(net127833) );
  CLKMX2X2 U1665 ( .A(n8740), .B(n8739), .S0(net107794), .Y(n8966) );
  CLKINVX1 U1666 ( .A(n8738), .Y(n9275) );
  INVX3 U1667 ( .A(n9154), .Y(n8167) );
  CLKINVX1 U1668 ( .A(n7967), .Y(n7827) );
  NAND2X4 U1669 ( .A(n8750), .B(n8730), .Y(n9140) );
  INVX3 U1670 ( .A(n8355), .Y(n8351) );
  NAND2X2 U1671 ( .A(\i_MIPS/ALUin1[18] ), .B(n6574), .Y(n8736) );
  AO22X1 U1672 ( .A0(net112008), .A1(n463), .B0(net112026), .B1(n2050), .Y(
        n9034) );
  AO22X1 U1673 ( .A0(net112008), .A1(n462), .B0(net112026), .B1(n2049), .Y(
        n9025) );
  NAND2X4 U1674 ( .A(n7060), .B(n4536), .Y(n8264) );
  OAI222X1 U1675 ( .A0(n9167), .A1(n9469), .B0(n9463), .B1(n8159), .C0(n8158), 
        .C1(net133688), .Y(n8161) );
  CLKINVX1 U1676 ( .A(n8172), .Y(n8174) );
  NAND2X1 U1677 ( .A(n11183), .B(n8150), .Y(n8175) );
  NAND2X1 U1678 ( .A(n7805), .B(n7154), .Y(n7171) );
  CLKAND2X3 U1679 ( .A(n9145), .B(n7610), .Y(n4172) );
  INVX3 U1680 ( .A(n7805), .Y(n7153) );
  AOI2BB1X2 U1681 ( .A0N(net112332), .A1N(\i_MIPS/n368 ), .B0(n4517), .Y(n6685) );
  INVX3 U1682 ( .A(n7227), .Y(n8348) );
  AOI2BB1X1 U1683 ( .A0N(\i_MIPS/ALUin1[15] ), .A1N(n3828), .B0(n4463), .Y(
        n7151) );
  AND2X2 U1684 ( .A(n4659), .B(\i_MIPS/n340 ), .Y(n4449) );
  INVX4 U1685 ( .A(n4659), .Y(n8349) );
  OAI211X1 U1686 ( .A0(\i_MIPS/ALUin1[16] ), .A1(net112350), .B0(n8251), .C0(
        n6923), .Y(net104868) );
  AOI2BB1X2 U1687 ( .A0N(net112368), .A1N(\i_MIPS/n368 ), .B0(net127829), .Y(
        n6484) );
  NAND2X4 U1688 ( .A(\i_MIPS/ALUin1[14] ), .B(n6576), .Y(n7609) );
  OAI221X1 U1689 ( .A0(net112304), .A1(n4320), .B0(n9481), .B1(net101257), 
        .C0(net112420), .Y(n7613) );
  OAI221X1 U1690 ( .A0(\i_MIPS/ALUin1[22] ), .A1(net112364), .B0(
        \i_MIPS/ALUin1[23] ), .B1(net112346), .C0(n8164), .Y(n9047) );
  NAND2X1 U1691 ( .A(n8852), .B(n8236), .Y(n6580) );
  CLKMX2X4 U1692 ( .A(n8352), .B(n4519), .S0(net107794), .Y(n8354) );
  AO21X1 U1693 ( .A0(n10078), .A1(n10077), .B0(n10076), .Y(n10084) );
  OA22X1 U1694 ( .A0(n4923), .A1(n767), .B0(n4949), .B1(n2329), .Y(n7349) );
  OA22X2 U1695 ( .A0(n4922), .A1(n3395), .B0(n4249), .B1(n1766), .Y(n7094) );
  INVX8 U1696 ( .A(n4950), .Y(n4248) );
  OA22X2 U1697 ( .A0(n4918), .A1(n2141), .B0(n4949), .B1(n561), .Y(n7345) );
  BUFX4 U1698 ( .A(n4800), .Y(n4799) );
  OAI222X1 U1699 ( .A0(net133471), .A1(n8970), .B0(n8969), .B1(n8968), .C0(
        n8967), .C1(net112420), .Y(n8971) );
  AO22X2 U1700 ( .A0(n9328), .A1(n8966), .B0(n8965), .B1(n9327), .Y(n8972) );
  INVX1 U1701 ( .A(n8964), .Y(n8965) );
  OA22X1 U1702 ( .A0(\i_MIPS/Register/register[6][28] ), .A1(n4682), .B0(
        \i_MIPS/Register/register[14][28] ), .B1(n4679), .Y(n8505) );
  INVX4 U1703 ( .A(n4675), .Y(n3761) );
  NOR4X1 U1704 ( .A(n8218), .B(n8217), .C(n8216), .D(n8215), .Y(n8219) );
  AO22X1 U1705 ( .A0(n4722), .A1(n475), .B0(n4719), .B1(n2067), .Y(n8216) );
  NOR4X1 U1706 ( .A(n8209), .B(n8208), .C(n8207), .D(n8206), .Y(n8210) );
  AO22X1 U1707 ( .A0(n4722), .A1(n476), .B0(n4719), .B1(n2068), .Y(n8207) );
  INVX3 U1708 ( .A(n8941), .Y(n6519) );
  NAND2X4 U1709 ( .A(n4522), .B(n4500), .Y(n9417) );
  NAND2X6 U1710 ( .A(n4505), .B(n4445), .Y(n9411) );
  CLKXOR2X2 U1711 ( .A(n259), .B(net107812), .Y(n6609) );
  AO22X1 U1712 ( .A0(n9531), .A1(n455), .B0(n4715), .B1(n2041), .Y(n9210) );
  NOR4X1 U1713 ( .A(n7761), .B(n7760), .C(n7759), .D(n7758), .Y(n7762) );
  AO22X1 U1714 ( .A0(n4722), .A1(n440), .B0(n4719), .B1(n2023), .Y(n7759) );
  NOR4X1 U1715 ( .A(n7770), .B(n7769), .C(n7768), .D(n7767), .Y(n7771) );
  AO22X1 U1716 ( .A0(n4722), .A1(n439), .B0(n4719), .B1(n2020), .Y(n7768) );
  OR2X2 U1717 ( .A(n7542), .B(n7541), .Y(n3856) );
  OA21XL U1718 ( .A0(net103917), .A1(net102253), .B0(net103919), .Y(n7489) );
  NAND2X1 U1719 ( .A(n10065), .B(n3783), .Y(n10178) );
  OAI221XL U1720 ( .A0(\i_MIPS/Register/register[2][3] ), .A1(net112078), .B0(
        \i_MIPS/Register/register[10][3] ), .B1(net112096), .C0(n8371), .Y(
        n8374) );
  AO22X1 U1721 ( .A0(net112000), .A1(n466), .B0(net112018), .B1(n2053), .Y(
        n6792) );
  AO22X1 U1722 ( .A0(net112000), .A1(n445), .B0(net112018), .B1(n2028), .Y(
        n6783) );
  AO22X1 U1723 ( .A0(net112000), .A1(n446), .B0(net112018), .B1(n2029), .Y(
        n6998) );
  AO22X1 U1724 ( .A0(net112000), .A1(n444), .B0(net112018), .B1(n2027), .Y(
        n6989) );
  NOR4X1 U1725 ( .A(n7927), .B(n7926), .C(n7925), .D(n7924), .Y(n7928) );
  NAND4X1 U1726 ( .A(n7922), .B(n7921), .C(n7920), .D(n7919), .Y(n7927) );
  OAI221XL U1727 ( .A0(\i_MIPS/Register/register[18][8] ), .A1(net112072), 
        .B0(\i_MIPS/Register/register[26][8] ), .B1(net112098), .C0(n7081), 
        .Y(n7084) );
  AO22X1 U1728 ( .A0(net112000), .A1(n467), .B0(net112018), .B1(n2054), .Y(
        n7082) );
  OAI221XL U1729 ( .A0(\i_MIPS/Register/register[2][8] ), .A1(net112072), .B0(
        \i_MIPS/Register/register[10][8] ), .B1(net112098), .C0(n7072), .Y(
        n7075) );
  NAND4X1 U1730 ( .A(n8666), .B(n8665), .C(n8664), .D(n8663), .Y(n8671) );
  OAI221XL U1731 ( .A0(\i_MIPS/Register/register[2][9] ), .A1(net112078), .B0(
        \i_MIPS/Register/register[10][9] ), .B1(net112096), .C0(n8667), .Y(
        n8670) );
  OA22X1 U1732 ( .A0(\i_MIPS/Register/register[1][12] ), .A1(net112258), .B0(
        \i_MIPS/Register/register[9][12] ), .B1(n150), .Y(n7383) );
  OAI221X1 U1733 ( .A0(\i_MIPS/Register/register[2][12] ), .A1(net112072), 
        .B0(\i_MIPS/Register/register[10][12] ), .B1(net112098), .C0(n7384), 
        .Y(n7387) );
  BUFX16 U1734 ( .A(n9506), .Y(n4250) );
  NAND4X4 U1735 ( .A(n10072), .B(\i_MIPS/EX_MEM_1 ), .C(DCACHE_ren), .D(n8), 
        .Y(n9506) );
  NAND4X4 U1736 ( .A(n6110), .B(n6109), .C(n6108), .D(n6107), .Y(n6122) );
  NOR2X2 U1737 ( .A(n6075), .B(n6074), .Y(n6108) );
  NOR2X2 U1738 ( .A(n6043), .B(n6042), .Y(n6109) );
  INVX16 U1739 ( .A(net112372), .Y(net112366) );
  OA22X2 U1740 ( .A0(n5202), .A1(n3012), .B0(n183), .B1(n1444), .Y(n9646) );
  BUFX6 U1741 ( .A(n5173), .Y(n5167) );
  BUFX6 U1742 ( .A(n5173), .Y(n5171) );
  CLKBUFX3 U1743 ( .A(n5215), .Y(n5214) );
  CLKBUFX3 U1744 ( .A(n5176), .Y(n5156) );
  OA22X2 U1745 ( .A0(n5100), .A1(n2179), .B0(n5089), .B1(n605), .Y(n5976) );
  OA22X1 U1746 ( .A0(n5387), .A1(n793), .B0(n5324), .B1(n2355), .Y(n5977) );
  OA22X2 U1747 ( .A0(n5378), .A1(n2151), .B0(n5325), .B1(n572), .Y(n5993) );
  OA22X1 U1748 ( .A0(n4971), .A1(n808), .B0(n5016), .B1(n2371), .Y(n8696) );
  CLKBUFX8 U1749 ( .A(n5036), .Y(n5026) );
  OA22X1 U1750 ( .A0(n4981), .A1(n666), .B0(n5027), .B1(n2236), .Y(n7194) );
  OA22X1 U1751 ( .A0(n4968), .A1(n773), .B0(n5031), .B1(n2335), .Y(n9184) );
  BUFX16 U1752 ( .A(n4950), .Y(n4947) );
  OR2X2 U1753 ( .A(n4762), .B(n2208), .Y(n4178) );
  OR2X2 U1754 ( .A(n4795), .B(n2018), .Y(n4179) );
  INVX4 U1755 ( .A(n6331), .Y(n11014) );
  INVX3 U1756 ( .A(n4989), .Y(n3777) );
  OA22X2 U1757 ( .A0(n4993), .A1(n2111), .B0(n5034), .B1(n524), .Y(n6338) );
  OR2X2 U1758 ( .A(n4952), .B(n2222), .Y(n4156) );
  OA22X1 U1759 ( .A0(n4924), .A1(n1771), .B0(n4955), .B1(n3401), .Y(n6406) );
  INVX3 U1760 ( .A(n4799), .Y(n4508) );
  CLKAND2X3 U1761 ( .A(n4159), .B(n4160), .Y(n6415) );
  OR2X1 U1762 ( .A(n5032), .B(n3209), .Y(n4160) );
  OA22X2 U1763 ( .A0(n4989), .A1(n628), .B0(n5034), .B1(n3360), .Y(n6347) );
  INVX4 U1764 ( .A(n6326), .Y(n11017) );
  AND3X6 U1765 ( .A(n3778), .B(n3779), .C(n6327), .Y(n3415) );
  OR2X4 U1766 ( .A(n4933), .B(n2221), .Y(n3778) );
  OR2X4 U1767 ( .A(n4946), .B(n2436), .Y(n3779) );
  NAND4BX1 U1768 ( .AN(n7030), .B(n7029), .C(n7028), .D(n7027), .Y(n7041) );
  CLKMX2X4 U1769 ( .A(n7890), .B(n7230), .S0(net107794), .Y(n8356) );
  MX3XL U1770 ( .A(n8358), .B(n8357), .C(n8359), .S0(net112764), .S1(net107796), .Y(n8362) );
  OAI221XL U1771 ( .A0(\i_MIPS/Register/register[2][0] ), .A1(n4692), .B0(
        \i_MIPS/Register/register[10][0] ), .B1(n4687), .C0(n7591), .Y(n7599)
         );
  OA22X1 U1772 ( .A0(\i_MIPS/Register/register[6][0] ), .A1(n4683), .B0(
        \i_MIPS/Register/register[14][0] ), .B1(n4680), .Y(n7591) );
  OA22X1 U1773 ( .A0(\i_MIPS/Register/register[22][0] ), .A1(n4683), .B0(
        \i_MIPS/Register/register[30][0] ), .B1(n4680), .Y(n7600) );
  NOR4X1 U1774 ( .A(n7604), .B(n7603), .C(n7602), .D(n7601), .Y(n7605) );
  AO22X2 U1775 ( .A0(n4722), .A1(n290), .B0(n4719), .B1(n2060), .Y(n7602) );
  NOR4X1 U1776 ( .A(n7962), .B(n7961), .C(n7960), .D(n7959), .Y(n7963) );
  NOR4X1 U1777 ( .A(n7953), .B(n7952), .C(n7951), .D(n7950), .Y(n7954) );
  OA22X1 U1778 ( .A0(\i_MIPS/Register/register[6][7] ), .A1(n4682), .B0(
        \i_MIPS/Register/register[14][7] ), .B1(n4679), .Y(n7949) );
  NOR4X1 U1779 ( .A(n7676), .B(n7675), .C(n7674), .D(n7673), .Y(n7677) );
  AO22X1 U1780 ( .A0(n4712), .A1(n273), .B0(n4708), .B1(n2046), .Y(n7676) );
  NOR4X1 U1781 ( .A(n7667), .B(n7666), .C(n7665), .D(n7664), .Y(n7668) );
  AO22X1 U1782 ( .A0(n9531), .A1(n326), .B0(n4716), .B1(n478), .Y(n7666) );
  NOR4X1 U1783 ( .A(n8620), .B(n8619), .C(n8618), .D(n8617), .Y(n8621) );
  AO22X1 U1784 ( .A0(n4720), .A1(n472), .B0(n4719), .B1(n2059), .Y(n9537) );
  AO22X1 U1785 ( .A0(n9531), .A1(n477), .B0(n4715), .B1(n2069), .Y(n8908) );
  OAI221XL U1786 ( .A0(\i_MIPS/Register/register[18][23] ), .A1(n4690), .B0(
        \i_MIPS/Register/register[26][23] ), .B1(n4686), .C0(n8905), .Y(n8913)
         );
  NOR4X1 U1787 ( .A(n8900), .B(n8899), .C(n8898), .D(n8897), .Y(n8901) );
  AO22X1 U1788 ( .A0(n9531), .A1(n644), .B0(n4714), .B1(n2219), .Y(n8899) );
  CLKINVX1 U1789 ( .A(n8873), .Y(n6690) );
  AOI222X1 U1790 ( .A0(net100583), .A1(n6695), .B0(net101082), .B1(n4455), 
        .C0(n4509), .C1(net100585), .Y(n6696) );
  NAND3X2 U1791 ( .A(n8246), .B(n8245), .C(n8852), .Y(n8259) );
  NAND2X1 U1792 ( .A(n8853), .B(n9457), .Y(n8242) );
  CLKINVX1 U1793 ( .A(net102573), .Y(net102555) );
  AOI32X1 U1794 ( .A0(n3838), .A1(net107804), .A2(n8250), .B0(n9058), .B1(
        n8249), .Y(n8257) );
  OA22X1 U1795 ( .A0(net133471), .A1(n8947), .B0(net102555), .B1(net112420), 
        .Y(n8268) );
  AOI32X1 U1796 ( .A0(n8263), .A1(n4662), .A2(n9165), .B0(n8262), .B1(n9328), 
        .Y(n8270) );
  NAND2X1 U1797 ( .A(n8265), .B(n9054), .Y(n8269) );
  NAND3X4 U1798 ( .A(n4306), .B(n4307), .C(n4308), .Y(n6980) );
  OR2X4 U1799 ( .A(net104864), .B(net103076), .Y(n4306) );
  CLKINVX1 U1800 ( .A(n7620), .Y(n6981) );
  OAI2BB1X2 U1801 ( .A0N(n4672), .A1N(\i_MIPS/ALU/N303 ), .B0(n6494), .Y(
        net103710) );
  NAND2X1 U1802 ( .A(n7874), .B(n7511), .Y(n6975) );
  NOR2X1 U1803 ( .A(n9468), .B(n3843), .Y(n3764) );
  AO22X1 U1804 ( .A0(n4721), .A1(n289), .B0(n4719), .B1(n2034), .Y(n7364) );
  CLKMX2X2 U1805 ( .A(n8046), .B(n8045), .S0(net107810), .Y(net102937) );
  NAND4BX1 U1806 ( .AN(n8035), .B(n8034), .C(n8033), .D(n8032), .Y(n8046) );
  NAND4BX1 U1807 ( .AN(n8044), .B(n8043), .C(n8042), .D(n8041), .Y(n8045) );
  INVX3 U1808 ( .A(n10178), .Y(n10138) );
  AND2X2 U1809 ( .A(n7312), .B(n7311), .Y(n3766) );
  AND2X2 U1810 ( .A(n7310), .B(n7309), .Y(n3767) );
  CLKINVX1 U1811 ( .A(n6976), .Y(n7302) );
  INVX6 U1812 ( .A(n10248), .Y(n10250) );
  CLKMX2X2 U1813 ( .A(n7644), .B(n7643), .S0(net107816), .Y(n7645) );
  NOR4X1 U1814 ( .A(n7642), .B(n7641), .C(n7640), .D(n7639), .Y(n7643) );
  NOR4X1 U1815 ( .A(n7633), .B(n7632), .C(n7631), .D(n7630), .Y(n7644) );
  AO21X1 U1816 ( .A0(n7662), .A1(n7661), .B0(n5546), .Y(net112786) );
  INVX3 U1817 ( .A(net98663), .Y(net98662) );
  CLKINVX6 U1818 ( .A(n10241), .Y(n10239) );
  NAND3X4 U1819 ( .A(ICACHE_addr[16]), .B(ICACHE_addr[15]), .C(n10250), .Y(
        n10226) );
  OAI2BB1X1 U1820 ( .A0N(n8504), .A1N(n8503), .B0(n3720), .Y(n4610) );
  NAND2X1 U1821 ( .A(net112400), .B(n10839), .Y(n10577) );
  AO21X2 U1822 ( .A0(n10563), .A1(n10562), .B0(net111902), .Y(n10678) );
  OR2X4 U1823 ( .A(n9663), .B(n4247), .Y(n4313) );
  OR2X4 U1824 ( .A(n9662), .B(n5427), .Y(n4314) );
  CLKMX2X2 U1825 ( .A(n6478), .B(n6477), .S0(\i_MIPS/IR_ID[25] ), .Y(n6603) );
  NAND4BX1 U1826 ( .AN(n6467), .B(n6466), .C(n6465), .D(n6464), .Y(n6478) );
  CLKINVX1 U1827 ( .A(n11077), .Y(n4302) );
  CLKINVX1 U1828 ( .A(n10846), .Y(n10847) );
  CLKMX2X2 U1829 ( .A(n6678), .B(n6677), .S0(\i_MIPS/IR_ID[25] ), .Y(n6679) );
  NAND2BX1 U1830 ( .AN(n4247), .B(n11288), .Y(n10111) );
  NAND2X4 U1831 ( .A(n10603), .B(n10601), .Y(n10404) );
  AND2X4 U1832 ( .A(n10605), .B(n10604), .Y(n4474) );
  NAND2BX2 U1833 ( .AN(n10402), .B(n10401), .Y(n10403) );
  AOI2BB1X2 U1834 ( .A0N(n10420), .A1N(n10400), .B0(n10399), .Y(n10402) );
  OAI221XL U1835 ( .A0(\i_MIPS/Register/register[18][8] ), .A1(n4692), .B0(
        \i_MIPS/Register/register[26][8] ), .B1(n4688), .C0(n7116), .Y(n7124)
         );
  CLKMX2X2 U1836 ( .A(n6961), .B(n6960), .S0(net107812), .Y(net104887) );
  NAND4BX1 U1837 ( .AN(n6959), .B(n6958), .C(n6957), .D(n6956), .Y(n6960) );
  OR2X1 U1838 ( .A(n10579), .B(net112404), .Y(n4230) );
  AO21X2 U1839 ( .A0(n10568), .A1(n4608), .B0(net111902), .Y(n10580) );
  MXI2X1 U1840 ( .A(n9241), .B(n9240), .S0(\i_MIPS/IR_ID[25] ), .Y(n3664) );
  NOR4X1 U1841 ( .A(n9230), .B(n9229), .C(n9228), .D(n9227), .Y(n9241) );
  NAND2X1 U1842 ( .A(n10465), .B(net97874), .Y(n10823) );
  CLKINVX3 U1843 ( .A(n10338), .Y(n10316) );
  CLKMX2X2 U1844 ( .A(n8938), .B(n8937), .S0(\i_MIPS/IR_ID[25] ), .Y(n8978) );
  INVX4 U1845 ( .A(net111962), .Y(n3653) );
  INVX3 U1846 ( .A(n10388), .Y(n10592) );
  CLKINVX4 U1847 ( .A(net103806), .Y(net98363) );
  CLKMX2X2 U1848 ( .A(n7571), .B(n7570), .S0(net107816), .Y(n7572) );
  CLKINVX6 U1849 ( .A(net103504), .Y(net98216) );
  CLKMX2X2 U1850 ( .A(n7737), .B(n7736), .S0(net107816), .Y(n7738) );
  NOR4X1 U1851 ( .A(n7726), .B(n7725), .C(n7724), .D(n7723), .Y(n7737) );
  NOR4X1 U1852 ( .A(n4107), .B(n4108), .C(n4109), .D(n4110), .Y(n4106) );
  NAND2X2 U1853 ( .A(n8763), .B(n8762), .Y(n4226) );
  NAND3BX1 U1854 ( .AN(n8760), .B(net111994), .C(n8746), .Y(n8763) );
  AO22X1 U1855 ( .A0(net100583), .A1(n8745), .B0(n9275), .B1(net100585), .Y(
        n8742) );
  NAND2X1 U1856 ( .A(\i_MIPS/ALUin1[13] ), .B(n6562), .Y(n7694) );
  AOI32X1 U1857 ( .A0(net100585), .A1(\i_MIPS/ALUin1[30] ), .A2(n6598), .B0(
        n9327), .B1(n6496), .Y(n6497) );
  NAND2X4 U1858 ( .A(\i_MIPS/ALUin1[15] ), .B(n6556), .Y(n7154) );
  CLKINVX1 U1859 ( .A(n9491), .Y(n9484) );
  NAND3X1 U1860 ( .A(n4224), .B(n4225), .C(n9466), .Y(n9471) );
  AO21X1 U1861 ( .A0(n8349), .A1(net104866), .B0(n4449), .Y(n7618) );
  CLKMX2X2 U1862 ( .A(net101082), .B(net112415), .S0(n7803), .Y(n7619) );
  CLKMX2X2 U1863 ( .A(net104868), .B(n7302), .S0(net107798), .Y(n7620) );
  NOR3X1 U1864 ( .A(\i_MIPS/Reg_W[1] ), .B(\i_MIPS/Reg_W[2] ), .C(
        \i_MIPS/Reg_W[0] ), .Y(\i_MIPS/Register/n119 ) );
  NOR3X1 U1865 ( .A(\i_MIPS/Reg_W[1] ), .B(\i_MIPS/Reg_W[2] ), .C(n415), .Y(
        \i_MIPS/Register/n117 ) );
  NOR3X1 U1866 ( .A(\i_MIPS/Reg_W[0] ), .B(\i_MIPS/Reg_W[1] ), .C(n4534), .Y(
        \i_MIPS/Register/n111 ) );
  NOR3X1 U1867 ( .A(n303), .B(\i_MIPS/Reg_W[0] ), .C(n4534), .Y(
        \i_MIPS/Register/n107 ) );
  OA22X1 U1868 ( .A0(n5281), .A1(n3325), .B0(n5240), .B1(n1723), .Y(n6116) );
  CLKBUFX3 U1869 ( .A(n11039), .Y(n5526) );
  CLKINVX1 U1870 ( .A(n11372), .Y(n10215) );
  INVX3 U1871 ( .A(n11371), .Y(n10673) );
  OA22X1 U1872 ( .A0(n4747), .A1(n2161), .B0(n4790), .B1(n585), .Y(n8502) );
  OA22X1 U1873 ( .A0(n4758), .A1(n798), .B0(n4788), .B1(n2361), .Y(n9397) );
  OA22X1 U1874 ( .A0(n4818), .A1(n797), .B0(n4857), .B1(n2360), .Y(n9396) );
  OA22X1 U1875 ( .A0(n4832), .A1(n2148), .B0(n4877), .B1(n568), .Y(n6894) );
  OA22X1 U1876 ( .A0(n4826), .A1(n2093), .B0(n4871), .B1(n506), .Y(n7652) );
  INVX4 U1877 ( .A(n11417), .Y(n10917) );
  INVX3 U1878 ( .A(n11415), .Y(n10908) );
  BUFX8 U1879 ( .A(n10994), .Y(n5500) );
  INVX3 U1880 ( .A(n11476), .Y(n10139) );
  CLKINVX1 U1881 ( .A(n11462), .Y(n10288) );
  NAND4X1 U1882 ( .A(n7649), .B(n7648), .C(n7647), .D(n7646), .Y(n11460) );
  NAND4X1 U1883 ( .A(n7267), .B(n7266), .C(n7265), .D(n7264), .Y(n11457) );
  BUFX8 U1884 ( .A(n4864), .Y(n263) );
  OA22X2 U1885 ( .A0(n10782), .A1(n4245), .B0(n10785), .B1(n4246), .Y(n8313)
         );
  OAI21X2 U1886 ( .A0(n3700), .A1(n3701), .B0(n3720), .Y(n10558) );
  OAI2BB1X2 U1887 ( .A0N(n7199), .A1N(n7198), .B0(n3690), .Y(net98386) );
  OA22X2 U1888 ( .A0(n10695), .A1(n4675), .B0(n10698), .B1(n4250), .Y(n8701)
         );
  NAND2X4 U1889 ( .A(n4152), .B(n4153), .Y(net98391) );
  OA22X2 U1890 ( .A0(n10893), .A1(n4676), .B0(n10896), .B1(n4250), .Y(n7106)
         );
  OA22X2 U1891 ( .A0(n10881), .A1(n4676), .B0(n10884), .B1(n4250), .Y(n7948)
         );
  OA22X2 U1892 ( .A0(n10978), .A1(n4675), .B0(n10981), .B1(n4250), .Y(n6816)
         );
  NOR3X1 U1893 ( .A(n415), .B(\i_MIPS/Reg_W[2] ), .C(n303), .Y(
        \i_MIPS/Register/n113 ) );
  NOR3X1 U1894 ( .A(n415), .B(\i_MIPS/Reg_W[1] ), .C(n4534), .Y(
        \i_MIPS/Register/n109 ) );
  NAND4BX1 U1895 ( .AN(n6621), .B(n6620), .C(n6619), .D(n6618), .Y(n6632) );
  INVX12 U1896 ( .A(n3400), .Y(n4245) );
  NAND4BX1 U1897 ( .AN(n9206), .B(n9205), .C(n9204), .D(n9203), .Y(n9217) );
  OA22X1 U1898 ( .A0(n10868), .A1(n4675), .B0(n10871), .B1(n4250), .Y(n6658)
         );
  NOR3BX2 U1899 ( .AN(\i_MIPS/Register/n120 ), .B(\i_MIPS/Reg_W[3] ), .C(
        \i_MIPS/Reg_W[4] ), .Y(\i_MIPS/Register/n140 ) );
  NOR3X1 U1900 ( .A(\i_MIPS/Reg_W[0] ), .B(\i_MIPS/Reg_W[2] ), .C(n303), .Y(
        \i_MIPS/Register/n115 ) );
  AO21X2 U1901 ( .A0(net98780), .A1(net98781), .B0(net111902), .Y(net97687) );
  AO21X2 U1902 ( .A0(n10561), .A1(n10560), .B0(net111902), .Y(n10584) );
  INVX3 U1903 ( .A(net111968), .Y(n3773) );
  CLKMX2X2 U1904 ( .A(n7263), .B(n7262), .S0(net107816), .Y(n3738) );
  INVX3 U1905 ( .A(net104495), .Y(net98530) );
  CLKMX2X2 U1906 ( .A(n7146), .B(n7145), .S0(net107816), .Y(n7181) );
  NAND2X2 U1907 ( .A(n2212), .B(n10188), .Y(n11189) );
  OAI22X1 U1908 ( .A0(n5121), .A1(n480), .B0(n167), .B1(n2070), .Y(n4338) );
  OA22X2 U1909 ( .A0(n5303), .A1(n630), .B0(n5257), .B1(n2983), .Y(n10033) );
  OA22X2 U1910 ( .A0(n5203), .A1(n2739), .B0(n5159), .B1(n1279), .Y(n9656) );
  NAND4BX2 U1911 ( .AN(n4344), .B(n9740), .C(n9739), .D(n9738), .Y(n11293) );
  NAND4BX2 U1912 ( .AN(n4346), .B(n9593), .C(n9592), .D(n9591), .Y(n11296) );
  NAND2X1 U1913 ( .A(n11317), .B(n11319), .Y(n11318) );
  NAND4X2 U1914 ( .A(n6003), .B(n6002), .C(n6001), .D(n6000), .Y(n11322) );
  OA22X1 U1915 ( .A0(n5281), .A1(n770), .B0(n5238), .B1(n2332), .Y(n6005) );
  OA22X1 U1916 ( .A0(n5375), .A1(n790), .B0(n5355), .B1(n2352), .Y(n6016) );
  NAND2X4 U1917 ( .A(n3326), .B(n6045), .Y(n11327) );
  OA22X1 U1918 ( .A0(n5286), .A1(n777), .B0(n5239), .B1(n2339), .Y(n6045) );
  NAND4X2 U1919 ( .A(n6055), .B(n6054), .C(n6053), .D(n6052), .Y(n11328) );
  NAND4X2 U1920 ( .A(n6027), .B(n6026), .C(n6025), .D(n6024), .Y(n11330) );
  OA22X1 U1921 ( .A0(n5380), .A1(n789), .B0(n5327), .B1(n2351), .Y(n6024) );
  OA22X1 U1922 ( .A0(n5287), .A1(n2157), .B0(n5255), .B1(n580), .Y(n6081) );
  OA22X1 U1923 ( .A0(n5193), .A1(n2177), .B0(n5170), .B1(n603), .Y(n5979) );
  OA22X2 U1924 ( .A0(n5278), .A1(n2178), .B0(n5234), .B1(n604), .Y(n5978) );
  OA22X2 U1925 ( .A0(n5100), .A1(n2176), .B0(n5067), .B1(n602), .Y(n5980) );
  NAND4X2 U1926 ( .A(n6079), .B(n6078), .C(n6077), .D(n6076), .Y(n11336) );
  OA22X1 U1927 ( .A0(n5287), .A1(n2159), .B0(n5258), .B1(n582), .Y(n6077) );
  OA22X1 U1928 ( .A0(n5368), .A1(n785), .B0(n5328), .B1(n2347), .Y(n6032) );
  NAND4X2 U1929 ( .A(n6067), .B(n6066), .C(n6065), .D(n6064), .Y(n11339) );
  NAND4X2 U1930 ( .A(n6059), .B(n6058), .C(n6057), .D(n6056), .Y(n11340) );
  NAND4X2 U1931 ( .A(n6071), .B(n6070), .C(n6069), .D(n6068), .Y(n11341) );
  NAND4X2 U1932 ( .A(n6039), .B(n6038), .C(n6037), .D(n6036), .Y(n11342) );
  OA22X1 U1933 ( .A0(n5287), .A1(n2202), .B0(n5255), .B1(n485), .Y(n6089) );
  OA22X1 U1934 ( .A0(n4979), .A1(n741), .B0(n5024), .B1(n2302), .Y(n7581) );
  OA22X1 U1935 ( .A0(n4976), .A1(n2129), .B0(n185), .B1(n543), .Y(n8017) );
  OA22X1 U1936 ( .A0(n4916), .A1(n758), .B0(n4947), .B1(n2319), .Y(n8018) );
  NAND4X2 U1937 ( .A(n6891), .B(n6890), .C(n6889), .D(n6888), .Y(n11354) );
  OA22X1 U1938 ( .A0(n4759), .A1(n822), .B0(n4796), .B1(n2385), .Y(n6891) );
  OA22X1 U1939 ( .A0(n4984), .A1(n821), .B0(n5030), .B1(n2384), .Y(n6888) );
  NAND4X2 U1940 ( .A(n6810), .B(n6809), .C(n6808), .D(n6807), .Y(n11355) );
  OA22X1 U1941 ( .A0(n4984), .A1(n2294), .B0(n5030), .B1(n732), .Y(n6807) );
  NAND4X2 U1942 ( .A(n7015), .B(n7014), .C(n7013), .D(n7012), .Y(n11356) );
  OA22X1 U1943 ( .A0(n4979), .A1(n743), .B0(n5024), .B1(n2304), .Y(n7653) );
  OA22X1 U1944 ( .A0(n4747), .A1(n820), .B0(n4790), .B1(n2383), .Y(n8598) );
  OA22X2 U1945 ( .A0(n4972), .A1(n2132), .B0(n5017), .B1(n546), .Y(n8595) );
  NAND4X2 U1946 ( .A(n9298), .B(n9297), .C(n9296), .D(n9295), .Y(n11370) );
  OA22X1 U1947 ( .A0(n4755), .A1(n2414), .B0(n4788), .B1(n728), .Y(n9298) );
  NAND4X2 U1948 ( .A(n9087), .B(n9086), .C(n9085), .D(n9084), .Y(n11375) );
  OA22X1 U1949 ( .A0(n4915), .A1(n2076), .B0(n4949), .B1(n488), .Y(n9085) );
  OA22X1 U1950 ( .A0(n4744), .A1(n2416), .B0(n4789), .B1(n730), .Y(n8990) );
  OA22X1 U1951 ( .A0(n4969), .A1(n712), .B0(n5014), .B1(n2280), .Y(n8987) );
  NAND4X4 U1952 ( .A(n9393), .B(n9392), .C(n9391), .D(n9390), .Y(n11377) );
  OA22X1 U1953 ( .A0(n4827), .A1(n704), .B0(n4874), .B1(n2272), .Y(n9392) );
  OA22X1 U1954 ( .A0(n4746), .A1(n2412), .B0(n4788), .B1(n727), .Y(n9393) );
  NAND4X2 U1955 ( .A(n8498), .B(n8497), .C(n8496), .D(n8495), .Y(n11378) );
  OA22X1 U1956 ( .A0(n4747), .A1(n2204), .B0(n4790), .B1(n587), .Y(n8498) );
  OA22X1 U1957 ( .A0(n4973), .A1(n2086), .B0(n5018), .B1(n498), .Y(n8495) );
  OA22X1 U1958 ( .A0(n4749), .A1(n825), .B0(n4791), .B1(n2388), .Y(n8198) );
  NAND4X2 U1959 ( .A(n6652), .B(n6651), .C(n6650), .D(n6649), .Y(n11381) );
  OA22X1 U1960 ( .A0(n4985), .A1(n823), .B0(n5031), .B1(n2386), .Y(n6649) );
  NAND4X2 U1961 ( .A(n7588), .B(n7587), .C(n7586), .D(n7585), .Y(n11382) );
  OA22X1 U1962 ( .A0(n4754), .A1(n2410), .B0(n4792), .B1(n849), .Y(n7588) );
  OA22X1 U1963 ( .A0(n4826), .A1(n744), .B0(n4871), .B1(n2305), .Y(n7587) );
  OA22X1 U1964 ( .A0(n4979), .A1(n654), .B0(n5024), .B1(n2229), .Y(n7585) );
  NAND4X2 U1965 ( .A(n6939), .B(n6938), .C(n6937), .D(n6936), .Y(n11384) );
  NAND4X2 U1966 ( .A(n6814), .B(n6813), .C(n6812), .D(n6811), .Y(n11387) );
  OA22X1 U1967 ( .A0(n4923), .A1(n2083), .B0(n4249), .B1(n495), .Y(n6812) );
  OA22X1 U1968 ( .A0(n4984), .A1(n713), .B0(n5030), .B1(n2281), .Y(n6811) );
  OA22X1 U1969 ( .A0(n4832), .A1(n700), .B0(n4877), .B1(n2269), .Y(n6813) );
  NAND4X2 U1970 ( .A(n7946), .B(n7945), .C(n7944), .D(n7943), .Y(n11389) );
  OA22X1 U1971 ( .A0(n4818), .A1(n809), .B0(n263), .B1(n2372), .Y(n8698) );
  OA22X1 U1972 ( .A0(n4822), .A1(n800), .B0(n4868), .B1(n2363), .Y(n8106) );
  OA22X1 U1973 ( .A0(n4750), .A1(n801), .B0(n4791), .B1(n2364), .Y(n8107) );
  OA22X1 U1974 ( .A0(n4910), .A1(n2088), .B0(n4947), .B1(n501), .Y(n8893) );
  INVX3 U1975 ( .A(n11409), .Y(n10310) );
  INVX3 U1976 ( .A(n11410), .Y(n10484) );
  CLKINVX1 U1977 ( .A(n11416), .Y(n10931) );
  OA22X1 U1978 ( .A0(n4984), .A1(n772), .B0(n5030), .B1(n2334), .Y(n6884) );
  INVX3 U1979 ( .A(n11421), .Y(n10884) );
  NAND4X2 U1980 ( .A(n7432), .B(n7431), .C(n7430), .D(n7429), .Y(n11426) );
  OA22X1 U1981 ( .A0(n4830), .A1(n2140), .B0(n4861), .B1(n560), .Y(n9186) );
  OA22X1 U1982 ( .A0(n4743), .A1(n746), .B0(n4788), .B1(n2307), .Y(n9187) );
  OA22X1 U1983 ( .A0(n4915), .A1(n745), .B0(n4947), .B1(n2306), .Y(n9185) );
  NAND4X1 U1984 ( .A(n6316), .B(n6315), .C(n6314), .D(n6313), .Y(n11444) );
  OA22X1 U1985 ( .A0(n4989), .A1(n2082), .B0(n5035), .B1(n494), .Y(n6313) );
  OA22X1 U1986 ( .A0(n4984), .A1(n719), .B0(n5030), .B1(n2287), .Y(n6880) );
  OA22X1 U1987 ( .A0(n4923), .A1(n681), .B0(n4249), .B1(n2253), .Y(n6881) );
  OA22X1 U1988 ( .A0(n4832), .A1(n680), .B0(n4877), .B1(n2252), .Y(n6882) );
  CLKINVX1 U1989 ( .A(n11457), .Y(n10707) );
  INVX3 U1990 ( .A(n11460), .Y(n10741) );
  OA22X2 U1991 ( .A0(n4976), .A1(n2135), .B0(n185), .B1(n550), .Y(n8092) );
  INVX3 U1992 ( .A(n11464), .Y(n10508) );
  OA22X1 U1993 ( .A0(n4747), .A1(n2411), .B0(n4790), .B1(n725), .Y(n8590) );
  OA22X2 U1994 ( .A0(n4972), .A1(n2081), .B0(n5017), .B1(n493), .Y(n8587) );
  INVX3 U1995 ( .A(n11467), .Y(n10667) );
  OAI22XL U1996 ( .A0(n4773), .A1(n650), .B0(n4788), .B1(n2227), .Y(n4347) );
  OA22X1 U1997 ( .A0(n4744), .A1(n840), .B0(n4789), .B1(n2403), .Y(n9079) );
  OA22X1 U1998 ( .A0(n4969), .A1(n839), .B0(n5014), .B1(n2402), .Y(n9076) );
  NAND4X2 U1999 ( .A(n8982), .B(n8981), .C(n8980), .D(n8979), .Y(n11472) );
  OA22X1 U2000 ( .A0(n4744), .A1(n702), .B0(n4789), .B1(n2357), .Y(n8982) );
  OA22X1 U2001 ( .A0(n4970), .A1(n2291), .B0(n5015), .B1(n726), .Y(n8979) );
  OA22X2 U2002 ( .A0(n4924), .A1(n2146), .B0(n4955), .B1(n566), .Y(n6400) );
  NAND4X4 U2003 ( .A(n6376), .B(n6375), .C(n6374), .D(n6373), .Y(n11489) );
  OA22X2 U2004 ( .A0(n4988), .A1(n3391), .B0(n5037), .B1(n1762), .Y(n6373) );
  OA22X2 U2005 ( .A0(n4844), .A1(n3389), .B0(n4881), .B1(n1760), .Y(n6375) );
  OA22X1 U2006 ( .A0(n4836), .A1(n3008), .B0(n4882), .B1(n584), .Y(n6345) );
  OA22X2 U2007 ( .A0(n4764), .A1(n3005), .B0(n4796), .B1(n577), .Y(n6346) );
  OA22X2 U2008 ( .A0(n4926), .A1(n2999), .B0(n4950), .B1(n557), .Y(n6344) );
  OA22X2 U2009 ( .A0(n4986), .A1(n635), .B0(n5032), .B1(n3353), .Y(n6405) );
  OA22X2 U2010 ( .A0(n4762), .A1(n2987), .B0(n4795), .B1(n540), .Y(n6408) );
  OA22X2 U2011 ( .A0(n4834), .A1(n2652), .B0(n4879), .B1(n590), .Y(n6407) );
  OA22X2 U2012 ( .A0(n4926), .A1(n3376), .B0(n4950), .B1(n1747), .Y(n6354) );
  OA22X2 U2013 ( .A0(n4764), .A1(n3366), .B0(n4796), .B1(n1737), .Y(n6356) );
  OA22X1 U2014 ( .A0(n4834), .A1(n2997), .B0(n4879), .B1(n555), .Y(n6434) );
  BUFX16 U2015 ( .A(n11511), .Y(n5551) );
  CLKINVX1 U2016 ( .A(n10368), .Y(n10378) );
  NAND4BX1 U2017 ( .AN(n7863), .B(n7862), .C(n7861), .D(n7860), .Y(net103252)
         );
  NAND4BX2 U2018 ( .AN(n7872), .B(n7871), .C(n7870), .D(n7869), .Y(net103253)
         );
  CLKMX2X2 U2019 ( .A(net104410), .B(net104411), .S0(net107812), .Y(net104407)
         );
  NAND4BX1 U2020 ( .AN(n7217), .B(n7216), .C(n7215), .D(n7214), .Y(net104411)
         );
  NAND4BX1 U2021 ( .AN(n8812), .B(n8811), .C(n8810), .D(n8809), .Y(n8823) );
  AOI2BB1X1 U2022 ( .A0N(n8658), .A1N(n9461), .B0(n8657), .Y(n8659) );
  NOR4X4 U2023 ( .A(n9174), .B(n9173), .C(n9172), .D(n9171), .Y(n9175) );
  INVX4 U2024 ( .A(n3913), .Y(n10652) );
  CLKMX2X2 U2025 ( .A(net105048), .B(net105049), .S0(net107812), .Y(net105045)
         );
  NAND4BX1 U2026 ( .AN(n6906), .B(n6905), .C(n6904), .D(n6903), .Y(net105048)
         );
  NAND4BX1 U2027 ( .AN(n6915), .B(n6914), .C(n6913), .D(n6912), .Y(net105049)
         );
  CLKMX2X2 U2028 ( .A(n9323), .B(n9322), .S0(net107810), .Y(n9325) );
  INVX3 U2029 ( .A(n10549), .Y(n10556) );
  CLKINVX1 U2030 ( .A(n11110), .Y(n11108) );
  NAND4X2 U2031 ( .A(n6283), .B(n6282), .C(n6281), .D(n6280), .Y(n9560) );
  INVX3 U2032 ( .A(n3818), .Y(n3819) );
  INVX3 U2033 ( .A(net98393), .Y(net104106) );
  CLKMX2X2 U2034 ( .A(net104254), .B(net104255), .S0(net107812), .Y(net104251)
         );
  NAND4BX1 U2035 ( .AN(n7290), .B(n7289), .C(n7288), .D(n7287), .Y(net104254)
         );
  INVX3 U2036 ( .A(n3783), .Y(n3784) );
  INVX3 U2037 ( .A(n10236), .Y(n10587) );
  INVX1 U2038 ( .A(n10406), .Y(n10412) );
  CLKINVX1 U2039 ( .A(n10828), .Y(n10340) );
  CLKINVX1 U2040 ( .A(n10804), .Y(n10802) );
  INVX3 U2041 ( .A(n10357), .Y(n10579) );
  CLKINVX1 U2042 ( .A(n10425), .Y(n10423) );
  CLKINVX1 U2043 ( .A(n10595), .Y(n10593) );
  XOR3X1 U2044 ( .A(net112400), .B(n10650), .C(n10634), .Y(n10645) );
  NAND2BX2 U2045 ( .AN(n5425), .B(n11252), .Y(n9948) );
  NAND2BX2 U2046 ( .AN(n5425), .B(n11254), .Y(n9908) );
  NAND4X4 U2047 ( .A(n10111), .B(n10110), .C(n10109), .D(n10108), .Y(n10368)
         );
  NAND2BX2 U2048 ( .AN(n5427), .B(n11192), .Y(n10109) );
  NAND2BX2 U2049 ( .AN(n5429), .B(n11224), .Y(n10108) );
  NAND2BX2 U2050 ( .AN(n5425), .B(n11256), .Y(n10110) );
  NAND2BX2 U2051 ( .AN(n5425), .B(n11255), .Y(n9932) );
  XOR3X1 U2052 ( .A(n10423), .B(n4386), .C(n10422), .Y(n10426) );
  XOR2X2 U2053 ( .A(n10254), .B(n10531), .Y(n10255) );
  CLKINVX1 U2054 ( .A(n10591), .Y(n10597) );
  OAI222X1 U2055 ( .A0(n7706), .A1(n7234), .B0(net133471), .B1(n6966), .C0(
        net103060), .C1(n7978), .Y(n6777) );
  BUFX16 U2056 ( .A(n4382), .Y(n4664) );
  INVX3 U2057 ( .A(n9979), .Y(n8429) );
  OR2X2 U2058 ( .A(net102790), .B(net111624), .Y(n3702) );
  AOI2BB2X2 U2059 ( .B0(n7886), .B1(n7885), .A0N(n7884), .A1N(n7883), .Y(n7909) );
  INVX3 U2060 ( .A(n4301), .Y(n10176) );
  AOI2BB1X1 U2061 ( .A0N(net137891), .A1N(n7420), .B0(n7419), .Y(n7421) );
  CLKINVX1 U2062 ( .A(n3725), .Y(n7422) );
  NAND3BX1 U2063 ( .AN(n8562), .B(n8561), .C(net111994), .Y(n8563) );
  CLKINVX1 U2064 ( .A(\i_MIPS/ID_EX[86] ), .Y(n6444) );
  OAI33X1 U2065 ( .A0(net101257), .A1(n9045), .A2(n9350), .B0(net101257), .B1(
        n9044), .B2(n9052), .Y(n9073) );
  AO22X2 U2066 ( .A0(n5528), .A1(DCACHE_addr[12]), .B0(n5526), .B1(n11490), 
        .Y(n11024) );
  AO22X2 U2067 ( .A0(n5544), .A1(ICACHE_addr[16]), .B0(n239), .B1(n11331), .Y(
        n11153) );
  AO22X2 U2068 ( .A0(n5544), .A1(ICACHE_addr[12]), .B0(n239), .B1(n11327), .Y(
        n11148) );
  AO22X2 U2069 ( .A0(n5544), .A1(ICACHE_addr[21]), .B0(n240), .B1(n11336), .Y(
        n11154) );
  AO22X2 U2070 ( .A0(n5544), .A1(ICACHE_addr[28]), .B0(n240), .B1(n11343), .Y(
        n11150) );
  AO22X2 U2071 ( .A0(n5544), .A1(ICACHE_addr[26]), .B0(n240), .B1(n11341), .Y(
        n11144) );
  AO22X2 U2072 ( .A0(n5544), .A1(ICACHE_addr[24]), .B0(n240), .B1(n11339), .Y(
        n11145) );
  AO22X2 U2073 ( .A0(n5543), .A1(ICACHE_addr[8]), .B0(n240), .B1(n11323), .Y(
        n11135) );
  AO22X2 U2074 ( .A0(n5543), .A1(ICACHE_addr[23]), .B0(n239), .B1(n11338), .Y(
        n11137) );
  AO22X2 U2075 ( .A0(n5543), .A1(n3781), .B0(n239), .B1(n11321), .Y(n11134) );
  AO22X2 U2076 ( .A0(n5543), .A1(ICACHE_addr[18]), .B0(n240), .B1(n11333), .Y(
        n11132) );
  AO22X2 U2077 ( .A0(mem_rdata_I[30]), .A1(n5542), .B0(n252), .B1(n11216), .Y(
        n6211) );
  AO22X2 U2078 ( .A0(mem_rdata_I[11]), .A1(n5539), .B0(n250), .B1(n11197), .Y(
        n9751) );
  AO22X2 U2079 ( .A0(mem_rdata_I[5]), .A1(n5537), .B0(n253), .B1(n11191), .Y(
        n9924) );
  AO22X2 U2080 ( .A0(mem_rdata_I[0]), .A1(n5543), .B0(n249), .B1(n11186), .Y(
        n6151) );
  AO22X2 U2081 ( .A0(mem_rdata_I[62]), .A1(n5542), .B0(n252), .B1(n11248), .Y(
        n6216) );
  AO22X2 U2082 ( .A0(mem_rdata_I[44]), .A1(n5539), .B0(n253), .B1(n11230), .Y(
        n9779) );
  AO22X2 U2083 ( .A0(mem_rdata_I[43]), .A1(n5539), .B0(n253), .B1(n11229), .Y(
        n9756) );
  AO22X2 U2084 ( .A0(mem_rdata_I[34]), .A1(n5536), .B0(n252), .B1(n11220), .Y(
        n11105) );
  AO22X2 U2085 ( .A0(mem_rdata_I[66]), .A1(n5536), .B0(n251), .B1(n11252), .Y(
        n11103) );
  AO22X2 U2086 ( .A0(mem_rdata_I[125]), .A1(n5542), .B0(n249), .B1(n11311), 
        .Y(n6221) );
  AO22X2 U2087 ( .A0(mem_rdata_I[107]), .A1(n5539), .B0(n249), .B1(n11293), 
        .Y(n9741) );
  AO22X2 U2088 ( .A0(mem_rdata_I[100]), .A1(n5543), .B0(n250), .B1(n11286), 
        .Y(n6131) );
  AO22X2 U2089 ( .A0(mem_rdata_I[96]), .A1(n5543), .B0(n252), .B1(n11282), .Y(
        n6141) );
  NAND2X1 U2090 ( .A(n4303), .B(n9974), .Y(n9983) );
  AO22X2 U2091 ( .A0(n5528), .A1(DCACHE_addr[28]), .B0(n5526), .B1(n11506), 
        .Y(n11021) );
  AO22X2 U2092 ( .A0(n5528), .A1(DCACHE_addr[27]), .B0(n5527), .B1(n11505), 
        .Y(n11029) );
  AO22X2 U2093 ( .A0(n5528), .A1(n12939), .B0(n5527), .B1(n11496), .Y(n11035)
         );
  INVX3 U2094 ( .A(n3833), .Y(n3834) );
  CLKINVX1 U2095 ( .A(n11036), .Y(n3833) );
  AO22X2 U2096 ( .A0(n5528), .A1(n12952), .B0(n5526), .B1(n11483), .Y(n11019)
         );
  AOI222X1 U2097 ( .A0(n5505), .A1(n11367), .B0(mem_rdata_D[17]), .B1(n235), 
        .C0(n12970), .C1(n5502), .Y(n10770) );
  AOI222X1 U2098 ( .A0(n5505), .A1(n11365), .B0(mem_rdata_D[15]), .B1(n232), 
        .C0(n12972), .C1(n5502), .Y(n10759) );
  MXI2X2 U2099 ( .A(n10702), .B(n10701), .S0(n5517), .Y(n10703) );
  NAND2X1 U2100 ( .A(n10148), .B(n5513), .Y(n4195) );
  NAND2X1 U2101 ( .A(n10149), .B(n4232), .Y(n4194) );
  NAND2X1 U2102 ( .A(n10690), .B(n5517), .Y(n4197) );
  NAND2X1 U2103 ( .A(n10500), .B(n5516), .Y(n4200) );
  NAND2X1 U2104 ( .A(n10501), .B(n4198), .Y(n4199) );
  NAND2X1 U2105 ( .A(n10786), .B(n4232), .Y(n4233) );
  AOI222XL U2106 ( .A0(n5511), .A1(n11406), .B0(mem_rdata_D[56]), .B1(n235), 
        .C0(n12963), .C1(n5507), .Y(n10786) );
  AOI222X1 U2107 ( .A0(n5510), .A1(n11404), .B0(mem_rdata_D[54]), .B1(n234), 
        .C0(n12965), .C1(n5506), .Y(n10219) );
  NAND2X1 U2108 ( .A(n10676), .B(n5517), .Y(n4236) );
  NAND2X1 U2109 ( .A(n10677), .B(n4232), .Y(n4235) );
  NAND2X1 U2110 ( .A(n10663), .B(n5516), .Y(n4203) );
  MXI2X2 U2111 ( .A(n11005), .B(n11004), .S0(n5523), .Y(n11006) );
  NAND2X1 U2112 ( .A(n10517), .B(n5516), .Y(n4239) );
  NAND2X1 U2113 ( .A(n10772), .B(n5519), .Y(n4206) );
  NAND2X1 U2114 ( .A(n10773), .B(n4204), .Y(n4205) );
  NAND2X1 U2115 ( .A(n10761), .B(n5519), .Y(n4209) );
  NAND2X1 U2116 ( .A(n10762), .B(n4207), .Y(n4208) );
  NAND2X1 U2117 ( .A(n10750), .B(n5519), .Y(n4241) );
  NAND2X1 U2118 ( .A(n10751), .B(n4190), .Y(n4240) );
  NAND2X1 U2119 ( .A(n10739), .B(n5518), .Y(n4211) );
  NAND2X1 U2120 ( .A(n10740), .B(n4232), .Y(n4210) );
  NAND2X1 U2121 ( .A(n10728), .B(n5518), .Y(n4213) );
  NAND2X1 U2122 ( .A(n10729), .B(n4232), .Y(n4212) );
  NAND2X1 U2123 ( .A(n10716), .B(n5518), .Y(n4243) );
  NAND2X1 U2124 ( .A(n10717), .B(n4190), .Y(n4242) );
  AOI222XL U2125 ( .A0(n5511), .A1(n11393), .B0(mem_rdata_D[43]), .B1(n232), 
        .C0(n12976), .C1(n5507), .Y(n10717) );
  NAND2X1 U2126 ( .A(n10086), .B(n5513), .Y(n4215) );
  NAND2X1 U2127 ( .A(n10087), .B(n4190), .Y(n4214) );
  AOI222X1 U2128 ( .A0(n5512), .A1(n11385), .B0(mem_rdata_D[35]), .B1(n233), 
        .C0(n12984), .C1(n5507), .Y(n10924) );
  AOI222X1 U2129 ( .A0(n5512), .A1(n11383), .B0(mem_rdata_D[33]), .B1(n233), 
        .C0(n12986), .C1(n5507), .Y(n10915) );
  AOI222X1 U2130 ( .A0(n5499), .A1(n11443), .B0(mem_rdata_D[93]), .B1(n233), 
        .C0(n12958), .C1(n5497), .Y(n10685) );
  AOI222X1 U2131 ( .A0(n5499), .A1(n11438), .B0(mem_rdata_D[88]), .B1(n236), 
        .C0(n12963), .C1(n5497), .Y(n10780) );
  AOI222X1 U2132 ( .A0(n5498), .A1(n11436), .B0(mem_rdata_D[86]), .B1(n236), 
        .C0(n12965), .C1(n4385), .Y(n10213) );
  AOI222X1 U2133 ( .A0(n5498), .A1(n11434), .B0(mem_rdata_D[84]), .B1(n235), 
        .C0(n12967), .C1(n4385), .Y(n10658) );
  MXI2X2 U2134 ( .A(n10512), .B(n10511), .S0(n5516), .Y(n10513) );
  AOI222X1 U2135 ( .A0(n5499), .A1(n11431), .B0(mem_rdata_D[81]), .B1(n234), 
        .C0(n12970), .C1(n5497), .Y(n10767) );
  AOI222X1 U2136 ( .A0(n5499), .A1(n11429), .B0(mem_rdata_D[79]), .B1(n234), 
        .C0(n12972), .C1(n5497), .Y(n10756) );
  AOI222X1 U2137 ( .A0(n5499), .A1(n11427), .B0(mem_rdata_D[77]), .B1(n235), 
        .C0(n12974), .C1(n5497), .Y(n10734) );
  CLKBUFX3 U2138 ( .A(n10711), .Y(n3709) );
  AOI222X1 U2139 ( .A0(n5499), .A1(n11423), .B0(mem_rdata_D[73]), .B1(n232), 
        .C0(n12978), .C1(n5497), .Y(n10699) );
  AOI222X1 U2140 ( .A0(n5498), .A1(n11420), .B0(mem_rdata_D[70]), .B1(n236), 
        .C0(n12981), .C1(n4385), .Y(n10074) );
  AOI222X1 U2141 ( .A0(n5495), .A1(n11469), .B0(mem_rdata_D[119]), .B1(n234), 
        .C0(n12964), .C1(n5494), .Y(n10941) );
  MXI2X2 U2142 ( .A(n10655), .B(n10654), .S0(n5516), .Y(n10656) );
  AOI222X1 U2143 ( .A0(n5496), .A1(n11458), .B0(mem_rdata_D[108]), .B1(n232), 
        .C0(n12975), .C1(n5493), .Y(n10720) );
  AOI222X1 U2144 ( .A0(n5495), .A1(n11448), .B0(mem_rdata_D[98]), .B1(n234), 
        .C0(n12985), .C1(n5494), .Y(n10929) );
  AOI222X1 U2145 ( .A0(n5496), .A1(n11447), .B0(mem_rdata_D[97]), .B1(n235), 
        .C0(n12986), .C1(n5494), .Y(n10906) );
  CLKMX2X2 U2146 ( .A(n9016), .B(n9015), .S0(net107810), .Y(n9018) );
  CLKMX2X2 U2147 ( .A(n8524), .B(n8523), .S0(net107810), .Y(n8527) );
  CLKMX2X2 U2148 ( .A(n9113), .B(n9112), .S0(net107810), .Y(n9116) );
  NAND4BX1 U2149 ( .AN(n9102), .B(n9101), .C(n9100), .D(n9099), .Y(n9113) );
  OR2X2 U2150 ( .A(n8226), .B(net111622), .Y(n3691) );
  NOR4X1 U2151 ( .A(n9346), .B(n9345), .C(n9344), .D(n9343), .Y(n9360) );
  NAND3BX2 U2152 ( .AN(n9430), .B(n5547), .C(net111646), .Y(n9431) );
  CLKMX2X2 U2153 ( .A(n9428), .B(n9427), .S0(net107810), .Y(n9429) );
  NAND2BX1 U2154 ( .AN(n5429), .B(n11248), .Y(n6284) );
  NAND2BX1 U2155 ( .AN(n4247), .B(n11312), .Y(n6287) );
  AO22X2 U2156 ( .A0(mem_rdata_I[59]), .A1(n5535), .B0(n251), .B1(n11245), .Y(
        n11160) );
  AO22X2 U2157 ( .A0(mem_rdata_I[54]), .A1(n5538), .B0(n253), .B1(n11240), .Y(
        n9877) );
  AO22X2 U2158 ( .A0(mem_rdata_I[49]), .A1(n5536), .B0(n250), .B1(n11235), .Y(
        n10172) );
  AO22X2 U2159 ( .A0(mem_rdata_I[91]), .A1(n5535), .B0(n249), .B1(n11277), .Y(
        n11158) );
  AO22X2 U2160 ( .A0(mem_rdata_I[88]), .A1(n5539), .B0(n251), .B1(n11274), .Y(
        n9793) );
  AO22X2 U2161 ( .A0(mem_rdata_I[81]), .A1(n5536), .B0(n250), .B1(n11267), .Y(
        n10162) );
  AO22X2 U2162 ( .A0(mem_rdata_I[123]), .A1(n5535), .B0(n250), .B1(n11309), 
        .Y(n11157) );
  AO22X2 U2163 ( .A0(mem_rdata_I[119]), .A1(n5539), .B0(n252), .B1(n11305), 
        .Y(n9829) );
  AO22X2 U2164 ( .A0(mem_rdata_I[118]), .A1(n5538), .B0(n253), .B1(n11304), 
        .Y(n9865) );
  AO22X2 U2165 ( .A0(mem_rdata_I[117]), .A1(n5538), .B0(n251), .B1(n11303), 
        .Y(n9849) );
  AO22X2 U2166 ( .A0(mem_rdata_I[112]), .A1(n5539), .B0(n252), .B1(n11298), 
        .Y(n9717) );
  NAND2X4 U2167 ( .A(\i_MIPS/BranchAddr[0] ), .B(n4315), .Y(n10524) );
  CLKINVX1 U2168 ( .A(n10604), .Y(n10603) );
  INVX4 U2169 ( .A(net107802), .Y(net107796) );
  AOI222X1 U2170 ( .A0(n4422), .A1(n4587), .B0(n6848), .B1(n6847), .C0(n6846), 
        .C1(n6845), .Y(n6857) );
  OAI222X1 U2171 ( .A0(n9248), .A1(n7234), .B0(net133471), .B1(n6844), .C0(
        net103060), .C1(n7062), .Y(n6858) );
  BUFX16 U2172 ( .A(n12932), .Y(DCACHE_addr[25]) );
  BUFX16 U2173 ( .A(n12930), .Y(DCACHE_addr[27]) );
  BUFX12 U2174 ( .A(n12927), .Y(mem_wdata_I[1]) );
  BUFX12 U2175 ( .A(n12926), .Y(mem_wdata_I[4]) );
  BUFX12 U2176 ( .A(n12925), .Y(mem_wdata_I[5]) );
  BUFX12 U2177 ( .A(n12924), .Y(mem_wdata_I[6]) );
  BUFX12 U2178 ( .A(n12923), .Y(mem_wdata_I[7]) );
  BUFX12 U2179 ( .A(n12922), .Y(mem_wdata_I[8]) );
  BUFX12 U2180 ( .A(n12921), .Y(mem_wdata_I[9]) );
  BUFX12 U2181 ( .A(n12920), .Y(mem_wdata_I[10]) );
  BUFX12 U2182 ( .A(n12919), .Y(mem_wdata_I[11]) );
  BUFX12 U2183 ( .A(n12918), .Y(mem_wdata_I[12]) );
  BUFX12 U2184 ( .A(n12917), .Y(mem_wdata_I[13]) );
  INVX12 U2185 ( .A(n3953), .Y(mem_wdata_I[16]) );
  OR2X1 U2186 ( .A(n4655), .B(n3954), .Y(n3953) );
  INVX12 U2187 ( .A(n3959), .Y(mem_wdata_I[17]) );
  OR2X1 U2188 ( .A(n4655), .B(n3960), .Y(n3959) );
  BUFX12 U2189 ( .A(n12916), .Y(mem_wdata_I[18]) );
  BUFX12 U2190 ( .A(n12915), .Y(mem_wdata_I[19]) );
  BUFX12 U2191 ( .A(n12914), .Y(mem_wdata_I[20]) );
  BUFX12 U2192 ( .A(n12913), .Y(mem_wdata_I[21]) );
  BUFX12 U2193 ( .A(n12912), .Y(mem_wdata_I[22]) );
  BUFX12 U2194 ( .A(n12911), .Y(mem_wdata_I[23]) );
  BUFX12 U2195 ( .A(n12910), .Y(mem_wdata_I[24]) );
  BUFX12 U2196 ( .A(n12909), .Y(mem_wdata_I[25]) );
  BUFX12 U2197 ( .A(n12908), .Y(mem_wdata_I[26]) );
  BUFX12 U2198 ( .A(n12907), .Y(mem_wdata_I[27]) );
  BUFX12 U2199 ( .A(n12906), .Y(mem_wdata_I[28]) );
  BUFX12 U2200 ( .A(n12905), .Y(mem_wdata_I[29]) );
  BUFX12 U2201 ( .A(n12904), .Y(mem_wdata_I[30]) );
  BUFX12 U2202 ( .A(n12903), .Y(mem_wdata_I[31]) );
  BUFX12 U2203 ( .A(n12902), .Y(mem_wdata_I[32]) );
  BUFX12 U2204 ( .A(n12901), .Y(mem_wdata_I[33]) );
  BUFX12 U2205 ( .A(n12900), .Y(mem_wdata_I[35]) );
  BUFX12 U2206 ( .A(n12899), .Y(mem_wdata_I[36]) );
  BUFX12 U2207 ( .A(n12898), .Y(mem_wdata_I[37]) );
  BUFX12 U2208 ( .A(n12897), .Y(mem_wdata_I[38]) );
  BUFX12 U2209 ( .A(n12896), .Y(mem_wdata_I[39]) );
  BUFX12 U2210 ( .A(n12895), .Y(mem_wdata_I[40]) );
  BUFX12 U2211 ( .A(n12894), .Y(mem_wdata_I[42]) );
  BUFX12 U2212 ( .A(n12893), .Y(mem_wdata_I[43]) );
  BUFX12 U2213 ( .A(n12892), .Y(mem_wdata_I[44]) );
  BUFX12 U2214 ( .A(n12891), .Y(mem_wdata_I[45]) );
  BUFX12 U2215 ( .A(n12890), .Y(mem_wdata_I[46]) );
  BUFX16 U2216 ( .A(n12889), .Y(mem_wdata_I[49]) );
  BUFX16 U2217 ( .A(n12888), .Y(mem_wdata_I[52]) );
  BUFX16 U2218 ( .A(n12887), .Y(mem_wdata_I[53]) );
  BUFX16 U2219 ( .A(n12886), .Y(mem_wdata_I[55]) );
  BUFX16 U2220 ( .A(n12885), .Y(mem_wdata_I[56]) );
  BUFX12 U2221 ( .A(n12884), .Y(mem_wdata_I[57]) );
  BUFX16 U2222 ( .A(n12883), .Y(mem_wdata_I[58]) );
  BUFX16 U2223 ( .A(n12882), .Y(mem_wdata_I[59]) );
  BUFX16 U2224 ( .A(n12881), .Y(mem_wdata_I[60]) );
  BUFX16 U2225 ( .A(n12880), .Y(mem_wdata_I[61]) );
  BUFX16 U2226 ( .A(n12879), .Y(mem_wdata_I[62]) );
  BUFX16 U2227 ( .A(n12878), .Y(mem_wdata_I[63]) );
  BUFX16 U2228 ( .A(n12877), .Y(mem_wdata_I[64]) );
  BUFX16 U2229 ( .A(n12876), .Y(mem_wdata_I[65]) );
  BUFX16 U2230 ( .A(n12875), .Y(mem_wdata_I[67]) );
  BUFX16 U2231 ( .A(n12874), .Y(mem_wdata_I[68]) );
  BUFX12 U2232 ( .A(n12873), .Y(mem_wdata_I[69]) );
  BUFX16 U2233 ( .A(n12872), .Y(mem_wdata_I[70]) );
  BUFX16 U2234 ( .A(n12871), .Y(mem_wdata_I[71]) );
  BUFX16 U2235 ( .A(n12869), .Y(mem_wdata_I[73]) );
  BUFX12 U2236 ( .A(n12867), .Y(mem_wdata_I[75]) );
  BUFX16 U2237 ( .A(n12866), .Y(mem_wdata_I[76]) );
  BUFX16 U2238 ( .A(n12865), .Y(mem_wdata_I[77]) );
  BUFX16 U2239 ( .A(n12863), .Y(mem_wdata_I[79]) );
  BUFX16 U2240 ( .A(n12862), .Y(mem_wdata_I[80]) );
  BUFX12 U2241 ( .A(n12861), .Y(mem_wdata_I[81]) );
  BUFX16 U2242 ( .A(n12860), .Y(mem_wdata_I[82]) );
  BUFX16 U2243 ( .A(n12859), .Y(mem_wdata_I[83]) );
  BUFX16 U2244 ( .A(n12857), .Y(mem_wdata_I[85]) );
  BUFX16 U2245 ( .A(n12856), .Y(mem_wdata_I[86]) );
  BUFX16 U2246 ( .A(n12854), .Y(mem_wdata_I[88]) );
  BUFX16 U2247 ( .A(n12853), .Y(mem_wdata_I[89]) );
  BUFX12 U2248 ( .A(n12852), .Y(mem_wdata_I[90]) );
  BUFX16 U2249 ( .A(n12851), .Y(mem_wdata_I[91]) );
  BUFX16 U2250 ( .A(n12850), .Y(mem_wdata_I[92]) );
  BUFX12 U2251 ( .A(n12849), .Y(mem_wdata_I[93]) );
  BUFX16 U2252 ( .A(n12848), .Y(mem_wdata_I[94]) );
  BUFX16 U2253 ( .A(n12847), .Y(mem_wdata_I[95]) );
  BUFX16 U2254 ( .A(n12845), .Y(mem_wdata_I[97]) );
  BUFX16 U2255 ( .A(n12844), .Y(mem_wdata_I[98]) );
  BUFX12 U2256 ( .A(n12843), .Y(mem_wdata_I[99]) );
  BUFX16 U2257 ( .A(n12842), .Y(mem_wdata_I[100]) );
  BUFX16 U2258 ( .A(n12840), .Y(mem_wdata_I[103]) );
  BUFX16 U2259 ( .A(n12839), .Y(mem_wdata_I[104]) );
  BUFX16 U2260 ( .A(n12837), .Y(mem_wdata_I[106]) );
  BUFX16 U2261 ( .A(n12836), .Y(mem_wdata_I[109]) );
  BUFX12 U2262 ( .A(n12835), .Y(mem_wdata_I[111]) );
  BUFX16 U2263 ( .A(n12834), .Y(mem_wdata_I[112]) );
  BUFX16 U2264 ( .A(n12833), .Y(mem_wdata_I[113]) );
  BUFX16 U2265 ( .A(n12831), .Y(mem_wdata_I[115]) );
  BUFX16 U2266 ( .A(n12830), .Y(mem_wdata_I[116]) );
  BUFX16 U2267 ( .A(n12828), .Y(mem_wdata_I[118]) );
  BUFX16 U2268 ( .A(n12827), .Y(mem_wdata_I[119]) );
  BUFX16 U2269 ( .A(n12825), .Y(mem_wdata_I[121]) );
  BUFX16 U2270 ( .A(n12824), .Y(mem_wdata_I[122]) );
  BUFX12 U2271 ( .A(n12823), .Y(mem_wdata_I[123]) );
  BUFX16 U2272 ( .A(n12822), .Y(mem_wdata_I[124]) );
  BUFX16 U2273 ( .A(n12821), .Y(mem_wdata_I[125]) );
  AOI22X1 U2274 ( .A0(n3781), .A1(n11512), .B0(mem_write_I), .B1(n11321), .Y(
        n410) );
  AOI22X1 U2275 ( .A0(ICACHE_addr[9]), .A1(n11512), .B0(n5556), .B1(n11324), 
        .Y(n411) );
  AOI22X1 U2276 ( .A0(ICACHE_addr[12]), .A1(n11512), .B0(mem_write_I), .B1(
        n11327), .Y(n412) );
  AO22X1 U2277 ( .A0(ICACHE_addr[14]), .A1(n11512), .B0(n4656), .B1(n11329), 
        .Y(n12819) );
  BUFX20 U2278 ( .A(n5554), .Y(mem_write_I) );
  INVX12 U2279 ( .A(n3867), .Y(mem_wdata_D[7]) );
  INVX12 U2280 ( .A(n3872), .Y(mem_wdata_D[11]) );
  INVX12 U2281 ( .A(n3882), .Y(mem_wdata_D[13]) );
  INVX12 U2282 ( .A(n3878), .Y(mem_wdata_D[15]) );
  INVX12 U2283 ( .A(n3742), .Y(mem_wdata_D[36]) );
  OR2X1 U2284 ( .A(n4649), .B(n10975), .Y(n3742) );
  INVX12 U2285 ( .A(n3871), .Y(mem_wdata_D[40]) );
  INVX12 U2286 ( .A(n3874), .Y(mem_wdata_D[46]) );
  INVX12 U2287 ( .A(n3668), .Y(mem_wdata_D[56]) );
  INVX12 U2288 ( .A(n3870), .Y(mem_wdata_D[58]) );
  INVX12 U2289 ( .A(n3670), .Y(mem_wdata_D[59]) );
  OR2X1 U2290 ( .A(n4649), .B(n10310), .Y(n3670) );
  INVX12 U2291 ( .A(n3669), .Y(mem_wdata_D[60]) );
  OR2X1 U2292 ( .A(n4649), .B(n10484), .Y(n3669) );
  INVX12 U2293 ( .A(n3877), .Y(mem_wdata_D[61]) );
  INVX12 U2294 ( .A(n3672), .Y(mem_wdata_D[62]) );
  OR2X1 U2295 ( .A(n4649), .B(n10148), .Y(n3672) );
  INVX12 U2296 ( .A(n3671), .Y(mem_wdata_D[63]) );
  INVX12 U2297 ( .A(n3883), .Y(mem_wdata_D[64]) );
  INVX12 U2298 ( .A(n3674), .Y(mem_wdata_D[65]) );
  INVX12 U2299 ( .A(n3673), .Y(mem_wdata_D[66]) );
  OR2X1 U2300 ( .A(n4649), .B(n10931), .Y(n3673) );
  INVX12 U2301 ( .A(n3710), .Y(mem_wdata_D[71]) );
  OR2X1 U2302 ( .A(n4649), .B(n10884), .Y(n3710) );
  INVX12 U2303 ( .A(n3675), .Y(mem_wdata_D[72]) );
  OR2X1 U2304 ( .A(n4649), .B(n10896), .Y(n3675) );
  INVX12 U2305 ( .A(n3717), .Y(mem_wdata_D[74]) );
  INVX12 U2306 ( .A(n3711), .Y(mem_wdata_D[75]) );
  INVX12 U2307 ( .A(n3723), .Y(mem_wdata_D[77]) );
  INVX12 U2308 ( .A(n3719), .Y(mem_wdata_D[78]) );
  INVX12 U2309 ( .A(n3724), .Y(mem_wdata_D[81]) );
  INVX12 U2310 ( .A(n3727), .Y(mem_wdata_D[83]) );
  INVX12 U2311 ( .A(n3739), .Y(mem_wdata_D[86]) );
  OR2X1 U2312 ( .A(n4649), .B(n10212), .Y(n3739) );
  INVX12 U2313 ( .A(n3728), .Y(mem_wdata_D[87]) );
  INVX12 U2314 ( .A(n3743), .Y(mem_wdata_D[89]) );
  INVX12 U2315 ( .A(n3740), .Y(mem_wdata_D[90]) );
  OR2X1 U2316 ( .A(n4649), .B(n10272), .Y(n3740) );
  INVX12 U2317 ( .A(n3868), .Y(mem_wdata_D[92]) );
  INVX12 U2318 ( .A(n3744), .Y(mem_wdata_D[93]) );
  INVX12 U2319 ( .A(n3873), .Y(mem_wdata_D[95]) );
  INVX12 U2320 ( .A(n3869), .Y(mem_wdata_D[96]) );
  INVX12 U2321 ( .A(n3881), .Y(mem_wdata_D[99]) );
  INVX12 U2322 ( .A(n3880), .Y(mem_wdata_D[101]) );
  INVX12 U2323 ( .A(n3876), .Y(mem_wdata_D[102]) );
  INVX12 U2324 ( .A(n1975), .Y(mem_wdata_D[105]) );
  INVX12 U2325 ( .A(n1976), .Y(mem_wdata_D[108]) );
  INVX12 U2326 ( .A(n1981), .Y(mem_wdata_D[111]) );
  INVX12 U2327 ( .A(n1982), .Y(mem_wdata_D[120]) );
  INVX12 U2328 ( .A(n1983), .Y(mem_wdata_D[123]) );
  INVX12 U2329 ( .A(n1984), .Y(mem_wdata_D[126]) );
  BUFX12 U2330 ( .A(n12795), .Y(mem_addr_D[11]) );
  BUFX12 U2331 ( .A(n12794), .Y(mem_addr_D[14]) );
  INVX12 U2332 ( .A(n3712), .Y(mem_addr_D[21]) );
  INVX12 U2333 ( .A(n3810), .Y(mem_addr_D[24]) );
  INVX12 U2334 ( .A(n3831), .Y(mem_addr_D[25]) );
  INVX12 U2335 ( .A(n3832), .Y(mem_addr_D[26]) );
  CLKMX2X2 U2336 ( .A(\I_cache/cache[4][152] ), .B(n11152), .S0(n5276), .Y(
        n11567) );
  CLKMX2X2 U2337 ( .A(\D_cache/cache[0][83] ), .B(n11006), .S0(n4738), .Y(
        \D_cache/n1132 ) );
  CLKMX2X2 U2338 ( .A(\D_cache/cache[2][83] ), .B(n11006), .S0(n4808), .Y(
        \D_cache/n1130 ) );
  CLKMX2X2 U2339 ( .A(\I_cache/cache[1][99] ), .B(n11169), .S0(n5051), .Y(
        n11994) );
  OAI2BB2XL U2340 ( .B0(\i_MIPS/n234 ), .B1(net108200), .A0N(n4072), .A1N(
        n10829), .Y(\i_MIPS/N82 ) );
  AO22X1 U2341 ( .A0(n4072), .A1(net97452), .B0(net112406), .B1(
        \i_MIPS/IF_ID[97] ), .Y(\i_MIPS/N123 ) );
  AO22X1 U2342 ( .A0(n5545), .A1(n10550), .B0(net112406), .B1(net107812), .Y(
        \i_MIPS/N78 ) );
  AOI2BB2X2 U2343 ( .B0(\i_MIPS/IF_ID[87] ), .B1(net108670), .A0N(net108674), 
        .A1N(\i_MIPS/n205 ), .Y(n10554) );
  AO21X1 U2344 ( .A0(\i_MIPS/ID_EX[102] ), .A1(n202), .B0(n4380), .Y(
        \i_MIPS/n483 ) );
  AOI2BB2X2 U2345 ( .B0(net98496), .B1(n3897), .A0N(net98495), .A1N(net108660), 
        .Y(n4145) );
  MXI2X1 U2346 ( .A(n4540), .B(\i_MIPS/n229 ), .S0(n219), .Y(\i_MIPS/n498 ) );
  NAND3BX2 U2347 ( .AN(n10620), .B(n10618), .C(n10619), .Y(\i_MIPS/PC/n50 ) );
  MXI2X1 U2348 ( .A(\i_MIPS/n329 ), .B(\i_MIPS/n328 ), .S0(n205), .Y(
        \i_MIPS/n521 ) );
  NAND3X2 U2349 ( .A(n3932), .B(n10799), .C(n10798), .Y(\i_MIPS/PC/n64 ) );
  AOI32X1 U2350 ( .A0(net97444), .A1(n10855), .A2(n10797), .B0(
        \i_MIPS/IF_ID_30 ), .B1(net108682), .Y(n10798) );
  INVX1 U2351 ( .A(n11125), .Y(n11122) );
  OAI2BB2XL U2352 ( .B0(\i_MIPS/n225 ), .B1(net108198), .A0N(n5545), .A1N(
        n10394), .Y(\i_MIPS/N68 ) );
  OAI2BB2XL U2353 ( .B0(\i_MIPS/n222 ), .B1(net108198), .A0N(n4315), .A1N(
        n10236), .Y(\i_MIPS/N65 ) );
  OAI2BB2XL U2354 ( .B0(\i_MIPS/n160 ), .B1(net108198), .A0N(n4315), .A1N(
        n10207), .Y(\i_MIPS/N100 ) );
  CLKINVX1 U2355 ( .A(n10830), .Y(n10827) );
  CLKINVX1 U2356 ( .A(n10841), .Y(n10837) );
  CLKINVX1 U2357 ( .A(n10411), .Y(n10409) );
  OAI2BB2XL U2358 ( .B0(\i_MIPS/n168 ), .B1(net108194), .A0N(n4073), .A1N(
        n10438), .Y(\i_MIPS/N108 ) );
  NAND3BX2 U2359 ( .AN(n10821), .B(n10820), .C(n10819), .Y(\i_MIPS/PC/n44 ) );
  NAND3BX2 U2360 ( .AN(n10398), .B(n10397), .C(n10396), .Y(\i_MIPS/PC/n46 ) );
  NAND3BX1 U2361 ( .AN(n4452), .B(n9971), .C(n9970), .Y(\i_MIPS/n470 ) );
  CLKMX2X2 U2362 ( .A(\I_cache/cache[3][15] ), .B(n9643), .S0(n5135), .Y(
        n12664) );
  CLKMX2X2 U2363 ( .A(\I_cache/cache[7][152] ), .B(n11152), .S0(n5321), .Y(
        n11564) );
  CLKMX2X2 U2364 ( .A(\I_cache/cache[5][152] ), .B(n11152), .S0(n5233), .Y(
        n11566) );
  CLKMX2X2 U2365 ( .A(\I_cache/cache[3][152] ), .B(n11152), .S0(n5143), .Y(
        n11568) );
  CLKMX2X2 U2366 ( .A(\I_cache/cache[6][152] ), .B(n11152), .S0(n5359), .Y(
        n11565) );
  CLKMX2X2 U2367 ( .A(\I_cache/cache[1][152] ), .B(n11152), .S0(n5048), .Y(
        n11570) );
  CLKMX2X2 U2368 ( .A(\I_cache/cache[2][152] ), .B(n11152), .S0(n5189), .Y(
        n11569) );
  CLKMX2X2 U2369 ( .A(\I_cache/cache[0][152] ), .B(n11152), .S0(n5098), .Y(
        n11571) );
  CLKMX2X2 U2370 ( .A(\D_cache/cache[2][141] ), .B(n11035), .S0(n4808), .Y(
        \D_cache/n666 ) );
  CLKMX2X2 U2371 ( .A(\D_cache/cache[3][119] ), .B(n10948), .S0(n4854), .Y(
        \D_cache/n841 ) );
  CLKMX2X2 U2372 ( .A(\D_cache/cache[1][119] ), .B(n10948), .S0(n4784), .Y(
        \D_cache/n843 ) );
  CLKMX2X2 U2373 ( .A(\D_cache/cache[5][107] ), .B(n10715), .S0(n4942), .Y(
        \D_cache/n935 ) );
  CLKMX2X2 U2374 ( .A(\D_cache/cache[7][105] ), .B(n10703), .S0(n5004), .Y(
        \D_cache/n949 ) );
  CLKMX2X2 U2375 ( .A(\D_cache/cache[6][105] ), .B(n10703), .S0(n4960), .Y(
        \D_cache/n950 ) );
  CLKMX2X2 U2376 ( .A(\D_cache/cache[5][105] ), .B(n10703), .S0(n4941), .Y(
        \D_cache/n951 ) );
  CLKMX2X2 U2377 ( .A(\D_cache/cache[4][105] ), .B(n10703), .S0(n4896), .Y(
        \D_cache/n952 ) );
  CLKMX2X2 U2378 ( .A(\D_cache/cache[7][95] ), .B(n10879), .S0(n5002), .Y(
        \D_cache/n1029 ) );
  CLKMX2X2 U2379 ( .A(\D_cache/cache[6][95] ), .B(n10879), .S0(n4958), .Y(
        \D_cache/n1030 ) );
  CLKMX2X2 U2380 ( .A(\D_cache/cache[5][95] ), .B(n10879), .S0(n4938), .Y(
        \D_cache/n1031 ) );
  CLKMX2X2 U2381 ( .A(\D_cache/cache[4][95] ), .B(n10879), .S0(n4895), .Y(
        \D_cache/n1032 ) );
  CLKMX2X2 U2382 ( .A(\D_cache/cache[3][95] ), .B(n10879), .S0(n4848), .Y(
        \D_cache/n1033 ) );
  CLKMX2X2 U2383 ( .A(\D_cache/cache[2][95] ), .B(n10879), .S0(n4804), .Y(
        \D_cache/n1034 ) );
  CLKMX2X2 U2384 ( .A(\D_cache/cache[1][95] ), .B(n10879), .S0(n4781), .Y(
        \D_cache/n1035 ) );
  CLKMX2X2 U2385 ( .A(\D_cache/cache[5][94] ), .B(n3342), .S0(n4941), .Y(
        \D_cache/n1039 ) );
  CLKMX2X2 U2386 ( .A(\D_cache/cache[4][94] ), .B(n3342), .S0(n4894), .Y(
        \D_cache/n1040 ) );
  CLKMX2X2 U2387 ( .A(\D_cache/cache[1][94] ), .B(n3342), .S0(n4780), .Y(
        \D_cache/n1043 ) );
  CLKMX2X2 U2388 ( .A(\D_cache/cache[7][89] ), .B(n3337), .S0(n5000), .Y(
        \D_cache/n1077 ) );
  CLKMX2X2 U2389 ( .A(\D_cache/cache[6][89] ), .B(n3337), .S0(n4956), .Y(
        \D_cache/n1078 ) );
  CLKMX2X2 U2390 ( .A(\D_cache/cache[5][89] ), .B(n3337), .S0(n4936), .Y(
        \D_cache/n1079 ) );
  CLKMX2X2 U2391 ( .A(\D_cache/cache[4][89] ), .B(n3337), .S0(n4892), .Y(
        \D_cache/n1080 ) );
  CLKMX2X2 U2392 ( .A(\D_cache/cache[3][89] ), .B(n3337), .S0(n4846), .Y(
        \D_cache/n1081 ) );
  CLKMX2X2 U2393 ( .A(\D_cache/cache[2][89] ), .B(n3337), .S0(n4801), .Y(
        \D_cache/n1082 ) );
  CLKMX2X2 U2394 ( .A(\D_cache/cache[1][89] ), .B(n3337), .S0(n4778), .Y(
        \D_cache/n1083 ) );
  CLKMX2X2 U2395 ( .A(\D_cache/cache[7][88] ), .B(n3327), .S0(n5003), .Y(
        \D_cache/n1085 ) );
  CLKMX2X2 U2396 ( .A(\D_cache/cache[6][88] ), .B(n3327), .S0(n4959), .Y(
        \D_cache/n1086 ) );
  CLKMX2X2 U2397 ( .A(\D_cache/cache[5][88] ), .B(n3327), .S0(n4940), .Y(
        \D_cache/n1087 ) );
  CLKMX2X2 U2398 ( .A(\D_cache/cache[4][88] ), .B(n3327), .S0(n4895), .Y(
        \D_cache/n1088 ) );
  CLKMX2X2 U2399 ( .A(\D_cache/cache[3][88] ), .B(n3327), .S0(n4849), .Y(
        \D_cache/n1089 ) );
  CLKMX2X2 U2400 ( .A(\D_cache/cache[2][88] ), .B(n3327), .S0(n4805), .Y(
        \D_cache/n1090 ) );
  CLKMX2X2 U2401 ( .A(\D_cache/cache[1][88] ), .B(n3327), .S0(n4783), .Y(
        \D_cache/n1091 ) );
  CLKMX2X2 U2402 ( .A(\D_cache/cache[0][88] ), .B(n3327), .S0(n4736), .Y(
        \D_cache/n1092 ) );
  CLKMX2X2 U2403 ( .A(\D_cache/cache[5][85] ), .B(n3341), .S0(n4936), .Y(
        \D_cache/n1111 ) );
  CLKMX2X2 U2404 ( .A(\D_cache/cache[4][85] ), .B(n3341), .S0(n4893), .Y(
        \D_cache/n1112 ) );
  CLKMX2X2 U2405 ( .A(\D_cache/cache[3][85] ), .B(n3341), .S0(n4847), .Y(
        \D_cache/n1113 ) );
  CLKMX2X2 U2406 ( .A(\D_cache/cache[2][85] ), .B(n3341), .S0(n4802), .Y(
        \D_cache/n1114 ) );
  CLKMX2X2 U2407 ( .A(\D_cache/cache[1][85] ), .B(n3341), .S0(n4779), .Y(
        \D_cache/n1115 ) );
  CLKMX2X2 U2408 ( .A(\D_cache/cache[5][84] ), .B(n3340), .S0(n4942), .Y(
        \D_cache/n1119 ) );
  CLKMX2X2 U2409 ( .A(\D_cache/cache[4][84] ), .B(n3340), .S0(n4893), .Y(
        \D_cache/n1120 ) );
  CLKMX2X2 U2410 ( .A(\D_cache/cache[3][84] ), .B(n3340), .S0(n4847), .Y(
        \D_cache/n1121 ) );
  CLKMX2X2 U2411 ( .A(\D_cache/cache[2][84] ), .B(n3340), .S0(n4802), .Y(
        \D_cache/n1122 ) );
  CLKMX2X2 U2412 ( .A(\D_cache/cache[1][84] ), .B(n3340), .S0(n4779), .Y(
        \D_cache/n1123 ) );
  CLKMX2X2 U2413 ( .A(\D_cache/cache[5][83] ), .B(n11006), .S0(n4942), .Y(
        \D_cache/n1127 ) );
  CLKMX2X2 U2414 ( .A(\D_cache/cache[4][83] ), .B(n11006), .S0(n4898), .Y(
        \D_cache/n1128 ) );
  CLKMX2X2 U2415 ( .A(\D_cache/cache[1][83] ), .B(n11006), .S0(n4784), .Y(
        \D_cache/n1131 ) );
  CLKMX2X2 U2416 ( .A(\D_cache/cache[6][82] ), .B(n3339), .S0(n4957), .Y(
        \D_cache/n1134 ) );
  CLKMX2X2 U2417 ( .A(\D_cache/cache[5][82] ), .B(n3339), .S0(n4942), .Y(
        \D_cache/n1135 ) );
  CLKMX2X2 U2418 ( .A(\D_cache/cache[4][82] ), .B(n3339), .S0(n4893), .Y(
        \D_cache/n1136 ) );
  CLKMX2X2 U2419 ( .A(\D_cache/cache[3][82] ), .B(n3339), .S0(n4847), .Y(
        \D_cache/n1137 ) );
  CLKMX2X2 U2420 ( .A(\D_cache/cache[2][82] ), .B(n3339), .S0(n4802), .Y(
        \D_cache/n1138 ) );
  CLKMX2X2 U2421 ( .A(\D_cache/cache[1][82] ), .B(n3339), .S0(n4779), .Y(
        \D_cache/n1139 ) );
  CLKMX2X2 U2422 ( .A(\D_cache/cache[7][81] ), .B(n3331), .S0(n5003), .Y(
        \D_cache/n1141 ) );
  CLKMX2X2 U2423 ( .A(\D_cache/cache[6][81] ), .B(n3331), .S0(n4959), .Y(
        \D_cache/n1142 ) );
  CLKMX2X2 U2424 ( .A(\D_cache/cache[5][81] ), .B(n3331), .S0(n4938), .Y(
        \D_cache/n1143 ) );
  CLKMX2X2 U2425 ( .A(\D_cache/cache[4][81] ), .B(n3331), .S0(n4896), .Y(
        \D_cache/n1144 ) );
  CLKMX2X2 U2426 ( .A(\D_cache/cache[3][81] ), .B(n3331), .S0(n4849), .Y(
        \D_cache/n1145 ) );
  CLKMX2X2 U2427 ( .A(\D_cache/cache[2][81] ), .B(n3331), .S0(n4805), .Y(
        \D_cache/n1146 ) );
  CLKMX2X2 U2428 ( .A(\D_cache/cache[1][81] ), .B(n3331), .S0(n4781), .Y(
        \D_cache/n1147 ) );
  CLKMX2X2 U2429 ( .A(\D_cache/cache[0][81] ), .B(n3331), .S0(n4736), .Y(
        \D_cache/n1148 ) );
  CLKMX2X2 U2430 ( .A(\D_cache/cache[7][79] ), .B(n3330), .S0(n5004), .Y(
        \D_cache/n1157 ) );
  CLKMX2X2 U2431 ( .A(\D_cache/cache[6][79] ), .B(n3330), .S0(n4960), .Y(
        \D_cache/n1158 ) );
  CLKMX2X2 U2432 ( .A(\D_cache/cache[5][79] ), .B(n3330), .S0(n4942), .Y(
        \D_cache/n1159 ) );
  CLKMX2X2 U2433 ( .A(\D_cache/cache[4][79] ), .B(n3330), .S0(n4896), .Y(
        \D_cache/n1160 ) );
  CLKMX2X2 U2434 ( .A(\D_cache/cache[3][79] ), .B(n3330), .S0(n4850), .Y(
        \D_cache/n1161 ) );
  CLKMX2X2 U2435 ( .A(\D_cache/cache[2][79] ), .B(n3330), .S0(n4806), .Y(
        \D_cache/n1162 ) );
  CLKMX2X2 U2436 ( .A(\D_cache/cache[1][79] ), .B(n3330), .S0(n4784), .Y(
        \D_cache/n1163 ) );
  CLKMX2X2 U2437 ( .A(\D_cache/cache[0][79] ), .B(n3330), .S0(n4736), .Y(
        \D_cache/n1164 ) );
  CLKMX2X2 U2438 ( .A(\D_cache/cache[5][78] ), .B(n3350), .S0(n4941), .Y(
        \D_cache/n1167 ) );
  CLKMX2X2 U2439 ( .A(\D_cache/cache[1][78] ), .B(n3350), .S0(n4784), .Y(
        \D_cache/n1171 ) );
  CLKMX2X2 U2440 ( .A(\D_cache/cache[0][78] ), .B(n3350), .S0(n4739), .Y(
        \D_cache/n1172 ) );
  CLKMX2X2 U2441 ( .A(\D_cache/cache[5][77] ), .B(n3351), .S0(n4942), .Y(
        \D_cache/n1175 ) );
  CLKMX2X2 U2442 ( .A(\D_cache/cache[1][77] ), .B(n3351), .S0(n4784), .Y(
        \D_cache/n1179 ) );
  CLKMX2X2 U2443 ( .A(\D_cache/cache[0][77] ), .B(n3351), .S0(n4739), .Y(
        \D_cache/n1180 ) );
  CLKMX2X2 U2444 ( .A(\D_cache/cache[5][76] ), .B(n3352), .S0(n4942), .Y(
        \D_cache/n1183 ) );
  CLKMX2X2 U2445 ( .A(\D_cache/cache[1][76] ), .B(n3352), .S0(n4785), .Y(
        \D_cache/n1187 ) );
  CLKMX2X2 U2446 ( .A(\D_cache/cache[0][76] ), .B(n3352), .S0(n4739), .Y(
        \D_cache/n1188 ) );
  CLKMX2X2 U2447 ( .A(\D_cache/cache[7][75] ), .B(n3332), .S0(n5004), .Y(
        \D_cache/n1189 ) );
  CLKMX2X2 U2448 ( .A(\D_cache/cache[6][75] ), .B(n3332), .S0(n4960), .Y(
        \D_cache/n1190 ) );
  CLKMX2X2 U2449 ( .A(\D_cache/cache[5][75] ), .B(n3332), .S0(n4941), .Y(
        \D_cache/n1191 ) );
  CLKMX2X2 U2450 ( .A(\D_cache/cache[4][75] ), .B(n3332), .S0(n4896), .Y(
        \D_cache/n1192 ) );
  CLKMX2X2 U2451 ( .A(\D_cache/cache[3][75] ), .B(n3332), .S0(n4850), .Y(
        \D_cache/n1193 ) );
  CLKMX2X2 U2452 ( .A(\D_cache/cache[2][75] ), .B(n3332), .S0(n4806), .Y(
        \D_cache/n1194 ) );
  CLKMX2X2 U2453 ( .A(\D_cache/cache[1][75] ), .B(n3332), .S0(n4785), .Y(
        \D_cache/n1195 ) );
  CLKMX2X2 U2454 ( .A(\D_cache/cache[0][75] ), .B(n3332), .S0(n4738), .Y(
        \D_cache/n1196 ) );
  CLKMX2X2 U2455 ( .A(\D_cache/cache[7][70] ), .B(n3338), .S0(n5001), .Y(
        \D_cache/n1229 ) );
  CLKMX2X2 U2456 ( .A(\D_cache/cache[6][70] ), .B(n3338), .S0(n4959), .Y(
        \D_cache/n1230 ) );
  CLKMX2X2 U2457 ( .A(\D_cache/cache[5][70] ), .B(n3338), .S0(n4936), .Y(
        \D_cache/n1231 ) );
  CLKMX2X2 U2458 ( .A(\D_cache/cache[4][70] ), .B(n3338), .S0(n4894), .Y(
        \D_cache/n1232 ) );
  CLKMX2X2 U2459 ( .A(\D_cache/cache[3][70] ), .B(n3338), .S0(n4846), .Y(
        \D_cache/n1233 ) );
  CLKMX2X2 U2460 ( .A(\D_cache/cache[2][70] ), .B(n3338), .S0(n4803), .Y(
        \D_cache/n1234 ) );
  CLKMX2X2 U2461 ( .A(\D_cache/cache[1][70] ), .B(n3338), .S0(n4780), .Y(
        \D_cache/n1235 ) );
  CLKMX2X2 U2462 ( .A(\D_cache/cache[7][64] ), .B(n10964), .S0(n5009), .Y(
        \D_cache/n1277 ) );
  CLKMX2X2 U2463 ( .A(\D_cache/cache[6][64] ), .B(n10964), .S0(n4965), .Y(
        \D_cache/n1278 ) );
  CLKMX2X2 U2464 ( .A(\D_cache/cache[5][64] ), .B(n10964), .S0(n4944), .Y(
        \D_cache/n1279 ) );
  CLKMX2X2 U2465 ( .A(\D_cache/cache[7][61] ), .B(n10686), .S0(n5001), .Y(
        \D_cache/n1301 ) );
  CLKMX2X2 U2466 ( .A(\D_cache/cache[6][61] ), .B(n10686), .S0(n4957), .Y(
        \D_cache/n1302 ) );
  CLKMX2X2 U2467 ( .A(\D_cache/cache[5][44] ), .B(n10724), .S0(n4941), .Y(
        \D_cache/n1439 ) );
  CLKMX2X2 U2468 ( .A(\D_cache/cache[7][21] ), .B(n10669), .S0(n5001), .Y(
        \D_cache/n1621 ) );
  CLKMX2X2 U2469 ( .A(\D_cache/cache[6][21] ), .B(n10669), .S0(n4957), .Y(
        \D_cache/n1622 ) );
  CLKMX2X2 U2470 ( .A(\D_cache/cache[0][11] ), .B(n10709), .S0(n4738), .Y(
        \D_cache/n1708 ) );
  CLKMX2X2 U2471 ( .A(\I_cache/cache[2][26] ), .B(n9561), .S0(n5184), .Y(
        n12577) );
  CLKMX2X2 U2472 ( .A(n11061), .B(n3606), .S0(net112691), .Y(n11062) );
  MXI2X1 U2473 ( .A(\i_MIPS/PHT_2/n4 ), .B(\i_MIPS/PHT_2/n3 ), .S0(n4530), .Y(
        \i_MIPS/PHT_2/n50 ) );
  CLKMX2X2 U2474 ( .A(n406), .B(\i_MIPS/PHT_2/current_state_3[0] ), .S0(n11050), .Y(\i_MIPS/PHT_2/n44 ) );
  NAND2X1 U2475 ( .A(n11056), .B(n11053), .Y(\i_MIPS/PHT_2/n47 ) );
  CLKMX2X2 U2476 ( .A(\i_MIPS/PHT_2/n6 ), .B(n11052), .S0(n4461), .Y(n11053)
         );
  NAND3BX2 U2477 ( .AN(n11166), .B(n11165), .C(n11164), .Y(\i_MIPS/PC/n39 ) );
  OAI2BB2X1 U2478 ( .B0(\i_MIPS/n233 ), .B1(net108200), .A0N(n4073), .A1N(
        n10469), .Y(\i_MIPS/N81 ) );
  MXI2X1 U2479 ( .A(n406), .B(\i_MIPS/PHT_2/n2 ), .S0(net112691), .Y(n11049)
         );
  NAND2BX1 U2480 ( .AN(\i_MIPS/PHT_2/current_state_2[0] ), .B(net112691), .Y(
        n11052) );
  BUFX16 U2481 ( .A(net97574), .Y(net112691) );
  INVX1 U2482 ( .A(net101771), .Y(n4126) );
  CLKBUFX3 U2483 ( .A(n5179), .Y(n5160) );
  INVX12 U2484 ( .A(n4151), .Y(n9350) );
  INVX3 U2485 ( .A(net97995), .Y(net103250) );
  INVX16 U2486 ( .A(net102405), .Y(net101910) );
  INVX4 U2487 ( .A(net97834), .Y(net103090) );
  OA22X1 U2488 ( .A0(n4971), .A1(n1116), .B0(n5016), .B1(n2654), .Y(n8692) );
  OA22X1 U2489 ( .A0(n4974), .A1(n1129), .B0(n5019), .B1(n2663), .Y(n8199) );
  AND3X2 U2490 ( .A(net112306), .B(net101257), .C(net112420), .Y(n7477) );
  INVX4 U2491 ( .A(n10693), .Y(n8723) );
  NAND2X4 U2492 ( .A(n6572), .B(\i_MIPS/n352 ), .Y(n8553) );
  MX2X6 U2493 ( .A(\i_MIPS/n271 ), .B(n4496), .S0(n5622), .Y(n6572) );
  INVX3 U2494 ( .A(n8969), .Y(n9054) );
  NAND2X4 U2495 ( .A(n8862), .B(n7822), .Y(n8969) );
  INVX3 U2496 ( .A(n8940), .Y(n6521) );
  XOR3X1 U2497 ( .A(n10802), .B(n10801), .C(n10800), .Y(n10805) );
  BUFX4 U2498 ( .A(n4931), .Y(n4909) );
  OA22X1 U2499 ( .A0(n4827), .A1(n1148), .B0(n4872), .B1(n2706), .Y(n7431) );
  INVX4 U2500 ( .A(n11426), .Y(n10722) );
  CLKINVX1 U2501 ( .A(n7406), .Y(n254) );
  OAI31X1 U2502 ( .A0(n9044), .A1(n11182), .A2(n8172), .B0(n6596), .Y(n256) );
  AOI2BB1X4 U2503 ( .A0N(n11182), .A1N(n6595), .B0(n7482), .Y(n6596) );
  OA22X1 U2504 ( .A0(n4908), .A1(n1149), .B0(n4947), .B1(n2707), .Y(n9391) );
  NAND4X4 U2505 ( .A(n8107), .B(n8106), .C(n8105), .D(n8104), .Y(n11398) );
  INVX6 U2506 ( .A(n11398), .Y(n10297) );
  INVX3 U2507 ( .A(n8939), .Y(n8942) );
  NAND2X2 U2508 ( .A(n3414), .B(net98598), .Y(n4100) );
  INVX3 U2509 ( .A(net98728), .Y(net102791) );
  MX2X4 U2510 ( .A(n8347), .B(n8352), .S0(net107794), .Y(n7892) );
  OAI221X4 U2511 ( .A0(n4668), .A1(\i_MIPS/n347 ), .B0(net112334), .B1(
        \i_MIPS/n348 ), .C0(n7148), .Y(n8347) );
  XOR2X4 U2512 ( .A(n257), .B(n4135), .Y(n3933) );
  OA22XL U2513 ( .A0(n4816), .A1(n2144), .B0(n4862), .B1(n564), .Y(n8993) );
  OA22XL U2514 ( .A0(n4816), .A1(n709), .B0(n4862), .B1(n2277), .Y(n9082) );
  OA22XL U2515 ( .A0(n4816), .A1(n1257), .B0(n4862), .B1(n2799), .Y(n9078) );
  OA22XL U2516 ( .A0(n4843), .A1(n1111), .B0(n4862), .B1(n2700), .Y(n9509) );
  OA22XL U2517 ( .A0(n4816), .A1(n692), .B0(n4862), .B1(n2261), .Y(n8985) );
  OA22XL U2518 ( .A0(n4816), .A1(n1109), .B0(n4862), .B1(n2698), .Y(n8989) );
  OA22X1 U2519 ( .A0(n4816), .A1(n1140), .B0(n4862), .B1(n2702), .Y(n9086) );
  CLKINVX6 U2520 ( .A(n3929), .Y(n3798) );
  AO22X1 U2521 ( .A0(n4419), .A1(net137952), .B0(net112296), .B1(n8340), .Y(
        n8343) );
  AND3X6 U2522 ( .A(n6706), .B(n7481), .C(net111992), .Y(n6712) );
  MX2X4 U2523 ( .A(n7812), .B(n3844), .S0(net107796), .Y(n9163) );
  NAND2X6 U2524 ( .A(net98216), .B(net98217), .Y(n4094) );
  AO21X2 U2525 ( .A0(net98776), .A1(net98777), .B0(net111904), .Y(net98231) );
  INVX1 U2526 ( .A(n8339), .Y(n7505) );
  NAND3X4 U2527 ( .A(n4168), .B(n4169), .C(net112420), .Y(n8645) );
  INVX3 U2528 ( .A(n7504), .Y(n7508) );
  AOI22X4 U2529 ( .A0(net111960), .A1(n7836), .B0(net111968), .B1(net97995), 
        .Y(n3321) );
  NAND2X1 U2530 ( .A(n10691), .B(n4190), .Y(n4196) );
  AO22X1 U2531 ( .A0(net100583), .A1(n9492), .B0(n9458), .B1(net100585), .Y(
        n9473) );
  NAND2X8 U2532 ( .A(n4322), .B(n8943), .Y(n9065) );
  MX2XL U2533 ( .A(net112415), .B(net101082), .S0(n254), .Y(n7318) );
  MXI2X1 U2534 ( .A(\i_MIPS/n369 ), .B(net129005), .S0(n222), .Y(\i_MIPS/n560 ) );
  NAND2X4 U2535 ( .A(n6770), .B(n4536), .Y(n9162) );
  NOR4X4 U2536 ( .A(n8880), .B(n8879), .C(n8878), .D(n8877), .Y(net101556) );
  INVX1 U2537 ( .A(net105034), .Y(net102431) );
  BUFX2 U2538 ( .A(n4994), .Y(n4968) );
  BUFX16 U2539 ( .A(n4990), .Y(n4994) );
  OAI221X4 U2540 ( .A0(n3405), .A1(net100682), .B0(n8606), .B1(net101978), 
        .C0(n8605), .Y(n10636) );
  NAND2X6 U2541 ( .A(n10859), .B(n4457), .Y(n10880) );
  OAI2BB1X1 U2542 ( .A0N(n6842), .A1N(n3685), .B0(n6844), .Y(n6759) );
  OAI221X4 U2543 ( .A0(net112304), .A1(n6842), .B0(n6843), .B1(net101257), 
        .C0(net112420), .Y(n6847) );
  AO22X1 U2544 ( .A0(n6843), .A1(net137952), .B0(net112296), .B1(n6842), .Y(
        n6846) );
  NAND2X2 U2545 ( .A(n6962), .B(n8341), .Y(n6842) );
  NOR2X4 U2546 ( .A(n4170), .B(n7063), .Y(n7065) );
  CLKMX2X2 U2547 ( .A(net101082), .B(net112415), .S0(n8633), .Y(n7063) );
  OAI211X2 U2548 ( .A0(n9481), .A1(n9269), .B0(n9268), .C0(n9267), .Y(n9280)
         );
  INVX12 U2549 ( .A(n9145), .Y(n9481) );
  INVXL U2550 ( .A(n6640), .Y(n258) );
  NAND3BX2 U2551 ( .AN(n9056), .B(n3641), .C(n8953), .Y(n8977) );
  NOR3X2 U2552 ( .A(n4531), .B(n4532), .C(n4533), .Y(n6607) );
  NAND2BX2 U2553 ( .AN(n8241), .B(n8240), .Y(n8243) );
  NAND3X4 U2554 ( .A(n3814), .B(n7412), .C(n4433), .Y(n8240) );
  BUFX2 U2555 ( .A(n4930), .Y(n4913) );
  OA22X1 U2556 ( .A0(n4907), .A1(n1302), .B0(n4947), .B1(n2832), .Y(n9504) );
  NAND2X8 U2557 ( .A(n8862), .B(n4444), .Y(n9467) );
  NOR3X8 U2558 ( .A(n8946), .B(n2442), .C(n6515), .Y(n6525) );
  OAI211X2 U2559 ( .A0(n3412), .A1(net100682), .B0(n9400), .C0(n9399), .Y(
        n10319) );
  CLKMX2X2 U2560 ( .A(n7682), .B(n7681), .S0(net107812), .Y(net103581) );
  CLKBUFX6 U2561 ( .A(\i_MIPS/IR_ID[20] ), .Y(net107812) );
  BUFX4 U2562 ( .A(n9882), .Y(n259) );
  BUFX3 U2563 ( .A(n4767), .Y(n4758) );
  NAND4X2 U2564 ( .A(n9945), .B(n9944), .C(n9943), .D(n9942), .Y(n11220) );
  OA22X1 U2565 ( .A0(n5210), .A1(n1613), .B0(n5167), .B1(n3190), .Y(n9944) );
  OAI22XL U2566 ( .A0(n5114), .A1(n646), .B0(n5062), .B1(n2224), .Y(n4344) );
  OA22XL U2567 ( .A0(n5102), .A1(n1238), .B0(n5066), .B1(n2779), .Y(n6047) );
  OA22X2 U2568 ( .A0(n5102), .A1(n1409), .B0(n5074), .B1(n2940), .Y(n6051) );
  OAI21X4 U2569 ( .A0(n9044), .A1(n3776), .B0(n9042), .Y(n3698) );
  MX2XL U2570 ( .A(n3594), .B(n4601), .S0(n217), .Y(\i_MIPS/n403 ) );
  NAND2X4 U2571 ( .A(\i_MIPS/ALUin1[15] ), .B(n3666), .Y(n7798) );
  NAND3X6 U2572 ( .A(n3650), .B(n3651), .C(net103418), .Y(net98044) );
  XNOR2X2 U2573 ( .A(ICACHE_addr[29]), .B(n11344), .Y(n6092) );
  AND2X2 U2574 ( .A(n11120), .B(n10544), .Y(n4219) );
  NAND3X4 U2575 ( .A(n3680), .B(n3681), .C(n10544), .Y(n10444) );
  MX2XL U2576 ( .A(n3595), .B(n4621), .S0(n214), .Y(\i_MIPS/n401 ) );
  CLKAND2X2 U2577 ( .A(n10383), .B(n10228), .Y(n4390) );
  NAND3X4 U2578 ( .A(n7705), .B(n3429), .C(n4147), .Y(n7711) );
  CLKBUFX6 U2579 ( .A(n9987), .Y(n4885) );
  MX2XL U2580 ( .A(n4378), .B(n4614), .S0(n214), .Y(\i_MIPS/n407 ) );
  CLKBUFX3 U2581 ( .A(n4886), .Y(n4864) );
  NAND2X2 U2582 ( .A(net97496), .B(n10637), .Y(n10326) );
  BUFX8 U2583 ( .A(n4476), .Y(n4672) );
  AND2X2 U2584 ( .A(\i_MIPS/n312 ), .B(\i_MIPS/n314 ), .Y(n4448) );
  CLKBUFX2 U2585 ( .A(n9990), .Y(n4998) );
  CLKBUFX3 U2586 ( .A(n4998), .Y(n4997) );
  AO21XL U2587 ( .A0(n9266), .A1(n9265), .B0(n9264), .Y(n9267) );
  CLKINVX1 U2588 ( .A(n7536), .Y(n9266) );
  INVX4 U2589 ( .A(net112246), .Y(net112244) );
  INVX8 U2590 ( .A(net112248), .Y(net112240) );
  INVX6 U2591 ( .A(net112250), .Y(net112236) );
  INVX4 U2592 ( .A(net112246), .Y(net112242) );
  BUFX6 U2593 ( .A(n4425), .Y(n264) );
  AOI22X4 U2594 ( .A0(net111960), .A1(n9499), .B0(net111968), .B1(n10557), .Y(
        n3417) );
  BUFX4 U2595 ( .A(n4766), .Y(n4763) );
  BUFX12 U2596 ( .A(n3840), .Y(n5033) );
  CLKBUFX2 U2597 ( .A(n5312), .Y(n5309) );
  BUFX4 U2598 ( .A(n4840), .Y(n4818) );
  CLKBUFX4 U2599 ( .A(n4334), .Y(n5152) );
  CLKBUFX3 U2600 ( .A(n5216), .Y(n5211) );
  CLKBUFX2 U2601 ( .A(n5132), .Y(n5131) );
  BUFX8 U2602 ( .A(n4838), .Y(n4835) );
  CLKBUFX3 U2603 ( .A(n5312), .Y(n5310) );
  BUFX4 U2604 ( .A(n4884), .Y(n4883) );
  CLKBUFX3 U2605 ( .A(n5176), .Y(n5154) );
  CLKBUFX3 U2606 ( .A(n5525), .Y(n5518) );
  BUFX3 U2607 ( .A(n4931), .Y(n4910) );
  CLKBUFX2 U2608 ( .A(n5268), .Y(n5266) );
  CLKBUFX3 U2609 ( .A(n5261), .Y(n5259) );
  BUFX4 U2610 ( .A(n4774), .Y(n4769) );
  BUFX3 U2611 ( .A(n4774), .Y(n4771) );
  BUFX4 U2612 ( .A(n4954), .Y(n4953) );
  CLKBUFX3 U2613 ( .A(n5037), .Y(n5021) );
  CLKBUFX3 U2614 ( .A(n5037), .Y(n5023) );
  CLKBUFX3 U2615 ( .A(n4885), .Y(n4871) );
  CLKBUFX2 U2616 ( .A(n5179), .Y(n5178) );
  BUFX2 U2617 ( .A(n5085), .Y(n5060) );
  CLKBUFX4 U2618 ( .A(n5357), .Y(n5344) );
  CLKBUFX2 U2619 ( .A(net108160), .Y(net108150) );
  BUFX3 U2620 ( .A(n4891), .Y(n4934) );
  BUFX12 U2621 ( .A(n5261), .Y(n5240) );
  CLKBUFX3 U2622 ( .A(n5040), .Y(n5039) );
  CLKBUFX3 U2623 ( .A(n5032), .Y(n5016) );
  CLKBUFX8 U2624 ( .A(n4766), .Y(n4764) );
  BUFX16 U2625 ( .A(n4951), .Y(n4949) );
  BUFX8 U2626 ( .A(n4953), .Y(n4946) );
  CLKBUFX3 U2627 ( .A(n4884), .Y(n4875) );
  CLKBUFX3 U2628 ( .A(n4885), .Y(n4870) );
  BUFX4 U2629 ( .A(n9986), .Y(n4845) );
  BUFX4 U2630 ( .A(n4838), .Y(n4837) );
  BUFX16 U2631 ( .A(n4928), .Y(n4924) );
  BUFX4 U2632 ( .A(n4935), .Y(n4929) );
  BUFX20 U2633 ( .A(n4800), .Y(n4796) );
  BUFX4 U2634 ( .A(n5268), .Y(n5262) );
  BUFX4 U2635 ( .A(n5264), .Y(n5247) );
  BUFX4 U2636 ( .A(n5262), .Y(n5256) );
  BUFX4 U2637 ( .A(n4766), .Y(n4765) );
  CLKBUFX3 U2638 ( .A(n5032), .Y(n5018) );
  CLKBUFX3 U2639 ( .A(n3840), .Y(n5030) );
  BUFX4 U2640 ( .A(n4955), .Y(n4951) );
  INVX12 U2641 ( .A(n4248), .Y(n4249) );
  CLKBUFX3 U2642 ( .A(n4838), .Y(n4825) );
  CLKBUFX2 U2643 ( .A(n4890), .Y(n4889) );
  BUFX2 U2644 ( .A(n4886), .Y(n4862) );
  CLKBUFX3 U2645 ( .A(n5525), .Y(n5517) );
  CLKBUFX3 U2646 ( .A(n3840), .Y(n5029) );
  CLKBUFX3 U2647 ( .A(n5132), .Y(n5129) );
  CLKBUFX3 U2648 ( .A(n4994), .Y(n4970) );
  CLKBUFX2 U2649 ( .A(n4890), .Y(n4888) );
  BUFX2 U2650 ( .A(n4886), .Y(n4861) );
  BUFX4 U2651 ( .A(n4845), .Y(n4840) );
  BUFX4 U2652 ( .A(n4838), .Y(n4830) );
  BUFX4 U2653 ( .A(n5313), .Y(n5308) );
  BUFX4 U2654 ( .A(n5173), .Y(n5166) );
  CLKBUFX3 U2655 ( .A(n5032), .Y(n5019) );
  BUFX3 U2656 ( .A(n4891), .Y(n4932) );
  BUFX4 U2657 ( .A(n10193), .Y(n5223) );
  CLKBUFX3 U2658 ( .A(n4844), .Y(n4824) );
  BUFX4 U2659 ( .A(n5305), .Y(n5303) );
  CLKBUFX2 U2660 ( .A(n4890), .Y(n4887) );
  CLKBUFX3 U2661 ( .A(n4886), .Y(n4863) );
  CLKBUFX3 U2662 ( .A(n5520), .Y(n5519) );
  BUFX12 U2663 ( .A(n4797), .Y(n4788) );
  CLKBUFX3 U2664 ( .A(n5040), .Y(n5038) );
  CLKBUFX3 U2665 ( .A(n5032), .Y(n5014) );
  CLKBUFX3 U2666 ( .A(n3840), .Y(n5015) );
  CLKBUFX3 U2667 ( .A(n4991), .Y(n4981) );
  CLKBUFX3 U2668 ( .A(n4934), .Y(n4933) );
  BUFX4 U2669 ( .A(n5356), .Y(n5351) );
  CLKBUFX3 U2670 ( .A(n5356), .Y(n5352) );
  CLKBUFX2 U2671 ( .A(n5350), .Y(n5342) );
  BUFX4 U2672 ( .A(n5224), .Y(n5215) );
  CLKBUFX3 U2673 ( .A(n5215), .Y(n5213) );
  CLKBUFX8 U2674 ( .A(n10194), .Y(n5261) );
  CLKBUFX3 U2675 ( .A(n4840), .Y(n4817) );
  CLKBUFX3 U2676 ( .A(n4884), .Y(n4874) );
  BUFX8 U2677 ( .A(n5530), .Y(n5540) );
  CLKBUFX3 U2678 ( .A(n5036), .Y(n5020) );
  BUFX8 U2679 ( .A(n4333), .Y(n4800) );
  BUFX2 U2680 ( .A(n5261), .Y(n5239) );
  BUFX16 U2681 ( .A(n9990), .Y(n4990) );
  BUFX4 U2682 ( .A(n9990), .Y(n4993) );
  BUFX8 U2683 ( .A(n4990), .Y(n4989) );
  CLKBUFX2 U2684 ( .A(n5132), .Y(n5130) );
  CLKBUFX3 U2685 ( .A(n5180), .Y(n5170) );
  CLKBUFX3 U2686 ( .A(n5312), .Y(n5311) );
  CLKBUFX3 U2687 ( .A(n5306), .Y(n5298) );
  CLKBUFX3 U2688 ( .A(n4838), .Y(n4827) );
  BUFX16 U2689 ( .A(n9989), .Y(n4950) );
  BUFX4 U2690 ( .A(n4928), .Y(n4925) );
  BUFX4 U2691 ( .A(n4930), .Y(n4912) );
  CLKBUFX4 U2692 ( .A(n5133), .Y(n5127) );
  BUFX4 U2693 ( .A(n9990), .Y(n4991) );
  BUFX12 U2694 ( .A(n4796), .Y(n4790) );
  BUFX6 U2695 ( .A(n9529), .Y(n4713) );
  BUFX4 U2696 ( .A(n9529), .Y(n4711) );
  BUFX6 U2697 ( .A(n9529), .Y(n4712) );
  CLKBUFX3 U2698 ( .A(n3840), .Y(n5025) );
  BUFX4 U2699 ( .A(n4767), .Y(n4761) );
  BUFX4 U2700 ( .A(n4928), .Y(n4927) );
  CLKBUFX3 U2701 ( .A(n5261), .Y(n5260) );
  CLKBUFX3 U2702 ( .A(n4993), .Y(n4973) );
  BUFX8 U2703 ( .A(n4798), .Y(n4791) );
  CLKBUFX4 U2704 ( .A(n5357), .Y(n5349) );
  BUFX4 U2705 ( .A(n5349), .Y(n5348) );
  BUFX4 U2706 ( .A(n5216), .Y(n5210) );
  CLKBUFX3 U2707 ( .A(n5223), .Y(n5220) );
  CLKBUFX3 U2708 ( .A(n5215), .Y(n5212) );
  CLKBUFX2 U2709 ( .A(n4955), .Y(n4952) );
  CLKBUFX8 U2710 ( .A(n4955), .Y(n4948) );
  AND2X1 U2711 ( .A(n10287), .B(n10286), .Y(n2211) );
  AND2X1 U2712 ( .A(n10559), .B(n10558), .Y(n1978) );
  AND2X2 U2713 ( .A(n4521), .B(n4446), .Y(net128160) );
  INVX6 U2714 ( .A(net112196), .Y(net112182) );
  BUFX4 U2715 ( .A(net108200), .Y(net108192) );
  BUFX4 U2716 ( .A(net133468), .Y(net112090) );
  BUFX4 U2717 ( .A(net133470), .Y(net112142) );
  CLKINVX3 U2718 ( .A(n4439), .Y(n5463) );
  CLKINVX3 U2719 ( .A(n4439), .Y(n5462) );
  AND2X2 U2720 ( .A(net98385), .B(net98386), .Y(n1996) );
  INVX4 U2721 ( .A(n4485), .Y(n10194) );
  CLKBUFX3 U2722 ( .A(n4998), .Y(n4995) );
  CLKBUFX3 U2723 ( .A(n4994), .Y(n4971) );
  BUFX4 U2724 ( .A(n3840), .Y(n5027) );
  CLKBUFX3 U2725 ( .A(n3840), .Y(n5031) );
  BUFX8 U2726 ( .A(n4334), .Y(n5179) );
  BUFX4 U2727 ( .A(n4335), .Y(n5357) );
  BUFX8 U2728 ( .A(n5313), .Y(n5307) );
  BUFX4 U2729 ( .A(n5307), .Y(n5295) );
  AND2X2 U2730 ( .A(\i_MIPS/PHT_2/history_state[1] ), .B(\i_MIPS/PHT_2/n13 ), 
        .Y(n270) );
  INVX4 U2731 ( .A(net112228), .Y(net112224) );
  BUFX4 U2732 ( .A(n9535), .Y(n4729) );
  BUFX4 U2733 ( .A(net112046), .Y(net112036) );
  BUFX4 U2734 ( .A(net133468), .Y(net112098) );
  INVX4 U2735 ( .A(n4477), .Y(n4698) );
  BUFX12 U2736 ( .A(net112300), .Y(net112304) );
  CLKAND2X8 U2737 ( .A(n10789), .B(n10788), .Y(n4439) );
  BUFX6 U2738 ( .A(n4724), .Y(n4726) );
  BUFX4 U2739 ( .A(n5532), .Y(n5531) );
  AND2XL U2740 ( .A(net98780), .B(net98781), .Y(n301) );
  AND2XL U2741 ( .A(n10526), .B(n10525), .Y(n302) );
  BUFX4 U2742 ( .A(n4774), .Y(n4770) );
  BUFX4 U2743 ( .A(n5041), .Y(n5037) );
  BUFX4 U2744 ( .A(n5262), .Y(n5255) );
  CLKBUFX3 U2745 ( .A(n5261), .Y(n5258) );
  CLKBUFX4 U2746 ( .A(n4935), .Y(n4931) );
  BUFX2 U2747 ( .A(n4928), .Y(n4915) );
  BUFX4 U2748 ( .A(n5134), .Y(n5126) );
  AND2X4 U2749 ( .A(n4661), .B(n3783), .Y(n4469) );
  CLKBUFX8 U2750 ( .A(n4884), .Y(n4873) );
  CLKBUFX4 U2751 ( .A(n4845), .Y(n4839) );
  INVX4 U2752 ( .A(n11511), .Y(n4652) );
  INVX6 U2753 ( .A(n4482), .Y(n4700) );
  AND2XL U2754 ( .A(n10563), .B(n10562), .Y(n1985) );
  AND2XL U2755 ( .A(n10565), .B(n10564), .Y(n1980) );
  AND2XL U2756 ( .A(n10561), .B(n10560), .Y(n1991) );
  AND2XL U2757 ( .A(n10322), .B(n10321), .Y(n1995) );
  AND2XL U2758 ( .A(n10489), .B(n10488), .Y(n1999) );
  AND2XL U2759 ( .A(net98340), .B(net98341), .Y(n1988) );
  AND2XL U2760 ( .A(net98776), .B(net98777), .Y(n1989) );
  AND2XL U2761 ( .A(net98758), .B(net98759), .Y(n1990) );
  AND2XL U2762 ( .A(net98335), .B(net98336), .Y(n1992) );
  AND2XL U2763 ( .A(net99164), .B(net99165), .Y(n1986) );
  AND2XL U2764 ( .A(n9978), .B(n9977), .Y(n2000) );
  AND2XL U2765 ( .A(net99002), .B(net99003), .Y(n1979) );
  AND2XL U2766 ( .A(net98366), .B(net98367), .Y(n1994) );
  CLKBUFX3 U2767 ( .A(n10639), .Y(n5425) );
  AND3X2 U2768 ( .A(net97452), .B(\i_MIPS/IF_ID[97] ), .C(\i_MIPS/n236 ), .Y(
        n324) );
  AND2X4 U2769 ( .A(n9242), .B(n9456), .Y(n325) );
  BUFX4 U2770 ( .A(net112046), .Y(net112038) );
  CLKBUFX3 U2771 ( .A(net112034), .Y(net112030) );
  BUFX4 U2772 ( .A(net112034), .Y(net112020) );
  BUFX8 U2773 ( .A(n4706), .Y(n4708) );
  BUFX6 U2774 ( .A(n4706), .Y(n4709) );
  BUFX4 U2775 ( .A(n4706), .Y(n4707) );
  BUFX4 U2776 ( .A(n4349), .Y(n4688) );
  CLKBUFX4 U2777 ( .A(n4349), .Y(n4687) );
  MXI2X2 U2778 ( .A(n10891), .B(n10890), .S0(n5520), .Y(n10892) );
  BUFX4 U2779 ( .A(net112084), .Y(net112072) );
  INVX1 U2780 ( .A(net100682), .Y(net100537) );
  BUFX12 U2781 ( .A(net97418), .Y(net108200) );
  BUFX4 U2782 ( .A(n9533), .Y(n4721) );
  BUFX8 U2783 ( .A(n4714), .Y(n4716) );
  BUFX12 U2784 ( .A(net101413), .Y(net112300) );
  CLKINVX3 U2785 ( .A(n9411), .Y(n9534) );
  BUFX4 U2786 ( .A(n4768), .Y(n4754) );
  BUFX6 U2787 ( .A(n9990), .Y(n4992) );
  CLKINVX3 U2788 ( .A(n4945), .Y(n4943) );
  CLKINVX3 U2789 ( .A(n4791), .Y(n4780) );
  BUFX4 U2790 ( .A(n5224), .Y(n5216) );
  OR2X1 U2791 ( .A(n3677), .B(n10511), .Y(n407) );
  NAND2X1 U2792 ( .A(DCACHE_addr[4]), .B(n11481), .Y(n408) );
  XNOR2X2 U2793 ( .A(n10234), .B(ICACHE_addr[10]), .Y(n409) );
  CLKINVX1 U2794 ( .A(n10317), .Y(n5409) );
  AND2XL U2795 ( .A(n7798), .B(n7527), .Y(n413) );
  AND2X2 U2796 ( .A(n11130), .B(n6121), .Y(n414) );
  BUFX4 U2797 ( .A(n9524), .Y(n4680) );
  BUFX16 U2798 ( .A(n12954), .Y(DCACHE_addr[1]) );
  INVX6 U2799 ( .A(net112160), .Y(net112152) );
  INVX4 U2800 ( .A(net128158), .Y(net112170) );
  CLKBUFX6 U2801 ( .A(net100537), .Y(net111966) );
  XNOR3X1 U2802 ( .A(n10603), .B(n10602), .C(n10601), .Y(n637) );
  INVX12 U2803 ( .A(n11480), .Y(n11511) );
  INVX6 U2804 ( .A(n4652), .Y(n4653) );
  INVX4 U2805 ( .A(n4652), .Y(n4654) );
  BUFX4 U2806 ( .A(n9527), .Y(n4690) );
  CLKBUFX8 U2807 ( .A(n4689), .Y(n4692) );
  CLKBUFX6 U2808 ( .A(n4689), .Y(n4691) );
  CLKBUFX8 U2809 ( .A(n3428), .Y(n5428) );
  NAND2XL U2810 ( .A(ICACHE_addr[1]), .B(n10176), .Y(n10639) );
  BUFX4 U2811 ( .A(net100599), .Y(net112034) );
  NAND2X2 U2812 ( .A(n6458), .B(n4446), .Y(net133496) );
  BUFX4 U2813 ( .A(net133496), .Y(net112084) );
  CLKINVX1 U2814 ( .A(n11346), .Y(n11003) );
  BUFX8 U2815 ( .A(n5503), .Y(n5505) );
  BUFX8 U2816 ( .A(n5503), .Y(n5504) );
  BUFX4 U2817 ( .A(net107808), .Y(net107804) );
  INVX4 U2818 ( .A(net128154), .Y(net112222) );
  INVX6 U2819 ( .A(net128160), .Y(net112188) );
  BUFX3 U2820 ( .A(n9534), .Y(n4724) );
  BUFX12 U2821 ( .A(n4725), .Y(n4727) );
  BUFX4 U2822 ( .A(n4714), .Y(n4717) );
  BUFX16 U2823 ( .A(n12951), .Y(DCACHE_addr[6]) );
  CLKBUFX3 U2824 ( .A(n11039), .Y(n5527) );
  BUFX12 U2825 ( .A(net133469), .Y(net112112) );
  BUFX20 U2826 ( .A(net128151), .Y(net112338) );
  INVX16 U2827 ( .A(net101257), .Y(net137952) );
  CLKINVX3 U2828 ( .A(n4742), .Y(n4739) );
  CLKINVX3 U2829 ( .A(n4948), .Y(n4936) );
  CLKINVX3 U2830 ( .A(n4948), .Y(n4937) );
  CLKINVX3 U2831 ( .A(n4788), .Y(n4784) );
  CLKINVX3 U2832 ( .A(n4788), .Y(n4785) );
  CLKINVX3 U2833 ( .A(n4913), .Y(n4900) );
  CLKINVX3 U2834 ( .A(n4904), .Y(n4898) );
  CLKBUFX2 U2835 ( .A(n5310), .Y(n5283) );
  CLKINVX3 U2836 ( .A(n5058), .Y(n5048) );
  NAND2X1 U2837 ( .A(n4653), .B(n11350), .Y(n1939) );
  NAND2X1 U2838 ( .A(n4653), .B(n11352), .Y(n1940) );
  NAND2X1 U2839 ( .A(n4653), .B(n11356), .Y(n1941) );
  NAND2X1 U2840 ( .A(n4653), .B(n11367), .Y(n1942) );
  NAND2X1 U2841 ( .A(n4653), .B(n11372), .Y(n1943) );
  NAND2X1 U2842 ( .A(n4653), .B(n11376), .Y(n1944) );
  NAND2X1 U2843 ( .A(n4654), .B(n11399), .Y(n1945) );
  NAND2X1 U2844 ( .A(n4654), .B(n11404), .Y(n1946) );
  NAND2X1 U2845 ( .A(n4653), .B(n11430), .Y(n1947) );
  AOI22X1 U2846 ( .A0(n12952), .A1(n11510), .B0(n4653), .B1(n11483), .Y(n1948)
         );
  AOI22X1 U2847 ( .A0(DCACHE_addr[8]), .A1(n11510), .B0(n4653), .B1(n11486), 
        .Y(n1949) );
  AOI22X1 U2848 ( .A0(n12947), .A1(n11510), .B0(n4654), .B1(n11488), .Y(n1950)
         );
  AOI22X1 U2849 ( .A0(n12941), .A1(n11510), .B0(n3737), .B1(n11494), .Y(n1951)
         );
  AOI22X1 U2850 ( .A0(n12940), .A1(n11510), .B0(n5551), .B1(n11495), .Y(n1952)
         );
  NAND2X1 U2851 ( .A(n5551), .B(n11382), .Y(n1953) );
  NAND2X1 U2852 ( .A(n5551), .B(n11384), .Y(n1954) );
  NAND2X1 U2853 ( .A(n5551), .B(n11388), .Y(n1955) );
  NAND2X1 U2854 ( .A(n5551), .B(n11393), .Y(n1956) );
  NAND2X1 U2855 ( .A(n5551), .B(n11394), .Y(n1957) );
  NAND2X1 U2856 ( .A(n4653), .B(n11441), .Y(n1958) );
  NAND2X1 U2857 ( .A(n4653), .B(n11444), .Y(n1959) );
  NAND2X1 U2858 ( .A(n4653), .B(n11447), .Y(n1960) );
  NAND2X1 U2859 ( .A(n4654), .B(n11450), .Y(n1961) );
  NAND2X1 U2860 ( .A(n4653), .B(n11454), .Y(n1962) );
  NAND2X1 U2861 ( .A(n4653), .B(n11462), .Y(n1963) );
  NAND2X1 U2862 ( .A(n4653), .B(n11466), .Y(n1964) );
  NAND2X1 U2863 ( .A(n4653), .B(n11468), .Y(n1965) );
  NAND2X1 U2864 ( .A(n4653), .B(n11469), .Y(n1966) );
  NAND2X1 U2865 ( .A(n4654), .B(n11471), .Y(n1967) );
  NAND2X1 U2866 ( .A(n4653), .B(n11474), .Y(n1968) );
  NAND2X1 U2867 ( .A(n4653), .B(n11477), .Y(n1969) );
  AOI22X2 U2868 ( .A0(ICACHE_addr[5]), .A1(n11512), .B0(n4656), .B1(n11320), 
        .Y(n1970) );
  AOI22X2 U2869 ( .A0(ICACHE_addr[7]), .A1(n11512), .B0(n4657), .B1(n11322), 
        .Y(n1971) );
  AOI22X2 U2870 ( .A0(ICACHE_addr[8]), .A1(n11512), .B0(n4656), .B1(n11323), 
        .Y(n1972) );
  AOI22X2 U2871 ( .A0(ICACHE_addr[10]), .A1(n11512), .B0(n4657), .B1(n11325), 
        .Y(n1973) );
  AOI22X2 U2872 ( .A0(ICACHE_addr[11]), .A1(n11512), .B0(n4656), .B1(n11326), 
        .Y(n1974) );
  BUFX12 U2873 ( .A(n5554), .Y(n5556) );
  INVX12 U2874 ( .A(n4655), .Y(n4657) );
  INVX12 U2875 ( .A(n4655), .Y(n4656) );
  NAND2X1 U2876 ( .A(n4654), .B(n11455), .Y(n1975) );
  NAND2X1 U2877 ( .A(n4654), .B(n11458), .Y(n1976) );
  NAND2X1 U2878 ( .A(n4654), .B(n11461), .Y(n1981) );
  NAND2X1 U2879 ( .A(n4654), .B(n11470), .Y(n1982) );
  NAND2X1 U2880 ( .A(n4654), .B(n11473), .Y(n1983) );
  NAND2X1 U2881 ( .A(n4654), .B(n11476), .Y(n1984) );
  AND2X2 U2882 ( .A(n10568), .B(n4608), .Y(n1993) );
  AND2X2 U2883 ( .A(net98390), .B(net98391), .Y(n1997) );
  AND2X2 U2884 ( .A(n10137), .B(n10136), .Y(n1998) );
  INVX6 U2885 ( .A(n11482), .Y(n11510) );
  XNOR3X1 U2886 ( .A(n11161), .B(n4387), .C(n11173), .Y(n2016) );
  BUFX16 U2887 ( .A(n12950), .Y(DCACHE_addr[7]) );
  CLKINVX1 U2888 ( .A(net137891), .Y(n3718) );
  AND2X2 U2889 ( .A(n8955), .B(n8970), .Y(n2209) );
  AND3X2 U2890 ( .A(n10187), .B(n10189), .C(n10190), .Y(n2212) );
  AND2X4 U2891 ( .A(n4521), .B(n4503), .Y(net128159) );
  BUFX4 U2892 ( .A(net128158), .Y(net112176) );
  OR2X1 U2893 ( .A(n9140), .B(n9142), .Y(n2442) );
  BUFX4 U2894 ( .A(n4440), .Y(n4705) );
  XNOR3X1 U2895 ( .A(net112400), .B(n10465), .C(n10822), .Y(n2649) );
  BUFX16 U2896 ( .A(n12955), .Y(net112962) );
  CLKBUFX3 U2897 ( .A(net128155), .Y(net112248) );
  BUFX16 U2898 ( .A(net128830), .Y(net111628) );
  INVX16 U2899 ( .A(net111628), .Y(net111624) );
  MXI2X2 U2900 ( .A(n10219), .B(n10218), .S0(n5515), .Y(n10220) );
  MXI2X2 U2901 ( .A(n10267), .B(n10266), .S0(n5515), .Y(n10268) );
  BUFX8 U2902 ( .A(n4383), .Y(n5494) );
  NAND2X2 U2903 ( .A(n6458), .B(n4504), .Y(net133468) );
  AOI22X2 U2904 ( .A0(net111966), .A1(n10965), .B0(net111962), .B1(n8387), .Y(
        n3324) );
  BUFX4 U2905 ( .A(n9525), .Y(n4681) );
  BUFX8 U2906 ( .A(n4681), .Y(n4684) );
  BUFX8 U2907 ( .A(n4681), .Y(n4683) );
  BUFX16 U2908 ( .A(\i_MIPS/ID_EX[82] ), .Y(n4662) );
  INVX6 U2909 ( .A(net112420), .Y(net100583) );
  AND3X2 U2910 ( .A(n6044), .B(n6047), .C(n6046), .Y(n3326) );
  NAND2X1 U2911 ( .A(n4524), .B(n11009), .Y(n11039) );
  AND2X2 U2912 ( .A(n4500), .B(n4448), .Y(n4477) );
  AND2X8 U2913 ( .A(n3745), .B(n10072), .Y(n4385) );
  AND2X4 U2914 ( .A(n4238), .B(n4239), .Y(n3339) );
  AND2X4 U2915 ( .A(n4202), .B(n4203), .Y(n3340) );
  AND2X4 U2916 ( .A(n4240), .B(n4241), .Y(n3350) );
  AND2X2 U2917 ( .A(n4210), .B(n4211), .Y(n3351) );
  AND2X2 U2918 ( .A(n4212), .B(n4213), .Y(n3352) );
  AND3X8 U2919 ( .A(n3678), .B(n3679), .C(n10451), .Y(n3357) );
  AND3X4 U2920 ( .A(n4155), .B(n4156), .C(n6338), .Y(n3359) );
  CLKBUFX3 U2921 ( .A(net133470), .Y(net112138) );
  BUFX4 U2922 ( .A(net112084), .Y(net112078) );
  AND4X8 U2923 ( .A(n4392), .B(\i_MIPS/EX_MEM_1 ), .C(DCACHE_ren), .D(n9), .Y(
        n3400) );
  CLKBUFX3 U2924 ( .A(net108156), .Y(net108128) );
  BUFX4 U2925 ( .A(n9535), .Y(n4728) );
  BUFX12 U2926 ( .A(n9534), .Y(n4725) );
  BUFX16 U2927 ( .A(n12945), .Y(DCACHE_addr[12]) );
  NAND2X6 U2928 ( .A(n4618), .B(n6500), .Y(n7046) );
  AND2X4 U2929 ( .A(n6353), .B(n6355), .Y(n3410) );
  AO21X2 U2930 ( .A0(net98366), .A1(net98367), .B0(net111904), .Y(net98364) );
  BUFX16 U2931 ( .A(n12929), .Y(DCACHE_addr[28]) );
  CLKBUFX3 U2932 ( .A(n10640), .Y(n5429) );
  BUFX12 U2933 ( .A(n10990), .Y(n5495) );
  BUFX8 U2934 ( .A(n10990), .Y(n5496) );
  AND2X4 U2935 ( .A(n7221), .B(n7045), .Y(n3413) );
  INVX1 U2936 ( .A(net102049), .Y(net100597) );
  CLKBUFX3 U2937 ( .A(net100597), .Y(net112014) );
  CLKMX2X4 U2938 ( .A(\i_MIPS/n275 ), .B(n4495), .S0(n5622), .Y(n6573) );
  AOI22X2 U2939 ( .A0(net97817), .A1(net111968), .B0(net111962), .B1(n7088), 
        .Y(n3414) );
  BUFX16 U2940 ( .A(n3927), .Y(net108708) );
  AOI22X4 U2941 ( .A0(net111960), .A1(n8187), .B0(net111968), .B1(n3830), .Y(
        n3416) );
  INVX3 U2942 ( .A(net112406), .Y(net97418) );
  AOI22X4 U2943 ( .A0(net111966), .A1(n10502), .B0(net111962), .B1(n8785), .Y(
        n3419) );
  AOI22X4 U2944 ( .A0(net111966), .A1(net97783), .B0(net111964), .B1(n4104), 
        .Y(n3420) );
  AOI22X4 U2945 ( .A0(net111968), .A1(net97770), .B0(net111964), .B1(n6879), 
        .Y(n3421) );
  AOI22X4 U2946 ( .A0(net111966), .A1(n10693), .B0(net111960), .B1(n8683), .Y(
        n3422) );
  AOI22X4 U2947 ( .A0(n10774), .A1(net111966), .B0(net111962), .B1(n8296), .Y(
        n3423) );
  NAND4X4 U2948 ( .A(\i_MIPS/EX_MEM_1 ), .B(DCACHE_ren), .C(n10071), .D(n11345), .Y(n3424) );
  BUFX4 U2949 ( .A(net128156), .Y(net112266) );
  BUFX4 U2950 ( .A(net101413), .Y(net112306) );
  INVX3 U2951 ( .A(n4652), .Y(n3737) );
  AND2X4 U2952 ( .A(n402), .B(n4503), .Y(net128154) );
  BUFX8 U2953 ( .A(net137952), .Y(net111994) );
  CLKBUFX3 U2954 ( .A(net111996), .Y(net111992) );
  AOI22X4 U2955 ( .A0(net111968), .A1(net98393), .B0(net111962), .B1(n7343), 
        .Y(n3425) );
  AOI22X4 U2956 ( .A0(net111968), .A1(net97684), .B0(net111962), .B1(n7004), 
        .Y(n3426) );
  OR3X4 U2957 ( .A(n7402), .B(n7403), .C(n7401), .Y(n3427) );
  CLKINVX16 U2958 ( .A(n5626), .Y(n5622) );
  CLKINVX1 U2959 ( .A(n9163), .Y(n7706) );
  CLKMX2X2 U2960 ( .A(\D_cache/cache[2][130] ), .B(n3834), .S0(n4808), .Y(
        \D_cache/n754 ) );
  NAND2X2 U2961 ( .A(n9487), .B(n9476), .Y(n8945) );
  INVX12 U2962 ( .A(net133471), .Y(net100585) );
  NAND2X4 U2963 ( .A(n6458), .B(n4503), .Y(net133469) );
  INVX3 U2964 ( .A(n6978), .Y(n9468) );
  INVX3 U2965 ( .A(\i_MIPS/ID_EX[81] ), .Y(net107808) );
  INVX4 U2966 ( .A(net111960), .Y(n3787) );
  BUFX16 U2967 ( .A(net100535), .Y(net111962) );
  AND3X8 U2968 ( .A(n3691), .B(n3692), .C(n8225), .Y(n3430) );
  BUFX2 U2969 ( .A(n4954), .Y(n4945) );
  AND2X2 U2970 ( .A(n11346), .B(mem_ready_D), .Y(n3431) );
  INVX3 U2971 ( .A(net97783), .Y(net104888) );
  AND4X6 U2972 ( .A(n8186), .B(n8185), .C(n8184), .D(n8183), .Y(n3714) );
  NAND4X2 U2973 ( .A(n6412), .B(n6411), .C(n6410), .D(n6409), .Y(n11498) );
  AND2X2 U2974 ( .A(\i_MIPS/IF_ID[64] ), .B(\i_MIPS/IF_ID[97] ), .Y(n3432) );
  INVX3 U2975 ( .A(n10601), .Y(n10605) );
  NAND4X6 U2976 ( .A(n9760), .B(n9759), .C(n9758), .D(n9757), .Y(n10601) );
  INVX16 U2977 ( .A(n4593), .Y(DCACHE_addr[18]) );
  INVX12 U2978 ( .A(n4666), .Y(n6298) );
  CLKINVX1 U2979 ( .A(mem_ready_D), .Y(n3854) );
  NAND2X1 U2980 ( .A(n8532), .B(n9268), .Y(n8560) );
  CLKAND2X12 U2981 ( .A(n4656), .B(n11293), .Y(mem_wdata_I[107]) );
  CLKAND2X12 U2982 ( .A(n4661), .B(n11318), .Y(mem_addr_I[5]) );
  CLKAND2X12 U2983 ( .A(n3785), .B(n11318), .Y(mem_addr_I[6]) );
  CLKAND2X12 U2984 ( .A(n4656), .B(n11236), .Y(mem_wdata_I[50]) );
  CLKAND2X12 U2985 ( .A(n4656), .B(n11287), .Y(mem_wdata_I[101]) );
  CLKAND2X12 U2986 ( .A(n4654), .B(n11419), .Y(mem_wdata_D[69]) );
  CLKAND2X12 U2987 ( .A(n4654), .B(n11434), .Y(mem_wdata_D[84]) );
  CLKAND2X12 U2988 ( .A(n4654), .B(n11407), .Y(mem_wdata_D[57]) );
  CLKAND2X12 U2989 ( .A(n4654), .B(n11401), .Y(mem_wdata_D[51]) );
  INVX12 U2990 ( .A(n3708), .Y(mem_addr_D[20]) );
  INVX12 U2991 ( .A(n3811), .Y(mem_addr_D[13]) );
  CLKAND2X12 U2992 ( .A(n4653), .B(n11400), .Y(mem_wdata_D[50]) );
  CLKAND2X12 U2993 ( .A(n4653), .B(n11403), .Y(mem_wdata_D[53]) );
  BUFX12 U2994 ( .A(n4665), .Y(DCACHE_addr[3]) );
  CLKAND2X12 U2995 ( .A(n4653), .B(n11374), .Y(mem_wdata_D[24]) );
  INVX12 U2996 ( .A(n1942), .Y(mem_wdata_D[17]) );
  INVX12 U2997 ( .A(n1939), .Y(mem_wdata_D[0]) );
  NAND2X1 U2998 ( .A(n3677), .B(n3803), .Y(n11481) );
  INVX1 U2999 ( .A(n11510), .Y(n3803) );
  CLKINVX1 U3000 ( .A(n11096), .Y(n11094) );
  XOR2X1 U3001 ( .A(n10066), .B(n3785), .Y(n11096) );
  NOR2BX1 U3002 ( .AN(net98380), .B(n4438), .Y(n4437) );
  NAND2X1 U3003 ( .A(DCACHE_addr[12]), .B(n4674), .Y(net98380) );
  NAND2X1 U3004 ( .A(n9138), .B(n9137), .Y(n9168) );
  XOR2X1 U3005 ( .A(n10178), .B(n4661), .Y(n11162) );
  INVX16 U3006 ( .A(n4057), .Y(DCACHE_addr[2]) );
  CLKINVX1 U3007 ( .A(n4663), .Y(n4057) );
  NAND2X1 U3008 ( .A(n4434), .B(n11060), .Y(n4530) );
  INVX3 U3009 ( .A(n5012), .Y(n5007) );
  CLKBUFX3 U3010 ( .A(n4934), .Y(n4904) );
  MX2XL U3011 ( .A(\D_cache/cache[7][83] ), .B(n11006), .S0(n5006), .Y(
        \D_cache/n1125 ) );
  MX2XL U3012 ( .A(\D_cache/cache[6][83] ), .B(n11006), .S0(n4962), .Y(
        \D_cache/n1126 ) );
  MX2XL U3013 ( .A(\D_cache/cache[3][83] ), .B(n11006), .S0(n4852), .Y(
        \D_cache/n1129 ) );
  INVX3 U3014 ( .A(n4742), .Y(n4732) );
  CLKINVX1 U3015 ( .A(n11202), .Y(n3954) );
  CLKINVX1 U3016 ( .A(n11203), .Y(n3960) );
  MX2XL U3017 ( .A(\D_cache/cache[0][119] ), .B(n10948), .S0(n4741), .Y(
        \D_cache/n844 ) );
  MX2XL U3018 ( .A(\D_cache/cache[0][0] ), .B(n182), .S0(n4741), .Y(
        \D_cache/n1795 ) );
  MX2XL U3019 ( .A(\D_cache/cache[0][23] ), .B(n10942), .S0(n4741), .Y(
        \D_cache/n1612 ) );
  INVX3 U3020 ( .A(n4811), .Y(n4808) );
  MX2XL U3021 ( .A(\D_cache/cache[0][39] ), .B(n10886), .S0(n4737), .Y(
        \D_cache/n1484 ) );
  MX2XL U3022 ( .A(\D_cache/cache[0][89] ), .B(n3337), .S0(n4737), .Y(
        \D_cache/n1084 ) );
  MX2X1 U3023 ( .A(\D_cache/cache[0][95] ), .B(n10879), .S0(n4737), .Y(
        \D_cache/n1036 ) );
  CLKINVX1 U3024 ( .A(n11499), .Y(n3733) );
  CLKINVX1 U3025 ( .A(n4413), .Y(n3860) );
  AND2X2 U3026 ( .A(net98351), .B(net98352), .Y(n4413) );
  INVX3 U3027 ( .A(n4967), .Y(n4958) );
  INVX3 U3028 ( .A(n4858), .Y(n4848) );
  INVX3 U3029 ( .A(n4812), .Y(n4804) );
  INVX3 U3030 ( .A(n5012), .Y(n5003) );
  INVX3 U3031 ( .A(n4966), .Y(n4959) );
  INVX3 U3032 ( .A(n263), .Y(n4849) );
  INVX3 U3033 ( .A(n4811), .Y(n4805) );
  INVX3 U3034 ( .A(n4787), .Y(n4781) );
  INVX3 U3035 ( .A(n4787), .Y(n4783) );
  INVX3 U3036 ( .A(n4946), .Y(n4938) );
  INVX3 U3037 ( .A(n4946), .Y(n4940) );
  INVX3 U3038 ( .A(n5015), .Y(n5002) );
  MX2XL U3039 ( .A(\D_cache/cache[0][82] ), .B(n3339), .S0(n4733), .Y(
        \D_cache/n1140 ) );
  MX2XL U3040 ( .A(\D_cache/cache[0][85] ), .B(n3341), .S0(n4733), .Y(
        \D_cache/n1116 ) );
  MX2XL U3041 ( .A(\D_cache/cache[0][84] ), .B(n3340), .S0(n4733), .Y(
        \D_cache/n1124 ) );
  MX2XL U3042 ( .A(\D_cache/cache[0][21] ), .B(n10669), .S0(n4733), .Y(
        \D_cache/n1628 ) );
  MX2XL U3043 ( .A(\D_cache/cache[0][50] ), .B(n10513), .S0(n4733), .Y(
        \D_cache/n1396 ) );
  INVX3 U3044 ( .A(n4856), .Y(n4854) );
  INVX3 U3045 ( .A(n5029), .Y(n5008) );
  INVX3 U3046 ( .A(n4997), .Y(n4964) );
  INVX3 U3047 ( .A(n4810), .Y(n4809) );
  INVX3 U3048 ( .A(n4857), .Y(n4850) );
  INVX3 U3049 ( .A(n4818), .Y(n4806) );
  INVX3 U3050 ( .A(n4860), .Y(n4846) );
  INVX3 U3051 ( .A(n4815), .Y(n4801) );
  BUFX16 U3052 ( .A(n12949), .Y(DCACHE_addr[8]) );
  CLKBUFX3 U3053 ( .A(n11510), .Y(n4637) );
  BUFX16 U3054 ( .A(n12928), .Y(DCACHE_addr[29]) );
  BUFX16 U3055 ( .A(n12935), .Y(DCACHE_addr[22]) );
  INVX3 U3056 ( .A(n5023), .Y(n5000) );
  INVX3 U3057 ( .A(n4967), .Y(n4956) );
  AO22X2 U3058 ( .A0(n5528), .A1(DCACHE_addr[13]), .B0(n5526), .B1(n11491), 
        .Y(n11020) );
  BUFX16 U3059 ( .A(n12944), .Y(DCACHE_addr[13]) );
  MX2XL U3060 ( .A(\D_cache/cache[4][14] ), .B(n10743), .S0(n4897), .Y(
        \D_cache/n1680 ) );
  MX2XL U3061 ( .A(\D_cache/cache[4][45] ), .B(n10735), .S0(n4897), .Y(
        \D_cache/n1432 ) );
  MX2XL U3062 ( .A(\D_cache/cache[4][78] ), .B(n3350), .S0(n4897), .Y(
        \D_cache/n1168 ) );
  MX2XL U3063 ( .A(\D_cache/cache[4][76] ), .B(n3352), .S0(n4897), .Y(
        \D_cache/n1184 ) );
  MX2XL U3064 ( .A(\D_cache/cache[4][77] ), .B(n3351), .S0(n4897), .Y(
        \D_cache/n1176 ) );
  MX2XL U3065 ( .A(\D_cache/cache[4][13] ), .B(n10732), .S0(n4897), .Y(
        \D_cache/n1688 ) );
  MX2XL U3066 ( .A(\D_cache/cache[7][14] ), .B(n10743), .S0(n5005), .Y(
        \D_cache/n1677 ) );
  MX2XL U3067 ( .A(\D_cache/cache[7][45] ), .B(n10735), .S0(n5005), .Y(
        \D_cache/n1429 ) );
  MX2XL U3068 ( .A(\D_cache/cache[7][78] ), .B(n3350), .S0(n5005), .Y(
        \D_cache/n1165 ) );
  MX2XL U3069 ( .A(\D_cache/cache[7][76] ), .B(n3352), .S0(n5005), .Y(
        \D_cache/n1181 ) );
  MX2XL U3070 ( .A(\D_cache/cache[7][77] ), .B(n3351), .S0(n5005), .Y(
        \D_cache/n1173 ) );
  MX2XL U3071 ( .A(\D_cache/cache[7][13] ), .B(n10732), .S0(n5005), .Y(
        \D_cache/n1685 ) );
  MX2XL U3072 ( .A(\D_cache/cache[6][14] ), .B(n10743), .S0(n4961), .Y(
        \D_cache/n1678 ) );
  MX2XL U3073 ( .A(\D_cache/cache[6][45] ), .B(n10735), .S0(n4961), .Y(
        \D_cache/n1430 ) );
  MX2XL U3074 ( .A(\D_cache/cache[6][78] ), .B(n3350), .S0(n4961), .Y(
        \D_cache/n1166 ) );
  MX2XL U3075 ( .A(\D_cache/cache[6][76] ), .B(n3352), .S0(n4961), .Y(
        \D_cache/n1182 ) );
  MX2XL U3076 ( .A(\D_cache/cache[6][77] ), .B(n3351), .S0(n4961), .Y(
        \D_cache/n1174 ) );
  MX2XL U3077 ( .A(\D_cache/cache[6][13] ), .B(n10732), .S0(n4961), .Y(
        \D_cache/n1686 ) );
  MX2XL U3078 ( .A(\D_cache/cache[3][14] ), .B(n10743), .S0(n4851), .Y(
        \D_cache/n1681 ) );
  MX2XL U3079 ( .A(\D_cache/cache[3][45] ), .B(n10735), .S0(n4851), .Y(
        \D_cache/n1433 ) );
  MX2XL U3080 ( .A(\D_cache/cache[3][78] ), .B(n3350), .S0(n4851), .Y(
        \D_cache/n1169 ) );
  MX2XL U3081 ( .A(\D_cache/cache[3][76] ), .B(n3352), .S0(n4851), .Y(
        \D_cache/n1185 ) );
  MX2XL U3082 ( .A(\D_cache/cache[3][77] ), .B(n3351), .S0(n4851), .Y(
        \D_cache/n1177 ) );
  MX2XL U3083 ( .A(\D_cache/cache[3][13] ), .B(n10732), .S0(n4851), .Y(
        \D_cache/n1689 ) );
  MX2XL U3084 ( .A(\D_cache/cache[2][14] ), .B(n10743), .S0(n4807), .Y(
        \D_cache/n1682 ) );
  MX2XL U3085 ( .A(\D_cache/cache[2][45] ), .B(n10735), .S0(n4807), .Y(
        \D_cache/n1434 ) );
  MX2XL U3086 ( .A(\D_cache/cache[2][78] ), .B(n3350), .S0(n4807), .Y(
        \D_cache/n1170 ) );
  MX2XL U3087 ( .A(\D_cache/cache[2][76] ), .B(n3352), .S0(n4807), .Y(
        \D_cache/n1186 ) );
  MX2XL U3088 ( .A(\D_cache/cache[2][77] ), .B(n3351), .S0(n4807), .Y(
        \D_cache/n1178 ) );
  MX2XL U3089 ( .A(\D_cache/cache[2][13] ), .B(n10732), .S0(n4807), .Y(
        \D_cache/n1690 ) );
  INVX3 U3090 ( .A(n4918), .Y(n4896) );
  INVX3 U3091 ( .A(n5012), .Y(n5004) );
  INVX3 U3092 ( .A(n4966), .Y(n4960) );
  INVX3 U3093 ( .A(n4859), .Y(n4847) );
  INVX3 U3094 ( .A(n4814), .Y(n4802) );
  MX2XL U3095 ( .A(\D_cache/cache[0][112] ), .B(n10296), .S0(n4734), .Y(
        \D_cache/n900 ) );
  MX2XL U3096 ( .A(\D_cache/cache[0][3] ), .B(n9992), .S0(n4734), .Y(
        \D_cache/n1772 ) );
  MX2XL U3097 ( .A(\D_cache/cache[0][6] ), .B(n10069), .S0(n4734), .Y(
        \D_cache/n1748 ) );
  MX2XL U3098 ( .A(\D_cache/cache[0][70] ), .B(n3338), .S0(n4734), .Y(
        \D_cache/n1236 ) );
  MX2XL U3099 ( .A(\D_cache/cache[0][94] ), .B(n3342), .S0(n4734), .Y(
        \D_cache/n1044 ) );
  MX2XL U3100 ( .A(\D_cache/cache[0][126] ), .B(n166), .S0(n4734), .Y(
        \D_cache/n788 ) );
  MX2XL U3101 ( .A(\D_cache/cache[0][48] ), .B(n10293), .S0(n4734), .Y(
        \D_cache/n1412 ) );
  MX2XL U3102 ( .A(\D_cache/cache[0][62] ), .B(n10144), .S0(n4734), .Y(
        \D_cache/n1300 ) );
  AO22X2 U3103 ( .A0(n5528), .A1(n12941), .B0(n5526), .B1(n11494), .Y(n11016)
         );
  AO22X2 U3104 ( .A0(n5528), .A1(n12940), .B0(n5526), .B1(n11495), .Y(n11010)
         );
  CLKMX2X2 U3105 ( .A(\D_cache/cache[7][94] ), .B(n3342), .S0(n5007), .Y(
        \D_cache/n1037 ) );
  CLKMX2X2 U3106 ( .A(\D_cache/cache[6][94] ), .B(n3342), .S0(n4960), .Y(
        \D_cache/n1038 ) );
  CLKMX2X2 U3107 ( .A(\D_cache/cache[3][94] ), .B(n3342), .S0(n4850), .Y(
        \D_cache/n1041 ) );
  CLKMX2X2 U3108 ( .A(\D_cache/cache[2][94] ), .B(n3342), .S0(n4803), .Y(
        \D_cache/n1042 ) );
  INVX3 U3109 ( .A(n4813), .Y(n4803) );
  MXI2X2 U3110 ( .A(n10988), .B(n10987), .S0(n5523), .Y(n10989) );
  MXI2X2 U3111 ( .A(n10996), .B(n10995), .S0(n5523), .Y(n10997) );
  MXI2X2 U3112 ( .A(n10985), .B(n10984), .S0(n5523), .Y(n10986) );
  MXI2X2 U3113 ( .A(n10932), .B(n10931), .S0(n5521), .Y(n10933) );
  MXI2X1 U3114 ( .A(n10903), .B(n10902), .S0(n5521), .Y(n10904) );
  MXI2X2 U3115 ( .A(n10912), .B(n10911), .S0(n5521), .Y(n10913) );
  MXI2X2 U3116 ( .A(n10909), .B(n10908), .S0(n5521), .Y(n10910) );
  MXI2X2 U3117 ( .A(n10906), .B(n10905), .S0(n5521), .Y(n10907) );
  MXI2X2 U3118 ( .A(n10915), .B(n10914), .S0(n5521), .Y(n10916) );
  MXI2X2 U3119 ( .A(n10929), .B(n10928), .S0(n5521), .Y(n10930) );
  CLKMX2X2 U3120 ( .A(\D_cache/cache[6][84] ), .B(n3340), .S0(n4957), .Y(
        \D_cache/n1118 ) );
  CLKMX2X2 U3121 ( .A(\D_cache/cache[6][85] ), .B(n3341), .S0(n4957), .Y(
        \D_cache/n1110 ) );
  INVX3 U3122 ( .A(n4966), .Y(n4957) );
  CLKMX2X2 U3123 ( .A(\D_cache/cache[7][84] ), .B(n3340), .S0(n5001), .Y(
        \D_cache/n1117 ) );
  CLKMX2X2 U3124 ( .A(\D_cache/cache[7][85] ), .B(n3341), .S0(n5001), .Y(
        \D_cache/n1109 ) );
  CLKMX2X2 U3125 ( .A(\D_cache/cache[7][82] ), .B(n3339), .S0(n5001), .Y(
        \D_cache/n1133 ) );
  INVX3 U3126 ( .A(n5030), .Y(n5001) );
  INVX12 U3127 ( .A(n407), .Y(mem_wdata_D[82]) );
  CLKAND2X12 U3128 ( .A(n5557), .B(n11233), .Y(mem_wdata_I[47]) );
  CLKAND2X12 U3129 ( .A(n4653), .B(n11423), .Y(mem_wdata_D[73]) );
  CLKAND2X12 U3130 ( .A(n4653), .B(n11429), .Y(mem_wdata_D[79]) );
  CLKAND2X12 U3131 ( .A(n5557), .B(n11201), .Y(mem_wdata_I[15]) );
  CLKAND2X12 U3132 ( .A(mem_write_I), .B(n11252), .Y(mem_wdata_I[66]) );
  CLKAND2X12 U3133 ( .A(n5557), .B(n11220), .Y(mem_wdata_I[34]) );
  BUFX12 U3134 ( .A(n5554), .Y(n5557) );
  CLKAND2X12 U3135 ( .A(n5556), .B(n11312), .Y(mem_wdata_I[126]) );
  BUFX4 U3136 ( .A(n5525), .Y(n5515) );
  CLKAND2X12 U3137 ( .A(n5551), .B(n11397), .Y(mem_wdata_D[47]) );
  CLKAND2X12 U3138 ( .A(n5551), .B(n11351), .Y(mem_wdata_D[1]) );
  CLKAND2X12 U3139 ( .A(n5551), .B(n11383), .Y(mem_wdata_D[33]) );
  CLKAND2X12 U3140 ( .A(n5551), .B(n11420), .Y(mem_wdata_D[70]) );
  CLKAND2X12 U3141 ( .A(n5551), .B(n11402), .Y(mem_wdata_D[52]) );
  CLKAND2X12 U3142 ( .A(n5551), .B(n11435), .Y(mem_wdata_D[85]) );
  CLKAND2X12 U3143 ( .A(n5551), .B(n11359), .Y(mem_wdata_D[9]) );
  CLKAND2X12 U3144 ( .A(n5551), .B(n11391), .Y(mem_wdata_D[41]) );
  CLKAND2X12 U3145 ( .A(n5551), .B(n11385), .Y(mem_wdata_D[35]) );
  CLKAND2X12 U3146 ( .A(n5551), .B(n11381), .Y(mem_wdata_D[31]) );
  BUFX12 U3147 ( .A(n11511), .Y(mem_write_D) );
  AO22X2 U3148 ( .A0(n5528), .A1(DCACHE_addr[20]), .B0(n5527), .B1(n11498), 
        .Y(n11034) );
  BUFX16 U3149 ( .A(n12937), .Y(DCACHE_addr[20]) );
  INVX12 U3150 ( .A(n1948), .Y(mem_addr_D[7]) );
  INVXL U3151 ( .A(n12797), .Y(n3619) );
  INVX12 U3152 ( .A(n3619), .Y(mem_addr_D[8]) );
  AO22X1 U3153 ( .A0(DCACHE_addr[6]), .A1(n11510), .B0(n4654), .B1(n11484), 
        .Y(n12797) );
  INVXL U3154 ( .A(n12796), .Y(n3621) );
  INVX12 U3155 ( .A(n3621), .Y(mem_addr_D[9]) );
  AO22X1 U3156 ( .A0(DCACHE_addr[7]), .A1(n11510), .B0(n4653), .B1(n11485), 
        .Y(n12796) );
  INVX12 U3157 ( .A(n1949), .Y(mem_addr_D[10]) );
  INVX12 U3158 ( .A(n1950), .Y(mem_addr_D[12]) );
  INVX12 U3159 ( .A(n1951), .Y(mem_addr_D[18]) );
  INVX12 U3160 ( .A(n1952), .Y(mem_addr_D[19]) );
  INVX12 U3161 ( .A(n1944), .Y(mem_wdata_D[26]) );
  CLKAND2X12 U3162 ( .A(n5551), .B(n11354), .Y(mem_wdata_D[4]) );
  CLKAND2X12 U3163 ( .A(n5551), .B(n11360), .Y(mem_wdata_D[10]) );
  CLKAND2X12 U3164 ( .A(n5551), .B(n11370), .Y(mem_wdata_D[20]) );
  CLKAND2X12 U3165 ( .A(n5551), .B(n11366), .Y(mem_wdata_D[16]) );
  CLKAND2X12 U3166 ( .A(n5551), .B(n11392), .Y(mem_wdata_D[42]) );
  CLKAND2X12 U3167 ( .A(n5551), .B(n11369), .Y(mem_wdata_D[19]) );
  CLKAND2X12 U3168 ( .A(n5551), .B(n11379), .Y(mem_wdata_D[29]) );
  CLKAND2X12 U3169 ( .A(n5551), .B(n11371), .Y(mem_wdata_D[21]) );
  CLKAND2X12 U3170 ( .A(n5551), .B(n11355), .Y(mem_wdata_D[5]) );
  CLKAND2X12 U3171 ( .A(n5551), .B(n11353), .Y(mem_wdata_D[3]) );
  CLKAND2X12 U3172 ( .A(n5551), .B(n11377), .Y(mem_wdata_D[27]) );
  INVX12 U3173 ( .A(n1947), .Y(mem_wdata_D[80]) );
  CLKAND2X12 U3174 ( .A(n4653), .B(n11475), .Y(mem_wdata_D[125]) );
  CLKAND2X12 U3175 ( .A(n4653), .B(n11472), .Y(mem_wdata_D[122]) );
  CLKAND2X12 U3176 ( .A(n4653), .B(n11418), .Y(mem_wdata_D[68]) );
  CLKAND2X12 U3177 ( .A(n4653), .B(n11448), .Y(mem_wdata_D[98]) );
  CLKAND2X12 U3178 ( .A(n5551), .B(n11405), .Y(mem_wdata_D[55]) );
  CLKAND2X12 U3179 ( .A(n11511), .B(n11398), .Y(mem_wdata_D[48]) );
  CLKAND2X12 U3180 ( .A(n11511), .B(n11438), .Y(mem_wdata_D[88]) );
  INVX12 U3181 ( .A(n1945), .Y(mem_wdata_D[49]) );
  CLKAND2X12 U3182 ( .A(n11511), .B(n11465), .Y(mem_wdata_D[115]) );
  INVX12 U3183 ( .A(n1940), .Y(mem_wdata_D[2]) );
  INVX12 U3184 ( .A(n1941), .Y(mem_wdata_D[6]) );
  CLKAND2X12 U3185 ( .A(n4653), .B(n11378), .Y(mem_wdata_D[28]) );
  INVX12 U3186 ( .A(n1943), .Y(mem_wdata_D[22]) );
  INVX12 U3187 ( .A(n1946), .Y(mem_wdata_D[54]) );
  CLKAND2X12 U3188 ( .A(n3737), .B(n11358), .Y(mem_wdata_D[8]) );
  CLKAND2X12 U3189 ( .A(n4654), .B(n11362), .Y(mem_wdata_D[12]) );
  CLKAND2X12 U3190 ( .A(n4654), .B(n11364), .Y(mem_wdata_D[14]) );
  CLKAND2X12 U3191 ( .A(n4654), .B(n11368), .Y(mem_wdata_D[18]) );
  CLKAND2X12 U3192 ( .A(n3737), .B(n11380), .Y(mem_wdata_D[30]) );
  BUFX16 U3193 ( .A(n4296), .Y(DCACHE_addr[4]) );
  INVX3 U3194 ( .A(n4948), .Y(n4941) );
  INVX3 U3195 ( .A(n4249), .Y(n4942) );
  INVX12 U3196 ( .A(n3735), .Y(net100573) );
  NOR3X6 U3197 ( .A(n4620), .B(n11003), .C(n9980), .Y(n11348) );
  BUFX20 U3198 ( .A(n5549), .Y(n4620) );
  CLKINVX3 U3199 ( .A(n3746), .Y(n3747) );
  NOR2X1 U3200 ( .A(n6545), .B(\i_MIPS/ALUin1[11] ), .Y(n3634) );
  NOR4X2 U3201 ( .A(n9211), .B(n9210), .C(n9209), .D(n9208), .Y(n9212) );
  CLKINVX1 U3202 ( .A(n10083), .Y(n10085) );
  INVX2 U3203 ( .A(n4163), .Y(n3635) );
  NAND2X4 U3204 ( .A(n6561), .B(\i_MIPS/n359 ), .Y(n7688) );
  CLKBUFX16 U3205 ( .A(net100424), .Y(net111634) );
  INVX6 U3206 ( .A(net133317), .Y(net100424) );
  CLKAND2X12 U3207 ( .A(net111640), .B(net111636), .Y(net128830) );
  INVX3 U3208 ( .A(n6604), .Y(n9883) );
  CLKMX2X4 U3209 ( .A(\i_MIPS/n319 ), .B(n4540), .S0(\i_MIPS/ID_EX_5 ), .Y(
        n6604) );
  CLKINVX16 U3210 ( .A(n5626), .Y(n5624) );
  INVX8 U3211 ( .A(net100399), .Y(net100397) );
  AND4X6 U3212 ( .A(n3935), .B(n3936), .C(n3934), .D(n3933), .Y(net102784) );
  INVX12 U3213 ( .A(net100401), .Y(net100396) );
  AND2X2 U3214 ( .A(net108658), .B(n3637), .Y(n4415) );
  AO22X1 U3215 ( .A0(n4720), .A1(n981), .B0(n4719), .B1(n2496), .Y(n9517) );
  CLKINVX1 U3216 ( .A(n7232), .Y(n3636) );
  CLKAND2X12 U3217 ( .A(n7702), .B(n7701), .Y(n4150) );
  BUFX2 U3218 ( .A(n5128), .Y(n5103) );
  INVX6 U3219 ( .A(n9153), .Y(n8862) );
  NOR2X4 U3220 ( .A(n6573), .B(\i_MIPS/ALUin1[17] ), .Y(n3638) );
  NAND2X4 U3221 ( .A(n4321), .B(n4570), .Y(n9141) );
  INVX12 U3222 ( .A(net112356), .Y(net112348) );
  BUFX2 U3223 ( .A(n5310), .Y(n5282) );
  NAND2X6 U3224 ( .A(n3891), .B(n10866), .Y(n6749) );
  BUFX12 U3225 ( .A(n12953), .Y(n4663) );
  AND3X4 U3226 ( .A(n6704), .B(n6705), .C(net112296), .Y(n6713) );
  BUFX6 U3227 ( .A(net128151), .Y(net112340) );
  INVX4 U3228 ( .A(net112340), .Y(net112332) );
  OAI221X2 U3229 ( .A0(net112366), .A1(\i_MIPS/n351 ), .B0(net112348), .B1(
        \i_MIPS/n352 ), .C0(n6766), .Y(n7813) );
  NAND4X4 U3230 ( .A(n6007), .B(n6006), .C(n6005), .D(n6004), .Y(n11323) );
  NAND2X2 U3231 ( .A(\i_MIPS/ALUin1[28] ), .B(n6589), .Y(n8432) );
  CLKMX2X12 U3232 ( .A(\i_MIPS/n273 ), .B(n4494), .S0(n5622), .Y(n6574) );
  CLKMX2X2 U3233 ( .A(net103721), .B(net103722), .S0(net107812), .Y(net103718)
         );
  OAI221XL U3234 ( .A0(n9116), .A1(net111622), .B0(net111634), .B1(n9115), 
        .C0(n9114), .Y(n4615) );
  AOI32X2 U3235 ( .A0(n8627), .A1(net111910), .A2(n3690), .B0(n8604), .B1(
        net111910), .Y(n8605) );
  NAND2X1 U3236 ( .A(\i_MIPS/ALUin1[8] ), .B(n7495), .Y(n7219) );
  NAND2X2 U3237 ( .A(net102427), .B(n8338), .Y(n3639) );
  AND2X8 U3238 ( .A(n6540), .B(n3640), .Y(n6969) );
  INVX3 U3239 ( .A(n3639), .Y(n3640) );
  NAND2X6 U3240 ( .A(n6539), .B(\i_MIPS/n368 ), .Y(n8338) );
  CLKMX2X2 U3241 ( .A(n8823), .B(n8822), .S0(net107812), .Y(n8826) );
  OA22X2 U3242 ( .A0(net133471), .A1(n7617), .B0(n7616), .B1(n7901), .Y(n7623)
         );
  CLKMX2X8 U3243 ( .A(n10), .B(n7314), .S0(net107798), .Y(n8959) );
  NAND2X1 U3244 ( .A(n7503), .B(n4381), .Y(n7507) );
  NAND2X4 U3245 ( .A(n8339), .B(n7503), .Y(n6968) );
  INVX6 U3246 ( .A(n11436), .Y(n10212) );
  OAI2BB2X1 U3247 ( .B0(net112306), .B1(n8946), .A0N(n9481), .A1N(net137952), 
        .Y(n7612) );
  INVX16 U3248 ( .A(net112300), .Y(net112296) );
  MXI2X2 U3249 ( .A(n10216), .B(n10215), .S0(n5513), .Y(n10217) );
  AOI222XL U3250 ( .A0(n5504), .A1(n11372), .B0(mem_rdata_D[22]), .B1(n232), 
        .C0(n12965), .C1(n5501), .Y(n10216) );
  NAND2X4 U3251 ( .A(n6573), .B(\i_MIPS/n354 ), .Y(n8750) );
  NAND2X4 U3252 ( .A(\i_MIPS/ALUin1[17] ), .B(n6573), .Y(n8539) );
  OA22X1 U3253 ( .A0(n4755), .A1(n1208), .B0(n4793), .B1(n2745), .Y(n7355) );
  BUFX12 U3254 ( .A(n4797), .Y(n4793) );
  NAND3X8 U3255 ( .A(n4311), .B(n4312), .C(n7045), .Y(n7218) );
  OR2X8 U3256 ( .A(n7047), .B(n7046), .Y(n4312) );
  AND3X8 U3257 ( .A(\i_MIPS/ALU_Control/n11 ), .B(\i_MIPS/n323 ), .C(
        \i_MIPS/ALU_Control/n18 ), .Y(n4379) );
  INVX8 U3258 ( .A(net105600), .Y(net103910) );
  NAND3X6 U3259 ( .A(n3706), .B(n6983), .C(n6982), .Y(net97684) );
  NAND2BX4 U3260 ( .AN(n8536), .B(n8738), .Y(n8537) );
  AOI2BB1X4 U3261 ( .A0N(n9044), .A1N(n8449), .B0(n8450), .Y(n8434) );
  CLKAND2X12 U3262 ( .A(n11067), .B(n10176), .Y(n4456) );
  OA22X2 U3263 ( .A0(n5390), .A1(n1458), .B0(n5332), .B1(n3032), .Y(n6147) );
  NAND3BX1 U3264 ( .AN(n9046), .B(n9065), .C(n9066), .Y(n3641) );
  INVX3 U3265 ( .A(n9041), .Y(n9046) );
  CLKINVX12 U3266 ( .A(n9269), .Y(n3825) );
  OA22XL U3267 ( .A0(n5302), .A1(n1287), .B0(n5256), .B1(n2820), .Y(n9999) );
  OA22XL U3268 ( .A0(n5302), .A1(n1288), .B0(n5256), .B1(n2821), .Y(n10018) );
  OA22XL U3269 ( .A0(n5302), .A1(n3217), .B0(n5256), .B1(n1420), .Y(n9994) );
  OA22X1 U3270 ( .A0(n5302), .A1(n1209), .B0(n5256), .B1(n2746), .Y(n10004) );
  OR2X4 U3271 ( .A(net104407), .B(net111624), .Y(n3642) );
  OR2X4 U3272 ( .A(net104408), .B(net111636), .Y(n3643) );
  CLKMX2X4 U3273 ( .A(n8439), .B(n8438), .S0(net107798), .Y(n9247) );
  CLKBUFX3 U3274 ( .A(net100535), .Y(net111964) );
  INVX12 U3275 ( .A(net101978), .Y(net100535) );
  NAND3X6 U3276 ( .A(n3789), .B(n3790), .C(net104889), .Y(net97755) );
  AND3X2 U3277 ( .A(n6449), .B(n6448), .C(n6447), .Y(n6450) );
  NAND4X4 U3278 ( .A(n9901), .B(n9900), .C(n9899), .D(n9898), .Y(n11190) );
  INVX3 U3279 ( .A(n8551), .Y(n8552) );
  INVX20 U3280 ( .A(n5548), .Y(n5546) );
  CLKINVX20 U3281 ( .A(n4671), .Y(n4669) );
  AND2X8 U3282 ( .A(n3426), .B(net99118), .Y(n3817) );
  NAND3X6 U3283 ( .A(n3644), .B(n3645), .C(n3646), .Y(n3647) );
  NAND2X6 U3284 ( .A(n3647), .B(n6522), .Y(n3905) );
  CLKINVX3 U3285 ( .A(n6524), .Y(n3645) );
  INVX3 U3286 ( .A(n6523), .Y(n3646) );
  NOR2X2 U3287 ( .A(n8227), .B(n8232), .Y(n3648) );
  NOR2X4 U3288 ( .A(n8232), .B(n8229), .Y(n3649) );
  OR3X6 U3289 ( .A(n3648), .B(n3649), .C(n8945), .Y(n8941) );
  AOI2BB1X4 U3290 ( .A0N(n8942), .A1N(n8941), .B0(n8940), .Y(n8943) );
  NAND4BX2 U3291 ( .AN(n9014), .B(n9013), .C(n9012), .D(n9011), .Y(n9015) );
  NOR4X4 U3292 ( .A(n9261), .B(n9260), .C(n9259), .D(n9258), .Y(n9287) );
  INVX6 U3293 ( .A(net97800), .Y(net102938) );
  MX2X6 U3294 ( .A(n7300), .B(n7317), .S0(net107796), .Y(n6978) );
  OR2X4 U3295 ( .A(n9462), .B(net101914), .Y(n4308) );
  NAND2X4 U3296 ( .A(n7495), .B(\i_MIPS/n363 ), .Y(n8636) );
  NAND3X6 U3297 ( .A(n3759), .B(n3760), .C(net103091), .Y(n4134) );
  AO22X1 U3298 ( .A0(n4713), .A1(n280), .B0(n4708), .B1(n2497), .Y(n7962) );
  NAND2X4 U3299 ( .A(n7410), .B(n3636), .Y(n7685) );
  OA22X1 U3300 ( .A0(n4828), .A1(n1078), .B0(n4873), .B1(n2656), .Y(n7278) );
  BUFX4 U3301 ( .A(n4991), .Y(n4980) );
  OAI211X4 U3302 ( .A0(n4416), .A1(n8751), .B0(n8750), .C0(n8749), .Y(n8755)
         );
  AOI2BB1X4 U3303 ( .A0N(n2210), .A1N(n9140), .B0(n9139), .Y(n9143) );
  CLKINVX12 U3304 ( .A(net100426), .Y(net111646) );
  NAND3BX4 U3305 ( .AN(n7520), .B(n7692), .C(n7798), .Y(n7525) );
  NAND2X6 U3306 ( .A(\i_MIPS/ALUin1[13] ), .B(n6547), .Y(n7692) );
  NAND2X6 U3307 ( .A(n10679), .B(n10678), .Y(n9221) );
  INVX3 U3308 ( .A(n9149), .Y(n9147) );
  XNOR2X1 U3309 ( .A(n6605), .B(\i_MIPS/IR_ID[16] ), .Y(n4532) );
  INVX20 U3310 ( .A(net111630), .Y(net111622) );
  INVX1 U3311 ( .A(n11474), .Y(n10475) );
  INVX20 U3312 ( .A(net108710), .Y(net108702) );
  CLKMX2X12 U3313 ( .A(n7815), .B(n9059), .S0(net107798), .Y(n6770) );
  NAND2X6 U3314 ( .A(n7306), .B(n7406), .Y(n4304) );
  AND2X8 U3315 ( .A(n4304), .B(n4305), .Y(n4484) );
  BUFX2 U3316 ( .A(n5128), .Y(n5102) );
  AO21X2 U3317 ( .A0(n10521), .A1(net98375), .B0(net111642), .Y(net103418) );
  NAND2X6 U3318 ( .A(n6555), .B(\i_MIPS/n357 ), .Y(n7610) );
  INVX3 U3319 ( .A(net112176), .Y(net112166) );
  NAND4X6 U3320 ( .A(n4329), .B(n6365), .C(n6364), .D(n6363), .Y(n11492) );
  BUFX4 U3321 ( .A(n4928), .Y(n4926) );
  INVX16 U3322 ( .A(n4570), .Y(n8946) );
  NAND3BX2 U3323 ( .AN(n6520), .B(n8231), .C(n8534), .Y(n6515) );
  NAND2X4 U3324 ( .A(n8553), .B(n9263), .Y(n9142) );
  AOI222X2 U3325 ( .A0(net101908), .A1(n4125), .B0(net103548), .B1(n4126), 
        .C0(net101402), .C1(net101401), .Y(net105007) );
  NAND2X6 U3326 ( .A(net101910), .B(n4536), .Y(n7234) );
  NAND2X6 U3327 ( .A(n9165), .B(n4536), .Y(n9336) );
  NAND2X1 U3328 ( .A(\i_MIPS/ID_EX[81] ), .B(n4536), .Y(n8651) );
  BUFX8 U3329 ( .A(net129024), .Y(net108662) );
  AOI22X2 U3330 ( .A0(n10601), .A1(n3897), .B0(n637), .B1(net108662), .Y(
        n10606) );
  OR2X2 U3331 ( .A(n9454), .B(n7901), .Y(n4307) );
  CLKAND2X2 U3332 ( .A(\i_MIPS/ALUin1[0] ), .B(net112338), .Y(n4520) );
  AND3X4 U3333 ( .A(\i_MIPS/ID_EX[78] ), .B(\i_MIPS/ID_EX[73] ), .C(
        \i_MIPS/ID_EX[75] ), .Y(n4541) );
  OA21X2 U3334 ( .A0(n7480), .A1(n7479), .B0(n9330), .Y(n7483) );
  NAND2X4 U3335 ( .A(n4505), .B(n4501), .Y(n9412) );
  BUFX4 U3336 ( .A(n9533), .Y(n4722) );
  AND2X8 U3337 ( .A(net98620), .B(n4146), .Y(n3652) );
  BUFX8 U3338 ( .A(net97444), .Y(net108686) );
  NAND2BX1 U3339 ( .AN(n4655), .B(n11200), .Y(n3952) );
  NAND2X1 U3340 ( .A(n6121), .B(n4060), .Y(n11315) );
  OA22X1 U3341 ( .A0(n4753), .A1(n1485), .B0(n4792), .B1(n3068), .Y(n4350) );
  BUFX8 U3342 ( .A(n4798), .Y(n4792) );
  MXI2X2 U3343 ( .A(n10734), .B(n10733), .S0(n5518), .Y(n10735) );
  NAND2BX1 U3344 ( .AN(n5428), .B(n11216), .Y(n6285) );
  CLKINVX8 U3345 ( .A(n5623), .Y(n4316) );
  NAND2X8 U3346 ( .A(net101910), .B(n8349), .Y(n7707) );
  OAI2BB2X4 U3347 ( .B0(n3653), .B1(n3654), .A0N(net111966), .A1N(net97800), 
        .Y(net103025) );
  MXI2X2 U3348 ( .A(n8008), .B(n8007), .S0(net107816), .Y(n3654) );
  OA22X4 U3349 ( .A0(n9463), .A1(net101771), .B0(n8732), .B1(n9469), .Y(n8733)
         );
  MX2X1 U3350 ( .A(net112438), .B(net100573), .S0(n8730), .Y(n8735) );
  MXI2X2 U3351 ( .A(n8847), .B(n8846), .S0(\i_MIPS/IR_ID[25] ), .Y(n3655) );
  CLKINVX8 U3352 ( .A(n3734), .Y(net127710) );
  CLKBUFX8 U3353 ( .A(net97444), .Y(net108690) );
  XOR3XL U3354 ( .A(n11094), .B(n11093), .C(n11092), .Y(n11097) );
  NAND2X4 U3355 ( .A(n11094), .B(n11092), .Y(n10363) );
  CLKMX2X2 U3356 ( .A(n7317), .B(net103710), .S0(net107794), .Y(n7316) );
  CLKAND2X12 U3357 ( .A(n5557), .B(n11188), .Y(mem_wdata_I[2]) );
  OA22X1 U3358 ( .A0(n5301), .A1(n1486), .B0(n5256), .B1(n3069), .Y(n9939) );
  CLKMX2X3 U3359 ( .A(n7041), .B(n7040), .S0(net107812), .Y(net104739) );
  NAND4BX2 U3360 ( .AN(n7039), .B(n7038), .C(n7037), .D(n7036), .Y(n7040) );
  INVX8 U3361 ( .A(n10431), .Y(n10434) );
  OA22X1 U3362 ( .A0(n5371), .A1(n1487), .B0(n5344), .B1(n3070), .Y(n9938) );
  NAND2X8 U3363 ( .A(n4618), .B(n7044), .Y(n7400) );
  MXI2X2 U3364 ( .A(n10767), .B(n10766), .S0(n5519), .Y(n10768) );
  CLKINVX2 U3365 ( .A(n9493), .Y(n9489) );
  AND3X2 U3366 ( .A(net103911), .B(n3823), .C(net103913), .Y(net103840) );
  NAND4X4 U3367 ( .A(n9613), .B(n9612), .C(n9611), .D(n9610), .Y(n10611) );
  NAND2BX2 U3368 ( .AN(n5428), .B(n11200), .Y(n9611) );
  NAND4X2 U3369 ( .A(n9598), .B(n9597), .C(n9596), .D(n9595), .Y(n11264) );
  OA22X1 U3370 ( .A0(n5293), .A1(n1080), .B0(n5246), .B1(n2673), .Y(n9596) );
  OA22XL U3371 ( .A0(n5370), .A1(n3071), .B0(n5337), .B1(n1183), .Y(n9595) );
  MXI2X6 U3372 ( .A(\i_MIPS/ID_EX[50] ), .B(n4662), .S0(n5624), .Y(n3686) );
  NOR4X2 U3373 ( .A(n8559), .B(n8558), .C(n8557), .D(n8556), .Y(n8564) );
  NAND2X4 U3374 ( .A(n8349), .B(n9165), .Y(n8555) );
  MX2X1 U3375 ( .A(net100573), .B(net112438), .S0(n9272), .Y(n8554) );
  NAND4X8 U3376 ( .A(n3656), .B(n3657), .C(n6437), .D(n6436), .Y(n11347) );
  AND4X8 U3377 ( .A(n6427), .B(n3906), .C(n6425), .D(n6426), .Y(n3657) );
  OAI2BB1X4 U3378 ( .A0N(n7442), .A1N(n7441), .B0(n3690), .Y(net98372) );
  INVX16 U3379 ( .A(n3697), .Y(n3690) );
  OA21X1 U3380 ( .A0(net112346), .A1(net103561), .B0(n6767), .Y(n6684) );
  NAND2X2 U3381 ( .A(\i_MIPS/ALUin1[8] ), .B(net112370), .Y(n6767) );
  BUFX16 U3382 ( .A(net127709), .Y(net112370) );
  NAND3X4 U3383 ( .A(n3774), .B(n3775), .C(n9114), .Y(n10490) );
  NAND2X4 U3384 ( .A(\i_MIPS/ALUin1[16] ), .B(n6551), .Y(n8753) );
  AO21X4 U3385 ( .A0(n10567), .A1(n10566), .B0(net111640), .Y(n8335) );
  NAND4X6 U3386 ( .A(n7551), .B(n7550), .C(n7549), .D(n7548), .Y(net97736) );
  AOI211X4 U3387 ( .A0(n4498), .A1(net100585), .B0(n7487), .C0(n7486), .Y(
        n7550) );
  NAND2X4 U3388 ( .A(n10065), .B(n9569), .Y(n10638) );
  BUFX4 U3389 ( .A(n5265), .Y(n5241) );
  CLKINVX1 U3390 ( .A(n10377), .Y(n10371) );
  NOR2X4 U3391 ( .A(n7223), .B(n7159), .Y(n7161) );
  AO22X4 U3392 ( .A0(n9161), .A1(n9160), .B0(n9159), .B1(n12), .Y(n9173) );
  XNOR2X2 U3393 ( .A(ICACHE_addr[17]), .B(n11332), .Y(n6093) );
  AO22X4 U3394 ( .A0(mem_rdata_I[39]), .A1(n5543), .B0(n252), .B1(n11225), .Y(
        n10131) );
  OA22X1 U3395 ( .A0(n5103), .A1(n1210), .B0(n5073), .B1(n2747), .Y(n6087) );
  CLKAND2X8 U3396 ( .A(n7053), .B(n7891), .Y(n6509) );
  NAND2X4 U3397 ( .A(\i_MIPS/ALUin1[8] ), .B(n7053), .Y(n8635) );
  CLKBUFX6 U3398 ( .A(n9987), .Y(n4886) );
  NAND2BX1 U3399 ( .AN(n7610), .B(n7798), .Y(n7528) );
  BUFX20 U3400 ( .A(n4296), .Y(n4666) );
  NAND3BX1 U3401 ( .AN(n8967), .B(net111994), .C(n3698), .Y(n8975) );
  NOR2X4 U3402 ( .A(n7404), .B(n3427), .Y(n7408) );
  NAND2X1 U3403 ( .A(n4389), .B(n10399), .Y(n3658) );
  OR2X8 U3404 ( .A(n10238), .B(n10237), .Y(n3659) );
  OR2X4 U3405 ( .A(n409), .B(n10394), .Y(n3660) );
  NAND2X6 U3406 ( .A(n10386), .B(n10389), .Y(n10237) );
  MXI2X2 U3407 ( .A(n6745), .B(n6744), .S0(net107810), .Y(n6746) );
  NAND4X2 U3408 ( .A(n6743), .B(n6742), .C(n6741), .D(n6740), .Y(n6744) );
  NAND2X2 U3409 ( .A(n6545), .B(\i_MIPS/n360 ), .Y(n7500) );
  NAND2X2 U3410 ( .A(n6544), .B(\i_MIPS/n361 ), .Y(n7492) );
  CLKINVX1 U3411 ( .A(n5625), .Y(n3801) );
  OR2X4 U3412 ( .A(net104887), .B(net111624), .Y(n3789) );
  OAI221X4 U3413 ( .A0(\i_MIPS/Register/register[18][2] ), .A1(n4691), .B0(
        \i_MIPS/Register/register[26][2] ), .B1(n4688), .C0(n6951), .Y(n6959)
         );
  OA22X4 U3414 ( .A0(n4997), .A1(n2100), .B0(n5020), .B1(n515), .Y(n9503) );
  OAI221X2 U3415 ( .A0(n9455), .A1(n8876), .B0(n9463), .B1(n8875), .C0(n4658), 
        .Y(n8877) );
  OR2X2 U3416 ( .A(\i_MIPS/n341 ), .B(net112364), .Y(n4161) );
  NAND4BX2 U3417 ( .AN(n4343), .B(n9509), .C(n9508), .D(n9507), .Y(n11372) );
  OA22XL U3418 ( .A0(n4927), .A1(n1574), .B0(n4950), .B1(n3156), .Y(n6314) );
  OA22XL U3419 ( .A0(n4927), .A1(n1456), .B0(n4950), .B1(n3026), .Y(n6322) );
  NAND4X4 U3420 ( .A(n6306), .B(n6305), .C(n6304), .D(n6303), .Y(n6312) );
  OA22X2 U3421 ( .A0(n4927), .A1(n1460), .B0(n4950), .B1(n3034), .Y(n6340) );
  CLKBUFX2 U3422 ( .A(n8737), .Y(n3661) );
  AOI2BB1X4 U3423 ( .A0N(net112306), .A1N(n7172), .B0(net100583), .Y(n7173) );
  CLKINVX12 U3424 ( .A(n3662), .Y(n8532) );
  INVX4 U3425 ( .A(n10621), .Y(n10624) );
  NAND4X4 U3426 ( .A(n10203), .B(n10202), .C(n10201), .D(n10200), .Y(n11173)
         );
  NAND2BX2 U3427 ( .AN(n5429), .B(n11221), .Y(n10200) );
  AOI2BB2X4 U3428 ( .B0(net111968), .B1(n10652), .A0N(n3787), .A1N(n3664), .Y(
        n3663) );
  INVX20 U3429 ( .A(n5547), .Y(n3665) );
  CLKBUFX3 U3430 ( .A(n5357), .Y(n5350) );
  BUFX3 U3431 ( .A(n5349), .Y(n5346) );
  OA22X2 U3432 ( .A0(n5370), .A1(n1461), .B0(n5347), .B1(n3035), .Y(n10117) );
  NOR4X4 U3433 ( .A(n8744), .B(n8743), .C(n8742), .D(n8741), .Y(n8764) );
  NAND2BX1 U3434 ( .AN(n4649), .B(n11406), .Y(n3668) );
  AO21X4 U3435 ( .A0(n8204), .A1(n8203), .B0(n3665), .Y(n4608) );
  OA22X1 U3436 ( .A0(n7618), .A1(net101914), .B0(n9468), .B1(net102404), .Y(
        n7622) );
  AO22X1 U3437 ( .A0(n4713), .A1(n982), .B0(n4708), .B1(n2498), .Y(n7953) );
  NAND2X4 U3438 ( .A(\i_MIPS/ALUin1[17] ), .B(n6553), .Y(n8752) );
  NAND4X2 U3439 ( .A(n6215), .B(n6214), .C(n6213), .D(n6212), .Y(n11248) );
  OA22XL U3440 ( .A0(n5392), .A1(n1575), .B0(n5334), .B1(n3157), .Y(n6212) );
  OA22XL U3441 ( .A0(n5198), .A1(n1576), .B0(n5155), .B1(n3158), .Y(n6214) );
  NAND2BX1 U3442 ( .AN(n4649), .B(n11413), .Y(n3671) );
  NAND2BX2 U3443 ( .AN(n5427), .B(n11194), .Y(n10014) );
  AO22X4 U3444 ( .A0(mem_rdata_I[8]), .A1(n5537), .B0(n252), .B1(n11194), .Y(
        n10007) );
  NAND4X4 U3445 ( .A(n10006), .B(n10005), .C(n10004), .D(n10003), .Y(n11194)
         );
  OA22X1 U3446 ( .A0(n5393), .A1(n1637), .B0(n5345), .B1(n3219), .Y(n10003) );
  NOR4X2 U3447 ( .A(n7035), .B(n7034), .C(n7033), .D(n7032), .Y(n7036) );
  NAND2X2 U3448 ( .A(n6530), .B(\i_MIPS/ALUin1[10] ), .Y(n7496) );
  CLKMX2X8 U3449 ( .A(n9160), .B(n7815), .S0(net107794), .Y(n9057) );
  INVX12 U3450 ( .A(net111646), .Y(net111642) );
  OA22XL U3451 ( .A0(n5195), .A1(n1680), .B0(n5152), .B1(n3271), .Y(n6134) );
  OA22XL U3452 ( .A0(n5195), .A1(n1577), .B0(n5152), .B1(n3159), .Y(n6125) );
  OA22XL U3453 ( .A0(n5195), .A1(n1681), .B0(n5152), .B1(n3272), .Y(n6129) );
  OA22XL U3454 ( .A0(n5195), .A1(n1289), .B0(n5169), .B1(n2822), .Y(n6101) );
  OA22XL U3455 ( .A0(n5195), .A1(n1728), .B0(n5146), .B1(n3335), .Y(n6117) );
  NAND2X2 U3456 ( .A(n4), .B(net105038), .Y(net102429) );
  NAND2X2 U3457 ( .A(n6917), .B(n6916), .Y(net102426) );
  AOI33X2 U3458 ( .A0(n9356), .A1(n9355), .A2(net112292), .B0(net111996), .B1(
        n9353), .B2(n9354), .Y(n9357) );
  NAND4X1 U3459 ( .A(n6324), .B(n6323), .C(n6322), .D(n6321), .Y(n11412) );
  NAND2X4 U3460 ( .A(n1774), .B(net100398), .Y(net100403) );
  INVX8 U3461 ( .A(n5551), .Y(n4649) );
  INVX3 U3462 ( .A(n7901), .Y(n7702) );
  INVX4 U3463 ( .A(n7401), .Y(n7221) );
  INVXL U3464 ( .A(n8641), .Y(n8656) );
  CLKINVX2 U3465 ( .A(n9353), .Y(n9351) );
  NAND2X2 U3466 ( .A(n3825), .B(n9242), .Y(n9483) );
  NAND2BX1 U3467 ( .AN(n4649), .B(n11415), .Y(n3674) );
  AND4X6 U3468 ( .A(n10376), .B(n10375), .C(net97444), .D(net97592), .Y(n3921)
         );
  CLKMX2X3 U3469 ( .A(n7929), .B(n7928), .S0(net107816), .Y(n7930) );
  NOR4X2 U3470 ( .A(n7918), .B(n7917), .C(n7916), .D(n7915), .Y(n7929) );
  AND2X8 U3471 ( .A(n4217), .B(n10246), .Y(n3676) );
  INVX20 U3472 ( .A(net108682), .Y(net108674) );
  OAI2BB2X1 U3473 ( .B0(\i_MIPS/n177 ), .B1(net108190), .A0N(n4072), .A1N(
        n10827), .Y(\i_MIPS/N117 ) );
  OAI221X4 U3474 ( .A0(net112366), .A1(\i_MIPS/n369 ), .B0(net112348), .B1(
        \i_MIPS/n368 ), .C0(n6769), .Y(n7815) );
  AO22X4 U3475 ( .A0(n3838), .A1(n9169), .B0(net100583), .B1(n9168), .Y(n9171)
         );
  INVX20 U3476 ( .A(n9469), .Y(n9328) );
  AND4X6 U3477 ( .A(n3929), .B(net133411), .C(net103923), .D(net105600), .Y(
        net128301) );
  XOR2X4 U3478 ( .A(n10344), .B(n10357), .Y(n10345) );
  NAND2X4 U3479 ( .A(n3690), .B(n8627), .Y(n10151) );
  INVX12 U3480 ( .A(n4620), .Y(n3697) );
  OAI221X2 U3481 ( .A0(n8428), .A1(net111622), .B0(n8427), .B1(net111634), 
        .C0(n8426), .Y(n9979) );
  INVX16 U3482 ( .A(n5546), .Y(n4153) );
  INVXL U3483 ( .A(n3737), .Y(n3677) );
  INVX3 U3484 ( .A(n10077), .Y(n10071) );
  NAND4BX4 U3485 ( .AN(n3820), .B(n3705), .C(net105783), .D(net127933), .Y(
        net105777) );
  OR2X8 U3486 ( .A(n10333), .B(n10334), .Y(n3678) );
  OR2X1 U3487 ( .A(n10448), .B(net112404), .Y(n3679) );
  OR2X8 U3488 ( .A(n10331), .B(n10335), .Y(n3680) );
  INVX3 U3489 ( .A(n10456), .Y(n10448) );
  BUFX4 U3490 ( .A(n5224), .Y(n5218) );
  NAND3BX2 U3491 ( .AN(n3858), .B(n4377), .C(n10359), .Y(\i_MIPS/PC/n62 ) );
  AOI21X2 U3492 ( .A0(n9274), .A1(n2210), .B0(n9140), .Y(n8536) );
  NAND2BX4 U3493 ( .AN(n10541), .B(n10540), .Y(n11120) );
  CLKBUFX2 U3494 ( .A(n5179), .Y(n5158) );
  OR2X4 U3495 ( .A(n4987), .B(n2206), .Y(n4183) );
  BUFX16 U3496 ( .A(n4990), .Y(n4987) );
  NAND4X6 U3497 ( .A(n6396), .B(n6395), .C(n6394), .D(n6393), .Y(n11497) );
  NAND2X6 U3498 ( .A(n9153), .B(n6753), .Y(n7468) );
  NOR3X6 U3499 ( .A(n3765), .B(n3766), .C(n3767), .Y(n7321) );
  INVX12 U3500 ( .A(net112438), .Y(net101082) );
  OA22X2 U3501 ( .A0(n10497), .A1(n4245), .B0(n10500), .B1(n4246), .Y(n9092)
         );
  NAND3X6 U3502 ( .A(n3795), .B(n3796), .C(net103251), .Y(n4135) );
  OA22XL U3503 ( .A0(\i_MIPS/Control_ID/n15 ), .A1(net112406), .B0(n220), .B1(
        n5625), .Y(n9970) );
  NAND2X2 U3504 ( .A(\i_MIPS/n295 ), .B(n5625), .Y(n4181) );
  NAND4X8 U3505 ( .A(n6372), .B(n6371), .C(n6370), .D(n6369), .Y(n11488) );
  BUFX3 U3506 ( .A(n5174), .Y(n5161) );
  AOI222X4 U3507 ( .A0(n5500), .A1(n11437), .B0(mem_rdata_D[87]), .B1(n236), 
        .C0(n12964), .C1(n4385), .Y(n10944) );
  INVX12 U3508 ( .A(n1953), .Y(mem_wdata_D[32]) );
  OR3X8 U3509 ( .A(n4412), .B(n7873), .C(n6537), .Y(n3683) );
  INVX3 U3510 ( .A(n7511), .Y(n7873) );
  INVX3 U3511 ( .A(n4381), .Y(n6537) );
  NAND3X6 U3512 ( .A(n6354), .B(n6356), .C(n3410), .Y(n11503) );
  NAND2X4 U3513 ( .A(n5547), .B(n11345), .Y(n10076) );
  AO22X1 U3514 ( .A0(DCACHE_addr[25]), .A1(n4637), .B0(n5551), .B1(n11503), 
        .Y(n12791) );
  OA22X2 U3515 ( .A0(n10514), .A1(n4245), .B0(n10517), .B1(n4246), .Y(n8802)
         );
  OA22X4 U3516 ( .A0(n10842), .A1(net133585), .B0(n10841), .B1(net108658), .Y(
        n10843) );
  BUFX4 U3517 ( .A(n4891), .Y(n4935) );
  OA22X4 U3518 ( .A0(n10534), .A1(net133585), .B0(n10533), .B1(net108660), .Y(
        n10535) );
  INVX12 U3519 ( .A(net133585), .Y(n3897) );
  NOR2X6 U3520 ( .A(n7), .B(n4379), .Y(net105787) );
  NAND4X6 U3521 ( .A(n10039), .B(n10038), .C(n10037), .D(n10036), .Y(n10591)
         );
  OA22X1 U3522 ( .A0(n237), .A1(n1638), .B0(n5346), .B1(n3220), .Y(n10022) );
  AO21XL U3523 ( .A0(n3720), .A1(n10315), .B0(n10314), .Y(n10317) );
  AO21X2 U3524 ( .A0(net98385), .A1(net98386), .B0(net111904), .Y(net98531) );
  NAND2XL U3525 ( .A(net98371), .B(net98372), .Y(n10718) );
  OAI221XL U3526 ( .A0(net104407), .A1(net111624), .B0(net104408), .B1(
        net111636), .C0(net104409), .Y(n4614) );
  AND2XL U3527 ( .A(net98571), .B(net98572), .Y(n4403) );
  AO21X2 U3528 ( .A0(net98390), .A1(net98391), .B0(net111904), .Y(net98598) );
  AND2XL U3529 ( .A(net98530), .B(net98531), .Y(n4400) );
  CLKINVX1 U3530 ( .A(n7709), .Y(n3684) );
  AND2X6 U3531 ( .A(n11163), .B(n11162), .Y(n4435) );
  NAND4X2 U3532 ( .A(n10199), .B(n10198), .C(n10197), .D(n10196), .Y(n11221)
         );
  CLKINVX1 U3533 ( .A(n6606), .Y(n9884) );
  NAND3X2 U3534 ( .A(n9356), .B(net111994), .C(n9351), .Y(n9359) );
  NAND2X2 U3535 ( .A(n6542), .B(\i_MIPS/n367 ), .Y(n6963) );
  MXI2X4 U3536 ( .A(\i_MIPS/ID_EX[50] ), .B(n4662), .S0(n5624), .Y(n3687) );
  MXI2X4 U3537 ( .A(\i_MIPS/ID_EX[50] ), .B(n4662), .S0(n5624), .Y(n6529) );
  OAI222X2 U3538 ( .A0(n9245), .A1(n8457), .B0(n9342), .B1(n8456), .C0(n9455), 
        .C1(n8455), .Y(n8458) );
  NAND2X2 U3539 ( .A(n6548), .B(\i_MIPS/n349 ), .Y(n9476) );
  CLKMX2X8 U3540 ( .A(\i_MIPS/n265 ), .B(n4375), .S0(n5624), .Y(n6548) );
  NAND2X4 U3541 ( .A(n6541), .B(\i_MIPS/n368 ), .Y(n8360) );
  AND4X8 U3542 ( .A(net133414), .B(\i_MIPS/n333 ), .C(\i_MIPS/n331 ), .D(n3704), .Y(\i_MIPS/ALU_Control/n11 ) );
  OAI221X1 U3543 ( .A0(net112304), .A1(n8634), .B0(n7052), .B1(net101257), 
        .C0(net112420), .Y(n7056) );
  OAI221X1 U3544 ( .A0(net112304), .A1(n7878), .B0(n6971), .B1(net101257), 
        .C0(net112420), .Y(n6974) );
  OAI2BB1X4 U3545 ( .A0N(n8996), .A1N(n8995), .B0(n3690), .Y(n10281) );
  INVX3 U3546 ( .A(n8159), .Y(n7704) );
  NAND2X1 U3547 ( .A(net107808), .B(n4536), .Y(n8649) );
  INVX16 U3548 ( .A(\i_MIPS/ID_EX[80] ), .Y(net102253) );
  INVX12 U3549 ( .A(net112338), .Y(net112334) );
  AO22X2 U3550 ( .A0(n7413), .A1(net137952), .B0(net112296), .B1(n7685), .Y(
        n7415) );
  AO21X2 U3551 ( .A0(n7021), .A1(n7020), .B0(n5546), .Y(net112799) );
  CLKBUFX2 U3552 ( .A(n7683), .Y(n3688) );
  NAND2X8 U3553 ( .A(n6533), .B(\i_MIPS/ALUin1[5] ), .Y(n6966) );
  AND3X8 U3554 ( .A(n9066), .B(n8939), .C(n6519), .Y(n6524) );
  MXI2X4 U3555 ( .A(n10723), .B(n10722), .S0(n5518), .Y(n10724) );
  OA22X2 U3556 ( .A0(n10673), .A1(n4245), .B0(n10676), .B1(n4246), .Y(n9196)
         );
  OAI221X2 U3557 ( .A0(n9481), .A1(n8538), .B0(n7800), .B1(n7799), .C0(n8071), 
        .Y(n7811) );
  OA22X2 U3558 ( .A0(n5130), .A1(n740), .B0(n5069), .B1(n2301), .Y(n6003) );
  NAND2X4 U3559 ( .A(n6009), .B(n6008), .Y(n6010) );
  CLKBUFX6 U3560 ( .A(net97418), .Y(net108198) );
  NOR2BX4 U3561 ( .AN(net112338), .B(\i_MIPS/n340 ), .Y(n4519) );
  OAI2BB1X4 U3562 ( .A0N(n6531), .A1N(\i_MIPS/n363 ), .B0(n8641), .Y(n6507) );
  AOI2BB1X1 U3563 ( .A0N(n3676), .A1N(n10445), .B0(n10444), .Y(n10447) );
  AOI2BB1X2 U3564 ( .A0N(n3676), .A1N(n3889), .B0(n10323), .Y(n10252) );
  AND3X8 U3565 ( .A(net133411), .B(net103924), .C(net105600), .Y(n3731) );
  AND2X8 U3566 ( .A(net103907), .B(net103924), .Y(n4394) );
  INVX12 U3567 ( .A(n3929), .Y(net103924) );
  NAND4X2 U3568 ( .A(n6130), .B(n6129), .C(n6128), .D(n6127), .Y(n11286) );
  NOR4X4 U3569 ( .A(n7026), .B(n7025), .C(n7024), .D(n7023), .Y(n7027) );
  NAND2X2 U3570 ( .A(n4522), .B(n4502), .Y(n9414) );
  INVX6 U3571 ( .A(n10839), .Y(n10836) );
  INVX4 U3572 ( .A(net112338), .Y(n3829) );
  INVX16 U3573 ( .A(net112338), .Y(net112336) );
  NAND4X2 U3574 ( .A(n7355), .B(n7354), .C(n7353), .D(n7352), .Y(n11360) );
  NOR2X6 U3575 ( .A(n4219), .B(n10543), .Y(n10545) );
  NAND4X4 U3576 ( .A(n9913), .B(n9912), .C(n9911), .D(n9910), .Y(n11287) );
  NAND4X2 U3577 ( .A(n6730), .B(n6729), .C(n6728), .D(n6727), .Y(n6745) );
  NOR3X1 U3578 ( .A(n6726), .B(n6725), .C(n6724), .Y(n6727) );
  INVXL U3579 ( .A(n3412), .Y(n3689) );
  AOI2BB2X1 U3580 ( .B0(n11457), .B1(n3761), .A0N(n10710), .A1N(n4250), .Y(
        n7281) );
  NAND3BX2 U3581 ( .AN(n10555), .B(n10554), .C(n10553), .Y(\i_MIPS/PC/n56 ) );
  CLKINVX2 U3582 ( .A(n7707), .Y(n7615) );
  XNOR2X4 U3583 ( .A(\i_MIPS/ID_EX[106] ), .B(\i_MIPS/ID_EX[107] ), .Y(
        \i_MIPS/ALU_Control/n18 ) );
  AOI222X2 U3584 ( .A0(n3848), .A1(net101401), .B0(net101402), .B1(n8960), 
        .C0(n9058), .C1(n8959), .Y(n8961) );
  NAND2X6 U3585 ( .A(net98351), .B(net98352), .Y(n4092) );
  OA22X2 U3586 ( .A0(n10920), .A1(n4245), .B0(n10923), .B1(n4246), .Y(n8404)
         );
  BUFX6 U3587 ( .A(net97701), .Y(n3918) );
  OA22X2 U3588 ( .A0(n10984), .A1(n4245), .B0(n10987), .B1(n4246), .Y(n6815)
         );
  XOR2X4 U3589 ( .A(n4138), .B(n3693), .Y(n3925) );
  INVX4 U3590 ( .A(n4478), .Y(n4695) );
  NAND4X2 U3591 ( .A(n6235), .B(n6234), .C(n6233), .D(n6232), .Y(n11247) );
  OAI21X4 U3592 ( .A0(n8977), .A1(n8976), .B0(n8975), .Y(n3895) );
  NAND2X1 U3593 ( .A(n9064), .B(n9041), .Y(n8953) );
  MXI2X4 U3594 ( .A(n3695), .B(n3694), .S0(n5622), .Y(n6530) );
  INVX12 U3595 ( .A(n4671), .Y(n4670) );
  OA22X4 U3596 ( .A0(\i_MIPS/ALUin1[25] ), .A1(n4670), .B0(\i_MIPS/ALUin1[26] ), .B1(n3828), .Y(n6482) );
  OA22X2 U3597 ( .A0(\i_MIPS/ALUin1[26] ), .A1(n4670), .B0(\i_MIPS/ALUin1[27] ), .B1(n3828), .Y(n6681) );
  OR2X2 U3598 ( .A(n8640), .B(net101257), .Y(n4169) );
  AND2X2 U3599 ( .A(n5557), .B(n11232), .Y(n12890) );
  NAND4X2 U3600 ( .A(n9608), .B(n9607), .C(n9606), .D(n9605), .Y(n11232) );
  BUFX20 U3601 ( .A(n5549), .Y(n5548) );
  OAI22X1 U3602 ( .A0(n10940), .A1(n4675), .B0(n10943), .B1(n4250), .Y(n3700)
         );
  OAI22X1 U3603 ( .A0(n10946), .A1(n4245), .B0(n10949), .B1(n4246), .Y(n3701)
         );
  INVX6 U3604 ( .A(n5546), .Y(n3720) );
  AOI222X4 U3605 ( .A0(n5503), .A1(n11350), .B0(mem_rdata_D[0]), .B1(n232), 
        .C0(n12987), .C1(n5502), .Y(n10960) );
  NAND3X2 U3606 ( .A(n4220), .B(n4221), .C(n4222), .Y(n10398) );
  OR2X4 U3607 ( .A(n4403), .B(net108704), .Y(n4222) );
  BUFX16 U3608 ( .A(n3927), .Y(net108710) );
  OA22X2 U3609 ( .A0(n10508), .A1(n4675), .B0(n10511), .B1(n4250), .Y(n8803)
         );
  NAND2X4 U3610 ( .A(n4539), .B(n5623), .Y(n4318) );
  CLKMX2X6 U3611 ( .A(n7126), .B(n7125), .S0(net107812), .Y(net104582) );
  NAND4BX2 U3612 ( .AN(n7115), .B(n7114), .C(n7113), .D(n7112), .Y(n7126) );
  NOR4X2 U3613 ( .A(n7111), .B(n7110), .C(n7109), .D(n7108), .Y(n7112) );
  NAND3X6 U3614 ( .A(n3702), .B(n3703), .C(net102792), .Y(net98722) );
  CLKMX2X2 U3615 ( .A(n8129), .B(n8128), .S0(net107810), .Y(net102790) );
  AOI21X1 U3616 ( .A0(net102426), .A1(net102427), .B0(net102428), .Y(n4419) );
  NAND2X4 U3617 ( .A(\i_MIPS/ALUin1[4] ), .B(n6542), .Y(n7503) );
  AOI2BB2X1 U3618 ( .B0(n4248), .B1(\D_cache/cache[5][147] ), .A0N(n4926), 
        .A1N(n3320), .Y(n6429) );
  NAND2X8 U3619 ( .A(net111902), .B(net100682), .Y(net101978) );
  XOR2X1 U3620 ( .A(n6604), .B(\i_MIPS/IR_ID[24] ), .Y(n6452) );
  AO21X4 U3621 ( .A0(n10559), .A1(n10558), .B0(net111640), .Y(n8916) );
  NAND2X4 U3622 ( .A(n4504), .B(n4447), .Y(net102049) );
  BUFX4 U3623 ( .A(net100597), .Y(net112002) );
  NAND4BX2 U3624 ( .AN(n7124), .B(n7123), .C(n7122), .D(n7121), .Y(n7125) );
  OA22X1 U3625 ( .A0(\i_MIPS/Register/register[20][8] ), .A1(n4699), .B0(
        \i_MIPS/Register/register[28][8] ), .B1(n4695), .Y(n7123) );
  NOR4X4 U3626 ( .A(n7120), .B(n7119), .C(n7118), .D(n7117), .Y(n7121) );
  AO22X1 U3627 ( .A0(n9531), .A1(n983), .B0(n4715), .B1(n2499), .Y(n7119) );
  OAI222X2 U3628 ( .A0(n7043), .A1(n7303), .B0(n7042), .B1(n7301), .C0(
        net101914), .C1(n8258), .Y(n7067) );
  OR2X4 U3629 ( .A(net102404), .B(net107796), .Y(n7301) );
  AO21X4 U3630 ( .A0(n6658), .A1(n6657), .B0(n3697), .Y(n10136) );
  OAI221X2 U3631 ( .A0(net104230), .A1(n8353), .B0(n4662), .B1(n6978), .C0(
        n8350), .Y(n9462) );
  CLKBUFX4 U3632 ( .A(n4934), .Y(n4902) );
  AO22X1 U3633 ( .A0(net108200), .A1(n9893), .B0(n202), .B1(n3704), .Y(
        \i_MIPS/n472 ) );
  NOR3X2 U3634 ( .A(n4173), .B(n4174), .C(n4175), .Y(n3706) );
  OAI2BB1X4 U3635 ( .A0N(net97496), .A1N(n10627), .B0(n3707), .Y(n10323) );
  BUFX8 U3636 ( .A(n9989), .Y(n4954) );
  INVX4 U3637 ( .A(n10862), .Y(n3756) );
  AOI22X1 U3638 ( .A0(n12939), .A1(n11510), .B0(n5551), .B1(n11496), .Y(n3708)
         );
  MXI2X2 U3639 ( .A(n10699), .B(n10698), .S0(n5517), .Y(n10700) );
  AOI211X2 U3640 ( .A0(n3838), .A1(n9251), .B0(n6855), .C0(n6854), .Y(n6856)
         );
  AND2X8 U3641 ( .A(n4484), .B(net112292), .Y(n4310) );
  MXI2X2 U3642 ( .A(n10897), .B(n10896), .S0(n5520), .Y(n10898) );
  AOI222X4 U3643 ( .A0(n5499), .A1(n11422), .B0(mem_rdata_D[72]), .B1(n233), 
        .C0(n12979), .C1(n5497), .Y(n10897) );
  CLKBUFX3 U3644 ( .A(n5033), .Y(n5017) );
  AND2X2 U3645 ( .A(net101910), .B(n3764), .Y(n4173) );
  BUFX6 U3646 ( .A(n10653), .Y(n3909) );
  NAND2BX1 U3647 ( .AN(n4649), .B(n11425), .Y(n3711) );
  AO22X4 U3648 ( .A0(n8640), .A1(net137952), .B0(net112296), .B1(n8639), .Y(
        n8644) );
  OA21X4 U3649 ( .A0(n9463), .A1(n8258), .B0(n8257), .Y(n3821) );
  OA22X1 U3650 ( .A0(n4970), .A1(n1081), .B0(n5015), .B1(n2674), .Y(n8892) );
  OAI211X2 U3651 ( .A0(n6969), .A1(n6968), .B0(n7502), .C0(n7509), .Y(n6970)
         );
  MX2X1 U3652 ( .A(net112415), .B(net101082), .S0(n3634), .Y(n7235) );
  NAND2X4 U3653 ( .A(n9243), .B(n9144), .Y(n9477) );
  OA22X1 U3654 ( .A0(n3716), .A1(n3804), .B0(n4649), .B1(n3815), .Y(n3715) );
  CLKINVX3 U3655 ( .A(n4637), .Y(n3804) );
  MXI2X4 U3656 ( .A(\i_MIPS/ID_EX[64] ), .B(\i_MIPS/ID_EX[96] ), .S0(n3801), 
        .Y(n6566) );
  NAND2X2 U3657 ( .A(n6978), .B(n9164), .Y(n4225) );
  NAND2X8 U3658 ( .A(n7822), .B(n6771), .Y(n9463) );
  INVX8 U3659 ( .A(n6753), .Y(n6771) );
  NAND2X2 U3660 ( .A(n4570), .B(n8534), .Y(n9274) );
  AOI2BB2XL U3661 ( .B0(net111962), .B1(n3738), .A0N(n3773), .A1N(net104252), 
        .Y(n3722) );
  INVX1 U3662 ( .A(n3824), .Y(n7406) );
  NAND2X2 U3663 ( .A(\i_MIPS/IR_ID[22] ), .B(\i_MIPS/n231 ), .Y(n6457) );
  XOR2X1 U3664 ( .A(n6606), .B(\i_MIPS/IR_ID[22] ), .Y(n6447) );
  AND2X4 U3665 ( .A(n402), .B(n4499), .Y(net128155) );
  NAND2BX1 U3666 ( .AN(n4649), .B(n11427), .Y(n3723) );
  NAND2BX1 U3667 ( .AN(n4649), .B(n11431), .Y(n3724) );
  CLKBUFX2 U3668 ( .A(n9991), .Y(n4999) );
  NAND2X8 U3669 ( .A(\i_MIPS/ALUin1[12] ), .B(n6561), .Y(n7683) );
  INVX4 U3670 ( .A(n9461), .Y(n3838) );
  AO22X2 U3671 ( .A0(net103548), .A1(n3726), .B0(n6850), .B1(net101908), .Y(
        n3725) );
  NAND2X6 U3672 ( .A(n4443), .B(n7468), .Y(net102404) );
  CLKINVX12 U3673 ( .A(net102404), .Y(net101908) );
  INVX2 U3674 ( .A(n7689), .Y(n7413) );
  NAND2X6 U3675 ( .A(\i_MIPS/n285 ), .B(n4316), .Y(n4317) );
  NAND2BX1 U3676 ( .AN(n4649), .B(n11433), .Y(n3727) );
  BUFX6 U3677 ( .A(n10193), .Y(n5224) );
  OA22X2 U3678 ( .A0(n5213), .A1(n1448), .B0(n5172), .B1(n3019), .Y(n10189) );
  NAND2BX1 U3679 ( .AN(n4649), .B(n11437), .Y(n3728) );
  NAND2BX2 U3680 ( .AN(net97798), .B(n4092), .Y(n4130) );
  INVX8 U3681 ( .A(n11432), .Y(n10511) );
  NAND4X4 U3682 ( .A(n8793), .B(n8792), .C(n8791), .D(n8790), .Y(n11432) );
  OA22X2 U3683 ( .A0(n4971), .A1(n678), .B0(n5016), .B1(n2249), .Y(n8790) );
  INVX12 U3684 ( .A(n6542), .Y(n6532) );
  CLKBUFX2 U3685 ( .A(n5309), .Y(n5285) );
  AOI2BB1X4 U3686 ( .A0N(n10339), .A1N(n10572), .B0(n10575), .Y(n10341) );
  INVX12 U3687 ( .A(net112306), .Y(net112292) );
  AOI21X2 U3688 ( .A0(n10451), .A1(net98487), .B0(n10450), .Y(n10452) );
  OA22X2 U3689 ( .A0(n5374), .A1(n1462), .B0(n5345), .B1(n3036), .Y(n9962) );
  NAND2BX4 U3690 ( .AN(n10447), .B(n10446), .Y(net98487) );
  INVX8 U3691 ( .A(n3842), .Y(net133411) );
  MXI2X2 U3692 ( .A(n10918), .B(n10917), .S0(n5521), .Y(n10919) );
  AOI222X4 U3693 ( .A0(n5500), .A1(n11417), .B0(mem_rdata_D[67]), .B1(n234), 
        .C0(n12984), .C1(n4385), .Y(n10918) );
  AO21X4 U3694 ( .A0(n10287), .A1(n10286), .B0(net111902), .Y(net98708) );
  OAI2BB1X4 U3695 ( .A0N(n10287), .A1N(n10286), .B0(net112782), .Y(net102792)
         );
  OR2X4 U3696 ( .A(n6640), .B(net111636), .Y(n4187) );
  NAND2X6 U3697 ( .A(n3420), .B(n4139), .Y(n4103) );
  AO21X4 U3698 ( .A0(net99002), .A1(net99003), .B0(net111644), .Y(net104889)
         );
  NOR4X2 U3699 ( .A(n7859), .B(n7858), .C(n7857), .D(n7856), .Y(n7860) );
  OA22X1 U3700 ( .A0(n4631), .A1(n3804), .B0(n4649), .B1(n3733), .Y(n3732) );
  NAND2BX4 U3701 ( .AN(net112764), .B(n3839), .Y(n3734) );
  BUFX20 U3702 ( .A(net127710), .Y(net112356) );
  AND3X8 U3703 ( .A(net133411), .B(net103923), .C(n4395), .Y(n3735) );
  INVX16 U3704 ( .A(n9455), .Y(n9165) );
  INVX8 U3705 ( .A(n9336), .Y(n9058) );
  NOR2X6 U3706 ( .A(n9455), .B(n3849), .Y(n3848) );
  OAI2BB1X4 U3707 ( .A0N(n8026), .A1N(n8025), .B0(n4153), .Y(n10525) );
  NAND4X2 U3708 ( .A(n6200), .B(n6199), .C(n6198), .D(n6197), .Y(n11312) );
  BUFX16 U3709 ( .A(n5090), .Y(n5133) );
  OA22XL U3710 ( .A0(n5198), .A1(n1578), .B0(n5155), .B1(n3160), .Y(n6199) );
  AND2X8 U3711 ( .A(n3839), .B(net102253), .Y(net128151) );
  INVX20 U3712 ( .A(net112338), .Y(n3828) );
  XNOR2X4 U3713 ( .A(n8918), .B(n3736), .Y(n3957) );
  NAND3X6 U3714 ( .A(n4176), .B(n4177), .C(n8916), .Y(n3736) );
  AO22XL U3715 ( .A0(n4298), .A1(net137952), .B0(net112296), .B1(n4498), .Y(
        n7980) );
  AO22X1 U3716 ( .A0(n4713), .A1(n279), .B0(n4708), .B1(n2500), .Y(n7868) );
  AO22X2 U3717 ( .A0(n4722), .A1(n642), .B0(n4719), .B1(n2217), .Y(n7866) );
  INVX2 U3718 ( .A(n7469), .Y(n7042) );
  OAI221X4 U3719 ( .A0(net112366), .A1(\i_MIPS/n352 ), .B0(net112348), .B1(
        \i_MIPS/n353 ), .C0(n6853), .Y(n7469) );
  AOI2BB2X4 U3720 ( .B0(net111960), .B1(n3738), .A0N(n3773), .A1N(net104252), 
        .Y(n3772) );
  NAND4X2 U3721 ( .A(n8986), .B(n8985), .C(n8984), .D(n8983), .Y(n11440) );
  MX2XL U3722 ( .A(DCACHE_addr[9]), .B(net112999), .S0(n214), .Y(\i_MIPS/n458 ) );
  MX2XL U3723 ( .A(DCACHE_addr[6]), .B(net97817), .S0(n222), .Y(\i_MIPS/n461 )
         );
  AOI2BB2X2 U3724 ( .B0(n11446), .B1(n3761), .A0N(n10956), .A1N(n4250), .Y(
        n7590) );
  NAND4X2 U3725 ( .A(n7576), .B(n7575), .C(n7574), .D(n7573), .Y(n11446) );
  NAND2X8 U3726 ( .A(n6532), .B(\i_MIPS/n367 ), .Y(n7509) );
  MXI2X2 U3727 ( .A(n10756), .B(n10755), .S0(n5519), .Y(n10757) );
  OAI221XL U3728 ( .A0(net103581), .A1(net111624), .B0(net103582), .B1(
        net111636), .C0(net103583), .Y(n3741) );
  INVX16 U3729 ( .A(net101914), .Y(net103548) );
  OA22X4 U3730 ( .A0(n4669), .A1(\i_MIPS/n344 ), .B0(net112330), .B1(
        \i_MIPS/n345 ), .Y(n6918) );
  OA22X4 U3731 ( .A0(n4669), .A1(n7696), .B0(n3828), .B1(\i_MIPS/n364 ), .Y(
        n6686) );
  NAND2X6 U3732 ( .A(net101908), .B(net107796), .Y(n7303) );
  AND3X2 U3733 ( .A(n8860), .B(n8871), .C(net137952), .Y(n8880) );
  OR2X1 U3734 ( .A(n4649), .B(n10684), .Y(n3744) );
  OR2X1 U3735 ( .A(n4649), .B(n10494), .Y(n3743) );
  NAND4X2 U3736 ( .A(n9083), .B(n9082), .C(n9081), .D(n9080), .Y(n11439) );
  NAND4X2 U3737 ( .A(n4356), .B(n8194), .C(n8193), .D(n8192), .Y(n11443) );
  INVX1 U3738 ( .A(n11443), .Y(n10684) );
  AO21X4 U3739 ( .A0(n6897), .A1(n6896), .B0(n3729), .Y(net99165) );
  MXI2X2 U3740 ( .A(n10685), .B(n10684), .S0(n5517), .Y(n10686) );
  NAND2X4 U3741 ( .A(n6612), .B(n4501), .Y(n9524) );
  CLKBUFX8 U3742 ( .A(n4677), .Y(n4679) );
  NAND2BX4 U3743 ( .AN(n5425), .B(n11257), .Y(n10134) );
  XOR3XL U3744 ( .A(n10227), .B(n4390), .C(n10236), .Y(n10586) );
  OAI2BB2X2 U3745 ( .B0(\i_MIPS/n179 ), .B1(net108192), .A0N(n4315), .A1N(
        n10354), .Y(\i_MIPS/N119 ) );
  CLKINVX12 U3746 ( .A(n6457), .Y(n6458) );
  BUFX4 U3747 ( .A(net112138), .Y(net112132) );
  OA22X2 U3748 ( .A0(n10269), .A1(n4675), .B0(n10272), .B1(n4250), .Y(n8996)
         );
  OR2X1 U3749 ( .A(n4649), .B(n10956), .Y(n3883) );
  OR2X1 U3750 ( .A(n4649), .B(n10871), .Y(n3873) );
  OR2X1 U3751 ( .A(n4649), .B(n10478), .Y(n3868) );
  NAND2BX1 U3752 ( .AN(n4649), .B(n11452), .Y(n3876) );
  NAND2BX1 U3753 ( .AN(n4649), .B(n11411), .Y(n3877) );
  NAND2BX1 U3754 ( .AN(n4649), .B(n11449), .Y(n3881) );
  OR2X1 U3755 ( .A(n4649), .B(n10978), .Y(n3880) );
  OR2X1 U3756 ( .A(n4649), .B(n10278), .Y(n3870) );
  OR2X1 U3757 ( .A(n4649), .B(n10887), .Y(n3867) );
  OR2X1 U3758 ( .A(n4649), .B(n10736), .Y(n3882) );
  OR2X1 U3759 ( .A(n4649), .B(n10750), .Y(n3874) );
  OR2X1 U3760 ( .A(n4649), .B(n10902), .Y(n3871) );
  OR2X1 U3761 ( .A(n4649), .B(n10758), .Y(n3878) );
  OR2X1 U3762 ( .A(n4649), .B(n10713), .Y(n3872) );
  OR2X1 U3763 ( .A(n4649), .B(n10953), .Y(n3869) );
  OR2X1 U3764 ( .A(n4649), .B(n10763), .Y(n4607) );
  AOI22X1 U3765 ( .A0(DCACHE_addr[13]), .A1(n11510), .B0(n4653), .B1(n11491), 
        .Y(n4636) );
  INVXL U3766 ( .A(n3845), .Y(n3846) );
  INVX4 U3767 ( .A(n10150), .Y(n3845) );
  NAND4X4 U3768 ( .A(n6023), .B(n6022), .C(n6021), .D(n6020), .Y(n11324) );
  OA22X4 U3769 ( .A0(n5379), .A1(n2101), .B0(n5326), .B1(n516), .Y(n6020) );
  BUFX4 U3770 ( .A(n5533), .Y(n5541) );
  XNOR2X2 U3771 ( .A(ICACHE_addr[9]), .B(n11324), .Y(n6029) );
  AOI222X2 U3772 ( .A0(n7980), .A1(n7979), .B0(n4459), .B1(net101908), .C0(
        net101402), .C1(n9059), .Y(n7986) );
  OR2X8 U3773 ( .A(n8167), .B(n7707), .Y(n4147) );
  BUFX12 U3774 ( .A(net127709), .Y(net112374) );
  OAI222X2 U3775 ( .A0(n9247), .A1(n9469), .B0(n9463), .B1(n8443), .C0(n8442), 
        .C1(net133688), .Y(n8446) );
  NAND2X1 U3776 ( .A(net112374), .B(\i_MIPS/n354 ), .Y(n8251) );
  BUFX4 U3777 ( .A(n4837), .Y(n4826) );
  CLKAND2X12 U3778 ( .A(n4303), .B(n9974), .Y(n3745) );
  AND2X4 U3779 ( .A(n4620), .B(n8), .Y(n4303) );
  CLKINVX1 U3780 ( .A(DCACHE_ren), .Y(n9974) );
  INVX4 U3781 ( .A(n10965), .Y(n8427) );
  OA21X4 U3782 ( .A0(n4670), .A1(\i_MIPS/n352 ), .B0(n6920), .Y(n6921) );
  NAND3X8 U3783 ( .A(n11348), .B(n3854), .C(n11349), .Y(n11480) );
  OA22X2 U3784 ( .A0(n10758), .A1(n4245), .B0(n10761), .B1(n4246), .Y(n7198)
         );
  INVX3 U3785 ( .A(n7807), .Y(n7809) );
  AO22X2 U3786 ( .A0(net100583), .A1(n8560), .B0(n9276), .B1(net100585), .Y(
        n8559) );
  AO22X4 U3787 ( .A0(net100583), .A1(n7820), .B0(n7819), .B1(net100585), .Y(
        n7829) );
  MXI2X4 U3788 ( .A(n10714), .B(n10713), .S0(n5517), .Y(n10715) );
  INVX8 U3789 ( .A(n7609), .Y(n7520) );
  OA22X2 U3790 ( .A0(n4917), .A1(n652), .B0(n4249), .B1(n2228), .Y(n8600) );
  OAI221X2 U3791 ( .A0(net112366), .A1(\i_MIPS/n361 ), .B0(net112348), .B1(
        \i_MIPS/n360 ), .C0(n7699), .Y(n9158) );
  BUFX3 U3792 ( .A(n9533), .Y(n4723) );
  NAND2X2 U3793 ( .A(n8237), .B(n8851), .Y(n3746) );
  NAND3X8 U3794 ( .A(n6565), .B(n8244), .C(n3747), .Y(n6583) );
  INVX1 U3795 ( .A(n6841), .Y(n6843) );
  MX2XL U3796 ( .A(\i_MIPS/ID_EX[73] ), .B(\i_MIPS/Sign_Extend_ID[0] ), .S0(
        n208), .Y(\i_MIPS/n512 ) );
  OAI221X4 U3797 ( .A0(\i_MIPS/Register/register[18][13] ), .A1(net112076), 
        .B0(\i_MIPS/Register/register[26][13] ), .B1(net112090), .C0(n7731), 
        .Y(n7734) );
  NAND4X2 U3798 ( .A(n6170), .B(n6169), .C(n6168), .D(n6167), .Y(n11214) );
  OA22X2 U3799 ( .A0(n5106), .A1(n3016), .B0(n5088), .B1(n722), .Y(n6170) );
  NAND4X1 U3800 ( .A(n10351), .B(n10350), .C(n10349), .D(n10348), .Y(n10374)
         );
  OAI2BB1X4 U3801 ( .A0N(n8405), .A1N(n8404), .B0(n4153), .Y(n9977) );
  NAND4X2 U3802 ( .A(n9385), .B(n9384), .C(n9383), .D(n9382), .Y(n11473) );
  AOI222X4 U3803 ( .A0(n5504), .A1(n11375), .B0(mem_rdata_D[25]), .B1(n232), 
        .C0(n12962), .C1(n5501), .Y(n10498) );
  AO21X2 U3804 ( .A0(n9978), .A1(n9977), .B0(net111902), .Y(n10926) );
  OAI2BB2XL U3805 ( .B0(\i_MIPS/n218 ), .B1(net108194), .A0N(n4315), .A1N(
        n11173), .Y(\i_MIPS/N61 ) );
  XOR3X1 U3806 ( .A(net112400), .B(n10437), .C(n10621), .Y(n10440) );
  NAND2X2 U3807 ( .A(n11161), .B(n11173), .Y(n11090) );
  OA22X1 U3808 ( .A0(n5124), .A1(n1639), .B0(n5070), .B1(n3221), .Y(n10199) );
  AOI222XL U3809 ( .A0(n5510), .A1(n11400), .B0(mem_rdata_D[50]), .B1(n233), 
        .C0(n12969), .C1(n5506), .Y(n10518) );
  INVX8 U3810 ( .A(n11400), .Y(n10517) );
  OA22X2 U3811 ( .A0(n4970), .A1(n661), .B0(n5015), .B1(n2250), .Y(n8798) );
  OA22X4 U3812 ( .A0(n10288), .A1(n4676), .B0(n10291), .B1(n4250), .Y(n8109)
         );
  NAND4X8 U3813 ( .A(n6384), .B(n6383), .C(n6382), .D(n6381), .Y(n11493) );
  NAND3X2 U3814 ( .A(n10082), .B(n10085), .C(n10084), .Y(n11002) );
  AOI222X4 U3815 ( .A0(n5510), .A1(n11410), .B0(mem_rdata_D[60]), .B1(n235), 
        .C0(n12959), .C1(n5506), .Y(n10485) );
  BUFX4 U3816 ( .A(n4421), .Y(n5506) );
  AOI2BB1X4 U3817 ( .A0N(net112304), .A1N(n8076), .B0(net100583), .Y(n8082) );
  OAI2BB1X4 U3818 ( .A0N(n7755), .A1N(n7756), .B0(n4153), .Y(n10521) );
  XNOR2X4 U3819 ( .A(n9019), .B(n4592), .Y(n3748) );
  XOR2X4 U3820 ( .A(n3797), .B(n10490), .Y(n3749) );
  XNOR2X4 U3821 ( .A(n9221), .B(n225), .Y(n3750) );
  XNOR2X4 U3822 ( .A(n9326), .B(n3909), .Y(n3751) );
  NAND3BX2 U3823 ( .AN(n3752), .B(n3793), .C(n3794), .Y(n11166) );
  NOR2X2 U3824 ( .A(\i_MIPS/PC/n7 ), .B(net108686), .Y(n3752) );
  CLKBUFX6 U3825 ( .A(n5036), .Y(n5028) );
  NAND4X4 U3826 ( .A(n8797), .B(n8796), .C(n8795), .D(n8794), .Y(n11368) );
  OA22X1 U3827 ( .A0(n4745), .A1(n2952), .B0(n4789), .B1(n1139), .Y(n8797) );
  OA22X2 U3828 ( .A0(n4971), .A1(n679), .B0(n5016), .B1(n2251), .Y(n8794) );
  OA22X4 U3829 ( .A0(n4986), .A1(n2102), .B0(n5032), .B1(n517), .Y(n6419) );
  AOI2BB2X4 U3830 ( .B0(n4508), .B1(\D_cache/cache[1][145] ), .A0N(n4762), 
        .A1N(n2019), .Y(n6422) );
  OA22X4 U3831 ( .A0(n4763), .A1(n2103), .B0(n4795), .B1(n518), .Y(n6396) );
  OA22X2 U3832 ( .A0(n5295), .A1(n1449), .B0(n5248), .B1(n3020), .Y(n9655) );
  BUFX8 U3833 ( .A(n5264), .Y(n5248) );
  NAND4X6 U3834 ( .A(n9657), .B(n9656), .C(n9655), .D(n9654), .Y(n11233) );
  OA22X2 U3835 ( .A0(n5214), .A1(n1463), .B0(n5171), .B1(n3037), .Y(n10124) );
  OA22X1 U3836 ( .A0(n5211), .A1(n1640), .B0(n5168), .B1(n3222), .Y(n10010) );
  OA22X2 U3837 ( .A0(n5211), .A1(n1465), .B0(n5168), .B1(n3039), .Y(n10005) );
  AOI222X4 U3838 ( .A0(n5496), .A1(n11459), .B0(mem_rdata_D[109]), .B1(n232), 
        .C0(n12974), .C1(n5493), .Y(n10731) );
  NAND3X8 U3839 ( .A(n6298), .B(n4663), .C(n4665), .Y(n9987) );
  AOI222X4 U3840 ( .A0(n5498), .A1(n11439), .B0(mem_rdata_D[89]), .B1(n233), 
        .C0(n12962), .C1(n4385), .Y(n10495) );
  NAND3X6 U3841 ( .A(n3756), .B(n10861), .C(n10860), .Y(\i_MIPS/PC/n65 ) );
  NAND3X6 U3842 ( .A(net100396), .B(net100397), .C(n3917), .Y(n4528) );
  OR2X2 U3843 ( .A(n8337), .B(net111622), .Y(n3757) );
  OR2X6 U3844 ( .A(n8336), .B(net111634), .Y(n3758) );
  NAND3X6 U3845 ( .A(n3757), .B(n3758), .C(n8335), .Y(n10775) );
  CLKMX2X2 U3846 ( .A(n8334), .B(n8333), .S0(net107810), .Y(n8337) );
  NAND4X8 U3847 ( .A(n6114), .B(n6113), .C(n6112), .D(n6111), .Y(n9569) );
  NAND3XL U3848 ( .A(n4313), .B(n4314), .C(n9661), .Y(n3865) );
  NAND4X2 U3849 ( .A(n9697), .B(n9696), .C(n9695), .D(n9694), .Y(n11199) );
  NAND4X6 U3850 ( .A(n9712), .B(n9711), .C(n9710), .D(n9709), .Y(n10422) );
  BUFX16 U3851 ( .A(net127709), .Y(net112372) );
  NAND2X6 U3852 ( .A(\i_MIPS/ALUin1[7] ), .B(n4616), .Y(n7891) );
  OA22X2 U3853 ( .A0(n10752), .A1(n4676), .B0(n10755), .B1(n4250), .Y(n7199)
         );
  NAND2X6 U3854 ( .A(n4154), .B(n7405), .Y(n7410) );
  NAND2X6 U3855 ( .A(net103070), .B(net105034), .Y(n6755) );
  OR2X2 U3856 ( .A(net103089), .B(net111624), .Y(n3759) );
  OR2X4 U3857 ( .A(net103090), .B(net111634), .Y(n3760) );
  AOI2BB2X1 U3858 ( .B0(n11471), .B1(n3761), .A0N(n10494), .A1N(n4250), .Y(
        n9093) );
  NAND4X2 U3859 ( .A(n9079), .B(n9078), .C(n9077), .D(n9076), .Y(n11471) );
  NAND4X4 U3860 ( .A(n6416), .B(n6417), .C(n6418), .D(n6415), .Y(n11505) );
  INVXL U3861 ( .A(n4536), .Y(n3843) );
  INVX4 U3862 ( .A(n5626), .Y(n4299) );
  CLKMX2X12 U3863 ( .A(\i_MIPS/n247 ), .B(n4490), .S0(n4299), .Y(n6693) );
  AOI2BB1XL U3864 ( .A0N(\i_MIPS/ALUin1[16] ), .A1N(net112334), .B0(n4464), 
        .Y(n8067) );
  AOI2BB1X1 U3865 ( .A0N(\i_MIPS/ALUin1[16] ), .A1N(net112368), .B0(n4472), 
        .Y(n6683) );
  AND2XL U3866 ( .A(n7313), .B(net100585), .Y(n3765) );
  NOR2X6 U3867 ( .A(n3894), .B(n3895), .Y(n3893) );
  AOI2BB1X1 U3868 ( .A0N(n9455), .A1N(n9454), .B0(n9453), .Y(n9474) );
  AO22X1 U3869 ( .A0(n3848), .A1(n9059), .B0(n9058), .B1(n9057), .Y(n9060) );
  OA22X2 U3870 ( .A0(n8356), .A1(n3762), .B0(n8547), .B1(net102405), .Y(n8364)
         );
  AOI211X2 U3871 ( .A0(net101908), .A1(n7712), .B0(n6774), .C0(n6773), .Y(
        n6775) );
  INVXL U3872 ( .A(n11497), .Y(n3769) );
  OA22X2 U3873 ( .A0(n10701), .A1(n4245), .B0(n10704), .B1(n4246), .Y(n8700)
         );
  CLKINVX1 U3874 ( .A(n3634), .Y(n7405) );
  NAND4X2 U3875 ( .A(n6435), .B(n6434), .C(n6433), .D(n6432), .Y(n11504) );
  NAND2X2 U3876 ( .A(n6553), .B(\i_MIPS/n354 ), .Y(n3770) );
  NOR4X6 U3877 ( .A(n7530), .B(n7536), .C(n9478), .D(n7529), .Y(n7531) );
  INVX1 U3878 ( .A(n9137), .Y(n9478) );
  OAI222X2 U3879 ( .A0(n7314), .A1(n8353), .B0(net101401), .B1(net103552), 
        .C0(n4662), .C1(n9464), .Y(n7616) );
  NAND4X2 U3880 ( .A(n6220), .B(n6219), .C(n6218), .D(n6217), .Y(n11311) );
  NAND2X4 U3881 ( .A(n8737), .B(n8532), .Y(n9264) );
  NAND2XL U3882 ( .A(n3661), .B(n8736), .Y(n8745) );
  NAND2X2 U3883 ( .A(net128301), .B(n7822), .Y(n7901) );
  OA22XL U3884 ( .A0(\i_MIPS/Register/register[5][21] ), .A1(net112224), .B0(
        \i_MIPS/Register/register[13][21] ), .B1(net112240), .Y(n9119) );
  OA22XL U3885 ( .A0(\i_MIPS/Register/register[21][21] ), .A1(net112224), .B0(
        \i_MIPS/Register/register[29][21] ), .B1(net112244), .Y(n9128) );
  OA22XL U3886 ( .A0(\i_MIPS/Register/register[5][20] ), .A1(net112224), .B0(
        \i_MIPS/Register/register[13][20] ), .B1(net112244), .Y(n9224) );
  OA22XL U3887 ( .A0(\i_MIPS/Register/register[21][20] ), .A1(net112224), .B0(
        \i_MIPS/Register/register[29][20] ), .B1(net112240), .Y(n9233) );
  OA22X1 U3888 ( .A0(\i_MIPS/Register/register[21][27] ), .A1(net112224), .B0(
        \i_MIPS/Register/register[29][27] ), .B1(net112242), .Y(n9372) );
  OA22X1 U3889 ( .A0(\i_MIPS/Register/register[5][27] ), .A1(net112224), .B0(
        \i_MIPS/Register/register[13][27] ), .B1(net112236), .Y(n9363) );
  OR2X2 U3890 ( .A(n9116), .B(net111622), .Y(n3774) );
  INVX3 U3891 ( .A(n10487), .Y(n9115) );
  OA22X4 U3892 ( .A0(n4987), .A1(n2104), .B0(n5033), .B1(n519), .Y(n6377) );
  NAND2X6 U3893 ( .A(n3731), .B(net103913), .Y(net101413) );
  AO22X2 U3894 ( .A0(n9166), .A1(n9165), .B0(n9164), .B1(n9163), .Y(n9172) );
  OA22X2 U3895 ( .A0(n10667), .A1(n4675), .B0(n10670), .B1(n4250), .Y(n9197)
         );
  INVX4 U3896 ( .A(n10419), .Y(n10245) );
  AOI33X2 U3897 ( .A0(net112292), .A1(n8560), .A2(n8545), .B0(n8543), .B1(
        n8544), .B2(net137952), .Y(n8566) );
  INVX12 U3898 ( .A(n3847), .Y(net137951) );
  OA22XL U3899 ( .A0(\i_MIPS/Register/register[6][24] ), .A1(net112112), .B0(
        \i_MIPS/Register/register[14][24] ), .B1(net112132), .Y(n8280) );
  AND2X4 U3900 ( .A(n4521), .B(n4499), .Y(net128158) );
  OAI32X1 U3901 ( .A0(n8085), .A1(n7822), .A2(n8084), .B0(n7477), .B1(n7476), 
        .Y(n7487) );
  INVX1 U3902 ( .A(n7468), .Y(n8085) );
  OA22X2 U3903 ( .A0(n10660), .A1(n4245), .B0(n10663), .B1(n4246), .Y(n9302)
         );
  NOR2X8 U3904 ( .A(n6413), .B(n6414), .Y(n6426) );
  OA22X2 U3905 ( .A0(n4762), .A1(n3028), .B0(n4795), .B1(n846), .Y(n6412) );
  BUFX8 U3906 ( .A(n5041), .Y(n5032) );
  NAND2X4 U3907 ( .A(n3359), .B(n4506), .Y(n3916) );
  NAND2X8 U3908 ( .A(n7877), .B(n7902), .Y(n7403) );
  NAND2BX2 U3909 ( .AN(n4247), .B(n11295), .Y(n9712) );
  INVX12 U3910 ( .A(n6535), .Y(n6533) );
  AO22X2 U3911 ( .A0(n5528), .A1(DCACHE_addr[8]), .B0(n5527), .B1(n11486), .Y(
        n11037) );
  INVX3 U3912 ( .A(n9042), .Y(n8951) );
  NAND2X6 U3913 ( .A(\i_MIPS/ALUin1[25] ), .B(n6590), .Y(n9042) );
  NAND2X8 U3914 ( .A(n6551), .B(\i_MIPS/n355 ), .Y(n8072) );
  AOI2BB2X4 U3915 ( .B0(n3777), .B1(\D_cache/cache[6][139] ), .A0N(n5034), 
        .A1N(n3345), .Y(n6330) );
  OA22X4 U3916 ( .A0(n4924), .A1(n3367), .B0(n4950), .B1(n1738), .Y(n6420) );
  NAND4X2 U3917 ( .A(n6883), .B(n6882), .C(n6881), .D(n6880), .Y(n11450) );
  OAI221X2 U3918 ( .A0(net104864), .A1(net103060), .B0(n4084), .B1(net103076), 
        .C0(n4085), .Y(n4083) );
  INVX1 U3919 ( .A(n7887), .Y(n8863) );
  OAI211X2 U3920 ( .A0(n7538), .A1(n3661), .B0(n8532), .C0(n7537), .Y(n7540)
         );
  INVX3 U3921 ( .A(n7407), .Y(n6512) );
  OR2X2 U3922 ( .A(\i_MIPS/PC/n14 ), .B(net108686), .Y(n4220) );
  OAI21X4 U3923 ( .A0(n7167), .A1(n7166), .B0(n7165), .Y(n7168) );
  AND2X2 U3924 ( .A(n4502), .B(n4448), .Y(n4482) );
  INVX4 U3925 ( .A(n4482), .Y(n4701) );
  OAI221X2 U3926 ( .A0(net102937), .A1(net111624), .B0(net102938), .B1(
        net111634), .C0(net102939), .Y(n3780) );
  AO21X2 U3927 ( .A0(n10565), .A1(n10564), .B0(net111902), .Y(n10530) );
  NAND2X8 U3928 ( .A(n6533), .B(\i_MIPS/n366 ), .Y(n7502) );
  CLKMX2X3 U3929 ( .A(n8626), .B(n8625), .S0(net107810), .Y(n8629) );
  BUFX20 U3930 ( .A(n4140), .Y(net108670) );
  MXI2X2 U3931 ( .A(n10671), .B(n10670), .S0(n5516), .Y(n10672) );
  AOI222X4 U3932 ( .A0(n5498), .A1(n11435), .B0(mem_rdata_D[85]), .B1(n233), 
        .C0(n12966), .C1(n4385), .Y(n10671) );
  OAI221X2 U3933 ( .A0(net102937), .A1(net111624), .B0(net102938), .B1(
        net111634), .C0(net102939), .Y(net97798) );
  OA22X2 U3934 ( .A0(n4909), .A1(n653), .B0(n4947), .B1(n2230), .Y(n9193) );
  AOI222X4 U3935 ( .A0(n5505), .A1(n11358), .B0(mem_rdata_D[8]), .B1(n236), 
        .C0(n12979), .C1(n5502), .Y(n10900) );
  AOI222X4 U3936 ( .A0(n5505), .A1(n11364), .B0(mem_rdata_D[14]), .B1(n234), 
        .C0(n12973), .C1(n5502), .Y(n10748) );
  OA22X2 U3937 ( .A0(n10654), .A1(n4675), .B0(n10657), .B1(n4250), .Y(n9303)
         );
  AOI2BB2X2 U3938 ( .B0(\i_MIPS/IF_ID[75] ), .B1(n3930), .A0N(net108676), 
        .A1N(\i_MIPS/n193 ), .Y(n10820) );
  AOI2BB2X2 U3939 ( .B0(\i_MIPS/IF_ID[65] ), .B1(net108670), .A0N(net108674), 
        .A1N(\i_MIPS/n183 ), .Y(n10523) );
  AOI2BB2X2 U3940 ( .B0(\i_MIPS/IF_ID[70] ), .B1(n3930), .A0N(net108678), 
        .A1N(\i_MIPS/n188 ), .Y(n11165) );
  BUFX20 U3941 ( .A(net97416), .Y(net112406) );
  CLKINVX1 U3942 ( .A(n3781), .Y(n3782) );
  NAND2BX4 U3943 ( .AN(n5427), .B(n11187), .Y(n9967) );
  BUFX20 U3944 ( .A(n4884), .Y(n4881) );
  MXI2X2 U3945 ( .A(n10737), .B(n10736), .S0(n5518), .Y(n10738) );
  AOI222X4 U3946 ( .A0(n5505), .A1(n11363), .B0(mem_rdata_D[13]), .B1(n235), 
        .C0(n12974), .C1(n5502), .Y(n10737) );
  OA22X2 U3947 ( .A0(n5384), .A1(n1466), .B0(n5347), .B1(n3040), .Y(n10122) );
  INVX6 U3948 ( .A(net108680), .Y(net108678) );
  AND3X8 U3949 ( .A(n3652), .B(n10358), .C(net97592), .Y(n3927) );
  OA22X1 U3950 ( .A0(n4912), .A1(n1211), .B0(n4249), .B1(n2748), .Y(n8596) );
  OAI2BB2X1 U3951 ( .B0(\i_MIPS/n187 ), .B1(net108198), .A0N(n11108), .A1N(
        n4315), .Y(\i_MIPS/N30 ) );
  BUFX20 U3952 ( .A(n3915), .Y(n4315) );
  BUFX16 U3953 ( .A(n5036), .Y(n5035) );
  OAI2BB2X1 U3954 ( .B0(\i_MIPS/n232 ), .B1(net108198), .A0N(n4315), .A1N(
        n10457), .Y(\i_MIPS/N80 ) );
  AOI2BB2X2 U3955 ( .B0(n2016), .B1(net108664), .A0N(n11163), .A1N(net133585), 
        .Y(n11164) );
  OAI222X1 U3956 ( .A0(\i_MIPS/PC/n15 ), .A1(net108690), .B0(n3637), .B1(
        n10604), .C0(n4402), .C1(net108704), .Y(n10608) );
  NAND3BX4 U3957 ( .AN(n4143), .B(n4145), .C(n4144), .Y(\i_MIPS/PC/n57 ) );
  OAI2BB2X4 U3958 ( .B0(n3787), .B1(n3788), .A0N(net111966), .A1N(net98063), 
        .Y(net104042) );
  MXI2X2 U3959 ( .A(n7399), .B(n7398), .S0(net107816), .Y(n3788) );
  OR2X8 U3960 ( .A(n7543), .B(n7544), .Y(n3855) );
  AND2X4 U3961 ( .A(n3745), .B(n4460), .Y(n4421) );
  OA22X2 U3962 ( .A0(n11112), .A1(net133585), .B0(n11111), .B1(net108658), .Y(
        n11113) );
  OA22X2 U3963 ( .A0(n10587), .A1(net133585), .B0(n10586), .B1(net108660), .Y(
        n10588) );
  OA22X2 U3964 ( .A0(n10412), .A1(net133585), .B0(n10411), .B1(net108660), .Y(
        n10413) );
  NAND3BX2 U3965 ( .AN(n10537), .B(n10536), .C(n10535), .Y(\i_MIPS/PC/n54 ) );
  NAND3BX4 U3966 ( .AN(n3798), .B(net103923), .C(n6480), .Y(net100574) );
  OA22X4 U3967 ( .A0(n4918), .A1(n2105), .B0(n4948), .B1(n482), .Y(n7658) );
  OA22X4 U3968 ( .A0(n4918), .A1(n2107), .B0(n4948), .B1(n520), .Y(n7654) );
  AOI222X4 U3969 ( .A0(n5500), .A1(n11433), .B0(mem_rdata_D[83]), .B1(n236), 
        .C0(n4385), .C1(n12968), .Y(n10996) );
  AND2X2 U3970 ( .A(n232), .B(n11346), .Y(n4486) );
  AOI222X1 U3971 ( .A0(n5495), .A1(n11451), .B0(mem_rdata_D[101]), .B1(n236), 
        .C0(n12982), .C1(n5494), .Y(n10979) );
  AOI222X4 U3972 ( .A0(n5498), .A1(n11444), .B0(mem_rdata_D[94]), .B1(n232), 
        .C0(n12957), .C1(n4385), .Y(n10143) );
  MXI2X4 U3973 ( .A(n10143), .B(n10142), .S0(n5513), .Y(n10144) );
  OR2X6 U3974 ( .A(net104888), .B(net111636), .Y(n3790) );
  OA22X1 U3975 ( .A0(n8874), .A1(net102404), .B0(net137891), .B1(n7896), .Y(
        n7179) );
  NAND3BX4 U3976 ( .AN(n10430), .B(n10428), .C(n10429), .Y(\i_MIPS/PC/n49 ) );
  NOR4X4 U3977 ( .A(n7237), .B(n7238), .C(n7236), .D(n7235), .Y(n7239) );
  OA22X1 U3978 ( .A0(n4910), .A1(n1212), .B0(n4949), .B1(n2749), .Y(n9077) );
  INVX12 U3979 ( .A(n1955), .Y(mem_wdata_D[38]) );
  NAND3BX4 U3980 ( .AN(n10633), .B(n10632), .C(n10631), .Y(\i_MIPS/PC/n52 ) );
  OAI222X1 U3981 ( .A0(\i_MIPS/PC/n20 ), .A1(net108690), .B0(n3637), .B1(
        n10627), .C0(n4399), .C1(net108702), .Y(n10633) );
  AOI222X4 U3982 ( .A0(n5504), .A1(n11360), .B0(mem_rdata_D[10]), .B1(n236), 
        .C0(n12977), .C1(n5501), .Y(n10264) );
  INVX12 U3983 ( .A(n1957), .Y(mem_wdata_D[44]) );
  NOR4X1 U3984 ( .A(\i_MIPS/PHT_2/n12 ), .B(\i_MIPS/PHT_2/n13 ), .C(net112406), 
        .D(net97592), .Y(n11050) );
  MXI2X4 U3985 ( .A(n10668), .B(n10667), .S0(n5516), .Y(n10669) );
  AOI222X2 U3986 ( .A0(\i_MIPS/IF_ID[96] ), .A1(net108670), .B0(
        \i_MIPS/IF_ID_31 ), .B1(net108682), .C0(net108710), .C1(n3808), .Y(
        n10860) );
  INVX4 U3987 ( .A(n8456), .Y(n8250) );
  NAND4X4 U3988 ( .A(n6155), .B(n6154), .C(n6153), .D(n6152), .Y(n11218) );
  AOI2BB2X2 U3989 ( .B0(n10394), .B1(n3897), .A0N(n10395), .A1N(net108660), 
        .Y(n10396) );
  CLKMX2X4 U3990 ( .A(\i_MIPS/PHT_2/history_state[0] ), .B(n11044), .S0(n11045), .Y(\i_MIPS/PHT_2/n52 ) );
  XOR2X2 U3991 ( .A(\i_MIPS/IF_ID[64] ), .B(net112691), .Y(n11044) );
  OR2X1 U3992 ( .A(net97445), .B(n11162), .Y(n3793) );
  OR2X4 U3993 ( .A(n4407), .B(net108704), .Y(n3794) );
  NAND2BX2 U3994 ( .AN(n4247), .B(n11285), .Y(n10203) );
  CLKMX2X6 U3995 ( .A(n260), .B(n7470), .S0(net107796), .Y(n6850) );
  CLKMX2X4 U3996 ( .A(n7470), .B(n4587), .S0(net107794), .Y(n7060) );
  OAI221X4 U3997 ( .A0(n4669), .A1(\i_MIPS/n346 ), .B0(net112334), .B1(
        \i_MIPS/n347 ), .C0(n6838), .Y(n7470) );
  OA22X2 U3998 ( .A0(n4817), .A1(n662), .B0(n4863), .B1(n2231), .Y(n8800) );
  MX2X1 U3999 ( .A(net101082), .B(net112415), .S0(n7684), .Y(n7419) );
  NAND2X1 U4000 ( .A(\i_MIPS/ALUin1[13] ), .B(net128151), .Y(n7698) );
  INVX8 U4001 ( .A(n3892), .Y(n9990) );
  OR2X2 U4002 ( .A(net103249), .B(net111624), .Y(n3795) );
  OR2X4 U4003 ( .A(net103250), .B(net111636), .Y(n3796) );
  CLKMX2X4 U4004 ( .A(net103252), .B(net103253), .S0(net107812), .Y(net103249)
         );
  XNOR2X4 U4005 ( .A(n3845), .B(n11176), .Y(net105349) );
  BUFX8 U4006 ( .A(n4332), .Y(n4774) );
  AOI222X1 U4007 ( .A0(n5505), .A1(n11359), .B0(mem_rdata_D[9]), .B1(n236), 
        .C0(n12978), .C1(n5502), .Y(n10702) );
  BUFX6 U4008 ( .A(n4840), .Y(n4816) );
  OA22X1 U4009 ( .A0(n7489), .A1(net103076), .B0(net103060), .B1(n7488), .Y(
        n7549) );
  OAI222X2 U4010 ( .A0(n9247), .A1(n9461), .B0(n9463), .B1(n9246), .C0(n9245), 
        .C1(n9459), .Y(n9260) );
  AND2X8 U4011 ( .A(n10467), .B(n10466), .Y(n3797) );
  OA22X4 U4012 ( .A0(n4669), .A1(\i_MIPS/n350 ), .B0(net112334), .B1(
        \i_MIPS/n351 ), .Y(n6837) );
  NAND2X2 U4013 ( .A(n6594), .B(n3358), .Y(n8166) );
  INVX16 U4014 ( .A(n4323), .Y(n5625) );
  BUFX20 U4015 ( .A(n4990), .Y(n4986) );
  NOR2X6 U4016 ( .A(n3713), .B(n11497), .Y(n3816) );
  OA22X4 U4017 ( .A0(n4835), .A1(n2109), .B0(n4880), .B1(n522), .Y(n6395) );
  INVX20 U4018 ( .A(net112370), .Y(net112368) );
  AOI2BB1X2 U4019 ( .A0N(net112368), .A1N(\i_MIPS/n344 ), .B0(n4510), .Y(n6838) );
  OAI221X2 U4020 ( .A0(net112368), .A1(\i_MIPS/n364 ), .B0(net112350), .B1(
        \i_MIPS/n363 ), .C0(n6486), .Y(n7315) );
  INVX4 U4021 ( .A(n9057), .Y(n8658) );
  INVX4 U4022 ( .A(n3844), .Y(n7814) );
  AOI2BB1X4 U4023 ( .A0N(net112368), .A1N(n7149), .B0(n4511), .Y(n6752) );
  AOI211X2 U4024 ( .A0(n10245), .A1(n10244), .B0(n10432), .C0(n10416), .Y(
        n10246) );
  OAI221X2 U4025 ( .A0(n8353), .A1(n8650), .B0(n4662), .B1(n9163), .C0(n8350), 
        .Y(n9151) );
  NAND4X6 U4026 ( .A(n7746), .B(n7745), .C(n7744), .D(n7743), .Y(n11427) );
  OA22X4 U4027 ( .A0(n4978), .A1(n2110), .B0(n5023), .B1(n523), .Y(n7743) );
  INVX8 U4028 ( .A(n11427), .Y(n10733) );
  NAND2X2 U4029 ( .A(\i_MIPS/ID_EX[88] ), .B(n5622), .Y(n4165) );
  OR2X4 U4030 ( .A(n4904), .B(n3014), .Y(n4155) );
  NOR2X4 U4031 ( .A(n3822), .B(n8254), .Y(n8256) );
  NAND3BX4 U4032 ( .AN(\i_MIPS/n340 ), .B(n6771), .C(\i_MIPS/ID_EX[83] ), .Y(
        n9339) );
  BUFX12 U4033 ( .A(n8533), .Y(n4570) );
  AND2X8 U4034 ( .A(n4178), .B(n4179), .Y(n3799) );
  OA22X4 U4035 ( .A0(n4835), .A1(n511), .B0(n4880), .B1(n2098), .Y(n3800) );
  OAI222X2 U4036 ( .A0(n8353), .A1(n7317), .B0(n4660), .B1(n7300), .C0(n6976), 
        .C1(n4659), .Y(net105012) );
  AOI2BB2X2 U4037 ( .B0(\i_MIPS/IF_ID[83] ), .B1(net108670), .A0N(net108676), 
        .A1N(\i_MIPS/n201 ), .Y(n10632) );
  NAND2X8 U4038 ( .A(n10363), .B(n10366), .Y(n10205) );
  NAND2X8 U4039 ( .A(n10802), .B(n10800), .Y(n10366) );
  INVXL U4040 ( .A(n9569), .Y(n4059) );
  OAI31X2 U4041 ( .A0(n6525), .A1(n6524), .A2(n6523), .B0(n6522), .Y(n8431) );
  MX2X1 U4042 ( .A(net101082), .B(net112415), .S0(n6964), .Y(n6773) );
  OR4X4 U4043 ( .A(\i_MIPS/ID_EX[73] ), .B(n3696), .C(\i_MIPS/ID_EX[77] ), .D(
        n3704), .Y(net127702) );
  AOI211X2 U4044 ( .A0(n7508), .A1(net102426), .B0(n7507), .C0(n7506), .Y(
        n7513) );
  AO21X4 U4045 ( .A0(n11184), .A1(n11183), .B0(n11182), .Y(n11546) );
  INVX4 U4046 ( .A(n8150), .Y(n11182) );
  NAND4X4 U4047 ( .A(n7428), .B(n7427), .C(n7426), .D(n7425), .Y(n11458) );
  OA22X1 U4048 ( .A0(n4824), .A1(n1213), .B0(n4869), .B1(n2750), .Y(n7941) );
  AOI222X4 U4049 ( .A0(n5496), .A1(n11463), .B0(mem_rdata_D[113]), .B1(n235), 
        .C0(n12970), .C1(n5493), .Y(n10764) );
  BUFX12 U4050 ( .A(n4383), .Y(n5493) );
  AOI222X4 U4051 ( .A0(n5498), .A1(n11442), .B0(mem_rdata_D[92]), .B1(n235), 
        .C0(n12959), .C1(n4385), .Y(n10479) );
  BUFX12 U4052 ( .A(n11510), .Y(mem_read_D) );
  INVX1 U4053 ( .A(n11479), .Y(n11009) );
  INVXL U4054 ( .A(net97444), .Y(net138001) );
  AND3X6 U4055 ( .A(n3926), .B(n3652), .C(n4223), .Y(net129024) );
  OA22X4 U4056 ( .A0(n4762), .A1(n2112), .B0(n4795), .B1(n525), .Y(n3805) );
  OA22X4 U4057 ( .A0(n4835), .A1(n2113), .B0(n4880), .B1(n526), .Y(n3806) );
  INVXL U4058 ( .A(net102791), .Y(n3807) );
  CLKBUFX3 U4059 ( .A(n4382), .Y(n4665) );
  NAND2BX2 U4060 ( .AN(n4247), .B(n11293), .Y(n9760) );
  OAI221X1 U4061 ( .A0(\i_MIPS/Register/register[2][27] ), .A1(net112078), 
        .B0(\i_MIPS/Register/register[10][27] ), .B1(net112100), .C0(n9365), 
        .Y(n9368) );
  CLKBUFX2 U4062 ( .A(n10880), .Y(n3808) );
  CLKAND2X12 U4063 ( .A(net103910), .B(n3798), .Y(n4395) );
  MXI2X2 U4064 ( .A(n10921), .B(n10920), .S0(n5521), .Y(n10922) );
  AOI222X4 U4065 ( .A0(n5503), .A1(n11353), .B0(mem_rdata_D[3]), .B1(n233), 
        .C0(n12984), .C1(n5502), .Y(n10921) );
  NAND2X6 U4066 ( .A(n6589), .B(n7149), .Y(n11181) );
  BUFX20 U4067 ( .A(n4800), .Y(n4795) );
  CLKMX2X4 U4068 ( .A(\i_MIPS/n313 ), .B(n4537), .S0(\i_MIPS/ID_EX_5 ), .Y(
        n6605) );
  MXI2X2 U4069 ( .A(\i_MIPS/ID_EX[115] ), .B(\i_MIPS/ID_EX[88] ), .S0(
        \i_MIPS/ID_EX_5 ), .Y(n9882) );
  NAND3BX4 U4070 ( .AN(n3783), .B(n4661), .C(n224), .Y(n10193) );
  INVXL U4071 ( .A(n3405), .Y(n3809) );
  OA22X1 U4072 ( .A0(n4826), .A1(n2953), .B0(n4871), .B1(n1290), .Y(n7655) );
  MX2X2 U4073 ( .A(n7796), .B(n7795), .S0(net107816), .Y(n7836) );
  AO22XL U4074 ( .A0(net112036), .A1(n888), .B0(net100603), .B1(n2582), .Y(
        n8145) );
  AO22XL U4075 ( .A0(net112036), .A1(n866), .B0(net100603), .B1(n2548), .Y(
        n8136) );
  AO22XL U4076 ( .A0(net112036), .A1(n889), .B0(net100603), .B1(n2583), .Y(
        n7925) );
  AO22XL U4077 ( .A0(net112036), .A1(n890), .B0(net100603), .B1(n2584), .Y(
        n7733) );
  AO22XL U4078 ( .A0(net112036), .A1(n891), .B0(net100603), .B1(n2585), .Y(
        n8062) );
  XOR2X1 U4079 ( .A(n9885), .B(\i_MIPS/IR_ID[23] ), .Y(n6449) );
  OA21X4 U4080 ( .A0(net112368), .A1(n7696), .B0(n7695), .Y(n7697) );
  AO22X1 U4081 ( .A0(DCACHE_addr[9]), .A1(n11510), .B0(n4654), .B1(n11487), 
        .Y(n12795) );
  AOI2BB1X4 U4082 ( .A0N(n3828), .A1N(n7149), .B0(n4516), .Y(n6840) );
  NOR4X6 U4083 ( .A(n9063), .B(n9062), .C(n9061), .D(n9060), .Y(n9072) );
  INVXL U4084 ( .A(n7308), .Y(n7313) );
  AND2X4 U4085 ( .A(\i_MIPS/ALUin1[25] ), .B(net112372), .Y(n4512) );
  BUFX2 U4086 ( .A(n5313), .Y(n5306) );
  AOI22X1 U4087 ( .A0(DCACHE_addr[22]), .A1(n11510), .B0(n5551), .B1(n11500), 
        .Y(n3810) );
  OR2X4 U4088 ( .A(n10385), .B(n10237), .Y(n10400) );
  OA22X2 U4089 ( .A0(n5285), .A1(n750), .B0(n5258), .B1(n2311), .Y(n10099) );
  AOI22X1 U4090 ( .A0(n12946), .A1(n11510), .B0(n4653), .B1(n11489), .Y(n3811)
         );
  NAND3BX2 U4091 ( .AN(n4661), .B(n3784), .C(n224), .Y(n10192) );
  INVX8 U4092 ( .A(net105777), .Y(n4080) );
  OAI221X2 U4093 ( .A0(net112304), .A1(n7306), .B0(n7307), .B1(net101257), 
        .C0(net112420), .Y(n7311) );
  AOI211X2 U4094 ( .A0(n7874), .A1(n7519), .B0(n7518), .C0(n7517), .Y(n7534)
         );
  OAI22X1 U4095 ( .A0(n4758), .A1(n648), .B0(n4788), .B1(n2225), .Y(n4341) );
  NAND2X4 U4096 ( .A(n6535), .B(\i_MIPS/n366 ), .Y(n6964) );
  OA22X2 U4097 ( .A0(n10818), .A1(net133585), .B0(n10817), .B1(net108658), .Y(
        n10819) );
  CLKINVX2 U4098 ( .A(n10812), .Y(n10818) );
  AO22X2 U4099 ( .A0(n4723), .A1(n417), .B0(n4719), .B1(n2001), .Y(n8618) );
  OAI211XL U4100 ( .A0(\i_MIPS/ID_EX[80] ), .A1(n8358), .B0(n7695), .C0(n6767), 
        .Y(n6768) );
  AO22X4 U4101 ( .A0(n4722), .A1(n456), .B0(n4719), .B1(n2042), .Y(n7951) );
  AO22X4 U4102 ( .A0(n4722), .A1(n457), .B0(n4719), .B1(n2043), .Y(n7857) );
  CLKINVX8 U4103 ( .A(net101552), .Y(net98499) );
  NAND3X6 U4104 ( .A(n7798), .B(n8071), .C(n7797), .Y(n6577) );
  NOR3X1 U4105 ( .A(n6739), .B(n6738), .C(n6737), .Y(n6740) );
  AOI221X2 U4106 ( .A0(net137952), .A1(n7691), .B0(n7690), .B1(net112292), 
        .C0(net100583), .Y(n7715) );
  AOI222XL U4107 ( .A0(n5510), .A1(n11402), .B0(mem_rdata_D[52]), .B1(n235), 
        .C0(n12967), .C1(n5506), .Y(n10664) );
  INVX8 U4108 ( .A(n11402), .Y(n10663) );
  OA22X2 U4109 ( .A0(n4909), .A1(n655), .B0(n4947), .B1(n2232), .Y(n9300) );
  OAI2BB1X4 U4110 ( .A0N(n3667), .A1N(n6512), .B0(n6504), .Y(n6513) );
  NAND3BX1 U4111 ( .AN(n9352), .B(net112294), .C(n3899), .Y(n9358) );
  AOI221X1 U4112 ( .A0(n4450), .A1(n7540), .B0(n7539), .B1(n9137), .C0(n9482), 
        .Y(n7542) );
  OAI221X2 U4113 ( .A0(n8356), .A1(net137891), .B0(n9334), .B1(n9249), .C0(
        n7233), .Y(n7237) );
  OA22XL U4114 ( .A0(n8652), .A1(n9249), .B0(n9053), .B1(net101914), .Y(n8661)
         );
  NAND2X6 U4115 ( .A(net97936), .B(net97937), .Y(n4093) );
  CLKINVX8 U4116 ( .A(net103177), .Y(net97936) );
  NAND3BX4 U4117 ( .AN(n6969), .B(n4420), .C(n4388), .Y(n3814) );
  INVXL U4118 ( .A(n11498), .Y(n3815) );
  INVX1 U4119 ( .A(n11437), .Y(n10943) );
  OAI221X2 U4120 ( .A0(net104230), .A1(n4660), .B0(n4659), .B1(n7317), .C0(
        n8648), .Y(n8964) );
  OAI221X4 U4121 ( .A0(n3358), .A1(net112364), .B0(net112348), .B1(n7149), 
        .C0(n6918), .Y(n7317) );
  OA22X1 U4122 ( .A0(\i_MIPS/Register/register[22][2] ), .A1(n4684), .B0(
        \i_MIPS/Register/register[30][2] ), .B1(n4680), .Y(n6951) );
  OR2X4 U4123 ( .A(n5033), .B(n2207), .Y(n4184) );
  NAND2X6 U4124 ( .A(n11017), .B(n3415), .Y(n4336) );
  NAND2XL U4125 ( .A(n3415), .B(n11017), .Y(n11507) );
  AOI222X4 U4126 ( .A0(n5496), .A1(n11460), .B0(mem_rdata_D[110]), .B1(n233), 
        .C0(n12973), .C1(n5493), .Y(n10742) );
  MXI2X2 U4127 ( .A(\i_MIPS/ID_EX[68] ), .B(\i_MIPS/ID_EX[100] ), .S0(n5624), 
        .Y(n6592) );
  MXI2X2 U4128 ( .A(\i_MIPS/ID_EX[67] ), .B(\i_MIPS/ID_EX[99] ), .S0(n5622), 
        .Y(n6591) );
  CLKMX2X8 U4129 ( .A(\i_MIPS/n249 ), .B(n4492), .S0(n5622), .Y(n11180) );
  AOI222X2 U4130 ( .A0(n6771), .A1(\i_MIPS/ALU/N303 ), .B0(n9328), .B1(n6690), 
        .C0(n6689), .C1(n9165), .Y(n6691) );
  INVX3 U4131 ( .A(n7147), .Y(n6689) );
  OA22X4 U4132 ( .A0(n8353), .A1(n7899), .B0(n8864), .B1(n4659), .Y(n6688) );
  BUFX3 U4133 ( .A(net127709), .Y(net112376) );
  OAI211X1 U4134 ( .A0(n8453), .A1(n8179), .B0(n8166), .C0(n6526), .Y(n6527)
         );
  BUFX8 U4135 ( .A(n4334), .Y(n5180) );
  BUFX20 U4136 ( .A(n5041), .Y(n3840) );
  NAND2X4 U4137 ( .A(n6570), .B(\i_MIPS/n351 ), .Y(n9263) );
  NAND2X4 U4138 ( .A(n3713), .B(n11497), .Y(n4229) );
  NAND4X4 U4139 ( .A(n9905), .B(n9904), .C(n9903), .D(n9902), .Y(n11222) );
  OA22X1 U4140 ( .A0(n5375), .A1(n1641), .B0(n5347), .B1(n3223), .Y(n9902) );
  CLKINVX8 U4141 ( .A(n6511), .Y(n6504) );
  MX2X1 U4142 ( .A(net101082), .B(net112415), .S0(n7877), .Y(n6979) );
  NAND2BX4 U4143 ( .AN(n5425), .B(n11260), .Y(n10062) );
  NAND2BX1 U4144 ( .AN(n5427), .B(n11196), .Y(n10061) );
  NAND4X2 U4145 ( .A(n10053), .B(n10052), .C(n10051), .D(n10050), .Y(n11196)
         );
  OA22XL U4146 ( .A0(n4989), .A1(n1141), .B0(n5035), .B1(n2703), .Y(n6317) );
  OA22XL U4147 ( .A0(n4989), .A1(n1142), .B0(n5035), .B1(n2704), .Y(n6321) );
  BUFX3 U4148 ( .A(n4830), .Y(n4833) );
  NAND2BX4 U4149 ( .AN(net111640), .B(n6747), .Y(n6748) );
  NAND4X2 U4150 ( .A(n6644), .B(n6643), .C(n6642), .D(n6641), .Y(n11477) );
  OA22X2 U4151 ( .A0(n4833), .A1(n682), .B0(n4878), .B1(n2254), .Y(n6643) );
  BUFX2 U4152 ( .A(n4931), .Y(n4911) );
  OA22X2 U4153 ( .A0(n4911), .A1(n683), .B0(n4947), .B1(n2255), .Y(n8795) );
  NAND2X2 U4154 ( .A(\i_MIPS/ALUin1[20] ), .B(n6570), .Y(n9243) );
  OA22X4 U4155 ( .A0(n4669), .A1(net103561), .B0(n3829), .B1(\i_MIPS/n361 ), 
        .Y(n6486) );
  BUFX16 U4156 ( .A(n9991), .Y(n5041) );
  XNOR2X4 U4157 ( .A(n3817), .B(net99151), .Y(n4102) );
  NAND2X2 U4158 ( .A(n8957), .B(n8960), .Y(n6488) );
  OAI221X4 U4159 ( .A0(\i_MIPS/ALUin1[23] ), .A1(net112364), .B0(
        \i_MIPS/ALUin1[24] ), .B1(net112346), .C0(n6482), .Y(n6483) );
  XOR2X4 U4160 ( .A(n4336), .B(n3928), .Y(n3850) );
  OA22X4 U4161 ( .A0(n4484), .A1(net112306), .B0(net101257), .B1(n7225), .Y(
        n7242) );
  NAND2X8 U4162 ( .A(n7474), .B(n7982), .Y(n6916) );
  NAND2X2 U4163 ( .A(\i_MIPS/ALUin1[29] ), .B(n6585), .Y(n8165) );
  CLKMX2X3 U4164 ( .A(net101082), .B(net112415), .S0(n4483), .Y(n7903) );
  BUFX20 U4165 ( .A(n3735), .Y(net112415) );
  NAND2X4 U4166 ( .A(n6748), .B(n6750), .Y(n3818) );
  NAND2X2 U4167 ( .A(net111630), .B(n6746), .Y(n6750) );
  MX2X1 U4168 ( .A(n3610), .B(n10867), .S0(n213), .Y(\i_MIPS/n375 ) );
  INVXL U4169 ( .A(n7890), .Y(n7895) );
  OAI221X4 U4170 ( .A0(\i_MIPS/ALUin1[12] ), .A1(n4668), .B0(
        \i_MIPS/ALUin1[11] ), .B1(n3828), .C0(n7229), .Y(n7890) );
  OAI32X2 U4171 ( .A0(n8180), .A1(n8179), .A2(n8152), .B0(n8178), .B1(n8152), 
        .Y(n8171) );
  OA22X4 U4172 ( .A0(n10831), .A1(net133585), .B0(n10830), .B1(net108658), .Y(
        n10832) );
  NOR4X2 U4173 ( .A(n7485), .B(net103923), .C(n3798), .D(n7484), .Y(n7486) );
  INVX3 U4174 ( .A(n7976), .Y(n7977) );
  OAI221X4 U4175 ( .A0(\i_MIPS/ALUin1[12] ), .A1(net112364), .B0(
        \i_MIPS/ALUin1[11] ), .B1(net112346), .C0(n6754), .Y(n7978) );
  OA22X1 U4176 ( .A0(\i_MIPS/ALUin1[10] ), .A1(n4670), .B0(\i_MIPS/ALUin1[9] ), 
        .B1(n3828), .Y(n6754) );
  AO21X2 U4177 ( .A0(n9146), .A1(n9145), .B0(n9477), .Y(n9149) );
  INVX4 U4178 ( .A(n9477), .Y(n9479) );
  AO21X2 U4179 ( .A0(n4393), .A1(n9145), .B0(n8070), .Y(n8073) );
  AO22X4 U4180 ( .A0(n9328), .A1(n9332), .B0(n8552), .B1(n9327), .Y(n8557) );
  OA22X4 U4181 ( .A0(n4824), .A1(n2114), .B0(n4889), .B1(n527), .Y(n9505) );
  INVX8 U4182 ( .A(n7403), .Y(n7045) );
  NOR3X2 U4183 ( .A(net105783), .B(n3820), .C(n3704), .Y(n4081) );
  AND3X6 U4184 ( .A(n4295), .B(n4664), .C(n4666), .Y(n3892) );
  AO21X2 U4185 ( .A0(n8255), .A1(n8957), .B0(n9453), .Y(n3822) );
  OAI221X4 U4186 ( .A0(n4660), .A1(n4587), .B0(n4659), .B1(n7470), .C0(n8648), 
        .Y(n8258) );
  INVX4 U4187 ( .A(n9342), .Y(n8957) );
  INVX16 U4188 ( .A(n4658), .Y(n9453) );
  MX2X1 U4189 ( .A(net101082), .B(net112415), .S0(n8253), .Y(n8254) );
  NAND2X4 U4190 ( .A(n6574), .B(\i_MIPS/n353 ), .Y(n8730) );
  CLKINVX2 U4191 ( .A(n9140), .Y(n9273) );
  INVXL U4192 ( .A(n3798), .Y(n3823) );
  NOR4X4 U4193 ( .A(n8706), .B(n8705), .C(n8704), .D(n8703), .Y(n8707) );
  AO22X2 U4194 ( .A0(n4723), .A1(n638), .B0(n4719), .B1(n2213), .Y(n8704) );
  BUFX12 U4195 ( .A(n9530), .Y(n4714) );
  AOI211X1 U4196 ( .A0(n8157), .A1(net102253), .B0(n4513), .C0(n4511), .Y(
        n8158) );
  INVX3 U4197 ( .A(n8156), .Y(n8157) );
  NAND3X8 U4198 ( .A(n3825), .B(n3826), .C(n325), .Y(n3827) );
  NAND2X8 U4199 ( .A(n3827), .B(n9457), .Y(n6565) );
  CLKINVX12 U4200 ( .A(n9138), .Y(n9482) );
  NAND2X6 U4201 ( .A(\i_MIPS/ALUin1[22] ), .B(n6548), .Y(n9457) );
  MX2X2 U4202 ( .A(n9136), .B(n9135), .S0(\i_MIPS/IR_ID[25] ), .Y(n9179) );
  OA22XL U4203 ( .A0(\i_MIPS/Register/register[3][20] ), .A1(net112188), .B0(
        \i_MIPS/Register/register[11][20] ), .B1(n199), .Y(n9223) );
  OA22XL U4204 ( .A0(\i_MIPS/Register/register[19][20] ), .A1(net112182), .B0(
        \i_MIPS/Register/register[27][20] ), .B1(n197), .Y(n9232) );
  OA22X1 U4205 ( .A0(\i_MIPS/Register/register[19][21] ), .A1(net112182), .B0(
        \i_MIPS/Register/register[27][21] ), .B1(n198), .Y(n9127) );
  NAND2BX4 U4206 ( .AN(n4092), .B(n3780), .Y(n4131) );
  INVX6 U4207 ( .A(n7305), .Y(n7307) );
  OA22X4 U4208 ( .A0(n4835), .A1(n2121), .B0(n4880), .B1(n534), .Y(n6391) );
  OA22X4 U4209 ( .A0(n4987), .A1(n2122), .B0(n5033), .B1(n535), .Y(n6389) );
  OR2X6 U4210 ( .A(n6639), .B(net111624), .Y(n4188) );
  CLKMX2X2 U4211 ( .A(n6632), .B(n6631), .S0(net107812), .Y(n6639) );
  AO22X1 U4212 ( .A0(n4711), .A1(n424), .B0(n4707), .B1(n2003), .Y(n6617) );
  NAND2X6 U4213 ( .A(n10076), .B(n11346), .Y(n11479) );
  OA22X2 U4214 ( .A0(n4993), .A1(n751), .B0(n5034), .B1(n2312), .Y(n6339) );
  INVX3 U4215 ( .A(net112340), .Y(net112330) );
  NAND2X1 U4216 ( .A(n8339), .B(n7050), .Y(n6841) );
  NAND2X2 U4217 ( .A(\i_MIPS/ALUin1[11] ), .B(n6549), .Y(n7497) );
  NAND2BX4 U4218 ( .AN(n6755), .B(net105038), .Y(n6502) );
  NAND2X4 U4219 ( .A(\i_MIPS/ALUin1[21] ), .B(n6558), .Y(n9152) );
  NAND2BX4 U4220 ( .AN(n5429), .B(n11226), .Y(n10013) );
  AO22X4 U4221 ( .A0(mem_rdata_I[40]), .A1(n5537), .B0(n249), .B1(n11226), .Y(
        n10012) );
  NAND4BX2 U4222 ( .AN(n8513), .B(n8512), .C(n8511), .D(n8510), .Y(n8524) );
  AO22XL U4223 ( .A0(n9531), .A1(n322), .B0(n4714), .B1(n2549), .Y(n8327) );
  AO22XL U4224 ( .A0(n9531), .A1(n337), .B0(n4714), .B1(n2550), .Y(n8816) );
  AO22XL U4225 ( .A0(n9531), .A1(n352), .B0(n4714), .B1(n2586), .Y(n8418) );
  AO22XL U4226 ( .A0(n9531), .A1(n353), .B0(n4714), .B1(n2587), .Y(n8517) );
  AO22XL U4227 ( .A0(n9531), .A1(n354), .B0(n4714), .B1(n2588), .Y(n8409) );
  AO22XL U4228 ( .A0(n9531), .A1(n355), .B0(n4714), .B1(n2589), .Y(n8705) );
  NAND2X2 U4229 ( .A(n4522), .B(n4501), .Y(n9416) );
  AO22X4 U4230 ( .A0(n6710), .A1(net112294), .B0(n6709), .B1(net111992), .Y(
        n6711) );
  NAND4XL U4231 ( .A(n7501), .B(n7500), .C(n9456), .D(n7499), .Y(n7535) );
  NOR2BX4 U4232 ( .AN(n4527), .B(n4661), .Y(n4485) );
  AOI2BB1X4 U4233 ( .A0N(n6704), .A1N(net112306), .B0(n6597), .Y(n6601) );
  NAND3X6 U4234 ( .A(n4161), .B(n4162), .C(n7150), .Y(n8352) );
  OR2X2 U4235 ( .A(n3358), .B(net112346), .Y(n4162) );
  OAI2BB1X1 U4236 ( .A0N(n256), .A1N(n6708), .B0(n7481), .Y(n6702) );
  NAND2X4 U4237 ( .A(n6531), .B(\i_MIPS/n364 ), .Y(n7902) );
  NAND3BX2 U4238 ( .AN(n9430), .B(n3690), .C(net111910), .Y(n9399) );
  NAND3BX4 U4239 ( .AN(n8182), .B(net111994), .C(n264), .Y(n8183) );
  OA22X4 U4240 ( .A0(n4987), .A1(n2124), .B0(n5033), .B1(n537), .Y(n6397) );
  OR3X6 U4241 ( .A(net102554), .B(net102555), .C(net112304), .Y(net138213) );
  NAND2X8 U4242 ( .A(n7683), .B(n7409), .Y(n6510) );
  AO22X1 U4243 ( .A0(ICACHE_addr[17]), .A1(n11512), .B0(mem_write_I), .B1(
        n11332), .Y(n12816) );
  NAND2BX1 U4244 ( .AN(n5427), .B(n11190), .Y(n9907) );
  AOI22X1 U4245 ( .A0(DCACHE_addr[23]), .A1(n4637), .B0(n5551), .B1(n11501), 
        .Y(n3831) );
  AOI22X1 U4246 ( .A0(n12933), .A1(n11510), .B0(n5551), .B1(n11502), .Y(n3832)
         );
  OA22XL U4247 ( .A0(\i_MIPS/Register/register[22][4] ), .A1(n4684), .B0(
        \i_MIPS/Register/register[30][4] ), .B1(n4680), .Y(n6907) );
  AND2XL U4248 ( .A(net98363), .B(net98364), .Y(n4432) );
  CLKMX2X2 U4249 ( .A(net101082), .B(net112415), .S0(n8360), .Y(n8361) );
  OAI2BB2XL U4250 ( .B0(n9417), .B1(\i_MIPS/Register/register[7][25] ), .A0N(
        n4713), .A1N(n2443), .Y(n9098) );
  BUFX3 U4251 ( .A(n9528), .Y(n4710) );
  AOI31X1 U4252 ( .A0(n7495), .A1(\i_MIPS/n363 ), .A2(n8630), .B0(n7494), .Y(
        n7498) );
  AOI222X2 U4253 ( .A0(n5495), .A1(n11452), .B0(mem_rdata_D[102]), .B1(n233), 
        .C0(n12981), .C1(n5494), .Y(n10068) );
  XOR2X4 U4254 ( .A(n3918), .B(n3835), .Y(n3920) );
  INVX8 U4255 ( .A(n4298), .Y(n7474) );
  CLKINVX8 U4256 ( .A(n11233), .Y(n9659) );
  OAI221X2 U4257 ( .A0(n4668), .A1(\i_MIPS/n348 ), .B0(net112336), .B1(
        \i_MIPS/n349 ), .C0(n6919), .Y(n7300) );
  AOI2BB1X4 U4258 ( .A0N(net112350), .A1N(\i_MIPS/n347 ), .B0(n4512), .Y(n6919) );
  NOR4X6 U4259 ( .A(n7831), .B(n7830), .C(n7829), .D(n7828), .Y(n7832) );
  MX2X1 U4260 ( .A(net101082), .B(net112415), .S0(n9487), .Y(n9174) );
  MX2XL U4261 ( .A(n3612), .B(net99151), .S0(n216), .Y(\i_MIPS/n425 ) );
  OAI2BB2X4 U4262 ( .B0(n4163), .B1(n3836), .A0N(\i_MIPS/ID_EX[43] ), .A1N(
        n5625), .Y(net105677) );
  OA22X4 U4263 ( .A0(n5112), .A1(n2984), .B0(n5084), .B1(n1428), .Y(n9652) );
  NAND4X8 U4264 ( .A(n9652), .B(n9651), .C(n9650), .D(n9649), .Y(n11265) );
  BUFX3 U4265 ( .A(n5134), .Y(n5112) );
  NAND4X2 U4266 ( .A(n10043), .B(n10042), .C(n10041), .D(n10040), .Y(n11292)
         );
  AO22X2 U4267 ( .A0(n8550), .A1(n9054), .B0(n4471), .B1(n3838), .Y(n8558) );
  CLKINVX1 U4268 ( .A(n8547), .Y(n8550) );
  NAND2X4 U4269 ( .A(n4388), .B(n7159), .Y(n7412) );
  NAND3BX4 U4270 ( .AN(n8436), .B(net112294), .C(n9347), .Y(n8437) );
  INVX6 U4271 ( .A(n8437), .Y(n8448) );
  NAND4X4 U4272 ( .A(n8662), .B(n8661), .C(n8660), .D(n8659), .Y(n10693) );
  NAND4X4 U4273 ( .A(n7624), .B(n7623), .C(n7622), .D(n7621), .Y(net98029) );
  AOI222X2 U4274 ( .A0(n7615), .A1(net103710), .B0(n7614), .B1(n7613), .C0(
        n7612), .C1(n7611), .Y(n7624) );
  INVX4 U4275 ( .A(n8637), .Y(n7052) );
  INVX8 U4276 ( .A(n6965), .Y(n6500) );
  OAI221X4 U4277 ( .A0(net112306), .A1(n6759), .B0(n6760), .B1(net101257), 
        .C0(net112420), .Y(n6763) );
  BUFX20 U4278 ( .A(n4774), .Y(n4766) );
  OA22X4 U4279 ( .A0(n5203), .A1(n2985), .B0(n5159), .B1(n1429), .Y(n9651) );
  OA22XL U4280 ( .A0(n5203), .A1(n1848), .B0(n5159), .B1(n3504), .Y(n9681) );
  CLKBUFX6 U4281 ( .A(n5218), .Y(n5203) );
  NAND3X6 U4282 ( .A(ICACHE_addr[14]), .B(ICACHE_addr[13]), .C(n10239), .Y(
        n10248) );
  INVX6 U4283 ( .A(n10637), .Y(n10650) );
  OA22X4 U4284 ( .A0(n4764), .A1(n3368), .B0(n4796), .B1(n1739), .Y(n4329) );
  BUFX6 U4285 ( .A(n4335), .Y(n5356) );
  OA22X2 U4286 ( .A0(n5389), .A1(n1450), .B0(n5348), .B1(n3021), .Y(n10187) );
  AO22X2 U4287 ( .A0(n6971), .A1(net137952), .B0(net112296), .B1(n7878), .Y(
        n6973) );
  INVX20 U4288 ( .A(n4323), .Y(n5626) );
  BUFX20 U4289 ( .A(net100574), .Y(net112438) );
  CLKMX2X4 U4290 ( .A(net100573), .B(net112438), .S0(n8754), .Y(n7818) );
  CLKMX2X4 U4291 ( .A(net100573), .B(net112438), .S0(n8865), .Y(n8868) );
  OAI221X2 U4292 ( .A0(net112306), .A1(net102429), .B0(n4090), .B1(net101257), 
        .C0(net112420), .Y(n4087) );
  AO22X1 U4293 ( .A0(n4728), .A1(n984), .B0(n4725), .B1(n2501), .Y(n8206) );
  AND2X4 U4294 ( .A(n10427), .B(n10425), .Y(n4465) );
  INVX3 U4295 ( .A(n10611), .Y(n10617) );
  NAND2BX2 U4296 ( .AN(n5426), .B(n11264), .Y(n9612) );
  NAND2X6 U4297 ( .A(\i_MIPS/ALUin1[19] ), .B(n6554), .Y(n8546) );
  OA21X1 U4298 ( .A0(\i_MIPS/ALUin1[19] ), .A1(net112350), .B0(n8153), .Y(
        n8154) );
  OAI221X2 U4299 ( .A0(\i_MIPS/ALUin1[18] ), .A1(n4668), .B0(
        \i_MIPS/ALUin1[19] ), .B1(n3828), .C0(n6683), .Y(n8549) );
  OA22X2 U4300 ( .A0(n4913), .A1(n752), .B0(n4249), .B1(n2313), .Y(n8401) );
  NAND4X6 U4301 ( .A(n8403), .B(n8402), .C(n8401), .D(n8400), .Y(n11385) );
  NOR4X4 U4302 ( .A(n9202), .B(n9201), .C(n9200), .D(n9199), .Y(n9203) );
  AO22X1 U4303 ( .A0(n4713), .A1(n937), .B0(n4710), .B1(n2444), .Y(n9202) );
  CLKINVX20 U4304 ( .A(net137951), .Y(net101257) );
  NAND2X6 U4305 ( .A(n3731), .B(net103923), .Y(n3847) );
  OA22X4 U4306 ( .A0(n4669), .A1(\i_MIPS/n368 ), .B0(n3829), .B1(\i_MIPS/n367 ), .Y(n6849) );
  NOR4BX4 U4307 ( .AN(n9474), .B(n9473), .C(n9472), .D(n9471), .Y(n9498) );
  OAI222X4 U4308 ( .A0(n9463), .A1(n9462), .B0(n9461), .B1(n9460), .C0(
        net100581), .C1(n9459), .Y(n9472) );
  NAND4X2 U4309 ( .A(n8399), .B(n8398), .C(n8397), .D(n8396), .Y(n11353) );
  OA22X2 U4310 ( .A0(n4913), .A1(n753), .B0(n4249), .B1(n2314), .Y(n8397) );
  AO21X2 U4311 ( .A0(n4423), .A1(n9350), .B0(n9349), .Y(n9353) );
  NOR4X4 U4312 ( .A(n9308), .B(n9307), .C(n9306), .D(n9305), .Y(n9309) );
  NAND2BX2 U4313 ( .AN(n5426), .B(n11262), .Y(n9782) );
  NAND4BX4 U4314 ( .AN(n4345), .B(n9763), .C(n9762), .D(n9761), .Y(n11294) );
  OAI22X1 U4315 ( .A0(n5115), .A1(n647), .B0(n5064), .B1(n2223), .Y(n4345) );
  OA22X2 U4316 ( .A0(n5206), .A1(n3017), .B0(n5162), .B1(n723), .Y(n9763) );
  NAND4X2 U4317 ( .A(n7347), .B(n7346), .C(n7345), .D(n7344), .Y(n11456) );
  OA22X2 U4318 ( .A0(n4756), .A1(n754), .B0(n4793), .B1(n2315), .Y(n7347) );
  NAND3X6 U4319 ( .A(n3855), .B(n3856), .C(n8851), .Y(n7545) );
  AO22X1 U4320 ( .A0(n4712), .A1(n284), .B0(n4709), .B1(n2502), .Y(n8218) );
  OA22X4 U4321 ( .A0(n4755), .A1(n2203), .B0(n4793), .B1(n513), .Y(n7436) );
  MX2XL U4322 ( .A(\i_MIPS/ID_EX[75] ), .B(\i_MIPS/Sign_Extend_ID[2] ), .S0(
        n210), .Y(\i_MIPS/n510 ) );
  AND4X2 U4323 ( .A(n4080), .B(n3812), .C(net127930), .D(n3836), .Y(n3842) );
  OA22X1 U4324 ( .A0(n4836), .A1(n3215), .B0(n4882), .B1(n1291), .Y(n6341) );
  OAI222X4 U4325 ( .A0(n9337), .A1(n9336), .B0(net133688), .B1(n9335), .C0(
        n9334), .C1(n9333), .Y(n9344) );
  OAI222X4 U4326 ( .A0(n8874), .A1(n9467), .B0(n8873), .B1(n9461), .C0(n8872), 
        .C1(net112420), .Y(n8878) );
  NOR2BX4 U4327 ( .AN(\i_MIPS/IR_ID[21] ), .B(\i_MIPS/n232 ), .Y(n4521) );
  NAND4BX4 U4328 ( .AN(n4342), .B(n9512), .C(n9511), .D(n9510), .Y(n11404) );
  NAND2BX4 U4329 ( .AN(n5428), .B(n11197), .Y(n9758) );
  OA22XL U4330 ( .A0(n5205), .A1(n1143), .B0(n5161), .B1(n2738), .Y(n9740) );
  INVX8 U4331 ( .A(n9242), .Y(n7539) );
  NAND3X8 U4332 ( .A(n4376), .B(n6479), .C(\i_MIPS/ALU_Control/n20 ), .Y(
        net103923) );
  NAND4BX2 U4333 ( .AN(\i_MIPS/ID_EX[106] ), .B(\i_MIPS/ID_EX[105] ), .C(
        \i_MIPS/ID_EX[107] ), .D(\i_MIPS/ALU_Control/n11 ), .Y(
        \i_MIPS/ALU_Control/n20 ) );
  AO22X4 U4334 ( .A0(n4713), .A1(n304), .B0(n4710), .B1(n2021), .Y(n9107) );
  NAND2X8 U4335 ( .A(n4317), .B(n4318), .Y(n6550) );
  CLKINVX6 U4336 ( .A(n11106), .Y(n11112) );
  NAND2BX2 U4337 ( .AN(n5429), .B(n11220), .Y(n9946) );
  INVX3 U4338 ( .A(n9460), .Y(n6493) );
  INVX16 U4339 ( .A(net112356), .Y(net112350) );
  INVX8 U4340 ( .A(n10422), .Y(n10427) );
  NAND2BX2 U4341 ( .AN(n5426), .B(n11263), .Y(n9710) );
  BUFX6 U4342 ( .A(n6566), .Y(n3841) );
  NAND3X6 U4343 ( .A(ICACHE_addr[24]), .B(ICACHE_addr[23]), .C(n10316), .Y(
        n10342) );
  NOR4BBX4 U4344 ( .AN(ICACHE_addr[7]), .BN(ICACHE_addr[5]), .C(n224), .D(
        n10223), .Y(n10224) );
  NAND2X8 U4345 ( .A(ICACHE_addr[1]), .B(n4301), .Y(n10223) );
  OAI221X2 U4346 ( .A0(n8866), .A1(n4660), .B0(net103552), .B1(n7898), .C0(
        n6688), .Y(n7147) );
  NAND2X4 U4347 ( .A(n8641), .B(n6505), .Y(n7401) );
  OAI222X2 U4348 ( .A0(n7304), .A1(n7303), .B0(n7302), .B1(n7301), .C0(
        net104248), .C1(n9249), .Y(n7322) );
  NAND2BX4 U4349 ( .AN(n5427), .B(n11189), .Y(n10201) );
  NOR2X2 U4350 ( .A(n7164), .B(n7163), .Y(n7165) );
  NAND4X4 U4351 ( .A(n10001), .B(n10000), .C(n9999), .D(n9998), .Y(n11258) );
  OA22X1 U4352 ( .A0(n5391), .A1(n1642), .B0(n5345), .B1(n3224), .Y(n9998) );
  OA22X1 U4353 ( .A0(n5211), .A1(n1643), .B0(n5168), .B1(n3225), .Y(n10000) );
  BUFX20 U4354 ( .A(n5173), .Y(n5168) );
  NAND2X2 U4355 ( .A(n10423), .B(n10422), .Y(n10609) );
  NAND2X8 U4356 ( .A(\i_MIPS/ALUin1[18] ), .B(n6552), .Y(n8738) );
  CLKBUFX2 U4357 ( .A(n4797), .Y(n4794) );
  OAI2BB2X4 U4358 ( .B0(n8655), .B1(n3843), .A0N(n7814), .A1N(n8958), .Y(n7821) );
  OA22X4 U4359 ( .A0(n4987), .A1(n2125), .B0(n5033), .B1(n538), .Y(n6399) );
  CLKMX2X4 U4360 ( .A(n8739), .B(n7315), .S0(net107796), .Y(n9464) );
  NAND4X4 U4361 ( .A(n8598), .B(n8597), .C(n8596), .D(n8595), .Y(n11369) );
  NAND4BBX4 U4362 ( .AN(n10348), .BN(n9565), .C(n10350), .D(n6297), .Y(
        net98630) );
  NAND2X4 U4363 ( .A(n7969), .B(\i_MIPS/ALUin1[1] ), .Y(n6917) );
  OA22X2 U4364 ( .A0(n4917), .A1(n755), .B0(n4948), .B1(n2316), .Y(n7846) );
  OAI221X2 U4365 ( .A0(n8353), .A1(n4587), .B0(n4662), .B1(n6850), .C0(n8350), 
        .Y(n9246) );
  MX2XL U4366 ( .A(n3613), .B(n10775), .S0(n216), .Y(\i_MIPS/n389 ) );
  BUFX4 U4367 ( .A(net133469), .Y(net112116) );
  OA22X1 U4368 ( .A0(\i_MIPS/Register/register[6][28] ), .A1(net112116), .B0(
        \i_MIPS/Register/register[14][28] ), .B1(net112134), .Y(n8469) );
  NAND4X6 U4369 ( .A(n4327), .B(n6359), .C(n6358), .D(n6357), .Y(n11487) );
  NAND2X1 U4370 ( .A(n8151), .B(n8432), .Y(n6526) );
  NAND2X2 U4371 ( .A(\i_MIPS/ALUin1[26] ), .B(n6587), .Y(n8970) );
  INVX4 U4372 ( .A(n261), .Y(n6587) );
  NAND3X4 U4373 ( .A(n6298), .B(n4295), .C(n4664), .Y(n9986) );
  AO22XL U4374 ( .A0(net112002), .A1(n853), .B0(net112020), .B1(n2434), .Y(
        n7337) );
  AOI21X2 U4375 ( .A0(n7231), .A1(n8349), .B0(n4449), .Y(n4418) );
  OA22X2 U4376 ( .A0(n4918), .A1(n2289), .B0(n4948), .B1(n724), .Y(n7744) );
  AO22X1 U4377 ( .A0(n9531), .A1(n382), .B0(n4717), .B1(n2503), .Y(n8714) );
  AO22X1 U4378 ( .A0(n9531), .A1(n383), .B0(n4714), .B1(n2504), .Y(n8508) );
  AO22X1 U4379 ( .A0(n9531), .A1(n323), .B0(n4714), .B1(n2445), .Y(n8318) );
  AO22X1 U4380 ( .A0(n9531), .A1(n367), .B0(n4714), .B1(n2446), .Y(n8807) );
  MXI2X4 U4381 ( .A(n3709), .B(n10710), .S0(n5517), .Y(n10712) );
  OR4X6 U4382 ( .A(n8974), .B(n8973), .C(n8972), .D(n8971), .Y(n3894) );
  INVX4 U4383 ( .A(n8749), .Y(n8079) );
  OAI221X2 U4384 ( .A0(n4668), .A1(\i_MIPS/n345 ), .B0(n3828), .B1(
        \i_MIPS/n346 ), .C0(n6752), .Y(n8653) );
  OA22X2 U4385 ( .A0(n10911), .A1(n4245), .B0(n10914), .B1(n4246), .Y(n8025)
         );
  CLKBUFX3 U4386 ( .A(n5264), .Y(n5246) );
  NAND4X2 U4387 ( .A(n9603), .B(n9602), .C(n9601), .D(n9600), .Y(n11200) );
  NAND4X2 U4388 ( .A(n9558), .B(n4060), .C(n9568), .D(n11479), .Y(net97416) );
  NAND2X2 U4389 ( .A(n11349), .B(n9), .Y(n11478) );
  CLKBUFX4 U4390 ( .A(n9528), .Y(n4706) );
  NAND2X8 U4391 ( .A(n6536), .B(n7696), .Y(n7874) );
  NAND2X4 U4392 ( .A(n6585), .B(n3358), .Y(n8150) );
  AOI222X2 U4393 ( .A0(n5503), .A1(n11352), .B0(mem_rdata_D[2]), .B1(n234), 
        .C0(n12985), .C1(n5502), .Y(n10935) );
  INVX8 U4394 ( .A(n11352), .Y(n10934) );
  NAND4X4 U4395 ( .A(n6935), .B(n6934), .C(n6933), .D(n6932), .Y(n11352) );
  NAND2X1 U4396 ( .A(n3812), .B(\i_MIPS/ID_EX[78] ), .Y(n4076) );
  NAND2BX2 U4397 ( .AN(n5425), .B(n11280), .Y(n6286) );
  AND2X2 U4398 ( .A(n4662), .B(n7822), .Y(n4443) );
  INVX8 U4399 ( .A(n11401), .Y(n11004) );
  AOI222X1 U4400 ( .A0(n5512), .A1(n11401), .B0(mem_rdata_D[51]), .B1(n234), 
        .C0(n12968), .C1(n5507), .Y(n11005) );
  NAND4X4 U4401 ( .A(n8602), .B(n8601), .C(n8600), .D(n8599), .Y(n11401) );
  NOR4X6 U4402 ( .A(n9317), .B(n9316), .C(n9315), .D(n9314), .Y(n9318) );
  OAI21X1 U4403 ( .A0(n11349), .A1(n4620), .B0(n11345), .Y(n9982) );
  NAND4X8 U4404 ( .A(n4514), .B(n4515), .C(\i_MIPS/EX_MEM_0 ), .D(net111634), 
        .Y(net100426) );
  XNOR2X1 U4405 ( .A(n6606), .B(\i_MIPS/IR_ID[17] ), .Y(n4533) );
  MX2X1 U4406 ( .A(net112415), .B(net101082), .S0(n7709), .Y(n7710) );
  AO22X4 U4407 ( .A0(n7827), .A1(n9054), .B0(n7826), .B1(n3838), .Y(n7828) );
  NAND3BX4 U4408 ( .AN(n9490), .B(net112294), .C(n9489), .Y(n9496) );
  NAND3BX2 U4409 ( .AN(n9485), .B(net111992), .C(n9484), .Y(n9497) );
  OA22X1 U4410 ( .A0(n4749), .A1(n1215), .B0(n4791), .B1(n2752), .Y(n4356) );
  OAI222X4 U4411 ( .A0(net133471), .A1(n9347), .B0(n9331), .B1(n9467), .C0(
        n9352), .C1(net112420), .Y(n9345) );
  NAND4X4 U4412 ( .A(n8870), .B(n8869), .C(n8868), .D(n8867), .Y(n8879) );
  INVX1 U4413 ( .A(n8849), .Y(n8865) );
  NAND2X4 U4414 ( .A(net108664), .B(n4326), .Y(n10861) );
  MX2XL U4415 ( .A(\i_MIPS/ID_EX[49] ), .B(n5), .S0(n214), .Y(\i_MIPS/n421 )
         );
  AO21X4 U4416 ( .A0(n8728), .A1(n9145), .B0(n8727), .Y(n8746) );
  INVX1 U4417 ( .A(n8746), .Y(n8729) );
  OA22X2 U4418 ( .A0(n4917), .A1(n663), .B0(n4948), .B1(n2233), .Y(n7850) );
  NAND3BX2 U4419 ( .AN(n9153), .B(n4443), .C(net107804), .Y(n9459) );
  BUFX20 U4420 ( .A(net129024), .Y(net108664) );
  OA22X4 U4421 ( .A0(n10552), .A1(net133585), .B0(n10551), .B1(net108660), .Y(
        n10553) );
  OA22X1 U4422 ( .A0(n5123), .A1(n1644), .B0(n5089), .B1(n3226), .Y(n10130) );
  AND3X8 U4423 ( .A(n4331), .B(n4663), .C(n4666), .Y(n4330) );
  INVX1 U4424 ( .A(n8852), .Y(n7544) );
  NAND2X8 U4425 ( .A(n6563), .B(\i_MIPS/n348 ), .Y(n8851) );
  NAND4X6 U4426 ( .A(n7545), .B(n7547), .C(n7546), .D(net103840), .Y(n7548) );
  NAND2BX1 U4427 ( .AN(n4247), .B(n11286), .Y(n9909) );
  XNOR2X4 U4428 ( .A(n3931), .B(net112400), .Y(n10795) );
  OAI221X2 U4429 ( .A0(net112366), .A1(\i_MIPS/n347 ), .B0(net112348), .B1(
        \i_MIPS/n348 ), .C0(n6751), .Y(n7812) );
  OA22X4 U4430 ( .A0(n4669), .A1(\i_MIPS/n349 ), .B0(net112334), .B1(
        \i_MIPS/n350 ), .Y(n6751) );
  OA22X4 U4431 ( .A0(n4762), .A1(n2127), .B0(n4795), .B1(n541), .Y(n6418) );
  INVX12 U4432 ( .A(n1954), .Y(mem_wdata_D[34]) );
  CLKINVX2 U4433 ( .A(n9282), .Y(n9279) );
  INVX6 U4434 ( .A(n3686), .Y(n6543) );
  AOI2BB2X2 U4435 ( .B0(n10422), .B1(n3897), .A0N(n10426), .A1N(net108660), 
        .Y(n10428) );
  NAND4X4 U4436 ( .A(n7818), .B(n7817), .C(n4658), .D(n7816), .Y(n7830) );
  NAND4X1 U4437 ( .A(net103913), .B(net133411), .C(n3929), .D(net105600), .Y(
        net100791) );
  OAI222X1 U4438 ( .A0(\i_MIPS/PC/n22 ), .A1(net108686), .B0(n3637), .B1(
        n10531), .C0(n4428), .C1(net108704), .Y(n10537) );
  OAI222X1 U4439 ( .A0(\i_MIPS/PC/n5 ), .A1(net108688), .B0(n3637), .B1(n11078), .C0(n4409), .C1(net108702), .Y(n11084) );
  OAI222X1 U4440 ( .A0(\i_MIPS/PC/n24 ), .A1(net108688), .B0(net97445), .B1(
        n10549), .C0(n4426), .C1(net108704), .Y(n10555) );
  MX2XL U4441 ( .A(DCACHE_addr[29]), .B(n10866), .S0(n223), .Y(\i_MIPS/n438 )
         );
  CLKBUFX6 U4442 ( .A(n4677), .Y(n4678) );
  NAND2BXL U4443 ( .AN(n4247), .B(n11313), .Y(n6283) );
  NAND4X2 U4444 ( .A(n6180), .B(n6179), .C(n6178), .D(n6177), .Y(n11313) );
  AOI2BB1X4 U4445 ( .A0N(n6569), .A1N(n6580), .B0(n6568), .Y(n6582) );
  CLKMX2X3 U4446 ( .A(n9217), .B(n9216), .S0(net107810), .Y(n9220) );
  CLKINVX8 U4447 ( .A(net103025), .Y(net98351) );
  AOI2BB2X2 U4448 ( .B0(\i_MIPS/IF_ID[78] ), .B1(net108670), .A0N(net108676), 
        .A1N(\i_MIPS/n196 ), .Y(n10607) );
  OAI221XL U4449 ( .A0(net103718), .A1(net111624), .B0(net103719), .B1(
        net111636), .C0(net103720), .Y(n4617) );
  AOI222X2 U4450 ( .A0(\i_MIPS/IF_ID_29 ), .A1(net108682), .B0(
        \i_MIPS/IF_ID[94] ), .B1(net108670), .C0(net108710), .C1(n10692), .Y(
        n10581) );
  NAND2X8 U4451 ( .A(n9170), .B(net107804), .Y(net133688) );
  BUFX20 U4452 ( .A(net112128), .Y(net112134) );
  OA22X2 U4453 ( .A0(net112400), .A1(net133585), .B0(n10440), .B1(net108660), 
        .Y(n10441) );
  OAI222X1 U4454 ( .A0(\i_MIPS/PC/n19 ), .A1(net108686), .B0(n3637), .B1(
        n10439), .C0(n4429), .C1(net108704), .Y(n10443) );
  OAI22X1 U4455 ( .A0(n4414), .A1(net108704), .B0(\i_MIPS/PC/n30 ), .B1(
        net97444), .Y(n3858) );
  BUFX12 U4456 ( .A(n12793), .Y(mem_addr_D[16]) );
  AO22XL U4457 ( .A0(n12943), .A1(n11510), .B0(n4653), .B1(n11492), .Y(n12793)
         );
  NAND3BX2 U4458 ( .AN(n10845), .B(n10844), .C(n10843), .Y(\i_MIPS/PC/n61 ) );
  OAI222X1 U4459 ( .A0(\i_MIPS/PC/n29 ), .A1(net108690), .B0(n3637), .B1(
        n10839), .C0(n10838), .C1(net108702), .Y(n10845) );
  NAND3BX2 U4460 ( .AN(n10834), .B(n10833), .C(n10832), .Y(\i_MIPS/PC/n60 ) );
  OAI222X1 U4461 ( .A0(\i_MIPS/PC/n28 ), .A1(net108690), .B0(n3637), .B1(
        n10828), .C0(n4397), .C1(net108702), .Y(n10834) );
  OAI222X1 U4462 ( .A0(\i_MIPS/PC/n18 ), .A1(net108686), .B0(n3637), .B1(
        n10615), .C0(net128955), .C1(net108702), .Y(n10620) );
  AOI2BB2X1 U4463 ( .B0(n3860), .B1(net108708), .A0N(\i_MIPS/PC/n3 ), .A1N(
        net108690), .Y(n10527) );
  BUFX12 U4464 ( .A(n12791), .Y(mem_addr_D[27]) );
  BUFX12 U4465 ( .A(n12792), .Y(mem_addr_D[17]) );
  AO22XL U4466 ( .A0(n12942), .A1(n4637), .B0(n4654), .B1(n11493), .Y(n12792)
         );
  OA22X4 U4467 ( .A0(n5210), .A1(n2988), .B0(n5167), .B1(n1431), .Y(n9956) );
  OA22X2 U4468 ( .A0(n5301), .A1(n1467), .B0(n5247), .B1(n3041), .Y(n9955) );
  BUFX12 U4469 ( .A(n12790), .Y(mem_addr_D[28]) );
  AO22XL U4470 ( .A0(n12931), .A1(n4637), .B0(n5551), .B1(n11504), .Y(n12790)
         );
  BUFX12 U4471 ( .A(n12788), .Y(mem_addr_D[30]) );
  AO22X1 U4472 ( .A0(DCACHE_addr[28]), .A1(n11510), .B0(n5551), .B1(n11506), 
        .Y(n12788) );
  OAI21X1 U4473 ( .A0(\i_MIPS/n237 ), .A1(net108190), .B0(n10524), .Y(
        \i_MIPS/N91 ) );
  OAI21X1 U4474 ( .A0(\i_MIPS/n183 ), .A1(net108190), .B0(n10524), .Y(
        \i_MIPS/N26 ) );
  MX2X1 U4475 ( .A(\D_cache/cache[0][46] ), .B(n10746), .S0(n4739), .Y(
        \D_cache/n1428 ) );
  CLKMX2X2 U4476 ( .A(\D_cache/cache[1][46] ), .B(n10746), .S0(n4785), .Y(
        \D_cache/n1427 ) );
  CLKMX2X2 U4477 ( .A(\D_cache/cache[2][46] ), .B(n10746), .S0(n4807), .Y(
        \D_cache/n1426 ) );
  CLKMX2X2 U4478 ( .A(\D_cache/cache[3][46] ), .B(n10746), .S0(n4851), .Y(
        \D_cache/n1425 ) );
  CLKMX2X2 U4479 ( .A(\D_cache/cache[4][46] ), .B(n10746), .S0(n4897), .Y(
        \D_cache/n1424 ) );
  CLKMX2X2 U4480 ( .A(\D_cache/cache[5][46] ), .B(n10746), .S0(n4942), .Y(
        \D_cache/n1423 ) );
  CLKMX2X2 U4481 ( .A(\D_cache/cache[6][46] ), .B(n10746), .S0(n4961), .Y(
        \D_cache/n1422 ) );
  CLKMX2X2 U4482 ( .A(\D_cache/cache[7][46] ), .B(n10746), .S0(n5005), .Y(
        \D_cache/n1421 ) );
  MXI2X4 U4483 ( .A(n10745), .B(n10744), .S0(n5518), .Y(n10746) );
  CLKMX2X2 U4484 ( .A(\D_cache/cache[0][45] ), .B(n10735), .S0(n4739), .Y(
        \D_cache/n1436 ) );
  CLKMX2X2 U4485 ( .A(\D_cache/cache[1][45] ), .B(n10735), .S0(n4784), .Y(
        \D_cache/n1435 ) );
  CLKMX2X2 U4486 ( .A(\D_cache/cache[5][45] ), .B(n10735), .S0(n4941), .Y(
        \D_cache/n1431 ) );
  CLKMX2X2 U4487 ( .A(\D_cache/cache[7][44] ), .B(n10724), .S0(n5004), .Y(
        \D_cache/n1437 ) );
  CLKMX2X2 U4488 ( .A(\D_cache/cache[6][44] ), .B(n10724), .S0(n4960), .Y(
        \D_cache/n1438 ) );
  CLKMX2X2 U4489 ( .A(\D_cache/cache[4][44] ), .B(n10724), .S0(n4896), .Y(
        \D_cache/n1440 ) );
  CLKMX2X2 U4490 ( .A(\D_cache/cache[3][44] ), .B(n10724), .S0(n4850), .Y(
        \D_cache/n1441 ) );
  CLKMX2X2 U4491 ( .A(\D_cache/cache[2][44] ), .B(n10724), .S0(n4806), .Y(
        \D_cache/n1442 ) );
  CLKMX2X2 U4492 ( .A(\D_cache/cache[1][44] ), .B(n10724), .S0(n4785), .Y(
        \D_cache/n1443 ) );
  MX2X1 U4493 ( .A(\D_cache/cache[0][44] ), .B(n10724), .S0(n4737), .Y(
        \D_cache/n1444 ) );
  NAND3BX4 U4494 ( .AN(n10462), .B(n10461), .C(n10460), .Y(\i_MIPS/PC/n58 ) );
  CLKMX2X2 U4495 ( .A(\D_cache/cache[7][107] ), .B(n10715), .S0(n5004), .Y(
        \D_cache/n933 ) );
  CLKMX2X2 U4496 ( .A(\D_cache/cache[6][107] ), .B(n10715), .S0(n4960), .Y(
        \D_cache/n934 ) );
  CLKMX2X2 U4497 ( .A(\D_cache/cache[4][107] ), .B(n10715), .S0(n4896), .Y(
        \D_cache/n936 ) );
  CLKMX2X2 U4498 ( .A(\D_cache/cache[3][107] ), .B(n10715), .S0(n4850), .Y(
        \D_cache/n937 ) );
  CLKMX2X2 U4499 ( .A(\D_cache/cache[2][107] ), .B(n10715), .S0(n4806), .Y(
        \D_cache/n938 ) );
  CLKMX2X2 U4500 ( .A(\D_cache/cache[1][107] ), .B(n10715), .S0(n4785), .Y(
        \D_cache/n939 ) );
  MX2X1 U4501 ( .A(\D_cache/cache[0][107] ), .B(n10715), .S0(n4738), .Y(
        \D_cache/n940 ) );
  MXI2X4 U4502 ( .A(n10748), .B(n10747), .S0(n5518), .Y(n10749) );
  MX2X1 U4503 ( .A(\D_cache/cache[1][108] ), .B(n10727), .S0(n4783), .Y(
        \D_cache/n931 ) );
  MX2X1 U4504 ( .A(\D_cache/cache[2][108] ), .B(n10727), .S0(n4803), .Y(
        \D_cache/n930 ) );
  MX2X1 U4505 ( .A(\D_cache/cache[3][108] ), .B(n10727), .S0(n4848), .Y(
        \D_cache/n929 ) );
  MX2X1 U4506 ( .A(\D_cache/cache[4][108] ), .B(n10727), .S0(n4898), .Y(
        \D_cache/n928 ) );
  MX2X1 U4507 ( .A(\D_cache/cache[5][108] ), .B(n10727), .S0(n4940), .Y(
        \D_cache/n927 ) );
  MX2X1 U4508 ( .A(\D_cache/cache[6][108] ), .B(n10727), .S0(n4958), .Y(
        \D_cache/n926 ) );
  MX2X1 U4509 ( .A(\D_cache/cache[7][108] ), .B(n10727), .S0(n5008), .Y(
        \D_cache/n925 ) );
  MXI2X4 U4510 ( .A(n10726), .B(n10725), .S0(n5518), .Y(n10727) );
  OA22X2 U4511 ( .A0(n5209), .A1(n1468), .B0(n5166), .B1(n3042), .Y(n9900) );
  AOI2BB2X2 U4512 ( .B0(\i_MIPS/IF_ID[81] ), .B1(net108670), .A0N(net108676), 
        .A1N(\i_MIPS/n199 ), .Y(n10619) );
  AOI2BB2X2 U4513 ( .B0(\i_MIPS/IF_ID[72] ), .B1(n3930), .A0N(net108676), 
        .A1N(\i_MIPS/n190 ), .Y(n10808) );
  AOI2BB2X2 U4514 ( .B0(\i_MIPS/IF_ID[68] ), .B1(n3930), .A0N(net108676), 
        .A1N(\i_MIPS/n186 ), .Y(n11083) );
  BUFX16 U4515 ( .A(n15), .Y(net108680) );
  MX2X1 U4516 ( .A(\D_cache/cache[1][51] ), .B(n10997), .S0(n4786), .Y(
        \D_cache/n1387 ) );
  MX2X1 U4517 ( .A(\D_cache/cache[0][51] ), .B(n10997), .S0(n4738), .Y(
        \D_cache/n1388 ) );
  NAND3BX4 U4518 ( .AN(n10381), .B(n10380), .C(n10379), .Y(\i_MIPS/PC/n42 ) );
  XOR3X2 U4519 ( .A(net112400), .B(net98502), .C(net98487), .Y(net98495) );
  AOI2BB2X2 U4520 ( .B0(n10611), .B1(n3897), .A0N(n10616), .A1N(net108658), 
        .Y(n10618) );
  OA22X2 U4521 ( .A0(n4432), .A1(net108704), .B0(\i_MIPS/PC/n2 ), .B1(
        net108686), .Y(n10522) );
  OA22X4 U4522 ( .A0(n10630), .A1(net133585), .B0(n10629), .B1(net108658), .Y(
        n10631) );
  OAI222X1 U4523 ( .A0(\i_MIPS/PC/n16 ), .A1(net108690), .B0(n3637), .B1(
        n10410), .C0(n4401), .C1(net108704), .Y(n10415) );
  BUFX12 U4524 ( .A(n5128), .Y(n5104) );
  CLKAND2X12 U4525 ( .A(DCACHE_addr[2]), .B(n11481), .Y(mem_addr_D[4]) );
  BUFX12 U4526 ( .A(n12798), .Y(mem_addr_D[5]) );
  AND2XL U4527 ( .A(DCACHE_addr[3]), .B(n11481), .Y(n12798) );
  NOR4X2 U4528 ( .A(n8410), .B(n8409), .C(n8408), .D(n8407), .Y(n8411) );
  AO22X1 U4529 ( .A0(n4729), .A1(n368), .B0(n4725), .B1(n1022), .Y(n8407) );
  NAND2X8 U4530 ( .A(n409), .B(n10394), .Y(n10401) );
  OAI221X2 U4531 ( .A0(net104251), .A1(net111624), .B0(net104252), .B1(
        net111636), .C0(net104253), .Y(n4137) );
  AOI33X2 U4532 ( .A0(n9070), .A1(n9069), .A2(net112292), .B0(n9068), .B1(
        n9067), .B2(net112292), .Y(n9071) );
  OAI222X1 U4533 ( .A0(\i_MIPS/PC/n9 ), .A1(net108688), .B0(n3637), .B1(n10804), .C0(n4405), .C1(net108702), .Y(n10809) );
  MX2XL U4534 ( .A(\i_MIPS/ALU/N303 ), .B(n3808), .S0(n222), .Y(\i_MIPS/n531 )
         );
  INVX2 U4535 ( .A(n11408), .Y(n10278) );
  NAND4X2 U4536 ( .A(n7275), .B(n7274), .C(n7273), .D(n7272), .Y(n11361) );
  INVX2 U4537 ( .A(n11361), .Y(n10713) );
  OAI222X1 U4538 ( .A0(\i_MIPS/PC/n21 ), .A1(net108686), .B0(n3637), .B1(
        n10637), .C0(n11007), .C1(net108702), .Y(n10649) );
  INVX4 U4539 ( .A(n11445), .Y(n10871) );
  INVX4 U4540 ( .A(n11396), .Y(n10750) );
  INVXL U4541 ( .A(net103719), .Y(n3875) );
  BUFX4 U4542 ( .A(n5533), .Y(n5538) );
  CLKBUFX4 U4543 ( .A(n5037), .Y(n5024) );
  NAND4X4 U4544 ( .A(n7656), .B(n7655), .C(n7654), .D(n7653), .Y(n11364) );
  INVX2 U4545 ( .A(n11365), .Y(n10758) );
  BUFX12 U4546 ( .A(n12799), .Y(mem_wdata_D[76]) );
  AND2XL U4547 ( .A(n4653), .B(n11426), .Y(n12799) );
  OA22X2 U4548 ( .A0(n10646), .A1(net133585), .B0(n10645), .B1(net108658), .Y(
        n10647) );
  OA22X2 U4549 ( .A0(n11126), .A1(net133585), .B0(n11125), .B1(net108658), .Y(
        n11127) );
  OAI22X1 U4550 ( .A0(n5103), .A1(n649), .B0(n5079), .B1(n2226), .Y(n4339) );
  BUFX20 U4551 ( .A(n5085), .Y(n5061) );
  INVX4 U4552 ( .A(n11451), .Y(n10978) );
  OA22X1 U4553 ( .A0(n5288), .A1(n1645), .B0(n5241), .B1(n3227), .Y(n6143) );
  OA22X1 U4554 ( .A0(n5395), .A1(n1646), .B0(n5332), .B1(n3228), .Y(n6142) );
  AND3X8 U4555 ( .A(n3926), .B(n3652), .C(n4218), .Y(net112676) );
  MX2XL U4556 ( .A(n3599), .B(n3741), .S0(n216), .Y(\i_MIPS/n409 ) );
  CLKMX2X2 U4557 ( .A(\D_cache/cache[7][50] ), .B(n10513), .S0(n5001), .Y(
        \D_cache/n1389 ) );
  CLKMX2X2 U4558 ( .A(\D_cache/cache[6][50] ), .B(n10513), .S0(n4957), .Y(
        \D_cache/n1390 ) );
  CLKMX2X2 U4559 ( .A(\D_cache/cache[5][50] ), .B(n10513), .S0(n4936), .Y(
        \D_cache/n1391 ) );
  CLKMX2X2 U4560 ( .A(\D_cache/cache[4][50] ), .B(n10513), .S0(n4893), .Y(
        \D_cache/n1392 ) );
  CLKMX2X2 U4561 ( .A(\D_cache/cache[3][50] ), .B(n10513), .S0(n4847), .Y(
        \D_cache/n1393 ) );
  CLKMX2X2 U4562 ( .A(\D_cache/cache[2][50] ), .B(n10513), .S0(n4802), .Y(
        \D_cache/n1394 ) );
  CLKMX2X2 U4563 ( .A(\D_cache/cache[1][50] ), .B(n10513), .S0(n4779), .Y(
        \D_cache/n1395 ) );
  NAND4X4 U4564 ( .A(n7580), .B(n7579), .C(n7578), .D(n7577), .Y(n11414) );
  INVX2 U4565 ( .A(n11414), .Y(n10956) );
  AOI2BB1X4 U4566 ( .A0N(net112764), .A1N(\i_MIPS/n340 ), .B0(n6772), .Y(n3884) );
  BUFX12 U4567 ( .A(n12803), .Y(mem_wdata_D[23]) );
  AND2XL U4568 ( .A(n5551), .B(n11373), .Y(n12803) );
  BUFX12 U4569 ( .A(n12802), .Y(mem_wdata_D[25]) );
  AND2XL U4570 ( .A(n5551), .B(n11375), .Y(n12802) );
  BUFX12 U4571 ( .A(n12801), .Y(mem_wdata_D[37]) );
  AND2XL U4572 ( .A(n5551), .B(n11387), .Y(n12801) );
  BUFX12 U4573 ( .A(n12800), .Y(mem_wdata_D[39]) );
  AND2XL U4574 ( .A(n5551), .B(n11389), .Y(n12800) );
  NAND4X4 U4575 ( .A(n7934), .B(n7933), .C(n7932), .D(n7931), .Y(n11453) );
  OA22X2 U4576 ( .A0(n4917), .A1(n757), .B0(n4948), .B1(n2318), .Y(n7932) );
  AOI2BB1X2 U4577 ( .A0N(net112346), .A1N(n7696), .B0(net127833), .Y(n7058) );
  INVX8 U4578 ( .A(n11442), .Y(n10478) );
  NAND4X4 U4579 ( .A(n9091), .B(n9090), .C(n9089), .D(n9088), .Y(n11407) );
  OA22X2 U4580 ( .A0(n4968), .A1(n664), .B0(n5027), .B1(n2234), .Y(n9088) );
  INVX8 U4581 ( .A(n11407), .Y(n10500) );
  AO22X1 U4582 ( .A0(DCACHE_addr[12]), .A1(n4637), .B0(n4654), .B1(n11490), 
        .Y(n12794) );
  CLKMX2X2 U4583 ( .A(\i_MIPS/n340 ), .B(\i_MIPS/n341 ), .S0(net112338), .Y(
        net104866) );
  NAND2XL U4584 ( .A(net112340), .B(\i_MIPS/ALUin1[30] ), .Y(n6494) );
  OAI211XL U4585 ( .A0(n10249), .A1(n10432), .B0(n10622), .C0(n10435), .Y(
        n3889) );
  CLKMX2X2 U4586 ( .A(\D_cache/cache[7][59] ), .B(n10306), .S0(n5000), .Y(
        \D_cache/n1317 ) );
  CLKMX2X2 U4587 ( .A(\D_cache/cache[6][59] ), .B(n10306), .S0(n4956), .Y(
        \D_cache/n1318 ) );
  CLKMX2X2 U4588 ( .A(\D_cache/cache[5][59] ), .B(n10306), .S0(n4936), .Y(
        \D_cache/n1319 ) );
  CLKMX2X2 U4589 ( .A(\D_cache/cache[4][59] ), .B(n10306), .S0(n4892), .Y(
        \D_cache/n1320 ) );
  CLKMX2X2 U4590 ( .A(\D_cache/cache[3][59] ), .B(n10306), .S0(n4846), .Y(
        \D_cache/n1321 ) );
  CLKMX2X2 U4591 ( .A(\D_cache/cache[2][59] ), .B(n10306), .S0(n4801), .Y(
        \D_cache/n1322 ) );
  CLKMX2X2 U4592 ( .A(\D_cache/cache[1][59] ), .B(n10306), .S0(n4778), .Y(
        \D_cache/n1323 ) );
  MX2X1 U4593 ( .A(\D_cache/cache[0][59] ), .B(n10306), .S0(n4732), .Y(
        \D_cache/n1324 ) );
  CLKMX2X2 U4594 ( .A(\D_cache/cache[7][57] ), .B(n10496), .S0(n5000), .Y(
        \D_cache/n1333 ) );
  CLKMX2X2 U4595 ( .A(\D_cache/cache[6][57] ), .B(n10496), .S0(n4956), .Y(
        \D_cache/n1334 ) );
  CLKMX2X2 U4596 ( .A(\D_cache/cache[5][57] ), .B(n10496), .S0(n4941), .Y(
        \D_cache/n1335 ) );
  CLKMX2X2 U4597 ( .A(\D_cache/cache[4][57] ), .B(n10496), .S0(n4892), .Y(
        \D_cache/n1336 ) );
  CLKMX2X2 U4598 ( .A(\D_cache/cache[3][57] ), .B(n10496), .S0(n4846), .Y(
        \D_cache/n1337 ) );
  CLKMX2X2 U4599 ( .A(\D_cache/cache[2][57] ), .B(n10496), .S0(n4801), .Y(
        \D_cache/n1338 ) );
  CLKMX2X2 U4600 ( .A(\D_cache/cache[1][57] ), .B(n10496), .S0(n4778), .Y(
        \D_cache/n1339 ) );
  MX2X1 U4601 ( .A(\D_cache/cache[0][57] ), .B(n10496), .S0(n4732), .Y(
        \D_cache/n1340 ) );
  INVXL U4602 ( .A(n7300), .Y(n7304) );
  AO22X4 U4603 ( .A0(n9054), .A1(net128963), .B0(n3838), .B1(n8966), .Y(n8741)
         );
  CLKMX2X2 U4604 ( .A(\D_cache/cache[7][62] ), .B(n10144), .S0(n5008), .Y(
        \D_cache/n1293 ) );
  CLKMX2X2 U4605 ( .A(\D_cache/cache[6][62] ), .B(n10144), .S0(n4964), .Y(
        \D_cache/n1294 ) );
  CLKMX2X2 U4606 ( .A(\D_cache/cache[5][62] ), .B(n10144), .S0(n4936), .Y(
        \D_cache/n1295 ) );
  CLKMX2X2 U4607 ( .A(\D_cache/cache[4][62] ), .B(n10144), .S0(n4894), .Y(
        \D_cache/n1296 ) );
  CLKMX2X2 U4608 ( .A(\D_cache/cache[3][62] ), .B(n10144), .S0(n4849), .Y(
        \D_cache/n1297 ) );
  CLKMX2X2 U4609 ( .A(\D_cache/cache[2][62] ), .B(n10144), .S0(n4803), .Y(
        \D_cache/n1298 ) );
  CLKMX2X2 U4610 ( .A(\D_cache/cache[1][62] ), .B(n10144), .S0(n4780), .Y(
        \D_cache/n1299 ) );
  AO22X4 U4611 ( .A0(mem_rdata_I[24]), .A1(n5541), .B0(n253), .B1(n11210), .Y(
        n9797) );
  AO22X4 U4612 ( .A0(mem_rdata_I[56]), .A1(n5541), .B0(n252), .B1(n11242), .Y(
        n9801) );
  AO22X4 U4613 ( .A0(mem_rdata_I[121]), .A1(n5541), .B0(n251), .B1(n11307), 
        .Y(n9809) );
  AO22X4 U4614 ( .A0(mem_rdata_I[57]), .A1(n5541), .B0(n249), .B1(n11243), .Y(
        n9821) );
  OAI2BB1X4 U4615 ( .A0N(n8637), .A1N(n8636), .B0(n8635), .Y(n8638) );
  INVX6 U4616 ( .A(n8638), .Y(n8640) );
  AOI222X2 U4617 ( .A0(n5495), .A1(n11476), .B0(mem_rdata_D[126]), .B1(n234), 
        .C0(n12957), .C1(n5494), .Y(n10140) );
  OA22X2 U4618 ( .A0(n4969), .A1(n685), .B0(n5014), .B1(n2257), .Y(n9084) );
  AOI31X2 U4619 ( .A0(n7411), .A1(n7412), .A2(n4433), .B0(n8241), .Y(n6584) );
  AND2X4 U4620 ( .A(net112356), .B(\i_MIPS/n354 ), .Y(n4472) );
  OAI221X2 U4621 ( .A0(\i_MIPS/ALUin1[11] ), .A1(net112364), .B0(
        \i_MIPS/ALUin1[10] ), .B1(net112348), .C0(n6839), .Y(n7062) );
  AO22X1 U4622 ( .A0(n4729), .A1(n384), .B0(n4725), .B1(n1034), .Y(n8416) );
  XOR2X4 U4623 ( .A(n259), .B(\i_MIPS/IR_ID[25] ), .Y(n6451) );
  OAI211X2 U4624 ( .A0(n3412), .A1(net111636), .B0(n9432), .C0(n9431), .Y(
        n3890) );
  OAI211XL U4625 ( .A0(n3412), .A1(net111636), .B0(n9432), .C0(n9431), .Y(
        n10318) );
  AO21X4 U4626 ( .A0(n10281), .A1(n10282), .B0(net111640), .Y(n9017) );
  AO22X1 U4627 ( .A0(n4729), .A1(n985), .B0(n4725), .B1(n2505), .Y(n8037) );
  NAND2X4 U4628 ( .A(net98502), .B(net112404), .Y(n10449) );
  INVX3 U4629 ( .A(net98497), .Y(net98502) );
  MXI2X2 U4630 ( .A(n10960), .B(n10959), .S0(n5522), .Y(n10961) );
  INVX3 U4631 ( .A(n11350), .Y(n10959) );
  OAI2BB1X4 U4632 ( .A0N(n10565), .A1N(n10564), .B0(net111646), .Y(n9324) );
  OA22X2 U4633 ( .A0(n4973), .A1(n686), .B0(n5018), .B1(n2258), .Y(n8487) );
  AO22X2 U4634 ( .A0(n5544), .A1(ICACHE_addr[29]), .B0(n240), .B1(n11344), .Y(
        n11152) );
  MX2X1 U4635 ( .A(\D_cache/cache[3][0] ), .B(n182), .S0(n4854), .Y(
        \D_cache/n1792 ) );
  MX2XL U4636 ( .A(n3601), .B(n2), .S0(n211), .Y(\i_MIPS/n413 ) );
  AO22X4 U4637 ( .A0(net112008), .A1(n441), .B0(net112026), .B1(n2024), .Y(
        n9236) );
  AO22X4 U4638 ( .A0(net112008), .A1(n274), .B0(net112026), .B1(n306), .Y(
        n9366) );
  MXI2X4 U4639 ( .A(n10479), .B(n10478), .S0(n5515), .Y(n10480) );
  OA22X2 U4640 ( .A0(n10806), .A1(net133585), .B0(n10805), .B1(net108658), .Y(
        n10807) );
  OA22X2 U4641 ( .A0(n11081), .A1(net133585), .B0(n11080), .B1(net108658), .Y(
        n11082) );
  OA22X2 U4642 ( .A0(n10378), .A1(net133585), .B0(n10377), .B1(net108658), .Y(
        n10379) );
  OA22X1 U4643 ( .A0(\i_MIPS/Register/register[22][6] ), .A1(n4683), .B0(
        \i_MIPS/Register/register[30][6] ), .B1(n4680), .Y(n7031) );
  OA22X1 U4644 ( .A0(\i_MIPS/Register/register[22][8] ), .A1(n4683), .B0(
        \i_MIPS/Register/register[30][8] ), .B1(n4680), .Y(n7116) );
  OA22X1 U4645 ( .A0(\i_MIPS/Register/register[22][13] ), .A1(n4683), .B0(
        \i_MIPS/Register/register[30][13] ), .B1(n4680), .Y(n7766) );
  OA22X1 U4646 ( .A0(\i_MIPS/Register/register[6][8] ), .A1(n4683), .B0(
        \i_MIPS/Register/register[14][8] ), .B1(n4680), .Y(n7107) );
  OA22X1 U4647 ( .A0(\i_MIPS/Register/register[6][13] ), .A1(n4683), .B0(
        \i_MIPS/Register/register[14][13] ), .B1(n4680), .Y(n7757) );
  OA22X1 U4648 ( .A0(\i_MIPS/Register/register[22][14] ), .A1(n4683), .B0(
        \i_MIPS/Register/register[30][14] ), .B1(n4680), .Y(n7672) );
  OA22X1 U4649 ( .A0(\i_MIPS/Register/register[6][14] ), .A1(n4683), .B0(
        \i_MIPS/Register/register[14][14] ), .B1(n4680), .Y(n7663) );
  OA22X1 U4650 ( .A0(\i_MIPS/Register/register[22][12] ), .A1(n4683), .B0(
        \i_MIPS/Register/register[30][12] ), .B1(n4680), .Y(n7452) );
  CLKMX2X2 U4651 ( .A(\I_cache/cache[0][79] ), .B(n9658), .S0(n5092), .Y(
        n12155) );
  MX2X1 U4652 ( .A(\I_cache/cache[1][79] ), .B(n9658), .S0(n5050), .Y(n12154)
         );
  MX2X1 U4653 ( .A(\I_cache/cache[2][118] ), .B(n9873), .S0(n5187), .Y(n11841)
         );
  INVX8 U4654 ( .A(n11357), .Y(n10887) );
  AOI222X2 U4655 ( .A0(n5505), .A1(n11357), .B0(mem_rdata_D[7]), .B1(n235), 
        .C0(n12980), .C1(n5502), .Y(n10888) );
  NAND4X4 U4656 ( .A(n7942), .B(n7941), .C(n7940), .D(n7939), .Y(n11357) );
  MXI2X4 U4657 ( .A(n10888), .B(n10887), .S0(n5520), .Y(n10889) );
  INVX8 U4658 ( .A(n7234), .Y(n7893) );
  INVX1 U4659 ( .A(n7219), .Y(n8632) );
  AO21X4 U4660 ( .A0(n8634), .A1(n8633), .B0(n8632), .Y(n8639) );
  OA22X4 U4661 ( .A0(n4970), .A1(n2078), .B0(n5015), .B1(n490), .Y(n8888) );
  NAND4X4 U4662 ( .A(n8891), .B(n8890), .C(n8889), .D(n8888), .Y(n11373) );
  OA22X2 U4663 ( .A0(n4817), .A1(n2408), .B0(n4863), .B1(n674), .Y(n8890) );
  AOI211X2 U4664 ( .A0(n7905), .A1(net101908), .B0(n7904), .C0(n7903), .Y(
        n7906) );
  INVX4 U4665 ( .A(n10464), .Y(n10339) );
  OAI2BB1X4 U4666 ( .A0N(n8874), .A1N(n4536), .B0(n8648), .Y(n8875) );
  INVX4 U4667 ( .A(n10822), .Y(n10825) );
  NAND4X6 U4668 ( .A(n10016), .B(n10015), .C(n10014), .D(n10013), .Y(n10812)
         );
  INVX3 U4669 ( .A(n11463), .Y(n10763) );
  OAI221XL U4670 ( .A0(n9548), .A1(net111622), .B0(n9547), .B1(net111634), 
        .C0(n9546), .Y(n10208) );
  NAND4X4 U4671 ( .A(n9195), .B(n9194), .C(n9193), .D(n9192), .Y(n11403) );
  OA22X1 U4672 ( .A0(n4968), .A1(n1082), .B0(n5027), .B1(n2675), .Y(n9192) );
  INVX8 U4673 ( .A(n11403), .Y(n10676) );
  AOI2BB2X2 U4674 ( .B0(\i_MIPS/IF_ID[77] ), .B1(n3930), .A0N(net108674), 
        .A1N(\i_MIPS/n195 ), .Y(n10397) );
  AO22X4 U4675 ( .A0(n7228), .A1(n7227), .B0(n7226), .B1(n8347), .Y(n7238) );
  INVX3 U4676 ( .A(n11471), .Y(n10491) );
  NAND4X4 U4677 ( .A(n6145), .B(n6144), .C(n6143), .D(n6142), .Y(n11250) );
  NAND2BX2 U4678 ( .AN(n5429), .B(n11218), .Y(n9950) );
  INVX2 U4679 ( .A(n9332), .Y(n9337) );
  AO22X2 U4680 ( .A0(n4471), .A1(n9328), .B0(n4418), .B1(n9327), .Y(n9346) );
  BUFX20 U4681 ( .A(n4476), .Y(n4671) );
  OA22X1 U4682 ( .A0(n5123), .A1(n1647), .B0(n5054), .B1(n3229), .Y(n10125) );
  MXI2X1 U4683 ( .A(\i_MIPS/n333 ), .B(\i_MIPS/n332 ), .S0(n208), .Y(
        \i_MIPS/n523 ) );
  AO21X4 U4684 ( .A0(net98391), .A1(net98390), .B0(net111642), .Y(net104584)
         );
  AO21X4 U4685 ( .A0(n10222), .A1(n10221), .B0(net111642), .Y(n9546) );
  NAND2X6 U4686 ( .A(n6963), .B(n6964), .Y(n7044) );
  BUFX6 U4687 ( .A(n5264), .Y(n5263) );
  NAND4X6 U4688 ( .A(n9389), .B(n9388), .C(n9387), .D(n9386), .Y(n11441) );
  OA22X4 U4689 ( .A0(n4966), .A1(n2079), .B0(n5012), .B1(n491), .Y(n9386) );
  OAI221X2 U4690 ( .A0(n4660), .A1(n9160), .B0(net103552), .B1(n9059), .C0(
        n7700), .Y(n8163) );
  AO22X2 U4691 ( .A0(\i_MIPS/ALUin1[1] ), .A1(net112338), .B0(
        \i_MIPS/ALUin1[0] ), .B1(n4672), .Y(n9059) );
  OA22X2 U4692 ( .A0(n10719), .A1(n4676), .B0(n10722), .B1(n4250), .Y(n7442)
         );
  XNOR2X4 U4693 ( .A(n3898), .B(n4133), .Y(n3946) );
  AO22XL U4694 ( .A0(n4731), .A1(n852), .B0(n4725), .B1(n2437), .Y(n7758) );
  AO22X2 U4695 ( .A0(net112000), .A1(n640), .B0(net112018), .B1(n2215), .Y(
        n4110) );
  AO22X4 U4696 ( .A0(net112000), .A1(n443), .B0(net112018), .B1(n2026), .Y(
        n4119) );
  NAND2X2 U4697 ( .A(n4470), .B(n7164), .Y(n8244) );
  NAND3BX4 U4698 ( .AN(n4664), .B(n6298), .C(n4295), .Y(n4332) );
  MXI2X2 U4699 ( .A(n3844), .B(n9154), .S0(net107794), .Y(n8654) );
  CLKAND2X8 U4700 ( .A(n7692), .B(n9457), .Y(n4470) );
  OAI221X2 U4701 ( .A0(\i_MIPS/ALUin1[21] ), .A1(net112364), .B0(
        \i_MIPS/ALUin1[22] ), .B1(net112346), .C0(n8248), .Y(n8456) );
  NAND2BX2 U4702 ( .AN(n5429), .B(n11223), .Y(n9930) );
  AO22X2 U4703 ( .A0(mem_rdata_I[37]), .A1(n5537), .B0(n249), .B1(n11223), .Y(
        n9929) );
  NAND4X2 U4704 ( .A(n9928), .B(n9927), .C(n9926), .D(n9925), .Y(n11223) );
  NAND2X8 U4705 ( .A(\i_MIPS/IF_ID[97] ), .B(n9559), .Y(n3926) );
  NAND4BX4 U4706 ( .AN(n4340), .B(n9301), .C(n9300), .D(n9299), .Y(n11402) );
  AOI222X2 U4707 ( .A0(n7895), .A1(net103224), .B0(n7894), .B1(net100585), 
        .C0(n7893), .C1(n7892), .Y(n7907) );
  OA22X2 U4708 ( .A0(n4756), .A1(n759), .B0(n4793), .B1(n2320), .Y(n7351) );
  BUFX2 U4709 ( .A(n4768), .Y(n4756) );
  OAI221X1 U4710 ( .A0(\i_MIPS/Register/register[18][12] ), .A1(net112072), 
        .B0(\i_MIPS/Register/register[26][12] ), .B1(net112098), .C0(n7393), 
        .Y(n7396) );
  MXI2X1 U4711 ( .A(\i_MIPS/n331 ), .B(\i_MIPS/n330 ), .S0(n205), .Y(
        \i_MIPS/n522 ) );
  MX2XL U4712 ( .A(n12952), .B(net97834), .S0(n207), .Y(\i_MIPS/n462 ) );
  NAND4BX4 U4713 ( .AN(n8464), .B(n3900), .C(n8463), .D(n8462), .Y(n10320) );
  BUFX12 U4714 ( .A(net97444), .Y(net108688) );
  OA22X4 U4715 ( .A0(n4972), .A1(n2080), .B0(n5017), .B1(n492), .Y(n8591) );
  OA22X4 U4716 ( .A0(n4972), .A1(n2131), .B0(n5017), .B1(n545), .Y(n8599) );
  OA22X4 U4717 ( .A0(n4972), .A1(n2133), .B0(n5017), .B1(n547), .Y(n8684) );
  CLKINVX1 U4718 ( .A(n10439), .Y(n10437) );
  CLKXOR2X2 U4719 ( .A(n10248), .B(ICACHE_addr[15]), .Y(n10439) );
  NAND2X4 U4720 ( .A(n10437), .B(n4571), .Y(n10622) );
  OAI2BB2X1 U4721 ( .B0(\i_MIPS/n200 ), .B1(net108194), .A0N(n10437), .A1N(
        n4073), .Y(\i_MIPS/N43 ) );
  NAND4X4 U4722 ( .A(n4354), .B(n9294), .C(n9293), .D(n9292), .Y(n11434) );
  INVX8 U4723 ( .A(n11434), .Y(n10657) );
  AND2X2 U4724 ( .A(n3884), .B(net103354), .Y(n4171) );
  OA22X4 U4725 ( .A0(n5296), .A1(n2989), .B0(n5249), .B1(n548), .Y(n9700) );
  OA22X4 U4726 ( .A0(n5296), .A1(n629), .B0(n5249), .B1(n2981), .Y(n9705) );
  OA22X4 U4727 ( .A0(n5296), .A1(n2134), .B0(n5249), .B1(n549), .Y(n9695) );
  OA22X2 U4728 ( .A0(n5296), .A1(n760), .B0(n5249), .B1(n2321), .Y(n9690) );
  OA22XL U4729 ( .A0(n5296), .A1(n1849), .B0(n5249), .B1(n3505), .Y(n9714) );
  OA22XL U4730 ( .A0(n5296), .A1(n1850), .B0(n5249), .B1(n3506), .Y(n9719) );
  XOR2X4 U4731 ( .A(n10330), .B(ICACHE_addr[20]), .Y(n10549) );
  OAI2BB2X1 U4732 ( .B0(\i_MIPS/n205 ), .B1(net108192), .A0N(n10556), .A1N(
        n5545), .Y(\i_MIPS/N48 ) );
  OAI221X4 U4733 ( .A0(\i_MIPS/ALUin1[20] ), .A1(net112364), .B0(
        \i_MIPS/ALUin1[21] ), .B1(net112346), .C0(n6682), .Y(n9341) );
  CLKMX2X4 U4734 ( .A(n9341), .B(n8549), .S0(net107798), .Y(n8873) );
  OA22X2 U4735 ( .A0(n4924), .A1(n1772), .B0(n4955), .B1(n3402), .Y(n6410) );
  OA22X2 U4736 ( .A0(n4924), .A1(n1469), .B0(n4950), .B1(n3043), .Y(n6416) );
  OA22X4 U4737 ( .A0(n5119), .A1(n2741), .B0(n5076), .B1(n1281), .Y(n9918) );
  OA22X4 U4738 ( .A0(n5119), .A1(n2742), .B0(n5080), .B1(n1282), .Y(n9913) );
  OA22X4 U4739 ( .A0(n5119), .A1(n2743), .B0(n5060), .B1(n1283), .Y(n9923) );
  OA22X2 U4740 ( .A0(n5122), .A1(n1470), .B0(n5077), .B1(n3044), .Y(n10106) );
  AO22X2 U4741 ( .A0(mem_rdata_I[76]), .A1(n5539), .B0(n249), .B1(n11262), .Y(
        n9769) );
  AO22X2 U4742 ( .A0(mem_rdata_I[48]), .A1(n5539), .B0(n251), .B1(n11234), .Y(
        n9732) );
  AO22X2 U4743 ( .A0(mem_rdata_I[80]), .A1(n5539), .B0(n253), .B1(n11266), .Y(
        n9722) );
  AO22X2 U4744 ( .A0(mem_rdata_I[16]), .A1(n5539), .B0(n252), .B1(n11202), .Y(
        n9727) );
  OAI32X4 U4745 ( .A0(n10858), .A1(n10857), .A2(net138001), .B0(
        \i_MIPS/PC/n33 ), .B1(net97444), .Y(n10862) );
  AO22X1 U4746 ( .A0(n4315), .A1(n11175), .B0(net112406), .B1(n11174), .Y(
        \i_MIPS/N75 ) );
  AO22X1 U4747 ( .A0(n4315), .A1(n10348), .B0(net112406), .B1(
        \i_MIPS/IR_ID[27] ), .Y(\i_MIPS/N85 ) );
  OAI2BB2XL U4748 ( .B0(\i_MIPS/n241 ), .B1(net108190), .A0N(n4315), .A1N(
        n11109), .Y(\i_MIPS/N95 ) );
  OAI2BB2XL U4749 ( .B0(\i_MIPS/n188 ), .B1(net108198), .A0N(n11161), .A1N(
        n4315), .Y(\i_MIPS/N31 ) );
  OAI2BB2XL U4750 ( .B0(\i_MIPS/n193 ), .B1(net108198), .A0N(n10814), .A1N(
        n4315), .Y(\i_MIPS/N36 ) );
  OAI2BB2XL U4751 ( .B0(\i_MIPS/n201 ), .B1(net108194), .A0N(n10505), .A1N(
        n4315), .Y(\i_MIPS/N44 ) );
  OAI2BB2XL U4752 ( .B0(\i_MIPS/n163 ), .B1(net108194), .A0N(n4315), .A1N(
        n10393), .Y(\i_MIPS/N103 ) );
  OAI2BB2XL U4753 ( .B0(\i_MIPS/n176 ), .B1(net108194), .A0N(n4315), .A1N(
        n2649), .Y(\i_MIPS/N116 ) );
  OAI2BB2XL U4754 ( .B0(\i_MIPS/n219 ), .B1(net108198), .A0N(n4315), .A1N(
        n11092), .Y(\i_MIPS/N62 ) );
  OAI2BB2XL U4755 ( .B0(\i_MIPS/n221 ), .B1(net108198), .A0N(n4315), .A1N(
        n10368), .Y(\i_MIPS/N64 ) );
  BUFX20 U4756 ( .A(n3915), .Y(n4072) );
  OA22X2 U4757 ( .A0(n10796), .A1(net108704), .B0(\i_MIPS/PC/n32 ), .B1(
        net108690), .Y(n10799) );
  AOI222X1 U4758 ( .A0(n5510), .A1(n11408), .B0(mem_rdata_D[58]), .B1(n233), 
        .C0(n12961), .C1(n5506), .Y(n10279) );
  AOI222X1 U4759 ( .A0(n5510), .A1(n11409), .B0(mem_rdata_D[59]), .B1(n233), 
        .C0(n12960), .C1(n5506), .Y(n10311) );
  AOI222X1 U4760 ( .A0(n5510), .A1(n11403), .B0(mem_rdata_D[53]), .B1(n232), 
        .C0(n12966), .C1(n5506), .Y(n10677) );
  AOI222X1 U4761 ( .A0(n5510), .A1(n11412), .B0(mem_rdata_D[62]), .B1(n235), 
        .C0(n12957), .C1(n5506), .Y(n10149) );
  OA22X4 U4762 ( .A0(n4974), .A1(n2136), .B0(n5019), .B1(n551), .Y(n8301) );
  OA22X2 U4763 ( .A0(n4914), .A1(n761), .B0(n4947), .B1(n2322), .Y(n8302) );
  OAI221X2 U4764 ( .A0(\i_MIPS/ALUin1[20] ), .A1(n4668), .B0(
        \i_MIPS/ALUin1[21] ), .B1(n3828), .C0(n8154), .Y(n9050) );
  OAI221X4 U4765 ( .A0(net112304), .A1(n7685), .B0(n7413), .B1(net101257), 
        .C0(net112420), .Y(n7416) );
  OAI22X1 U4766 ( .A0(n5110), .A1(n1446), .B0(n5079), .B1(n3015), .Y(n4346) );
  NAND2BX2 U4767 ( .AN(n4247), .B(n11296), .Y(n9613) );
  OAI221X2 U4768 ( .A0(n5624), .A1(\i_MIPS/n293 ), .B0(n3837), .B1(n5625), 
        .C0(\i_MIPS/n363 ), .Y(n6505) );
  NAND2XL U4769 ( .A(n8949), .B(n8948), .Y(n8950) );
  OA21X4 U4770 ( .A0(n7490), .A1(n7478), .B0(n8949), .Y(n7479) );
  OAI2BB1X4 U4771 ( .A0N(n8450), .A1N(n11181), .B0(n8433), .Y(n8173) );
  NAND4X4 U4772 ( .A(n7750), .B(n7749), .C(n7748), .D(n7747), .Y(n11363) );
  OA22X4 U4773 ( .A0(n10736), .A1(n4245), .B0(n10739), .B1(n4246), .Y(n7755)
         );
  INVX8 U4774 ( .A(n11363), .Y(n10736) );
  OAI221X2 U4775 ( .A0(net104582), .A1(net111624), .B0(net104583), .B1(
        net111636), .C0(net104584), .Y(net97815) );
  AO22X1 U4776 ( .A0(n4720), .A1(n986), .B0(n4719), .B1(n2506), .Y(n9209) );
  AO22X1 U4777 ( .A0(n4720), .A1(n987), .B0(n4719), .B1(n2507), .Y(n9200) );
  AO22X4 U4778 ( .A0(n4723), .A1(n447), .B0(n4719), .B1(n2030), .Y(n9105) );
  AO22X4 U4779 ( .A0(n4723), .A1(n448), .B0(n4719), .B1(n2031), .Y(n9096) );
  AO22X4 U4780 ( .A0(n4723), .A1(n470), .B0(n4719), .B1(n2057), .Y(n9008) );
  AO22X4 U4781 ( .A0(n4720), .A1(n471), .B0(n4719), .B1(n2058), .Y(n8999) );
  INVXL U4782 ( .A(net101465), .Y(n3902) );
  CLKINVX1 U4783 ( .A(n3902), .Y(n3903) );
  OA22X2 U4784 ( .A0(n4976), .A1(n738), .B0(n5025), .B1(n2297), .Y(n7433) );
  NAND4X4 U4785 ( .A(n7436), .B(n7435), .C(n7434), .D(n7433), .Y(n11362) );
  MX2XL U4786 ( .A(DCACHE_addr[22]), .B(n16), .S0(n208), .Y(\i_MIPS/n445 ) );
  NAND4X2 U4787 ( .A(n6210), .B(n6209), .C(n6208), .D(n6207), .Y(n11216) );
  NAND4X4 U4788 ( .A(n6287), .B(n6286), .C(n6285), .D(n6284), .Y(n10346) );
  OA22X4 U4789 ( .A0(n8353), .A1(n7815), .B0(n9158), .B1(n4659), .Y(n7700) );
  AO22X4 U4790 ( .A0(n9486), .A1(net100585), .B0(n9155), .B1(n9154), .Y(n9156)
         );
  NAND2X6 U4791 ( .A(\i_MIPS/ALUin1[19] ), .B(n6572), .Y(n9268) );
  AND4X4 U4792 ( .A(n6487), .B(n6489), .C(n6488), .D(n4658), .Y(n3908) );
  OA21X4 U4793 ( .A0(\i_MIPS/ALUin1[15] ), .A1(net112368), .B0(n8068), .Y(
        n6852) );
  NAND3BX2 U4794 ( .AN(n4473), .B(n8068), .C(n8067), .Y(n8438) );
  MX2XL U4795 ( .A(n12936), .B(n3902), .S0(n213), .Y(\i_MIPS/n446 ) );
  OA22XL U4796 ( .A0(n5295), .A1(n1851), .B0(n5248), .B1(n3507), .Y(n9680) );
  OA22XL U4797 ( .A0(n5295), .A1(n1852), .B0(n5248), .B1(n3508), .Y(n9670) );
  OA22X4 U4798 ( .A0(n5295), .A1(n2993), .B0(n5248), .B1(n1435), .Y(n9650) );
  AO22X4 U4799 ( .A0(mem_rdata_I[32]), .A1(n5543), .B0(n249), .B1(n11218), .Y(
        n6156) );
  AO22X4 U4800 ( .A0(mem_rdata_I[64]), .A1(n5543), .B0(n250), .B1(n11250), .Y(
        n6146) );
  AO22X1 U4801 ( .A0(n4722), .A1(n299), .B0(n4719), .B1(n2447), .Y(n7593) );
  AO22X4 U4802 ( .A0(n4722), .A1(n287), .B0(n4719), .B1(n2032), .Y(n7674) );
  AO22X4 U4803 ( .A0(n4722), .A1(n288), .B0(n4719), .B1(n2033), .Y(n7665) );
  AO22X4 U4804 ( .A0(n4722), .A1(n293), .B0(n4719), .B1(n2063), .Y(n7202) );
  AO22X4 U4805 ( .A0(n4721), .A1(n294), .B0(n4719), .B1(n2064), .Y(n7211) );
  NOR4X2 U4806 ( .A(n7595), .B(n7594), .C(n7593), .D(n7592), .Y(n7596) );
  NAND2X2 U4807 ( .A(\i_MIPS/ALUin1[7] ), .B(net112356), .Y(n7695) );
  INVX20 U4808 ( .A(n5556), .Y(n4655) );
  INVX12 U4809 ( .A(n3952), .Y(mem_wdata_I[14]) );
  MX2XL U4810 ( .A(n3602), .B(n3909), .S0(n208), .Y(\i_MIPS/n397 ) );
  CLKAND2X12 U4811 ( .A(n5557), .B(n11186), .Y(mem_wdata_I[0]) );
  NAND4X4 U4812 ( .A(n6150), .B(n6149), .C(n6148), .D(n6147), .Y(n11186) );
  NAND4X4 U4813 ( .A(n6927), .B(n6926), .C(n6925), .D(n6924), .Y(n11448) );
  INVX8 U4814 ( .A(n11448), .Y(n10928) );
  OAI2BB2X4 U4815 ( .B0(n8347), .B1(n4660), .A0N(n8349), .A1N(n8348), .Y(n8355) );
  MXI2X4 U4816 ( .A(n10900), .B(n10899), .S0(n5520), .Y(n10901) );
  INVX6 U4817 ( .A(n11358), .Y(n10899) );
  OA22X1 U4818 ( .A0(n6495), .A1(net133688), .B0(net133688), .B1(n6494), .Y(
        n6498) );
  NAND4X4 U4819 ( .A(n8594), .B(n8593), .C(n8592), .D(n8591), .Y(n11433) );
  INVX8 U4820 ( .A(n11395), .Y(n10739) );
  NAND4X4 U4821 ( .A(n7754), .B(n7753), .C(n7752), .D(n7751), .Y(n11395) );
  MX2XL U4822 ( .A(n3607), .B(net98044), .S0(n213), .Y(\i_MIPS/n411 ) );
  AO22X4 U4823 ( .A0(n5537), .A1(ICACHE_addr[20]), .B0(n240), .B1(n11335), .Y(
        n11133) );
  AO22X4 U4824 ( .A0(n5537), .A1(ICACHE_addr[11]), .B0(n239), .B1(n11326), .Y(
        n11142) );
  AO22X4 U4825 ( .A0(n5537), .A1(ICACHE_addr[15]), .B0(n239), .B1(n11330), .Y(
        n11140) );
  AO22X4 U4826 ( .A0(n5537), .A1(ICACHE_addr[9]), .B0(n239), .B1(n11324), .Y(
        n11143) );
  AO22X4 U4827 ( .A0(n5537), .A1(ICACHE_addr[22]), .B0(n240), .B1(n11337), .Y(
        n11139) );
  AO22X4 U4828 ( .A0(n5537), .A1(ICACHE_addr[13]), .B0(n240), .B1(n11328), .Y(
        n11149) );
  AO22X4 U4829 ( .A0(n5537), .A1(ICACHE_addr[7]), .B0(n239), .B1(n11322), .Y(
        n11136) );
  AO22X4 U4830 ( .A0(n5537), .A1(ICACHE_addr[10]), .B0(n239), .B1(n11325), .Y(
        n11141) );
  AO22X4 U4831 ( .A0(n5537), .A1(ICACHE_addr[14]), .B0(n240), .B1(n11329), .Y(
        n11147) );
  AO22X4 U4832 ( .A0(n5537), .A1(ICACHE_addr[27]), .B0(n240), .B1(n11342), .Y(
        n11138) );
  OA22X1 U4833 ( .A0(n5211), .A1(n1648), .B0(n5168), .B1(n3230), .Y(n9995) );
  NAND2BX4 U4834 ( .AN(n4247), .B(n11290), .Y(n10016) );
  OAI221X2 U4835 ( .A0(n8826), .A1(net111622), .B0(n8825), .B1(net111634), 
        .C0(n8824), .Y(n10507) );
  NAND4X2 U4836 ( .A(n8312), .B(n8311), .C(n8310), .D(n8309), .Y(n11406) );
  NAND2XL U4837 ( .A(n10785), .B(n5520), .Y(n4234) );
  INVX8 U4838 ( .A(\i_MIPS/ALUin1[28] ), .Y(n7149) );
  AOI33X2 U4839 ( .A0(net112292), .A1(n9168), .A2(n9148), .B0(n9147), .B1(
        n9150), .B2(net137952), .Y(n9178) );
  NAND3BX4 U4840 ( .AN(n6777), .B(n6776), .C(n6775), .Y(net97703) );
  OA22X1 U4841 ( .A0(n4824), .A1(n1216), .B0(n4869), .B1(n2753), .Y(n7937) );
  AOI222X2 U4842 ( .A0(n5499), .A1(n11421), .B0(mem_rdata_D[71]), .B1(n232), 
        .C0(n12980), .C1(n5497), .Y(n10885) );
  NAND2X1 U4843 ( .A(n10791), .B(net112404), .Y(n10852) );
  NAND4X4 U4844 ( .A(n8801), .B(n8800), .C(n8799), .D(n8798), .Y(n11400) );
  AOI222X2 U4845 ( .A0(n5505), .A1(n11379), .B0(mem_rdata_D[29]), .B1(n236), 
        .C0(n12958), .C1(n5502), .Y(n10688) );
  NAND4X2 U4846 ( .A(n8198), .B(n8197), .C(n8196), .D(n8195), .Y(n11379) );
  AOI33X2 U4847 ( .A0(net112292), .A1(n9494), .A2(n9493), .B0(net137952), .B1(
        n9492), .B2(n9491), .Y(n9495) );
  OAI222X4 U4848 ( .A0(n9463), .A1(n9053), .B0(n9052), .B1(net112420), .C0(
        n9469), .C1(n9051), .Y(n9062) );
  AO22X2 U4849 ( .A0(n9056), .A1(net100585), .B0(n9055), .B1(n9054), .Y(n9061)
         );
  OAI211X4 U4850 ( .A0(n9342), .A1(n9050), .B0(n9049), .C0(n9048), .Y(n9063)
         );
  AOI222X1 U4851 ( .A0(n5511), .A1(n11394), .B0(mem_rdata_D[44]), .B1(n232), 
        .C0(n12975), .C1(n5507), .Y(n10729) );
  INVX8 U4852 ( .A(n11394), .Y(n10728) );
  NAND4X6 U4853 ( .A(n7440), .B(n7439), .C(n7438), .D(n7437), .Y(n11394) );
  AOI222X1 U4854 ( .A0(n5495), .A1(n11465), .B0(mem_rdata_D[115]), .B1(n232), 
        .C0(n5494), .C1(n12968), .Y(n10992) );
  NAND4X2 U4855 ( .A(n8590), .B(n8589), .C(n8588), .D(n8587), .Y(n11465) );
  OAI31X2 U4856 ( .A0(n6525), .A1(n6524), .A2(n6523), .B0(n6522), .Y(n3910) );
  OAI211X4 U4857 ( .A0(n6521), .A1(n6520), .B0(n8947), .C0(n9040), .Y(n6523)
         );
  INVXL U4858 ( .A(n11505), .Y(n4625) );
  NAND4X4 U4859 ( .A(n7660), .B(n7659), .C(n7658), .D(n7657), .Y(n11396) );
  OAI211X2 U4860 ( .A0(net112304), .A1(net101554), .B0(net101555), .C0(
        net101556), .Y(net97753) );
  INVXL U4861 ( .A(n3721), .Y(n3911) );
  INVXL U4862 ( .A(net102938), .Y(n3912) );
  OAI221X2 U4863 ( .A0(n9325), .A1(net111622), .B0(n3913), .B1(net111634), 
        .C0(n9324), .Y(n10653) );
  INVXL U4864 ( .A(n8526), .Y(n3914) );
  MX2XL U4865 ( .A(\i_MIPS/EX_MEM[6] ), .B(n3912), .S0(n216), .Y(\i_MIPS/n468 ) );
  INVX3 U4866 ( .A(n8555), .Y(n8731) );
  AO22X4 U4867 ( .A0(n4723), .A1(n449), .B0(n4719), .B1(n2035), .Y(n8507) );
  AO22X4 U4868 ( .A0(n4723), .A1(n416), .B0(n4719), .B1(n1977), .Y(n8609) );
  AO22X4 U4869 ( .A0(n4723), .A1(n450), .B0(n4719), .B1(n2036), .Y(n8815) );
  NOR4X2 U4870 ( .A(n8518), .B(n8517), .C(n8516), .D(n8515), .Y(n8519) );
  MX2XL U4871 ( .A(n12933), .B(n3911), .S0(n217), .Y(\i_MIPS/n443 ) );
  NAND4X4 U4872 ( .A(n7852), .B(n7851), .C(n7850), .D(n7849), .Y(n11399) );
  OA22X2 U4873 ( .A0(n4977), .A1(n665), .B0(n4999), .B1(n2235), .Y(n7849) );
  BUFX20 U4874 ( .A(net112002), .Y(net112004) );
  NOR4X2 U4875 ( .A(n8006), .B(n8005), .C(n8004), .D(n8003), .Y(n8007) );
  OA22X4 U4876 ( .A0(n5296), .A1(n2137), .B0(n5240), .B1(n552), .Y(n6100) );
  OA22X4 U4877 ( .A0(n10475), .A1(n4675), .B0(n10478), .B1(n4250), .Y(n8504)
         );
  MX2XL U4878 ( .A(n12942), .B(net97995), .S0(n213), .Y(\i_MIPS/n452 ) );
  OA22X4 U4879 ( .A0(n4836), .A1(n3369), .B0(n4882), .B1(n1740), .Y(n6333) );
  AOI33X2 U4880 ( .A0(net112292), .A1(n9283), .A2(n9282), .B0(net111994), .B1(
        n9281), .B2(n4251), .Y(n9284) );
  AND3X6 U4881 ( .A(n10375), .B(net97444), .C(net97592), .Y(n3915) );
  OAI2BB2X1 U4882 ( .B0(\i_MIPS/n231 ), .B1(net108198), .A0N(n5545), .A1N(
        net98496), .Y(\i_MIPS/N79 ) );
  BUFX12 U4883 ( .A(n5134), .Y(n5125) );
  AOI222X4 U4884 ( .A0(n5512), .A1(n11382), .B0(mem_rdata_D[32]), .B1(n232), 
        .C0(n12987), .C1(n5507), .Y(n10963) );
  OAI2BB2X1 U4885 ( .B0(\i_MIPS/n235 ), .B1(net108198), .A0N(n4072), .A1N(
        n10840), .Y(\i_MIPS/N83 ) );
  AO22X4 U4886 ( .A0(mem_rdata_I[116]), .A1(n5541), .B0(n252), .B1(n11302), 
        .Y(n9619) );
  AO22X4 U4887 ( .A0(mem_rdata_I[110]), .A1(n5541), .B0(n249), .B1(n11296), 
        .Y(n9594) );
  AO22X4 U4888 ( .A0(mem_rdata_I[61]), .A1(n5541), .B0(n251), .B1(n11247), .Y(
        n6236) );
  NAND4X4 U4889 ( .A(n9178), .B(n9177), .C(n9176), .D(n9175), .Y(n10665) );
  CLKINVX8 U4890 ( .A(n9180), .Y(n10679) );
  AND2X8 U4891 ( .A(\i_MIPS/ID_EX[79] ), .B(net102253), .Y(n4476) );
  NAND4X4 U4892 ( .A(n8695), .B(n8694), .C(n8693), .D(n8692), .Y(n11359) );
  OA22X2 U4893 ( .A0(n4746), .A1(n2409), .B0(n4790), .B1(n847), .Y(n8695) );
  INVX8 U4894 ( .A(n11359), .Y(n10701) );
  NAND2X4 U4895 ( .A(net107794), .B(n9170), .Y(n9342) );
  NAND4X2 U4896 ( .A(n8012), .B(n8011), .C(n8010), .D(n8009), .Y(n11447) );
  OA22X4 U4897 ( .A0(n10905), .A1(n4676), .B0(n10908), .B1(n4250), .Y(n8026)
         );
  NAND2X4 U4898 ( .A(\i_MIPS/ALUin1[27] ), .B(n6592), .Y(n9329) );
  OA22X4 U4899 ( .A0(n4834), .A1(n2138), .B0(n4879), .B1(n553), .Y(n6417) );
  OA22X4 U4900 ( .A0(n4834), .A1(n2996), .B0(n4879), .B1(n554), .Y(n6411) );
  CLKBUFX8 U4901 ( .A(n4845), .Y(n4834) );
  OA22X1 U4902 ( .A0(n4922), .A1(n1083), .B0(n4249), .B1(n2676), .Y(n7090) );
  BUFX2 U4903 ( .A(n4927), .Y(n4922) );
  OA22X1 U4904 ( .A0(n4978), .A1(n1217), .B0(n5023), .B1(n2754), .Y(n7837) );
  OA22X2 U4905 ( .A0(n10763), .A1(n4676), .B0(n10766), .B1(n4250), .Y(n7854)
         );
  MXI2X4 U4906 ( .A(n10947), .B(n10946), .S0(n5522), .Y(n10948) );
  OAI31X4 U4907 ( .A0(\i_MIPS/ALUin1[30] ), .A1(n11180), .A2(n11179), .B0(
        n11178), .Y(n11547) );
  INVXL U4908 ( .A(n11177), .Y(n11179) );
  AOI2BB1X4 U4909 ( .A0N(n7483), .A1N(net103914), .B0(n4337), .Y(n7484) );
  OA22X4 U4910 ( .A0(n10215), .A1(n4245), .B0(n10218), .B1(n4246), .Y(n9513)
         );
  AND3X8 U4911 ( .A(n4129), .B(n3919), .C(n3920), .Y(net102781) );
  XNOR2X4 U4912 ( .A(n4132), .B(n4127), .Y(n3919) );
  AO22X4 U4913 ( .A0(mem_rdata_I[106]), .A1(n5537), .B0(n251), .B1(n11292), 
        .Y(n10044) );
  AO22X4 U4914 ( .A0(mem_rdata_I[104]), .A1(n5537), .B0(n251), .B1(n11290), 
        .Y(n9997) );
  AO22X4 U4915 ( .A0(mem_rdata_I[9]), .A1(n5537), .B0(n253), .B1(n11195), .Y(
        n10031) );
  AO22X4 U4916 ( .A0(mem_rdata_I[73]), .A1(n5537), .B0(n251), .B1(n11259), .Y(
        n10026) );
  AO22X4 U4917 ( .A0(mem_rdata_I[105]), .A1(n5537), .B0(n249), .B1(n11291), 
        .Y(n10021) );
  AO22X4 U4918 ( .A0(mem_rdata_I[41]), .A1(n5537), .B0(n252), .B1(n11227), .Y(
        n10035) );
  AO22X4 U4919 ( .A0(mem_rdata_I[72]), .A1(n5537), .B0(n250), .B1(n11258), .Y(
        n10002) );
  NAND2BX4 U4920 ( .AN(n4247), .B(n11289), .Y(n10135) );
  AOI2BB1X2 U4921 ( .A0N(n3676), .A1N(n10539), .B0(n4071), .Y(n10541) );
  CLKINVX8 U4922 ( .A(n9075), .Y(n10467) );
  OAI222X4 U4923 ( .A0(\i_MIPS/PC/n26 ), .A1(net108688), .B0(net97445), .B1(
        n10456), .C0(n4410), .C1(net108704), .Y(n10462) );
  OAI222X4 U4924 ( .A0(n3784), .A1(net108688), .B0(net97445), .B1(n11110), 
        .C0(n4408), .C1(net108702), .Y(n11115) );
  NAND3BX4 U4925 ( .AN(n11115), .B(n11114), .C(n11113), .Y(\i_MIPS/PC/n38 ) );
  CLKMX2X2 U4926 ( .A(\D_cache/cache[7][69] ), .B(n10989), .S0(n5009), .Y(
        \D_cache/n1237 ) );
  CLKMX2X2 U4927 ( .A(\D_cache/cache[6][69] ), .B(n10989), .S0(n4965), .Y(
        \D_cache/n1238 ) );
  CLKMX2X2 U4928 ( .A(\D_cache/cache[5][69] ), .B(n10989), .S0(n4944), .Y(
        \D_cache/n1239 ) );
  CLKMX2X2 U4929 ( .A(\D_cache/cache[4][69] ), .B(n10989), .S0(n4901), .Y(
        \D_cache/n1240 ) );
  CLKMX2X2 U4930 ( .A(\D_cache/cache[3][69] ), .B(n10989), .S0(n4855), .Y(
        \D_cache/n1241 ) );
  CLKMX2X2 U4931 ( .A(\D_cache/cache[2][69] ), .B(n10989), .S0(n4808), .Y(
        \D_cache/n1242 ) );
  CLKMX2X2 U4932 ( .A(\D_cache/cache[1][69] ), .B(n10989), .S0(n4786), .Y(
        \D_cache/n1243 ) );
  MX2X1 U4933 ( .A(\D_cache/cache[0][69] ), .B(n10989), .S0(n4739), .Y(
        \D_cache/n1244 ) );
  CLKMX2X2 U4934 ( .A(\D_cache/cache[2][51] ), .B(n10997), .S0(n4809), .Y(
        \D_cache/n1386 ) );
  CLKMX2X2 U4935 ( .A(\D_cache/cache[3][51] ), .B(n10997), .S0(n4855), .Y(
        \D_cache/n1385 ) );
  CLKMX2X2 U4936 ( .A(\D_cache/cache[4][51] ), .B(n10997), .S0(n4901), .Y(
        \D_cache/n1384 ) );
  CLKMX2X2 U4937 ( .A(\D_cache/cache[5][51] ), .B(n10997), .S0(n4944), .Y(
        \D_cache/n1383 ) );
  CLKMX2X2 U4938 ( .A(\D_cache/cache[6][51] ), .B(n10997), .S0(n4965), .Y(
        \D_cache/n1382 ) );
  CLKMX2X2 U4939 ( .A(\D_cache/cache[7][51] ), .B(n10997), .S0(n5009), .Y(
        \D_cache/n1381 ) );
  INVX20 U4940 ( .A(net108708), .Y(net108704) );
  NAND3BX4 U4941 ( .AN(n10590), .B(n10589), .C(n10588), .Y(\i_MIPS/PC/n43 ) );
  OAI222X4 U4942 ( .A0(\i_MIPS/PC/n25 ), .A1(net108688), .B0(net97445), .B1(
        net98497), .C0(net129017), .C1(net108704), .Y(n4143) );
  AOI222X1 U4943 ( .A0(n5511), .A1(n11391), .B0(mem_rdata_D[41]), .B1(n234), 
        .C0(n12978), .C1(n5507), .Y(n10705) );
  AND4X8 U4944 ( .A(n8528), .B(n8531), .C(n8530), .D(n8529), .Y(net129200) );
  NAND4BX4 U4945 ( .AN(n4347), .B(n9502), .C(n9501), .D(n9500), .Y(n11468) );
  INVX8 U4946 ( .A(n11468), .Y(n10209) );
  INVXL U4947 ( .A(n8740), .Y(n6492) );
  OAI2BB2X1 U4948 ( .B0(\i_MIPS/n202 ), .B1(net108192), .A0N(n10650), .A1N(
        n4315), .Y(\i_MIPS/N45 ) );
  OAI2BB2X1 U4949 ( .B0(\i_MIPS/n204 ), .B1(net108192), .A0N(n11121), .A1N(
        n4315), .Y(\i_MIPS/N47 ) );
  AO22X4 U4950 ( .A0(mem_rdata_I[42]), .A1(n5543), .B0(n253), .B1(n11228), .Y(
        n10059) );
  AO22X4 U4951 ( .A0(mem_rdata_I[10]), .A1(n5543), .B0(n250), .B1(n11196), .Y(
        n10054) );
  AO22X4 U4952 ( .A0(mem_rdata_I[102]), .A1(n5535), .B0(n253), .B1(n11288), 
        .Y(n10092) );
  AO22X4 U4953 ( .A0(mem_rdata_I[103]), .A1(n5543), .B0(n249), .B1(n11289), 
        .Y(n10116) );
  AO22X4 U4954 ( .A0(mem_rdata_I[71]), .A1(n5543), .B0(n249), .B1(n11257), .Y(
        n10121) );
  AO22X4 U4955 ( .A0(mem_rdata_I[38]), .A1(n5543), .B0(n252), .B1(n11224), .Y(
        n10107) );
  AO22X4 U4956 ( .A0(mem_rdata_I[6]), .A1(n5544), .B0(n250), .B1(n11192), .Y(
        n10102) );
  AO22X4 U4957 ( .A0(mem_rdata_I[70]), .A1(n5543), .B0(n253), .B1(n11256), .Y(
        n10097) );
  AO22X4 U4958 ( .A0(mem_rdata_I[74]), .A1(n5541), .B0(n250), .B1(n11260), .Y(
        n10049) );
  OAI21X1 U4959 ( .A0(\i_MIPS/n184 ), .A1(net108190), .B0(n10529), .Y(
        \i_MIPS/N27 ) );
  NAND2X4 U4960 ( .A(\i_MIPS/PC_o[1] ), .B(n5545), .Y(n10529) );
  OA22X4 U4961 ( .A0(n4926), .A1(n3000), .B0(n4950), .B1(n558), .Y(n6348) );
  NAND4X4 U4962 ( .A(n8789), .B(n8788), .C(n8787), .D(n8786), .Y(n11464) );
  OA22XL U4963 ( .A0(n4746), .A1(n1292), .B0(n4789), .B1(n2823), .Y(n8789) );
  NAND4X4 U4964 ( .A(n10125), .B(n10124), .C(n10123), .D(n10122), .Y(n11193)
         );
  OA22X1 U4965 ( .A0(n5304), .A1(n1218), .B0(n5259), .B1(n2755), .Y(n10123) );
  AO22X4 U4966 ( .A0(mem_rdata_I[7]), .A1(n5535), .B0(n251), .B1(n11193), .Y(
        n10126) );
  NAND2X8 U4967 ( .A(net101906), .B(net107798), .Y(net103060) );
  INVX6 U4968 ( .A(net107808), .Y(net107798) );
  MX2XL U4969 ( .A(\i_MIPS/ID_EX[69] ), .B(n262), .S0(n216), .Y(\i_MIPS/n381 )
         );
  OA22X4 U4970 ( .A0(n10481), .A1(n4245), .B0(n10484), .B1(n4246), .Y(n8503)
         );
  NOR4X2 U4971 ( .A(n6626), .B(n6625), .C(n6624), .D(n6623), .Y(n6627) );
  AO22X1 U4972 ( .A0(n4721), .A1(n423), .B0(n4719), .B1(n2002), .Y(n6624) );
  NAND4X4 U4973 ( .A(n9778), .B(n9777), .C(n9776), .D(n9775), .Y(n11230) );
  NAND2BX2 U4974 ( .AN(n5430), .B(n11230), .Y(n9780) );
  AO22X4 U4975 ( .A0(n4723), .A1(n451), .B0(n4719), .B1(n2037), .Y(n8806) );
  AO22X4 U4976 ( .A0(n4723), .A1(n473), .B0(n4719), .B1(n2065), .Y(n8417) );
  AO22X4 U4977 ( .A0(n4723), .A1(n452), .B0(n4719), .B1(n2038), .Y(n8408) );
  AO22X4 U4978 ( .A0(n4723), .A1(n453), .B0(n4719), .B1(n2039), .Y(n8317) );
  AO22X4 U4979 ( .A0(n4723), .A1(n454), .B0(n4719), .B1(n2040), .Y(n8713) );
  OA22X4 U4980 ( .A0(n7984), .A1(net103060), .B0(n7983), .B1(n7982), .Y(n7985)
         );
  MXI2X4 U4981 ( .A(\i_MIPS/ID_EX[112] ), .B(\i_MIPS/ID_EX[85] ), .S0(
        \i_MIPS/ID_EX_5 ), .Y(n6606) );
  AO21X4 U4982 ( .A0(net103354), .A1(net104866), .B0(net105012), .Y(net101771)
         );
  AND2X4 U4983 ( .A(n4671), .B(\i_MIPS/n356 ), .Y(n4464) );
  AOI222X2 U4984 ( .A0(n5504), .A1(n11378), .B0(mem_rdata_D[28]), .B1(n235), 
        .C0(n12959), .C1(n5501), .Y(n10482) );
  OA22X1 U4985 ( .A0(n4831), .A1(n1219), .B0(n4876), .B1(n2756), .Y(n6938) );
  NAND2BX1 U4986 ( .AN(n8956), .B(n8957), .Y(n8962) );
  INVXL U4987 ( .A(n8630), .Y(n7521) );
  AO22X4 U4988 ( .A0(n4722), .A1(n474), .B0(n4719), .B1(n2066), .Y(n7960) );
  NOR4X4 U4989 ( .A(n8040), .B(n8039), .C(n8038), .D(n8037), .Y(n8041) );
  INVX3 U4990 ( .A(n10152), .Y(n8604) );
  OA22X2 U4991 ( .A0(n5210), .A1(n1471), .B0(n5167), .B1(n3045), .Y(n9960) );
  OA22X2 U4992 ( .A0(n5301), .A1(n1472), .B0(n5247), .B1(n3046), .Y(n9959) );
  INVX8 U4993 ( .A(n11367), .Y(n10769) );
  NAND4X4 U4994 ( .A(n7848), .B(n7847), .C(n7846), .D(n7845), .Y(n11367) );
  CLKMX2X2 U4995 ( .A(\D_cache/cache[7][87] ), .B(n10951), .S0(n5008), .Y(
        \D_cache/n1093 ) );
  CLKMX2X2 U4996 ( .A(\D_cache/cache[6][87] ), .B(n10951), .S0(n4964), .Y(
        \D_cache/n1094 ) );
  CLKMX2X2 U4997 ( .A(\D_cache/cache[5][87] ), .B(n10951), .S0(n4943), .Y(
        \D_cache/n1095 ) );
  CLKMX2X2 U4998 ( .A(\D_cache/cache[4][87] ), .B(n10951), .S0(n4900), .Y(
        \D_cache/n1096 ) );
  CLKMX2X2 U4999 ( .A(\D_cache/cache[3][87] ), .B(n10951), .S0(n4854), .Y(
        \D_cache/n1097 ) );
  CLKMX2X2 U5000 ( .A(\D_cache/cache[2][87] ), .B(n10951), .S0(n4809), .Y(
        \D_cache/n1098 ) );
  CLKMX2X2 U5001 ( .A(\D_cache/cache[1][87] ), .B(n10951), .S0(n4786), .Y(
        \D_cache/n1099 ) );
  MX2X1 U5002 ( .A(\D_cache/cache[0][87] ), .B(n10951), .S0(n4741), .Y(
        \D_cache/n1100 ) );
  MX2X1 U5003 ( .A(\D_cache/cache[4][64] ), .B(n10964), .S0(n4901), .Y(
        \D_cache/n1280 ) );
  CLKMX2X2 U5004 ( .A(\D_cache/cache[7][55] ), .B(n10945), .S0(n5008), .Y(
        \D_cache/n1349 ) );
  CLKMX2X2 U5005 ( .A(\D_cache/cache[6][55] ), .B(n10945), .S0(n4964), .Y(
        \D_cache/n1350 ) );
  CLKMX2X2 U5006 ( .A(\D_cache/cache[5][55] ), .B(n10945), .S0(n4943), .Y(
        \D_cache/n1351 ) );
  CLKMX2X2 U5007 ( .A(\D_cache/cache[4][55] ), .B(n10945), .S0(n4900), .Y(
        \D_cache/n1352 ) );
  CLKMX2X2 U5008 ( .A(\D_cache/cache[3][55] ), .B(n10945), .S0(n4854), .Y(
        \D_cache/n1353 ) );
  CLKMX2X2 U5009 ( .A(\D_cache/cache[2][55] ), .B(n10945), .S0(n4809), .Y(
        \D_cache/n1354 ) );
  CLKMX2X2 U5010 ( .A(\D_cache/cache[1][55] ), .B(n10945), .S0(n4778), .Y(
        \D_cache/n1355 ) );
  MX2X1 U5011 ( .A(\D_cache/cache[0][55] ), .B(n10945), .S0(n4741), .Y(
        \D_cache/n1356 ) );
  CLKMX2X2 U5012 ( .A(\D_cache/cache[7][32] ), .B(n10958), .S0(n5007), .Y(
        \D_cache/n1533 ) );
  CLKMX2X2 U5013 ( .A(\D_cache/cache[6][32] ), .B(n10958), .S0(n4963), .Y(
        \D_cache/n1534 ) );
  CLKMX2X2 U5014 ( .A(\D_cache/cache[5][32] ), .B(n10958), .S0(n4937), .Y(
        \D_cache/n1535 ) );
  CLKMX2X2 U5015 ( .A(\D_cache/cache[4][32] ), .B(n10958), .S0(n4899), .Y(
        \D_cache/n1536 ) );
  CLKMX2X2 U5016 ( .A(\D_cache/cache[3][32] ), .B(n10958), .S0(n4853), .Y(
        \D_cache/n1537 ) );
  CLKMX2X2 U5017 ( .A(\D_cache/cache[2][32] ), .B(n10958), .S0(n4808), .Y(
        \D_cache/n1538 ) );
  CLKMX2X2 U5018 ( .A(\D_cache/cache[1][32] ), .B(n10958), .S0(n4783), .Y(
        \D_cache/n1539 ) );
  MX2X1 U5019 ( .A(\D_cache/cache[0][32] ), .B(n10958), .S0(n4740), .Y(
        \D_cache/n1540 ) );
  NAND2X2 U5020 ( .A(n9475), .B(n8848), .Y(n8940) );
  NAND4X4 U5021 ( .A(n9745), .B(n9744), .C(n9743), .D(n9742), .Y(n11261) );
  OA22X2 U5022 ( .A0(n5297), .A1(n687), .B0(n5250), .B1(n2298), .Y(n9743) );
  AO21X4 U5023 ( .A0(n7875), .A1(n7874), .B0(n7873), .Y(n7889) );
  BUFX2 U5024 ( .A(n4929), .Y(n4920) );
  INVX1 U5025 ( .A(net102426), .Y(n4090) );
  AO21X4 U5026 ( .A0(n8850), .A1(n8849), .B0(n8861), .Y(net102554) );
  NAND3X2 U5027 ( .A(n9281), .B(net112294), .C(n9279), .Y(n9285) );
  INVX8 U5028 ( .A(n11385), .Y(n10923) );
  OA21X4 U5029 ( .A0(n7687), .A1(n7525), .B0(n7524), .Y(n7526) );
  CLKMX2X2 U5030 ( .A(\i_MIPS/ALUin1[29] ), .B(n10692), .S0(n222), .Y(
        \i_MIPS/n533 ) );
  NAND2X2 U5031 ( .A(\i_MIPS/ALUin1[29] ), .B(n6594), .Y(n11183) );
  AO21X4 U5032 ( .A0(n9331), .A1(n4662), .B0(n8355), .Y(n8547) );
  NOR2X2 U5033 ( .A(n4662), .B(n8654), .Y(n9055) );
  XNOR2X4 U5034 ( .A(n4100), .B(n5), .Y(n3923) );
  XNOR2X4 U5035 ( .A(n4099), .B(n4136), .Y(n3924) );
  OA22X1 U5036 ( .A0(n5123), .A1(n1649), .B0(n5077), .B1(n3231), .Y(n10120) );
  BUFX4 U5037 ( .A(n5125), .Y(n5123) );
  NAND4X4 U5038 ( .A(n10120), .B(n10119), .C(n10118), .D(n10117), .Y(n11257)
         );
  OA22X1 U5039 ( .A0(n5304), .A1(n1220), .B0(n5259), .B1(n2757), .Y(n10118) );
  INVX4 U5040 ( .A(n6334), .Y(n11012) );
  OAI222X4 U5041 ( .A0(\i_MIPS/PC/n17 ), .A1(net108688), .B0(net97445), .B1(
        n10425), .C0(n4400), .C1(net108704), .Y(n10430) );
  XOR2X2 U5042 ( .A(n10846), .B(ICACHE_addr[28]), .Y(n10849) );
  NAND2BX4 U5043 ( .AN(n10793), .B(ICACHE_addr[27]), .Y(n10846) );
  INVX6 U5044 ( .A(n10849), .Y(n10855) );
  AND2X1 U5045 ( .A(n11177), .B(n7481), .Y(n4454) );
  NAND2X2 U5046 ( .A(\i_MIPS/ALUin1[30] ), .B(n11180), .Y(n7481) );
  OA22X2 U5047 ( .A0(n11547), .A1(n11546), .B0(n4454), .B1(n11547), .Y(n4337)
         );
  CLKAND2X6 U5048 ( .A(\i_MIPS/ALUin1[4] ), .B(net127710), .Y(net127829) );
  NAND2X2 U5049 ( .A(n6977), .B(n4536), .Y(n9454) );
  NAND4X4 U5050 ( .A(n9755), .B(n9754), .C(n9753), .D(n9752), .Y(n11229) );
  OA22X2 U5051 ( .A0(n5297), .A1(n688), .B0(n5250), .B1(n2299), .Y(n9753) );
  XNOR2X4 U5052 ( .A(n3716), .B(n11498), .Y(n6413) );
  NOR4X8 U5053 ( .A(n8542), .B(n7800), .C(n3638), .D(n3662), .Y(n6557) );
  NAND2X8 U5054 ( .A(n6557), .B(n4393), .Y(n9269) );
  AO22X4 U5055 ( .A0(mem_rdata_I[111]), .A1(n5540), .B0(n250), .B1(n11297), 
        .Y(n9643) );
  OA22X2 U5056 ( .A0(n10725), .A1(n4245), .B0(n10728), .B1(n4246), .Y(n7441)
         );
  NAND4X4 U5057 ( .A(n6392), .B(n6391), .C(n6390), .D(n6389), .Y(n11484) );
  NAND2BX4 U5058 ( .AN(n4247), .B(n11283), .Y(n9969) );
  NAND4X2 U5059 ( .A(n6135), .B(n6134), .C(n6133), .D(n6132), .Y(n11283) );
  OA22X4 U5060 ( .A0(n10459), .A1(net133585), .B0(n10458), .B1(net108660), .Y(
        n10460) );
  BUFX12 U5061 ( .A(n4074), .Y(n3929) );
  OAI211X2 U5062 ( .A0(n4075), .A1(n4076), .B0(n4078), .C0(n4077), .Y(n4074)
         );
  NAND2XL U5063 ( .A(n7509), .B(n7503), .Y(n6848) );
  NOR2X6 U5064 ( .A(n7051), .B(n6968), .Y(n4420) );
  NAND4X2 U5065 ( .A(n6656), .B(n6655), .C(n6654), .D(n6653), .Y(n11413) );
  OA22XL U5066 ( .A0(n4985), .A1(n1127), .B0(n5031), .B1(n2658), .Y(n6653) );
  OA22X4 U5067 ( .A0(n4987), .A1(n2139), .B0(n5033), .B1(n559), .Y(n6381) );
  MX2X1 U5068 ( .A(\D_cache/cache[1][49] ), .B(n10768), .S0(n4783), .Y(
        \D_cache/n1403 ) );
  MX2X1 U5069 ( .A(\D_cache/cache[2][49] ), .B(n10768), .S0(n4805), .Y(
        \D_cache/n1402 ) );
  MX2X1 U5070 ( .A(\D_cache/cache[3][49] ), .B(n10768), .S0(n4849), .Y(
        \D_cache/n1401 ) );
  MX2X1 U5071 ( .A(\D_cache/cache[4][49] ), .B(n10768), .S0(n4894), .Y(
        \D_cache/n1400 ) );
  MX2X1 U5072 ( .A(\D_cache/cache[5][49] ), .B(n10768), .S0(n4940), .Y(
        \D_cache/n1399 ) );
  MX2X1 U5073 ( .A(\D_cache/cache[6][49] ), .B(n10768), .S0(n4959), .Y(
        \D_cache/n1398 ) );
  MX2X1 U5074 ( .A(\D_cache/cache[7][49] ), .B(n10768), .S0(n5003), .Y(
        \D_cache/n1397 ) );
  MX2X1 U5075 ( .A(\D_cache/cache[0][63] ), .B(n10873), .S0(n4735), .Y(
        \D_cache/n1292 ) );
  CLKMX2X2 U5076 ( .A(\D_cache/cache[1][63] ), .B(n10873), .S0(n4783), .Y(
        \D_cache/n1291 ) );
  CLKMX2X2 U5077 ( .A(\D_cache/cache[2][63] ), .B(n10873), .S0(n4805), .Y(
        \D_cache/n1290 ) );
  CLKMX2X2 U5078 ( .A(\D_cache/cache[3][63] ), .B(n10873), .S0(n4849), .Y(
        \D_cache/n1289 ) );
  CLKMX2X2 U5079 ( .A(\D_cache/cache[4][63] ), .B(n10873), .S0(n4898), .Y(
        \D_cache/n1288 ) );
  CLKMX2X2 U5080 ( .A(\D_cache/cache[5][63] ), .B(n10873), .S0(n4940), .Y(
        \D_cache/n1287 ) );
  CLKMX2X2 U5081 ( .A(\D_cache/cache[6][63] ), .B(n10873), .S0(n4959), .Y(
        \D_cache/n1286 ) );
  CLKMX2X2 U5082 ( .A(\D_cache/cache[7][63] ), .B(n10873), .S0(n5003), .Y(
        \D_cache/n1285 ) );
  MXI2X4 U5083 ( .A(n10872), .B(n10871), .S0(n5520), .Y(n10873) );
  AOI222X4 U5084 ( .A0(n5495), .A1(n11449), .B0(mem_rdata_D[99]), .B1(n233), 
        .C0(n12984), .C1(n5494), .Y(n9985) );
  MXI2X6 U5085 ( .A(n9985), .B(n9984), .S0(n5513), .Y(n9992) );
  NAND2BX2 U5086 ( .AN(n5430), .B(n11232), .Y(n9610) );
  XOR3X2 U5087 ( .A(n10613), .B(n10612), .C(n10611), .Y(n10616) );
  BUFX20 U5088 ( .A(n3915), .Y(n4073) );
  INVX4 U5089 ( .A(n11423), .Y(n10698) );
  NAND4X4 U5090 ( .A(n8691), .B(n8690), .C(n8689), .D(n8688), .Y(n11423) );
  AO22X1 U5091 ( .A0(n4731), .A1(n385), .B0(n4724), .B1(n2508), .Y(n7601) );
  OAI2BB2X1 U5092 ( .B0(\i_MIPS/n213 ), .B1(net108192), .A0N(n10855), .A1N(
        n4073), .Y(\i_MIPS/N56 ) );
  OAI2BB2X1 U5093 ( .B0(\i_MIPS/n196 ), .B1(net108192), .A0N(n10603), .A1N(
        n4072), .Y(\i_MIPS/N39 ) );
  NOR2X8 U5094 ( .A(n6423), .B(n6424), .Y(n6425) );
  CLKMX2X2 U5095 ( .A(\D_cache/cache[7][119] ), .B(n10948), .S0(n5008), .Y(
        \D_cache/n837 ) );
  CLKMX2X2 U5096 ( .A(\D_cache/cache[6][119] ), .B(n10948), .S0(n4964), .Y(
        \D_cache/n838 ) );
  CLKMX2X2 U5097 ( .A(\D_cache/cache[5][119] ), .B(n10948), .S0(n4943), .Y(
        \D_cache/n839 ) );
  CLKMX2X2 U5098 ( .A(\D_cache/cache[4][119] ), .B(n10948), .S0(n4900), .Y(
        \D_cache/n840 ) );
  CLKMX2X2 U5099 ( .A(\D_cache/cache[2][119] ), .B(n10948), .S0(n4809), .Y(
        \D_cache/n842 ) );
  CLKINVX1 U5100 ( .A(n7044), .Y(n7049) );
  MXI2X2 U5101 ( .A(n10289), .B(n10288), .S0(n5514), .Y(n10290) );
  CLKMX2X2 U5102 ( .A(\D_cache/cache[7][141] ), .B(n11035), .S0(n5007), .Y(
        \D_cache/n661 ) );
  OA22X2 U5103 ( .A0(n4757), .A1(n689), .B0(n4793), .B1(n2323), .Y(n7189) );
  INVX8 U5104 ( .A(n11429), .Y(n10755) );
  AOI222X2 U5105 ( .A0(n5505), .A1(n11381), .B0(mem_rdata_D[31]), .B1(n232), 
        .C0(n12956), .C1(n5502), .Y(n10875) );
  OAI21X4 U5106 ( .A0(n4541), .A1(net105781), .B0(n4080), .Y(n4376) );
  AOI222X2 U5107 ( .A0(n5504), .A1(n11356), .B0(mem_rdata_D[6]), .B1(n235), 
        .C0(n12981), .C1(n5501), .Y(n10080) );
  NAND3BX4 U5108 ( .AN(n8079), .B(n7805), .C(n7803), .Y(n8228) );
  OA22X1 U5109 ( .A0(n4968), .A1(n1076), .B0(n5027), .B1(n2653), .Y(n9181) );
  NAND2BX1 U5110 ( .AN(\i_MIPS/ALUOp[1] ), .B(n3704), .Y(n6479) );
  OA22X1 U5111 ( .A0(n5400), .A1(n1650), .B0(n5344), .B1(n3232), .Y(n9954) );
  XOR3X2 U5112 ( .A(n10370), .B(n10369), .C(n10368), .Y(n10377) );
  OA22X1 U5113 ( .A0(n4820), .A1(n1221), .B0(n4866), .B1(n2758), .Y(n8398) );
  OA22X2 U5114 ( .A0(n4973), .A1(n762), .B0(n5018), .B1(n2324), .Y(n8396) );
  OA22X2 U5115 ( .A0(n4748), .A1(n763), .B0(n4790), .B1(n2325), .Y(n8399) );
  AOI222X4 U5116 ( .A0(n5511), .A1(n11389), .B0(mem_rdata_D[39]), .B1(n232), 
        .C0(n12980), .C1(n5507), .Y(n10891) );
  NAND2X6 U5117 ( .A(\i_MIPS/ALUin1[4] ), .B(n6532), .Y(n6844) );
  AO22X4 U5118 ( .A0(mem_rdata_I[29]), .A1(n5541), .B0(n250), .B1(n11215), .Y(
        n6231) );
  NAND4X2 U5119 ( .A(n6230), .B(n6229), .C(n6228), .D(n6227), .Y(n11215) );
  INVX4 U5120 ( .A(n9566), .Y(n10349) );
  INVX8 U5121 ( .A(n11461), .Y(n10752) );
  AOI222X2 U5122 ( .A0(n5496), .A1(n11461), .B0(mem_rdata_D[111]), .B1(n235), 
        .C0(n12972), .C1(n5493), .Y(n10753) );
  NAND4X4 U5123 ( .A(n7185), .B(n7184), .C(n7183), .D(n7182), .Y(n11461) );
  INVX8 U5124 ( .A(n11420), .Y(n10073) );
  NAND4X4 U5125 ( .A(n7011), .B(n7010), .C(n7009), .D(n7008), .Y(n11420) );
  XNOR2X4 U5126 ( .A(n10794), .B(n10849), .Y(n3931) );
  CLKBUFX4 U5127 ( .A(n4927), .Y(n4923) );
  INVX3 U5128 ( .A(n11475), .Y(n10681) );
  NAND4X2 U5129 ( .A(n8191), .B(n8190), .C(n8189), .D(n8188), .Y(n11475) );
  XNOR2X4 U5130 ( .A(n4093), .B(n4134), .Y(n3934) );
  XOR2X4 U5131 ( .A(net128955), .B(net98722), .Y(n3936) );
  OA22X4 U5132 ( .A0(n5124), .A1(n1721), .B0(n5080), .B1(n3322), .Y(n10190) );
  OA22X1 U5133 ( .A0(n5122), .A1(n1651), .B0(n5083), .B1(n3233), .Y(n10091) );
  BUFX4 U5134 ( .A(n5125), .Y(n5122) );
  OA22X1 U5135 ( .A0(n5213), .A1(n1652), .B0(n5170), .B1(n3234), .Y(n10090) );
  AND2X8 U5136 ( .A(n8642), .B(n7308), .Y(n6506) );
  AO22X4 U5137 ( .A0(mem_rdata_I[4]), .A1(n5536), .B0(n253), .B1(n11190), .Y(
        n11086) );
  AO22X4 U5138 ( .A0(mem_rdata_I[1]), .A1(n5536), .B0(n252), .B1(n11187), .Y(
        n11074) );
  AO22X4 U5139 ( .A0(mem_rdata_I[36]), .A1(n5536), .B0(n253), .B1(n11222), .Y(
        n11087) );
  AO22X4 U5140 ( .A0(mem_rdata_I[33]), .A1(n5536), .B0(n253), .B1(n11219), .Y(
        n11075) );
  AO22X4 U5141 ( .A0(mem_rdata_I[68]), .A1(n5536), .B0(n249), .B1(n11254), .Y(
        n11085) );
  CLKMX2X2 U5142 ( .A(n7230), .B(n8348), .S0(net107798), .Y(n7896) );
  INVX8 U5143 ( .A(n11388), .Y(n10086) );
  AOI222X1 U5144 ( .A0(n5510), .A1(n11388), .B0(mem_rdata_D[38]), .B1(n236), 
        .C0(n12981), .C1(n5506), .Y(n10087) );
  NAND4X4 U5145 ( .A(n7019), .B(n7018), .C(n7017), .D(n7016), .Y(n11388) );
  BUFX16 U5146 ( .A(n5508), .Y(n5510) );
  OA22X4 U5147 ( .A0(n4997), .A1(n2085), .B0(n5025), .B1(n497), .Y(n7577) );
  INVX8 U5148 ( .A(n11377), .Y(n10307) );
  AOI222X2 U5149 ( .A0(n5504), .A1(n11377), .B0(mem_rdata_D[27]), .B1(n233), 
        .C0(n12960), .C1(n5501), .Y(n10308) );
  NAND4X2 U5150 ( .A(n8300), .B(n8299), .C(n8298), .D(n8297), .Y(n11470) );
  OA22X2 U5151 ( .A0(n10776), .A1(n4675), .B0(n10779), .B1(n4250), .Y(n8314)
         );
  INVX6 U5152 ( .A(n11438), .Y(n10779) );
  OAI221X2 U5153 ( .A0(net105045), .A1(net111624), .B0(net105046), .B1(
        net111636), .C0(net105047), .Y(n4132) );
  NAND4X4 U5154 ( .A(n8099), .B(n8098), .C(n8097), .D(n8096), .Y(n11430) );
  INVX8 U5155 ( .A(n11430), .Y(n10291) );
  AO22X4 U5156 ( .A0(n4072), .A1(n9560), .B0(net112406), .B1(
        \i_MIPS/IR_ID[31] ), .Y(\i_MIPS/N89 ) );
  OA22X2 U5157 ( .A0(n5212), .A1(n1473), .B0(n5169), .B1(n3047), .Y(n10024) );
  NAND2X4 U5158 ( .A(n10593), .B(n10591), .Y(n10389) );
  CLKAND2X12 U5159 ( .A(n10401), .B(n10404), .Y(n4389) );
  OA22X2 U5160 ( .A0(n10275), .A1(n4245), .B0(n10278), .B1(n4246), .Y(n8995)
         );
  NOR2BX4 U5161 ( .AN(\i_MIPS/IR_ID[16] ), .B(\i_MIPS/n314 ), .Y(n4522) );
  NOR4X4 U5162 ( .A(n8031), .B(n8030), .C(n8029), .D(n8028), .Y(n8032) );
  AOI222X1 U5163 ( .A0(n5495), .A1(n11466), .B0(mem_rdata_D[116]), .B1(n236), 
        .C0(n12967), .C1(n5494), .Y(n10655) );
  OA22X2 U5164 ( .A0(n4921), .A1(n764), .B0(n4949), .B1(n2326), .Y(n7191) );
  BUFX2 U5165 ( .A(n4929), .Y(n4921) );
  OA22X1 U5166 ( .A0(n4757), .A1(n1222), .B0(n4793), .B1(n2759), .Y(n7193) );
  NAND3X6 U5167 ( .A(n3770), .B(n6577), .C(n8072), .Y(n9265) );
  AND2XL U5168 ( .A(n5557), .B(n11190), .Y(n12926) );
  AND2XL U5169 ( .A(n5557), .B(n11191), .Y(n12925) );
  AND2XL U5170 ( .A(n5557), .B(n11192), .Y(n12924) );
  AOI222X2 U5171 ( .A0(n5504), .A1(n11370), .B0(mem_rdata_D[20]), .B1(n236), 
        .C0(n12967), .C1(n5501), .Y(n10661) );
  AND2XL U5172 ( .A(n5557), .B(n11193), .Y(n12923) );
  AND2XL U5173 ( .A(n5557), .B(n11194), .Y(n12922) );
  AND2XL U5174 ( .A(n5557), .B(n11195), .Y(n12921) );
  AND2XL U5175 ( .A(n5557), .B(n11196), .Y(n12920) );
  XNOR2X4 U5176 ( .A(net98061), .B(n4096), .Y(n3945) );
  XNOR2X4 U5177 ( .A(n4095), .B(net98027), .Y(n3947) );
  XNOR2X4 U5178 ( .A(n4094), .B(net98044), .Y(n3948) );
  AND2XL U5179 ( .A(n5557), .B(n11197), .Y(n12919) );
  AND2XL U5180 ( .A(n5557), .B(n11198), .Y(n12918) );
  OAI221X2 U5181 ( .A0(net104105), .A1(net111624), .B0(net104106), .B1(
        net111636), .C0(net104107), .Y(n4138) );
  AND2XL U5182 ( .A(n5557), .B(n11199), .Y(n12917) );
  NAND2BX4 U5183 ( .AN(n5429), .B(n11225), .Y(n10132) );
  NAND4X4 U5184 ( .A(n10130), .B(n10129), .C(n10128), .D(n10127), .Y(n11225)
         );
  OAI2BB1X4 U5185 ( .A0N(n10577), .A1N(n10835), .B0(n10573), .Y(n10344) );
  AOI222X1 U5186 ( .A0(n5495), .A1(n11450), .B0(mem_rdata_D[100]), .B1(n234), 
        .C0(n12983), .C1(n5494), .Y(n10967) );
  OA22X2 U5187 ( .A0(n10966), .A1(n4675), .B0(n10969), .B1(n4250), .Y(n6897)
         );
  AO21X4 U5188 ( .A0(n10322), .A1(n10321), .B0(net111640), .Y(n8525) );
  NOR4X2 U5189 ( .A(n7997), .B(n7996), .C(n7995), .D(n7994), .Y(n8008) );
  AO22XL U5190 ( .A0(net112004), .A1(n338), .B0(net112032), .B1(n1053), .Y(
        n7994) );
  NAND3BX4 U5191 ( .AN(n9482), .B(n8851), .C(n9456), .Y(n8239) );
  INVX1 U5192 ( .A(n9456), .Y(n7532) );
  NAND3X2 U5193 ( .A(n9456), .B(n9138), .C(n8854), .Y(n8855) );
  NAND2X4 U5194 ( .A(\i_MIPS/ALUin1[23] ), .B(n3841), .Y(n8852) );
  AOI222X1 U5195 ( .A0(n5511), .A1(n11395), .B0(mem_rdata_D[45]), .B1(n233), 
        .C0(n12974), .C1(n5507), .Y(n10740) );
  CLKMX2X2 U5196 ( .A(\I_cache/cache[2][99] ), .B(n11169), .S0(n5189), .Y(
        n11993) );
  CLKMX2X2 U5197 ( .A(\I_cache/cache[0][99] ), .B(n11169), .S0(n5098), .Y(
        n11995) );
  CLKMX2X2 U5198 ( .A(\I_cache/cache[5][99] ), .B(n11169), .S0(n5233), .Y(
        n11990) );
  CLKMX2X2 U5199 ( .A(\I_cache/cache[4][99] ), .B(n11169), .S0(n5276), .Y(
        n11991) );
  CLKMX2X2 U5200 ( .A(\I_cache/cache[3][99] ), .B(n11169), .S0(n5143), .Y(
        n11992) );
  CLKMX2X2 U5201 ( .A(\I_cache/cache[7][99] ), .B(n11169), .S0(n5321), .Y(
        n11988) );
  CLKMX2X2 U5202 ( .A(\I_cache/cache[6][99] ), .B(n11169), .S0(n5358), .Y(
        n11989) );
  AO22X2 U5203 ( .A0(mem_rdata_I[3]), .A1(n5535), .B0(n253), .B1(n11189), .Y(
        n11169) );
  XNOR2X4 U5204 ( .A(n10636), .B(n14), .Y(n3955) );
  XNOR2X4 U5205 ( .A(n8725), .B(n10694), .Y(n3956) );
  XNOR2X4 U5206 ( .A(n10507), .B(n8827), .Y(n3958) );
  CLKAND2X12 U5207 ( .A(n4657), .B(n11234), .Y(mem_wdata_I[48]) );
  AND2XL U5208 ( .A(n5557), .B(n11204), .Y(n12916) );
  AND2XL U5209 ( .A(n4657), .B(n11235), .Y(n12889) );
  AND2XL U5210 ( .A(n5557), .B(n11205), .Y(n12915) );
  CLKAND2X12 U5211 ( .A(mem_write_I), .B(n11237), .Y(mem_wdata_I[51]) );
  AND2XL U5212 ( .A(n4657), .B(n11238), .Y(n12888) );
  AND2XL U5213 ( .A(n5557), .B(n11206), .Y(n12914) );
  AND2XL U5214 ( .A(n5557), .B(n11207), .Y(n12913) );
  AND2XL U5215 ( .A(n5557), .B(n11208), .Y(n12912) );
  AND2XL U5216 ( .A(n5557), .B(n11209), .Y(n12911) );
  AND2XL U5217 ( .A(n5557), .B(n11210), .Y(n12910) );
  AND2XL U5218 ( .A(n5557), .B(n11211), .Y(n12909) );
  AND2XL U5219 ( .A(n5557), .B(n11212), .Y(n12908) );
  AND2XL U5220 ( .A(n5557), .B(n11213), .Y(n12907) );
  AND2XL U5221 ( .A(n5557), .B(n11214), .Y(n12906) );
  AND2XL U5222 ( .A(n5557), .B(n11216), .Y(n12904) );
  AND2XL U5223 ( .A(n5557), .B(n11217), .Y(n12903) );
  AND2XL U5224 ( .A(n5557), .B(n11218), .Y(n12902) );
  AOI222X2 U5225 ( .A0(n3838), .A1(n9332), .B0(n7232), .B1(net100585), .C0(
        net103548), .C1(n4418), .Y(n7233) );
  AND2XL U5226 ( .A(n5557), .B(n11219), .Y(n12901) );
  AND2XL U5227 ( .A(n5557), .B(n11221), .Y(n12900) );
  OA22X2 U5228 ( .A0(n4908), .A1(n693), .B0(n4947), .B1(n2262), .Y(n9081) );
  AND2XL U5229 ( .A(n5557), .B(n11222), .Y(n12899) );
  AND2XL U5230 ( .A(n5557), .B(n11223), .Y(n12898) );
  NAND2X1 U5231 ( .A(n4651), .B(n6120), .Y(n11130) );
  AND2XL U5232 ( .A(n5557), .B(n11224), .Y(n12897) );
  AND2XL U5233 ( .A(n5557), .B(n11225), .Y(n12896) );
  AND2XL U5234 ( .A(n5557), .B(n11226), .Y(n12895) );
  AND2XL U5235 ( .A(n4657), .B(n11241), .Y(n12886) );
  AND2XL U5236 ( .A(n5556), .B(n11243), .Y(n12884) );
  AND2XL U5237 ( .A(n4656), .B(n11239), .Y(n12887) );
  AND2XL U5238 ( .A(n5557), .B(n11228), .Y(n12894) );
  AND2XL U5239 ( .A(n4657), .B(n11244), .Y(n12883) );
  AND2XL U5240 ( .A(n4656), .B(n11246), .Y(n12881) );
  AND2XL U5241 ( .A(n4656), .B(n11242), .Y(n12885) );
  AND2XL U5242 ( .A(n5557), .B(n11229), .Y(n12893) );
  AND2XL U5243 ( .A(n4657), .B(n11247), .Y(n12880) );
  AND2XL U5244 ( .A(n4657), .B(n11249), .Y(n12878) );
  AND2XL U5245 ( .A(n4656), .B(n11245), .Y(n12882) );
  AND2XL U5246 ( .A(n5557), .B(n11230), .Y(n12892) );
  AND2XL U5247 ( .A(n4657), .B(n11250), .Y(n12877) );
  INVX8 U5248 ( .A(n11360), .Y(n10263) );
  AND2XL U5249 ( .A(n5556), .B(n11255), .Y(n12873) );
  AND2XL U5250 ( .A(n4656), .B(n11248), .Y(n12879) );
  AND2XL U5251 ( .A(n5557), .B(n11231), .Y(n12891) );
  AND2XL U5252 ( .A(n4657), .B(n11253), .Y(n12875) );
  AND2XL U5253 ( .A(mem_write_I), .B(n11258), .Y(n12870) );
  AND2XL U5254 ( .A(n4656), .B(n11251), .Y(n12876) );
  AND2XL U5255 ( .A(n4657), .B(n11256), .Y(n12872) );
  AND2XL U5256 ( .A(n5556), .B(n11261), .Y(n12867) );
  AND2XL U5257 ( .A(n4656), .B(n11254), .Y(n12874) );
  NAND4X4 U5258 ( .A(n9191), .B(n9190), .C(n9189), .D(n9188), .Y(n11371) );
  AOI222X2 U5259 ( .A0(n5504), .A1(n11371), .B0(mem_rdata_D[21]), .B1(n236), 
        .C0(n12966), .C1(n5501), .Y(n10674) );
  AND2XL U5260 ( .A(n4657), .B(n11259), .Y(n12869) );
  AND2XL U5261 ( .A(mem_write_I), .B(n11264), .Y(n12864) );
  AND2XL U5262 ( .A(n4656), .B(n11257), .Y(n12871) );
  AND2XL U5263 ( .A(n4657), .B(n11262), .Y(n12866) );
  AND2XL U5264 ( .A(n5556), .B(n11267), .Y(n12861) );
  AND2XL U5265 ( .A(n4656), .B(n11260), .Y(n12868) );
  AND2XL U5266 ( .A(n4657), .B(n11265), .Y(n12863) );
  AND2XL U5267 ( .A(mem_write_I), .B(n11270), .Y(n12858) );
  AND2XL U5268 ( .A(n4656), .B(n11263), .Y(n12865) );
  AOI2BB1X4 U5269 ( .A0N(n10391), .A1N(n10592), .B0(n10390), .Y(n10392) );
  AND2XL U5270 ( .A(n4657), .B(n11268), .Y(n12860) );
  AND2XL U5271 ( .A(mem_write_I), .B(n11273), .Y(n12855) );
  AND2XL U5272 ( .A(n4656), .B(n11266), .Y(n12862) );
  AND2XL U5273 ( .A(n4657), .B(n11271), .Y(n12857) );
  AND2XL U5274 ( .A(n5556), .B(n11276), .Y(n12852) );
  AND2XL U5275 ( .A(n4656), .B(n11269), .Y(n12859) );
  AND2XL U5276 ( .A(n4657), .B(n11274), .Y(n12854) );
  AND2XL U5277 ( .A(n5556), .B(n11279), .Y(n12849) );
  AND2XL U5278 ( .A(n4656), .B(n11272), .Y(n12856) );
  AND2XL U5279 ( .A(n4657), .B(n11277), .Y(n12851) );
  AND2XL U5280 ( .A(mem_write_I), .B(n11282), .Y(n12846) );
  AND2XL U5281 ( .A(n4656), .B(n11275), .Y(n12853) );
  AND2XL U5282 ( .A(n4657), .B(n11280), .Y(n12848) );
  AND2XL U5283 ( .A(n5556), .B(n11285), .Y(n12843) );
  AND2XL U5284 ( .A(n4656), .B(n11278), .Y(n12850) );
  AOI222X1 U5285 ( .A0(n5503), .A1(n11354), .B0(mem_rdata_D[4]), .B1(n236), 
        .C0(n12983), .C1(n5502), .Y(n10973) );
  OA22X2 U5286 ( .A0(n10972), .A1(n4245), .B0(n10975), .B1(n4246), .Y(n6896)
         );
  AND2XL U5287 ( .A(n4657), .B(n11283), .Y(n12845) );
  AND2XL U5288 ( .A(mem_write_I), .B(n11288), .Y(n12841) );
  CLKINVX8 U5289 ( .A(n9249), .Y(n9159) );
  AND2XL U5290 ( .A(n4656), .B(n11281), .Y(n12847) );
  AND2XL U5291 ( .A(n4657), .B(n11286), .Y(n12842) );
  AND2XL U5292 ( .A(mem_write_I), .B(n11291), .Y(n12838) );
  AND2XL U5293 ( .A(n4656), .B(n11284), .Y(n12844) );
  AND2XL U5294 ( .A(n4657), .B(n11289), .Y(n12840) );
  AND2XL U5295 ( .A(n5556), .B(n11297), .Y(n12835) );
  AND2XL U5296 ( .A(n4656), .B(n11290), .Y(n12839) );
  AND2XL U5297 ( .A(n4657), .B(n11292), .Y(n12837) );
  AND2XL U5298 ( .A(mem_write_I), .B(n11300), .Y(n12832) );
  AND2XL U5299 ( .A(n4656), .B(n11299), .Y(n12833) );
  AND2XL U5300 ( .A(n4657), .B(n11295), .Y(n12836) );
  AND2XL U5301 ( .A(mem_write_I), .B(n11303), .Y(n12829) );
  AND2XL U5302 ( .A(n4656), .B(n11302), .Y(n12830) );
  AND2XL U5303 ( .A(n4657), .B(n11298), .Y(n12834) );
  AND2XL U5304 ( .A(mem_write_I), .B(n11306), .Y(n12826) );
  AND2XL U5305 ( .A(n4656), .B(n11305), .Y(n12827) );
  AND2XL U5306 ( .A(n4657), .B(n11301), .Y(n12831) );
  AND2XL U5307 ( .A(n5556), .B(n11309), .Y(n12823) );
  AND2XL U5308 ( .A(n4657), .B(n11304), .Y(n12828) );
  AND2XL U5309 ( .A(n4656), .B(n11311), .Y(n12821) );
  AND2XL U5310 ( .A(n4657), .B(n11307), .Y(n12825) );
  AND2XL U5311 ( .A(n4657), .B(n11310), .Y(n12822) );
  OA22X4 U5312 ( .A0(\i_MIPS/Register/register[1][13] ), .A1(net112258), .B0(
        \i_MIPS/Register/register[9][13] ), .B1(n151), .Y(n7721) );
  OA22X2 U5313 ( .A0(n5120), .A1(n1474), .B0(n5082), .B1(n3048), .Y(n9957) );
  AND3X2 U5314 ( .A(n8729), .B(net137952), .C(n8747), .Y(n8744) );
  CLKMX2X2 U5315 ( .A(\I_cache/cache[6][79] ), .B(n9658), .S0(n5359), .Y(
        n12149) );
  CLKMX2X2 U5316 ( .A(\I_cache/cache[7][79] ), .B(n9658), .S0(n5318), .Y(
        n12148) );
  CLKMX2X2 U5317 ( .A(\I_cache/cache[2][79] ), .B(n9658), .S0(n5186), .Y(
        n12153) );
  CLKMX2X2 U5318 ( .A(\I_cache/cache[3][79] ), .B(n9658), .S0(n5140), .Y(
        n12152) );
  CLKMX2X2 U5319 ( .A(\I_cache/cache[4][79] ), .B(n9658), .S0(n5272), .Y(
        n12151) );
  CLKMX2X2 U5320 ( .A(\I_cache/cache[5][79] ), .B(n9658), .S0(n5229), .Y(
        n12150) );
  AO22X2 U5321 ( .A0(mem_rdata_I[47]), .A1(n5540), .B0(n250), .B1(n11233), .Y(
        n9658) );
  INVX4 U5322 ( .A(n8173), .Y(n6595) );
  AO22X4 U5323 ( .A0(n4090), .A1(net137952), .B0(net112296), .B1(net102429), 
        .Y(n4088) );
  XOR2X4 U5324 ( .A(n10319), .B(n3890), .Y(n9551) );
  NOR4X1 U5325 ( .A(net103907), .B(n7491), .C(n7490), .D(n8951), .Y(n7546) );
  OA21X4 U5326 ( .A0(n8951), .A1(n8237), .B0(n9043), .Y(n7478) );
  NOR2BX4 U5327 ( .AN(net108200), .B(\i_MIPS/Control_ID/n12 ), .Y(n4452) );
  NAND4X2 U5328 ( .A(\i_MIPS/IR_ID[29] ), .B(\i_MIPS/IR_ID[31] ), .C(n4544), 
        .D(n9570), .Y(n9971) );
  AND2X1 U5329 ( .A(n10467), .B(n10466), .Y(n4398) );
  AO21X2 U5330 ( .A0(n10489), .A1(n10488), .B0(net111902), .Y(n10466) );
  AO22X4 U5331 ( .A0(n241), .A1(net111966), .B0(net111962), .B1(n7738), .Y(
        net103504) );
  AOI32X2 U5332 ( .A0(n10852), .A1(n10851), .A2(n10850), .B0(net112400), .B1(
        n10849), .Y(n10854) );
  NAND2X1 U5333 ( .A(n10579), .B(net112404), .Y(n10850) );
  NAND2X2 U5334 ( .A(n6970), .B(n4381), .Y(n7875) );
  NAND2X6 U5335 ( .A(\i_MIPS/ALUin1[5] ), .B(n6535), .Y(n4381) );
  OAI2BB1X4 U5336 ( .A0N(n7305), .A1N(n7492), .B0(n7496), .Y(n7225) );
  INVX3 U5337 ( .A(n7301), .Y(n7228) );
  NAND3BX4 U5338 ( .AN(n9482), .B(n3825), .C(n325), .Y(n8853) );
  AOI222X1 U5339 ( .A0(n5504), .A1(n11376), .B0(mem_rdata_D[26]), .B1(n232), 
        .C0(n12961), .C1(n5501), .Y(n10276) );
  NAND4X2 U5340 ( .A(n8990), .B(n8989), .C(n8988), .D(n8987), .Y(n11376) );
  AND4X4 U5341 ( .A(n6610), .B(n6609), .C(n6608), .D(n6607), .Y(net133317) );
  NAND4X4 U5342 ( .A(n6887), .B(n6886), .C(n6885), .D(n6884), .Y(n11418) );
  INVX8 U5343 ( .A(n11418), .Y(n10969) );
  AOI222X1 U5344 ( .A0(n5500), .A1(n11418), .B0(mem_rdata_D[68]), .B1(n232), 
        .C0(n12983), .C1(n4385), .Y(n10970) );
  NOR4X2 U5345 ( .A(n7735), .B(n7734), .C(n7733), .D(n7732), .Y(n7736) );
  AOI222X4 U5346 ( .A0(n5511), .A1(n11390), .B0(mem_rdata_D[40]), .B1(n233), 
        .C0(n12979), .C1(n5507), .Y(n10903) );
  AO22X4 U5347 ( .A0(mem_rdata_I[15]), .A1(n5540), .B0(n250), .B1(n11201), .Y(
        n9648) );
  NAND4X6 U5348 ( .A(n9647), .B(n9646), .C(n9645), .D(n9644), .Y(n11201) );
  NAND2X2 U5349 ( .A(n11121), .B(n3865), .Y(n10542) );
  INVX4 U5350 ( .A(n7485), .Y(n6480) );
  NAND2X4 U5351 ( .A(net103910), .B(net133411), .Y(n7485) );
  CLKMX2X2 U5352 ( .A(\D_cache/cache[7][30] ), .B(n10141), .S0(n5002), .Y(
        \D_cache/n1549 ) );
  CLKMX2X2 U5353 ( .A(\D_cache/cache[6][30] ), .B(n10141), .S0(n4960), .Y(
        \D_cache/n1550 ) );
  CLKMX2X2 U5354 ( .A(\D_cache/cache[5][30] ), .B(n10141), .S0(n4943), .Y(
        \D_cache/n1551 ) );
  CLKMX2X2 U5355 ( .A(\D_cache/cache[4][30] ), .B(n10141), .S0(n4894), .Y(
        \D_cache/n1552 ) );
  CLKMX2X2 U5356 ( .A(\D_cache/cache[3][30] ), .B(n10141), .S0(n4847), .Y(
        \D_cache/n1553 ) );
  CLKMX2X2 U5357 ( .A(\D_cache/cache[2][30] ), .B(n10141), .S0(n4803), .Y(
        \D_cache/n1554 ) );
  CLKMX2X2 U5358 ( .A(\D_cache/cache[1][30] ), .B(n10141), .S0(n4780), .Y(
        \D_cache/n1555 ) );
  MX2X1 U5359 ( .A(\D_cache/cache[0][30] ), .B(n10141), .S0(n4734), .Y(
        \D_cache/n1556 ) );
  NAND2X6 U5360 ( .A(\i_MIPS/ALUin1[27] ), .B(n6588), .Y(n9347) );
  BUFX16 U5361 ( .A(n4884), .Y(n4880) );
  AOI222X4 U5362 ( .A0(n5510), .A1(n11392), .B0(mem_rdata_D[42]), .B1(n236), 
        .C0(n12977), .C1(n5506), .Y(n10267) );
  NAND4X4 U5363 ( .A(n7359), .B(n7358), .C(n7357), .D(n7356), .Y(n11392) );
  INVX8 U5364 ( .A(n11392), .Y(n10266) );
  MX2X6 U5365 ( .A(n8866), .B(n7899), .S0(net107796), .Y(n9332) );
  CLKMX2X4 U5366 ( .A(n7899), .B(n7898), .S0(net107796), .Y(n7900) );
  OAI221X4 U5367 ( .A0(net112368), .A1(\i_MIPS/n367 ), .B0(net112348), .B1(
        \i_MIPS/n366 ), .C0(n6686), .Y(n7899) );
  MX2X1 U5368 ( .A(\D_cache/cache[5][20] ), .B(n10656), .S0(n4936), .Y(
        \D_cache/n1631 ) );
  CLKMX2X2 U5369 ( .A(\D_cache/cache[6][20] ), .B(n10656), .S0(n4957), .Y(
        \D_cache/n1630 ) );
  CLKMX2X2 U5370 ( .A(\D_cache/cache[7][20] ), .B(n10656), .S0(n5001), .Y(
        \D_cache/n1629 ) );
  NOR4X2 U5371 ( .A(n7331), .B(n7330), .C(n7329), .D(n7328), .Y(n7342) );
  NAND2X1 U5372 ( .A(n8730), .B(n8738), .Y(n8747) );
  AO21X4 U5373 ( .A0(n10152), .A1(n10151), .B0(net111640), .Y(n8628) );
  BUFX20 U5374 ( .A(n4384), .Y(n5501) );
  NAND4X4 U5375 ( .A(n8103), .B(n8102), .C(n8101), .D(n8100), .Y(n11366) );
  OA22X2 U5376 ( .A0(n4975), .A1(n694), .B0(n5020), .B1(n2263), .Y(n8100) );
  BUFX12 U5377 ( .A(net100424), .Y(net111636) );
  OAI211X2 U5378 ( .A0(n7973), .A1(net103076), .B0(n7971), .C0(n7972), .Y(
        n7988) );
  OA21X4 U5379 ( .A0(n7408), .A1(n4070), .B0(n7406), .Y(n4154) );
  OAI31X4 U5380 ( .A0(n6509), .A1(n6508), .A2(n6507), .B0(n6506), .Y(n4070) );
  INVX2 U5381 ( .A(n10229), .Y(n10230) );
  NAND3X4 U5382 ( .A(n3781), .B(ICACHE_addr[5]), .C(n10174), .Y(n10229) );
  AOI222X2 U5383 ( .A0(n5496), .A1(n11457), .B0(mem_rdata_D[107]), .B1(n235), 
        .C0(n12976), .C1(n5493), .Y(n10708) );
  NAND2X4 U5384 ( .A(n4423), .B(n9330), .Y(n8449) );
  NAND2BX2 U5385 ( .AN(n8449), .B(n11181), .Y(n8172) );
  AOI222X4 U5386 ( .A0(n5505), .A1(n11355), .B0(mem_rdata_D[5]), .B1(n235), 
        .C0(n12982), .C1(n5502), .Y(n10985) );
  INVX3 U5387 ( .A(n10403), .Y(n10602) );
  NAND4X4 U5388 ( .A(n6140), .B(n6139), .C(n6138), .D(n6137), .Y(n11282) );
  OA22X2 U5389 ( .A0(n4980), .A1(n695), .B0(n5025), .B1(n2264), .Y(n7429) );
  OAI2BB1X4 U5390 ( .A0N(n10563), .A1N(n10562), .B0(net112782), .Y(n9218) );
  OA22X4 U5391 ( .A0(n4910), .A1(n2145), .B0(n4949), .B1(n565), .Y(n8992) );
  INVX8 U5392 ( .A(n11383), .Y(n10914) );
  NAND4X6 U5393 ( .A(n8024), .B(n8023), .C(n8022), .D(n8021), .Y(n11383) );
  CLKMX2X2 U5394 ( .A(\D_cache/cache[0][28] ), .B(n10477), .S0(n4732), .Y(
        \D_cache/n1572 ) );
  CLKMX2X2 U5395 ( .A(\D_cache/cache[1][28] ), .B(n10477), .S0(n4778), .Y(
        \D_cache/n1571 ) );
  CLKMX2X2 U5396 ( .A(\D_cache/cache[2][28] ), .B(n10477), .S0(n4801), .Y(
        \D_cache/n1570 ) );
  CLKMX2X2 U5397 ( .A(\D_cache/cache[3][28] ), .B(n10477), .S0(n4846), .Y(
        \D_cache/n1569 ) );
  CLKMX2X2 U5398 ( .A(\D_cache/cache[4][28] ), .B(n10477), .S0(n4892), .Y(
        \D_cache/n1568 ) );
  CLKMX2X2 U5399 ( .A(\D_cache/cache[5][28] ), .B(n10477), .S0(n4936), .Y(
        \D_cache/n1567 ) );
  CLKMX2X2 U5400 ( .A(\D_cache/cache[6][28] ), .B(n10477), .S0(n4956), .Y(
        \D_cache/n1566 ) );
  CLKMX2X2 U5401 ( .A(\D_cache/cache[7][28] ), .B(n10477), .S0(n5000), .Y(
        \D_cache/n1565 ) );
  AO21X4 U5402 ( .A0(n9488), .A1(n9487), .B0(n9486), .Y(n9493) );
  INVX20 U5403 ( .A(n1970), .Y(mem_addr_I[7]) );
  INVX20 U5404 ( .A(n1971), .Y(mem_addr_I[9]) );
  AOI221XL U5405 ( .A0(n4507), .A1(\D_cache/cache[0][140] ), .B0(n4508), .B1(
        \D_cache/cache[1][140] ), .C0(n3403), .Y(n4064) );
  INVX20 U5406 ( .A(n1972), .Y(mem_addr_I[10]) );
  NAND2X2 U5407 ( .A(n6592), .B(\i_MIPS/n344 ), .Y(n9348) );
  OAI211X1 U5408 ( .A0(n9342), .A1(n9341), .B0(n9340), .C0(n4658), .Y(n9343)
         );
  CLKMX2X4 U5409 ( .A(net100573), .B(net112438), .S0(n9338), .Y(n9340) );
  INVX20 U5410 ( .A(n1973), .Y(mem_addr_I[12]) );
  AOI222X4 U5411 ( .A0(n5495), .A1(n11472), .B0(mem_rdata_D[122]), .B1(n234), 
        .C0(n12961), .C1(n5494), .Y(n10270) );
  INVX20 U5412 ( .A(n1974), .Y(mem_addr_I[13]) );
  CLKMX2X2 U5413 ( .A(\D_cache/cache[0][19] ), .B(n10993), .S0(n4736), .Y(
        \D_cache/n1644 ) );
  CLKMX2X2 U5414 ( .A(\D_cache/cache[1][19] ), .B(n10993), .S0(n4786), .Y(
        \D_cache/n1643 ) );
  CLKMX2X2 U5415 ( .A(\D_cache/cache[2][19] ), .B(n10993), .S0(n4809), .Y(
        \D_cache/n1642 ) );
  CLKMX2X2 U5416 ( .A(\D_cache/cache[3][19] ), .B(n10993), .S0(n4855), .Y(
        \D_cache/n1641 ) );
  CLKMX2X2 U5417 ( .A(\D_cache/cache[4][19] ), .B(n10993), .S0(n4901), .Y(
        \D_cache/n1640 ) );
  CLKMX2X2 U5418 ( .A(\D_cache/cache[5][19] ), .B(n10993), .S0(n4944), .Y(
        \D_cache/n1639 ) );
  CLKMX2X2 U5419 ( .A(\D_cache/cache[6][19] ), .B(n10993), .S0(n4965), .Y(
        \D_cache/n1638 ) );
  CLKMX2X2 U5420 ( .A(\D_cache/cache[7][19] ), .B(n10993), .S0(n5009), .Y(
        \D_cache/n1637 ) );
  MXI2X1 U5421 ( .A(\i_MIPS/n288 ), .B(\i_MIPS/n289 ), .S0(n219), .Y(
        \i_MIPS/n416 ) );
  CLKMX2X2 U5422 ( .A(\D_cache/cache[7][23] ), .B(n10942), .S0(n5008), .Y(
        \D_cache/n1605 ) );
  CLKMX2X2 U5423 ( .A(\D_cache/cache[6][23] ), .B(n10942), .S0(n4964), .Y(
        \D_cache/n1606 ) );
  CLKMX2X2 U5424 ( .A(\D_cache/cache[5][23] ), .B(n10942), .S0(n4943), .Y(
        \D_cache/n1607 ) );
  CLKMX2X2 U5425 ( .A(\D_cache/cache[4][23] ), .B(n10942), .S0(n4900), .Y(
        \D_cache/n1608 ) );
  CLKMX2X2 U5426 ( .A(\D_cache/cache[3][23] ), .B(n10942), .S0(n4854), .Y(
        \D_cache/n1609 ) );
  CLKMX2X2 U5427 ( .A(\D_cache/cache[2][23] ), .B(n10942), .S0(n4809), .Y(
        \D_cache/n1610 ) );
  CLKMX2X2 U5428 ( .A(\D_cache/cache[1][23] ), .B(n10942), .S0(n4779), .Y(
        \D_cache/n1611 ) );
  CLKMX2X2 U5429 ( .A(\D_cache/cache[7][4] ), .B(n10968), .S0(n5009), .Y(
        \D_cache/n1757 ) );
  CLKMX2X2 U5430 ( .A(\D_cache/cache[6][4] ), .B(n10968), .S0(n4965), .Y(
        \D_cache/n1758 ) );
  CLKMX2X2 U5431 ( .A(\D_cache/cache[5][4] ), .B(n10968), .S0(n4944), .Y(
        \D_cache/n1759 ) );
  CLKMX2X2 U5432 ( .A(\D_cache/cache[4][4] ), .B(n10968), .S0(n4901), .Y(
        \D_cache/n1760 ) );
  CLKMX2X2 U5433 ( .A(\D_cache/cache[3][4] ), .B(n10968), .S0(n4855), .Y(
        \D_cache/n1761 ) );
  CLKMX2X2 U5434 ( .A(\D_cache/cache[2][4] ), .B(n10968), .S0(n4808), .Y(
        \D_cache/n1762 ) );
  CLKMX2X2 U5435 ( .A(\D_cache/cache[1][4] ), .B(n10968), .S0(n4786), .Y(
        \D_cache/n1763 ) );
  MX2X1 U5436 ( .A(\D_cache/cache[0][4] ), .B(n10968), .S0(n4732), .Y(
        \D_cache/n1764 ) );
  CLKMX2X2 U5437 ( .A(\D_cache/cache[7][0] ), .B(n182), .S0(n5008), .Y(
        \D_cache/n1796 ) );
  CLKMX2X2 U5438 ( .A(\D_cache/cache[6][0] ), .B(n182), .S0(n4964), .Y(
        \D_cache/n1789 ) );
  CLKMX2X2 U5439 ( .A(\D_cache/cache[5][0] ), .B(n182), .S0(n4943), .Y(
        \D_cache/n1790 ) );
  CLKMX2X2 U5440 ( .A(\D_cache/cache[4][0] ), .B(n182), .S0(n4900), .Y(
        \D_cache/n1791 ) );
  CLKMX2X2 U5441 ( .A(\D_cache/cache[2][0] ), .B(n182), .S0(n4809), .Y(
        \D_cache/n1793 ) );
  CLKMX2X2 U5442 ( .A(\D_cache/cache[1][0] ), .B(n182), .S0(n4785), .Y(
        \D_cache/n1794 ) );
  CLKMX2X2 U5443 ( .A(\D_cache/cache[1][8] ), .B(n169), .S0(n4781), .Y(
        \D_cache/n1731 ) );
  CLKMX2X2 U5444 ( .A(\D_cache/cache[2][8] ), .B(n169), .S0(n4804), .Y(
        \D_cache/n1730 ) );
  CLKMX2X2 U5445 ( .A(\D_cache/cache[3][8] ), .B(n169), .S0(n4854), .Y(
        \D_cache/n1729 ) );
  CLKMX2X2 U5446 ( .A(\D_cache/cache[4][8] ), .B(n169), .S0(n4892), .Y(
        \D_cache/n1728 ) );
  CLKMX2X2 U5447 ( .A(\D_cache/cache[5][8] ), .B(n169), .S0(n4938), .Y(
        \D_cache/n1727 ) );
  CLKMX2X2 U5448 ( .A(\D_cache/cache[6][8] ), .B(n169), .S0(n4957), .Y(
        \D_cache/n1726 ) );
  CLKMX2X2 U5449 ( .A(\D_cache/cache[7][8] ), .B(n169), .S0(n5000), .Y(
        \D_cache/n1725 ) );
  OAI2BB1X4 U5450 ( .A0N(n7221), .A1N(n7220), .B0(n8642), .Y(n7306) );
  MXI2X1 U5451 ( .A(\i_MIPS/n272 ), .B(\i_MIPS/n273 ), .S0(n219), .Y(
        \i_MIPS/n400 ) );
  NAND3BX2 U5452 ( .AN(n8760), .B(n8759), .C(net112294), .Y(n8761) );
  AO22X4 U5453 ( .A0(mem_rdata_I[122]), .A1(n5541), .B0(n250), .B1(n11308), 
        .Y(n9561) );
  AOI222X1 U5454 ( .A0(n5504), .A1(n11369), .B0(mem_rdata_D[19]), .B1(n234), 
        .C0(n5502), .C1(n12968), .Y(n11000) );
  AO22X4 U5455 ( .A0(net111966), .A1(net97834), .B0(net111962), .B1(n7930), 
        .Y(net103177) );
  AO22X4 U5456 ( .A0(net97736), .A1(net111966), .B0(net111962), .B1(n7572), 
        .Y(net103806) );
  AO22X2 U5457 ( .A0(net111966), .A1(n10320), .B0(net111962), .B1(n8485), .Y(
        n8486) );
  OAI32X2 U5458 ( .A0(n7534), .A1(n7535), .A2(n7533), .B0(n7532), .B1(n7531), 
        .Y(n7543) );
  CLKMX2X2 U5459 ( .A(\D_cache/cache[7][58] ), .B(n10274), .S0(n5002), .Y(
        \D_cache/n1325 ) );
  CLKMX2X2 U5460 ( .A(\D_cache/cache[6][58] ), .B(n10274), .S0(n4958), .Y(
        \D_cache/n1326 ) );
  CLKMX2X2 U5461 ( .A(\D_cache/cache[5][58] ), .B(n10274), .S0(n4938), .Y(
        \D_cache/n1327 ) );
  CLKMX2X2 U5462 ( .A(\D_cache/cache[4][58] ), .B(n10274), .S0(n4895), .Y(
        \D_cache/n1328 ) );
  CLKMX2X2 U5463 ( .A(\D_cache/cache[3][58] ), .B(n10274), .S0(n4848), .Y(
        \D_cache/n1329 ) );
  CLKMX2X2 U5464 ( .A(\D_cache/cache[2][58] ), .B(n10274), .S0(n4804), .Y(
        \D_cache/n1330 ) );
  CLKMX2X2 U5465 ( .A(\D_cache/cache[1][58] ), .B(n10274), .S0(n4781), .Y(
        \D_cache/n1331 ) );
  MX2X1 U5466 ( .A(\D_cache/cache[0][58] ), .B(n10274), .S0(n4735), .Y(
        \D_cache/n1332 ) );
  CLKMX2X2 U5467 ( .A(\D_cache/cache[7][48] ), .B(n10293), .S0(n5002), .Y(
        \D_cache/n1405 ) );
  CLKMX2X2 U5468 ( .A(\D_cache/cache[6][48] ), .B(n10293), .S0(n4958), .Y(
        \D_cache/n1406 ) );
  CLKMX2X2 U5469 ( .A(\D_cache/cache[5][48] ), .B(n10293), .S0(n4940), .Y(
        \D_cache/n1407 ) );
  CLKMX2X2 U5470 ( .A(\D_cache/cache[4][48] ), .B(n10293), .S0(n4895), .Y(
        \D_cache/n1408 ) );
  CLKMX2X2 U5471 ( .A(\D_cache/cache[3][48] ), .B(n10293), .S0(n4848), .Y(
        \D_cache/n1409 ) );
  CLKMX2X2 U5472 ( .A(\D_cache/cache[2][48] ), .B(n10293), .S0(n4804), .Y(
        \D_cache/n1410 ) );
  CLKMX2X2 U5473 ( .A(\D_cache/cache[1][48] ), .B(n10293), .S0(n4783), .Y(
        \D_cache/n1411 ) );
  INVXL U5474 ( .A(n10331), .Y(n4071) );
  AOI222X1 U5475 ( .A0(n5510), .A1(n11398), .B0(mem_rdata_D[48]), .B1(n235), 
        .C0(n12971), .C1(n5506), .Y(n10298) );
  MX2XL U5476 ( .A(n3600), .B(net98722), .S0(n214), .Y(\i_MIPS/n405 ) );
  OA22X2 U5477 ( .A0(n5303), .A1(n1475), .B0(n5257), .B1(n3049), .Y(n10041) );
  OA22X2 U5478 ( .A0(n5303), .A1(n765), .B0(n5257), .B1(n2327), .Y(n10023) );
  OA22X2 U5479 ( .A0(n5303), .A1(n1476), .B0(n5257), .B1(n3050), .Y(n10051) );
  OA22X2 U5480 ( .A0(n5303), .A1(n1451), .B0(n5257), .B1(n3024), .Y(n10046) );
  CLKBUFX3 U5481 ( .A(n5261), .Y(n5257) );
  CLKMX2X2 U5482 ( .A(\D_cache/cache[7][126] ), .B(n166), .S0(n5000), .Y(
        \D_cache/n781 ) );
  CLKMX2X2 U5483 ( .A(\D_cache/cache[6][126] ), .B(n166), .S0(n4959), .Y(
        \D_cache/n782 ) );
  CLKMX2X2 U5484 ( .A(\D_cache/cache[5][126] ), .B(n166), .S0(n4936), .Y(
        \D_cache/n783 ) );
  CLKMX2X2 U5485 ( .A(\D_cache/cache[4][126] ), .B(n166), .S0(n4894), .Y(
        \D_cache/n784 ) );
  CLKMX2X2 U5486 ( .A(\D_cache/cache[3][126] ), .B(n166), .S0(n4846), .Y(
        \D_cache/n785 ) );
  CLKMX2X2 U5487 ( .A(\D_cache/cache[2][126] ), .B(n166), .S0(n4803), .Y(
        \D_cache/n786 ) );
  CLKMX2X2 U5488 ( .A(\D_cache/cache[1][126] ), .B(n166), .S0(n4780), .Y(
        \D_cache/n787 ) );
  CLKMX2X2 U5489 ( .A(\D_cache/cache[7][118] ), .B(n10217), .S0(n5003), .Y(
        \D_cache/n845 ) );
  CLKMX2X2 U5490 ( .A(\D_cache/cache[6][118] ), .B(n10217), .S0(n4964), .Y(
        \D_cache/n846 ) );
  CLKMX2X2 U5491 ( .A(\D_cache/cache[5][118] ), .B(n10217), .S0(n4936), .Y(
        \D_cache/n847 ) );
  CLKMX2X2 U5492 ( .A(\D_cache/cache[4][118] ), .B(n10217), .S0(n4894), .Y(
        \D_cache/n848 ) );
  CLKMX2X2 U5493 ( .A(\D_cache/cache[3][118] ), .B(n10217), .S0(n4854), .Y(
        \D_cache/n849 ) );
  CLKMX2X2 U5494 ( .A(\D_cache/cache[2][118] ), .B(n10217), .S0(n4803), .Y(
        \D_cache/n850 ) );
  CLKMX2X2 U5495 ( .A(\D_cache/cache[1][118] ), .B(n10217), .S0(n4780), .Y(
        \D_cache/n851 ) );
  MX2X1 U5496 ( .A(\D_cache/cache[0][118] ), .B(n10217), .S0(n4735), .Y(
        \D_cache/n852 ) );
  CLKMX2X2 U5497 ( .A(\D_cache/cache[7][102] ), .B(n10081), .S0(n5004), .Y(
        \D_cache/n973 ) );
  CLKMX2X2 U5498 ( .A(\D_cache/cache[6][102] ), .B(n10081), .S0(n4959), .Y(
        \D_cache/n974 ) );
  CLKMX2X2 U5499 ( .A(\D_cache/cache[5][102] ), .B(n10081), .S0(n4944), .Y(
        \D_cache/n975 ) );
  CLKMX2X2 U5500 ( .A(\D_cache/cache[4][102] ), .B(n10081), .S0(n4894), .Y(
        \D_cache/n976 ) );
  CLKMX2X2 U5501 ( .A(\D_cache/cache[3][102] ), .B(n10081), .S0(n4848), .Y(
        \D_cache/n977 ) );
  CLKMX2X2 U5502 ( .A(\D_cache/cache[2][102] ), .B(n10081), .S0(n4803), .Y(
        \D_cache/n978 ) );
  CLKMX2X2 U5503 ( .A(\D_cache/cache[1][102] ), .B(n10081), .S0(n4780), .Y(
        \D_cache/n979 ) );
  MX2X1 U5504 ( .A(\D_cache/cache[0][102] ), .B(n10081), .S0(n4734), .Y(
        \D_cache/n980 ) );
  NAND3BX2 U5505 ( .AN(n10583), .B(n10582), .C(n10581), .Y(\i_MIPS/PC/n63 ) );
  MX2X1 U5506 ( .A(\D_cache/cache[6][117] ), .B(n10675), .S0(n4957), .Y(
        \D_cache/n854 ) );
  CLKMX2X2 U5507 ( .A(\D_cache/cache[7][117] ), .B(n10675), .S0(n5001), .Y(
        \D_cache/n853 ) );
  MXI2X4 U5508 ( .A(n10674), .B(n10673), .S0(n5516), .Y(n10675) );
  CLKMX2X2 U5509 ( .A(\D_cache/cache[7][116] ), .B(n10662), .S0(n5001), .Y(
        \D_cache/n861 ) );
  CLKMX2X2 U5510 ( .A(\D_cache/cache[6][116] ), .B(n10662), .S0(n4957), .Y(
        \D_cache/n862 ) );
  CLKMX2X2 U5511 ( .A(\D_cache/cache[5][116] ), .B(n10662), .S0(n4936), .Y(
        \D_cache/n863 ) );
  CLKMX2X2 U5512 ( .A(\D_cache/cache[4][116] ), .B(n10662), .S0(n4893), .Y(
        \D_cache/n864 ) );
  CLKMX2X2 U5513 ( .A(\D_cache/cache[3][116] ), .B(n10662), .S0(n4847), .Y(
        \D_cache/n865 ) );
  CLKMX2X2 U5514 ( .A(\D_cache/cache[2][116] ), .B(n10662), .S0(n4802), .Y(
        \D_cache/n866 ) );
  CLKMX2X2 U5515 ( .A(\D_cache/cache[1][116] ), .B(n10662), .S0(n4779), .Y(
        \D_cache/n867 ) );
  MX2X1 U5516 ( .A(\D_cache/cache[0][116] ), .B(n10662), .S0(n4733), .Y(
        \D_cache/n868 ) );
  CLKMX2X2 U5517 ( .A(\D_cache/cache[7][114] ), .B(n10516), .S0(n5001), .Y(
        \D_cache/n877 ) );
  CLKMX2X2 U5518 ( .A(\D_cache/cache[6][114] ), .B(n10516), .S0(n4957), .Y(
        \D_cache/n878 ) );
  CLKMX2X2 U5519 ( .A(\D_cache/cache[5][114] ), .B(n10516), .S0(n4943), .Y(
        \D_cache/n879 ) );
  CLKMX2X2 U5520 ( .A(\D_cache/cache[4][114] ), .B(n10516), .S0(n4893), .Y(
        \D_cache/n880 ) );
  CLKMX2X2 U5521 ( .A(\D_cache/cache[3][114] ), .B(n10516), .S0(n4847), .Y(
        \D_cache/n881 ) );
  CLKMX2X2 U5522 ( .A(\D_cache/cache[2][114] ), .B(n10516), .S0(n4802), .Y(
        \D_cache/n882 ) );
  CLKMX2X2 U5523 ( .A(\D_cache/cache[1][114] ), .B(n10516), .S0(n4779), .Y(
        \D_cache/n883 ) );
  MX2X1 U5524 ( .A(\D_cache/cache[0][114] ), .B(n10516), .S0(n4733), .Y(
        \D_cache/n884 ) );
  AO21X4 U5525 ( .A0(n9278), .A1(n9277), .B0(n9276), .Y(n9282) );
  AO22X4 U5526 ( .A0(mem_rdata_I[109]), .A1(n5540), .B0(n251), .B1(n11295), 
        .Y(n9693) );
  AO22X4 U5527 ( .A0(mem_rdata_I[13]), .A1(n5540), .B0(n252), .B1(n11199), .Y(
        n9698) );
  AO22X4 U5528 ( .A0(mem_rdata_I[45]), .A1(n5539), .B0(n253), .B1(n11231), .Y(
        n9708) );
  AO22X4 U5529 ( .A0(mem_rdata_I[77]), .A1(n5539), .B0(n249), .B1(n11263), .Y(
        n9703) );
  AO22X4 U5530 ( .A0(mem_rdata_I[79]), .A1(n5540), .B0(n251), .B1(n11265), .Y(
        n9653) );
  AOI2BB1X2 U5531 ( .A0N(net112336), .A1N(\i_MIPS/n356 ), .B0(n4523), .Y(n6687) );
  NAND2X8 U5532 ( .A(n8539), .B(n8736), .Y(n7536) );
  NAND2X2 U5533 ( .A(n8539), .B(n9265), .Y(n8727) );
  AOI21X2 U5534 ( .A0(\i_MIPS/ID_EX[78] ), .A1(n3813), .B0(n4082), .Y(
        net105781) );
  NAND2X8 U5535 ( .A(net128301), .B(n4444), .Y(n9461) );
  AOI211X4 U5536 ( .A0(net101908), .A1(n7467), .B0(n7466), .C0(n7465), .Y(
        n7551) );
  AO21X4 U5537 ( .A0(net99002), .A1(net99003), .B0(net111904), .Y(n4139) );
  AO21X4 U5538 ( .A0(n10526), .A1(n10525), .B0(net111904), .Y(net98352) );
  AO21X4 U5539 ( .A0(net99157), .A1(net112799), .B0(net111904), .Y(net99118)
         );
  AO21X4 U5540 ( .A0(n10222), .A1(n10221), .B0(net111904), .Y(n10548) );
  AO21X4 U5541 ( .A0(net98375), .A1(net112736), .B0(net111904), .Y(net98217)
         );
  AO21X4 U5542 ( .A0(net98380), .A1(net112786), .B0(net111904), .Y(net98550)
         );
  CLKMX2X2 U5543 ( .A(\D_cache/cache[6][124] ), .B(n10483), .S0(n4956), .Y(
        \D_cache/n798 ) );
  CLKMX2X2 U5544 ( .A(\D_cache/cache[7][124] ), .B(n10483), .S0(n5000), .Y(
        \D_cache/n797 ) );
  MXI2X4 U5545 ( .A(n10482), .B(n10481), .S0(n5514), .Y(n10483) );
  CLKMX2X2 U5546 ( .A(\D_cache/cache[7][123] ), .B(n10309), .S0(n5000), .Y(
        \D_cache/n805 ) );
  CLKMX2X2 U5547 ( .A(\D_cache/cache[6][123] ), .B(n10309), .S0(n4956), .Y(
        \D_cache/n806 ) );
  CLKMX2X2 U5548 ( .A(\D_cache/cache[5][123] ), .B(n10309), .S0(n4936), .Y(
        \D_cache/n807 ) );
  CLKMX2X2 U5549 ( .A(\D_cache/cache[4][123] ), .B(n10309), .S0(n4892), .Y(
        \D_cache/n808 ) );
  CLKMX2X2 U5550 ( .A(\D_cache/cache[3][123] ), .B(n10309), .S0(n4846), .Y(
        \D_cache/n809 ) );
  CLKMX2X2 U5551 ( .A(\D_cache/cache[2][123] ), .B(n10309), .S0(n4801), .Y(
        \D_cache/n810 ) );
  CLKMX2X2 U5552 ( .A(\D_cache/cache[1][123] ), .B(n10309), .S0(n4778), .Y(
        \D_cache/n811 ) );
  MX2X1 U5553 ( .A(\D_cache/cache[0][123] ), .B(n10309), .S0(n4732), .Y(
        \D_cache/n812 ) );
  CLKMX2X2 U5554 ( .A(\D_cache/cache[7][121] ), .B(n10499), .S0(n5000), .Y(
        \D_cache/n821 ) );
  CLKMX2X2 U5555 ( .A(\D_cache/cache[6][121] ), .B(n10499), .S0(n4956), .Y(
        \D_cache/n822 ) );
  CLKMX2X2 U5556 ( .A(\D_cache/cache[5][121] ), .B(n10499), .S0(n4944), .Y(
        \D_cache/n823 ) );
  CLKMX2X2 U5557 ( .A(\D_cache/cache[4][121] ), .B(n10499), .S0(n4892), .Y(
        \D_cache/n824 ) );
  CLKMX2X2 U5558 ( .A(\D_cache/cache[3][121] ), .B(n10499), .S0(n4846), .Y(
        \D_cache/n825 ) );
  CLKMX2X2 U5559 ( .A(\D_cache/cache[2][121] ), .B(n10499), .S0(n4801), .Y(
        \D_cache/n826 ) );
  CLKMX2X2 U5560 ( .A(\D_cache/cache[1][121] ), .B(n10499), .S0(n4778), .Y(
        \D_cache/n827 ) );
  MX2X1 U5561 ( .A(\D_cache/cache[0][121] ), .B(n10499), .S0(n4732), .Y(
        \D_cache/n828 ) );
  NAND2BX2 U5562 ( .AN(n5427), .B(n11191), .Y(n9931) );
  MX2X1 U5563 ( .A(\D_cache/cache[0][31] ), .B(n10870), .S0(n4736), .Y(
        \D_cache/n1548 ) );
  CLKMX2X2 U5564 ( .A(\D_cache/cache[1][31] ), .B(n10870), .S0(n4781), .Y(
        \D_cache/n1547 ) );
  CLKMX2X2 U5565 ( .A(\D_cache/cache[2][31] ), .B(n10870), .S0(n4805), .Y(
        \D_cache/n1546 ) );
  CLKMX2X2 U5566 ( .A(\D_cache/cache[3][31] ), .B(n10870), .S0(n4849), .Y(
        \D_cache/n1545 ) );
  CLKMX2X2 U5567 ( .A(\D_cache/cache[4][31] ), .B(n10870), .S0(n4900), .Y(
        \D_cache/n1544 ) );
  CLKMX2X2 U5568 ( .A(\D_cache/cache[5][31] ), .B(n10870), .S0(n4938), .Y(
        \D_cache/n1543 ) );
  CLKMX2X2 U5569 ( .A(\D_cache/cache[6][31] ), .B(n10870), .S0(n4959), .Y(
        \D_cache/n1542 ) );
  CLKMX2X2 U5570 ( .A(\D_cache/cache[7][31] ), .B(n10870), .S0(n5003), .Y(
        \D_cache/n1541 ) );
  MX2X1 U5571 ( .A(\D_cache/cache[0][14] ), .B(n10743), .S0(n4739), .Y(
        \D_cache/n1684 ) );
  CLKMX2X2 U5572 ( .A(\D_cache/cache[1][14] ), .B(n10743), .S0(n4784), .Y(
        \D_cache/n1683 ) );
  CLKMX2X2 U5573 ( .A(\D_cache/cache[5][14] ), .B(n10743), .S0(n4942), .Y(
        \D_cache/n1679 ) );
  MXI2X4 U5574 ( .A(n10742), .B(n10741), .S0(n5518), .Y(n10743) );
  MX2X1 U5575 ( .A(\D_cache/cache[1][13] ), .B(n10732), .S0(n4785), .Y(
        \D_cache/n1691 ) );
  MX2X1 U5576 ( .A(\D_cache/cache[5][13] ), .B(n10732), .S0(n4941), .Y(
        \D_cache/n1687 ) );
  MXI2X4 U5577 ( .A(n10731), .B(n10730), .S0(n5518), .Y(n10732) );
  CLKMX2X2 U5578 ( .A(\I_cache/cache[0][8] ), .B(n9997), .S0(n5095), .Y(n12723) );
  AO22X4 U5579 ( .A0(mem_rdata_I[35]), .A1(n5539), .B0(n250), .B1(n11221), .Y(
        n11172) );
  AO22X4 U5580 ( .A0(mem_rdata_I[67]), .A1(n5535), .B0(n251), .B1(n11253), .Y(
        n11168) );
  AO22X4 U5581 ( .A0(mem_rdata_I[99]), .A1(n5535), .B0(n252), .B1(n11285), .Y(
        n11167) );
  AOI222X2 U5582 ( .A0(net102431), .A1(net100585), .B0(n4086), .B1(n4087), 
        .C0(n4088), .C1(n4089), .Y(n4085) );
  OAI211X2 U5583 ( .A0(n4415), .A1(\i_MIPS/PC/n2 ), .B0(n10523), .C0(n10522), 
        .Y(\i_MIPS/PC/n34 ) );
  CLKMX2X2 U5584 ( .A(\D_cache/cache[7][122] ), .B(n10277), .S0(n5002), .Y(
        \D_cache/n813 ) );
  CLKMX2X2 U5585 ( .A(\D_cache/cache[6][122] ), .B(n10277), .S0(n4958), .Y(
        \D_cache/n814 ) );
  CLKMX2X2 U5586 ( .A(\D_cache/cache[5][122] ), .B(n10277), .S0(n4940), .Y(
        \D_cache/n815 ) );
  CLKMX2X2 U5587 ( .A(\D_cache/cache[4][122] ), .B(n10277), .S0(n4895), .Y(
        \D_cache/n816 ) );
  CLKMX2X2 U5588 ( .A(\D_cache/cache[3][122] ), .B(n10277), .S0(n4848), .Y(
        \D_cache/n817 ) );
  CLKMX2X2 U5589 ( .A(\D_cache/cache[2][122] ), .B(n10277), .S0(n4804), .Y(
        \D_cache/n818 ) );
  CLKMX2X2 U5590 ( .A(\D_cache/cache[1][122] ), .B(n10277), .S0(n4783), .Y(
        \D_cache/n819 ) );
  MX2X1 U5591 ( .A(\D_cache/cache[0][122] ), .B(n10277), .S0(n4735), .Y(
        \D_cache/n820 ) );
  CLKMX2X2 U5592 ( .A(\D_cache/cache[1][112] ), .B(n10296), .S0(n4780), .Y(
        \D_cache/n899 ) );
  CLKMX2X2 U5593 ( .A(\D_cache/cache[2][112] ), .B(n10296), .S0(n4803), .Y(
        \D_cache/n898 ) );
  CLKMX2X2 U5594 ( .A(\D_cache/cache[3][112] ), .B(n10296), .S0(n4847), .Y(
        \D_cache/n897 ) );
  CLKMX2X2 U5595 ( .A(\D_cache/cache[4][112] ), .B(n10296), .S0(n4894), .Y(
        \D_cache/n896 ) );
  CLKMX2X2 U5596 ( .A(\D_cache/cache[5][112] ), .B(n10296), .S0(n4937), .Y(
        \D_cache/n895 ) );
  CLKMX2X2 U5597 ( .A(\D_cache/cache[6][112] ), .B(n10296), .S0(n4960), .Y(
        \D_cache/n894 ) );
  CLKMX2X2 U5598 ( .A(\D_cache/cache[7][112] ), .B(n10296), .S0(n5002), .Y(
        \D_cache/n893 ) );
  CLKMX2X2 U5599 ( .A(\D_cache/cache[5][21] ), .B(n10669), .S0(n4936), .Y(
        \D_cache/n1623 ) );
  CLKMX2X2 U5600 ( .A(\D_cache/cache[4][21] ), .B(n10669), .S0(n4893), .Y(
        \D_cache/n1624 ) );
  CLKMX2X2 U5601 ( .A(\D_cache/cache[3][21] ), .B(n10669), .S0(n4847), .Y(
        \D_cache/n1625 ) );
  CLKMX2X2 U5602 ( .A(\D_cache/cache[2][21] ), .B(n10669), .S0(n4802), .Y(
        \D_cache/n1626 ) );
  CLKMX2X2 U5603 ( .A(\D_cache/cache[1][21] ), .B(n10669), .S0(n4779), .Y(
        \D_cache/n1627 ) );
  AO22X4 U5604 ( .A0(mem_rdata_I[26]), .A1(n5541), .B0(n253), .B1(n11212), .Y(
        n9563) );
  AO22X4 U5605 ( .A0(mem_rdata_I[14]), .A1(n5541), .B0(n250), .B1(n11200), .Y(
        n9604) );
  AO22X4 U5606 ( .A0(mem_rdata_I[58]), .A1(n5541), .B0(n251), .B1(n11244), .Y(
        n9564) );
  AO22X4 U5607 ( .A0(mem_rdata_I[46]), .A1(n5541), .B0(n249), .B1(n11232), .Y(
        n9609) );
  AO22X4 U5608 ( .A0(mem_rdata_I[90]), .A1(n5541), .B0(n253), .B1(n11276), .Y(
        n9562) );
  AO22X4 U5609 ( .A0(mem_rdata_I[84]), .A1(n5541), .B0(n251), .B1(n11270), .Y(
        n9624) );
  AO22X4 U5610 ( .A0(mem_rdata_I[78]), .A1(n5541), .B0(n252), .B1(n11264), .Y(
        n9599) );
  NAND2BX4 U5611 ( .AN(n8538), .B(n3770), .Y(n8726) );
  NAND4BX4 U5612 ( .AN(n4341), .B(n9505), .C(n9504), .D(n9503), .Y(n11436) );
  OAI211X2 U5613 ( .A0(n4415), .A1(\i_MIPS/PC/n3 ), .B0(n10528), .C0(n10527), 
        .Y(\i_MIPS/PC/n35 ) );
  NAND3BX2 U5614 ( .AN(n10809), .B(n10808), .C(n10807), .Y(\i_MIPS/PC/n41 ) );
  NAND4X2 U5615 ( .A(n9768), .B(n9767), .C(n9766), .D(n9765), .Y(n11262) );
  OA22XL U5616 ( .A0(n5300), .A1(n1579), .B0(n5255), .B1(n3161), .Y(n9916) );
  OAI21X4 U5617 ( .A0(net127702), .A1(net127703), .B0(net105787), .Y(net105600) );
  AOI32X2 U5618 ( .A0(n4079), .A1(net127933), .A2(n4081), .B0(n4080), .B1(
        \i_MIPS/ID_EX[75] ), .Y(n4075) );
  NAND4X2 U5619 ( .A(n4079), .B(n4080), .C(net127930), .D(n3813), .Y(n4078) );
  OAI221X4 U5620 ( .A0(\i_MIPS/ALUin1[9] ), .A1(net112364), .B0(
        \i_MIPS/ALUin1[8] ), .B1(net112346), .C0(net105043), .Y(net104864) );
  AOI211XL U5621 ( .A0(n4091), .A1(net102253), .B0(net127829), .C0(net127833), 
        .Y(n4084) );
  INVX1 U5622 ( .A(net103917), .Y(n4091) );
  MX2XL U5623 ( .A(\i_MIPS/n369 ), .B(\i_MIPS/n368 ), .S0(\i_MIPS/ID_EX[79] ), 
        .Y(net103917) );
  NAND2X8 U5624 ( .A(net101906), .B(net107804), .Y(net103076) );
  NAND2XL U5625 ( .A(net102427), .B(net103889), .Y(n4086) );
  NAND2XL U5626 ( .A(net102430), .B(net105034), .Y(n4089) );
  NAND4BX4 U5627 ( .AN(n4083), .B(net105006), .C(net105007), .D(net105008), 
        .Y(net97783) );
  NAND4X8 U5628 ( .A(net102782), .B(net102781), .C(net102784), .D(net102783), 
        .Y(net100399) );
  AO21X4 U5629 ( .A0(net99164), .A1(net99165), .B0(net111644), .Y(net105047)
         );
  XOR2X4 U5630 ( .A(n4103), .B(net97755), .Y(n4101) );
  CLKINVX8 U5631 ( .A(net105282), .Y(net97686) );
  OAI221X2 U5632 ( .A0(net105194), .A1(net111624), .B0(net105195), .B1(
        net111636), .C0(net105196), .Y(net97701) );
  NOR2X8 U5633 ( .A(n3922), .B(n4097), .Y(net102782) );
  XOR2X4 U5634 ( .A(n4098), .B(n4137), .Y(n4097) );
  AO21X4 U5635 ( .A0(net98776), .A1(net98777), .B0(net111642), .Y(net104253)
         );
  CLKMX2X3 U5636 ( .A(net104108), .B(net104109), .S0(net107812), .Y(net104105)
         );
  AO21X4 U5637 ( .A0(net98758), .A1(net98759), .B0(net111642), .Y(net104107)
         );
  AO21X4 U5638 ( .A0(net98758), .A1(net98759), .B0(net111904), .Y(net98755) );
  AO21X4 U5639 ( .A0(net98386), .A1(net98385), .B0(net111642), .Y(net104409)
         );
  CLKINVX6 U5640 ( .A(net104042), .Y(net98571) );
  AO21X4 U5641 ( .A0(net98340), .A1(net98341), .B0(net111904), .Y(net98514) );
  AO21X4 U5642 ( .A0(net98340), .A1(net98341), .B0(net111642), .Y(net103251)
         );
  AO21X4 U5643 ( .A0(net98335), .A1(net98336), .B0(net111642), .Y(net103091)
         );
  OAI31X2 U5644 ( .A0(n11), .A1(net100403), .A2(net100399), .B0(net100404), 
        .Y(net100402) );
  NAND3BX4 U5645 ( .AN(net100399), .B(net100396), .C(n3917), .Y(net100400) );
  CLKMX2X2 U5646 ( .A(n4105), .B(n4106), .S0(\i_MIPS/IR_ID[25] ), .Y(n4104) );
  NOR4X1 U5647 ( .A(n4116), .B(n4117), .C(n4118), .D(n4119), .Y(n4105) );
  NAND4X1 U5648 ( .A(n4121), .B(n4122), .C(n4123), .D(n4124), .Y(n4116) );
  OA22X1 U5649 ( .A0(\i_MIPS/Register/register[1][2] ), .A1(net112258), .B0(
        \i_MIPS/Register/register[9][2] ), .B1(n147), .Y(n4121) );
  OA22X1 U5650 ( .A0(\i_MIPS/Register/register[5][2] ), .A1(n192), .B0(
        \i_MIPS/Register/register[13][2] ), .B1(net112236), .Y(n4122) );
  OA22XL U5651 ( .A0(\i_MIPS/Register/register[3][2] ), .A1(net112182), .B0(
        \i_MIPS/Register/register[11][2] ), .B1(n197), .Y(n4123) );
  OA22X1 U5652 ( .A0(\i_MIPS/Register/register[7][2] ), .A1(net112152), .B0(
        \i_MIPS/Register/register[15][2] ), .B1(net112164), .Y(n4124) );
  INVX8 U5653 ( .A(net112178), .Y(net112164) );
  OAI221XL U5654 ( .A0(\i_MIPS/Register/register[2][2] ), .A1(net112072), .B0(
        \i_MIPS/Register/register[10][2] ), .B1(net112090), .C0(n4120), .Y(
        n4117) );
  OA22X1 U5655 ( .A0(\i_MIPS/Register/register[6][2] ), .A1(net112110), .B0(
        \i_MIPS/Register/register[14][2] ), .B1(net112128), .Y(n4120) );
  BUFX8 U5656 ( .A(net112112), .Y(net112110) );
  BUFX8 U5657 ( .A(net112138), .Y(net112128) );
  AO22X1 U5658 ( .A0(net112036), .A1(n938), .B0(net100603), .B1(n2448), .Y(
        n4118) );
  BUFX8 U5659 ( .A(net112032), .Y(net112018) );
  NAND4X1 U5660 ( .A(n4112), .B(n4113), .C(n4114), .D(n4115), .Y(n4107) );
  OA22X1 U5661 ( .A0(\i_MIPS/Register/register[17][2] ), .A1(net112254), .B0(
        \i_MIPS/Register/register[25][2] ), .B1(n151), .Y(n4112) );
  OA22X1 U5662 ( .A0(\i_MIPS/Register/register[21][2] ), .A1(n192), .B0(
        \i_MIPS/Register/register[29][2] ), .B1(net112240), .Y(n4113) );
  OA22XL U5663 ( .A0(\i_MIPS/Register/register[19][2] ), .A1(net112182), .B0(
        \i_MIPS/Register/register[27][2] ), .B1(n200), .Y(n4114) );
  OA22X1 U5664 ( .A0(\i_MIPS/Register/register[23][2] ), .A1(net112152), .B0(
        \i_MIPS/Register/register[31][2] ), .B1(net112164), .Y(n4115) );
  OAI221XL U5665 ( .A0(\i_MIPS/Register/register[18][2] ), .A1(net112072), 
        .B0(\i_MIPS/Register/register[26][2] ), .B1(net112090), .C0(n4111), 
        .Y(n4108) );
  OA22X1 U5666 ( .A0(\i_MIPS/Register/register[22][2] ), .A1(net112110), .B0(
        \i_MIPS/Register/register[30][2] ), .B1(net112128), .Y(n4111) );
  AO22X1 U5667 ( .A0(net112036), .A1(n939), .B0(net100603), .B1(n2449), .Y(
        n4109) );
  AND2XL U5668 ( .A(n3420), .B(n4139), .Y(net129005) );
  INVX1 U5669 ( .A(net104229), .Y(n4125) );
  OAI221X4 U5670 ( .A0(net112350), .A1(\i_MIPS/n371 ), .B0(net112334), .B1(
        \i_MIPS/n369 ), .C0(net103919), .Y(net101401) );
  CLKMX2X2 U5671 ( .A(net100573), .B(net112438), .S0(n4128), .Y(net105008) );
  AND2XL U5672 ( .A(net105676), .B(\i_MIPS/n369 ), .Y(n4128) );
  MX2XL U5673 ( .A(net112962), .B(net97783), .S0(n216), .Y(\i_MIPS/n467 ) );
  AND2XL U5674 ( .A(net98499), .B(net98500), .Y(net129017) );
  NAND4X1 U5675 ( .A(net99633), .B(net99634), .C(net99635), .D(net99636), .Y(
        net98496) );
  CLKAND2X12 U5676 ( .A(net97444), .B(\i_MIPS/n236 ), .Y(n4141) );
  NOR2X8 U5677 ( .A(net105349), .B(net105350), .Y(net100398) );
  NAND4X8 U5678 ( .A(net129200), .B(net100415), .C(net100416), .D(net100417), 
        .Y(net100401) );
  AOI31X2 U5679 ( .A0(net97452), .A1(\i_MIPS/n567 ), .A2(\i_MIPS/IF_ID[97] ), 
        .B0(net112406), .Y(net100404) );
  OA22X2 U5680 ( .A0(n10747), .A1(n4245), .B0(n10750), .B1(n4246), .Y(n7661)
         );
  INVX3 U5681 ( .A(n11364), .Y(n10747) );
  NAND2X2 U5682 ( .A(\i_MIPS/ALUin1[1] ), .B(n4671), .Y(net103919) );
  BUFX20 U5683 ( .A(n9987), .Y(n4884) );
  AOI222X1 U5684 ( .A0(n5512), .A1(n11384), .B0(mem_rdata_D[34]), .B1(n232), 
        .C0(n12985), .C1(n5507), .Y(n10938) );
  OR2X8 U5685 ( .A(n4439), .B(net111640), .Y(n4189) );
  NAND4X2 U5686 ( .A(n8244), .B(n8243), .C(n8851), .D(n8242), .Y(n8245) );
  NAND2X4 U5687 ( .A(\i_MIPS/ALUin1[23] ), .B(n6563), .Y(n8848) );
  OA22X1 U5688 ( .A0(\i_MIPS/ALUin1[23] ), .A1(n4670), .B0(\i_MIPS/ALUin1[24] ), .B1(n3829), .Y(n8248) );
  INVX4 U5689 ( .A(n6520), .Y(n9066) );
  OR3X8 U5690 ( .A(n3676), .B(n10334), .C(n10445), .Y(n10570) );
  XNOR2X4 U5691 ( .A(n11502), .B(n12933), .Y(n6437) );
  OAI221X4 U5692 ( .A0(n4660), .A1(n8650), .B0(n4659), .B1(n3844), .C0(n8648), 
        .Y(n9053) );
  NOR4X1 U5693 ( .A(n11065), .B(n11051), .C(n270), .D(n11060), .Y(n11048) );
  NAND2X6 U5694 ( .A(n10814), .B(n10812), .Y(n10386) );
  XOR3X2 U5695 ( .A(n10814), .B(n10813), .C(n10812), .Y(n10817) );
  OA22X4 U5696 ( .A0(n10687), .A1(n4245), .B0(n10690), .B1(n4246), .Y(n8203)
         );
  NAND3BX4 U5697 ( .AN(n6969), .B(n4420), .C(n4388), .Y(n7411) );
  NAND2X6 U5698 ( .A(\i_MIPS/ALUin1[7] ), .B(n6531), .Y(n7880) );
  NAND2X4 U5699 ( .A(n7106), .B(n7105), .Y(n4152) );
  NAND4X4 U5700 ( .A(n7351), .B(n7350), .C(n7349), .D(n7348), .Y(n11424) );
  OA22X2 U5701 ( .A0(n4980), .A1(n766), .B0(n5026), .B1(n2328), .Y(n7348) );
  MX2X2 U5702 ( .A(n8915), .B(n8914), .S0(net107810), .Y(n8917) );
  NAND4BX2 U5703 ( .AN(n8904), .B(n8903), .C(n8902), .D(n8901), .Y(n8915) );
  NAND4BX2 U5704 ( .AN(n8913), .B(n8912), .C(n8911), .D(n8910), .Y(n8914) );
  NAND4X4 U5705 ( .A(n8366), .B(n8365), .C(n8364), .D(n8363), .Y(n10965) );
  AOI222X2 U5706 ( .A0(n8346), .A1(net100585), .B0(n8345), .B1(n8344), .C0(
        n8343), .C1(n8342), .Y(n8366) );
  OAI211X4 U5707 ( .A0(n8180), .A1(n8179), .B0(n8178), .C0(n8177), .Y(n8184)
         );
  AO21X4 U5708 ( .A0(n7021), .A1(n7020), .B0(n5546), .Y(n10064) );
  NAND4X6 U5709 ( .A(n6015), .B(n6014), .C(n6013), .D(n6012), .Y(n11326) );
  CLKMX2X2 U5710 ( .A(\D_cache/cache[0][101] ), .B(n10986), .S0(n4739), .Y(
        \D_cache/n988 ) );
  CLKMX2X2 U5711 ( .A(\D_cache/cache[7][101] ), .B(n10986), .S0(n5009), .Y(
        \D_cache/n981 ) );
  BUFX4 U5712 ( .A(n4839), .Y(n4832) );
  AOI2BB1X4 U5713 ( .A0N(n10434), .A1N(n10433), .B0(n10432), .Y(n10436) );
  NAND4X4 U5714 ( .A(n6087), .B(n6086), .C(n6085), .D(n6084), .Y(n11332) );
  CLKAND2X12 U5715 ( .A(n4657), .B(n11313), .Y(mem_wdata_I[127]) );
  BUFX12 U5716 ( .A(n10998), .Y(n5503) );
  NAND3BX4 U5717 ( .AN(n4295), .B(n4664), .C(n4666), .Y(n9991) );
  NAND3BX4 U5718 ( .AN(n8161), .B(n4658), .C(n8160), .Y(n8170) );
  AO21X4 U5719 ( .A0(n3884), .A1(n8349), .B0(n4449), .Y(n8159) );
  NAND4X4 U5720 ( .A(n7906), .B(n7908), .C(n7907), .D(n7909), .Y(net97834) );
  OAI221X2 U5721 ( .A0(net112366), .A1(\i_MIPS/n371 ), .B0(net112350), .B1(
        \i_MIPS/n370 ), .C0(n6685), .Y(n7898) );
  AO21X4 U5722 ( .A0(n7803), .A1(n4570), .B0(n7806), .Y(n7172) );
  OA22X2 U5723 ( .A0(n4765), .A1(n3029), .B0(n4796), .B1(n848), .Y(n6342) );
  NAND4X4 U5724 ( .A(n6342), .B(n6341), .C(n6340), .D(n6339), .Y(n11483) );
  MXI2X4 U5725 ( .A(n10264), .B(n10263), .S0(n5514), .Y(n10265) );
  AND3X2 U5726 ( .A(net111994), .B(net102573), .C(n8259), .Y(n8272) );
  OAI221X4 U5727 ( .A0(n9663), .A1(n4247), .B0(n9662), .B1(n5427), .C0(n9661), 
        .Y(n4571) );
  AOI2BB1X2 U5728 ( .A0N(\i_MIPS/ALUin1[17] ), .A1N(n3828), .B0(n4463), .Y(
        n7823) );
  AND2X4 U5729 ( .A(n4672), .B(\i_MIPS/n355 ), .Y(n4463) );
  OAI211X4 U5730 ( .A0(\i_MIPS/ALUin1[15] ), .A1(net112350), .B0(n7824), .C0(
        n7823), .Y(n8155) );
  INVXL U5731 ( .A(n7694), .Y(n7703) );
  NAND3BX4 U5732 ( .AN(n6503), .B(n7708), .C(n7684), .Y(n6511) );
  OAI221X2 U5733 ( .A0(n8629), .A1(net111622), .B0(n3405), .B1(net111634), 
        .C0(n8628), .Y(n10651) );
  OA22X2 U5734 ( .A0(n4835), .A1(n768), .B0(n4880), .B1(n2330), .Y(n6379) );
  AOI222X2 U5735 ( .A0(n5498), .A1(n11424), .B0(mem_rdata_D[74]), .B1(n234), 
        .C0(n12977), .C1(n4385), .Y(n10261) );
  AO21X4 U5736 ( .A0(net112400), .A1(n10828), .B0(n4467), .Y(n10575) );
  OA22X2 U5737 ( .A0(n4970), .A1(n696), .B0(n5015), .B1(n2265), .Y(n8881) );
  OA22X2 U5738 ( .A0(n4817), .A1(n697), .B0(n4863), .B1(n2266), .Y(n8883) );
  AO21X4 U5739 ( .A0(n7361), .A1(n7360), .B0(n3697), .Y(net98759) );
  BUFX20 U5740 ( .A(n4774), .Y(n4767) );
  CLKAND2X4 U5741 ( .A(n3745), .B(n4392), .Y(n4384) );
  AOI32X2 U5742 ( .A0(net103079), .A1(\i_MIPS/ALUin1[1] ), .A2(net112338), 
        .B0(n7970), .B1(\i_MIPS/ALUin1[1] ), .Y(n7971) );
  OA22X4 U5743 ( .A0(n4669), .A1(\i_MIPS/n353 ), .B0(net112332), .B1(
        \i_MIPS/n354 ), .Y(n6766) );
  OA22X4 U5744 ( .A0(net101914), .A1(n7968), .B0(net102405), .B1(n7967), .Y(
        n7972) );
  NAND4X4 U5745 ( .A(n8016), .B(n8015), .C(n8014), .D(n8013), .Y(n11415) );
  BUFX4 U5746 ( .A(n4799), .Y(n4787) );
  AOI222X2 U5747 ( .A0(n5495), .A1(n11468), .B0(mem_rdata_D[118]), .B1(n236), 
        .C0(n12965), .C1(n5494), .Y(n10210) );
  MXI2X4 U5748 ( .A(n10210), .B(n10209), .S0(n5513), .Y(n10211) );
  INVX3 U5749 ( .A(n3841), .Y(n6563) );
  INVX4 U5750 ( .A(net111642), .Y(net112782) );
  AO22X1 U5751 ( .A0(net100583), .A1(n9281), .B0(n9244), .B1(net100585), .Y(
        n9261) );
  OA22X4 U5752 ( .A0(n4763), .A1(n2150), .B0(n4795), .B1(n571), .Y(n6392) );
  AOI32X4 U5753 ( .A0(net97444), .A1(n10579), .A2(n10797), .B0(
        \i_MIPS/IF_ID_28 ), .B1(net108682), .Y(n10359) );
  AOI2BB1X4 U5754 ( .A0N(n4467), .A1N(n10825), .B0(n10824), .Y(n10826) );
  OA22X2 U5755 ( .A0(n5372), .A1(n769), .B0(n5348), .B1(n2331), .Y(n10179) );
  OAI221X1 U5756 ( .A0(\i_MIPS/Register/register[2][23] ), .A1(n4690), .B0(
        \i_MIPS/Register/register[10][23] ), .B1(n4685), .C0(n8896), .Y(n8904)
         );
  OAI221X2 U5757 ( .A0(n7717), .A1(n7716), .B0(n7715), .B1(n7714), .C0(n7713), 
        .Y(net98046) );
  NAND2BX4 U5758 ( .AN(n5425), .B(n11253), .Y(n10202) );
  NAND4X4 U5759 ( .A(n10186), .B(n10185), .C(n10184), .D(n10183), .Y(n11253)
         );
  OA22X1 U5760 ( .A0(n5392), .A1(n1225), .B0(n5348), .B1(n2762), .Y(n10183) );
  OA22X4 U5761 ( .A0(n10899), .A1(n4245), .B0(n10902), .B1(n4246), .Y(n7105)
         );
  NAND4X2 U5762 ( .A(n7100), .B(n7099), .C(n7098), .D(n7097), .Y(n11358) );
  OA22X1 U5763 ( .A0(n4982), .A1(n1226), .B0(n5028), .B1(n2763), .Y(n7097) );
  NAND4X4 U5764 ( .A(n8494), .B(n8493), .C(n8492), .D(n8491), .Y(n11442) );
  NAND2X4 U5765 ( .A(n9568), .B(n4060), .Y(n6120) );
  AO22X1 U5766 ( .A0(ICACHE_addr[25]), .A1(n11512), .B0(mem_write_I), .B1(
        n11340), .Y(n12808) );
  AO22X1 U5767 ( .A0(ICACHE_addr[16]), .A1(n11512), .B0(mem_write_I), .B1(
        n11331), .Y(n12817) );
  AO22X1 U5768 ( .A0(ICACHE_addr[21]), .A1(n11512), .B0(mem_write_I), .B1(
        n11336), .Y(n12812) );
  NAND4X1 U5769 ( .A(n7807), .B(n7820), .C(net112292), .D(n8753), .Y(n7834) );
  BUFX12 U5770 ( .A(n5509), .Y(n5512) );
  CLKMX2X3 U5771 ( .A(n7342), .B(n7341), .S0(net107816), .Y(n7343) );
  NAND4X4 U5772 ( .A(n9783), .B(n9782), .C(n9781), .D(n9780), .Y(n10406) );
  NAND2BX1 U5773 ( .AN(n4247), .B(n11294), .Y(n9783) );
  OA22X2 U5774 ( .A0(n5115), .A1(n698), .B0(n5081), .B1(n2267), .Y(n9778) );
  NAND4X8 U5775 ( .A(n5996), .B(n5995), .C(n5994), .D(n5993), .Y(n11338) );
  OAI221X2 U5776 ( .A0(\i_MIPS/n340 ), .A1(net112366), .B0(\i_MIPS/n341 ), 
        .B1(net112346), .C0(n6840), .Y(n7472) );
  CLKINVX4 U5777 ( .A(n8228), .Y(n8534) );
  OA21X4 U5778 ( .A0(n10420), .A1(n10419), .B0(n3658), .Y(n4319) );
  XNOR2X4 U5779 ( .A(ICACHE_addr[8]), .B(n11323), .Y(n6008) );
  AO22X4 U5780 ( .A0(mem_rdata_I[98]), .A1(n5535), .B0(n252), .B1(n11284), .Y(
        n11102) );
  OA22X4 U5781 ( .A0(n4669), .A1(\i_MIPS/n367 ), .B0(net112336), .B1(
        \i_MIPS/n366 ), .Y(n6769) );
  AO21X4 U5782 ( .A0(n7854), .A1(n7853), .B0(n3729), .Y(net98341) );
  CLKMX2X2 U5783 ( .A(\D_cache/cache[0][47] ), .B(n10757), .S0(n4739), .Y(
        \D_cache/n1420 ) );
  BUFX8 U5784 ( .A(n4385), .Y(n5497) );
  AO21X4 U5785 ( .A0(net112356), .A1(\i_MIPS/ALU/N303 ), .B0(n6772), .Y(n9154)
         );
  INVX8 U5786 ( .A(n11454), .Y(n10893) );
  NAND4X4 U5787 ( .A(n7092), .B(n7091), .C(n7090), .D(n7089), .Y(n11454) );
  INVX2 U5788 ( .A(n7172), .Y(n7156) );
  OAI222X2 U5789 ( .A0(n4439), .A1(net111902), .B0(n6603), .B1(net101978), 
        .C0(n6640), .C1(net100682), .Y(n10150) );
  AO21X4 U5790 ( .A0(n6439), .A1(n6438), .B0(n3665), .Y(n10788) );
  OA22X4 U5791 ( .A0(n4835), .A1(n2154), .B0(n4880), .B1(n575), .Y(n6383) );
  AOI222X2 U5792 ( .A0(n5495), .A1(n11473), .B0(mem_rdata_D[123]), .B1(n234), 
        .C0(n12960), .C1(n5494), .Y(n10302) );
  MXI2X4 U5793 ( .A(n10302), .B(n10301), .S0(n5515), .Y(n10303) );
  NAND2X2 U5794 ( .A(n7900), .B(n4536), .Y(n8876) );
  CLKMX2X4 U5795 ( .A(n7087), .B(n7086), .S0(net107816), .Y(n7088) );
  OA22X4 U5796 ( .A0(n4764), .A1(n3370), .B0(n4796), .B1(n1741), .Y(n4327) );
  OA22X4 U5797 ( .A0(n4764), .A1(n3371), .B0(n4796), .B1(n1742), .Y(n4328) );
  OA22X4 U5798 ( .A0(n4764), .A1(n3004), .B0(n4796), .B1(n576), .Y(n6350) );
  AO22X2 U5799 ( .A0(n9531), .A1(n645), .B0(n4715), .B1(n2220), .Y(n9201) );
  AO22X1 U5800 ( .A0(n9531), .A1(n988), .B0(n4716), .B1(n2509), .Y(n9106) );
  AO22X1 U5801 ( .A0(n9531), .A1(n989), .B0(n4714), .B1(n2510), .Y(n9097) );
  BUFX20 U5802 ( .A(n11513), .Y(n5554) );
  NAND2BX1 U5803 ( .AN(n4247), .B(n11292), .Y(n10063) );
  NAND2X6 U5804 ( .A(n4499), .B(n4447), .Y(net102051) );
  AOI2BB1X1 U5805 ( .A0N(\i_MIPS/IF_ID[97] ), .A1N(net97452), .B0(net112406), 
        .Y(n11042) );
  MXI2X4 U5806 ( .A(n10068), .B(n10067), .S0(n5513), .Y(n10069) );
  NAND2X6 U5807 ( .A(n4505), .B(n4502), .Y(n9410) );
  NAND4X2 U5808 ( .A(n9750), .B(n9749), .C(n9748), .D(n9747), .Y(n11197) );
  CLKMX2X2 U5809 ( .A(\D_cache/cache[0][26] ), .B(n10271), .S0(n4735), .Y(
        \D_cache/n1588 ) );
  CLKMX2X2 U5810 ( .A(\D_cache/cache[7][26] ), .B(n10271), .S0(n5002), .Y(
        \D_cache/n1581 ) );
  MXI2X4 U5811 ( .A(n10270), .B(n10269), .S0(n5514), .Y(n10271) );
  AOI222X4 U5812 ( .A0(n5495), .A1(n11464), .B0(mem_rdata_D[114]), .B1(n234), 
        .C0(n12969), .C1(n5494), .Y(n10509) );
  MXI2X6 U5813 ( .A(n10509), .B(n10508), .S0(n5516), .Y(n10510) );
  CLKMX2X2 U5814 ( .A(\D_cache/cache[0][16] ), .B(n10290), .S0(n4735), .Y(
        \D_cache/n1668 ) );
  OA22X4 U5815 ( .A0(n4763), .A1(n2155), .B0(n4796), .B1(n578), .Y(n6380) );
  INVX3 U5816 ( .A(n8860), .Y(n8858) );
  NOR2X4 U5817 ( .A(n8853), .B(n9481), .Y(n8856) );
  NOR2X2 U5818 ( .A(n7164), .B(n4451), .Y(n7158) );
  NAND2X4 U5819 ( .A(\i_MIPS/ALUin1[12] ), .B(n6550), .Y(n7523) );
  AOI222X4 U5820 ( .A0(n5495), .A1(n11471), .B0(mem_rdata_D[121]), .B1(n233), 
        .C0(n12962), .C1(n5494), .Y(n10492) );
  MXI2X6 U5821 ( .A(n10492), .B(n10491), .S0(n5515), .Y(n10493) );
  INVX4 U5822 ( .A(n8353), .Y(n8958) );
  INVX8 U5823 ( .A(n11390), .Y(n10902) );
  AOI222X4 U5824 ( .A0(n5495), .A1(n11456), .B0(mem_rdata_D[106]), .B1(n236), 
        .C0(n12977), .C1(n5494), .Y(n10258) );
  MXI2X6 U5825 ( .A(n10258), .B(n10257), .S0(n5515), .Y(n10259) );
  OAI31X2 U5826 ( .A0(n7514), .A1(n7513), .A2(n7512), .B0(n7511), .Y(n7519) );
  OAI221X2 U5827 ( .A0(n9220), .A1(net111622), .B0(n9219), .B1(net111634), 
        .C0(n9218), .Y(n10666) );
  OAI31X4 U5828 ( .A0(n7522), .A1(n7521), .A2(n7881), .B0(n7524), .Y(n7533) );
  AOI2BB1X2 U5829 ( .A0N(net102428), .A1N(n7505), .B0(n7504), .Y(n7506) );
  AOI222X2 U5830 ( .A0(n5496), .A1(n11470), .B0(mem_rdata_D[120]), .B1(n232), 
        .C0(n12963), .C1(n5493), .Y(n10777) );
  MXI2X4 U5831 ( .A(n10777), .B(n10776), .S0(n5519), .Y(n10778) );
  NAND4X4 U5832 ( .A(n6310), .B(n6309), .C(n6308), .D(n6307), .Y(n6311) );
  AOI222X4 U5833 ( .A0(n5500), .A1(n11416), .B0(mem_rdata_D[66]), .B1(n235), 
        .C0(n12985), .C1(n4385), .Y(n10932) );
  OA22X1 U5834 ( .A0(n5372), .A1(n1227), .B0(n5329), .B1(n2764), .Y(n6048) );
  XNOR2X4 U5835 ( .A(ICACHE_addr[10]), .B(n11325), .Y(n6030) );
  CLKMX2X2 U5836 ( .A(\D_cache/cache[0][17] ), .B(n10765), .S0(n4736), .Y(
        \D_cache/n1660 ) );
  MXI2X4 U5837 ( .A(n10764), .B(n10763), .S0(n5519), .Y(n10765) );
  OA22X4 U5838 ( .A0(n5287), .A1(n2156), .B0(n5255), .B1(n579), .Y(n6085) );
  OA22X4 U5839 ( .A0(n5287), .A1(n2158), .B0(n5255), .B1(n581), .Y(n6097) );
  NAND2X1 U5840 ( .A(n6612), .B(n4500), .Y(n9525) );
  INVX1 U5841 ( .A(n7523), .Y(n7687) );
  XOR2X4 U5842 ( .A(n10342), .B(ICACHE_addr[25]), .Y(n10839) );
  NAND2X4 U5843 ( .A(n10228), .B(n10810), .Y(n10385) );
  OAI33X2 U5844 ( .A0(n3899), .A1(n9338), .A2(n8435), .B0(n8436), .B1(n8434), 
        .B2(net101257), .Y(n8464) );
  XNOR2X4 U5845 ( .A(n11504), .B(n12931), .Y(n6436) );
  OA22X4 U5846 ( .A0(n4836), .A1(n3007), .B0(n4882), .B1(n583), .Y(n6349) );
  MXI2X4 U5847 ( .A(n10753), .B(n10752), .S0(n5519), .Y(n10754) );
  AO21X4 U5848 ( .A0(n6757), .A1(net105038), .B0(n6756), .Y(n6962) );
  AOI2BB1X4 U5849 ( .A0N(n3771), .A1N(n3824), .B0(n6510), .Y(n6503) );
  AOI2BB2X4 U5850 ( .B0(n6582), .B1(n6581), .A0N(n6584), .A1N(n6583), .Y(n4151) );
  XNOR2X4 U5851 ( .A(ICACHE_addr[11]), .B(n11326), .Y(n6031) );
  AOI222X2 U5852 ( .A0(n5496), .A1(n11453), .B0(mem_rdata_D[103]), .B1(n233), 
        .C0(n12980), .C1(n5493), .Y(n10882) );
  MXI2X4 U5853 ( .A(n10882), .B(n10881), .S0(n5520), .Y(n10883) );
  OA22X4 U5854 ( .A0(n10934), .A1(n4245), .B0(n10937), .B1(n4246), .Y(n6940)
         );
  OA22X2 U5855 ( .A0(n4983), .A1(n774), .B0(n5029), .B1(n2336), .Y(n6936) );
  NAND3BX2 U5856 ( .AN(n10443), .B(n10442), .C(n10441), .Y(\i_MIPS/PC/n51 ) );
  NAND2BX1 U5857 ( .AN(n4247), .B(n11287), .Y(n9933) );
  OAI211X2 U5858 ( .A0(n8079), .A1(n6517), .B0(n6516), .C0(n4436), .Y(n8939)
         );
  XNOR2X1 U5859 ( .A(ICACHE_addr[28]), .B(n11343), .Y(n6103) );
  NAND4X2 U5860 ( .A(n6102), .B(n6101), .C(n6100), .D(n6099), .Y(n11343) );
  NAND2X2 U5861 ( .A(n7516), .B(n8630), .Y(n7518) );
  NAND2X4 U5862 ( .A(\i_MIPS/ALUin1[9] ), .B(n3687), .Y(n8630) );
  NAND2X4 U5863 ( .A(\i_MIPS/ALUin1[3] ), .B(n6541), .Y(n8339) );
  NAND2X6 U5864 ( .A(n6586), .B(\i_MIPS/n346 ), .Y(n9043) );
  MXI2X4 U5865 ( .A(\i_MIPS/ID_EX[66] ), .B(\i_MIPS/ID_EX[98] ), .S0(n3635), 
        .Y(n6590) );
  OAI221X2 U5866 ( .A0(n4498), .A1(net101413), .B0(net101257), .B1(n4298), 
        .C0(net112420), .Y(n7981) );
  AOI222X2 U5867 ( .A0(n5496), .A1(n11475), .B0(mem_rdata_D[125]), .B1(n232), 
        .C0(n12958), .C1(n5493), .Y(n10682) );
  MXI2X4 U5868 ( .A(n10682), .B(n10681), .S0(n5517), .Y(n10683) );
  MXI2X4 U5869 ( .A(n10708), .B(n10707), .S0(n5517), .Y(n10709) );
  NAND4X4 U5870 ( .A(n7104), .B(n7103), .C(n7102), .D(n7101), .Y(n11390) );
  XNOR2X2 U5871 ( .A(ICACHE_addr[21]), .B(n11336), .Y(n6095) );
  OA22X2 U5872 ( .A0(n5101), .A1(n776), .B0(n5060), .B1(n2338), .Y(n6023) );
  XNOR2X4 U5873 ( .A(n4325), .B(n3802), .Y(n8531) );
  XNOR2X2 U5874 ( .A(ICACHE_addr[16]), .B(n11331), .Y(n6094) );
  NAND4X4 U5875 ( .A(n5990), .B(n5989), .C(n5988), .D(n5987), .Y(n11335) );
  NAND3BX4 U5876 ( .AN(net105600), .B(n4394), .C(net103913), .Y(n6753) );
  AO21X4 U5877 ( .A0(n10561), .A1(n10560), .B0(net111640), .Y(n8722) );
  NAND4X4 U5878 ( .A(n8687), .B(n8686), .C(n8685), .D(n8684), .Y(n11455) );
  OA22XL U5879 ( .A0(n4746), .A1(n1293), .B0(n4790), .B1(n2824), .Y(n8687) );
  XNOR2X4 U5880 ( .A(ICACHE_addr[25]), .B(n11340), .Y(n6060) );
  MX2XL U5881 ( .A(net112415), .B(net101082), .S0(n8656), .Y(n8657) );
  OAI2BB1X4 U5882 ( .A0N(n7685), .A1N(n7684), .B0(n7683), .Y(n7686) );
  AOI21X4 U5883 ( .A0(n6502), .A1(n6501), .B0(n7046), .Y(n7404) );
  AO21X4 U5884 ( .A0(n9349), .A1(n9330), .B0(n7480), .Y(n8450) );
  NAND2X4 U5885 ( .A(n6588), .B(\i_MIPS/n344 ), .Y(n9330) );
  OA22X4 U5886 ( .A0(n10681), .A1(n4675), .B0(n10684), .B1(n4250), .Y(n8204)
         );
  XOR2X4 U5887 ( .A(n10332), .B(ICACHE_addr[22]), .Y(n10456) );
  NAND2X2 U5888 ( .A(net98662), .B(ICACHE_addr[21]), .Y(n10332) );
  AO21X4 U5889 ( .A0(n10504), .A1(n10503), .B0(net111902), .Y(n10519) );
  OAI221X2 U5890 ( .A0(n3690), .A1(n4524), .B0(mem_ready_D), .B1(n9), .C0(
        n9981), .Y(n10083) );
  NAND3BX2 U5891 ( .AN(n9980), .B(n5548), .C(DCACHE_ren), .Y(n9981) );
  AOI211X4 U5892 ( .A0(n4436), .A1(n8535), .B0(n9142), .C0(n8230), .Y(n8233)
         );
  NOR4X2 U5893 ( .A(n7569), .B(n7568), .C(n7567), .D(n7566), .Y(n7570) );
  OA22XL U5894 ( .A0(\i_MIPS/Register/register[22][8] ), .A1(net112112), .B0(
        \i_MIPS/Register/register[30][8] ), .B1(net112142), .Y(n7081) );
  OA22XL U5895 ( .A0(\i_MIPS/Register/register[6][10] ), .A1(net112112), .B0(
        \i_MIPS/Register/register[14][10] ), .B1(net112142), .Y(n7327) );
  OA22XL U5896 ( .A0(\i_MIPS/Register/register[22][10] ), .A1(net112112), .B0(
        \i_MIPS/Register/register[30][10] ), .B1(net112142), .Y(n7336) );
  NAND3BX4 U5897 ( .AN(n8090), .B(n8088), .C(n8089), .Y(net98728) );
  AOI211X2 U5898 ( .A0(n9157), .A1(n9327), .B0(n9156), .C0(n9453), .Y(n9176)
         );
  INVX2 U5899 ( .A(n9151), .Y(n9157) );
  AO21X4 U5900 ( .A0(n6816), .A1(n6815), .B0(n3697), .Y(net98781) );
  BUFX20 U5901 ( .A(n5088), .Y(n5085) );
  AOI222X2 U5902 ( .A0(n5500), .A1(n11415), .B0(mem_rdata_D[65]), .B1(n236), 
        .C0(n12986), .C1(n4385), .Y(n10909) );
  NOR2BX4 U5903 ( .AN(\i_MIPS/IR_ID[23] ), .B(\i_MIPS/n234 ), .Y(n4499) );
  OA22X1 U5904 ( .A0(n5103), .A1(n1228), .B0(n5055), .B1(n2765), .Y(n6071) );
  NAND2BX4 U5905 ( .AN(n10387), .B(n10386), .Y(n10388) );
  AOI2BB1X4 U5906 ( .A0N(n10420), .A1N(n10385), .B0(n10384), .Y(n10387) );
  INVX2 U5907 ( .A(n10800), .Y(n10806) );
  NAND4X2 U5908 ( .A(n9923), .B(n9922), .C(n9921), .D(n9920), .Y(n11191) );
  OR2X2 U5909 ( .A(n8917), .B(net111622), .Y(n4176) );
  NAND4BX2 U5910 ( .AN(n7379), .B(n7378), .C(n7377), .D(n7376), .Y(net104109)
         );
  BUFX20 U5911 ( .A(n4728), .Y(n4731) );
  AOI222X2 U5912 ( .A0(n4422), .A1(net103710), .B0(n6975), .B1(n6974), .C0(
        n6973), .C1(n6972), .Y(n6983) );
  NAND2X4 U5913 ( .A(n4447), .B(n4446), .Y(net102048) );
  OA22X2 U5914 ( .A0(n4669), .A1(n7149), .B0(net112332), .B1(\i_MIPS/n344 ), 
        .Y(n7150) );
  AOI22X2 U5915 ( .A0(net108664), .A1(n10354), .B0(\i_MIPS/IF_ID[93] ), .B1(
        n3930), .Y(n4377) );
  NAND3BX4 U5916 ( .AN(n8228), .B(n9273), .C(n8227), .Y(n8944) );
  INVX3 U5917 ( .A(n9142), .Y(n8227) );
  OA22X4 U5918 ( .A0(n9984), .A1(n4675), .B0(n10917), .B1(n4250), .Y(n8405) );
  CLKAND2X12 U5919 ( .A(n5551), .B(n11417), .Y(mem_wdata_D[67]) );
  NAND4X4 U5920 ( .A(n8395), .B(n8394), .C(n8393), .D(n8392), .Y(n11417) );
  OAI221X2 U5921 ( .A0(net112368), .A1(\i_MIPS/n360 ), .B0(net112350), .B1(
        \i_MIPS/n359 ), .C0(n6485), .Y(n8739) );
  OA22X4 U5922 ( .A0(n4669), .A1(\i_MIPS/n358 ), .B0(net112336), .B1(
        \i_MIPS/n357 ), .Y(n6485) );
  AOI2BB1X4 U5923 ( .A0N(n4474), .A1N(n10602), .B0(n10405), .Y(n10407) );
  NAND2BX4 U5924 ( .AN(n5427), .B(n11186), .Y(n9951) );
  OAI221X2 U5925 ( .A0(n8724), .A1(net111622), .B0(n8723), .B1(net111634), 
        .C0(n8722), .Y(n10694) );
  AOI21X2 U5926 ( .A0(n10326), .A1(n10634), .B0(n10253), .Y(n10254) );
  AO21X4 U5927 ( .A0(n7590), .A1(n7589), .B0(n5546), .Y(net98367) );
  BUFX6 U5928 ( .A(n4800), .Y(n4798) );
  OAI222X4 U5929 ( .A0(net133471), .A1(n8165), .B0(n8163), .B1(n9455), .C0(
        n8162), .C1(net112420), .Y(n8169) );
  NAND4X4 U5930 ( .A(n6095), .B(n6094), .C(n6093), .D(n6092), .Y(n6106) );
  NAND4X4 U5931 ( .A(n6031), .B(n6030), .C(n6029), .D(n6028), .Y(n6043) );
  OA22X4 U5932 ( .A0(n5376), .A1(n2163), .B0(n5355), .B1(n588), .Y(n9649) );
  OAI2BB1X4 U5933 ( .A0N(n10853), .A1N(n10792), .B0(n10852), .Y(n10794) );
  NAND2X2 U5934 ( .A(n4527), .B(n4661), .Y(n4335) );
  AO21X4 U5935 ( .A0(net98780), .A1(net98781), .B0(net111640), .Y(net105196)
         );
  OAI221X4 U5936 ( .A0(n9257), .A1(n9336), .B0(n9256), .B1(n9255), .C0(n9254), 
        .Y(n9258) );
  INVX2 U5937 ( .A(n9255), .Y(n9161) );
  NAND3BX4 U5938 ( .AN(n6858), .B(n6856), .C(n6857), .Y(net97770) );
  INVX6 U5939 ( .A(n6693), .Y(n6694) );
  XNOR2X4 U5940 ( .A(ICACHE_addr[15]), .B(n11330), .Y(n6028) );
  AOI211X2 U5941 ( .A0(n8461), .A1(n8460), .B0(n8458), .C0(n8459), .Y(n8462)
         );
  OAI221X4 U5942 ( .A0(\i_MIPS/ALUin1[19] ), .A1(n4668), .B0(
        \i_MIPS/ALUin1[20] ), .B1(n3828), .C0(n8252), .Y(n8439) );
  OA21X2 U5943 ( .A0(\i_MIPS/ALUin1[18] ), .A1(net112350), .B0(n8251), .Y(
        n8252) );
  NAND4X6 U5944 ( .A(n5986), .B(n5985), .C(n5984), .D(n5983), .Y(n11321) );
  AO21X2 U5945 ( .A0(n7688), .A1(n7693), .B0(n7525), .Y(n7524) );
  AOI211X2 U5946 ( .A0(n3718), .A1(n7712), .B0(n7711), .C0(n7710), .Y(n7713)
         );
  OAI221X2 U5947 ( .A0(n4668), .A1(\i_MIPS/n363 ), .B0(n3828), .B1(net103561), 
        .C0(n7697), .Y(n9160) );
  XNOR3X4 U5948 ( .A(net112400), .B(n10863), .C(n10856), .Y(n4326) );
  NAND2BX4 U5949 ( .AN(n5427), .B(n11195), .Y(n10037) );
  AO22X4 U5950 ( .A0(net111960), .A1(n7181), .B0(net111968), .B1(net98012), 
        .Y(net104495) );
  OA22X1 U5951 ( .A0(n10874), .A1(n4245), .B0(n10877), .B1(n4246), .Y(n6657)
         );
  AOI21X2 U5952 ( .A0(n9268), .A1(n9264), .B0(n7539), .Y(n6578) );
  BUFX4 U5953 ( .A(n4800), .Y(n4797) );
  AOI33X4 U5954 ( .A0(n8074), .A1(n8077), .A2(net137952), .B0(n8073), .B1(
        n8075), .B2(net137952), .Y(n8089) );
  AO22X4 U5955 ( .A0(n10855), .A1(net112404), .B0(n10853), .B1(n10854), .Y(
        n10856) );
  XOR2X4 U5956 ( .A(n10284), .B(ICACHE_addr[24]), .Y(n10828) );
  NAND2X4 U5957 ( .A(n10340), .B(net112404), .Y(n10574) );
  OAI2BB1X4 U5958 ( .A0N(n9514), .A1N(n9513), .B0(n3720), .Y(n10221) );
  BUFX20 U5959 ( .A(n4990), .Y(n4988) );
  MXI2X4 U5960 ( .A(n10696), .B(n10695), .S0(n5517), .Y(n10697) );
  AOI222X2 U5961 ( .A0(n5496), .A1(n11455), .B0(mem_rdata_D[105]), .B1(n234), 
        .C0(n12978), .C1(n5493), .Y(n10696) );
  NAND4BX4 U5962 ( .AN(n7988), .B(n7987), .C(n7986), .D(n7985), .Y(net97800)
         );
  OA22X4 U5963 ( .A0(n4834), .A1(n2164), .B0(n4879), .B1(n589), .Y(n6421) );
  BUFX20 U5964 ( .A(n9339), .Y(n4658) );
  AOI2BB1X2 U5965 ( .A0N(net133688), .A1N(n9047), .B0(n9453), .Y(n9048) );
  BUFX20 U5966 ( .A(n5353), .Y(n5331) );
  INVX20 U5967 ( .A(net108664), .Y(net108658) );
  NAND2BX4 U5968 ( .AN(n10341), .B(n10574), .Y(n10835) );
  MXI2X4 U5969 ( .A(n10885), .B(n10884), .S0(n5520), .Y(n10886) );
  NAND3BX2 U5970 ( .AN(n10415), .B(n10413), .C(n10414), .Y(\i_MIPS/PC/n48 ) );
  OAI221X2 U5971 ( .A0(\i_MIPS/PHT_2/n8 ), .A1(n11065), .B0(\i_MIPS/PHT_2/n8 ), 
        .B1(n11064), .C0(n11063), .Y(n11508) );
  AO21X4 U5972 ( .A0(n10559), .A1(n10558), .B0(net111902), .Y(net98500) );
  BUFX20 U5973 ( .A(n4796), .Y(n4789) );
  OAI221X2 U5974 ( .A0(\i_MIPS/PHT_2/n4 ), .A1(n11060), .B0(\i_MIPS/PHT_2/n4 ), 
        .B1(n11064), .C0(n11059), .Y(n11509) );
  NAND2X4 U5975 ( .A(n11108), .B(n11106), .Y(n11089) );
  NAND4X4 U5976 ( .A(n9949), .B(n9948), .C(n9947), .D(n9946), .Y(n11106) );
  AOI222X4 U5977 ( .A0(n3718), .A1(n4459), .B0(net101908), .B1(n8655), .C0(
        net101910), .C1(n9055), .Y(n8660) );
  NAND2X4 U5978 ( .A(n7218), .B(n7891), .Y(n8634) );
  OAI2BB1X4 U5979 ( .A0N(n7878), .A1N(n7877), .B0(n7876), .Y(n7882) );
  CLKAND2X8 U5980 ( .A(n11064), .B(net112691), .Y(n4434) );
  NAND2X2 U5981 ( .A(n10505), .B(n4571), .Y(n10325) );
  AO21X4 U5982 ( .A0(n8314), .A1(n8313), .B0(n3697), .Y(n10566) );
  XOR2X4 U5983 ( .A(n8430), .B(n8429), .Y(n8529) );
  AO21X4 U5984 ( .A0(n9978), .A1(n9977), .B0(net111640), .Y(n8426) );
  CLKAND2X6 U5985 ( .A(\i_MIPS/ALUin1[26] ), .B(net112370), .Y(n4513) );
  INVX12 U5986 ( .A(n4671), .Y(n4668) );
  AOI2BB1X4 U5987 ( .A0N(net112350), .A1N(\i_MIPS/n346 ), .B0(n4513), .Y(n7148) );
  BUFX20 U5988 ( .A(n15), .Y(net108682) );
  NOR2BX4 U5989 ( .AN(\i_MIPS/IR_ID[18] ), .B(\i_MIPS/n318 ), .Y(n4501) );
  OAI211X2 U5990 ( .A0(n8082), .A1(n8083), .B0(n8081), .C0(n8080), .Y(n8087)
         );
  AO22X4 U5991 ( .A0(n4073), .A1(n10346), .B0(net112406), .B1(
        \i_MIPS/IR_ID[30] ), .Y(\i_MIPS/N88 ) );
  OA22X4 U5992 ( .A0(n10741), .A1(n4676), .B0(n10744), .B1(n4250), .Y(n7662)
         );
  BUFX20 U5993 ( .A(n3424), .Y(n4676) );
  NAND3BX2 U5994 ( .AN(n10608), .B(n10606), .C(n10607), .Y(\i_MIPS/PC/n47 ) );
  AO21X4 U5995 ( .A0(n8167), .A1(net103354), .B0(n7821), .Y(n7967) );
  AO21X4 U5996 ( .A0(n7948), .A1(n7947), .B0(n3729), .Y(net98336) );
  OA22X4 U5997 ( .A0(n10887), .A1(n4245), .B0(n10890), .B1(n4246), .Y(n7947)
         );
  XNOR2X2 U5998 ( .A(ICACHE_addr[13]), .B(n11328), .Y(n6061) );
  AO22X4 U5999 ( .A0(n5537), .A1(ICACHE_addr[25]), .B0(n239), .B1(n11340), .Y(
        n11146) );
  AND2X4 U6000 ( .A(\i_MIPS/ALUin1[26] ), .B(net127710), .Y(n4510) );
  NAND4X4 U6001 ( .A(n7424), .B(n7423), .C(n7422), .D(n7421), .Y(net98063) );
  AOI2BB1X4 U6002 ( .A0N(n4465), .A1N(n4386), .B0(n10610), .Y(n10612) );
  NAND4X2 U6003 ( .A(n6091), .B(n6090), .C(n6089), .D(n6088), .Y(n11344) );
  XNOR2X1 U6004 ( .A(ICACHE_addr[5]), .B(n11320), .Y(n6104) );
  NAND4BX4 U6005 ( .AN(n4339), .B(n6098), .C(n6097), .D(n6096), .Y(n11320) );
  XOR2X4 U6006 ( .A(n9549), .B(n3896), .Y(n9550) );
  NAND2X2 U6007 ( .A(n9161), .B(n8866), .Y(n8867) );
  NAND3BX2 U6008 ( .AN(n11084), .B(n11083), .C(n11082), .Y(\i_MIPS/PC/n37 ) );
  OAI221X4 U6009 ( .A0(n4668), .A1(\i_MIPS/n361 ), .B0(n3828), .B1(
        \i_MIPS/n360 ), .C0(n6684), .Y(n8866) );
  NAND4X2 U6010 ( .A(n6051), .B(n6050), .C(n6049), .D(n6048), .Y(n11329) );
  NAND2BX2 U6011 ( .AN(n5428), .B(n11198), .Y(n9781) );
  OR2X8 U6012 ( .A(n10335), .B(n10539), .Y(n10445) );
  OAI222X4 U6013 ( .A0(n8069), .A1(n4659), .B0(n4660), .B1(n9252), .C0(n4536), 
        .C1(n9251), .Y(n8455) );
  OA22X2 U6014 ( .A0(net133471), .A1(n3688), .B0(n8455), .B1(n7901), .Y(n7423)
         );
  AO21X4 U6015 ( .A0(n9303), .A1(n9302), .B0(n5546), .Y(n10564) );
  OAI221X2 U6016 ( .A0(n7243), .A1(n7242), .B0(n7241), .B1(n7240), .C0(n7239), 
        .Y(net98080) );
  AO22X1 U6017 ( .A0(n4073), .A1(n10347), .B0(net112406), .B1(
        \i_MIPS/IR_ID[28] ), .Y(\i_MIPS/N86 ) );
  XNOR2X4 U6018 ( .A(n4324), .B(n262), .Y(n8528) );
  AO21X4 U6019 ( .A0(n9066), .A1(n9065), .B0(n9064), .Y(n9068) );
  INVX3 U6020 ( .A(n9483), .Y(n9146) );
  OA22X2 U6021 ( .A0(n5385), .A1(n701), .B0(n5352), .B1(n2270), .Y(n9654) );
  XOR2X4 U6022 ( .A(n10345), .B(net112400), .Y(n10354) );
  NAND4X4 U6023 ( .A(n3781), .B(ICACHE_addr[8]), .C(n4469), .D(n10224), .Y(
        n10232) );
  NAND2X2 U6024 ( .A(n4462), .B(n10084), .Y(n10998) );
  OA22X4 U6025 ( .A0(n4924), .A1(n2165), .B0(n4955), .B1(n591), .Y(n6398) );
  NAND3BX2 U6026 ( .AN(n10649), .B(n10648), .C(n10647), .Y(\i_MIPS/PC/n53 ) );
  AOI211X2 U6027 ( .A0(n6981), .A1(net101908), .B0(n6980), .C0(n6979), .Y(
        n6982) );
  NAND2BX4 U6028 ( .AN(n10244), .B(n10247), .Y(n10383) );
  NAND2BX4 U6029 ( .AN(n10436), .B(n10435), .Y(n10621) );
  OAI32X2 U6030 ( .A0(n10362), .A1(n10361), .A2(n10205), .B0(n10204), .B1(
        n10205), .Y(n10206) );
  NAND2BX4 U6031 ( .AN(n11185), .B(n11314), .Y(n11317) );
  INVX6 U6032 ( .A(n11317), .Y(n11513) );
  NAND4X2 U6033 ( .A(n6083), .B(n6082), .C(n6081), .D(n6080), .Y(n11331) );
  OA22X4 U6034 ( .A0(n8457), .A1(net100581), .B0(n7616), .B1(n9455), .Y(n6487)
         );
  INVX4 U6035 ( .A(n6446), .Y(n6608) );
  INVX20 U6036 ( .A(net111910), .Y(net111902) );
  XNOR2X4 U6037 ( .A(ICACHE_addr[12]), .B(n11327), .Y(n6063) );
  OR2X1 U6038 ( .A(n4986), .B(n2951), .Y(n4159) );
  OAI211X2 U6039 ( .A0(n8353), .A1(n8352), .B0(n8351), .C0(n8350), .Y(n8551)
         );
  OR2X1 U6040 ( .A(net112366), .B(\i_MIPS/n349 ), .Y(n4166) );
  AOI222X2 U6041 ( .A0(n8647), .A1(net100585), .B0(n8646), .B1(n8645), .C0(
        n8644), .C1(n8643), .Y(n8662) );
  NAND3BX4 U6042 ( .AN(n7067), .B(n7066), .C(n7065), .Y(net97817) );
  OA22X2 U6043 ( .A0(n9463), .A1(n7968), .B0(n8658), .B1(n9469), .Y(n7816) );
  NOR2X2 U6044 ( .A(n4172), .B(n7520), .Y(n4441) );
  NOR2XL U6045 ( .A(net133471), .B(n7876), .Y(n4174) );
  NOR2X1 U6046 ( .A(net103060), .B(net104885), .Y(n4175) );
  NAND2X8 U6047 ( .A(n4395), .B(net133411), .Y(net133471) );
  NAND2X6 U6048 ( .A(\i_MIPS/ALUin1[6] ), .B(n6536), .Y(n7876) );
  BUFX16 U6049 ( .A(n4766), .Y(n4762) );
  NAND2X8 U6050 ( .A(net112764), .B(n5624), .Y(n4180) );
  NAND2X8 U6051 ( .A(n4180), .B(n4181), .Y(n4182) );
  CLKINVX12 U6052 ( .A(n4182), .Y(n4616) );
  NAND2X6 U6053 ( .A(n4616), .B(\i_MIPS/n364 ), .Y(n7881) );
  NAND3X6 U6054 ( .A(n4187), .B(n4188), .C(n4189), .Y(n11176) );
  NAND2X2 U6055 ( .A(n10878), .B(n4190), .Y(n4191) );
  NAND2X2 U6056 ( .A(n10877), .B(n5520), .Y(n4192) );
  NAND2X6 U6057 ( .A(n4191), .B(n4192), .Y(n4193) );
  CLKINVX1 U6058 ( .A(n5520), .Y(n4190) );
  INVX12 U6059 ( .A(n4193), .Y(n10879) );
  INVX4 U6060 ( .A(n11413), .Y(n10877) );
  INVX4 U6061 ( .A(n11412), .Y(n10148) );
  INVX3 U6062 ( .A(n11411), .Y(n10690) );
  CLKMX2X3 U6063 ( .A(\D_cache/cache[0][93] ), .B(n3329), .S0(n4738), .Y(
        \D_cache/n1052 ) );
  MX2X2 U6064 ( .A(\D_cache/cache[1][93] ), .B(n3329), .S0(n4785), .Y(
        \D_cache/n1051 ) );
  MX2X2 U6065 ( .A(\D_cache/cache[2][93] ), .B(n3329), .S0(n4806), .Y(
        \D_cache/n1050 ) );
  MX2X2 U6066 ( .A(\D_cache/cache[3][93] ), .B(n3329), .S0(n4850), .Y(
        \D_cache/n1049 ) );
  MX2X2 U6067 ( .A(\D_cache/cache[4][93] ), .B(n3329), .S0(n4896), .Y(
        \D_cache/n1048 ) );
  MX2X2 U6068 ( .A(\D_cache/cache[5][93] ), .B(n3329), .S0(n4941), .Y(
        \D_cache/n1047 ) );
  MX2X2 U6069 ( .A(\D_cache/cache[6][93] ), .B(n3329), .S0(n4960), .Y(
        \D_cache/n1046 ) );
  MX2X2 U6070 ( .A(\D_cache/cache[7][93] ), .B(n3329), .S0(n5004), .Y(
        \D_cache/n1045 ) );
  CLKINVX1 U6071 ( .A(n5516), .Y(n4198) );
  CLKINVX1 U6072 ( .A(n5516), .Y(n4201) );
  CLKINVX1 U6073 ( .A(n5519), .Y(n4204) );
  INVX4 U6074 ( .A(n11399), .Y(n10772) );
  CLKINVX1 U6075 ( .A(n5519), .Y(n4207) );
  INVX4 U6076 ( .A(n11397), .Y(n10761) );
  OA21X4 U6077 ( .A0(n8431), .A1(n6528), .B0(n6527), .Y(n4216) );
  NAND2XL U6078 ( .A(n8166), .B(n6526), .Y(n6528) );
  OA21X4 U6079 ( .A0(n10247), .A1(n10419), .B0(n10418), .Y(n4217) );
  NAND2BX4 U6080 ( .AN(n10400), .B(n4389), .Y(n10419) );
  OA22XL U6081 ( .A0(n5293), .A1(n1580), .B0(n5260), .B1(n3162), .Y(n10188) );
  CLKAND2X12 U6082 ( .A(n5557), .B(n11189), .Y(mem_wdata_I[3]) );
  CLKAND2X2 U6083 ( .A(n10372), .B(n4453), .Y(n4218) );
  AO21X4 U6084 ( .A0(n10353), .A1(n10352), .B0(net98630), .Y(n10372) );
  XOR2X4 U6085 ( .A(n10545), .B(n10549), .Y(n10546) );
  AND2X1 U6086 ( .A(n11041), .B(n4453), .Y(n4223) );
  INVX1 U6087 ( .A(n10372), .Y(n11041) );
  OR2X1 U6088 ( .A(n9470), .B(n9469), .Y(n4224) );
  INVXL U6089 ( .A(n9464), .Y(n9470) );
  MX2XL U6090 ( .A(net100573), .B(net112438), .S0(n9465), .Y(n9466) );
  NAND3X6 U6091 ( .A(n8764), .B(n8761), .C(n4227), .Y(n10502) );
  INVX3 U6092 ( .A(n4226), .Y(n4227) );
  BUFX16 U6093 ( .A(n12938), .Y(DCACHE_addr[19]) );
  CLKINVX1 U6094 ( .A(n5520), .Y(n4232) );
  BUFX4 U6095 ( .A(n5524), .Y(n5520) );
  CLKINVX1 U6096 ( .A(n5516), .Y(n4237) );
  BUFX4 U6097 ( .A(n5525), .Y(n5516) );
  INVX4 U6098 ( .A(n11393), .Y(n10716) );
  BUFX8 U6099 ( .A(n10904), .Y(n4244) );
  OAI221X4 U6100 ( .A0(net112366), .A1(\i_MIPS/n370 ), .B0(net112348), .B1(
        \i_MIPS/n369 ), .C0(n6849), .Y(n7059) );
  XOR3X2 U6101 ( .A(net112400), .B(n10826), .C(n10828), .Y(n10830) );
  XOR3X2 U6102 ( .A(n10408), .B(n10407), .C(n10406), .Y(n10411) );
  NOR2X2 U6103 ( .A(n7163), .B(n7164), .Y(n7162) );
  OA22X4 U6104 ( .A0(n10067), .A1(n4676), .B0(n10073), .B1(n4250), .Y(n7021)
         );
  AOI211X2 U6105 ( .A0(n9328), .A1(n8249), .B0(n8087), .C0(n8086), .Y(n8088)
         );
  CLKINVX4 U6106 ( .A(n10395), .Y(n10393) );
  XOR3X2 U6107 ( .A(n409), .B(n10392), .C(n10394), .Y(n10395) );
  MX2X6 U6108 ( .A(n9252), .B(n7059), .S0(net107796), .Y(n8249) );
  OAI221X4 U6109 ( .A0(n4668), .A1(\i_MIPS/n364 ), .B0(n3828), .B1(
        \i_MIPS/n363 ), .C0(n7058), .Y(n9252) );
  NAND2XL U6110 ( .A(n8631), .B(n8630), .Y(n8646) );
  INVX1 U6111 ( .A(n8631), .Y(n7494) );
  BUFX8 U6112 ( .A(n4884), .Y(n4879) );
  AND3X2 U6113 ( .A(n7811), .B(n7820), .C(net111994), .Y(n7831) );
  INVX3 U6114 ( .A(n7811), .Y(n7801) );
  NAND3BX4 U6115 ( .AN(n9073), .B(n9072), .C(n9071), .Y(n10487) );
  OAI221X4 U6116 ( .A0(net112366), .A1(\i_MIPS/n359 ), .B0(net112350), .B1(
        \i_MIPS/n358 ), .C0(n6687), .Y(n8864) );
  AOI211X4 U6117 ( .A0(n3838), .A1(n8959), .B0(n7319), .C0(n7318), .Y(n7320)
         );
  OAI2BB1X4 U6118 ( .A0N(net103891), .A1N(n8339), .B0(n8338), .Y(n7504) );
  NAND2X1 U6119 ( .A(n8339), .B(n8338), .Y(n8345) );
  OAI211X2 U6120 ( .A0(n6706), .A1(net101257), .B0(n3907), .C0(net112420), .Y(
        n6597) );
  AO21X4 U6121 ( .A0(n9245), .A1(n8349), .B0(n4449), .Y(n8443) );
  INVX4 U6122 ( .A(n4587), .Y(n9245) );
  OA22X4 U6123 ( .A0(n10079), .A1(n4245), .B0(n10086), .B1(n4246), .Y(n7020)
         );
  AO21X4 U6124 ( .A0(n9197), .A1(n9196), .B0(n3665), .Y(n10562) );
  OAI2BB1X2 U6125 ( .A0N(n6841), .A1N(n7509), .B0(n7503), .Y(n6758) );
  OA22X4 U6126 ( .A0(n4911), .A1(n2089), .B0(n4946), .B1(n502), .Y(n8889) );
  OA22X4 U6127 ( .A0(n4911), .A1(n2090), .B0(n4947), .B1(n503), .Y(n8882) );
  OA22X4 U6128 ( .A0(n4911), .A1(n2071), .B0(n4946), .B1(n486), .Y(n8799) );
  OAI221X2 U6129 ( .A0(n8756), .A1(n8755), .B0(n8754), .B1(n8753), .C0(n8752), 
        .Y(n8758) );
  AND2X4 U6130 ( .A(\i_MIPS/ALUin1[27] ), .B(net112356), .Y(n4511) );
  NAND3BX4 U6131 ( .AN(n7322), .B(n7321), .C(n7320), .Y(net98393) );
  NAND4X4 U6132 ( .A(n9933), .B(n9932), .C(n9931), .D(n9930), .Y(n10800) );
  XNOR2X4 U6133 ( .A(n10546), .B(net112404), .Y(n10551) );
  AOI21X4 U6134 ( .A0(n4303), .A1(n4460), .B0(n10083), .Y(n4462) );
  INVX8 U6135 ( .A(n11051), .Y(n11064) );
  OA21X4 U6136 ( .A0(n4670), .A1(\i_MIPS/n359 ), .B0(n7698), .Y(n7699) );
  OA22X4 U6137 ( .A0(n4921), .A1(n2075), .B0(n4949), .B1(n487), .Y(n7195) );
  OA22X2 U6138 ( .A0(n4920), .A1(n739), .B0(n4949), .B1(n2300), .Y(n7434) );
  OA22X4 U6139 ( .A0(n4921), .A1(n2167), .B0(n4949), .B1(n593), .Y(n7187) );
  OAI33X2 U6140 ( .A0(n8954), .A1(n2209), .A2(net112300), .B0(n3698), .B1(
        n2209), .B2(net101257), .Y(n8974) );
  AO21X4 U6141 ( .A0(n11112), .A1(n11110), .B0(n11107), .Y(n11088) );
  OAI221X4 U6142 ( .A0(n4668), .A1(\i_MIPS/n366 ), .B0(n3828), .B1(n7696), 
        .C0(n6484), .Y(n7314) );
  AOI2BB1X4 U6143 ( .A0N(n4297), .A1N(n10624), .B0(n10623), .Y(n10625) );
  AO21X4 U6144 ( .A0(n7281), .A1(n7280), .B0(n3665), .Y(net98777) );
  AO21X4 U6145 ( .A0(n8108), .A1(n8109), .B0(n3665), .Y(n10286) );
  AO21X4 U6146 ( .A0(n7662), .A1(n7661), .B0(n5546), .Y(n10520) );
  AO21X4 U6147 ( .A0(net112338), .A1(\i_MIPS/ALUin1[29] ), .B0(n4518), .Y(
        n6772) );
  NOR2BX2 U6148 ( .AN(n4672), .B(\i_MIPS/n341 ), .Y(n4518) );
  AO21X4 U6149 ( .A0(n8803), .A1(n8802), .B0(n3665), .Y(n10503) );
  AO21X4 U6150 ( .A0(n8701), .A1(n8700), .B0(n3665), .Y(n10560) );
  AO21X4 U6151 ( .A0(n8504), .A1(n8503), .B0(n3665), .Y(n10321) );
  AO21X4 U6152 ( .A0(n9093), .A1(n9092), .B0(n3665), .Y(n10488) );
  NAND3BX4 U6153 ( .AN(n8078), .B(n8077), .C(net112294), .Y(n8081) );
  NAND2X2 U6154 ( .A(net112294), .B(n8181), .Y(n8176) );
  NAND2X2 U6155 ( .A(\i_MIPS/ALUin1[21] ), .B(n6571), .Y(n9137) );
  AOI222X2 U6156 ( .A0(n7615), .A1(n4587), .B0(n7417), .B1(n7416), .C0(n7415), 
        .C1(n7414), .Y(n7424) );
  OAI2BB1X4 U6157 ( .A0N(n6579), .A1N(n9265), .B0(n6578), .Y(n9144) );
  OA21X2 U6158 ( .A0(\i_MIPS/ALUin1[13] ), .A1(net112350), .B0(n7824), .Y(
        n7229) );
  OAI221X4 U6159 ( .A0(\i_MIPS/ALUin1[13] ), .A1(n4668), .B0(
        \i_MIPS/ALUin1[12] ), .B1(n3828), .C0(n6852), .Y(n7061) );
  AOI2BB2X2 U6160 ( .B0(\i_MIPS/IF_ID[69] ), .B1(net108670), .A0N(net108678), 
        .A1N(\i_MIPS/n187 ), .Y(n11114) );
  AOI2BB2X2 U6161 ( .B0(\i_MIPS/IF_ID[74] ), .B1(net108670), .A0N(net108676), 
        .A1N(\i_MIPS/n192 ), .Y(n10589) );
  NAND3BX2 U6162 ( .AN(n11129), .B(n11128), .C(n11127), .Y(\i_MIPS/PC/n55 ) );
  OAI222X4 U6163 ( .A0(n9342), .A1(n9047), .B0(n8176), .B1(n8432), .C0(n8167), 
        .C1(n8457), .Y(n8168) );
  NAND4X4 U6164 ( .A(n9909), .B(n9908), .C(n9907), .D(n9906), .Y(n11092) );
  CLKMX2X2 U6165 ( .A(\D_cache/cache[7][139] ), .B(n11016), .S0(n5006), .Y(
        \D_cache/n677 ) );
  CLKMX2X2 U6166 ( .A(\D_cache/cache[6][139] ), .B(n11016), .S0(n4962), .Y(
        \D_cache/n678 ) );
  CLKMX2X2 U6167 ( .A(\D_cache/cache[5][139] ), .B(n11016), .S0(n4941), .Y(
        \D_cache/n679 ) );
  CLKMX2X2 U6168 ( .A(\D_cache/cache[4][139] ), .B(n11016), .S0(n4898), .Y(
        \D_cache/n680 ) );
  CLKMX2X2 U6169 ( .A(\D_cache/cache[3][139] ), .B(n11016), .S0(n4852), .Y(
        \D_cache/n681 ) );
  CLKMX2X2 U6170 ( .A(\D_cache/cache[2][139] ), .B(n11016), .S0(n4802), .Y(
        \D_cache/n682 ) );
  AO22X2 U6171 ( .A0(n5528), .A1(n12943), .B0(n5526), .B1(n11492), .Y(n11025)
         );
  AO22X2 U6172 ( .A0(n5528), .A1(n12936), .B0(n5526), .B1(n11499), .Y(n11013)
         );
  CLKAND2X12 U6173 ( .A(n3783), .B(n11318), .Y(mem_addr_I[4]) );
  CLKAND2X12 U6174 ( .A(n4656), .B(n11296), .Y(mem_wdata_I[110]) );
  CLKAND2X12 U6175 ( .A(mem_write_I), .B(n11294), .Y(mem_wdata_I[108]) );
  CLKAND2X12 U6176 ( .A(n5557), .B(n11227), .Y(mem_wdata_I[41]) );
  INVX12 U6177 ( .A(\i_MIPS/n310 ), .Y(DCACHE_wen) );
  INVXL U6178 ( .A(n12988), .Y(n9557) );
  INVX12 U6179 ( .A(\i_MIPS/n246 ), .Y(DCACHE_wdata[31]) );
  INVX12 U6180 ( .A(\i_MIPS/n248 ), .Y(DCACHE_wdata[30]) );
  INVX12 U6181 ( .A(\i_MIPS/n250 ), .Y(DCACHE_wdata[29]) );
  INVX12 U6182 ( .A(\i_MIPS/n254 ), .Y(DCACHE_wdata[27]) );
  INVX12 U6183 ( .A(\i_MIPS/n258 ), .Y(DCACHE_wdata[25]) );
  INVX12 U6184 ( .A(\i_MIPS/n260 ), .Y(DCACHE_wdata[24]) );
  INVX12 U6185 ( .A(\i_MIPS/n262 ), .Y(DCACHE_wdata[23]) );
  INVX12 U6186 ( .A(\i_MIPS/n264 ), .Y(DCACHE_wdata[22]) );
  INVX12 U6187 ( .A(\i_MIPS/n266 ), .Y(DCACHE_wdata[21]) );
  INVX12 U6188 ( .A(\i_MIPS/n268 ), .Y(DCACHE_wdata[20]) );
  INVX12 U6189 ( .A(\i_MIPS/n272 ), .Y(DCACHE_wdata[18]) );
  INVX12 U6190 ( .A(\i_MIPS/n274 ), .Y(DCACHE_wdata[17]) );
  INVX12 U6191 ( .A(\i_MIPS/n276 ), .Y(DCACHE_wdata[16]) );
  INVX12 U6192 ( .A(\i_MIPS/n278 ), .Y(DCACHE_wdata[15]) );
  INVX12 U6193 ( .A(\i_MIPS/n280 ), .Y(DCACHE_wdata[14]) );
  INVX12 U6194 ( .A(\i_MIPS/n282 ), .Y(DCACHE_wdata[13]) );
  INVX12 U6195 ( .A(\i_MIPS/n284 ), .Y(DCACHE_wdata[12]) );
  INVX12 U6196 ( .A(\i_MIPS/n286 ), .Y(DCACHE_wdata[11]) );
  INVX12 U6197 ( .A(\i_MIPS/n288 ), .Y(DCACHE_wdata[10]) );
  INVX12 U6198 ( .A(\i_MIPS/n290 ), .Y(DCACHE_wdata[9]) );
  INVX12 U6199 ( .A(\i_MIPS/n292 ), .Y(DCACHE_wdata[8]) );
  INVX12 U6200 ( .A(\i_MIPS/n294 ), .Y(DCACHE_wdata[7]) );
  INVX12 U6201 ( .A(\i_MIPS/n296 ), .Y(DCACHE_wdata[6]) );
  INVX12 U6202 ( .A(\i_MIPS/n298 ), .Y(DCACHE_wdata[5]) );
  INVX12 U6203 ( .A(\i_MIPS/n300 ), .Y(DCACHE_wdata[4]) );
  INVX12 U6204 ( .A(\i_MIPS/n302 ), .Y(DCACHE_wdata[3]) );
  INVX12 U6205 ( .A(\i_MIPS/n306 ), .Y(DCACHE_wdata[1]) );
  INVX12 U6206 ( .A(\i_MIPS/n308 ), .Y(DCACHE_wdata[0]) );
  INVX12 U6207 ( .A(\i_MIPS/n252 ), .Y(DCACHE_wdata[28]) );
  INVX12 U6208 ( .A(\i_MIPS/n256 ), .Y(DCACHE_wdata[26]) );
  INVX12 U6209 ( .A(\i_MIPS/n304 ), .Y(DCACHE_wdata[2]) );
  INVX12 U6210 ( .A(\i_MIPS/n270 ), .Y(DCACHE_wdata[19]) );
  BUFX12 U6211 ( .A(n12943), .Y(DCACHE_addr[14]) );
  INVX12 U6212 ( .A(n4289), .Y(DCACHE_addr[5]) );
  INVX12 U6213 ( .A(n4291), .Y(DCACHE_addr[26]) );
  INVX12 U6214 ( .A(n4293), .Y(DCACHE_addr[24]) );
  AND2XL U6215 ( .A(net112400), .B(n10439), .Y(n4297) );
  AOI221X4 U6216 ( .A0(net137684), .A1(n4299), .B0(\i_MIPS/n309 ), .B1(n5625), 
        .C0(\i_MIPS/ALUin1[0] ), .Y(n4298) );
  AO22X4 U6217 ( .A0(n7307), .A1(net137952), .B0(net112296), .B1(n7306), .Y(
        n7310) );
  AO22X4 U6218 ( .A0(n7879), .A1(net111994), .B0(net112296), .B1(n7882), .Y(
        n7886) );
  AOI2BB2X4 U6219 ( .B0(n4456), .B1(n10177), .A0N(n11081), .A1N(n4302), .Y(
        n11107) );
  INVXL U6220 ( .A(n7313), .Y(n4305) );
  CLKBUFX2 U6221 ( .A(n5524), .Y(n5523) );
  BUFX8 U6222 ( .A(n4728), .Y(n4730) );
  BUFX8 U6223 ( .A(n4714), .Y(n4715) );
  BUFX4 U6224 ( .A(n5180), .Y(n5177) );
  INVX4 U6225 ( .A(n4477), .Y(n4697) );
  BUFX2 U6226 ( .A(n4844), .Y(n4842) );
  CLKBUFX3 U6227 ( .A(n5223), .Y(n5221) );
  CLKBUFX2 U6228 ( .A(n4998), .Y(n4996) );
  BUFX4 U6229 ( .A(n9524), .Y(n4677) );
  AO21X4 U6230 ( .A0(n10504), .A1(n10503), .B0(net111640), .Y(n8824) );
  OA22XL U6231 ( .A0(n5397), .A1(n1581), .B0(n5339), .B1(n3275), .Y(n9694) );
  OA22XL U6232 ( .A0(n5204), .A1(n1582), .B0(n5160), .B1(n3276), .Y(n9696) );
  OA22XL U6233 ( .A0(n5113), .A1(n1583), .B0(n5080), .B1(n3163), .Y(n9697) );
  OA22X1 U6234 ( .A0(n4744), .A1(n2954), .B0(n4789), .B1(n1144), .Y(n8895) );
  OA22X1 U6235 ( .A0(n4817), .A1(n1084), .B0(n4863), .B1(n2678), .Y(n8894) );
  OA22X2 U6236 ( .A0(n4759), .A1(n779), .B0(n4796), .B1(n2341), .Y(n6931) );
  OA22X2 U6237 ( .A0(n4983), .A1(n780), .B0(n5029), .B1(n2342), .Y(n6928) );
  OA22X2 U6238 ( .A0(n4831), .A1(n781), .B0(n4876), .B1(n2343), .Y(n6930) );
  OA22XL U6239 ( .A0(n4759), .A1(n1294), .B0(n4796), .B1(n2825), .Y(n6939) );
  OAI211X2 U6240 ( .A0(n6514), .A1(n7404), .B0(n6513), .C0(n7694), .Y(n8533)
         );
  CLKMX2X4 U6241 ( .A(n8155), .B(n7825), .S0(net107798), .Y(n9051) );
  OR2X4 U6242 ( .A(n7049), .B(n7048), .Y(n4311) );
  AO22XL U6243 ( .A0(n4721), .A1(n892), .B0(n4719), .B1(n2590), .Y(n7118) );
  AO22XL U6244 ( .A0(n4721), .A1(n867), .B0(n4719), .B1(n2551), .Y(n7109) );
  AO22XL U6245 ( .A0(n4721), .A1(n868), .B0(n4719), .B1(n2552), .Y(n6909) );
  AO22XL U6246 ( .A0(n4721), .A1(n869), .B0(n4719), .B1(n2553), .Y(n6900) );
  AO22XL U6247 ( .A0(n4721), .A1(n893), .B0(n4719), .B1(n2591), .Y(n6828) );
  AO22XL U6248 ( .A0(n4721), .A1(n870), .B0(n4719), .B1(n2554), .Y(n6819) );
  AO22XL U6249 ( .A0(n4721), .A1(n420), .B0(n4719), .B1(n2010), .Y(n6615) );
  AND2X2 U6250 ( .A(net112962), .B(n437), .Y(n4460) );
  NAND2XL U6251 ( .A(DCACHE_addr[4]), .B(n4673), .Y(net99157) );
  OA22X2 U6252 ( .A0(n4910), .A1(n782), .B0(n4249), .B1(n2344), .Y(n6929) );
  OA22X2 U6253 ( .A0(n4915), .A1(n783), .B0(n4947), .B1(n2345), .Y(n8022) );
  OA22X2 U6254 ( .A0(n5371), .A1(n1477), .B0(n5344), .B1(n3051), .Y(n9958) );
  OA22XL U6255 ( .A0(n4908), .A1(n1295), .B0(n4249), .B1(n2826), .Y(n6937) );
  NAND3X2 U6256 ( .A(ICACHE_addr[26]), .B(ICACHE_addr[25]), .C(n10569), .Y(
        n10793) );
  OA22X1 U6257 ( .A0(n5290), .A1(n3059), .B0(n5243), .B1(n1145), .Y(n6218) );
  CLKMX2X2 U6258 ( .A(\I_cache/cache[4][74] ), .B(n10059), .S0(n5272), .Y(
        n12191) );
  OA22XL U6259 ( .A0(\i_MIPS/Register/register[20][18] ), .A1(n4697), .B0(
        \i_MIPS/Register/register[28][18] ), .B1(n4693), .Y(n8820) );
  AO22XL U6260 ( .A0(net112004), .A1(n339), .B0(net112030), .B1(n1054), .Y(
        n8052) );
  AO22XL U6261 ( .A0(net112004), .A1(n340), .B0(net112030), .B1(n1055), .Y(
        n8061) );
  AO22XL U6262 ( .A0(net112002), .A1(n894), .B0(net112020), .B1(n2592), .Y(
        n7639) );
  AO22XL U6263 ( .A0(net112002), .A1(n895), .B0(net112020), .B1(n2593), .Y(
        n7249) );
  AO22XL U6264 ( .A0(net112002), .A1(n896), .B0(net112020), .B1(n2594), .Y(
        n7258) );
  AO22XL U6265 ( .A0(net112002), .A1(n897), .B0(net112020), .B1(n2595), .Y(
        n7132) );
  AO22XL U6266 ( .A0(net112002), .A1(n898), .B0(net112020), .B1(n2596), .Y(
        n7141) );
  AO22XL U6267 ( .A0(net112004), .A1(n341), .B0(net112030), .B1(n1056), .Y(
        n7723) );
  AO22XL U6268 ( .A0(net112002), .A1(n899), .B0(net112020), .B1(n2597), .Y(
        n7557) );
  AO22XL U6269 ( .A0(net112002), .A1(n900), .B0(net112020), .B1(n2598), .Y(
        n7566) );
  AO22XL U6270 ( .A0(net112004), .A1(n356), .B0(net112032), .B1(n1064), .Y(
        n7732) );
  AO22XL U6271 ( .A0(net112004), .A1(n357), .B0(net112030), .B1(n1065), .Y(
        n7915) );
  AO22XL U6272 ( .A0(net112004), .A1(n358), .B0(net112030), .B1(n1066), .Y(
        n7924) );
  AO22XL U6273 ( .A0(net112004), .A1(n359), .B0(net112030), .B1(n1067), .Y(
        n7791) );
  OA22XL U6274 ( .A0(\i_MIPS/Register/register[16][18] ), .A1(n4702), .B0(
        \i_MIPS/Register/register[24][18] ), .B1(n4700), .Y(n8819) );
  OA22XL U6275 ( .A0(n5290), .A1(n3074), .B0(n5243), .B1(n1184), .Y(n6208) );
  MX2XL U6276 ( .A(\I_cache/cache[5][74] ), .B(n10059), .S0(n5229), .Y(n12190)
         );
  OA22X2 U6277 ( .A0(n5122), .A1(n1478), .B0(n5083), .B1(n3052), .Y(n10115) );
  CLKINVX16 U6278 ( .A(net111646), .Y(net111640) );
  NAND2X1 U6279 ( .A(net112962), .B(DCACHE_addr[1]), .Y(n10077) );
  OA22X2 U6280 ( .A0(n5292), .A1(n3030), .B0(n5258), .B1(n850), .Y(n10113) );
  AO22X4 U6281 ( .A0(\i_MIPS/ID_EX[42] ), .A1(n5625), .B0(n5624), .B1(n3812), 
        .Y(n6538) );
  CLKBUFX3 U6282 ( .A(n5263), .Y(n5250) );
  BUFX4 U6283 ( .A(n4685), .Y(n4686) );
  INVX3 U6284 ( .A(n10585), .Y(n10227) );
  AO22X4 U6285 ( .A0(net111966), .A1(net97703), .B0(net111960), .B1(n6798), 
        .Y(net105282) );
  OA22X2 U6286 ( .A0(n5401), .A1(n1479), .B0(n5344), .B1(n3053), .Y(n10112) );
  AND2X2 U6287 ( .A(n6638), .B(n6637), .Y(n4515) );
  BUFX2 U6288 ( .A(n4844), .Y(n4841) );
  AO21X4 U6289 ( .A0(n10489), .A1(n10488), .B0(net111640), .Y(n9114) );
  MX2X2 U6290 ( .A(n9050), .B(n8155), .S0(net107798), .Y(n9167) );
  BUFX2 U6291 ( .A(\i_MIPS/n336 ), .Y(n4673) );
  OA22XL U6292 ( .A0(n4915), .A1(n1146), .B0(n4947), .B1(n2705), .Y(n8097) );
  OA22XL U6293 ( .A0(n4915), .A1(n1296), .B0(n4947), .B1(n2827), .Y(n8105) );
  OA22XL U6294 ( .A0(\i_MIPS/Register/register[5][16] ), .A1(net112222), .B0(
        \i_MIPS/Register/register[13][16] ), .B1(net112240), .Y(n8049) );
  OA22XL U6295 ( .A0(\i_MIPS/Register/register[17][27] ), .A1(net112258), .B0(
        \i_MIPS/Register/register[25][27] ), .B1(n147), .Y(n9373) );
  OA22XL U6296 ( .A0(\i_MIPS/Register/register[19][27] ), .A1(net112188), .B0(
        \i_MIPS/Register/register[27][27] ), .B1(n197), .Y(n9371) );
  OA22XL U6297 ( .A0(\i_MIPS/Register/register[23][27] ), .A1(net112152), .B0(
        \i_MIPS/Register/register[31][27] ), .B1(net112172), .Y(n9370) );
  INVX3 U6298 ( .A(n5044), .Y(n5043) );
  CLKBUFX2 U6299 ( .A(n5223), .Y(n5222) );
  NAND2BX2 U6300 ( .AN(n5429), .B(n11222), .Y(n9906) );
  AO21X4 U6301 ( .A0(n8951), .A1(n8949), .B0(n7490), .Y(n9349) );
  NAND2BX2 U6302 ( .AN(n5425), .B(n11258), .Y(n10015) );
  INVXL U6303 ( .A(n9494), .Y(n9485) );
  OA22X2 U6304 ( .A0(n4746), .A1(n784), .B0(n4790), .B1(n2346), .Y(n8691) );
  OA22X1 U6305 ( .A0(n4753), .A1(n2955), .B0(n4792), .B1(n1147), .Y(n7746) );
  OA22XL U6306 ( .A0(n4825), .A1(n1297), .B0(n4870), .B1(n2828), .Y(n7745) );
  INVX3 U6307 ( .A(n10373), .Y(n10370) );
  AO22X1 U6308 ( .A0(net112036), .A1(n940), .B0(net100603), .B1(n2450), .Y(
        n6999) );
  OAI221XL U6309 ( .A0(\i_MIPS/Register/register[18][6] ), .A1(net112072), 
        .B0(\i_MIPS/Register/register[26][6] ), .B1(net112090), .C0(n6997), 
        .Y(n7000) );
  NAND2X1 U6310 ( .A(n4434), .B(n11065), .Y(n4529) );
  OA22X1 U6311 ( .A0(\i_MIPS/Register/register[5][8] ), .A1(n192), .B0(
        \i_MIPS/Register/register[13][8] ), .B1(net112236), .Y(n7070) );
  OA22X1 U6312 ( .A0(\i_MIPS/Register/register[16][16] ), .A1(n4703), .B0(
        \i_MIPS/Register/register[24][16] ), .B1(n4701), .Y(n8125) );
  AO22X1 U6313 ( .A0(n4728), .A1(n369), .B0(n4727), .B1(n1023), .Y(n8906) );
  NAND3BX4 U6314 ( .AN(n4664), .B(n6298), .C(n4663), .Y(n4333) );
  CLKBUFX2 U6315 ( .A(n5266), .Y(n5234) );
  BUFX2 U6316 ( .A(n5259), .Y(n5235) );
  BUFX8 U6317 ( .A(net128830), .Y(net111630) );
  BUFX8 U6318 ( .A(n5180), .Y(n5173) );
  CLKBUFX2 U6319 ( .A(n4844), .Y(n4843) );
  INVX3 U6320 ( .A(n8561), .Y(n8543) );
  AO22X4 U6321 ( .A0(net111960), .A1(n9179), .B0(net111966), .B1(n10665), .Y(
        n9180) );
  AO22XL U6322 ( .A0(n9531), .A1(n901), .B0(n4717), .B1(n2599), .Y(n7961) );
  AO22XL U6323 ( .A0(n9531), .A1(n902), .B0(n4717), .B1(n2600), .Y(n7952) );
  AO22XL U6324 ( .A0(n4712), .A1(n871), .B0(n4709), .B1(n2555), .Y(n8808) );
  AO22XL U6325 ( .A0(n4712), .A1(n276), .B0(n4709), .B1(n2601), .Y(n8715) );
  AO22XL U6326 ( .A0(n4712), .A1(n872), .B0(n4709), .B1(n2556), .Y(n8706) );
  OA22XL U6327 ( .A0(n5384), .A1(n3075), .B0(n5339), .B1(n1421), .Y(n9689) );
  OA22XL U6328 ( .A0(n5204), .A1(n1584), .B0(n5160), .B1(n3164), .Y(n9691) );
  OA22XL U6329 ( .A0(n5113), .A1(n1585), .B0(n5072), .B1(n3165), .Y(n9692) );
  OA22XL U6330 ( .A0(n4755), .A1(n2959), .B0(n4793), .B1(n1185), .Y(n7432) );
  OA22XL U6331 ( .A0(n4753), .A1(n1298), .B0(n4792), .B1(n2829), .Y(n7750) );
  OA22XL U6332 ( .A0(n4978), .A1(n1299), .B0(n5023), .B1(n2830), .Y(n7747) );
  OA22XL U6333 ( .A0(n5126), .A1(n1684), .B0(n5087), .B1(n3277), .Y(n10001) );
  AO22XL U6334 ( .A0(net128155), .A1(n423), .B0(net112232), .B1(n2002), .Y(
        n6470) );
  AO22XL U6335 ( .A0(net128155), .A1(n420), .B0(net112232), .B1(n2010), .Y(
        n6461) );
  AO22XL U6336 ( .A0(net128155), .A1(n416), .B0(net112232), .B1(n1977), .Y(
        n8569) );
  AO22XL U6337 ( .A0(net128155), .A1(n417), .B0(net112232), .B1(n2001), .Y(
        n8578) );
  AO22XL U6338 ( .A0(n9531), .A1(n903), .B0(n4714), .B1(n2602), .Y(n9538) );
  AO22XL U6339 ( .A0(n4713), .A1(n266), .B0(n4710), .B1(n2603), .Y(n9539) );
  AO22XL U6340 ( .A0(n9531), .A1(n904), .B0(n4714), .B1(n2604), .Y(n9518) );
  AO22XL U6341 ( .A0(n4713), .A1(n905), .B0(n4710), .B1(n2605), .Y(n9519) );
  AO22XL U6342 ( .A0(n9531), .A1(n906), .B0(n4717), .B1(n2606), .Y(n7867) );
  AO22XL U6343 ( .A0(n9531), .A1(n907), .B0(n4717), .B1(n2607), .Y(n7858) );
  AO22XL U6344 ( .A0(n4713), .A1(n908), .B0(n4708), .B1(n2608), .Y(n7859) );
  AO22XL U6345 ( .A0(n4713), .A1(n873), .B0(n4710), .B1(n2557), .Y(n8900) );
  AO22XL U6346 ( .A0(n9531), .A1(n909), .B0(n4717), .B1(n2609), .Y(n8217) );
  AO22XL U6347 ( .A0(n9531), .A1(n910), .B0(n4717), .B1(n2610), .Y(n8208) );
  AO22XL U6348 ( .A0(n4713), .A1(n911), .B0(n4708), .B1(n2611), .Y(n8209) );
  AO22XL U6349 ( .A0(n9531), .A1(n912), .B0(n4714), .B1(n2612), .Y(n9009) );
  AO22XL U6350 ( .A0(n4713), .A1(n267), .B0(n4710), .B1(n2613), .Y(n9010) );
  AO22XL U6351 ( .A0(n9531), .A1(n913), .B0(n4714), .B1(n2614), .Y(n9000) );
  AO22XL U6352 ( .A0(n4713), .A1(n914), .B0(n4710), .B1(n2615), .Y(n9001) );
  AO22XL U6353 ( .A0(n9531), .A1(n422), .B0(n4715), .B1(n2013), .Y(n6616) );
  AO22XL U6354 ( .A0(n9531), .A1(n421), .B0(n4715), .B1(n2012), .Y(n6625) );
  AO22XL U6355 ( .A0(n4711), .A1(n265), .B0(n4707), .B1(n2011), .Y(n6626) );
  AO22XL U6356 ( .A0(n4712), .A1(n268), .B0(n4709), .B1(n2616), .Y(n8419) );
  AO22XL U6357 ( .A0(n4712), .A1(n874), .B0(n4709), .B1(n2558), .Y(n8410) );
  AO22XL U6358 ( .A0(n4711), .A1(n309), .B0(n4707), .B1(n2617), .Y(n7120) );
  AO22XL U6359 ( .A0(n9531), .A1(n915), .B0(n4715), .B1(n2618), .Y(n7110) );
  AO22XL U6360 ( .A0(n4711), .A1(n916), .B0(n4707), .B1(n2619), .Y(n7111) );
  AO22XL U6361 ( .A0(n4712), .A1(n875), .B0(n4709), .B1(n2559), .Y(n8509) );
  AO22XL U6362 ( .A0(n4711), .A1(n271), .B0(n4709), .B1(n2560), .Y(n8328) );
  AO22XL U6363 ( .A0(n4712), .A1(n432), .B0(n4709), .B1(n2561), .Y(n8319) );
  AO22XL U6364 ( .A0(n4713), .A1(n278), .B0(n4709), .B1(n2620), .Y(n8518) );
  AO22XL U6365 ( .A0(n9531), .A1(n917), .B0(n4715), .B1(n2621), .Y(n6910) );
  AO22XL U6366 ( .A0(n4711), .A1(n310), .B0(n4707), .B1(n2622), .Y(n6911) );
  AO22XL U6367 ( .A0(n9531), .A1(n918), .B0(n4715), .B1(n2623), .Y(n6901) );
  AO22XL U6368 ( .A0(n4711), .A1(n876), .B0(n4707), .B1(n2562), .Y(n6902) );
  AO22XL U6369 ( .A0(n9531), .A1(n919), .B0(n4715), .B1(n2624), .Y(n6829) );
  AO22XL U6370 ( .A0(n4711), .A1(n277), .B0(n4707), .B1(n2625), .Y(n6830) );
  AO22XL U6371 ( .A0(n9531), .A1(n920), .B0(n4715), .B1(n2626), .Y(n6820) );
  AO22XL U6372 ( .A0(n4711), .A1(n877), .B0(n4707), .B1(n2563), .Y(n6821) );
  INVXL U6373 ( .A(n8439), .Y(n8255) );
  AO22XL U6374 ( .A0(n4730), .A1(n426), .B0(n4726), .B1(n2008), .Y(n6623) );
  AO22XL U6375 ( .A0(n4730), .A1(n427), .B0(n4726), .B1(n2009), .Y(n6614) );
  OA22XL U6376 ( .A0(\i_MIPS/Register/register[6][8] ), .A1(net112110), .B0(
        \i_MIPS/Register/register[14][8] ), .B1(net112128), .Y(n7072) );
  NAND3BX4 U6377 ( .AN(n9883), .B(n259), .C(n9885), .Y(n6445) );
  CLKMX2X2 U6378 ( .A(n3593), .B(n4611), .S0(n208), .Y(\i_MIPS/n429 ) );
  OA22XL U6379 ( .A0(\i_MIPS/Register/register[20][16] ), .A1(n4698), .B0(
        \i_MIPS/Register/register[28][16] ), .B1(n4694), .Y(n8126) );
  OA22XL U6380 ( .A0(n4912), .A1(n1300), .B0(n4249), .B1(n2980), .Y(n8689) );
  AO22XL U6381 ( .A0(n4729), .A1(n342), .B0(n4725), .B1(n1057), .Y(n8712) );
  AO22XL U6382 ( .A0(n4729), .A1(n343), .B0(n4725), .B1(n1058), .Y(n8703) );
  OA22XL U6383 ( .A0(n5293), .A1(n1586), .B0(n5246), .B1(n3166), .Y(n9601) );
  OA22XL U6384 ( .A0(\i_MIPS/Register/register[6][16] ), .A1(net112112), .B0(
        \i_MIPS/Register/register[14][16] ), .B1(net112132), .Y(n8051) );
  OA22XL U6385 ( .A0(\i_MIPS/Register/register[7][16] ), .A1(net112150), .B0(
        \i_MIPS/Register/register[15][16] ), .B1(net112170), .Y(n8047) );
  OA22XL U6386 ( .A0(\i_MIPS/Register/register[16][13] ), .A1(n4703), .B0(
        \i_MIPS/Register/register[24][13] ), .B1(n4701), .Y(n7772) );
  AO22XL U6387 ( .A0(n4729), .A1(n360), .B0(n4725), .B1(n1068), .Y(n8515) );
  AO22XL U6388 ( .A0(n4729), .A1(n344), .B0(n4725), .B1(n1059), .Y(n8506) );
  AO22XL U6389 ( .A0(n4729), .A1(n345), .B0(n4725), .B1(n1060), .Y(n8325) );
  AO22XL U6390 ( .A0(n4729), .A1(n346), .B0(n4725), .B1(n1061), .Y(n8316) );
  OA22XL U6391 ( .A0(\i_MIPS/Register/register[19][16] ), .A1(net112188), .B0(
        \i_MIPS/Register/register[27][16] ), .B1(n197), .Y(n8057) );
  AO22XL U6392 ( .A0(n4728), .A1(n921), .B0(n4725), .B1(n2627), .Y(n7865) );
  AO22XL U6393 ( .A0(n4731), .A1(n922), .B0(n4725), .B1(n2628), .Y(n7856) );
  AO22XL U6394 ( .A0(n4731), .A1(n923), .B0(n4725), .B1(n2629), .Y(n8215) );
  AO22XL U6395 ( .A0(n9535), .A1(n295), .B0(n4727), .B1(n404), .Y(n8897) );
  AO22XL U6396 ( .A0(n4728), .A1(n361), .B0(n4727), .B1(n1069), .Y(n9536) );
  AO22XL U6397 ( .A0(n4728), .A1(n362), .B0(n4727), .B1(n1070), .Y(n9516) );
  AO22XL U6398 ( .A0(n4728), .A1(n347), .B0(n4727), .B1(n1062), .Y(n9104) );
  AO22XL U6399 ( .A0(n4729), .A1(n348), .B0(n4727), .B1(n1063), .Y(n9095) );
  AO22XL U6400 ( .A0(n4728), .A1(n363), .B0(n4727), .B1(n1071), .Y(n9007) );
  AO22XL U6401 ( .A0(n4728), .A1(n364), .B0(n4727), .B1(n1072), .Y(n8998) );
  AO22XL U6402 ( .A0(n4730), .A1(n924), .B0(n4726), .B1(n2630), .Y(n7117) );
  AO22XL U6403 ( .A0(n4730), .A1(n925), .B0(n4726), .B1(n2631), .Y(n7108) );
  AO22XL U6404 ( .A0(n4730), .A1(n878), .B0(n4726), .B1(n2564), .Y(n6908) );
  AO22XL U6405 ( .A0(n4730), .A1(n879), .B0(n4726), .B1(n2565), .Y(n6899) );
  AO22XL U6406 ( .A0(n4730), .A1(n926), .B0(n4726), .B1(n2632), .Y(n6827) );
  AO22XL U6407 ( .A0(n4730), .A1(n880), .B0(n4726), .B1(n2566), .Y(n6818) );
  OA22XL U6408 ( .A0(\i_MIPS/Register/register[23][16] ), .A1(net112150), .B0(
        \i_MIPS/Register/register[31][16] ), .B1(net112170), .Y(n8056) );
  OA22XL U6409 ( .A0(\i_MIPS/Register/register[17][16] ), .A1(net112254), .B0(
        \i_MIPS/Register/register[25][16] ), .B1(n148), .Y(n8059) );
  OA22XL U6410 ( .A0(\i_MIPS/Register/register[21][16] ), .A1(net112222), .B0(
        \i_MIPS/Register/register[29][16] ), .B1(net112244), .Y(n8058) );
  OA22XL U6411 ( .A0(\i_MIPS/Register/register[19][13] ), .A1(net112188), .B0(
        \i_MIPS/Register/register[27][13] ), .B1(n198), .Y(n7728) );
  OA22XL U6412 ( .A0(\i_MIPS/Register/register[21][8] ), .A1(n192), .B0(
        \i_MIPS/Register/register[29][8] ), .B1(net112242), .Y(n7079) );
  OA22XL U6413 ( .A0(\i_MIPS/Register/register[22][16] ), .A1(net112112), .B0(
        \i_MIPS/Register/register[30][16] ), .B1(net112132), .Y(n8060) );
  MX2XL U6414 ( .A(\I_cache/cache[5][106] ), .B(n10054), .S0(n5229), .Y(n11934) );
  NOR2XL U6415 ( .A(\i_MIPS/Reg_W[4] ), .B(\i_MIPS/Reg_W[3] ), .Y(
        \i_MIPS/forward_unit/n25 ) );
  CLKBUFX2 U6416 ( .A(n5265), .Y(n5242) );
  CLKBUFX3 U6417 ( .A(n5357), .Y(n5354) );
  INVX3 U6418 ( .A(net112158), .Y(net112150) );
  INVX1 U6419 ( .A(n11079), .Y(n11080) );
  NAND2BX2 U6420 ( .AN(n5430), .B(n11231), .Y(n9709) );
  NAND2BX1 U6421 ( .AN(n5425), .B(n11259), .Y(n10038) );
  CLKINVX1 U6422 ( .A(n7171), .Y(n7155) );
  BUFX6 U6423 ( .A(n10194), .Y(n5268) );
  NAND2X1 U6424 ( .A(n9348), .B(n8444), .Y(n8151) );
  INVX1 U6425 ( .A(n7898), .Y(n9334) );
  CLKINVX1 U6426 ( .A(n9283), .Y(n9271) );
  INVX1 U6427 ( .A(n9069), .Y(n9052) );
  CLKINVX1 U6428 ( .A(n6705), .Y(n6481) );
  INVXL U6429 ( .A(n7888), .Y(n7884) );
  INVXL U6430 ( .A(n10520), .Y(n4438) );
  AND2XL U6431 ( .A(net99157), .B(net112799), .Y(n4391) );
  XNOR2X4 U6432 ( .A(n11501), .B(DCACHE_addr[23]), .Y(n6386) );
  OAI211X2 U6433 ( .A0(n7810), .A1(n7809), .B0(n7808), .C0(net112292), .Y(
        n7833) );
  BUFX8 U6434 ( .A(n10192), .Y(n5090) );
  INVX3 U6435 ( .A(n8432), .Y(n8453) );
  AO22X1 U6436 ( .A0(n4712), .A1(n990), .B0(n4708), .B1(n2511), .Y(n7447) );
  AO22X1 U6437 ( .A0(n9531), .A1(n386), .B0(n4716), .B1(n1035), .Y(n7446) );
  AO22X1 U6438 ( .A0(n4712), .A1(n313), .B0(n4708), .B1(n2512), .Y(n7295) );
  AO22X1 U6439 ( .A0(n4712), .A1(n941), .B0(n4708), .B1(n2451), .Y(n7286) );
  AO22X1 U6440 ( .A0(n9531), .A1(n387), .B0(n4716), .B1(n1036), .Y(n7285) );
  AO22X1 U6441 ( .A0(n4712), .A1(n314), .B0(n4708), .B1(n2452), .Y(n7375) );
  AO22X1 U6442 ( .A0(n9531), .A1(n370), .B0(n4716), .B1(n1024), .Y(n7374) );
  AO22X1 U6443 ( .A0(n4712), .A1(n312), .B0(n4708), .B1(n2513), .Y(n7213) );
  AO22X1 U6444 ( .A0(n9531), .A1(n388), .B0(n4716), .B1(n1037), .Y(n7212) );
  AO22X1 U6445 ( .A0(n4712), .A1(n942), .B0(n4708), .B1(n2453), .Y(n7366) );
  AO22X1 U6446 ( .A0(n9531), .A1(n371), .B0(n4716), .B1(n1025), .Y(n7365) );
  AO22X1 U6447 ( .A0(n4712), .A1(n991), .B0(n4708), .B1(n2514), .Y(n7204) );
  AO22X1 U6448 ( .A0(n9531), .A1(n389), .B0(n4716), .B1(n1038), .Y(n7203) );
  AO22X1 U6449 ( .A0(n4712), .A1(n315), .B0(n4708), .B1(n2515), .Y(n7604) );
  AO22X1 U6450 ( .A0(n9531), .A1(n390), .B0(n4716), .B1(n1039), .Y(n7603) );
  AO22X1 U6451 ( .A0(n4712), .A1(n943), .B0(n4708), .B1(n2454), .Y(n7595) );
  AO22X1 U6452 ( .A0(n9531), .A1(n391), .B0(n4716), .B1(n1040), .Y(n7594) );
  OA22XL U6453 ( .A0(n4820), .A1(n1301), .B0(n4866), .B1(n2831), .Y(n8493) );
  NAND2XL U6454 ( .A(n8947), .B(n8253), .Y(n8238) );
  NAND2X1 U6455 ( .A(n6590), .B(\i_MIPS/n346 ), .Y(n9041) );
  OA22X1 U6456 ( .A0(n5204), .A1(n1490), .B0(n5160), .B1(n3235), .Y(n9701) );
  OA22X1 U6457 ( .A0(n5113), .A1(n1491), .B0(n5078), .B1(n3236), .Y(n9702) );
  OA22X1 U6458 ( .A0(n5393), .A1(n1653), .B0(n5339), .B1(n3237), .Y(n9699) );
  OA22XL U6459 ( .A0(n5214), .A1(n1685), .B0(n5171), .B1(n3278), .Y(n10129) );
  OA22XL U6460 ( .A0(n5213), .A1(n1686), .B0(n5170), .B1(n3279), .Y(n10105) );
  OA22XL U6461 ( .A0(n5398), .A1(n1687), .B0(n5348), .B1(n3280), .Y(n10103) );
  OA22XL U6462 ( .A0(n5204), .A1(n1587), .B0(n5160), .B1(n3281), .Y(n9706) );
  OA22XL U6463 ( .A0(n5113), .A1(n1588), .B0(n5069), .B1(n3282), .Y(n9707) );
  OA22XL U6464 ( .A0(n5399), .A1(n1688), .B0(n5339), .B1(n3283), .Y(n9704) );
  OAI22XL U6465 ( .A0(n4754), .A1(n1051), .B0(n4788), .B1(n2646), .Y(n4340) );
  NAND2XL U6466 ( .A(n261), .B(\i_MIPS/n345 ), .Y(n8955) );
  NAND2X1 U6467 ( .A(n8166), .B(n8165), .Y(n8181) );
  INVXL U6468 ( .A(n7692), .Y(n7157) );
  INVX1 U6469 ( .A(n11181), .Y(n11184) );
  CLKAND2X3 U6470 ( .A(n9243), .B(n9137), .Y(n4450) );
  AO22X1 U6471 ( .A0(n4713), .A1(n311), .B0(n4710), .B1(n2455), .Y(n9211) );
  OA22X4 U6472 ( .A0(n5297), .A1(n2169), .B0(n5237), .B1(n595), .Y(n6021) );
  OA22X2 U6473 ( .A0(n230), .A1(n1480), .B0(n5247), .B1(n3054), .Y(n9645) );
  AOI2BB1X1 U6474 ( .A0N(\i_MIPS/ALUin1[14] ), .A1N(n3828), .B0(n4464), .Y(
        n6923) );
  XOR2X4 U6475 ( .A(n10251), .B(ICACHE_addr[16]), .Y(n10627) );
  NAND2X8 U6476 ( .A(n6771), .B(\i_MIPS/ID_EX[83] ), .Y(net101914) );
  MXI2XL U6477 ( .A(n4538), .B(\i_MIPS/n228 ), .S0(n207), .Y(\i_MIPS/n499 ) );
  XNOR2XL U6478 ( .A(\i_MIPS/Reg_W[1] ), .B(\i_MIPS/IR_ID[22] ), .Y(n6443) );
  XNOR2XL U6479 ( .A(\i_MIPS/Reg_W[0] ), .B(\i_MIPS/IR_ID[21] ), .Y(n6441) );
  AO22X1 U6480 ( .A0(net112004), .A1(n392), .B0(net112030), .B1(n1041), .Y(
        n8003) );
  AO22X1 U6481 ( .A0(n4731), .A1(n333), .B0(n4724), .B1(n2435), .Y(n7453) );
  AO22X1 U6482 ( .A0(net112002), .A1(n944), .B0(net112020), .B1(n2456), .Y(
        n7385) );
  AO22X1 U6483 ( .A0(net112002), .A1(n992), .B0(net112020), .B1(n2516), .Y(
        n7394) );
  OA22X1 U6484 ( .A0(n4908), .A1(n1085), .B0(n4947), .B1(n2679), .Y(n9387) );
  OA22X2 U6485 ( .A0(n5297), .A1(n3018), .B0(n5250), .B1(n845), .Y(n9748) );
  OA22X1 U6486 ( .A0(n5398), .A1(n1654), .B0(n5354), .B1(n3238), .Y(n9898) );
  OAI2BB1XL U6487 ( .A0N(n202), .A1N(n3614), .B0(n9971), .Y(\i_MIPS/n480 ) );
  OA22XL U6488 ( .A0(n5394), .A1(n1589), .B0(n5344), .B1(n3167), .Y(n9942) );
  AO21XL U6489 ( .A0(\i_MIPS/ID_EX[88] ), .A1(n202), .B0(n4380), .Y(
        \i_MIPS/n497 ) );
  OA22XL U6490 ( .A0(n5304), .A1(n1303), .B0(n5259), .B1(n3285), .Y(n10128) );
  OA22XL U6491 ( .A0(n4925), .A1(n1773), .B0(n4950), .B1(n3404), .Y(n6433) );
  OA22XL U6492 ( .A0(n4923), .A1(n1304), .B0(n4950), .B1(n2833), .Y(n6804) );
  MX2XL U6493 ( .A(\i_MIPS/ID_EX[43] ), .B(net97755), .S0(n220), .Y(
        \i_MIPS/n433 ) );
  OA22XL U6494 ( .A0(n4922), .A1(n1113), .B0(n4249), .B1(n2659), .Y(n7017) );
  OA22XL U6495 ( .A0(n4915), .A1(n1114), .B0(n4947), .B1(n2660), .Y(n9089) );
  AO22X1 U6496 ( .A0(net112008), .A1(n993), .B0(net112026), .B1(n2517), .Y(
        n9438) );
  AO22X1 U6497 ( .A0(n4729), .A1(n372), .B0(n4725), .B1(n1026), .Y(n8814) );
  AO22X1 U6498 ( .A0(n4729), .A1(n373), .B0(n4725), .B1(n1027), .Y(n8805) );
  AO22X1 U6499 ( .A0(net112008), .A1(n945), .B0(net112026), .B1(n2457), .Y(
        n9447) );
  AO22X1 U6500 ( .A0(n9535), .A1(n300), .B0(n4727), .B1(n403), .Y(n9208) );
  AO22X1 U6501 ( .A0(n4729), .A1(n374), .B0(n4727), .B1(n1028), .Y(n9199) );
  AO22X1 U6502 ( .A0(net112008), .A1(n946), .B0(net112026), .B1(n2458), .Y(
        n8924) );
  OA22X1 U6503 ( .A0(n5291), .A1(n3060), .B0(n5244), .B1(n1150), .Y(n6228) );
  MX2XL U6504 ( .A(\I_cache/cache[4][13] ), .B(n9693), .S0(n5269), .Y(n12679)
         );
  MX2XL U6505 ( .A(\I_cache/cache[4][109] ), .B(n9698), .S0(n5269), .Y(n11911)
         );
  MX2XL U6506 ( .A(\I_cache/cache[3][109] ), .B(n9698), .S0(n5136), .Y(n11912)
         );
  MX2XL U6507 ( .A(\I_cache/cache[4][77] ), .B(n9708), .S0(n5269), .Y(n12167)
         );
  MX2XL U6508 ( .A(\I_cache/cache[3][77] ), .B(n9708), .S0(n5136), .Y(n12168)
         );
  MX2XL U6509 ( .A(\I_cache/cache[4][45] ), .B(n9703), .S0(n5269), .Y(n12423)
         );
  MX2XL U6510 ( .A(\I_cache/cache[3][45] ), .B(n9703), .S0(n5136), .Y(n12424)
         );
  MX2XL U6511 ( .A(\I_cache/cache[6][77] ), .B(n9708), .S0(n5364), .Y(n12165)
         );
  MX2XL U6512 ( .A(\I_cache/cache[6][45] ), .B(n9703), .S0(n5365), .Y(n12421)
         );
  MX2XL U6513 ( .A(\I_cache/cache[1][77] ), .B(n9708), .S0(n5053), .Y(n12170)
         );
  MX2XL U6514 ( .A(\I_cache/cache[1][45] ), .B(n9703), .S0(n5047), .Y(n12426)
         );
  CLKMX2X2 U6515 ( .A(\I_cache/cache[7][12] ), .B(n9764), .S0(n5319), .Y(
        n12684) );
  MX2XL U6516 ( .A(\I_cache/cache[7][13] ), .B(n9693), .S0(n5315), .Y(n12676)
         );
  MX2XL U6517 ( .A(\I_cache/cache[7][109] ), .B(n9698), .S0(n5315), .Y(n11908)
         );
  MX2XL U6518 ( .A(\I_cache/cache[7][77] ), .B(n9708), .S0(n5315), .Y(n12164)
         );
  MX2XL U6519 ( .A(\I_cache/cache[7][45] ), .B(n9703), .S0(n5315), .Y(n12420)
         );
  CLKMX2X2 U6520 ( .A(\I_cache/cache[7][14] ), .B(n9594), .S0(n5314), .Y(
        n12668) );
  MX2XL U6521 ( .A(\I_cache/cache[5][13] ), .B(n9693), .S0(n5226), .Y(n12678)
         );
  MX2XL U6522 ( .A(\I_cache/cache[0][67] ), .B(n11172), .S0(n5092), .Y(n12251)
         );
  MX2XL U6523 ( .A(\I_cache/cache[4][100] ), .B(n11086), .S0(n5277), .Y(n11983) );
  MX2XL U6524 ( .A(\I_cache/cache[3][100] ), .B(n11086), .S0(n5142), .Y(n11984) );
  MX2XL U6525 ( .A(\I_cache/cache[2][100] ), .B(n11086), .S0(n5183), .Y(n11985) );
  MX2XL U6526 ( .A(\I_cache/cache[4][68] ), .B(n11087), .S0(n5277), .Y(n12239)
         );
  MX2XL U6527 ( .A(\I_cache/cache[3][68] ), .B(n11087), .S0(n5135), .Y(n12240)
         );
  MX2XL U6528 ( .A(\I_cache/cache[2][68] ), .B(n11087), .S0(n5186), .Y(n12241)
         );
  MX2XL U6529 ( .A(\I_cache/cache[4][36] ), .B(n11085), .S0(n5277), .Y(n12495)
         );
  MX2XL U6530 ( .A(\I_cache/cache[3][36] ), .B(n11085), .S0(n5140), .Y(n12496)
         );
  MX2XL U6531 ( .A(\I_cache/cache[2][36] ), .B(n11085), .S0(n5181), .Y(n12497)
         );
  MX2XL U6532 ( .A(\I_cache/cache[6][100] ), .B(n11086), .S0(n5362), .Y(n11981) );
  MX2XL U6533 ( .A(\I_cache/cache[6][68] ), .B(n11087), .S0(n5365), .Y(n12237)
         );
  MX2XL U6534 ( .A(\I_cache/cache[6][36] ), .B(n11085), .S0(n5360), .Y(n12493)
         );
  MX2XL U6535 ( .A(\I_cache/cache[5][2] ), .B(n11102), .S0(n5227), .Y(n12766)
         );
  MX2XL U6536 ( .A(\I_cache/cache[7][2] ), .B(n11102), .S0(n5322), .Y(n12764)
         );
  MX2XL U6537 ( .A(\I_cache/cache[5][100] ), .B(n11086), .S0(n5226), .Y(n11982) );
  MX2XL U6538 ( .A(\I_cache/cache[5][68] ), .B(n11087), .S0(n5233), .Y(n12238)
         );
  MX2XL U6539 ( .A(\I_cache/cache[5][36] ), .B(n11085), .S0(n5227), .Y(n12494)
         );
  MX2XL U6540 ( .A(\I_cache/cache[7][100] ), .B(n11086), .S0(n5322), .Y(n11980) );
  MX2XL U6541 ( .A(\I_cache/cache[7][68] ), .B(n11087), .S0(n5322), .Y(n12236)
         );
  MX2XL U6542 ( .A(\I_cache/cache[7][36] ), .B(n11085), .S0(n5322), .Y(n12492)
         );
  MX2XL U6543 ( .A(\I_cache/cache[2][10] ), .B(n10044), .S0(n5186), .Y(n12705)
         );
  MX2XL U6544 ( .A(\I_cache/cache[2][3] ), .B(n11167), .S0(n5189), .Y(n12761)
         );
  MX2XL U6545 ( .A(\I_cache/cache[0][3] ), .B(n11167), .S0(n5098), .Y(n12763)
         );
  MX2XL U6546 ( .A(\I_cache/cache[2][35] ), .B(n11168), .S0(n5189), .Y(n12505)
         );
  MX2XL U6547 ( .A(\I_cache/cache[0][35] ), .B(n11168), .S0(n5098), .Y(n12507)
         );
  MX2XL U6548 ( .A(\I_cache/cache[1][100] ), .B(n11086), .S0(n5045), .Y(n11986) );
  MX2XL U6549 ( .A(\I_cache/cache[1][68] ), .B(n11087), .S0(n5052), .Y(n12242)
         );
  MX2XL U6550 ( .A(\I_cache/cache[1][36] ), .B(n11085), .S0(n5051), .Y(n12498)
         );
  MX2XL U6551 ( .A(\I_cache/cache[6][3] ), .B(n11167), .S0(n5360), .Y(n12757)
         );
  MX2XL U6552 ( .A(\I_cache/cache[6][35] ), .B(n11168), .S0(n5363), .Y(n12501)
         );
  MX2XL U6553 ( .A(\I_cache/cache[4][3] ), .B(n11167), .S0(n5276), .Y(n12759)
         );
  MX2XL U6554 ( .A(\I_cache/cache[4][106] ), .B(n10054), .S0(n5272), .Y(n11935) );
  MX2XL U6555 ( .A(\I_cache/cache[4][10] ), .B(n10044), .S0(n5272), .Y(n12703)
         );
  MX2XL U6556 ( .A(\I_cache/cache[0][100] ), .B(n11086), .S0(n5099), .Y(n11987) );
  MX2XL U6557 ( .A(\I_cache/cache[0][68] ), .B(n11087), .S0(n5099), .Y(n12243)
         );
  MX2XL U6558 ( .A(\I_cache/cache[0][36] ), .B(n11085), .S0(n5099), .Y(n12499)
         );
  MX2XL U6559 ( .A(\I_cache/cache[3][106] ), .B(n10054), .S0(n5140), .Y(n11936) );
  MX2XL U6560 ( .A(\I_cache/cache[6][10] ), .B(n10044), .S0(n5366), .Y(n12701)
         );
  MX2XL U6561 ( .A(\I_cache/cache[1][106] ), .B(n10054), .S0(n5051), .Y(n11938) );
  MX2XL U6562 ( .A(\I_cache/cache[1][10] ), .B(n10044), .S0(n5046), .Y(n12706)
         );
  MX2XL U6563 ( .A(\I_cache/cache[7][106] ), .B(n10054), .S0(n5318), .Y(n11932) );
  OA22XL U6564 ( .A0(n5386), .A1(n1305), .B0(n5330), .B1(n2834), .Y(n6096) );
  OA22XL U6565 ( .A0(n5291), .A1(n3076), .B0(n5244), .B1(n1186), .Y(n6233) );
  OA22XL U6566 ( .A0(n5379), .A1(n3077), .B0(n5333), .B1(n1187), .Y(n6172) );
  CLKINVX2 U6567 ( .A(n4903), .Y(n4899) );
  CLKINVX2 U6568 ( .A(n4909), .Y(n4897) );
  CLKINVX2 U6569 ( .A(n4902), .Y(n4901) );
  CLKINVX3 U6570 ( .A(n5147), .Y(n5138) );
  CLKINVX3 U6571 ( .A(n5208), .Y(n5184) );
  CLKINVX3 U6572 ( .A(n5150), .Y(n5135) );
  CLKINVX3 U6573 ( .A(n5208), .Y(n5181) );
  CLKINVX3 U6574 ( .A(n5117), .Y(n5091) );
  CLKINVX3 U6575 ( .A(n5116), .Y(n5092) );
  CLKINVX3 U6576 ( .A(n5163), .Y(n5141) );
  CLKINVX3 U6577 ( .A(n5208), .Y(n5187) );
  CLKINVX3 U6578 ( .A(n5149), .Y(n5136) );
  CLKINVX3 U6579 ( .A(n5207), .Y(n5182) );
  CLKINVX3 U6580 ( .A(n5117), .Y(n5095) );
  CLKINVX3 U6581 ( .A(n5116), .Y(n5094) );
  CLKINVX3 U6582 ( .A(n5163), .Y(n5140) );
  CLKINVX3 U6583 ( .A(n5208), .Y(n5186) );
  CLKINVX3 U6584 ( .A(n5254), .Y(n5227) );
  CLKINVX3 U6585 ( .A(n5148), .Y(n5137) );
  CLKINVX3 U6586 ( .A(n5207), .Y(n5183) );
  CLKINVX3 U6587 ( .A(n5073), .Y(n5047) );
  CLKINVX3 U6588 ( .A(n5101), .Y(n5093) );
  CLKINVX2 U6589 ( .A(n5010), .Y(n5005) );
  CLKINVX2 U6590 ( .A(n5020), .Y(n5006) );
  CLKINVX2 U6591 ( .A(n5025), .Y(n5009) );
  CLKINVX2 U6592 ( .A(n4787), .Y(n4782) );
  CLKINVX2 U6593 ( .A(n4970), .Y(n4963) );
  CLKINVX2 U6594 ( .A(n4862), .Y(n4853) );
  CLKINVX2 U6595 ( .A(n4760), .Y(n4740) );
  CLKINVX2 U6596 ( .A(n4742), .Y(n4733) );
  CLKINVX2 U6597 ( .A(n4946), .Y(n4939) );
  CLKINVX2 U6598 ( .A(n4981), .Y(n4961) );
  CLKINVX2 U6599 ( .A(n4861), .Y(n4851) );
  CLKINVX2 U6600 ( .A(n4823), .Y(n4807) );
  CLKINVX2 U6601 ( .A(n4966), .Y(n4962) );
  CLKINVX2 U6602 ( .A(n4871), .Y(n4852) );
  CLKINVX2 U6603 ( .A(n4742), .Y(n4734) );
  CLKINVX2 U6604 ( .A(n4742), .Y(n4737) );
  CLKINVX2 U6605 ( .A(n4773), .Y(n4741) );
  CLKINVX2 U6606 ( .A(n4998), .Y(n4965) );
  CLKINVX2 U6607 ( .A(n4870), .Y(n4855) );
  BUFX12 U6608 ( .A(n5085), .Y(n5062) );
  CLKBUFX2 U6609 ( .A(n5264), .Y(n5249) );
  INVX1 U6610 ( .A(n7303), .Y(n7226) );
  CLKBUFX2 U6611 ( .A(n5265), .Y(n5243) );
  CLKBUFX2 U6612 ( .A(n5265), .Y(n5244) );
  CLKBUFX2 U6613 ( .A(n5265), .Y(n5245) );
  CLKBUFX2 U6614 ( .A(n5266), .Y(n5238) );
  CLKBUFX2 U6615 ( .A(n5267), .Y(n5236) );
  BUFX2 U6616 ( .A(n5524), .Y(n5525) );
  CLKBUFX2 U6617 ( .A(n5263), .Y(n5252) );
  CLKBUFX2 U6618 ( .A(n5262), .Y(n5254) );
  CLKBUFX2 U6619 ( .A(n5263), .Y(n5253) );
  CLKINVX3 U6620 ( .A(n5284), .Y(n5271) );
  CLKINVX3 U6621 ( .A(n5282), .Y(n5273) );
  CLKINVX3 U6622 ( .A(n5299), .Y(n5269) );
  CLKINVX3 U6623 ( .A(n5283), .Y(n5272) );
  CLKINVX3 U6624 ( .A(n5290), .Y(n5270) );
  BUFX8 U6625 ( .A(n5133), .Y(n5128) );
  BUFX12 U6626 ( .A(n4681), .Y(n4682) );
  BUFX8 U6627 ( .A(net112014), .Y(net112008) );
  NAND2X2 U6628 ( .A(n4303), .B(n4392), .Y(n10082) );
  INVX3 U6629 ( .A(n7892), .Y(n8874) );
  INVX1 U6630 ( .A(n8073), .Y(n8074) );
  INVXL U6631 ( .A(n8176), .Y(n8177) );
  CLKBUFX2 U6632 ( .A(n5179), .Y(n5175) );
  CLKBUFX2 U6633 ( .A(n5180), .Y(n5174) );
  CLKBUFX2 U6634 ( .A(n5224), .Y(n5217) );
  CLKBUFX2 U6635 ( .A(n4771), .Y(n4772) );
  CLKBUFX2 U6636 ( .A(n4769), .Y(n4773) );
  INVX3 U6637 ( .A(net102048), .Y(net100599) );
  INVXL U6638 ( .A(n8264), .Y(n8265) );
  AND2X2 U6639 ( .A(n3745), .B(n10071), .Y(n4383) );
  INVX4 U6640 ( .A(n4477), .Y(n4699) );
  OR2XL U6641 ( .A(n4649), .B(n10739), .Y(n4622) );
  OR2XL U6642 ( .A(n4649), .B(n10257), .Y(n4606) );
  OR2XL U6643 ( .A(n4649), .B(n10741), .Y(n4604) );
  OR2XL U6644 ( .A(n4649), .B(n10667), .Y(n4605) );
  OR2XL U6645 ( .A(n4649), .B(n10881), .Y(n4603) );
  OR2XL U6646 ( .A(n4649), .B(n10707), .Y(n4600) );
  OR2XL U6647 ( .A(n4649), .B(n10508), .Y(n4602) );
  INVX2 U6648 ( .A(net112176), .Y(net112172) );
  BUFX4 U6649 ( .A(n5532), .Y(n5544) );
  CLKBUFX2 U6650 ( .A(n5179), .Y(n5176) );
  CLKBUFX2 U6651 ( .A(n5223), .Y(n5219) );
  CLKBUFX2 U6652 ( .A(n5356), .Y(n5355) );
  CLKBUFX2 U6653 ( .A(net133468), .Y(net112100) );
  INVXL U6654 ( .A(n11067), .Y(n11069) );
  INVX1 U6655 ( .A(n10550), .Y(n10552) );
  INVX1 U6656 ( .A(n10532), .Y(n10534) );
  INVX1 U6657 ( .A(n11124), .Y(n11126) );
  INVX1 U6658 ( .A(n11175), .Y(n10646) );
  INVX1 U6659 ( .A(n10628), .Y(n10630) );
  INVX1 U6660 ( .A(n10457), .Y(n10459) );
  INVX1 U6661 ( .A(n10840), .Y(n10842) );
  INVX1 U6662 ( .A(n10829), .Y(n10831) );
  INVX1 U6663 ( .A(n10469), .Y(n10470) );
  NAND3BX4 U6664 ( .AN(net103913), .B(n4394), .C(net103910), .Y(n9153) );
  OAI211X2 U6665 ( .A0(n10249), .A1(n10432), .B0(n10622), .C0(n10435), .Y(
        n10336) );
  INVX3 U6666 ( .A(n10433), .Y(n10249) );
  NAND2XL U6667 ( .A(net112294), .B(n8950), .Y(n8976) );
  NAND2BX2 U6668 ( .AN(n5426), .B(n11261), .Y(n9759) );
  NAND2BX2 U6669 ( .AN(n5430), .B(n11229), .Y(n9757) );
  NAND2X2 U6670 ( .A(n4450), .B(n9144), .Y(n8854) );
  AO21X4 U6671 ( .A0(n10567), .A1(n10566), .B0(net111902), .Y(n10455) );
  INVX3 U6672 ( .A(n10858), .Y(n10797) );
  INVX3 U6673 ( .A(n11439), .Y(n10494) );
  INVXL U6674 ( .A(n7708), .Y(n7709) );
  CLKBUFX2 U6675 ( .A(n10639), .Y(n5426) );
  CLKBUFX2 U6676 ( .A(n10640), .Y(n5430) );
  CLKINVX6 U6677 ( .A(n10078), .Y(n10072) );
  NAND2X1 U6678 ( .A(n8731), .B(net101401), .Y(n8734) );
  INVX3 U6679 ( .A(n11380), .Y(n10145) );
  INVX3 U6680 ( .A(n11449), .Y(n9984) );
  INVX3 U6681 ( .A(n11444), .Y(n10142) );
  INVX3 U6682 ( .A(n11431), .Y(n10766) );
  INVX3 U6683 ( .A(n11425), .Y(n10710) );
  MX2X2 U6684 ( .A(n7314), .B(net101401), .S0(net107796), .Y(n6977) );
  NAND2BX4 U6685 ( .AN(n11315), .B(n6122), .Y(n11185) );
  INVX3 U6686 ( .A(n11456), .Y(n10257) );
  INVX3 U6687 ( .A(n11453), .Y(n10881) );
  INVX3 U6688 ( .A(n11441), .Y(n10304) );
  INVX3 U6689 ( .A(n11354), .Y(n10972) );
  INVX3 U6690 ( .A(n11458), .Y(n10719) );
  INVX3 U6691 ( .A(n11450), .Y(n10966) );
  INVX3 U6692 ( .A(n11470), .Y(n10776) );
  INVX3 U6693 ( .A(n11447), .Y(n10905) );
  INVX3 U6694 ( .A(n11455), .Y(n10695) );
  INVXL U6695 ( .A(n8553), .Y(n9272) );
  NAND2BXL U6696 ( .AN(n5427), .B(n11213), .Y(n6257) );
  INVX3 U6697 ( .A(n11440), .Y(n10272) );
  INVXL U6698 ( .A(n7502), .Y(n7514) );
  INVX3 U6699 ( .A(n9412), .Y(n9533) );
  INVX3 U6700 ( .A(n9410), .Y(n9535) );
  INVX3 U6701 ( .A(n9415), .Y(n9530) );
  INVX3 U6702 ( .A(n9416), .Y(n9529) );
  INVX3 U6703 ( .A(n9417), .Y(n9528) );
  INVX3 U6704 ( .A(net102051), .Y(net100601) );
  MX2XL U6705 ( .A(net112438), .B(net100573), .S0(n8166), .Y(n8160) );
  INVXL U6706 ( .A(n10319), .Y(n10838) );
  NAND2BXL U6707 ( .AN(n5428), .B(n11212), .Y(n6277) );
  INVX1 U6708 ( .A(n6708), .Y(n6709) );
  AND2XL U6709 ( .A(n10222), .B(n10221), .Y(n4411) );
  INVXL U6710 ( .A(n7896), .Y(n7905) );
  INVX1 U6711 ( .A(n7808), .Y(n7802) );
  INVXL U6712 ( .A(n8747), .Y(n8757) );
  AND2XL U6713 ( .A(net97686), .B(net97687), .Y(n4407) );
  AND2XL U6714 ( .A(n3421), .B(net99161), .Y(n4408) );
  AND2XL U6715 ( .A(n3426), .B(net99118), .Y(n4406) );
  AND2XL U6716 ( .A(n3422), .B(n10584), .Y(n4404) );
  AND2XL U6717 ( .A(n3722), .B(net98231), .Y(n4396) );
  AND2XL U6718 ( .A(n3425), .B(net98755), .Y(n4430) );
  AND2XL U6719 ( .A(n3419), .B(n10519), .Y(n4399) );
  NAND2BXL U6720 ( .AN(n5426), .B(n11270), .Y(n9637) );
  NAND2BXL U6721 ( .AN(n5430), .B(n11238), .Y(n9635) );
  NAND2BXL U6722 ( .AN(n5426), .B(n11268), .Y(n9686) );
  NAND2BXL U6723 ( .AN(n5430), .B(n11236), .Y(n9684) );
  NAND2BXL U6724 ( .AN(n5425), .B(n11269), .Y(n9589) );
  NAND2BXL U6725 ( .AN(n5429), .B(n11237), .Y(n9587) );
  NAND2BXL U6726 ( .AN(n5426), .B(n11267), .Y(n10643) );
  NAND2BXL U6727 ( .AN(n5430), .B(n11235), .Y(n10641) );
  NAND2BXL U6728 ( .AN(n5426), .B(n11266), .Y(n9735) );
  NAND2BXL U6729 ( .AN(n5430), .B(n11234), .Y(n9733) );
  NAND2BXL U6730 ( .AN(n5426), .B(n11272), .Y(n9880) );
  NAND2BXL U6731 ( .AN(n5430), .B(n11240), .Y(n9878) );
  NAND2BXL U6732 ( .AN(n5426), .B(n11271), .Y(net99634) );
  NAND2BXL U6733 ( .AN(n5430), .B(n11239), .Y(net99636) );
  NAND2BXL U6734 ( .AN(n5426), .B(n11275), .Y(n9824) );
  NAND2BXL U6735 ( .AN(n5430), .B(n11243), .Y(n9822) );
  NAND2BXL U6736 ( .AN(n5426), .B(n11274), .Y(n9804) );
  NAND2BXL U6737 ( .AN(n5430), .B(n11242), .Y(n9802) );
  NAND2BXL U6738 ( .AN(n5426), .B(n11273), .Y(n9844) );
  NAND2BXL U6739 ( .AN(n5430), .B(n11241), .Y(n9842) );
  INVXL U6740 ( .A(n10313), .Y(n10314) );
  INVX1 U6741 ( .A(n9891), .Y(n9887) );
  CLKBUFX2 U6742 ( .A(n4478), .Y(n4696) );
  NAND2XL U6743 ( .A(n6966), .B(n7876), .Y(n7048) );
  AO21X4 U6744 ( .A0(net98372), .A1(net98371), .B0(net111642), .Y(net103956)
         );
  OAI2BB1X4 U6745 ( .A0N(n10526), .A1N(n10525), .B0(net112782), .Y(net102939)
         );
  OAI31X2 U6746 ( .A0(n6509), .A1(n6508), .A2(n6507), .B0(n6506), .Y(n7407) );
  OA22X1 U6747 ( .A0(n4984), .A1(n1229), .B0(n5030), .B1(n2766), .Y(n6892) );
  OA22XL U6748 ( .A0(n4759), .A1(n1306), .B0(n4796), .B1(n2835), .Y(n6895) );
  OA22XL U6749 ( .A0(n4819), .A1(n2960), .B0(n4865), .B1(n1422), .Y(n8601) );
  INVXL U6750 ( .A(n8642), .Y(n8647) );
  NAND2XL U6751 ( .A(n8642), .B(n8641), .Y(n8643) );
  INVXL U6752 ( .A(n8341), .Y(n8346) );
  AO21X4 U6753 ( .A0(n10568), .A1(n4608), .B0(net111642), .Y(n8225) );
  XOR2X4 U6754 ( .A(n11505), .B(DCACHE_addr[27]), .Y(n6424) );
  AO21X4 U6755 ( .A0(n10412), .A1(n10410), .B0(n4474), .Y(n10416) );
  AO21X4 U6756 ( .A0(n10378), .A1(n10373), .B0(n4475), .Y(n10244) );
  AO21X4 U6757 ( .A0(n10818), .A1(n10816), .B0(n4466), .Y(n10384) );
  NOR4X1 U6758 ( .A(n6667), .B(n6666), .C(n6665), .D(n6664), .Y(n6678) );
  AO21X4 U6759 ( .A0(n10617), .A1(n10615), .B0(n4465), .Y(n10432) );
  AO22X4 U6760 ( .A0(net111960), .A1(n9074), .B0(net111968), .B1(n10487), .Y(
        n9075) );
  AO21X4 U6761 ( .A0(n10520), .A1(net98380), .B0(net111642), .Y(net103583) );
  OA21XL U6762 ( .A0(n8542), .A1(n8540), .B0(n8736), .Y(n8541) );
  AO21X4 U6763 ( .A0(n11098), .A1(n11096), .B0(n4435), .Y(n10360) );
  MX2XL U6764 ( .A(net100573), .B(net112438), .S0(n6481), .Y(n6489) );
  NAND4BX2 U6765 ( .AN(n6476), .B(n6475), .C(n6474), .D(n6473), .Y(n6477) );
  NAND4BX2 U6766 ( .AN(n8575), .B(n8574), .C(n8573), .D(n8572), .Y(n8586) );
  MX2X2 U6767 ( .A(n8586), .B(n8585), .S0(\i_MIPS/IR_ID[25] ), .Y(n8606) );
  NAND3BX4 U6768 ( .AN(n4664), .B(n4295), .C(n4666), .Y(n9988) );
  INVX1 U6769 ( .A(n8070), .Y(n7799) );
  NAND2X2 U6770 ( .A(n6694), .B(\i_MIPS/n340 ), .Y(n11177) );
  INVX3 U6771 ( .A(net111646), .Y(net111644) );
  NAND4X2 U6772 ( .A(n6019), .B(n6018), .C(n6017), .D(n6016), .Y(n11325) );
  NAND4BX2 U6773 ( .AN(n4338), .B(n10034), .C(n10033), .D(n10032), .Y(n11227)
         );
  OA22XL U6774 ( .A0(n5111), .A1(n1690), .B0(n5061), .B1(n3286), .Y(n10011) );
  OA22XL U6775 ( .A0(n5388), .A1(n1691), .B0(n5345), .B1(n3287), .Y(n10008) );
  NAND4X2 U6776 ( .A(n10025), .B(n10024), .C(n10023), .D(n10022), .Y(n11259)
         );
  OA22XL U6777 ( .A0(n5212), .A1(n1693), .B0(n5169), .B1(n3289), .Y(n10029) );
  OA22XL U6778 ( .A0(n5121), .A1(n1694), .B0(n5071), .B1(n3290), .Y(n10030) );
  OA22XL U6779 ( .A0(n5373), .A1(n1695), .B0(n5346), .B1(n3291), .Y(n10027) );
  OA22XL U6780 ( .A0(n5214), .A1(n1696), .B0(n5171), .B1(n3292), .Y(n10119) );
  OA22XL U6781 ( .A0(n5126), .A1(n1697), .B0(n5065), .B1(n3293), .Y(n10006) );
  NAND4X2 U6782 ( .A(n10115), .B(n10114), .C(n10113), .D(n10112), .Y(n11289)
         );
  OA22XL U6783 ( .A0(n5213), .A1(n1698), .B0(n5170), .B1(n3294), .Y(n10100) );
  OA22XL U6784 ( .A0(n5122), .A1(n1699), .B0(n5063), .B1(n3295), .Y(n10101) );
  OA22XL U6785 ( .A0(n5368), .A1(n1700), .B0(n5348), .B1(n3296), .Y(n10098) );
  NAND4X2 U6786 ( .A(n10096), .B(n10095), .C(n10094), .D(n10093), .Y(n11256)
         );
  OA22XL U6787 ( .A0(n5213), .A1(n1701), .B0(n5170), .B1(n3297), .Y(n10095) );
  OA22XL U6788 ( .A0(n5122), .A1(n1702), .B0(n5085), .B1(n3298), .Y(n10096) );
  OA22XL U6789 ( .A0(n5367), .A1(n1703), .B0(n5348), .B1(n3299), .Y(n10093) );
  NAND4X2 U6790 ( .A(n9707), .B(n9706), .C(n9705), .D(n9704), .Y(n11231) );
  NAND4X2 U6791 ( .A(n9702), .B(n9701), .C(n9700), .D(n9699), .Y(n11263) );
  NAND4X2 U6792 ( .A(n9692), .B(n9691), .C(n9690), .D(n9689), .Y(n11295) );
  NAND4X2 U6793 ( .A(n10058), .B(n10057), .C(n10056), .D(n10055), .Y(n11228)
         );
  OA22XL U6794 ( .A0(n5213), .A1(n1590), .B0(n5170), .B1(n3168), .Y(n10057) );
  OA22XL U6795 ( .A0(n5122), .A1(n1591), .B0(n5072), .B1(n3169), .Y(n10058) );
  OA22XL U6796 ( .A0(n5378), .A1(n1592), .B0(n5348), .B1(n3170), .Y(n10055) );
  OA22XL U6797 ( .A0(n4830), .A1(n1128), .B0(n4861), .B1(n2661), .Y(n9194) );
  OA22XL U6798 ( .A0(n4754), .A1(n2767), .B0(n4788), .B1(n1121), .Y(n9195) );
  OA22XL U6799 ( .A0(n4757), .A1(n1307), .B0(n4796), .B1(n2836), .Y(n7104) );
  OA22X1 U6800 ( .A0(n4980), .A1(n1230), .B0(n5026), .B1(n2768), .Y(n7356) );
  OA22X1 U6801 ( .A0(n4828), .A1(n1231), .B0(n4873), .B1(n2769), .Y(n7358) );
  OA22XL U6802 ( .A0(n4755), .A1(n1308), .B0(n4793), .B1(n2837), .Y(n7359) );
  OA22XL U6803 ( .A0(n4968), .A1(n2729), .B0(n5027), .B1(n1188), .Y(n9188) );
  OA22XL U6804 ( .A0(n4830), .A1(n1309), .B0(n4861), .B1(n2838), .Y(n9190) );
  OA22XL U6805 ( .A0(n4743), .A1(n2961), .B0(n4788), .B1(n1423), .Y(n9191) );
  NAND4X2 U6806 ( .A(n8895), .B(n8894), .C(n8893), .D(n8892), .Y(n11405) );
  OA22XL U6807 ( .A0(n4832), .A1(n1310), .B0(n4877), .B1(n2839), .Y(n6886) );
  OA22XL U6808 ( .A0(n4760), .A1(n1311), .B0(n4796), .B1(n2840), .Y(n6887) );
  OA22XL U6809 ( .A0(n4828), .A1(n1312), .B0(n4873), .B1(n2841), .Y(n7350) );
  OA22XL U6810 ( .A0(n4743), .A1(n2962), .B0(n4789), .B1(n1189), .Y(n9087) );
  OA22XL U6811 ( .A0(n4821), .A1(n1313), .B0(n4867), .B1(n2842), .Y(n8303) );
  OA22XL U6812 ( .A0(n4974), .A1(n1314), .B0(n5019), .B1(n2843), .Y(n8305) );
  OA22XL U6813 ( .A0(n4821), .A1(n1315), .B0(n4867), .B1(n2844), .Y(n8307) );
  OA22XL U6814 ( .A0(n4749), .A1(n1316), .B0(n4790), .B1(n2845), .Y(n8308) );
  OA22XL U6815 ( .A0(n4745), .A1(n2770), .B0(n4789), .B1(n1122), .Y(n8801) );
  OA22XL U6816 ( .A0(n4830), .A1(n1317), .B0(n4875), .B1(n2846), .Y(n7099) );
  OA22XL U6817 ( .A0(n4757), .A1(n1318), .B0(n4796), .B1(n2847), .Y(n7100) );
  OA22XL U6818 ( .A0(n4752), .A1(n1115), .B0(n4792), .B1(n2662), .Y(n7852) );
  OA22XL U6819 ( .A0(n4818), .A1(n1151), .B0(n263), .B1(n2708), .Y(n8792) );
  OA22XL U6820 ( .A0(n4745), .A1(n2963), .B0(n4789), .B1(n1190), .Y(n8793) );
  OA22XL U6821 ( .A0(n4976), .A1(n1319), .B0(n185), .B1(n2848), .Y(n8013) );
  OA22XL U6822 ( .A0(n4751), .A1(n1320), .B0(n4791), .B1(n2849), .Y(n8016) );
  OA22XL U6823 ( .A0(n4976), .A1(n1321), .B0(n185), .B1(n2850), .Y(n7943) );
  OA22XL U6824 ( .A0(n4751), .A1(n1322), .B0(n4791), .B1(n2851), .Y(n7946) );
  OA22XL U6825 ( .A0(n4980), .A1(n1323), .B0(n5026), .B1(n2852), .Y(n7352) );
  OA22XL U6826 ( .A0(n4828), .A1(n1324), .B0(n4873), .B1(n2853), .Y(n7354) );
  OA22XL U6827 ( .A0(n4973), .A1(n1325), .B0(n5018), .B1(n2854), .Y(n8392) );
  OA22XL U6828 ( .A0(n4820), .A1(n1326), .B0(n4866), .B1(n2855), .Y(n8394) );
  OA22XL U6829 ( .A0(n4748), .A1(n1327), .B0(n4790), .B1(n2856), .Y(n8395) );
  OA22XL U6830 ( .A0(n4981), .A1(n1328), .B0(n5027), .B1(n2857), .Y(n7190) );
  OA22XL U6831 ( .A0(n4829), .A1(n1329), .B0(n4874), .B1(n2858), .Y(n7192) );
  OA22XL U6832 ( .A0(n4754), .A1(n2964), .B0(n4792), .B1(n1191), .Y(n7580) );
  OA22XL U6833 ( .A0(n4980), .A1(n1152), .B0(n5026), .B1(n2709), .Y(n7272) );
  OA22XL U6834 ( .A0(n4828), .A1(n1153), .B0(n4873), .B1(n2710), .Y(n7274) );
  OA22XL U6835 ( .A0(n4756), .A1(n2965), .B0(n4793), .B1(n1192), .Y(n7275) );
  OA22XL U6836 ( .A0(n4745), .A1(n2966), .B0(n4789), .B1(n1123), .Y(n8891) );
  OA22XL U6837 ( .A0(n4744), .A1(n1330), .B0(n4789), .B1(n2859), .Y(n8994) );
  OA22XL U6838 ( .A0(n4818), .A1(n1154), .B0(n263), .B1(n2711), .Y(n8796) );
  OA22XL U6839 ( .A0(n4818), .A1(n1331), .B0(n263), .B1(n2860), .Y(n8694) );
  OA22XL U6840 ( .A0(n4751), .A1(n1332), .B0(n4791), .B1(n2861), .Y(n8020) );
  OA22XL U6841 ( .A0(n4977), .A1(n1333), .B0(n5022), .B1(n2862), .Y(n7935) );
  OA22XL U6842 ( .A0(n4751), .A1(n1334), .B0(n4791), .B1(n2863), .Y(n7938) );
  NAND4X2 U6843 ( .A(n7584), .B(n7583), .C(n7582), .D(n7581), .Y(n11350) );
  OA22XL U6844 ( .A0(n4826), .A1(n1335), .B0(n4871), .B1(n2864), .Y(n7583) );
  OA22XL U6845 ( .A0(n4754), .A1(n1336), .B0(n4792), .B1(n2865), .Y(n7584) );
  NAND4X2 U6846 ( .A(n6931), .B(n6930), .C(n6929), .D(n6928), .Y(n11416) );
  OAI22XL U6847 ( .A0(n4773), .A1(n1052), .B0(n4788), .B1(n2650), .Y(n4342) );
  OA22XL U6848 ( .A0(n4977), .A1(n1337), .B0(n5022), .B1(n2866), .Y(n7939) );
  OA22XL U6849 ( .A0(n4751), .A1(n1338), .B0(n4791), .B1(n2867), .Y(n7942) );
  OA22XL U6850 ( .A0(n4819), .A1(n1339), .B0(n4865), .B1(n2868), .Y(n8501) );
  OA22XL U6851 ( .A0(n4750), .A1(n2967), .B0(n4791), .B1(n1193), .Y(n8099) );
  OA22XL U6852 ( .A0(n4982), .A1(n1155), .B0(n5028), .B1(n2712), .Y(n7012) );
  OA22XL U6853 ( .A0(n4830), .A1(n1156), .B0(n4875), .B1(n2713), .Y(n7014) );
  OA22XL U6854 ( .A0(n4758), .A1(n2968), .B0(n4796), .B1(n1194), .Y(n7015) );
  OA22XL U6855 ( .A0(n4983), .A1(n1340), .B0(n5029), .B1(n2869), .Y(n6924) );
  OA22XL U6856 ( .A0(n4831), .A1(n1341), .B0(n4876), .B1(n2870), .Y(n6926) );
  OA22XL U6857 ( .A0(n4759), .A1(n1342), .B0(n4796), .B1(n2871), .Y(n6927) );
  OA22XL U6858 ( .A0(n4825), .A1(n1343), .B0(n4870), .B1(n2872), .Y(n7749) );
  OAI22XL U6859 ( .A0(n4773), .A1(n2647), .B0(n4788), .B1(n1074), .Y(n4343) );
  OA22XL U6860 ( .A0(n4753), .A1(n1344), .B0(n4792), .B1(n2873), .Y(n7656) );
  OA22XL U6861 ( .A0(n4820), .A1(n1345), .B0(n4866), .B1(n2874), .Y(n8497) );
  OA22XL U6862 ( .A0(n4983), .A1(n1346), .B0(n5029), .B1(n2875), .Y(n6932) );
  OA22XL U6863 ( .A0(n4831), .A1(n1347), .B0(n4876), .B1(n2876), .Y(n6934) );
  OA22XL U6864 ( .A0(n4759), .A1(n1348), .B0(n4796), .B1(n2877), .Y(n6935) );
  NAND4X2 U6865 ( .A(n8202), .B(n8201), .C(n8200), .D(n8199), .Y(n11411) );
  OA22XL U6866 ( .A0(n4821), .A1(n1130), .B0(n4867), .B1(n2664), .Y(n8201) );
  OA22XL U6867 ( .A0(n4749), .A1(n1117), .B0(n4791), .B1(n2665), .Y(n8202) );
  OA22XL U6868 ( .A0(n5211), .A1(n1704), .B0(n5168), .B1(n3300), .Y(n10019) );
  OA22XL U6869 ( .A0(n5114), .A1(n1705), .B0(n181), .B1(n3301), .Y(n10020) );
  OA22XL U6870 ( .A0(n5126), .A1(n1593), .B0(n5081), .B1(n3303), .Y(n9996) );
  OA22XL U6871 ( .A0(n5394), .A1(n1707), .B0(n5345), .B1(n3304), .Y(n9993) );
  OA22XL U6872 ( .A0(n4968), .A1(n1157), .B0(n5027), .B1(n2714), .Y(n9288) );
  OA22XL U6873 ( .A0(n4830), .A1(n1349), .B0(n4861), .B1(n2878), .Y(n9290) );
  OA22XL U6874 ( .A0(n4754), .A1(n2970), .B0(n4788), .B1(n1424), .Y(n9291) );
  NAND4X2 U6875 ( .A(n7279), .B(n7278), .C(n7277), .D(n7276), .Y(n11393) );
  OA22XL U6876 ( .A0(n4980), .A1(n1131), .B0(n5026), .B1(n2666), .Y(n7276) );
  OA22XL U6877 ( .A0(n4756), .A1(n1118), .B0(n4793), .B1(n2667), .Y(n7279) );
  OA22XL U6878 ( .A0(n4745), .A1(n2971), .B0(n4789), .B1(n1196), .Y(n8884) );
  OA22XL U6879 ( .A0(n4820), .A1(n1158), .B0(n4866), .B1(n2715), .Y(n8489) );
  NAND2XL U6880 ( .A(n9457), .B(n8852), .Y(n7541) );
  INVXL U6881 ( .A(n7409), .Y(n7232) );
  NAND4X2 U6882 ( .A(n7840), .B(n7839), .C(n7838), .D(n7837), .Y(n11463) );
  AO22XL U6883 ( .A0(n4711), .A1(n418), .B0(n4709), .B1(n2567), .Y(n8817) );
  AO22XL U6884 ( .A0(n4713), .A1(n308), .B0(n4710), .B1(n2568), .Y(n8909) );
  AO22XL U6885 ( .A0(n4720), .A1(n881), .B0(n4719), .B1(n2569), .Y(n8907) );
  AO22XL U6886 ( .A0(n4712), .A1(n419), .B0(n4708), .B1(n2633), .Y(n7456) );
  AO22XL U6887 ( .A0(n9531), .A1(n365), .B0(n4716), .B1(n1073), .Y(n7455) );
  AO22XL U6888 ( .A0(n4721), .A1(n296), .B0(n4719), .B1(n2570), .Y(n7293) );
  AO22XL U6889 ( .A0(n4722), .A1(n297), .B0(n4719), .B1(n2571), .Y(n7284) );
  AO22XL U6890 ( .A0(n4722), .A1(n298), .B0(n4719), .B1(n2572), .Y(n7373) );
  INVX3 U6891 ( .A(n10410), .Y(n10408) );
  NAND2XL U6892 ( .A(n9041), .B(n9040), .Y(n9067) );
  INVX3 U6893 ( .A(n10615), .Y(n10613) );
  NAND2X2 U6894 ( .A(n10138), .B(n4525), .Y(n10173) );
  OA22XL U6895 ( .A0(n4744), .A1(n2972), .B0(n4789), .B1(n1197), .Y(n8986) );
  OA22XL U6896 ( .A0(n4752), .A1(n2973), .B0(n4792), .B1(n1285), .Y(n7844) );
  OA22XL U6897 ( .A0(n4748), .A1(n1350), .B0(n4790), .B1(n2880), .Y(n8391) );
  OA22XL U6898 ( .A0(n4821), .A1(n1351), .B0(n4867), .B1(n2881), .Y(n8390) );
  OA22XL U6899 ( .A0(n4754), .A1(n3333), .B0(n4793), .B1(n1198), .Y(n7576) );
  OA22XL U6900 ( .A0(n4827), .A1(n3078), .B0(n4872), .B1(n1427), .Y(n7575) );
  NAND2X1 U6901 ( .A(n6612), .B(n4502), .Y(n4349) );
  OA22XL U6902 ( .A0(n4825), .A1(n1594), .B0(n4870), .B1(n3171), .Y(n4351) );
  INVXL U6903 ( .A(n9040), .Y(n9056) );
  CLKMX2X4 U6904 ( .A(n7059), .B(n4520), .S0(net107794), .Y(n9251) );
  AO22XL U6905 ( .A0(n4720), .A1(n882), .B0(n4719), .B1(n2573), .Y(n8898) );
  OA22XL U6906 ( .A0(n4754), .A1(n2974), .B0(n4792), .B1(n1199), .Y(n4352) );
  NAND4X2 U6907 ( .A(n4353), .B(n8887), .C(n8886), .D(n8885), .Y(n11437) );
  OA22XL U6908 ( .A0(n4745), .A1(n2975), .B0(n4789), .B1(n1200), .Y(n4353) );
  OA22XL U6909 ( .A0(n4754), .A1(n1352), .B0(n4788), .B1(n2882), .Y(n4354) );
  NAND4X2 U6910 ( .A(n4355), .B(n7007), .C(n7006), .D(n7005), .Y(n11452) );
  OA22XL U6911 ( .A0(n4758), .A1(n1353), .B0(n4796), .B1(n2883), .Y(n4355) );
  OA22X4 U6912 ( .A0(n5118), .A1(n2170), .B0(n5059), .B1(n596), .Y(n6015) );
  OA22X4 U6913 ( .A0(n5193), .A1(n2171), .B0(n5146), .B1(n597), .Y(n6014) );
  OA22X4 U6914 ( .A0(n5283), .A1(n2172), .B0(n5237), .B1(n598), .Y(n6013) );
  OA22X4 U6915 ( .A0(n5130), .A1(n2173), .B0(n5083), .B1(n599), .Y(n5990) );
  OA22X4 U6916 ( .A0(n5191), .A1(n2174), .B0(n5144), .B1(n600), .Y(n5989) );
  OA22X4 U6917 ( .A0(n5280), .A1(n2175), .B0(n5257), .B1(n601), .Y(n5988) );
  OA22X4 U6918 ( .A0(n5191), .A1(n2180), .B0(n5165), .B1(n606), .Y(n5975) );
  OA22X4 U6919 ( .A0(n5298), .A1(n2181), .B0(n5234), .B1(n607), .Y(n5974) );
  OA22X4 U6920 ( .A0(n5130), .A1(n2182), .B0(n5059), .B1(n608), .Y(n5986) );
  OA22X4 U6921 ( .A0(n5190), .A1(n2183), .B0(n5144), .B1(n609), .Y(n5985) );
  OA22X4 U6922 ( .A0(n5279), .A1(n2184), .B0(n5235), .B1(n610), .Y(n5984) );
  MX2XL U6923 ( .A(net100573), .B(net112438), .S0(n9046), .Y(n9049) );
  AND2XL U6924 ( .A(n7497), .B(n7500), .Y(n7240) );
  AND2XL U6925 ( .A(n3636), .B(n7405), .Y(n7243) );
  NAND2XL U6926 ( .A(DCACHE_addr[27]), .B(\i_MIPS/n336 ), .Y(n10568) );
  NAND2XL U6927 ( .A(n11178), .B(n11177), .Y(n6695) );
  NAND2XL U6928 ( .A(n7053), .B(\i_MIPS/n363 ), .Y(n8633) );
  NAND2XL U6929 ( .A(n4664), .B(n4673), .Y(net98780) );
  NAND2XL U6930 ( .A(DCACHE_addr[6]), .B(n4673), .Y(net98390) );
  NAND2XL U6931 ( .A(DCACHE_addr[22]), .B(\i_MIPS/n336 ), .Y(n10567) );
  NAND2XL U6932 ( .A(DCACHE_addr[8]), .B(n4673), .Y(net98758) );
  NAND2XL U6933 ( .A(DCACHE_addr[13]), .B(n4673), .Y(net98385) );
  NAND2XL U6934 ( .A(DCACHE_addr[9]), .B(n4673), .Y(net98776) );
  NAND2XL U6935 ( .A(DCACHE_addr[7]), .B(\i_MIPS/n336 ), .Y(n10561) );
  AO22XL U6936 ( .A0(net112178), .A1(n265), .B0(net112160), .B1(n2011), .Y(
        n6472) );
  AO22XL U6937 ( .A0(n195), .A1(n421), .B0(net112196), .B1(n2012), .Y(n6471)
         );
  AO22XL U6938 ( .A0(net112178), .A1(n424), .B0(net112160), .B1(n2003), .Y(
        n6463) );
  AO22XL U6939 ( .A0(n195), .A1(n422), .B0(net112196), .B1(n2013), .Y(n6462)
         );
  AO22XL U6940 ( .A0(n195), .A1(n318), .B0(net112196), .B1(n2005), .Y(n8579)
         );
  AO22XL U6941 ( .A0(net112178), .A1(n425), .B0(net112160), .B1(n2006), .Y(
        n8571) );
  AO22XL U6942 ( .A0(n195), .A1(n319), .B0(net112196), .B1(n2007), .Y(n8570)
         );
  CLKBUFX2 U6943 ( .A(\i_MIPS/n336 ), .Y(n4674) );
  INVX3 U6944 ( .A(n11078), .Y(n11077) );
  NAND2XL U6945 ( .A(n8753), .B(n8749), .Y(n8077) );
  NAND2XL U6946 ( .A(n6612), .B(n4445), .Y(n9527) );
  AOI2BB1XL U6947 ( .A0N(n8440), .A1N(net102253), .B0(n4516), .Y(n6495) );
  AND2XL U6948 ( .A(n10281), .B(n10282), .Y(n4442) );
  AND2XL U6949 ( .A(n10152), .B(n10151), .Y(n4458) );
  NAND2XL U6950 ( .A(n8633), .B(n7219), .Y(n7054) );
  OA22X4 U6951 ( .A0(n5130), .A1(n2185), .B0(n5086), .B1(n611), .Y(n5996) );
  OA22X4 U6952 ( .A0(n5192), .A1(n2186), .B0(n5145), .B1(n612), .Y(n5995) );
  OA22X4 U6953 ( .A0(n5281), .A1(n2187), .B0(n5236), .B1(n613), .Y(n5994) );
  INVXL U6954 ( .A(n8753), .Y(n7810) );
  NOR3X1 U6955 ( .A(n303), .B(n415), .C(n4534), .Y(\i_MIPS/Register/n105 ) );
  OA22XL U6956 ( .A0(n5293), .A1(n1853), .B0(n5246), .B1(n3509), .Y(n9584) );
  OA22XL U6957 ( .A0(n5109), .A1(n1854), .B0(n5083), .B1(n3510), .Y(n9578) );
  OA22XL U6958 ( .A0(n5292), .A1(n1855), .B0(n5245), .B1(n3511), .Y(n9576) );
  OA22XL U6959 ( .A0(n5200), .A1(n1856), .B0(n5164), .B1(n3512), .Y(n9577) );
  NAND4BX1 U6960 ( .AN(n4357), .B(n9820), .C(n9819), .D(n9818), .Y(n11243) );
  OAI22XL U6961 ( .A0(n5116), .A1(n1777), .B0(n5066), .B1(n3433), .Y(n4357) );
  NAND4BX1 U6962 ( .AN(n4358), .B(n9812), .C(n9811), .D(n9810), .Y(n11275) );
  OAI22XL U6963 ( .A0(n5116), .A1(n1778), .B0(n5082), .B1(n3434), .Y(n4358) );
  NAND4BX1 U6964 ( .AN(n4359), .B(n9800), .C(n9799), .D(n9798), .Y(n11242) );
  OAI22XL U6965 ( .A0(n5116), .A1(n1779), .B0(n5074), .B1(n3435), .Y(n4359) );
  OA22XL U6966 ( .A0(n5298), .A1(n1857), .B0(n5251), .B1(n3513), .Y(n9790) );
  NAND4BX1 U6967 ( .AN(n4360), .B(n9840), .C(n9839), .D(n9838), .Y(n11241) );
  OAI22XL U6968 ( .A0(n5117), .A1(n1780), .B0(n5078), .B1(n3436), .Y(n4360) );
  NAND4BX1 U6969 ( .AN(n4361), .B(n9832), .C(n9831), .D(n9830), .Y(n11273) );
  OAI22XL U6970 ( .A0(n5117), .A1(n1781), .B0(n5075), .B1(n3437), .Y(n4361) );
  NAND4BX1 U6971 ( .AN(n4362), .B(n9876), .C(n9875), .D(n9874), .Y(n11240) );
  OAI22XL U6972 ( .A0(n5118), .A1(n1782), .B0(n5071), .B1(n3438), .Y(n4362) );
  NAND4BX1 U6973 ( .AN(n4363), .B(n9868), .C(n9867), .D(n9866), .Y(n11272) );
  OAI22XL U6974 ( .A0(n5118), .A1(n1783), .B0(n5064), .B1(n3439), .Y(n4363) );
  NAND4BX1 U6975 ( .AN(n4364), .B(n9860), .C(n9859), .D(n9858), .Y(n11239) );
  OAI22XL U6976 ( .A0(n5118), .A1(n1784), .B0(n5054), .B1(n3440), .Y(n4364) );
  NAND4BX1 U6977 ( .AN(n4365), .B(n9852), .C(n9851), .D(n9850), .Y(n11271) );
  OAI22XL U6978 ( .A0(n5117), .A1(n1785), .B0(n5070), .B1(n3441), .Y(n4365) );
  OA22XL U6979 ( .A0(n5297), .A1(n1858), .B0(n5250), .B1(n3514), .Y(n9729) );
  OA22XL U6980 ( .A0(n5295), .A1(n1859), .B0(n5248), .B1(n3515), .Y(n9675) );
  OA22XL U6981 ( .A0(n5203), .A1(n1860), .B0(n5159), .B1(n3516), .Y(n9676) );
  OA22XL U6982 ( .A0(n5295), .A1(n1861), .B0(n5248), .B1(n3517), .Y(n9665) );
  OA22XL U6983 ( .A0(n5203), .A1(n1862), .B0(n5159), .B1(n3518), .Y(n9666) );
  OA22XL U6984 ( .A0(n5293), .A1(n1863), .B0(n5246), .B1(n3519), .Y(n9580) );
  OA22XL U6985 ( .A0(n5109), .A1(n1864), .B0(n5067), .B1(n3520), .Y(n9574) );
  OA22XL U6986 ( .A0(n5292), .A1(n1865), .B0(n5245), .B1(n3521), .Y(n9572) );
  OA22XL U6987 ( .A0(n5200), .A1(n1866), .B0(n5164), .B1(n3522), .Y(n9573) );
  NAND4BX1 U6988 ( .AN(n4366), .B(n9816), .C(n9815), .D(n9814), .Y(n11211) );
  OAI22XL U6989 ( .A0(n5116), .A1(n1786), .B0(n5076), .B1(n3442), .Y(n4366) );
  NAND4BX1 U6990 ( .AN(n4367), .B(n9808), .C(n9807), .D(n9806), .Y(n11307) );
  OAI22XL U6991 ( .A0(n5116), .A1(n1787), .B0(n5060), .B1(n3443), .Y(n4367) );
  NAND4BX1 U6992 ( .AN(n4368), .B(n9796), .C(n9795), .D(n9794), .Y(n11210) );
  OAI22XL U6993 ( .A0(n5116), .A1(n1788), .B0(n5058), .B1(n3444), .Y(n4368) );
  OA22XL U6994 ( .A0(n5298), .A1(n1867), .B0(n5251), .B1(n3523), .Y(n9785) );
  NAND4BX1 U6995 ( .AN(n4369), .B(n9836), .C(n9835), .D(n9834), .Y(n11209) );
  OAI22XL U6996 ( .A0(n5117), .A1(n1789), .B0(n181), .B1(n3445), .Y(n4369) );
  NAND4BX1 U6997 ( .AN(n4370), .B(n9828), .C(n9827), .D(n9826), .Y(n11305) );
  OAI22XL U6998 ( .A0(n5117), .A1(n1790), .B0(n5069), .B1(n3446), .Y(n4370) );
  NAND4BX1 U6999 ( .AN(n4371), .B(n9872), .C(n9871), .D(n9870), .Y(n11208) );
  OAI22XL U7000 ( .A0(n5118), .A1(n1791), .B0(n5072), .B1(n3447), .Y(n4371) );
  NAND4BX1 U7001 ( .AN(n4372), .B(n9864), .C(n9863), .D(n9862), .Y(n11304) );
  OAI22XL U7002 ( .A0(n5118), .A1(n1934), .B0(n5065), .B1(n3588), .Y(n4372) );
  NAND4BX1 U7003 ( .AN(n4373), .B(n9856), .C(n9855), .D(n9854), .Y(n11207) );
  OAI22XL U7004 ( .A0(n5118), .A1(n1792), .B0(n5055), .B1(n3448), .Y(n4373) );
  NAND4BX1 U7005 ( .AN(n4374), .B(n9848), .C(n9847), .D(n9846), .Y(n11303) );
  OAI22XL U7006 ( .A0(n5117), .A1(n1793), .B0(n5084), .B1(n3449), .Y(n4374) );
  OA22XL U7007 ( .A0(n5297), .A1(n1868), .B0(n5250), .B1(n3524), .Y(n9724) );
  NAND2XL U7008 ( .A(DCACHE_addr[28]), .B(n4673), .Y(n10789) );
  NAND2XL U7009 ( .A(DCACHE_addr[29]), .B(n4673), .Y(n10137) );
  INVX1 U7010 ( .A(n10375), .Y(n10358) );
  NAND2X1 U7011 ( .A(\i_MIPS/Register/n117 ), .B(\i_MIPS/Register/n104 ), .Y(
        \i_MIPS/Register/n116 ) );
  NAND2X1 U7012 ( .A(\i_MIPS/Register/n115 ), .B(\i_MIPS/Register/n104 ), .Y(
        \i_MIPS/Register/n114 ) );
  NAND2X1 U7013 ( .A(\i_MIPS/Register/n113 ), .B(\i_MIPS/Register/n104 ), .Y(
        \i_MIPS/Register/n112 ) );
  NAND2X1 U7014 ( .A(\i_MIPS/Register/n111 ), .B(\i_MIPS/Register/n104 ), .Y(
        \i_MIPS/Register/n110 ) );
  NAND2X1 U7015 ( .A(\i_MIPS/Register/n109 ), .B(\i_MIPS/Register/n104 ), .Y(
        \i_MIPS/Register/n108 ) );
  NAND2X1 U7016 ( .A(\i_MIPS/Register/n107 ), .B(\i_MIPS/Register/n104 ), .Y(
        \i_MIPS/Register/n106 ) );
  NAND2X1 U7017 ( .A(\i_MIPS/Register/n119 ), .B(\i_MIPS/Register/n104 ), .Y(
        \i_MIPS/Register/n118 ) );
  NAND2X1 U7018 ( .A(\i_MIPS/Register/n131 ), .B(\i_MIPS/Register/n119 ), .Y(
        \i_MIPS/Register/n138 ) );
  NAND2X1 U7019 ( .A(\i_MIPS/Register/n131 ), .B(\i_MIPS/Register/n117 ), .Y(
        \i_MIPS/Register/n137 ) );
  NAND2X1 U7020 ( .A(\i_MIPS/Register/n131 ), .B(\i_MIPS/Register/n115 ), .Y(
        \i_MIPS/Register/n136 ) );
  NAND2X1 U7021 ( .A(\i_MIPS/Register/n131 ), .B(\i_MIPS/Register/n113 ), .Y(
        \i_MIPS/Register/n135 ) );
  NAND2X1 U7022 ( .A(\i_MIPS/Register/n131 ), .B(\i_MIPS/Register/n111 ), .Y(
        \i_MIPS/Register/n134 ) );
  NAND2X1 U7023 ( .A(\i_MIPS/Register/n131 ), .B(\i_MIPS/Register/n109 ), .Y(
        \i_MIPS/Register/n133 ) );
  NAND2X1 U7024 ( .A(\i_MIPS/Register/n131 ), .B(\i_MIPS/Register/n107 ), .Y(
        \i_MIPS/Register/n132 ) );
  NAND2X1 U7025 ( .A(\i_MIPS/Register/n131 ), .B(\i_MIPS/Register/n105 ), .Y(
        \i_MIPS/Register/n130 ) );
  NAND2X1 U7026 ( .A(\i_MIPS/Register/n122 ), .B(\i_MIPS/Register/n119 ), .Y(
        \i_MIPS/Register/n129 ) );
  NAND2X1 U7027 ( .A(\i_MIPS/Register/n122 ), .B(\i_MIPS/Register/n117 ), .Y(
        \i_MIPS/Register/n128 ) );
  NAND2X1 U7028 ( .A(\i_MIPS/Register/n122 ), .B(\i_MIPS/Register/n115 ), .Y(
        \i_MIPS/Register/n127 ) );
  NAND2X1 U7029 ( .A(\i_MIPS/Register/n122 ), .B(\i_MIPS/Register/n113 ), .Y(
        \i_MIPS/Register/n126 ) );
  NAND2X1 U7030 ( .A(\i_MIPS/Register/n122 ), .B(\i_MIPS/Register/n111 ), .Y(
        \i_MIPS/Register/n125 ) );
  NAND2X1 U7031 ( .A(\i_MIPS/Register/n122 ), .B(\i_MIPS/Register/n109 ), .Y(
        \i_MIPS/Register/n124 ) );
  NAND2X1 U7032 ( .A(\i_MIPS/Register/n122 ), .B(\i_MIPS/Register/n107 ), .Y(
        \i_MIPS/Register/n123 ) );
  NAND2X1 U7033 ( .A(\i_MIPS/Register/n122 ), .B(\i_MIPS/Register/n105 ), .Y(
        \i_MIPS/Register/n121 ) );
  AO21X1 U7034 ( .A0(\i_MIPS/Register/n104 ), .A1(\i_MIPS/Register/n105 ), 
        .B0(n4488), .Y(n10865) );
  NAND2XL U7035 ( .A(\i_MIPS/Control_ID/n15 ), .B(\i_MIPS/Control_ID/n10 ), 
        .Y(\i_MIPS/control_out[7] ) );
  NAND2X1 U7036 ( .A(\i_MIPS/Register/n140 ), .B(\i_MIPS/Register/n119 ), .Y(
        \i_MIPS/Register/n147 ) );
  NAND2X1 U7037 ( .A(\i_MIPS/Register/n140 ), .B(\i_MIPS/Register/n111 ), .Y(
        \i_MIPS/Register/n143 ) );
  NAND2X1 U7038 ( .A(\i_MIPS/Register/n140 ), .B(\i_MIPS/Register/n109 ), .Y(
        \i_MIPS/Register/n142 ) );
  NAND2X1 U7039 ( .A(\i_MIPS/Register/n140 ), .B(\i_MIPS/Register/n107 ), .Y(
        \i_MIPS/Register/n141 ) );
  NAND2X1 U7040 ( .A(\i_MIPS/Register/n140 ), .B(\i_MIPS/Register/n117 ), .Y(
        \i_MIPS/Register/n146 ) );
  NAND2X1 U7041 ( .A(\i_MIPS/Register/n140 ), .B(\i_MIPS/Register/n115 ), .Y(
        \i_MIPS/Register/n145 ) );
  NAND2X1 U7042 ( .A(\i_MIPS/Register/n140 ), .B(\i_MIPS/Register/n113 ), .Y(
        \i_MIPS/Register/n144 ) );
  NAND2X1 U7043 ( .A(\i_MIPS/Register/n140 ), .B(\i_MIPS/Register/n105 ), .Y(
        \i_MIPS/Register/n139 ) );
  CLKXOR2X2 U7044 ( .A(n10226), .B(ICACHE_addr[17]), .Y(n10637) );
  INVXL U7045 ( .A(n10586), .Y(n10207) );
  INVXL U7046 ( .A(n10805), .Y(n10803) );
  INVXL U7047 ( .A(n10817), .Y(n10815) );
  NAND2BX4 U7048 ( .AN(n5035), .B(\D_cache/cache[7][154] ), .Y(n6303) );
  NAND2BX4 U7049 ( .AN(n4883), .B(\D_cache/cache[3][154] ), .Y(n6307) );
  NAND2X2 U7050 ( .A(n10250), .B(ICACHE_addr[15]), .Y(n10251) );
  OA22X2 U7051 ( .A0(n5381), .A1(n1481), .B0(n5338), .B1(n3055), .Y(n9639) );
  OA22XL U7052 ( .A0(n4907), .A1(n1354), .B0(n4249), .B1(n2884), .Y(n6893) );
  OA22XL U7053 ( .A0(n4922), .A1(n1355), .B0(n4249), .B1(n2885), .Y(n7009) );
  OA22XL U7054 ( .A0(n4912), .A1(n1160), .B0(n4249), .B1(n2716), .Y(n8588) );
  INVXL U7055 ( .A(\i_MIPS/n314 ), .Y(n11174) );
  AOI2BB1XL U7056 ( .A0N(n8156), .A1N(net102253), .B0(n4518), .Y(n6692) );
  BUFX20 U7057 ( .A(n12934), .Y(DCACHE_addr[23]) );
  OA22XL U7058 ( .A0(\i_MIPS/Register/register[22][27] ), .A1(n4684), .B0(
        \i_MIPS/Register/register[30][27] ), .B1(n4678), .Y(n9422) );
  OA22XL U7059 ( .A0(\i_MIPS/Register/register[6][27] ), .A1(n4684), .B0(
        \i_MIPS/Register/register[14][27] ), .B1(n4678), .Y(n9405) );
  OA22XL U7060 ( .A0(\i_MIPS/Register/register[6][3] ), .A1(net112116), .B0(
        \i_MIPS/Register/register[14][3] ), .B1(net112134), .Y(n8371) );
  OA22XL U7061 ( .A0(\i_MIPS/Register/register[6][9] ), .A1(net112116), .B0(
        \i_MIPS/Register/register[14][9] ), .B1(net112134), .Y(n8667) );
  OA22XL U7062 ( .A0(\i_MIPS/Register/register[6][23] ), .A1(net112116), .B0(
        \i_MIPS/Register/register[14][23] ), .B1(net112134), .Y(n8832) );
  OA22XL U7063 ( .A0(\i_MIPS/Register/register[6][14] ), .A1(net112112), .B0(
        \i_MIPS/Register/register[14][14] ), .B1(net112142), .Y(n7629) );
  OA22XL U7064 ( .A0(\i_MIPS/Register/register[6][13] ), .A1(net112112), .B0(
        \i_MIPS/Register/register[14][13] ), .B1(net112132), .Y(n7722) );
  OA22XL U7065 ( .A0(\i_MIPS/Register/register[6][1] ), .A1(net112112), .B0(
        \i_MIPS/Register/register[14][1] ), .B1(net112132), .Y(n7993) );
  OA22XL U7066 ( .A0(\i_MIPS/Register/register[6][7] ), .A1(net112112), .B0(
        \i_MIPS/Register/register[14][7] ), .B1(net112132), .Y(n7914) );
  OA22XL U7067 ( .A0(\i_MIPS/Register/register[6][5] ), .A1(net112110), .B0(
        \i_MIPS/Register/register[14][5] ), .B1(net112128), .Y(n6782) );
  OA22XL U7068 ( .A0(\i_MIPS/Register/register[6][29] ), .A1(net112112), .B0(
        \i_MIPS/Register/register[14][29] ), .B1(net112132), .Y(n8134) );
  OA22XL U7069 ( .A0(\i_MIPS/Register/register[6][11] ), .A1(net112112), .B0(
        \i_MIPS/Register/register[14][11] ), .B1(net112142), .Y(n7248) );
  OA22XL U7070 ( .A0(\i_MIPS/Register/register[6][17] ), .A1(net112112), .B0(
        \i_MIPS/Register/register[14][17] ), .B1(net112132), .Y(n7781) );
  OA22XL U7071 ( .A0(\i_MIPS/Register/register[6][15] ), .A1(net112112), .B0(
        \i_MIPS/Register/register[14][15] ), .B1(net112142), .Y(n7131) );
  MXI2X1 U7072 ( .A(\i_MIPS/n345 ), .B(n4397), .S0(n214), .Y(\i_MIPS/n536 ) );
  MXI2X1 U7073 ( .A(\i_MIPS/n348 ), .B(net129017), .S0(n211), .Y(\i_MIPS/n539 ) );
  MXI2X1 U7074 ( .A(\i_MIPS/n370 ), .B(n4413), .S0(n220), .Y(\i_MIPS/n561 ) );
  MXI2X1 U7075 ( .A(\i_MIPS/n351 ), .B(n4428), .S0(n211), .Y(\i_MIPS/n542 ) );
  MXI2X1 U7076 ( .A(\i_MIPS/n349 ), .B(n4426), .S0(n204), .Y(\i_MIPS/n540 ) );
  MXI2X1 U7077 ( .A(\i_MIPS/n347 ), .B(n4410), .S0(n223), .Y(\i_MIPS/n538 ) );
  MXI2X1 U7078 ( .A(\i_MIPS/n346 ), .B(n4398), .S0(n217), .Y(\i_MIPS/n537 ) );
  OA22XL U7079 ( .A0(\i_MIPS/Register/register[22][23] ), .A1(n4683), .B0(
        \i_MIPS/Register/register[30][23] ), .B1(n4678), .Y(n8905) );
  OA22XL U7080 ( .A0(\i_MIPS/Register/register[6][25] ), .A1(n4684), .B0(
        \i_MIPS/Register/register[14][25] ), .B1(n4678), .Y(n9094) );
  OA22XL U7081 ( .A0(\i_MIPS/Register/register[6][19] ), .A1(net112116), .B0(
        \i_MIPS/Register/register[14][19] ), .B1(net112134), .Y(n8567) );
  MXI2X1 U7082 ( .A(\i_MIPS/n321 ), .B(\i_MIPS/n320 ), .S0(n211), .Y(
        \i_MIPS/n517 ) );
  MXI2X1 U7083 ( .A(\i_MIPS/n317 ), .B(\i_MIPS/n316 ), .S0(n211), .Y(
        \i_MIPS/n515 ) );
  MXI2X1 U7084 ( .A(\i_MIPS/n315 ), .B(\i_MIPS/n314 ), .S0(n217), .Y(
        \i_MIPS/n514 ) );
  MXI2X1 U7085 ( .A(\i_MIPS/n327 ), .B(\i_MIPS/n326 ), .S0(n213), .Y(
        \i_MIPS/n520 ) );
  MXI2X1 U7086 ( .A(\i_MIPS/n323 ), .B(\i_MIPS/n322 ), .S0(n210), .Y(
        \i_MIPS/n518 ) );
  NAND2XL U7087 ( .A(n10233), .B(ICACHE_addr[9]), .Y(n10234) );
  MXI2XL U7088 ( .A(n4535), .B(\i_MIPS/n225 ), .S0(n220), .Y(\i_MIPS/n502 ) );
  MXI2XL U7089 ( .A(\i_MIPS/n302 ), .B(\i_MIPS/n303 ), .S0(n223), .Y(
        \i_MIPS/n430 ) );
  MXI2XL U7090 ( .A(\i_MIPS/n300 ), .B(\i_MIPS/n301 ), .S0(n204), .Y(
        \i_MIPS/n428 ) );
  MXI2XL U7091 ( .A(\i_MIPS/n284 ), .B(\i_MIPS/n285 ), .S0(n205), .Y(
        \i_MIPS/n412 ) );
  MXI2XL U7092 ( .A(\i_MIPS/n282 ), .B(\i_MIPS/n283 ), .S0(n207), .Y(
        \i_MIPS/n410 ) );
  MXI2XL U7093 ( .A(\i_MIPS/n278 ), .B(\i_MIPS/n279 ), .S0(n204), .Y(
        \i_MIPS/n406 ) );
  MXI2XL U7094 ( .A(\i_MIPS/n276 ), .B(\i_MIPS/n277 ), .S0(n222), .Y(
        \i_MIPS/n404 ) );
  MXI2XL U7095 ( .A(\i_MIPS/n274 ), .B(\i_MIPS/n275 ), .S0(n208), .Y(
        \i_MIPS/n402 ) );
  MXI2XL U7096 ( .A(\i_MIPS/n260 ), .B(\i_MIPS/n261 ), .S0(n219), .Y(
        \i_MIPS/n388 ) );
  MXI2XL U7097 ( .A(\i_MIPS/n248 ), .B(\i_MIPS/n249 ), .S0(n220), .Y(
        \i_MIPS/n376 ) );
  MXI2XL U7098 ( .A(\i_MIPS/n246 ), .B(\i_MIPS/n247 ), .S0(n219), .Y(
        \i_MIPS/n374 ) );
  MXI2XL U7099 ( .A(\i_MIPS/n286 ), .B(\i_MIPS/n287 ), .S0(n214), .Y(
        \i_MIPS/n414 ) );
  MXI2XL U7100 ( .A(\i_MIPS/n268 ), .B(\i_MIPS/n269 ), .S0(n216), .Y(
        \i_MIPS/n396 ) );
  MXI2XL U7101 ( .A(\i_MIPS/n266 ), .B(\i_MIPS/n267 ), .S0(n214), .Y(
        \i_MIPS/n394 ) );
  MXI2XL U7102 ( .A(\i_MIPS/n250 ), .B(\i_MIPS/n251 ), .S0(n213), .Y(
        \i_MIPS/n378 ) );
  MXI2XL U7103 ( .A(\i_MIPS/n310 ), .B(\i_MIPS/n311 ), .S0(n211), .Y(
        \i_MIPS/n479 ) );
  MXI2XL U7104 ( .A(\i_MIPS/n258 ), .B(\i_MIPS/n259 ), .S0(n208), .Y(
        \i_MIPS/n386 ) );
  MXI2XL U7105 ( .A(\i_MIPS/n298 ), .B(\i_MIPS/n299 ), .S0(n208), .Y(
        \i_MIPS/n426 ) );
  MXI2XL U7106 ( .A(\i_MIPS/n270 ), .B(\i_MIPS/n271 ), .S0(n220), .Y(
        \i_MIPS/n398 ) );
  MXI2XL U7107 ( .A(\i_MIPS/n368 ), .B(n4409), .S0(n204), .Y(\i_MIPS/n559 ) );
  INVX1 U7108 ( .A(n7618), .Y(n6496) );
  AOI2BB1XL U7109 ( .A0N(n8357), .A1N(net102253), .B0(n4517), .Y(n7973) );
  OR2XL U7110 ( .A(n10176), .B(ICACHE_addr[1]), .Y(n10640) );
  OR3XL U7111 ( .A(n9891), .B(\i_MIPS/n326 ), .C(\i_MIPS/IR_ID[29] ), .Y(n9892) );
  INVXL U7112 ( .A(\i_MIPS/Control_ID/n10 ), .Y(n9614) );
  CLKMX2X2 U7113 ( .A(n3699), .B(n4613), .S0(n204), .Y(\i_MIPS/n415 ) );
  CLKMX2X2 U7114 ( .A(n3596), .B(n4623), .S0(n207), .Y(\i_MIPS/n423 ) );
  CLKMX2X2 U7115 ( .A(\i_MIPS/ID_EX[64] ), .B(n4619), .S0(n222), .Y(
        \i_MIPS/n391 ) );
  CLKMX2X2 U7116 ( .A(n3695), .B(n4627), .S0(n219), .Y(\i_MIPS/n417 ) );
  CLKMX2X2 U7117 ( .A(n10952), .B(n4617), .S0(n223), .Y(\i_MIPS/n437 ) );
  CLKMX2X2 U7118 ( .A(\i_MIPS/ID_EX[50] ), .B(n4612), .S0(n205), .Y(
        \i_MIPS/n419 ) );
  AO21X1 U7119 ( .A0(\i_MIPS/ID_EX[91] ), .A1(n202), .B0(n4380), .Y(
        \i_MIPS/n494 ) );
  AO21X1 U7120 ( .A0(\i_MIPS/ID_EX[92] ), .A1(n202), .B0(n4380), .Y(
        \i_MIPS/n493 ) );
  AO21X1 U7121 ( .A0(\i_MIPS/ID_EX[90] ), .A1(n202), .B0(n4380), .Y(
        \i_MIPS/n495 ) );
  OA22XL U7122 ( .A0(\i_MIPS/Register/register[0][22] ), .A1(n4702), .B0(
        \i_MIPS/Register/register[8][22] ), .B1(n4700), .Y(n9521) );
  OA22XL U7123 ( .A0(\i_MIPS/Register/register[4][22] ), .A1(n4697), .B0(
        \i_MIPS/Register/register[12][22] ), .B1(n4693), .Y(n9522) );
  OA22XL U7124 ( .A0(\i_MIPS/Register/register[0][21] ), .A1(n4702), .B0(
        \i_MIPS/Register/register[8][21] ), .B1(n4700), .Y(n9204) );
  OA22XL U7125 ( .A0(\i_MIPS/Register/register[4][21] ), .A1(n4697), .B0(
        \i_MIPS/Register/register[12][21] ), .B1(n4693), .Y(n9205) );
  OA22XL U7126 ( .A0(\i_MIPS/Register/register[4][8] ), .A1(n4699), .B0(
        \i_MIPS/Register/register[12][8] ), .B1(n4695), .Y(n7114) );
  OA22XL U7127 ( .A0(\i_MIPS/Register/register[0][8] ), .A1(n4704), .B0(
        \i_MIPS/Register/register[8][8] ), .B1(n4700), .Y(n7113) );
  OA22XL U7128 ( .A0(\i_MIPS/Register/register[16][21] ), .A1(n4702), .B0(
        \i_MIPS/Register/register[24][21] ), .B1(n4700), .Y(n9213) );
  OA22XL U7129 ( .A0(\i_MIPS/Register/register[20][21] ), .A1(n4697), .B0(
        \i_MIPS/Register/register[28][21] ), .B1(n4693), .Y(n9214) );
  OA22XL U7130 ( .A0(\i_MIPS/Register/register[16][19] ), .A1(n4702), .B0(
        \i_MIPS/Register/register[24][19] ), .B1(n4700), .Y(n8622) );
  OA22XL U7131 ( .A0(\i_MIPS/Register/register[20][5] ), .A1(n4698), .B0(
        \i_MIPS/Register/register[28][5] ), .B1(n4695), .Y(n6833) );
  OA22XL U7132 ( .A0(\i_MIPS/Register/register[16][5] ), .A1(n4704), .B0(
        \i_MIPS/Register/register[24][5] ), .B1(n4700), .Y(n6832) );
  OA22XL U7133 ( .A0(\i_MIPS/Register/register[20][3] ), .A1(n4698), .B0(
        \i_MIPS/Register/register[28][3] ), .B1(n4694), .Y(n8422) );
  OA22XL U7134 ( .A0(\i_MIPS/Register/register[16][3] ), .A1(n4703), .B0(
        \i_MIPS/Register/register[24][3] ), .B1(n4701), .Y(n8421) );
  OA22XL U7135 ( .A0(\i_MIPS/Register/register[20][1] ), .A1(n4698), .B0(
        \i_MIPS/Register/register[28][1] ), .B1(n4694), .Y(n8043) );
  OA22XL U7136 ( .A0(\i_MIPS/Register/register[16][1] ), .A1(n4703), .B0(
        \i_MIPS/Register/register[24][1] ), .B1(n4701), .Y(n8042) );
  OA22XL U7137 ( .A0(\i_MIPS/Register/register[20][24] ), .A1(n4698), .B0(
        \i_MIPS/Register/register[28][24] ), .B1(n4694), .Y(n8331) );
  OA22XL U7138 ( .A0(\i_MIPS/Register/register[16][24] ), .A1(n4703), .B0(
        \i_MIPS/Register/register[24][24] ), .B1(n4701), .Y(n8330) );
  OA22XL U7139 ( .A0(\i_MIPS/Register/register[20][13] ), .A1(n4699), .B0(
        \i_MIPS/Register/register[28][13] ), .B1(n4695), .Y(n7773) );
  OA22XL U7140 ( .A0(\i_MIPS/Register/register[20][14] ), .A1(n4699), .B0(
        \i_MIPS/Register/register[28][14] ), .B1(n4695), .Y(n7679) );
  OA22XL U7141 ( .A0(\i_MIPS/Register/register[16][14] ), .A1(n4703), .B0(
        \i_MIPS/Register/register[24][14] ), .B1(n4701), .Y(n7678) );
  OA22XL U7142 ( .A0(\i_MIPS/Register/register[20][29] ), .A1(n4698), .B0(
        \i_MIPS/Register/register[28][29] ), .B1(n4694), .Y(n8221) );
  OA22XL U7143 ( .A0(\i_MIPS/Register/register[16][29] ), .A1(n4703), .B0(
        \i_MIPS/Register/register[24][29] ), .B1(n4701), .Y(n8220) );
  OA22XL U7144 ( .A0(\i_MIPS/Register/register[16][8] ), .A1(n4704), .B0(
        \i_MIPS/Register/register[24][8] ), .B1(n4700), .Y(n7122) );
  OA22XL U7145 ( .A0(\i_MIPS/Register/register[20][12] ), .A1(n4699), .B0(
        \i_MIPS/Register/register[28][12] ), .B1(n4695), .Y(n7459) );
  OA22XL U7146 ( .A0(\i_MIPS/Register/register[16][12] ), .A1(n4704), .B0(
        \i_MIPS/Register/register[24][12] ), .B1(n4700), .Y(n7458) );
  OA22XL U7147 ( .A0(n4922), .A1(n1162), .B0(n4249), .B1(n2718), .Y(n7013) );
  OA22XL U7148 ( .A0(n4923), .A1(n1356), .B0(n4249), .B1(n2886), .Y(n6885) );
  OA22XL U7149 ( .A0(n4908), .A1(n1357), .B0(n4249), .B1(n2887), .Y(n6889) );
  OA22XL U7150 ( .A0(n4921), .A1(n1358), .B0(n4249), .B1(n2888), .Y(n7102) );
  OA22XL U7151 ( .A0(n4910), .A1(n1359), .B0(n4249), .B1(n2889), .Y(n6925) );
  OA22XL U7152 ( .A0(n4918), .A1(n1360), .B0(n4249), .B1(n2890), .Y(n6933) );
  OA22XL U7153 ( .A0(n4921), .A1(n1361), .B0(n4249), .B1(n2891), .Y(n7098) );
  OA22XL U7154 ( .A0(n4917), .A1(n2771), .B0(n4948), .B1(n1137), .Y(n7752) );
  AO22XL U7155 ( .A0(n4728), .A1(n927), .B0(n4725), .B1(n2634), .Y(n8028) );
  AO22XL U7156 ( .A0(net112006), .A1(n928), .B0(net112020), .B1(n2635), .Y(
        n8833) );
  AO22XL U7157 ( .A0(net112006), .A1(n929), .B0(net112020), .B1(n2636), .Y(
        n8842) );
  AO22XL U7158 ( .A0(net112006), .A1(n883), .B0(net112020), .B1(n2574), .Y(
        n8470) );
  AO22XL U7159 ( .A0(net112006), .A1(n884), .B0(net112020), .B1(n2575), .Y(
        n8668) );
  AO22XL U7160 ( .A0(net112006), .A1(n930), .B0(net112020), .B1(n2637), .Y(
        n8677) );
  AO22XL U7161 ( .A0(net112006), .A1(n885), .B0(net112020), .B1(n2576), .Y(
        n8372) );
  AO22XL U7162 ( .A0(net112006), .A1(n886), .B0(net112020), .B1(n2577), .Y(
        n8479) );
  AO22XL U7163 ( .A0(n4731), .A1(n329), .B0(n4724), .B1(n2438), .Y(n7444) );
  AO22XL U7164 ( .A0(net112006), .A1(n931), .B0(net112020), .B1(n2638), .Y(
        n8381) );
  AO22XL U7165 ( .A0(net112006), .A1(n887), .B0(net112020), .B1(n2578), .Y(
        n8281) );
  AO22XL U7166 ( .A0(net112006), .A1(n932), .B0(net112020), .B1(n2639), .Y(
        n8290) );
  AO22XL U7167 ( .A0(net112000), .A1(n933), .B0(net112018), .B1(n2640), .Y(
        n7073) );
  OA22XL U7168 ( .A0(n4903), .A1(n1132), .B0(n4949), .B1(n2668), .Y(n7277) );
  OA22XL U7169 ( .A0(n4910), .A1(n1163), .B0(n4947), .B1(n2719), .Y(n8988) );
  OA22XL U7170 ( .A0(n4910), .A1(n1363), .B0(n4947), .B1(n2893), .Y(n8980) );
  OA22XL U7171 ( .A0(n4907), .A1(n2681), .B0(n4949), .B1(n1125), .Y(n7273) );
  OA22XL U7172 ( .A0(n4921), .A1(n1364), .B0(n4949), .B1(n2894), .Y(n7183) );
  OA22XL U7173 ( .A0(n4913), .A1(n1133), .B0(n4249), .B1(n2669), .Y(n8310) );
  OA22XL U7174 ( .A0(n4912), .A1(n1366), .B0(n4249), .B1(n2896), .Y(n8500) );
  OA22XL U7175 ( .A0(n4912), .A1(n1367), .B0(n4249), .B1(n2897), .Y(n8492) );
  OA22XL U7176 ( .A0(n4912), .A1(n1368), .B0(n4249), .B1(n2898), .Y(n8496) );
  OA22XL U7177 ( .A0(n4916), .A1(n1369), .B0(n4947), .B1(n2899), .Y(n7944) );
  OA22XL U7178 ( .A0(n4917), .A1(n1119), .B0(n4249), .B1(n2655), .Y(n8693) );
  OA22XL U7179 ( .A0(n4913), .A1(n1370), .B0(n4249), .B1(n2900), .Y(n8393) );
  OA22XL U7180 ( .A0(n4914), .A1(n1371), .B0(n4249), .B1(n2901), .Y(n8306) );
  OA22XL U7181 ( .A0(n4915), .A1(n1164), .B0(n4947), .B1(n2720), .Y(n8101) );
  OA22XL U7182 ( .A0(n4916), .A1(n1372), .B0(n4947), .B1(n2902), .Y(n7936) );
  OA22XL U7183 ( .A0(n4916), .A1(n1373), .B0(n4947), .B1(n2903), .Y(n8014) );
  OA22XL U7184 ( .A0(n4914), .A1(n1134), .B0(n4947), .B1(n2670), .Y(n8200) );
  OA22XL U7185 ( .A0(n4914), .A1(n1374), .B0(n4947), .B1(n2904), .Y(n8298) );
  OA22XL U7186 ( .A0(n4916), .A1(n1375), .B0(n4947), .B1(n2905), .Y(n7940) );
  OA22XL U7187 ( .A0(n4912), .A1(n1376), .B0(n4249), .B1(n2906), .Y(n8685) );
  OA22XL U7188 ( .A0(n4916), .A1(n1377), .B0(n4947), .B1(n2907), .Y(n8010) );
  OA22XL U7189 ( .A0(n4914), .A1(n1378), .B0(n4947), .B1(n2908), .Y(n8196) );
  OA22XL U7190 ( .A0(n4915), .A1(n1379), .B0(n4947), .B1(n2909), .Y(n8189) );
  OA22XL U7191 ( .A0(n4909), .A1(n1165), .B0(n4947), .B1(n2721), .Y(n9296) );
  OA22XL U7192 ( .A0(n4909), .A1(n1380), .B0(n4947), .B1(n2910), .Y(n9383) );
  OA22XL U7193 ( .A0(n5302), .A1(n1381), .B0(n5256), .B1(n2911), .Y(n10009) );
  OA22XL U7194 ( .A0(n5303), .A1(n1382), .B0(n5258), .B1(n2912), .Y(n10104) );
  OA22XL U7195 ( .A0(n5303), .A1(n1383), .B0(n5258), .B1(n2913), .Y(n10094) );
  OA22XL U7196 ( .A0(n5298), .A1(n1166), .B0(n5251), .B1(n2722), .Y(n9776) );
  OA22XL U7197 ( .A0(n5293), .A1(n1167), .B0(n5246), .B1(n2723), .Y(n9606) );
  OA22XL U7198 ( .A0(n5298), .A1(n1168), .B0(n5251), .B1(n2724), .Y(n9771) );
  OA22XL U7199 ( .A0(n5298), .A1(n1169), .B0(n5251), .B1(n2725), .Y(n9766) );
  OA22XL U7200 ( .A0(n5303), .A1(n1384), .B0(n5257), .B1(n2914), .Y(n10028) );
  OA22XL U7201 ( .A0(n5387), .A1(n1385), .B0(n5331), .B1(n2915), .Y(n6099) );
  OA22XL U7202 ( .A0(n5386), .A1(n1386), .B0(n5329), .B1(n2916), .Y(n6052) );
  OA22XL U7203 ( .A0(n5401), .A1(n1387), .B0(n5329), .B1(n2917), .Y(n6056) );
  OA22XL U7204 ( .A0(n5383), .A1(n1708), .B0(n5354), .B1(n3305), .Y(n9894) );
  OA22XL U7205 ( .A0(n269), .A1(n1595), .B0(n5354), .B1(n3172), .Y(n9920) );
  OA22XL U7206 ( .A0(n5385), .A1(n1596), .B0(n5329), .B1(n3173), .Y(n9915) );
  OA22X2 U7207 ( .A0(n5368), .A1(n786), .B0(n5323), .B1(n2348), .Y(n5983) );
  OA22XL U7208 ( .A0(\i_MIPS/Register/register[22][28] ), .A1(n4682), .B0(
        \i_MIPS/Register/register[30][28] ), .B1(n4679), .Y(n8514) );
  OA22XL U7209 ( .A0(\i_MIPS/Register/register[22][19] ), .A1(n4682), .B0(
        \i_MIPS/Register/register[30][19] ), .B1(n4679), .Y(n8616) );
  OA22XL U7210 ( .A0(\i_MIPS/Register/register[6][29] ), .A1(n4682), .B0(
        \i_MIPS/Register/register[14][29] ), .B1(n4679), .Y(n8205) );
  OA22XL U7211 ( .A0(\i_MIPS/Register/register[6][21] ), .A1(n4684), .B0(
        \i_MIPS/Register/register[14][21] ), .B1(n4678), .Y(n9198) );
  OA22XL U7212 ( .A0(\i_MIPS/Register/register[22][21] ), .A1(n4684), .B0(
        \i_MIPS/Register/register[30][21] ), .B1(n4678), .Y(n9207) );
  OA22XL U7213 ( .A0(\i_MIPS/Register/register[6][20] ), .A1(n4684), .B0(
        \i_MIPS/Register/register[14][20] ), .B1(n4678), .Y(n9304) );
  OA22XL U7214 ( .A0(\i_MIPS/Register/register[22][20] ), .A1(n4684), .B0(
        \i_MIPS/Register/register[30][20] ), .B1(n4678), .Y(n9313) );
  OA22XL U7215 ( .A0(\i_MIPS/Register/register[22][25] ), .A1(n4684), .B0(
        \i_MIPS/Register/register[30][25] ), .B1(n4678), .Y(n9103) );
  OA22XL U7216 ( .A0(\i_MIPS/Register/register[6][22] ), .A1(n4684), .B0(
        \i_MIPS/Register/register[14][22] ), .B1(n4678), .Y(n9515) );
  OA22XL U7217 ( .A0(\i_MIPS/Register/register[22][4] ), .A1(net112110), .B0(
        \i_MIPS/Register/register[30][4] ), .B1(net112128), .Y(n6872) );
  OA22XL U7218 ( .A0(\i_MIPS/Register/register[6][4] ), .A1(net112110), .B0(
        \i_MIPS/Register/register[14][4] ), .B1(net112128), .Y(n6863) );
  OA22XL U7219 ( .A0(\i_MIPS/Register/register[22][9] ), .A1(net112116), .B0(
        \i_MIPS/Register/register[30][9] ), .B1(net112134), .Y(n8676) );
  OA22XL U7220 ( .A0(\i_MIPS/Register/register[22][23] ), .A1(net112116), .B0(
        \i_MIPS/Register/register[30][23] ), .B1(net112134), .Y(n8841) );
  OA22XL U7221 ( .A0(\i_MIPS/Register/register[22][24] ), .A1(net112116), .B0(
        \i_MIPS/Register/register[30][24] ), .B1(net112134), .Y(n8289) );
  OA22XL U7222 ( .A0(\i_MIPS/Register/register[22][3] ), .A1(net112116), .B0(
        \i_MIPS/Register/register[30][3] ), .B1(net112134), .Y(n8380) );
  OA22XL U7223 ( .A0(\i_MIPS/Register/register[22][13] ), .A1(net112112), .B0(
        \i_MIPS/Register/register[30][13] ), .B1(net112132), .Y(n7731) );
  OA22XL U7224 ( .A0(\i_MIPS/Register/register[22][1] ), .A1(net112112), .B0(
        \i_MIPS/Register/register[30][1] ), .B1(net112132), .Y(n8002) );
  OA22XL U7225 ( .A0(\i_MIPS/Register/register[22][14] ), .A1(net112112), .B0(
        \i_MIPS/Register/register[30][14] ), .B1(net112142), .Y(n7638) );
  OA22XL U7226 ( .A0(\i_MIPS/Register/register[22][7] ), .A1(net112112), .B0(
        \i_MIPS/Register/register[30][7] ), .B1(net112132), .Y(n7923) );
  OA22XL U7227 ( .A0(\i_MIPS/Register/register[22][5] ), .A1(net112110), .B0(
        \i_MIPS/Register/register[30][5] ), .B1(net112128), .Y(n6791) );
  OA22XL U7228 ( .A0(\i_MIPS/Register/register[22][19] ), .A1(net112116), .B0(
        \i_MIPS/Register/register[30][19] ), .B1(net112134), .Y(n8576) );
  OA22XL U7229 ( .A0(\i_MIPS/Register/register[22][29] ), .A1(net112112), .B0(
        \i_MIPS/Register/register[30][29] ), .B1(net112132), .Y(n8143) );
  OA22XL U7230 ( .A0(\i_MIPS/Register/register[22][11] ), .A1(net112112), .B0(
        \i_MIPS/Register/register[30][11] ), .B1(net112142), .Y(n7257) );
  OA22XL U7231 ( .A0(\i_MIPS/Register/register[22][17] ), .A1(net112112), .B0(
        \i_MIPS/Register/register[30][17] ), .B1(net112132), .Y(n7790) );
  OA22XL U7232 ( .A0(\i_MIPS/Register/register[22][15] ), .A1(net112112), .B0(
        \i_MIPS/Register/register[30][15] ), .B1(net112142), .Y(n7140) );
  OA22XL U7233 ( .A0(\i_MIPS/Register/register[22][12] ), .A1(net112112), .B0(
        \i_MIPS/Register/register[30][12] ), .B1(net112142), .Y(n7393) );
  OA22XL U7234 ( .A0(\i_MIPS/Register/register[6][12] ), .A1(net112112), .B0(
        \i_MIPS/Register/register[14][12] ), .B1(net112142), .Y(n7384) );
  OA22XL U7235 ( .A0(\i_MIPS/Register/register[6][21] ), .A1(net112116), .B0(
        \i_MIPS/Register/register[14][21] ), .B1(net112142), .Y(n9121) );
  OA22XL U7236 ( .A0(\i_MIPS/Register/register[22][21] ), .A1(net112110), .B0(
        \i_MIPS/Register/register[30][21] ), .B1(net112142), .Y(n9130) );
  OA22XL U7237 ( .A0(\i_MIPS/Register/register[22][25] ), .A1(net112110), .B0(
        \i_MIPS/Register/register[30][25] ), .B1(net112142), .Y(n9033) );
  OA22XL U7238 ( .A0(\i_MIPS/Register/register[6][25] ), .A1(net112116), .B0(
        \i_MIPS/Register/register[14][25] ), .B1(net112142), .Y(n9024) );
  OA22XL U7239 ( .A0(\i_MIPS/Register/register[22][26] ), .A1(net112116), .B0(
        \i_MIPS/Register/register[30][26] ), .B1(net112142), .Y(n8932) );
  OA22XL U7240 ( .A0(\i_MIPS/Register/register[6][26] ), .A1(net112116), .B0(
        \i_MIPS/Register/register[14][26] ), .B1(net112142), .Y(n8923) );
  OA22XL U7241 ( .A0(\i_MIPS/Register/register[22][22] ), .A1(net112116), .B0(
        \i_MIPS/Register/register[30][22] ), .B1(net112142), .Y(n9446) );
  OA22XL U7242 ( .A0(\i_MIPS/Register/register[6][22] ), .A1(net112112), .B0(
        \i_MIPS/Register/register[14][22] ), .B1(net112142), .Y(n9437) );
  OA22XL U7243 ( .A0(\i_MIPS/Register/register[6][27] ), .A1(net112112), .B0(
        \i_MIPS/Register/register[14][27] ), .B1(net112142), .Y(n9365) );
  OA22XL U7244 ( .A0(\i_MIPS/Register/register[4][11] ), .A1(n4699), .B0(
        \i_MIPS/Register/register[12][11] ), .B1(n4695), .Y(n7289) );
  OA22XL U7245 ( .A0(\i_MIPS/Register/register[4][7] ), .A1(n4698), .B0(
        \i_MIPS/Register/register[12][7] ), .B1(n4694), .Y(n7956) );
  OA22XL U7246 ( .A0(\i_MIPS/Register/register[4][10] ), .A1(n4699), .B0(
        \i_MIPS/Register/register[12][10] ), .B1(n4695), .Y(n7369) );
  OA22XL U7247 ( .A0(\i_MIPS/Register/register[4][15] ), .A1(n4699), .B0(
        \i_MIPS/Register/register[12][15] ), .B1(n4695), .Y(n7207) );
  OA22XL U7248 ( .A0(\i_MIPS/Register/register[4][4] ), .A1(n4698), .B0(
        \i_MIPS/Register/register[12][4] ), .B1(n4695), .Y(n6905) );
  OA22XL U7249 ( .A0(\i_MIPS/Register/register[0][18] ), .A1(n4702), .B0(
        \i_MIPS/Register/register[8][18] ), .B1(n4700), .Y(n8810) );
  OA22XL U7250 ( .A0(\i_MIPS/Register/register[0][25] ), .A1(n4702), .B0(
        \i_MIPS/Register/register[8][25] ), .B1(n4700), .Y(n9100) );
  OA22XL U7251 ( .A0(\i_MIPS/Register/register[0][23] ), .A1(n4702), .B0(
        \i_MIPS/Register/register[8][23] ), .B1(n4700), .Y(n8902) );
  XNOR2X4 U7252 ( .A(ICACHE_addr[26]), .B(n11341), .Y(n6072) );
  XNOR2X4 U7253 ( .A(ICACHE_addr[24]), .B(n11339), .Y(n6073) );
  XNOR2X4 U7254 ( .A(ICACHE_addr[27]), .B(n11342), .Y(n6040) );
  XNOR2X4 U7255 ( .A(ICACHE_addr[22]), .B(n11337), .Y(n6041) );
  MX2XL U7256 ( .A(\D_cache/cache[7][60] ), .B(n10480), .S0(n5000), .Y(
        \D_cache/n1309 ) );
  MX2XL U7257 ( .A(\D_cache/cache[7][54] ), .B(n10214), .S0(n5002), .Y(
        \D_cache/n1357 ) );
  MX2XL U7258 ( .A(\D_cache/cache[7][53] ), .B(n10672), .S0(n5001), .Y(
        \D_cache/n1365 ) );
  MX2XL U7259 ( .A(\D_cache/cache[7][52] ), .B(n10659), .S0(n5001), .Y(
        \D_cache/n1373 ) );
  MX2XL U7260 ( .A(\D_cache/cache[7][42] ), .B(n10262), .S0(n5002), .Y(
        \D_cache/n1453 ) );
  MX2XL U7261 ( .A(\D_cache/cache[7][38] ), .B(n10075), .S0(n5004), .Y(
        \D_cache/n1485 ) );
  MX2XL U7262 ( .A(\D_cache/cache[7][27] ), .B(n10303), .S0(n5000), .Y(
        \D_cache/n1573 ) );
  MX2XL U7263 ( .A(\D_cache/cache[7][25] ), .B(n10493), .S0(n5000), .Y(
        \D_cache/n1589 ) );
  MX2XL U7264 ( .A(\D_cache/cache[7][22] ), .B(n10211), .S0(n5007), .Y(
        \D_cache/n1613 ) );
  MX2XL U7265 ( .A(\D_cache/cache[7][18] ), .B(n10510), .S0(n5003), .Y(
        \D_cache/n1645 ) );
  MX2XL U7266 ( .A(\D_cache/cache[7][16] ), .B(n10290), .S0(n5002), .Y(
        \D_cache/n1661 ) );
  MX2XL U7267 ( .A(\D_cache/cache[7][10] ), .B(n10259), .S0(n5002), .Y(
        \D_cache/n1709 ) );
  MX2XL U7268 ( .A(\D_cache/cache[7][6] ), .B(n10069), .S0(n5000), .Y(
        \D_cache/n1741 ) );
  MX2XL U7269 ( .A(\D_cache/cache[7][3] ), .B(n9992), .S0(n5006), .Y(
        \D_cache/n1765 ) );
  MX2XL U7270 ( .A(\D_cache/cache[7][127] ), .B(n10876), .S0(n5002), .Y(
        \D_cache/n773 ) );
  MX2XL U7271 ( .A(\D_cache/cache[7][125] ), .B(n10689), .S0(n5004), .Y(
        \D_cache/n789 ) );
  MX2XL U7272 ( .A(\D_cache/cache[7][120] ), .B(n10784), .S0(n5003), .Y(
        \D_cache/n829 ) );
  MX2XL U7273 ( .A(\D_cache/cache[7][113] ), .B(n10771), .S0(n5003), .Y(
        \D_cache/n885 ) );
  MX2XL U7274 ( .A(\D_cache/cache[7][111] ), .B(n10760), .S0(n5005), .Y(
        \D_cache/n901 ) );
  MX2XL U7275 ( .A(\D_cache/cache[7][110] ), .B(n10749), .S0(n5005), .Y(
        \D_cache/n909 ) );
  MX2XL U7276 ( .A(\D_cache/cache[7][109] ), .B(n10738), .S0(n5005), .Y(
        \D_cache/n917 ) );
  MX2XL U7277 ( .A(\D_cache/cache[7][106] ), .B(n10265), .S0(n5002), .Y(
        \D_cache/n941 ) );
  MX2XL U7278 ( .A(\D_cache/cache[7][104] ), .B(n10901), .S0(n5008), .Y(
        \D_cache/n957 ) );
  MX2XL U7279 ( .A(\D_cache/cache[7][103] ), .B(n10889), .S0(n5004), .Y(
        \D_cache/n965 ) );
  MX2XL U7280 ( .A(\D_cache/cache[7][56] ), .B(n10781), .S0(n5003), .Y(
        \D_cache/n1341 ) );
  MX2XL U7281 ( .A(\D_cache/cache[7][47] ), .B(n10757), .S0(n5005), .Y(
        \D_cache/n1413 ) );
  MX2XL U7282 ( .A(\D_cache/cache[7][43] ), .B(n10712), .S0(n5004), .Y(
        \D_cache/n1445 ) );
  MX2XL U7283 ( .A(\D_cache/cache[7][41] ), .B(n10700), .S0(n5004), .Y(
        \D_cache/n1461 ) );
  MX2XL U7284 ( .A(\D_cache/cache[7][40] ), .B(n10898), .S0(n5007), .Y(
        \D_cache/n1469 ) );
  MX2XL U7285 ( .A(\D_cache/cache[7][39] ), .B(n10886), .S0(n5007), .Y(
        \D_cache/n1477 ) );
  MX2XL U7286 ( .A(\D_cache/cache[7][92] ), .B(n10486), .S0(n5000), .Y(
        \D_cache/n1053 ) );
  MX2XL U7287 ( .A(\D_cache/cache[7][91] ), .B(n10312), .S0(n5000), .Y(
        \D_cache/n1061 ) );
  MX2XL U7288 ( .A(\D_cache/cache[7][90] ), .B(n10280), .S0(n5002), .Y(
        \D_cache/n1069 ) );
  MX2XL U7289 ( .A(\D_cache/cache[7][86] ), .B(n10220), .S0(n5002), .Y(
        \D_cache/n1101 ) );
  MX2XL U7290 ( .A(\D_cache/cache[7][80] ), .B(n10299), .S0(n5001), .Y(
        \D_cache/n1149 ) );
  MX2XL U7291 ( .A(\D_cache/cache[7][74] ), .B(n10268), .S0(n5002), .Y(
        \D_cache/n1197 ) );
  MX2XL U7292 ( .A(\D_cache/cache[7][73] ), .B(n10706), .S0(n5004), .Y(
        \D_cache/n1205 ) );
  MX2XL U7293 ( .A(\D_cache/cache[7][72] ), .B(n4244), .S0(n5002), .Y(
        \D_cache/n1213 ) );
  MX2XL U7294 ( .A(\D_cache/cache[7][71] ), .B(n10892), .S0(n5004), .Y(
        \D_cache/n1221 ) );
  MX2XL U7295 ( .A(\D_cache/cache[7][29] ), .B(n10683), .S0(n5001), .Y(
        \D_cache/n1557 ) );
  MX2XL U7296 ( .A(\D_cache/cache[7][24] ), .B(n10778), .S0(n5003), .Y(
        \D_cache/n1597 ) );
  MX2XL U7297 ( .A(\D_cache/cache[7][17] ), .B(n10765), .S0(n5003), .Y(
        \D_cache/n1653 ) );
  MX2XL U7298 ( .A(\D_cache/cache[7][15] ), .B(n10754), .S0(n5005), .Y(
        \D_cache/n1669 ) );
  MX2XL U7299 ( .A(\D_cache/cache[7][12] ), .B(n10721), .S0(n5004), .Y(
        \D_cache/n1693 ) );
  MX2XL U7300 ( .A(\D_cache/cache[7][11] ), .B(n10709), .S0(n5004), .Y(
        \D_cache/n1701 ) );
  MX2XL U7301 ( .A(\D_cache/cache[7][9] ), .B(n10697), .S0(n5004), .Y(
        \D_cache/n1717 ) );
  MX2XL U7302 ( .A(\D_cache/cache[7][7] ), .B(n10883), .S0(n5003), .Y(
        \D_cache/n1733 ) );
  MX2XL U7303 ( .A(\D_cache/cache[7][36] ), .B(n10971), .S0(n5009), .Y(
        \D_cache/n1501 ) );
  MX2XL U7304 ( .A(\D_cache/cache[7][35] ), .B(n10919), .S0(n5003), .Y(
        \D_cache/n1509 ) );
  MX2XL U7305 ( .A(\D_cache/cache[7][34] ), .B(n10933), .S0(n5008), .Y(
        \D_cache/n1517 ) );
  MX2XL U7306 ( .A(\D_cache/cache[7][33] ), .B(n10910), .S0(n5007), .Y(
        \D_cache/n1525 ) );
  MX2XL U7307 ( .A(\D_cache/cache[7][2] ), .B(n10930), .S0(n5008), .Y(
        \D_cache/n1773 ) );
  MX2XL U7308 ( .A(\D_cache/cache[7][1] ), .B(n10907), .S0(n5003), .Y(
        \D_cache/n1781 ) );
  MX2XL U7309 ( .A(\D_cache/cache[7][100] ), .B(n10974), .S0(n5009), .Y(
        \D_cache/n989 ) );
  MX2XL U7310 ( .A(\D_cache/cache[7][99] ), .B(n10922), .S0(n5008), .Y(
        \D_cache/n997 ) );
  MX2XL U7311 ( .A(\D_cache/cache[7][98] ), .B(n10936), .S0(n5008), .Y(
        \D_cache/n1005 ) );
  MX2XL U7312 ( .A(\D_cache/cache[7][97] ), .B(n190), .S0(n5008), .Y(
        \D_cache/n1013 ) );
  MX2XL U7313 ( .A(\D_cache/cache[7][96] ), .B(n10961), .S0(n5000), .Y(
        \D_cache/n1021 ) );
  MX2XL U7314 ( .A(\D_cache/cache[7][68] ), .B(n10977), .S0(n5009), .Y(
        \D_cache/n1245 ) );
  MX2XL U7315 ( .A(\D_cache/cache[7][67] ), .B(n10925), .S0(n5008), .Y(
        \D_cache/n1253 ) );
  MX2XL U7316 ( .A(\D_cache/cache[7][66] ), .B(n10939), .S0(n5008), .Y(
        \D_cache/n1261 ) );
  MX2XL U7317 ( .A(\D_cache/cache[7][65] ), .B(n10916), .S0(n5003), .Y(
        \D_cache/n1269 ) );
  MX2XL U7318 ( .A(\D_cache/cache[7][37] ), .B(n10983), .S0(n5009), .Y(
        \D_cache/n1493 ) );
  MX2XL U7319 ( .A(\D_cache/cache[7][5] ), .B(n10980), .S0(n5009), .Y(
        \D_cache/n1749 ) );
  MX2XL U7320 ( .A(\D_cache/cache[7][115] ), .B(n11001), .S0(n5008), .Y(
        \D_cache/n869 ) );
  MX2XL U7321 ( .A(\D_cache/cache[7][148] ), .B(n11026), .S0(n5005), .Y(
        \D_cache/n605 ) );
  MX2XL U7322 ( .A(\D_cache/cache[7][146] ), .B(n11033), .S0(n5007), .Y(
        \D_cache/n621 ) );
  MX2XL U7323 ( .A(\D_cache/cache[7][145] ), .B(n11028), .S0(n5007), .Y(
        \D_cache/n629 ) );
  MX2XL U7324 ( .A(\D_cache/cache[7][129] ), .B(n11038), .S0(n5007), .Y(
        \D_cache/n757 ) );
  MX2XL U7325 ( .A(\D_cache/cache[7][143] ), .B(n11034), .S0(n5007), .Y(
        \D_cache/n645 ) );
  MX2XL U7326 ( .A(\D_cache/cache[7][132] ), .B(n11027), .S0(n5007), .Y(
        \D_cache/n733 ) );
  MX2XL U7327 ( .A(\D_cache/cache[7][138] ), .B(n11032), .S0(n5007), .Y(
        \D_cache/n685 ) );
  MX2XL U7328 ( .A(\D_cache/cache[7][134] ), .B(n11030), .S0(n5007), .Y(
        \D_cache/n717 ) );
  MX2XL U7329 ( .A(\D_cache/cache[7][133] ), .B(n11031), .S0(n5007), .Y(
        \D_cache/n725 ) );
  MX2XL U7330 ( .A(\D_cache/cache[7][131] ), .B(n11037), .S0(n5007), .Y(
        \D_cache/n741 ) );
  MX2XL U7331 ( .A(\D_cache/cache[7][130] ), .B(n3834), .S0(n5007), .Y(
        \D_cache/n749 ) );
  MX2XL U7332 ( .A(\D_cache/cache[7][135] ), .B(n11024), .S0(n5006), .Y(
        \D_cache/n709 ) );
  MX2XL U7333 ( .A(\D_cache/cache[7][149] ), .B(n11023), .S0(n5006), .Y(
        \D_cache/n597 ) );
  MX2XL U7334 ( .A(\D_cache/cache[7][147] ), .B(n11022), .S0(n5006), .Y(
        \D_cache/n613 ) );
  MX2XL U7335 ( .A(\D_cache/cache[7][128] ), .B(n11019), .S0(n5006), .Y(
        \D_cache/n765 ) );
  MX2XL U7336 ( .A(\D_cache/cache[7][151] ), .B(n11021), .S0(n5006), .Y(
        \D_cache/n581 ) );
  MX2XL U7337 ( .A(\D_cache/cache[7][136] ), .B(n11020), .S0(n5006), .Y(
        \D_cache/n701 ) );
  AND4X4 U7338 ( .A(n6636), .B(n6635), .C(n6634), .D(n6633), .Y(n4514) );
  OA22XL U7339 ( .A0(\i_MIPS/Register/register[6][31] ), .A1(net112110), .B0(
        \i_MIPS/Register/register[14][31] ), .B1(net112128), .Y(n6663) );
  BUFX20 U7340 ( .A(n12948), .Y(DCACHE_addr[9]) );
  OA22XL U7341 ( .A0(\i_MIPS/Register/register[6][10] ), .A1(n4683), .B0(
        \i_MIPS/Register/register[14][10] ), .B1(n4680), .Y(n7362) );
  OA22XL U7342 ( .A0(\i_MIPS/Register/register[6][11] ), .A1(n4683), .B0(
        \i_MIPS/Register/register[14][11] ), .B1(n4680), .Y(n7282) );
  OA22XL U7343 ( .A0(\i_MIPS/Register/register[6][15] ), .A1(n4683), .B0(
        \i_MIPS/Register/register[14][15] ), .B1(n4680), .Y(n7200) );
  OAI221XL U7344 ( .A0(\i_MIPS/ALUin1[7] ), .A1(net112364), .B0(
        \i_MIPS/ALUin1[6] ), .B1(net112346), .C0(n6851), .Y(n7488) );
  NAND2XL U7345 ( .A(\i_MIPS/ALUin1[30] ), .B(n6598), .Y(n6707) );
  NAND2XL U7346 ( .A(\i_MIPS/EX_MEM[6] ), .B(n4674), .Y(n10526) );
  NAND2XL U7347 ( .A(n12946), .B(\i_MIPS/n336 ), .Y(net98375) );
  NAND2XL U7348 ( .A(n12947), .B(n4673), .Y(net98371) );
  NAND2XL U7349 ( .A(\i_MIPS/EX_MEM[5] ), .B(n4673), .Y(net98366) );
  NAND2XL U7350 ( .A(n12942), .B(\i_MIPS/n336 ), .Y(net98340) );
  NAND2XL U7351 ( .A(n12941), .B(n4674), .Y(n10504) );
  NAND2XL U7352 ( .A(n12939), .B(n4674), .Y(n10565) );
  XNOR2XL U7353 ( .A(\i_MIPS/Reg_W[4] ), .B(net107810), .Y(n6638) );
  NOR2XL U7354 ( .A(n4700), .B(\i_MIPS/Register/register[8][31] ), .Y(n6723)
         );
  NOR2XL U7355 ( .A(n4702), .B(\i_MIPS/Register/register[0][31] ), .Y(n6722)
         );
  NOR2XL U7356 ( .A(n4700), .B(\i_MIPS/Register/register[24][31] ), .Y(n6736)
         );
  NOR2XL U7357 ( .A(n4702), .B(\i_MIPS/Register/register[16][31] ), .Y(n6735)
         );
  OA22XL U7358 ( .A0(\i_MIPS/Register/register[5][26] ), .A1(net112224), .B0(
        \i_MIPS/Register/register[13][26] ), .B1(net112240), .Y(n8921) );
  OA22XL U7359 ( .A0(\i_MIPS/Register/register[1][26] ), .A1(net112258), .B0(
        \i_MIPS/Register/register[9][26] ), .B1(n148), .Y(n8922) );
  OA22XL U7360 ( .A0(\i_MIPS/Register/register[7][26] ), .A1(net112152), .B0(
        \i_MIPS/Register/register[15][26] ), .B1(net112170), .Y(n8919) );
  OA22XL U7361 ( .A0(\i_MIPS/Register/register[5][29] ), .A1(net112222), .B0(
        \i_MIPS/Register/register[13][29] ), .B1(net112236), .Y(n8132) );
  OA22XL U7362 ( .A0(\i_MIPS/Register/register[1][29] ), .A1(net112254), .B0(
        \i_MIPS/Register/register[9][29] ), .B1(n148), .Y(n8133) );
  OA22XL U7363 ( .A0(\i_MIPS/Register/register[7][29] ), .A1(net112150), .B0(
        \i_MIPS/Register/register[15][29] ), .B1(net112170), .Y(n8130) );
  OA22XL U7364 ( .A0(\i_MIPS/Register/register[1][8] ), .A1(net112258), .B0(
        \i_MIPS/Register/register[9][8] ), .B1(n148), .Y(n7071) );
  OA22XL U7365 ( .A0(\i_MIPS/Register/register[7][8] ), .A1(net112152), .B0(
        \i_MIPS/Register/register[15][8] ), .B1(net112164), .Y(n7068) );
  OA22XL U7366 ( .A0(\i_MIPS/Register/register[5][12] ), .A1(net112222), .B0(
        \i_MIPS/Register/register[13][12] ), .B1(net112240), .Y(n7382) );
  OA22XL U7367 ( .A0(\i_MIPS/Register/register[7][12] ), .A1(net112148), .B0(
        \i_MIPS/Register/register[15][12] ), .B1(net112166), .Y(n7380) );
  OA22XL U7368 ( .A0(\i_MIPS/Register/register[5][15] ), .A1(n192), .B0(
        \i_MIPS/Register/register[13][15] ), .B1(net112240), .Y(n7129) );
  OA22XL U7369 ( .A0(\i_MIPS/Register/register[1][15] ), .A1(net112254), .B0(
        \i_MIPS/Register/register[9][15] ), .B1(n150), .Y(n7130) );
  OA22XL U7370 ( .A0(\i_MIPS/Register/register[7][15] ), .A1(net112152), .B0(
        \i_MIPS/Register/register[15][15] ), .B1(net112164), .Y(n7127) );
  OA22XL U7371 ( .A0(\i_MIPS/Register/register[5][1] ), .A1(net112222), .B0(
        \i_MIPS/Register/register[13][1] ), .B1(net112240), .Y(n7991) );
  OA22XL U7372 ( .A0(\i_MIPS/Register/register[1][1] ), .A1(net112254), .B0(
        \i_MIPS/Register/register[9][1] ), .B1(n147), .Y(n7992) );
  OA22XL U7373 ( .A0(\i_MIPS/Register/register[7][1] ), .A1(net112150), .B0(
        \i_MIPS/Register/register[15][1] ), .B1(net112170), .Y(n7989) );
  OA22XL U7374 ( .A0(\i_MIPS/Register/register[1][16] ), .A1(net112254), .B0(
        \i_MIPS/Register/register[9][16] ), .B1(n150), .Y(n8050) );
  OA22XL U7375 ( .A0(\i_MIPS/Register/register[5][17] ), .A1(net112222), .B0(
        \i_MIPS/Register/register[13][17] ), .B1(net112244), .Y(n7779) );
  OA22XL U7376 ( .A0(\i_MIPS/Register/register[1][17] ), .A1(net112258), .B0(
        \i_MIPS/Register/register[9][17] ), .B1(n147), .Y(n7780) );
  OA22XL U7377 ( .A0(\i_MIPS/Register/register[7][17] ), .A1(net112150), .B0(
        \i_MIPS/Register/register[15][17] ), .B1(net112170), .Y(n7777) );
  OA22XL U7378 ( .A0(\i_MIPS/Register/register[5][22] ), .A1(net112224), .B0(
        \i_MIPS/Register/register[13][22] ), .B1(net112244), .Y(n9435) );
  OA22XL U7379 ( .A0(\i_MIPS/Register/register[1][22] ), .A1(net112254), .B0(
        \i_MIPS/Register/register[9][22] ), .B1(n147), .Y(n9436) );
  OA22XL U7380 ( .A0(\i_MIPS/Register/register[7][22] ), .A1(net112148), .B0(
        \i_MIPS/Register/register[15][22] ), .B1(net112172), .Y(n9433) );
  OA22XL U7381 ( .A0(\i_MIPS/Register/register[20][30] ), .A1(n4698), .B0(
        \i_MIPS/Register/register[28][30] ), .B1(n4695), .Y(n6629) );
  OA22XL U7382 ( .A0(\i_MIPS/Register/register[16][30] ), .A1(n4704), .B0(
        \i_MIPS/Register/register[24][30] ), .B1(n4700), .Y(n6628) );
  AO22XL U7383 ( .A0(net112000), .A1(n433), .B0(net112018), .B1(n2644), .Y(
        n6664) );
  OA22XL U7384 ( .A0(\i_MIPS/Register/register[20][7] ), .A1(n4698), .B0(
        \i_MIPS/Register/register[28][7] ), .B1(n4694), .Y(n7965) );
  OA22XL U7385 ( .A0(\i_MIPS/Register/register[20][10] ), .A1(n4699), .B0(
        \i_MIPS/Register/register[28][10] ), .B1(n4695), .Y(n7378) );
  OA22XL U7386 ( .A0(\i_MIPS/Register/register[20][11] ), .A1(n4699), .B0(
        \i_MIPS/Register/register[28][11] ), .B1(n4695), .Y(n7298) );
  OA22XL U7387 ( .A0(\i_MIPS/Register/register[20][17] ), .A1(n4698), .B0(
        \i_MIPS/Register/register[28][17] ), .B1(n4694), .Y(n7871) );
  OA22XL U7388 ( .A0(\i_MIPS/Register/register[20][15] ), .A1(n4699), .B0(
        \i_MIPS/Register/register[28][15] ), .B1(n4695), .Y(n7216) );
  OA22XL U7389 ( .A0(\i_MIPS/Register/register[20][0] ), .A1(n4699), .B0(
        \i_MIPS/Register/register[28][0] ), .B1(n4695), .Y(n7607) );
  AO22XL U7390 ( .A0(net112000), .A1(n936), .B0(net112018), .B1(n2645), .Y(
        n6673) );
  AO22XL U7391 ( .A0(n4731), .A1(n349), .B0(n4726), .B1(n2579), .Y(n7292) );
  AO22XL U7392 ( .A0(n4731), .A1(n350), .B0(n4724), .B1(n2580), .Y(n7283) );
  AO22XL U7393 ( .A0(n4731), .A1(n934), .B0(n4725), .B1(n2641), .Y(n7959) );
  AO22XL U7394 ( .A0(n4731), .A1(n935), .B0(n4725), .B1(n2642), .Y(n7950) );
  AO22XL U7395 ( .A0(n4731), .A1(n330), .B0(n4727), .B1(n2439), .Y(n7372) );
  AO22XL U7396 ( .A0(n4731), .A1(n331), .B0(n4724), .B1(n2440), .Y(n7363) );
  AO22XL U7397 ( .A0(n4731), .A1(n332), .B0(n4724), .B1(n2441), .Y(n7210) );
  AO22XL U7398 ( .A0(n4731), .A1(n366), .B0(n4724), .B1(n2643), .Y(n7201) );
  AO22XL U7399 ( .A0(n4731), .A1(n351), .B0(n4724), .B1(n2581), .Y(n7592) );
  OA22XL U7400 ( .A0(\i_MIPS/Register/register[4][30] ), .A1(n4697), .B0(
        \i_MIPS/Register/register[12][30] ), .B1(n4693), .Y(n6620) );
  OA22XL U7401 ( .A0(\i_MIPS/Register/register[4][25] ), .A1(n4697), .B0(
        \i_MIPS/Register/register[12][25] ), .B1(n4693), .Y(n9101) );
  OA22XL U7402 ( .A0(\i_MIPS/Register/register[20][25] ), .A1(n4697), .B0(
        \i_MIPS/Register/register[28][25] ), .B1(n4693), .Y(n9110) );
  OA22XL U7403 ( .A0(\i_MIPS/Register/register[4][23] ), .A1(n4697), .B0(
        \i_MIPS/Register/register[12][23] ), .B1(n4693), .Y(n8903) );
  OA22XL U7404 ( .A0(\i_MIPS/Register/register[20][23] ), .A1(n4697), .B0(
        \i_MIPS/Register/register[28][23] ), .B1(n4693), .Y(n8912) );
  OA22XL U7405 ( .A0(\i_MIPS/Register/register[4][18] ), .A1(n4697), .B0(
        \i_MIPS/Register/register[12][18] ), .B1(n4693), .Y(n8811) );
  OA22XL U7406 ( .A0(\i_MIPS/Register/register[4][9] ), .A1(n4697), .B0(
        \i_MIPS/Register/register[12][9] ), .B1(n4693), .Y(n8709) );
  OA22XL U7407 ( .A0(\i_MIPS/Register/register[20][9] ), .A1(n4697), .B0(
        \i_MIPS/Register/register[28][9] ), .B1(n4693), .Y(n8718) );
  OA22XL U7408 ( .A0(\i_MIPS/Register/register[0][4] ), .A1(n4704), .B0(
        \i_MIPS/Register/register[8][4] ), .B1(n4700), .Y(n6904) );
  OA22XL U7409 ( .A0(\i_MIPS/Register/register[16][4] ), .A1(n4704), .B0(
        \i_MIPS/Register/register[24][4] ), .B1(n4700), .Y(n6913) );
  OA22XL U7410 ( .A0(\i_MIPS/Register/register[0][7] ), .A1(n4703), .B0(
        \i_MIPS/Register/register[8][7] ), .B1(n4701), .Y(n7955) );
  OA22XL U7411 ( .A0(\i_MIPS/Register/register[0][10] ), .A1(n4704), .B0(
        \i_MIPS/Register/register[8][10] ), .B1(n4700), .Y(n7368) );
  OA22XL U7412 ( .A0(\i_MIPS/Register/register[0][11] ), .A1(n4704), .B0(
        \i_MIPS/Register/register[8][11] ), .B1(n4700), .Y(n7288) );
  OA22XL U7413 ( .A0(\i_MIPS/Register/register[16][7] ), .A1(n4703), .B0(
        \i_MIPS/Register/register[24][7] ), .B1(n4701), .Y(n7964) );
  OA22XL U7414 ( .A0(\i_MIPS/Register/register[16][10] ), .A1(n4704), .B0(
        \i_MIPS/Register/register[24][10] ), .B1(n4700), .Y(n7377) );
  OA22XL U7415 ( .A0(\i_MIPS/Register/register[16][11] ), .A1(n4704), .B0(
        \i_MIPS/Register/register[24][11] ), .B1(n4700), .Y(n7297) );
  OA22XL U7416 ( .A0(\i_MIPS/Register/register[0][15] ), .A1(n4704), .B0(
        \i_MIPS/Register/register[8][15] ), .B1(n4700), .Y(n7206) );
  OA22XL U7417 ( .A0(\i_MIPS/Register/register[0][17] ), .A1(n4703), .B0(
        \i_MIPS/Register/register[8][17] ), .B1(n4701), .Y(n7861) );
  OA22XL U7418 ( .A0(\i_MIPS/Register/register[16][15] ), .A1(n4704), .B0(
        \i_MIPS/Register/register[24][15] ), .B1(n4700), .Y(n7215) );
  OA22XL U7419 ( .A0(\i_MIPS/Register/register[16][17] ), .A1(n4703), .B0(
        \i_MIPS/Register/register[24][17] ), .B1(n4701), .Y(n7870) );
  OA22XL U7420 ( .A0(\i_MIPS/Register/register[0][0] ), .A1(n4704), .B0(
        \i_MIPS/Register/register[8][0] ), .B1(n4700), .Y(n7597) );
  OA22XL U7421 ( .A0(\i_MIPS/Register/register[16][0] ), .A1(n4704), .B0(
        \i_MIPS/Register/register[24][0] ), .B1(n4700), .Y(n7606) );
  OA22XL U7422 ( .A0(\i_MIPS/Register/register[0][30] ), .A1(n4702), .B0(
        \i_MIPS/Register/register[8][30] ), .B1(n4700), .Y(n6619) );
  OA22XL U7423 ( .A0(\i_MIPS/Register/register[16][25] ), .A1(n4702), .B0(
        \i_MIPS/Register/register[24][25] ), .B1(n4700), .Y(n9109) );
  OA22XL U7424 ( .A0(\i_MIPS/Register/register[0][19] ), .A1(n4702), .B0(
        \i_MIPS/Register/register[8][19] ), .B1(n4700), .Y(n8613) );
  OA22XL U7425 ( .A0(\i_MIPS/Register/register[16][23] ), .A1(n4702), .B0(
        \i_MIPS/Register/register[24][23] ), .B1(n4700), .Y(n8911) );
  OA22XL U7426 ( .A0(\i_MIPS/Register/register[16][9] ), .A1(n4702), .B0(
        \i_MIPS/Register/register[24][9] ), .B1(n4700), .Y(n8717) );
  OA22XL U7427 ( .A0(\i_MIPS/Register/register[5][31] ), .A1(n192), .B0(
        \i_MIPS/Register/register[13][31] ), .B1(net112242), .Y(n6661) );
  OA22XL U7428 ( .A0(\i_MIPS/Register/register[1][31] ), .A1(net112260), .B0(
        \i_MIPS/Register/register[9][31] ), .B1(n150), .Y(n6662) );
  OA22XL U7429 ( .A0(\i_MIPS/Register/register[7][31] ), .A1(net112152), .B0(
        \i_MIPS/Register/register[15][31] ), .B1(net112164), .Y(n6659) );
  OA22XL U7430 ( .A0(\i_MIPS/Register/register[17][28] ), .A1(net112254), .B0(
        \i_MIPS/Register/register[25][28] ), .B1(n151), .Y(n8477) );
  OA22XL U7431 ( .A0(\i_MIPS/Register/register[17][26] ), .A1(net112258), .B0(
        \i_MIPS/Register/register[25][26] ), .B1(n151), .Y(n8931) );
  OA22XL U7432 ( .A0(\i_MIPS/Register/register[17][3] ), .A1(net112260), .B0(
        \i_MIPS/Register/register[25][3] ), .B1(n148), .Y(n8379) );
  OA22XL U7433 ( .A0(\i_MIPS/Register/register[17][8] ), .A1(net112260), .B0(
        \i_MIPS/Register/register[25][8] ), .B1(n147), .Y(n7080) );
  OA22XL U7434 ( .A0(\i_MIPS/Register/register[17][5] ), .A1(net112258), .B0(
        \i_MIPS/Register/register[25][5] ), .B1(n150), .Y(n6790) );
  OA22XL U7435 ( .A0(\i_MIPS/Register/register[17][0] ), .A1(net112254), .B0(
        \i_MIPS/Register/register[25][0] ), .B1(n151), .Y(n7564) );
  OA22XL U7436 ( .A0(\i_MIPS/Register/register[17][1] ), .A1(net112254), .B0(
        \i_MIPS/Register/register[25][1] ), .B1(n148), .Y(n8001) );
  OA22XL U7437 ( .A0(\i_MIPS/Register/register[17][7] ), .A1(net112260), .B0(
        \i_MIPS/Register/register[25][7] ), .B1(n150), .Y(n7922) );
  OA22XL U7438 ( .A0(\i_MIPS/Register/register[5][7] ), .A1(net112222), .B0(
        \i_MIPS/Register/register[13][7] ), .B1(net112242), .Y(n7912) );
  OA22XL U7439 ( .A0(\i_MIPS/Register/register[1][7] ), .A1(net112258), .B0(
        \i_MIPS/Register/register[9][7] ), .B1(n150), .Y(n7913) );
  OA22XL U7440 ( .A0(\i_MIPS/Register/register[7][7] ), .A1(net112150), .B0(
        \i_MIPS/Register/register[15][7] ), .B1(net112170), .Y(n7910) );
  OA22XL U7441 ( .A0(\i_MIPS/Register/register[17][29] ), .A1(net112254), .B0(
        \i_MIPS/Register/register[25][29] ), .B1(n147), .Y(n8142) );
  OA22XL U7442 ( .A0(\i_MIPS/Register/register[17][17] ), .A1(net112254), .B0(
        \i_MIPS/Register/register[25][17] ), .B1(n148), .Y(n7789) );
  OA22XL U7443 ( .A0(\i_MIPS/Register/register[17][31] ), .A1(net112258), .B0(
        \i_MIPS/Register/register[25][31] ), .B1(n151), .Y(n6671) );
  OA22XL U7444 ( .A0(\i_MIPS/Register/register[19][4] ), .A1(net112182), .B0(
        \i_MIPS/Register/register[27][4] ), .B1(n197), .Y(n6869) );
  OA22XL U7445 ( .A0(\i_MIPS/Register/register[3][4] ), .A1(net112182), .B0(
        \i_MIPS/Register/register[11][4] ), .B1(n200), .Y(n6860) );
  OA22XL U7446 ( .A0(\i_MIPS/Register/register[19][5] ), .A1(net112182), .B0(
        \i_MIPS/Register/register[27][5] ), .B1(n198), .Y(n6788) );
  OA22XL U7447 ( .A0(\i_MIPS/Register/register[3][5] ), .A1(net112182), .B0(
        \i_MIPS/Register/register[11][5] ), .B1(n200), .Y(n6779) );
  OA22XL U7448 ( .A0(\i_MIPS/Register/register[19][25] ), .A1(net112188), .B0(
        \i_MIPS/Register/register[27][25] ), .B1(n198), .Y(n9030) );
  OA22XL U7449 ( .A0(\i_MIPS/Register/register[3][25] ), .A1(net112188), .B0(
        \i_MIPS/Register/register[11][25] ), .B1(n199), .Y(n9021) );
  OA22XL U7450 ( .A0(\i_MIPS/Register/register[19][28] ), .A1(net112188), .B0(
        \i_MIPS/Register/register[27][28] ), .B1(n199), .Y(n8475) );
  OA22XL U7451 ( .A0(\i_MIPS/Register/register[3][28] ), .A1(net112188), .B0(
        \i_MIPS/Register/register[11][28] ), .B1(n197), .Y(n8466) );
  OA22XL U7452 ( .A0(\i_MIPS/Register/register[19][9] ), .A1(net112188), .B0(
        \i_MIPS/Register/register[27][9] ), .B1(n199), .Y(n8673) );
  OA22XL U7453 ( .A0(\i_MIPS/Register/register[3][9] ), .A1(net112188), .B0(
        \i_MIPS/Register/register[11][9] ), .B1(n198), .Y(n8664) );
  OA22XL U7454 ( .A0(\i_MIPS/Register/register[19][23] ), .A1(net112188), .B0(
        \i_MIPS/Register/register[27][23] ), .B1(n197), .Y(n8838) );
  OA22XL U7455 ( .A0(\i_MIPS/Register/register[3][23] ), .A1(net112188), .B0(
        \i_MIPS/Register/register[11][23] ), .B1(n198), .Y(n8829) );
  OA22XL U7456 ( .A0(\i_MIPS/Register/register[19][26] ), .A1(net112188), .B0(
        \i_MIPS/Register/register[27][26] ), .B1(n199), .Y(n8929) );
  OA22XL U7457 ( .A0(\i_MIPS/Register/register[19][3] ), .A1(net112188), .B0(
        \i_MIPS/Register/register[27][3] ), .B1(n198), .Y(n8377) );
  OA22XL U7458 ( .A0(\i_MIPS/Register/register[3][26] ), .A1(net112188), .B0(
        \i_MIPS/Register/register[11][26] ), .B1(n200), .Y(n8920) );
  OA22XL U7459 ( .A0(\i_MIPS/Register/register[3][3] ), .A1(net112188), .B0(
        \i_MIPS/Register/register[11][3] ), .B1(n200), .Y(n8368) );
  OA22XL U7460 ( .A0(\i_MIPS/Register/register[19][29] ), .A1(net112188), .B0(
        \i_MIPS/Register/register[27][29] ), .B1(n197), .Y(n8140) );
  OA22XL U7461 ( .A0(\i_MIPS/Register/register[3][29] ), .A1(net112188), .B0(
        \i_MIPS/Register/register[11][29] ), .B1(n198), .Y(n8131) );
  OA22XL U7462 ( .A0(\i_MIPS/Register/register[19][8] ), .A1(net112182), .B0(
        \i_MIPS/Register/register[27][8] ), .B1(n199), .Y(n7078) );
  OA22XL U7463 ( .A0(\i_MIPS/Register/register[3][8] ), .A1(net112182), .B0(
        \i_MIPS/Register/register[11][8] ), .B1(n200), .Y(n7069) );
  OA22XL U7464 ( .A0(\i_MIPS/Register/register[3][15] ), .A1(net112182), .B0(
        \i_MIPS/Register/register[11][15] ), .B1(n198), .Y(n7128) );
  OA22XL U7465 ( .A0(\i_MIPS/Register/register[19][0] ), .A1(net112188), .B0(
        \i_MIPS/Register/register[27][0] ), .B1(n198), .Y(n7562) );
  OA22XL U7466 ( .A0(\i_MIPS/Register/register[3][0] ), .A1(net112188), .B0(
        \i_MIPS/Register/register[11][0] ), .B1(n198), .Y(n7553) );
  OA22XL U7467 ( .A0(\i_MIPS/Register/register[3][13] ), .A1(net112188), .B0(
        \i_MIPS/Register/register[11][13] ), .B1(n200), .Y(n7719) );
  OA22XL U7468 ( .A0(\i_MIPS/Register/register[19][1] ), .A1(net112188), .B0(
        \i_MIPS/Register/register[27][1] ), .B1(n200), .Y(n7999) );
  OA22XL U7469 ( .A0(\i_MIPS/Register/register[3][1] ), .A1(net112188), .B0(
        \i_MIPS/Register/register[11][1] ), .B1(n199), .Y(n7990) );
  OA22XL U7470 ( .A0(\i_MIPS/Register/register[19][11] ), .A1(net112188), .B0(
        \i_MIPS/Register/register[27][11] ), .B1(n199), .Y(n7254) );
  OA22XL U7471 ( .A0(\i_MIPS/Register/register[3][11] ), .A1(net112188), .B0(
        \i_MIPS/Register/register[11][11] ), .B1(n200), .Y(n7245) );
  OA22XL U7472 ( .A0(\i_MIPS/Register/register[19][14] ), .A1(net112188), .B0(
        \i_MIPS/Register/register[27][14] ), .B1(n197), .Y(n7635) );
  OA22XL U7473 ( .A0(\i_MIPS/Register/register[3][14] ), .A1(net112188), .B0(
        \i_MIPS/Register/register[11][14] ), .B1(n199), .Y(n7626) );
  OA22XL U7474 ( .A0(\i_MIPS/Register/register[19][7] ), .A1(net112188), .B0(
        \i_MIPS/Register/register[27][7] ), .B1(n197), .Y(n7920) );
  OA22XL U7475 ( .A0(\i_MIPS/Register/register[3][7] ), .A1(net112188), .B0(
        \i_MIPS/Register/register[11][7] ), .B1(n197), .Y(n7911) );
  OA22XL U7476 ( .A0(\i_MIPS/Register/register[3][16] ), .A1(net112188), .B0(
        \i_MIPS/Register/register[11][16] ), .B1(n199), .Y(n8048) );
  OA22XL U7477 ( .A0(\i_MIPS/Register/register[19][17] ), .A1(net112182), .B0(
        \i_MIPS/Register/register[27][17] ), .B1(n200), .Y(n7787) );
  OA22XL U7478 ( .A0(\i_MIPS/Register/register[3][17] ), .A1(net112182), .B0(
        \i_MIPS/Register/register[11][17] ), .B1(n200), .Y(n7778) );
  OA22XL U7479 ( .A0(\i_MIPS/Register/register[19][15] ), .A1(net112188), .B0(
        \i_MIPS/Register/register[27][15] ), .B1(n199), .Y(n7137) );
  OA22XL U7480 ( .A0(\i_MIPS/Register/register[19][12] ), .A1(net112188), .B0(
        \i_MIPS/Register/register[27][12] ), .B1(n198), .Y(n7390) );
  OA22XL U7481 ( .A0(\i_MIPS/Register/register[3][12] ), .A1(net112188), .B0(
        \i_MIPS/Register/register[11][12] ), .B1(n197), .Y(n7381) );
  OA22XL U7482 ( .A0(\i_MIPS/Register/register[19][31] ), .A1(net112182), .B0(
        \i_MIPS/Register/register[27][31] ), .B1(n199), .Y(n6669) );
  OA22XL U7483 ( .A0(\i_MIPS/Register/register[3][31] ), .A1(net112182), .B0(
        \i_MIPS/Register/register[11][31] ), .B1(n197), .Y(n6660) );
  OA22XL U7484 ( .A0(\i_MIPS/Register/register[21][28] ), .A1(net112224), .B0(
        \i_MIPS/Register/register[29][28] ), .B1(net112240), .Y(n8476) );
  OA22XL U7485 ( .A0(\i_MIPS/Register/register[21][26] ), .A1(net112224), .B0(
        \i_MIPS/Register/register[29][26] ), .B1(net112244), .Y(n8930) );
  OA22XL U7486 ( .A0(\i_MIPS/Register/register[21][3] ), .A1(net112224), .B0(
        \i_MIPS/Register/register[29][3] ), .B1(net112242), .Y(n8378) );
  OA22XL U7487 ( .A0(\i_MIPS/Register/register[21][5] ), .A1(n192), .B0(
        \i_MIPS/Register/register[29][5] ), .B1(net112240), .Y(n6789) );
  OA22XL U7488 ( .A0(\i_MIPS/Register/register[21][0] ), .A1(net112222), .B0(
        \i_MIPS/Register/register[29][0] ), .B1(net112240), .Y(n7563) );
  OA22XL U7489 ( .A0(\i_MIPS/Register/register[21][1] ), .A1(net112222), .B0(
        \i_MIPS/Register/register[29][1] ), .B1(net112240), .Y(n8000) );
  OA22XL U7490 ( .A0(\i_MIPS/Register/register[21][7] ), .A1(net112222), .B0(
        \i_MIPS/Register/register[29][7] ), .B1(net112236), .Y(n7921) );
  OA22XL U7491 ( .A0(\i_MIPS/Register/register[21][15] ), .A1(net112222), .B0(
        \i_MIPS/Register/register[29][15] ), .B1(net112240), .Y(n7138) );
  OA22XL U7492 ( .A0(\i_MIPS/Register/register[21][29] ), .A1(net112222), .B0(
        \i_MIPS/Register/register[29][29] ), .B1(net112240), .Y(n8141) );
  OA22XL U7493 ( .A0(\i_MIPS/Register/register[21][17] ), .A1(net112222), .B0(
        \i_MIPS/Register/register[29][17] ), .B1(net112242), .Y(n7788) );
  OA22XL U7494 ( .A0(\i_MIPS/Register/register[21][12] ), .A1(net112222), .B0(
        \i_MIPS/Register/register[29][12] ), .B1(net112240), .Y(n7391) );
  OA22XL U7495 ( .A0(\i_MIPS/Register/register[21][31] ), .A1(n192), .B0(
        \i_MIPS/Register/register[29][31] ), .B1(net112240), .Y(n6670) );
  OA22XL U7496 ( .A0(\i_MIPS/Register/register[20][4] ), .A1(n4698), .B0(
        \i_MIPS/Register/register[28][4] ), .B1(n4695), .Y(n6914) );
  OA22XL U7497 ( .A0(\i_MIPS/Register/register[17][22] ), .A1(net112258), .B0(
        \i_MIPS/Register/register[25][22] ), .B1(n150), .Y(n9445) );
  OA22XL U7498 ( .A0(\i_MIPS/Register/register[1][27] ), .A1(net112260), .B0(
        \i_MIPS/Register/register[9][27] ), .B1(n151), .Y(n9364) );
  OA22XL U7499 ( .A0(\i_MIPS/Register/register[3][21] ), .A1(net112188), .B0(
        \i_MIPS/Register/register[11][21] ), .B1(n198), .Y(n9118) );
  OA22XL U7500 ( .A0(\i_MIPS/Register/register[19][22] ), .A1(net112188), .B0(
        \i_MIPS/Register/register[27][22] ), .B1(n200), .Y(n9443) );
  OA22XL U7501 ( .A0(\i_MIPS/Register/register[3][22] ), .A1(net112188), .B0(
        \i_MIPS/Register/register[11][22] ), .B1(n197), .Y(n9434) );
  OA22XL U7502 ( .A0(\i_MIPS/Register/register[21][22] ), .A1(net112224), .B0(
        \i_MIPS/Register/register[29][22] ), .B1(net112236), .Y(n9444) );
  OA22XL U7503 ( .A0(\i_MIPS/Register/register[3][27] ), .A1(net112188), .B0(
        \i_MIPS/Register/register[11][27] ), .B1(n198), .Y(n9362) );
  OA22XL U7504 ( .A0(\i_MIPS/Register/register[23][4] ), .A1(net112152), .B0(
        \i_MIPS/Register/register[31][4] ), .B1(net112164), .Y(n6868) );
  OA22XL U7505 ( .A0(\i_MIPS/Register/register[23][5] ), .A1(net112148), .B0(
        \i_MIPS/Register/register[31][5] ), .B1(net112164), .Y(n6787) );
  OA22XL U7506 ( .A0(\i_MIPS/Register/register[23][28] ), .A1(net112152), .B0(
        \i_MIPS/Register/register[31][28] ), .B1(net112170), .Y(n8474) );
  OA22XL U7507 ( .A0(\i_MIPS/Register/register[23][9] ), .A1(net112152), .B0(
        \i_MIPS/Register/register[31][9] ), .B1(net112170), .Y(n8672) );
  OA22XL U7508 ( .A0(\i_MIPS/Register/register[23][26] ), .A1(net112152), .B0(
        \i_MIPS/Register/register[31][26] ), .B1(net112170), .Y(n8928) );
  OA22XL U7509 ( .A0(\i_MIPS/Register/register[23][3] ), .A1(net112152), .B0(
        \i_MIPS/Register/register[31][3] ), .B1(net112170), .Y(n8376) );
  OA22XL U7510 ( .A0(\i_MIPS/Register/register[23][29] ), .A1(net112150), .B0(
        \i_MIPS/Register/register[31][29] ), .B1(net112170), .Y(n8139) );
  OA22XL U7511 ( .A0(\i_MIPS/Register/register[23][8] ), .A1(net112152), .B0(
        \i_MIPS/Register/register[31][8] ), .B1(net112164), .Y(n7077) );
  OA22XL U7512 ( .A0(\i_MIPS/Register/register[23][0] ), .A1(net112148), .B0(
        \i_MIPS/Register/register[31][0] ), .B1(net112166), .Y(n7561) );
  OA22XL U7513 ( .A0(\i_MIPS/Register/register[23][1] ), .A1(net112150), .B0(
        \i_MIPS/Register/register[31][1] ), .B1(net112170), .Y(n7998) );
  OA22XL U7514 ( .A0(\i_MIPS/Register/register[23][11] ), .A1(net112148), .B0(
        \i_MIPS/Register/register[31][11] ), .B1(net112166), .Y(n7253) );
  OA22XL U7515 ( .A0(\i_MIPS/Register/register[23][14] ), .A1(net112148), .B0(
        \i_MIPS/Register/register[31][14] ), .B1(net112166), .Y(n7634) );
  OA22XL U7516 ( .A0(\i_MIPS/Register/register[23][7] ), .A1(net112150), .B0(
        \i_MIPS/Register/register[31][7] ), .B1(net112170), .Y(n7919) );
  OA22XL U7517 ( .A0(\i_MIPS/Register/register[23][17] ), .A1(net112150), .B0(
        \i_MIPS/Register/register[31][17] ), .B1(net112170), .Y(n7786) );
  OA22XL U7518 ( .A0(\i_MIPS/Register/register[23][15] ), .A1(net112148), .B0(
        \i_MIPS/Register/register[31][15] ), .B1(net112166), .Y(n7136) );
  OA22XL U7519 ( .A0(\i_MIPS/Register/register[23][12] ), .A1(net112148), .B0(
        \i_MIPS/Register/register[31][12] ), .B1(net112166), .Y(n7389) );
  OA22XL U7520 ( .A0(\i_MIPS/Register/register[23][31] ), .A1(net112152), .B0(
        \i_MIPS/Register/register[31][31] ), .B1(net112164), .Y(n6668) );
  OA22XL U7521 ( .A0(n5290), .A1(n1597), .B0(n5243), .B1(n3174), .Y(n6213) );
  OA22XL U7522 ( .A0(n5290), .A1(n1598), .B0(n5243), .B1(n3175), .Y(n6203) );
  OA22XL U7523 ( .A0(n5290), .A1(n1599), .B0(n5243), .B1(n3176), .Y(n6223) );
  OA22XL U7524 ( .A0(n5290), .A1(n1600), .B0(n5243), .B1(n3177), .Y(n6198) );
  OA22XL U7525 ( .A0(n5289), .A1(n1601), .B0(n5242), .B1(n3178), .Y(n6193) );
  OA22XL U7526 ( .A0(n5289), .A1(n1602), .B0(n5242), .B1(n3179), .Y(n6188) );
  OA22XL U7527 ( .A0(n5289), .A1(n1603), .B0(n5242), .B1(n3180), .Y(n6183) );
  OA22XL U7528 ( .A0(n5291), .A1(n1604), .B0(n5244), .B1(n3181), .Y(n6241) );
  OA22XL U7529 ( .A0(n5289), .A1(n1605), .B0(n5242), .B1(n3182), .Y(n6178) );
  OA22XL U7530 ( .A0(n5291), .A1(n1606), .B0(n5244), .B1(n3183), .Y(n6249) );
  OA22XL U7531 ( .A0(n5291), .A1(n1607), .B0(n5244), .B1(n3184), .Y(n6253) );
  OA22XL U7532 ( .A0(n5291), .A1(n1608), .B0(n5244), .B1(n3185), .Y(n6245) );
  OA22XL U7533 ( .A0(\i_MIPS/Register/register[7][27] ), .A1(net112152), .B0(
        \i_MIPS/Register/register[15][27] ), .B1(net112172), .Y(n9361) );
  OA22XL U7534 ( .A0(\i_MIPS/Register/register[23][22] ), .A1(net112150), .B0(
        \i_MIPS/Register/register[31][22] ), .B1(net112172), .Y(n9442) );
  OA22X2 U7535 ( .A0(n237), .A1(n787), .B0(n5325), .B1(n2349), .Y(n6004) );
  OA22X2 U7536 ( .A0(n5396), .A1(n788), .B0(n5324), .B1(n2350), .Y(n6000) );
  OA22X2 U7537 ( .A0(n5372), .A1(n791), .B0(n5325), .B1(n2353), .Y(n6012) );
  OA22X2 U7538 ( .A0(n5396), .A1(n792), .B0(n5323), .B1(n2354), .Y(n5987) );
  OA22X2 U7539 ( .A0(n269), .A1(n794), .B0(n5327), .B1(n2356), .Y(n5973) );
  OA22XL U7540 ( .A0(\i_MIPS/Register/register[22][29] ), .A1(n4682), .B0(
        \i_MIPS/Register/register[30][29] ), .B1(n4679), .Y(n8214) );
  OA22XL U7541 ( .A0(\i_MIPS/Register/register[6][12] ), .A1(n4683), .B0(
        \i_MIPS/Register/register[14][12] ), .B1(n4680), .Y(n7443) );
  OA22XL U7542 ( .A0(\i_MIPS/Register/register[22][7] ), .A1(n4682), .B0(
        \i_MIPS/Register/register[30][7] ), .B1(n4679), .Y(n7958) );
  OA22XL U7543 ( .A0(\i_MIPS/Register/register[22][10] ), .A1(n4683), .B0(
        \i_MIPS/Register/register[30][10] ), .B1(n4680), .Y(n7371) );
  OA22XL U7544 ( .A0(\i_MIPS/Register/register[22][11] ), .A1(n4683), .B0(
        \i_MIPS/Register/register[30][11] ), .B1(n4680), .Y(n7291) );
  OA22XL U7545 ( .A0(\i_MIPS/Register/register[6][17] ), .A1(n4683), .B0(
        \i_MIPS/Register/register[14][17] ), .B1(n4680), .Y(n7855) );
  OA22XL U7546 ( .A0(\i_MIPS/Register/register[22][15] ), .A1(n4683), .B0(
        \i_MIPS/Register/register[30][15] ), .B1(n4680), .Y(n7209) );
  OA22XL U7547 ( .A0(\i_MIPS/Register/register[22][17] ), .A1(n4683), .B0(
        \i_MIPS/Register/register[30][17] ), .B1(n4680), .Y(n7864) );
  OA22XL U7548 ( .A0(\i_MIPS/Register/register[4][0] ), .A1(n4699), .B0(
        \i_MIPS/Register/register[12][0] ), .B1(n4695), .Y(n7598) );
  OA22XL U7549 ( .A0(\i_MIPS/Register/register[6][30] ), .A1(net112110), .B0(
        \i_MIPS/Register/register[14][30] ), .B1(net112128), .Y(n6459) );
  OA22XL U7550 ( .A0(\i_MIPS/Register/register[22][30] ), .A1(net112110), .B0(
        \i_MIPS/Register/register[30][30] ), .B1(net112128), .Y(n6468) );
  OA22XL U7551 ( .A0(\i_MIPS/Register/register[22][31] ), .A1(net112110), .B0(
        \i_MIPS/Register/register[30][31] ), .B1(net112128), .Y(n6672) );
  OA22XL U7552 ( .A0(\i_MIPS/Register/register[6][2] ), .A1(n4684), .B0(
        \i_MIPS/Register/register[14][2] ), .B1(n4680), .Y(n6942) );
  OA22XL U7553 ( .A0(\i_MIPS/Register/register[6][5] ), .A1(n4684), .B0(
        \i_MIPS/Register/register[14][5] ), .B1(n4680), .Y(n6817) );
  OA22XL U7554 ( .A0(\i_MIPS/Register/register[22][5] ), .A1(n4684), .B0(
        \i_MIPS/Register/register[30][5] ), .B1(n4680), .Y(n6826) );
  OA22XL U7555 ( .A0(\i_MIPS/Register/register[22][30] ), .A1(n4684), .B0(
        \i_MIPS/Register/register[30][30] ), .B1(n4680), .Y(n6622) );
  OA22XL U7556 ( .A0(\i_MIPS/Register/register[4][17] ), .A1(n4698), .B0(
        \i_MIPS/Register/register[12][17] ), .B1(n4694), .Y(n7862) );
  OA22XL U7557 ( .A0(n5390), .A1(n1388), .B0(n5329), .B1(n2918), .Y(n6064) );
  OA22XL U7558 ( .A0(n5370), .A1(n1389), .B0(n5329), .B1(n2919), .Y(n6036) );
  OA22XL U7559 ( .A0(n5396), .A1(n1390), .B0(n5330), .B1(n2920), .Y(n6068) );
  MX2XL U7560 ( .A(\D_cache/cache[7][142] ), .B(n11040), .S0(n5003), .Y(
        \D_cache/n653 ) );
  MX2XL U7561 ( .A(\I_cache/cache[5][109] ), .B(n9698), .S0(n5226), .Y(n11910)
         );
  MX2X1 U7562 ( .A(\I_cache/cache[7][107] ), .B(n9751), .S0(n5319), .Y(n11924)
         );
  MX2X1 U7563 ( .A(\I_cache/cache[5][107] ), .B(n9751), .S0(n5230), .Y(n11926)
         );
  MX2X1 U7564 ( .A(\I_cache/cache[3][107] ), .B(n9751), .S0(n5141), .Y(n11928)
         );
  MX2XL U7565 ( .A(\I_cache/cache[7][105] ), .B(n10031), .S0(n5317), .Y(n11940) );
  MX2XL U7566 ( .A(\I_cache/cache[6][105] ), .B(n10031), .S0(n5366), .Y(n11941) );
  MX2XL U7567 ( .A(\I_cache/cache[5][105] ), .B(n10031), .S0(n5228), .Y(n11942) );
  MX2XL U7568 ( .A(\I_cache/cache[4][105] ), .B(n10031), .S0(n5271), .Y(n11943) );
  MX2XL U7569 ( .A(\I_cache/cache[3][105] ), .B(n10031), .S0(n5138), .Y(n11944) );
  MX2XL U7570 ( .A(\I_cache/cache[2][105] ), .B(n10031), .S0(n5184), .Y(n11945) );
  MX2XL U7571 ( .A(\I_cache/cache[1][105] ), .B(n10031), .S0(n5048), .Y(n11946) );
  MX2XL U7572 ( .A(\I_cache/cache[0][105] ), .B(n10031), .S0(n5091), .Y(n11947) );
  MX2XL U7573 ( .A(\I_cache/cache[7][104] ), .B(n10007), .S0(n5322), .Y(n11948) );
  MX2XL U7574 ( .A(\I_cache/cache[6][104] ), .B(n10007), .S0(n5360), .Y(n11949) );
  MX2XL U7575 ( .A(\I_cache/cache[5][104] ), .B(n10007), .S0(n5228), .Y(n11950) );
  MX2XL U7576 ( .A(\I_cache/cache[4][104] ), .B(n10007), .S0(n5269), .Y(n11951) );
  MX2XL U7577 ( .A(\I_cache/cache[3][104] ), .B(n10007), .S0(n5139), .Y(n11952) );
  MX2XL U7578 ( .A(\I_cache/cache[2][104] ), .B(n10007), .S0(n5185), .Y(n11953) );
  MX2XL U7579 ( .A(\I_cache/cache[1][104] ), .B(n10007), .S0(n5045), .Y(n11954) );
  MX2XL U7580 ( .A(\I_cache/cache[0][104] ), .B(n10007), .S0(n5094), .Y(n11955) );
  MX2XL U7581 ( .A(\I_cache/cache[7][103] ), .B(n10126), .S0(n5321), .Y(n11956) );
  MX2XL U7582 ( .A(\I_cache/cache[6][103] ), .B(n10126), .S0(n5359), .Y(n11957) );
  MX2XL U7583 ( .A(\I_cache/cache[5][103] ), .B(n10126), .S0(n5228), .Y(n11958) );
  MX2XL U7584 ( .A(\I_cache/cache[4][103] ), .B(n10126), .S0(n5270), .Y(n11959) );
  MX2XL U7585 ( .A(\I_cache/cache[3][103] ), .B(n10126), .S0(n5139), .Y(n11960) );
  MX2XL U7586 ( .A(\I_cache/cache[2][103] ), .B(n10126), .S0(n5185), .Y(n11961) );
  MX2XL U7587 ( .A(\I_cache/cache[1][103] ), .B(n10126), .S0(n5045), .Y(n11962) );
  MX2XL U7588 ( .A(\I_cache/cache[0][103] ), .B(n10126), .S0(n5099), .Y(n11963) );
  MX2XL U7589 ( .A(\I_cache/cache[5][102] ), .B(n10102), .S0(n5229), .Y(n11966) );
  MX2XL U7590 ( .A(\I_cache/cache[4][102] ), .B(n10102), .S0(n5272), .Y(n11967) );
  MX2XL U7591 ( .A(\I_cache/cache[3][102] ), .B(n10102), .S0(n5140), .Y(n11968) );
  MX2XL U7592 ( .A(\I_cache/cache[2][102] ), .B(n10102), .S0(n5186), .Y(n11969) );
  MX2XL U7593 ( .A(\I_cache/cache[1][102] ), .B(n10102), .S0(n5049), .Y(n11970) );
  MX2XL U7594 ( .A(\I_cache/cache[0][102] ), .B(n10102), .S0(n5092), .Y(n11971) );
  MX2XL U7595 ( .A(\I_cache/cache[5][97] ), .B(n11074), .S0(n5232), .Y(n12006)
         );
  MX2XL U7596 ( .A(\I_cache/cache[4][97] ), .B(n11074), .S0(n5277), .Y(n12007)
         );
  MX2XL U7597 ( .A(\I_cache/cache[3][97] ), .B(n11074), .S0(n5142), .Y(n12008)
         );
  MX2XL U7598 ( .A(\I_cache/cache[2][97] ), .B(n11074), .S0(n5184), .Y(n12009)
         );
  MX2XL U7599 ( .A(\I_cache/cache[1][97] ), .B(n11074), .S0(n5045), .Y(n12010)
         );
  MX2XL U7600 ( .A(\I_cache/cache[0][97] ), .B(n11074), .S0(n5099), .Y(n12011)
         );
  MX2XL U7601 ( .A(\I_cache/cache[5][77] ), .B(n9708), .S0(n5226), .Y(n12166)
         );
  MX2X1 U7602 ( .A(\I_cache/cache[7][75] ), .B(n9756), .S0(n5319), .Y(n12180)
         );
  MX2X1 U7603 ( .A(\I_cache/cache[5][75] ), .B(n9756), .S0(n5230), .Y(n12182)
         );
  MX2X1 U7604 ( .A(\I_cache/cache[3][75] ), .B(n9756), .S0(n5141), .Y(n12184)
         );
  MX2X1 U7605 ( .A(\I_cache/cache[1][75] ), .B(n9756), .S0(n5053), .Y(n12186)
         );
  MX2XL U7606 ( .A(\I_cache/cache[5][73] ), .B(n10035), .S0(n5229), .Y(n12198)
         );
  MX2XL U7607 ( .A(\I_cache/cache[4][73] ), .B(n10035), .S0(n5272), .Y(n12199)
         );
  MX2XL U7608 ( .A(\I_cache/cache[3][73] ), .B(n10035), .S0(n5140), .Y(n12200)
         );
  MX2XL U7609 ( .A(\I_cache/cache[2][73] ), .B(n10035), .S0(n5186), .Y(n12201)
         );
  MX2XL U7610 ( .A(\I_cache/cache[1][73] ), .B(n10035), .S0(n5052), .Y(n12202)
         );
  MX2XL U7611 ( .A(\I_cache/cache[0][73] ), .B(n10035), .S0(n5098), .Y(n12203)
         );
  MX2XL U7612 ( .A(\I_cache/cache[7][72] ), .B(n10012), .S0(n5315), .Y(n12204)
         );
  MX2XL U7613 ( .A(\I_cache/cache[6][72] ), .B(n10012), .S0(n5363), .Y(n12205)
         );
  MX2XL U7614 ( .A(\I_cache/cache[5][72] ), .B(n10012), .S0(n5228), .Y(n12206)
         );
  MX2XL U7615 ( .A(\I_cache/cache[4][72] ), .B(n10012), .S0(n5277), .Y(n12207)
         );
  MX2XL U7616 ( .A(\I_cache/cache[3][72] ), .B(n10012), .S0(n5139), .Y(n12208)
         );
  MX2XL U7617 ( .A(\I_cache/cache[2][72] ), .B(n10012), .S0(n5185), .Y(n12209)
         );
  MX2XL U7618 ( .A(\I_cache/cache[1][72] ), .B(n10012), .S0(n5045), .Y(n12210)
         );
  MX2XL U7619 ( .A(\I_cache/cache[0][72] ), .B(n10012), .S0(n5094), .Y(n12211)
         );
  MX2XL U7620 ( .A(\I_cache/cache[7][71] ), .B(n10131), .S0(n5322), .Y(n12212)
         );
  MX2XL U7621 ( .A(\I_cache/cache[6][71] ), .B(n10131), .S0(n5362), .Y(n12213)
         );
  MX2XL U7622 ( .A(\I_cache/cache[5][71] ), .B(n10131), .S0(n5228), .Y(n12214)
         );
  MX2XL U7623 ( .A(\I_cache/cache[4][71] ), .B(n10131), .S0(n5272), .Y(n12215)
         );
  MX2XL U7624 ( .A(\I_cache/cache[3][71] ), .B(n10131), .S0(n5139), .Y(n12216)
         );
  MX2XL U7625 ( .A(\I_cache/cache[2][71] ), .B(n10131), .S0(n5185), .Y(n12217)
         );
  MX2XL U7626 ( .A(\I_cache/cache[1][71] ), .B(n10131), .S0(n5046), .Y(n12218)
         );
  MX2XL U7627 ( .A(\I_cache/cache[0][71] ), .B(n10131), .S0(n5099), .Y(n12219)
         );
  MX2XL U7628 ( .A(\I_cache/cache[5][70] ), .B(n10107), .S0(n5229), .Y(n12222)
         );
  MX2XL U7629 ( .A(\I_cache/cache[4][70] ), .B(n10107), .S0(n5272), .Y(n12223)
         );
  MX2XL U7630 ( .A(\I_cache/cache[3][70] ), .B(n10107), .S0(n5140), .Y(n12224)
         );
  MX2XL U7631 ( .A(\I_cache/cache[2][70] ), .B(n10107), .S0(n5186), .Y(n12225)
         );
  MX2XL U7632 ( .A(\I_cache/cache[1][70] ), .B(n10107), .S0(n5052), .Y(n12226)
         );
  MX2XL U7633 ( .A(\I_cache/cache[0][70] ), .B(n10107), .S0(n5093), .Y(n12227)
         );
  MX2XL U7634 ( .A(\I_cache/cache[5][65] ), .B(n11075), .S0(n5229), .Y(n12262)
         );
  MX2XL U7635 ( .A(\I_cache/cache[4][65] ), .B(n11075), .S0(n5277), .Y(n12263)
         );
  MX2XL U7636 ( .A(\I_cache/cache[3][65] ), .B(n11075), .S0(n5137), .Y(n12264)
         );
  MX2XL U7637 ( .A(\I_cache/cache[2][65] ), .B(n11075), .S0(n5188), .Y(n12265)
         );
  MX2XL U7638 ( .A(\I_cache/cache[1][65] ), .B(n11075), .S0(n5046), .Y(n12266)
         );
  MX2XL U7639 ( .A(\I_cache/cache[0][65] ), .B(n11075), .S0(n5099), .Y(n12267)
         );
  MX2XL U7640 ( .A(\I_cache/cache[5][45] ), .B(n9703), .S0(n5226), .Y(n12422)
         );
  MX2X1 U7641 ( .A(\I_cache/cache[7][43] ), .B(n9746), .S0(n5319), .Y(n12436)
         );
  MX2X1 U7642 ( .A(\I_cache/cache[5][43] ), .B(n9746), .S0(n5230), .Y(n12438)
         );
  MX2X1 U7643 ( .A(\I_cache/cache[5][42] ), .B(n10049), .S0(n5229), .Y(n12446)
         );
  MX2X1 U7644 ( .A(\I_cache/cache[3][42] ), .B(n10049), .S0(n5140), .Y(n12448)
         );
  MX2X1 U7645 ( .A(\I_cache/cache[1][42] ), .B(n10049), .S0(n5053), .Y(n12450)
         );
  MX2XL U7646 ( .A(\I_cache/cache[7][41] ), .B(n10026), .S0(n5317), .Y(n12452)
         );
  MX2XL U7647 ( .A(\I_cache/cache[6][41] ), .B(n10026), .S0(n5359), .Y(n12453)
         );
  MX2XL U7648 ( .A(\I_cache/cache[5][41] ), .B(n10026), .S0(n5226), .Y(n12454)
         );
  MX2XL U7649 ( .A(\I_cache/cache[4][41] ), .B(n10026), .S0(n5271), .Y(n12455)
         );
  MX2XL U7650 ( .A(\I_cache/cache[3][41] ), .B(n10026), .S0(n5138), .Y(n12456)
         );
  MX2XL U7651 ( .A(\I_cache/cache[2][41] ), .B(n10026), .S0(n5184), .Y(n12457)
         );
  MX2XL U7652 ( .A(\I_cache/cache[1][41] ), .B(n10026), .S0(n5049), .Y(n12458)
         );
  MX2XL U7653 ( .A(\I_cache/cache[0][41] ), .B(n10026), .S0(n5091), .Y(n12459)
         );
  MX2XL U7654 ( .A(\I_cache/cache[7][40] ), .B(n10002), .S0(n5316), .Y(n12460)
         );
  MX2XL U7655 ( .A(\I_cache/cache[6][40] ), .B(n10002), .S0(n5361), .Y(n12461)
         );
  MX2XL U7656 ( .A(\I_cache/cache[5][40] ), .B(n10002), .S0(n5228), .Y(n12462)
         );
  MX2XL U7657 ( .A(\I_cache/cache[4][40] ), .B(n10002), .S0(n5271), .Y(n12463)
         );
  MX2XL U7658 ( .A(\I_cache/cache[3][40] ), .B(n10002), .S0(n5139), .Y(n12464)
         );
  MX2XL U7659 ( .A(\I_cache/cache[2][40] ), .B(n10002), .S0(n5185), .Y(n12465)
         );
  MX2XL U7660 ( .A(\I_cache/cache[1][40] ), .B(n10002), .S0(n5046), .Y(n12466)
         );
  MX2XL U7661 ( .A(\I_cache/cache[0][40] ), .B(n10002), .S0(n5099), .Y(n12467)
         );
  MX2XL U7662 ( .A(\I_cache/cache[5][39] ), .B(n10121), .S0(n5229), .Y(n12470)
         );
  MX2XL U7663 ( .A(\I_cache/cache[4][39] ), .B(n10121), .S0(n5272), .Y(n12471)
         );
  MX2XL U7664 ( .A(\I_cache/cache[3][39] ), .B(n10121), .S0(n5140), .Y(n12472)
         );
  MX2XL U7665 ( .A(\I_cache/cache[2][39] ), .B(n10121), .S0(n5186), .Y(n12473)
         );
  MX2XL U7666 ( .A(\I_cache/cache[1][39] ), .B(n10121), .S0(n5052), .Y(n12474)
         );
  MX2XL U7667 ( .A(\I_cache/cache[0][39] ), .B(n10121), .S0(n5098), .Y(n12475)
         );
  MX2XL U7668 ( .A(\I_cache/cache[5][38] ), .B(n10097), .S0(n5229), .Y(n12478)
         );
  MX2XL U7669 ( .A(\I_cache/cache[4][38] ), .B(n10097), .S0(n5272), .Y(n12479)
         );
  MX2XL U7670 ( .A(\I_cache/cache[3][38] ), .B(n10097), .S0(n5140), .Y(n12480)
         );
  MX2XL U7671 ( .A(\I_cache/cache[2][38] ), .B(n10097), .S0(n5186), .Y(n12481)
         );
  MX2XL U7672 ( .A(\I_cache/cache[1][38] ), .B(n10097), .S0(n5048), .Y(n12482)
         );
  MX2XL U7673 ( .A(\I_cache/cache[0][38] ), .B(n10097), .S0(n5092), .Y(n12483)
         );
  MX2XL U7674 ( .A(\I_cache/cache[2][33] ), .B(n11073), .S0(n5189), .Y(n12521)
         );
  MX2X1 U7675 ( .A(\I_cache/cache[7][11] ), .B(n9741), .S0(n5315), .Y(n12692)
         );
  MX2X1 U7676 ( .A(\I_cache/cache[5][11] ), .B(n9741), .S0(n5226), .Y(n12694)
         );
  MX2X1 U7677 ( .A(\I_cache/cache[3][11] ), .B(n9741), .S0(n5136), .Y(n12696)
         );
  MX2X1 U7678 ( .A(\I_cache/cache[1][11] ), .B(n9741), .S0(n5049), .Y(n12698)
         );
  MX2XL U7679 ( .A(\I_cache/cache[5][10] ), .B(n10044), .S0(n5229), .Y(n12702)
         );
  MX2XL U7680 ( .A(\I_cache/cache[3][10] ), .B(n10044), .S0(n5140), .Y(n12704)
         );
  MX2XL U7681 ( .A(\I_cache/cache[7][9] ), .B(n10021), .S0(n5318), .Y(n12708)
         );
  MX2XL U7682 ( .A(\I_cache/cache[6][9] ), .B(n10021), .S0(n5362), .Y(n12709)
         );
  MX2XL U7683 ( .A(\I_cache/cache[5][9] ), .B(n10021), .S0(n5228), .Y(n12710)
         );
  MX2XL U7684 ( .A(\I_cache/cache[4][9] ), .B(n10021), .S0(n5276), .Y(n12711)
         );
  MX2XL U7685 ( .A(\I_cache/cache[3][9] ), .B(n10021), .S0(n5139), .Y(n12712)
         );
  MX2XL U7686 ( .A(\I_cache/cache[2][9] ), .B(n10021), .S0(n5185), .Y(n12713)
         );
  MX2XL U7687 ( .A(\I_cache/cache[1][9] ), .B(n10021), .S0(n5051), .Y(n12714)
         );
  MX2XL U7688 ( .A(\I_cache/cache[0][9] ), .B(n10021), .S0(n5094), .Y(n12715)
         );
  MX2XL U7689 ( .A(\I_cache/cache[7][8] ), .B(n9997), .S0(n5320), .Y(n12716)
         );
  MX2XL U7690 ( .A(\I_cache/cache[6][8] ), .B(n9997), .S0(n5364), .Y(n12717)
         );
  MX2XL U7691 ( .A(\I_cache/cache[5][8] ), .B(n9997), .S0(n5228), .Y(n12718)
         );
  MX2XL U7692 ( .A(\I_cache/cache[4][8] ), .B(n9997), .S0(n5269), .Y(n12719)
         );
  MX2XL U7693 ( .A(\I_cache/cache[3][8] ), .B(n9997), .S0(n5139), .Y(n12720)
         );
  MX2XL U7694 ( .A(\I_cache/cache[2][8] ), .B(n9997), .S0(n5185), .Y(n12721)
         );
  MX2XL U7695 ( .A(\I_cache/cache[1][8] ), .B(n9997), .S0(n5048), .Y(n12722)
         );
  MX2XL U7696 ( .A(\I_cache/cache[5][7] ), .B(n10116), .S0(n5229), .Y(n12726)
         );
  MX2XL U7697 ( .A(\I_cache/cache[4][7] ), .B(n10116), .S0(n5272), .Y(n12727)
         );
  MX2XL U7698 ( .A(\I_cache/cache[3][7] ), .B(n10116), .S0(n5140), .Y(n12728)
         );
  MX2XL U7699 ( .A(\I_cache/cache[2][7] ), .B(n10116), .S0(n5186), .Y(n12729)
         );
  MX2XL U7700 ( .A(\I_cache/cache[1][7] ), .B(n10116), .S0(n5052), .Y(n12730)
         );
  MX2XL U7701 ( .A(\I_cache/cache[0][7] ), .B(n10116), .S0(n5093), .Y(n12731)
         );
  MX2XL U7702 ( .A(\I_cache/cache[5][6] ), .B(n10092), .S0(n5229), .Y(n12734)
         );
  MX2XL U7703 ( .A(\I_cache/cache[4][6] ), .B(n10092), .S0(n5272), .Y(n12735)
         );
  MX2XL U7704 ( .A(\I_cache/cache[3][6] ), .B(n10092), .S0(n5140), .Y(n12736)
         );
  MX2XL U7705 ( .A(\I_cache/cache[2][6] ), .B(n10092), .S0(n5186), .Y(n12737)
         );
  MX2XL U7706 ( .A(\I_cache/cache[1][6] ), .B(n10092), .S0(n5048), .Y(n12738)
         );
  MX2XL U7707 ( .A(\I_cache/cache[0][6] ), .B(n10092), .S0(n5094), .Y(n12739)
         );
  MX2XL U7708 ( .A(\I_cache/cache[2][15] ), .B(n9643), .S0(n5181), .Y(n12665)
         );
  MX2XL U7709 ( .A(\I_cache/cache[1][15] ), .B(n9643), .S0(n5047), .Y(n12666)
         );
  MX2XL U7710 ( .A(\I_cache/cache[0][15] ), .B(n9643), .S0(n5091), .Y(n12667)
         );
  MX2XL U7711 ( .A(\I_cache/cache[3][111] ), .B(n9648), .S0(n5135), .Y(n11896)
         );
  MX2XL U7712 ( .A(\I_cache/cache[2][111] ), .B(n9648), .S0(n5181), .Y(n11897)
         );
  MX2XL U7713 ( .A(\I_cache/cache[1][111] ), .B(n9648), .S0(n5046), .Y(n11898)
         );
  MX2XL U7714 ( .A(\I_cache/cache[0][111] ), .B(n9648), .S0(n5099), .Y(n11899)
         );
  MX2XL U7715 ( .A(\I_cache/cache[3][47] ), .B(n9653), .S0(n5135), .Y(n12408)
         );
  MX2XL U7716 ( .A(\I_cache/cache[2][47] ), .B(n9653), .S0(n5181), .Y(n12409)
         );
  MX2XL U7717 ( .A(\I_cache/cache[1][47] ), .B(n9653), .S0(n5049), .Y(n12410)
         );
  MX2XL U7718 ( .A(\I_cache/cache[0][47] ), .B(n9653), .S0(n5092), .Y(n12411)
         );
  MX2XL U7719 ( .A(\I_cache/cache[7][96] ), .B(n6151), .S0(n5316), .Y(n12012)
         );
  MX2XL U7720 ( .A(\I_cache/cache[6][96] ), .B(n6151), .S0(n5364), .Y(n12013)
         );
  MX2XL U7721 ( .A(\I_cache/cache[5][96] ), .B(n6151), .S0(n5227), .Y(n12014)
         );
  MX2XL U7722 ( .A(\I_cache/cache[4][96] ), .B(n6151), .S0(n5270), .Y(n12015)
         );
  MX2XL U7723 ( .A(\I_cache/cache[3][96] ), .B(n6151), .S0(n5137), .Y(n12016)
         );
  MX2XL U7724 ( .A(\I_cache/cache[2][96] ), .B(n6151), .S0(n5183), .Y(n12017)
         );
  MX2XL U7725 ( .A(\I_cache/cache[1][96] ), .B(n6151), .S0(n5047), .Y(n12018)
         );
  MX2XL U7726 ( .A(\I_cache/cache[0][96] ), .B(n6151), .S0(n5093), .Y(n12019)
         );
  MX2XL U7727 ( .A(\I_cache/cache[7][64] ), .B(n6156), .S0(n5316), .Y(n12268)
         );
  MX2XL U7728 ( .A(\I_cache/cache[6][64] ), .B(n6156), .S0(n5358), .Y(n12269)
         );
  MX2XL U7729 ( .A(\I_cache/cache[5][64] ), .B(n6156), .S0(n5227), .Y(n12270)
         );
  MX2XL U7730 ( .A(\I_cache/cache[4][64] ), .B(n6156), .S0(n5270), .Y(n12271)
         );
  MX2XL U7731 ( .A(\I_cache/cache[3][64] ), .B(n6156), .S0(n5137), .Y(n12272)
         );
  MX2XL U7732 ( .A(\I_cache/cache[2][64] ), .B(n6156), .S0(n5183), .Y(n12273)
         );
  MX2XL U7733 ( .A(\I_cache/cache[1][64] ), .B(n6156), .S0(n5047), .Y(n12274)
         );
  MX2XL U7734 ( .A(\I_cache/cache[0][64] ), .B(n6156), .S0(n5093), .Y(n12275)
         );
  MX2XL U7735 ( .A(\I_cache/cache[7][32] ), .B(n6146), .S0(n5316), .Y(n12524)
         );
  MX2XL U7736 ( .A(\I_cache/cache[6][32] ), .B(n6146), .S0(n5360), .Y(n12525)
         );
  MX2XL U7737 ( .A(\I_cache/cache[5][32] ), .B(n6146), .S0(n5227), .Y(n12526)
         );
  MX2XL U7738 ( .A(\I_cache/cache[4][32] ), .B(n6146), .S0(n5270), .Y(n12527)
         );
  MX2XL U7739 ( .A(\I_cache/cache[3][32] ), .B(n6146), .S0(n5137), .Y(n12528)
         );
  MX2XL U7740 ( .A(\I_cache/cache[2][32] ), .B(n6146), .S0(n5183), .Y(n12529)
         );
  MX2XL U7741 ( .A(\I_cache/cache[1][32] ), .B(n6146), .S0(n5049), .Y(n12530)
         );
  MX2XL U7742 ( .A(\I_cache/cache[0][32] ), .B(n6146), .S0(n5093), .Y(n12531)
         );
  MX2XL U7743 ( .A(\I_cache/cache[5][4] ), .B(n6131), .S0(n5232), .Y(n12750)
         );
  MX2XL U7744 ( .A(\I_cache/cache[4][4] ), .B(n6131), .S0(n5275), .Y(n12751)
         );
  MX2XL U7745 ( .A(\I_cache/cache[3][4] ), .B(n6131), .S0(n5139), .Y(n12752)
         );
  MX2XL U7746 ( .A(\I_cache/cache[2][4] ), .B(n6131), .S0(n5181), .Y(n12753)
         );
  MX2XL U7747 ( .A(\I_cache/cache[1][4] ), .B(n6131), .S0(n5049), .Y(n12754)
         );
  MX2XL U7748 ( .A(\I_cache/cache[0][4] ), .B(n6131), .S0(n5093), .Y(n12755)
         );
  MX2XL U7749 ( .A(\I_cache/cache[7][1] ), .B(n6136), .S0(n5316), .Y(n12772)
         );
  MX2XL U7750 ( .A(\I_cache/cache[6][1] ), .B(n6136), .S0(n5359), .Y(n12773)
         );
  MX2XL U7751 ( .A(\I_cache/cache[5][1] ), .B(n6136), .S0(n5227), .Y(n12774)
         );
  MX2XL U7752 ( .A(\I_cache/cache[4][1] ), .B(n6136), .S0(n5270), .Y(n12775)
         );
  MX2XL U7753 ( .A(\I_cache/cache[3][1] ), .B(n6136), .S0(n5137), .Y(n12776)
         );
  MX2XL U7754 ( .A(\I_cache/cache[2][1] ), .B(n6136), .S0(n5183), .Y(n12777)
         );
  MX2XL U7755 ( .A(\I_cache/cache[1][1] ), .B(n6136), .S0(n5053), .Y(n12778)
         );
  MX2XL U7756 ( .A(\I_cache/cache[0][1] ), .B(n6136), .S0(n5093), .Y(n12779)
         );
  MX2XL U7757 ( .A(\I_cache/cache[7][0] ), .B(n6141), .S0(n5316), .Y(n12787)
         );
  MX2XL U7758 ( .A(\I_cache/cache[6][0] ), .B(n6141), .S0(n5358), .Y(n12780)
         );
  MX2XL U7759 ( .A(\I_cache/cache[5][0] ), .B(n6141), .S0(n5227), .Y(n12781)
         );
  MX2XL U7760 ( .A(\I_cache/cache[4][0] ), .B(n6141), .S0(n5270), .Y(n12782)
         );
  MX2XL U7761 ( .A(\I_cache/cache[3][0] ), .B(n6141), .S0(n5137), .Y(n12783)
         );
  MX2XL U7762 ( .A(\I_cache/cache[2][0] ), .B(n6141), .S0(n5183), .Y(n12784)
         );
  MX2XL U7763 ( .A(\I_cache/cache[1][0] ), .B(n6141), .S0(n5047), .Y(n12785)
         );
  MX2XL U7764 ( .A(\I_cache/cache[0][0] ), .B(n6141), .S0(n5093), .Y(n12786)
         );
  MX2XL U7765 ( .A(\I_cache/cache[7][67] ), .B(n11172), .S0(n5314), .Y(n12244)
         );
  MX2XL U7766 ( .A(\I_cache/cache[6][67] ), .B(n11172), .S0(n5366), .Y(n12245)
         );
  MX2XL U7767 ( .A(\I_cache/cache[5][67] ), .B(n11172), .S0(n5228), .Y(n12246)
         );
  MX2XL U7768 ( .A(\I_cache/cache[4][67] ), .B(n11172), .S0(n5270), .Y(n12247)
         );
  MX2XL U7769 ( .A(\I_cache/cache[3][67] ), .B(n11172), .S0(n5139), .Y(n12248)
         );
  MX2XL U7770 ( .A(\I_cache/cache[2][67] ), .B(n11172), .S0(n5185), .Y(n12249)
         );
  MX2XL U7771 ( .A(\I_cache/cache[1][67] ), .B(n11172), .S0(n5047), .Y(n12250)
         );
  MX2XL U7772 ( .A(\I_cache/cache[5][35] ), .B(n11168), .S0(n5233), .Y(n12502)
         );
  MX2XL U7773 ( .A(\I_cache/cache[4][35] ), .B(n11168), .S0(n5276), .Y(n12503)
         );
  MX2XL U7774 ( .A(\I_cache/cache[3][35] ), .B(n11168), .S0(n5143), .Y(n12504)
         );
  MX2XL U7775 ( .A(\I_cache/cache[1][35] ), .B(n11168), .S0(n5045), .Y(n12506)
         );
  MX2XL U7776 ( .A(\I_cache/cache[5][3] ), .B(n11167), .S0(n5233), .Y(n12758)
         );
  MX2XL U7777 ( .A(\I_cache/cache[3][3] ), .B(n11167), .S0(n5143), .Y(n12760)
         );
  MX2XL U7778 ( .A(\I_cache/cache[1][3] ), .B(n11167), .S0(n5049), .Y(n12762)
         );
  MX2XL U7779 ( .A(\I_cache/cache[5][144] ), .B(n11154), .S0(n5233), .Y(n11630) );
  MX2XL U7780 ( .A(\I_cache/cache[4][144] ), .B(n11154), .S0(n5276), .Y(n11631) );
  MX2XL U7781 ( .A(\I_cache/cache[3][144] ), .B(n11154), .S0(n5143), .Y(n11632) );
  MX2XL U7782 ( .A(\I_cache/cache[2][144] ), .B(n11154), .S0(n5189), .Y(n11633) );
  MX2XL U7783 ( .A(\I_cache/cache[1][144] ), .B(n11154), .S0(n5045), .Y(n11634) );
  MX2XL U7784 ( .A(\I_cache/cache[0][144] ), .B(n11154), .S0(n5098), .Y(n11635) );
  MX2XL U7785 ( .A(\I_cache/cache[5][151] ), .B(n11150), .S0(n5231), .Y(n11574) );
  MX2XL U7786 ( .A(\I_cache/cache[4][151] ), .B(n11150), .S0(n5274), .Y(n11575) );
  MX2XL U7787 ( .A(\I_cache/cache[3][151] ), .B(n11150), .S0(n5142), .Y(n11576) );
  MX2XL U7788 ( .A(\I_cache/cache[2][151] ), .B(n11150), .S0(n5188), .Y(n11577) );
  MX2XL U7789 ( .A(\I_cache/cache[1][151] ), .B(n11150), .S0(n5053), .Y(n11578) );
  MX2XL U7790 ( .A(\I_cache/cache[0][151] ), .B(n11150), .S0(n5096), .Y(n11579) );
  MX2XL U7791 ( .A(\I_cache/cache[5][150] ), .B(n11138), .S0(n5232), .Y(n11582) );
  MX2XL U7792 ( .A(\I_cache/cache[4][150] ), .B(n11138), .S0(n5275), .Y(n11583) );
  MX2XL U7793 ( .A(\I_cache/cache[3][150] ), .B(n11138), .S0(n5141), .Y(n11584) );
  MX2XL U7794 ( .A(\I_cache/cache[2][150] ), .B(n11138), .S0(n5185), .Y(n11585) );
  MX2XL U7795 ( .A(\I_cache/cache[1][150] ), .B(n11138), .S0(n5053), .Y(n11586) );
  MX2XL U7796 ( .A(\I_cache/cache[0][150] ), .B(n11138), .S0(n5097), .Y(n11587) );
  MX2XL U7797 ( .A(\I_cache/cache[5][149] ), .B(n11144), .S0(n5232), .Y(n11590) );
  MX2XL U7798 ( .A(\I_cache/cache[4][149] ), .B(n11144), .S0(n5275), .Y(n11591) );
  MX2XL U7799 ( .A(\I_cache/cache[3][149] ), .B(n11144), .S0(n5143), .Y(n11592) );
  MX2XL U7800 ( .A(\I_cache/cache[2][149] ), .B(n11144), .S0(n5184), .Y(n11593) );
  MX2XL U7801 ( .A(\I_cache/cache[1][149] ), .B(n11144), .S0(n5048), .Y(n11594) );
  MX2XL U7802 ( .A(\I_cache/cache[0][149] ), .B(n11144), .S0(n5097), .Y(n11595) );
  MX2XL U7803 ( .A(\I_cache/cache[5][148] ), .B(n11146), .S0(n5232), .Y(n11598) );
  MX2XL U7804 ( .A(\I_cache/cache[4][148] ), .B(n11146), .S0(n5275), .Y(n11599) );
  MX2XL U7805 ( .A(\I_cache/cache[3][148] ), .B(n11146), .S0(n5138), .Y(n11600) );
  MX2XL U7806 ( .A(\I_cache/cache[2][148] ), .B(n11146), .S0(n5188), .Y(n11601) );
  MX2XL U7807 ( .A(\I_cache/cache[1][148] ), .B(n11146), .S0(n5045), .Y(n11602) );
  MX2XL U7808 ( .A(\I_cache/cache[0][148] ), .B(n11146), .S0(n5097), .Y(n11603) );
  MX2XL U7809 ( .A(\I_cache/cache[5][147] ), .B(n11145), .S0(n5232), .Y(n11606) );
  MX2XL U7810 ( .A(\I_cache/cache[4][147] ), .B(n11145), .S0(n5275), .Y(n11607) );
  MX2XL U7811 ( .A(\I_cache/cache[3][147] ), .B(n11145), .S0(n5136), .Y(n11608) );
  MX2XL U7812 ( .A(\I_cache/cache[2][147] ), .B(n11145), .S0(n5181), .Y(n11609) );
  MX2XL U7813 ( .A(\I_cache/cache[1][147] ), .B(n11145), .S0(n5052), .Y(n11610) );
  MX2XL U7814 ( .A(\I_cache/cache[0][147] ), .B(n11145), .S0(n5097), .Y(n11611) );
  MX2XL U7815 ( .A(\I_cache/cache[5][146] ), .B(n11137), .S0(n5226), .Y(n11614) );
  MX2XL U7816 ( .A(\I_cache/cache[4][146] ), .B(n11137), .S0(n5277), .Y(n11615) );
  MX2XL U7817 ( .A(\I_cache/cache[3][146] ), .B(n11137), .S0(n5137), .Y(n11616) );
  MX2XL U7818 ( .A(\I_cache/cache[2][146] ), .B(n11137), .S0(n5187), .Y(n11617) );
  MX2XL U7819 ( .A(\I_cache/cache[1][146] ), .B(n11137), .S0(n5051), .Y(n11618) );
  MX2XL U7820 ( .A(\I_cache/cache[0][146] ), .B(n11137), .S0(n5099), .Y(n11619) );
  MX2XL U7821 ( .A(\I_cache/cache[5][145] ), .B(n11139), .S0(n5232), .Y(n11622) );
  MX2XL U7822 ( .A(\I_cache/cache[4][145] ), .B(n11139), .S0(n5275), .Y(n11623) );
  MX2XL U7823 ( .A(\I_cache/cache[3][145] ), .B(n11139), .S0(n5135), .Y(n11624) );
  MX2XL U7824 ( .A(\I_cache/cache[2][145] ), .B(n11139), .S0(n5185), .Y(n11625) );
  MX2XL U7825 ( .A(\I_cache/cache[1][145] ), .B(n11139), .S0(n5046), .Y(n11626) );
  MX2XL U7826 ( .A(\I_cache/cache[0][145] ), .B(n11139), .S0(n5097), .Y(n11627) );
  MX2XL U7827 ( .A(\I_cache/cache[5][139] ), .B(n11153), .S0(n5233), .Y(n11670) );
  MX2XL U7828 ( .A(\I_cache/cache[4][139] ), .B(n11153), .S0(n5276), .Y(n11671) );
  MX2XL U7829 ( .A(\I_cache/cache[3][139] ), .B(n11153), .S0(n5143), .Y(n11672) );
  MX2XL U7830 ( .A(\I_cache/cache[2][139] ), .B(n11153), .S0(n5189), .Y(n11673) );
  MX2XL U7831 ( .A(\I_cache/cache[1][139] ), .B(n11153), .S0(n5050), .Y(n11674) );
  MX2XL U7832 ( .A(\I_cache/cache[0][139] ), .B(n11153), .S0(n5098), .Y(n11675) );
  MX2XL U7833 ( .A(\I_cache/cache[5][138] ), .B(n11140), .S0(n5232), .Y(n11678) );
  MX2XL U7834 ( .A(\I_cache/cache[4][138] ), .B(n11140), .S0(n5275), .Y(n11679) );
  MX2XL U7835 ( .A(\I_cache/cache[3][138] ), .B(n11140), .S0(n5139), .Y(n11680) );
  MX2XL U7836 ( .A(\I_cache/cache[2][138] ), .B(n11140), .S0(n5183), .Y(n11681) );
  MX2XL U7837 ( .A(\I_cache/cache[1][138] ), .B(n11140), .S0(n5046), .Y(n11682) );
  MX2XL U7838 ( .A(\I_cache/cache[0][138] ), .B(n11140), .S0(n5097), .Y(n11683) );
  MX2XL U7839 ( .A(\I_cache/cache[5][137] ), .B(n11147), .S0(n5232), .Y(n11686) );
  MX2XL U7840 ( .A(\I_cache/cache[4][137] ), .B(n11147), .S0(n5275), .Y(n11687) );
  MX2XL U7841 ( .A(\I_cache/cache[3][137] ), .B(n11147), .S0(n5137), .Y(n11688) );
  MX2XL U7842 ( .A(\I_cache/cache[2][137] ), .B(n11147), .S0(n5184), .Y(n11689) );
  MX2XL U7843 ( .A(\I_cache/cache[1][137] ), .B(n11147), .S0(n5047), .Y(n11690) );
  MX2XL U7844 ( .A(\I_cache/cache[0][137] ), .B(n11147), .S0(n5097), .Y(n11691) );
  MX2XL U7845 ( .A(\I_cache/cache[5][136] ), .B(n11149), .S0(n5232), .Y(n11694) );
  MX2XL U7846 ( .A(\I_cache/cache[4][136] ), .B(n11149), .S0(n5275), .Y(n11695) );
  MX2XL U7847 ( .A(\I_cache/cache[3][136] ), .B(n11149), .S0(n5141), .Y(n11696) );
  MX2XL U7848 ( .A(\I_cache/cache[2][136] ), .B(n11149), .S0(n5186), .Y(n11697) );
  MX2XL U7849 ( .A(\I_cache/cache[1][136] ), .B(n11149), .S0(n5047), .Y(n11698) );
  MX2XL U7850 ( .A(\I_cache/cache[0][136] ), .B(n11149), .S0(n5097), .Y(n11699) );
  MX2XL U7851 ( .A(\I_cache/cache[5][135] ), .B(n11148), .S0(n5232), .Y(n11702) );
  MX2XL U7852 ( .A(\I_cache/cache[4][135] ), .B(n11148), .S0(n5275), .Y(n11703) );
  MX2XL U7853 ( .A(\I_cache/cache[3][135] ), .B(n11148), .S0(n5140), .Y(n11704) );
  MX2XL U7854 ( .A(\I_cache/cache[2][135] ), .B(n11148), .S0(n5188), .Y(n11705) );
  MX2XL U7855 ( .A(\I_cache/cache[1][135] ), .B(n11148), .S0(n5050), .Y(n11706) );
  MX2XL U7856 ( .A(\I_cache/cache[0][135] ), .B(n11148), .S0(n5097), .Y(n11707) );
  MX2XL U7857 ( .A(\I_cache/cache[5][134] ), .B(n11142), .S0(n5232), .Y(n11710) );
  MX2XL U7858 ( .A(\I_cache/cache[4][134] ), .B(n11142), .S0(n5275), .Y(n11711) );
  MX2XL U7859 ( .A(\I_cache/cache[3][134] ), .B(n11142), .S0(n5143), .Y(n11712) );
  MX2XL U7860 ( .A(\I_cache/cache[2][134] ), .B(n11142), .S0(n5187), .Y(n11713) );
  MX2XL U7861 ( .A(\I_cache/cache[1][134] ), .B(n11142), .S0(n5053), .Y(n11714) );
  MX2XL U7862 ( .A(\I_cache/cache[0][134] ), .B(n11142), .S0(n5097), .Y(n11715) );
  MX2XL U7863 ( .A(\I_cache/cache[5][133] ), .B(n11141), .S0(n5232), .Y(n11718) );
  MX2XL U7864 ( .A(\I_cache/cache[4][133] ), .B(n11141), .S0(n5275), .Y(n11719) );
  MX2XL U7865 ( .A(\I_cache/cache[3][133] ), .B(n11141), .S0(n5142), .Y(n11720) );
  MX2XL U7866 ( .A(\I_cache/cache[2][133] ), .B(n11141), .S0(n5189), .Y(n11721) );
  MX2XL U7867 ( .A(\I_cache/cache[1][133] ), .B(n11141), .S0(n5045), .Y(n11722) );
  MX2XL U7868 ( .A(\I_cache/cache[0][133] ), .B(n11141), .S0(n5097), .Y(n11723) );
  MX2XL U7869 ( .A(\I_cache/cache[5][132] ), .B(n11143), .S0(n5232), .Y(n11726) );
  MX2XL U7870 ( .A(\I_cache/cache[4][132] ), .B(n11143), .S0(n5275), .Y(n11727) );
  MX2XL U7871 ( .A(\I_cache/cache[3][132] ), .B(n11143), .S0(n5141), .Y(n11728) );
  MX2XL U7872 ( .A(\I_cache/cache[2][132] ), .B(n11143), .S0(n5185), .Y(n11729) );
  MX2XL U7873 ( .A(\I_cache/cache[1][132] ), .B(n11143), .S0(n5047), .Y(n11730) );
  MX2XL U7874 ( .A(\I_cache/cache[0][132] ), .B(n11143), .S0(n5097), .Y(n11731) );
  MX2XL U7875 ( .A(\I_cache/cache[5][128] ), .B(n11151), .S0(n5233), .Y(n11758) );
  MX2XL U7876 ( .A(\I_cache/cache[4][128] ), .B(n11151), .S0(n5276), .Y(n11759) );
  MX2XL U7877 ( .A(\I_cache/cache[3][128] ), .B(n11151), .S0(n5143), .Y(n11760) );
  MX2XL U7878 ( .A(\I_cache/cache[2][128] ), .B(n11151), .S0(n5189), .Y(n11761) );
  MX2XL U7879 ( .A(\I_cache/cache[1][128] ), .B(n11151), .S0(n5050), .Y(n11762) );
  MX2XL U7880 ( .A(\I_cache/cache[0][128] ), .B(n11151), .S0(n5098), .Y(n11763) );
  MX2XL U7881 ( .A(\I_cache/cache[5][140] ), .B(n11156), .S0(n5233), .Y(n11662) );
  MX2XL U7882 ( .A(\I_cache/cache[4][140] ), .B(n11156), .S0(n5276), .Y(n11663) );
  MX2XL U7883 ( .A(\I_cache/cache[3][140] ), .B(n11156), .S0(n5143), .Y(n11664) );
  MX2XL U7884 ( .A(\I_cache/cache[2][140] ), .B(n11156), .S0(n5189), .Y(n11665) );
  MX2XL U7885 ( .A(\I_cache/cache[1][140] ), .B(n11156), .S0(n5047), .Y(n11666) );
  MX2XL U7886 ( .A(\I_cache/cache[0][140] ), .B(n11156), .S0(n5098), .Y(n11667) );
  MX2XL U7887 ( .A(\I_cache/cache[7][102] ), .B(n10102), .S0(n5318), .Y(n11964) );
  MX2XL U7888 ( .A(\I_cache/cache[6][102] ), .B(n10102), .S0(n5363), .Y(n11965) );
  MX2XL U7889 ( .A(\I_cache/cache[7][97] ), .B(n11074), .S0(n5322), .Y(n12004)
         );
  MX2XL U7890 ( .A(\I_cache/cache[6][97] ), .B(n11074), .S0(n5359), .Y(n12005)
         );
  MX2XL U7891 ( .A(\I_cache/cache[7][73] ), .B(n10035), .S0(n5318), .Y(n12196)
         );
  MX2XL U7892 ( .A(\I_cache/cache[6][73] ), .B(n10035), .S0(n5366), .Y(n12197)
         );
  MX2XL U7893 ( .A(\I_cache/cache[7][70] ), .B(n10107), .S0(n5318), .Y(n12220)
         );
  MX2XL U7894 ( .A(\I_cache/cache[6][70] ), .B(n10107), .S0(n5359), .Y(n12221)
         );
  MX2XL U7895 ( .A(\I_cache/cache[7][65] ), .B(n11075), .S0(n5322), .Y(n12260)
         );
  MX2XL U7896 ( .A(\I_cache/cache[6][65] ), .B(n11075), .S0(n5363), .Y(n12261)
         );
  MX2X1 U7897 ( .A(\I_cache/cache[7][42] ), .B(n10049), .S0(n5318), .Y(n12444)
         );
  MX2XL U7898 ( .A(\I_cache/cache[7][39] ), .B(n10121), .S0(n5318), .Y(n12468)
         );
  MX2XL U7899 ( .A(\I_cache/cache[6][39] ), .B(n10121), .S0(n5360), .Y(n12469)
         );
  MX2XL U7900 ( .A(\I_cache/cache[7][38] ), .B(n10097), .S0(n5318), .Y(n12476)
         );
  MX2XL U7901 ( .A(\I_cache/cache[6][38] ), .B(n10097), .S0(n5359), .Y(n12477)
         );
  MX2XL U7902 ( .A(\I_cache/cache[7][33] ), .B(n11073), .S0(n5322), .Y(n12516)
         );
  MX2XL U7903 ( .A(\I_cache/cache[7][10] ), .B(n10044), .S0(n5318), .Y(n12700)
         );
  MX2XL U7904 ( .A(\I_cache/cache[7][7] ), .B(n10116), .S0(n5318), .Y(n12724)
         );
  MX2XL U7905 ( .A(\I_cache/cache[6][7] ), .B(n10116), .S0(n5366), .Y(n12725)
         );
  MX2XL U7906 ( .A(\I_cache/cache[7][6] ), .B(n10092), .S0(n5318), .Y(n12732)
         );
  MX2XL U7907 ( .A(\I_cache/cache[6][6] ), .B(n10092), .S0(n5361), .Y(n12733)
         );
  MX2XL U7908 ( .A(\I_cache/cache[6][15] ), .B(n9643), .S0(n5363), .Y(n12661)
         );
  MX2XL U7909 ( .A(\I_cache/cache[5][15] ), .B(n9643), .S0(n5225), .Y(n12662)
         );
  MX2XL U7910 ( .A(\I_cache/cache[4][15] ), .B(n9643), .S0(n5276), .Y(n12663)
         );
  MX2XL U7911 ( .A(\I_cache/cache[6][111] ), .B(n9648), .S0(n5361), .Y(n11893)
         );
  MX2XL U7912 ( .A(\I_cache/cache[5][47] ), .B(n9653), .S0(n5225), .Y(n12406)
         );
  MX2XL U7913 ( .A(\I_cache/cache[4][47] ), .B(n9653), .S0(n5269), .Y(n12407)
         );
  MX2XL U7914 ( .A(\I_cache/cache[7][111] ), .B(n9648), .S0(n5314), .Y(n11892)
         );
  MX2XL U7915 ( .A(\I_cache/cache[7][35] ), .B(n11168), .S0(n5321), .Y(n12500)
         );
  MX2XL U7916 ( .A(\I_cache/cache[7][3] ), .B(n11167), .S0(n5321), .Y(n12756)
         );
  MX2XL U7917 ( .A(\I_cache/cache[5][142] ), .B(n11131), .S0(n5230), .Y(n11646) );
  MX2XL U7918 ( .A(\I_cache/cache[4][142] ), .B(n11131), .S0(n5275), .Y(n11647) );
  MX2XL U7919 ( .A(\I_cache/cache[3][142] ), .B(n11131), .S0(n5137), .Y(n11648) );
  MX2XL U7920 ( .A(\I_cache/cache[2][142] ), .B(n11131), .S0(n5182), .Y(n11649) );
  MX2XL U7921 ( .A(\I_cache/cache[1][142] ), .B(n11131), .S0(n5048), .Y(n11650) );
  MX2XL U7922 ( .A(\I_cache/cache[0][142] ), .B(n11131), .S0(n5097), .Y(n11651) );
  MX2XL U7923 ( .A(\I_cache/cache[5][143] ), .B(n11133), .S0(n5229), .Y(n11638) );
  MX2XL U7924 ( .A(\I_cache/cache[4][143] ), .B(n11133), .S0(n5275), .Y(n11639) );
  MX2XL U7925 ( .A(\I_cache/cache[3][143] ), .B(n11133), .S0(n5139), .Y(n11640) );
  MX2XL U7926 ( .A(\I_cache/cache[2][143] ), .B(n11133), .S0(n5182), .Y(n11641) );
  MX2XL U7927 ( .A(\I_cache/cache[1][143] ), .B(n11133), .S0(n5051), .Y(n11642) );
  MX2XL U7928 ( .A(\I_cache/cache[0][143] ), .B(n11133), .S0(n5099), .Y(n11643) );
  MX2XL U7929 ( .A(\I_cache/cache[5][141] ), .B(n11132), .S0(n5230), .Y(n11654) );
  MX2XL U7930 ( .A(\I_cache/cache[4][141] ), .B(n11132), .S0(n5277), .Y(n11655) );
  MX2XL U7931 ( .A(\I_cache/cache[3][141] ), .B(n11132), .S0(n5136), .Y(n11656) );
  MX2XL U7932 ( .A(\I_cache/cache[2][141] ), .B(n11132), .S0(n5183), .Y(n11657) );
  MX2XL U7933 ( .A(\I_cache/cache[1][141] ), .B(n11132), .S0(n5052), .Y(n11658) );
  MX2XL U7934 ( .A(\I_cache/cache[0][141] ), .B(n11132), .S0(n5097), .Y(n11659) );
  MX2XL U7935 ( .A(\I_cache/cache[5][131] ), .B(n11135), .S0(n5229), .Y(n11734) );
  MX2XL U7936 ( .A(\I_cache/cache[4][131] ), .B(n11135), .S0(n5276), .Y(n11735) );
  MX2XL U7937 ( .A(\I_cache/cache[3][131] ), .B(n11135), .S0(n5138), .Y(n11736) );
  MX2XL U7938 ( .A(\I_cache/cache[2][131] ), .B(n11135), .S0(n5182), .Y(n11737) );
  MX2XL U7939 ( .A(\I_cache/cache[1][131] ), .B(n11135), .S0(n5049), .Y(n11738) );
  MX2XL U7940 ( .A(\I_cache/cache[0][131] ), .B(n11135), .S0(n5098), .Y(n11739) );
  MX2XL U7941 ( .A(\I_cache/cache[5][130] ), .B(n11136), .S0(n5232), .Y(n11742) );
  MX2XL U7942 ( .A(\I_cache/cache[4][130] ), .B(n11136), .S0(n5275), .Y(n11743) );
  MX2XL U7943 ( .A(\I_cache/cache[3][130] ), .B(n11136), .S0(n5135), .Y(n11744) );
  MX2XL U7944 ( .A(\I_cache/cache[2][130] ), .B(n11136), .S0(n5181), .Y(n11745) );
  MX2XL U7945 ( .A(\I_cache/cache[1][130] ), .B(n11136), .S0(n5048), .Y(n11746) );
  MX2XL U7946 ( .A(\I_cache/cache[0][130] ), .B(n11136), .S0(n5099), .Y(n11747) );
  MX2XL U7947 ( .A(\I_cache/cache[5][129] ), .B(n11134), .S0(n5230), .Y(n11750) );
  MX2XL U7948 ( .A(\I_cache/cache[4][129] ), .B(n11134), .S0(n5277), .Y(n11751) );
  MX2XL U7949 ( .A(\I_cache/cache[3][129] ), .B(n11134), .S0(n5141), .Y(n11752) );
  MX2XL U7950 ( .A(\I_cache/cache[2][129] ), .B(n11134), .S0(n5185), .Y(n11753) );
  MX2XL U7951 ( .A(\I_cache/cache[1][129] ), .B(n11134), .S0(n5049), .Y(n11754) );
  MX2XL U7952 ( .A(\I_cache/cache[0][129] ), .B(n11134), .S0(n5097), .Y(n11755) );
  MX2XL U7953 ( .A(\D_cache/cache[6][142] ), .B(n11040), .S0(n4959), .Y(
        \D_cache/n654 ) );
  MX2XL U7954 ( .A(\D_cache/cache[3][142] ), .B(n11040), .S0(n4849), .Y(
        \D_cache/n657 ) );
  MX2XL U7955 ( .A(\D_cache/cache[2][142] ), .B(n11040), .S0(n4805), .Y(
        \D_cache/n658 ) );
  MX2XL U7956 ( .A(\D_cache/cache[1][142] ), .B(n11040), .S0(n4782), .Y(
        \D_cache/n659 ) );
  MX2XL U7957 ( .A(\D_cache/cache[0][142] ), .B(n11040), .S0(n4736), .Y(
        \D_cache/n660 ) );
  MX2XL U7958 ( .A(\I_cache/cache[7][4] ), .B(n6131), .S0(n5320), .Y(n12748)
         );
  MX2XL U7959 ( .A(\I_cache/cache[6][4] ), .B(n6131), .S0(n5366), .Y(n12749)
         );
  XOR2XL U7960 ( .A(n11067), .B(n4301), .Y(n11068) );
  OA22XL U7961 ( .A0(n5392), .A1(n1869), .B0(n5336), .B1(n3525), .Y(n9571) );
  OA22XL U7962 ( .A0(n5396), .A1(n1870), .B0(n5336), .B1(n3526), .Y(n9575) );
  AO21XL U7963 ( .A0(n3431), .A1(n5009), .B0(\D_cache/cache[7][154] ), .Y(
        \D_cache/n557 ) );
  AO21XL U7964 ( .A0(n3431), .A1(n4965), .B0(\D_cache/cache[6][154] ), .Y(
        \D_cache/n558 ) );
  AO21XL U7965 ( .A0(n3431), .A1(n4944), .B0(\D_cache/cache[5][154] ), .Y(
        \D_cache/n559 ) );
  AO21XL U7966 ( .A0(n3431), .A1(n4901), .B0(\D_cache/cache[4][154] ), .Y(
        \D_cache/n560 ) );
  AO21XL U7967 ( .A0(n3431), .A1(n4855), .B0(\D_cache/cache[3][154] ), .Y(
        \D_cache/n561 ) );
  AO21XL U7968 ( .A0(n3431), .A1(n4809), .B0(\D_cache/cache[2][154] ), .Y(
        \D_cache/n562 ) );
  AO21XL U7969 ( .A0(n3431), .A1(n4786), .B0(\D_cache/cache[1][154] ), .Y(
        \D_cache/n563 ) );
  AO21XL U7970 ( .A0(n3431), .A1(n4735), .B0(\D_cache/cache[0][154] ), .Y(
        \D_cache/n564 ) );
  MX2X1 U7971 ( .A(\I_cache/cache[0][153] ), .B(n414), .S0(n5097), .Y(n11563)
         );
  MX2X1 U7972 ( .A(\I_cache/cache[5][153] ), .B(n414), .S0(n5229), .Y(n11558)
         );
  MX2X1 U7973 ( .A(\I_cache/cache[4][153] ), .B(n414), .S0(n5273), .Y(n11559)
         );
  MX2X1 U7974 ( .A(\I_cache/cache[3][153] ), .B(n414), .S0(n5137), .Y(n11560)
         );
  MX2X1 U7975 ( .A(\I_cache/cache[2][153] ), .B(n414), .S0(n5187), .Y(n11561)
         );
  MX2X1 U7976 ( .A(\I_cache/cache[1][153] ), .B(n414), .S0(n5051), .Y(n11562)
         );
  MX2X1 U7977 ( .A(\I_cache/cache[7][153] ), .B(n414), .S0(n5319), .Y(n11556)
         );
  MX2X1 U7978 ( .A(\I_cache/cache[6][153] ), .B(n414), .S0(n5365), .Y(n11557)
         );
  AOI2BB1XL U7979 ( .A0N(\i_MIPS/n322 ), .A1N(\i_MIPS/n332 ), .B0(
        \i_MIPS/IR_ID[30] ), .Y(n9889) );
  XOR2XL U7980 ( .A(n9888), .B(n9887), .Y(n9890) );
  NAND2XL U7981 ( .A(\i_MIPS/IR_ID[31] ), .B(n4487), .Y(
        \i_MIPS/Control_ID/n12 ) );
  BUFX20 U7982 ( .A(n3915), .Y(n5545) );
  OA22X4 U7983 ( .A0(n4925), .A1(n2188), .B0(n4955), .B1(n614), .Y(n6390) );
  OA22X4 U7984 ( .A0(n4925), .A1(n2189), .B0(n4955), .B1(n615), .Y(n6394) );
  INVX3 U7985 ( .A(net108150), .Y(net108098) );
  CLKBUFX3 U7986 ( .A(n5524), .Y(n5514) );
  CLKBUFX3 U7987 ( .A(n5524), .Y(n5521) );
  CLKBUFX3 U7988 ( .A(n10864), .Y(n5465) );
  CLKBUFX3 U7989 ( .A(n10864), .Y(n5466) );
  INVX3 U7990 ( .A(n4791), .Y(n4778) );
  INVX3 U7991 ( .A(n4791), .Y(n4779) );
  INVX3 U7992 ( .A(n5116), .Y(n5097) );
  INVX3 U7993 ( .A(n5192), .Y(n5188) );
  INVX3 U7994 ( .A(n5116), .Y(n5096) );
  INVX3 U7995 ( .A(n5100), .Y(n5099) );
  INVX3 U7996 ( .A(n5193), .Y(n5185) );
  INVX3 U7997 ( .A(n5190), .Y(n5189) );
  INVX3 U7998 ( .A(n5117), .Y(n5098) );
  INVX3 U7999 ( .A(n4908), .Y(n4892) );
  INVX3 U8000 ( .A(n4910), .Y(n4893) );
  INVX3 U8001 ( .A(n4763), .Y(n4736) );
  INVX3 U8002 ( .A(n4916), .Y(n4895) );
  INVX3 U8003 ( .A(n4758), .Y(n4735) );
  INVX3 U8004 ( .A(n4750), .Y(n4738) );
  INVX3 U8005 ( .A(n4907), .Y(n4894) );
  INVX3 U8006 ( .A(n5343), .Y(n5317) );
  INVX3 U8007 ( .A(n5236), .Y(n5231) );
  INVX3 U8008 ( .A(n5145), .Y(n5142) );
  INVX3 U8009 ( .A(n5055), .Y(n5052) );
  INVX3 U8010 ( .A(n5328), .Y(n5314) );
  INVX3 U8011 ( .A(n5238), .Y(n5225) );
  INVX3 U8012 ( .A(n5059), .Y(n5045) );
  INVX3 U8013 ( .A(n5324), .Y(n5319) );
  INVX3 U8014 ( .A(n5254), .Y(n5230) );
  INVX3 U8015 ( .A(n5327), .Y(n5315) );
  INVX3 U8016 ( .A(n5254), .Y(n5226) );
  INVX3 U8017 ( .A(n5325), .Y(n5318) );
  INVX3 U8018 ( .A(n5253), .Y(n5229) );
  INVX3 U8019 ( .A(n5237), .Y(n5228) );
  INVX3 U8020 ( .A(n5146), .Y(n5139) );
  INVX3 U8021 ( .A(n5343), .Y(n5320) );
  INVX3 U8022 ( .A(n5252), .Y(n5232) );
  INVX3 U8023 ( .A(n5323), .Y(n5321) );
  INVX3 U8024 ( .A(n5235), .Y(n5233) );
  INVX3 U8025 ( .A(n5144), .Y(n5143) );
  INVX3 U8026 ( .A(n5343), .Y(n5322) );
  INVX3 U8027 ( .A(n5326), .Y(n5316) );
  INVX3 U8028 ( .A(n4705), .Y(n4702) );
  INVX3 U8029 ( .A(n4705), .Y(n4704) );
  INVX3 U8030 ( .A(n4705), .Y(n4703) );
  CLKBUFX3 U8031 ( .A(n4932), .Y(n4903) );
  CLKBUFX3 U8032 ( .A(n4841), .Y(n4815) );
  CLKBUFX3 U8033 ( .A(n4995), .Y(n4967) );
  CLKBUFX3 U8034 ( .A(n5129), .Y(n5101) );
  CLKBUFX3 U8035 ( .A(n5221), .Y(n5193) );
  CLKBUFX3 U8036 ( .A(n5131), .Y(n5100) );
  CLKBUFX3 U8037 ( .A(n5222), .Y(n5190) );
  CLKBUFX3 U8038 ( .A(n5222), .Y(n5191) );
  CLKBUFX3 U8039 ( .A(n5221), .Y(n5192) );
  CLKBUFX3 U8040 ( .A(n4932), .Y(n4907) );
  CLKBUFX3 U8041 ( .A(n4842), .Y(n4811) );
  CLKBUFX3 U8042 ( .A(n4841), .Y(n4813) );
  CLKBUFX3 U8043 ( .A(n4772), .Y(n4742) );
  CLKBUFX3 U8044 ( .A(n4841), .Y(n4812) );
  CLKBUFX3 U8045 ( .A(n4932), .Y(n4908) );
  CLKBUFX3 U8046 ( .A(n4841), .Y(n4814) );
  CLKBUFX3 U8047 ( .A(n4843), .Y(n4810) );
  CLKBUFX3 U8048 ( .A(n4933), .Y(n4905) );
  CLKBUFX3 U8049 ( .A(n4933), .Y(n4906) );
  CLKBUFX3 U8050 ( .A(n4996), .Y(n4966) );
  CLKBUFX3 U8051 ( .A(n4887), .Y(n4860) );
  CLKBUFX3 U8052 ( .A(n5177), .Y(n5150) );
  CLKBUFX3 U8053 ( .A(n5354), .Y(n5326) );
  CLKBUFX3 U8054 ( .A(n5177), .Y(n5148) );
  CLKBUFX3 U8055 ( .A(n5354), .Y(n5327) );
  CLKBUFX3 U8056 ( .A(n5177), .Y(n5149) );
  CLKBUFX3 U8057 ( .A(n5177), .Y(n5147) );
  CLKBUFX3 U8058 ( .A(n5178), .Y(n5146) );
  CLKBUFX3 U8059 ( .A(n5267), .Y(n5237) );
  CLKBUFX3 U8060 ( .A(n5355), .Y(n5325) );
  CLKBUFX3 U8061 ( .A(n5344), .Y(n5323) );
  CLKBUFX3 U8062 ( .A(n5166), .Y(n5144) );
  CLKBUFX3 U8063 ( .A(n5354), .Y(n5328) );
  CLKBUFX3 U8064 ( .A(n5355), .Y(n5324) );
  CLKBUFX3 U8065 ( .A(n5178), .Y(n5145) );
  CLKBUFX3 U8066 ( .A(n5039), .Y(n5011) );
  CLKBUFX3 U8067 ( .A(n5039), .Y(n5012) );
  CLKBUFX3 U8068 ( .A(n5038), .Y(n5013) );
  CLKBUFX3 U8069 ( .A(n4888), .Y(n4857) );
  CLKBUFX3 U8070 ( .A(n4887), .Y(n4858) );
  CLKBUFX3 U8071 ( .A(n4887), .Y(n4859) );
  CLKBUFX3 U8072 ( .A(n5039), .Y(n5010) );
  CLKBUFX3 U8073 ( .A(n4889), .Y(n4856) );
  CLKBUFX3 U8074 ( .A(n4769), .Y(n4753) );
  CLKBUFX3 U8075 ( .A(n4992), .Y(n4978) );
  CLKBUFX3 U8076 ( .A(n4838), .Y(n4829) );
  CLKBUFX3 U8077 ( .A(n4838), .Y(n4831) );
  CLKBUFX3 U8078 ( .A(n4771), .Y(n4744) );
  CLKBUFX3 U8079 ( .A(n4771), .Y(n4745) );
  CLKBUFX3 U8080 ( .A(n4770), .Y(n4749) );
  CLKBUFX3 U8081 ( .A(n4770), .Y(n4748) );
  CLKBUFX3 U8082 ( .A(n4769), .Y(n4752) );
  CLKBUFX3 U8083 ( .A(n4930), .Y(n4914) );
  CLKBUFX3 U8084 ( .A(n4924), .Y(n4917) );
  CLKBUFX3 U8085 ( .A(n4991), .Y(n4982) );
  CLKBUFX3 U8086 ( .A(n4992), .Y(n4983) );
  CLKBUFX3 U8087 ( .A(n4993), .Y(n4975) );
  CLKBUFX3 U8088 ( .A(n5216), .Y(n5194) );
  CLKBUFX3 U8089 ( .A(n4993), .Y(n4974) );
  CLKBUFX3 U8090 ( .A(n4992), .Y(n4977) );
  CLKBUFX3 U8091 ( .A(n5218), .Y(n5202) );
  CLKBUFX3 U8092 ( .A(n5134), .Y(n5113) );
  CLKBUFX3 U8093 ( .A(n4770), .Y(n4746) );
  CLKBUFX3 U8094 ( .A(n5218), .Y(n5204) );
  CLKBUFX3 U8095 ( .A(n5128), .Y(n5105) );
  CLKBUFX3 U8096 ( .A(n4838), .Y(n4828) );
  CLKBUFX3 U8097 ( .A(n5224), .Y(n5196) );
  CLKBUFX3 U8098 ( .A(n4767), .Y(n4759) );
  CLKBUFX3 U8099 ( .A(n4769), .Y(n4751) );
  CLKBUFX3 U8100 ( .A(n4768), .Y(n4757) );
  CLKBUFX3 U8101 ( .A(n4770), .Y(n4747) );
  CLKBUFX3 U8102 ( .A(n5127), .Y(n5110) );
  CLKBUFX3 U8103 ( .A(n5126), .Y(n5115) );
  CLKBUFX3 U8104 ( .A(n5217), .Y(n5205) );
  CLKBUFX3 U8105 ( .A(n5218), .Y(n5201) );
  CLKBUFX3 U8106 ( .A(n5217), .Y(n5206) );
  CLKBUFX3 U8107 ( .A(n4993), .Y(n4972) );
  CLKBUFX3 U8108 ( .A(n4992), .Y(n4976) );
  CLKBUFX3 U8109 ( .A(n5125), .Y(n5119) );
  CLKBUFX3 U8110 ( .A(n5216), .Y(n5209) );
  CLKBUFX3 U8111 ( .A(n4992), .Y(n4984) );
  CLKBUFX3 U8112 ( .A(n4991), .Y(n4985) );
  CLKBUFX3 U8113 ( .A(n5127), .Y(n5107) );
  CLKBUFX3 U8114 ( .A(n5219), .Y(n5198) );
  CLKBUFX3 U8115 ( .A(n5127), .Y(n5108) );
  CLKBUFX3 U8116 ( .A(n5219), .Y(n5199) );
  CLKBUFX3 U8117 ( .A(n5127), .Y(n5106) );
  CLKBUFX3 U8118 ( .A(n5219), .Y(n5197) );
  CLKBUFX3 U8119 ( .A(n5217), .Y(n5207) );
  CLKBUFX3 U8120 ( .A(n5126), .Y(n5116) );
  CLKBUFX3 U8121 ( .A(n5125), .Y(n5118) );
  CLKBUFX3 U8122 ( .A(n5217), .Y(n5208) );
  CLKBUFX3 U8123 ( .A(n5126), .Y(n5117) );
  CLKBUFX3 U8124 ( .A(n5219), .Y(n5200) );
  CLKBUFX3 U8125 ( .A(n5127), .Y(n5109) );
  CLKBUFX3 U8126 ( .A(n5037), .Y(n5022) );
  CLKBUFX3 U8127 ( .A(n4884), .Y(n4876) );
  CLKBUFX3 U8128 ( .A(n4885), .Y(n4868) );
  CLKBUFX3 U8129 ( .A(n4890), .Y(n4867) );
  CLKBUFX3 U8130 ( .A(n5177), .Y(n5151) );
  CLKBUFX3 U8131 ( .A(n5353), .Y(n5330) );
  CLKBUFX3 U8132 ( .A(n5353), .Y(n5329) );
  CLKBUFX3 U8133 ( .A(n5179), .Y(n5159) );
  CLKBUFX3 U8134 ( .A(n5351), .Y(n5338) );
  CLKBUFX3 U8135 ( .A(n5179), .Y(n5153) );
  CLKBUFX3 U8136 ( .A(n5356), .Y(n5345) );
  CLKBUFX3 U8137 ( .A(n5349), .Y(n5347) );
  CLKBUFX3 U8138 ( .A(n5180), .Y(n5169) );
  CLKBUFX3 U8139 ( .A(n5351), .Y(n5339) );
  CLKBUFX3 U8140 ( .A(n5350), .Y(n5340) );
  CLKBUFX3 U8141 ( .A(n5351), .Y(n5337) );
  CLKBUFX3 U8142 ( .A(n5350), .Y(n5341) );
  CLKBUFX3 U8143 ( .A(n4890), .Y(n4866) );
  CLKBUFX3 U8144 ( .A(n5263), .Y(n5251) );
  CLKBUFX3 U8145 ( .A(n5175), .Y(n5157) );
  CLKBUFX3 U8146 ( .A(n5174), .Y(n5162) );
  CLKBUFX3 U8147 ( .A(n4890), .Y(n4877) );
  CLKBUFX3 U8148 ( .A(n4886), .Y(n4878) );
  CLKBUFX3 U8149 ( .A(n5352), .Y(n5334) );
  CLKBUFX3 U8150 ( .A(n5352), .Y(n5335) );
  CLKBUFX3 U8151 ( .A(n5352), .Y(n5333) );
  CLKBUFX3 U8152 ( .A(n5174), .Y(n5163) );
  CLKBUFX3 U8153 ( .A(n5173), .Y(n5165) );
  CLKBUFX3 U8154 ( .A(n5350), .Y(n5343) );
  CLKBUFX3 U8155 ( .A(n5174), .Y(n5164) );
  CLKBUFX3 U8156 ( .A(n5352), .Y(n5336) );
  CLKINVX1 U8157 ( .A(n8229), .Y(n8230) );
  CLKBUFX3 U8158 ( .A(net112034), .Y(net112032) );
  CLKBUFX3 U8159 ( .A(n11003), .Y(n5524) );
  INVX3 U8160 ( .A(n4945), .Y(n4944) );
  INVX3 U8161 ( .A(n4790), .Y(n4786) );
  CLKBUFX3 U8162 ( .A(n10864), .Y(n5464) );
  INVX3 U8163 ( .A(n5281), .Y(n5274) );
  INVX3 U8164 ( .A(n5280), .Y(n5275) );
  INVX3 U8165 ( .A(n5279), .Y(n5276) );
  INVX3 U8166 ( .A(n5278), .Y(n5277) );
  CLKBUFX3 U8167 ( .A(n5954), .Y(n5837) );
  CLKBUFX3 U8168 ( .A(n5954), .Y(n5838) );
  CLKBUFX3 U8169 ( .A(n5953), .Y(n5839) );
  CLKBUFX3 U8170 ( .A(n5953), .Y(n5840) );
  CLKBUFX3 U8171 ( .A(n5953), .Y(n5841) );
  CLKBUFX3 U8172 ( .A(n5953), .Y(n5842) );
  CLKBUFX3 U8173 ( .A(n5953), .Y(n5843) );
  CLKBUFX3 U8174 ( .A(n5953), .Y(n5844) );
  CLKBUFX3 U8175 ( .A(n5953), .Y(n5845) );
  CLKBUFX3 U8176 ( .A(n5954), .Y(n5827) );
  CLKBUFX3 U8177 ( .A(n5954), .Y(n5828) );
  CLKBUFX3 U8178 ( .A(n5954), .Y(n5829) );
  CLKBUFX3 U8179 ( .A(n5954), .Y(n5830) );
  CLKBUFX3 U8180 ( .A(n5954), .Y(n5831) );
  CLKBUFX3 U8181 ( .A(n5954), .Y(n5832) );
  CLKBUFX3 U8182 ( .A(n5954), .Y(n5833) );
  CLKBUFX3 U8183 ( .A(n5954), .Y(n5834) );
  CLKBUFX3 U8184 ( .A(n5954), .Y(n5835) );
  CLKBUFX3 U8185 ( .A(n5954), .Y(n5836) );
  CLKBUFX3 U8186 ( .A(n5952), .Y(n5857) );
  CLKBUFX3 U8187 ( .A(n5952), .Y(n5858) );
  CLKBUFX3 U8188 ( .A(n5952), .Y(n5859) );
  CLKBUFX3 U8189 ( .A(n5952), .Y(n5860) );
  CLKBUFX3 U8190 ( .A(n5952), .Y(n5861) );
  CLKBUFX3 U8191 ( .A(n5952), .Y(n5862) );
  CLKBUFX3 U8192 ( .A(n5951), .Y(n5863) );
  CLKBUFX3 U8193 ( .A(n5951), .Y(n5864) );
  CLKBUFX3 U8194 ( .A(n5951), .Y(n5865) );
  CLKBUFX3 U8195 ( .A(n5953), .Y(n5846) );
  CLKBUFX3 U8196 ( .A(n5953), .Y(n5847) );
  CLKBUFX3 U8197 ( .A(n5953), .Y(n5848) );
  CLKBUFX3 U8198 ( .A(n5953), .Y(n5849) );
  CLKBUFX3 U8199 ( .A(n5953), .Y(n5850) );
  CLKBUFX3 U8200 ( .A(n5952), .Y(n5851) );
  CLKBUFX3 U8201 ( .A(n5952), .Y(n5852) );
  CLKBUFX3 U8202 ( .A(n5952), .Y(n5853) );
  CLKBUFX3 U8203 ( .A(n5952), .Y(n5854) );
  CLKBUFX3 U8204 ( .A(n5952), .Y(n5855) );
  CLKBUFX3 U8205 ( .A(n5952), .Y(n5856) );
  CLKBUFX3 U8206 ( .A(n5957), .Y(n5797) );
  CLKBUFX3 U8207 ( .A(n5957), .Y(n5798) );
  CLKBUFX3 U8208 ( .A(n5957), .Y(n5799) );
  CLKBUFX3 U8209 ( .A(n5957), .Y(n5800) );
  CLKBUFX3 U8210 ( .A(n5957), .Y(n5801) );
  CLKBUFX3 U8211 ( .A(n5957), .Y(n5802) );
  CLKBUFX3 U8212 ( .A(n5956), .Y(n5803) );
  CLKBUFX3 U8213 ( .A(n5956), .Y(n5804) );
  CLKBUFX3 U8214 ( .A(n5956), .Y(n5805) );
  CLKBUFX3 U8215 ( .A(n5958), .Y(n5787) );
  CLKBUFX3 U8216 ( .A(n5958), .Y(n5788) );
  CLKBUFX3 U8217 ( .A(n5958), .Y(n5789) );
  CLKBUFX3 U8218 ( .A(n5958), .Y(n5790) );
  CLKBUFX3 U8219 ( .A(n5957), .Y(n5791) );
  CLKBUFX3 U8220 ( .A(n5957), .Y(n5792) );
  CLKBUFX3 U8221 ( .A(n5957), .Y(n5793) );
  CLKBUFX3 U8222 ( .A(n5957), .Y(n5794) );
  CLKBUFX3 U8223 ( .A(n5957), .Y(n5795) );
  CLKBUFX3 U8224 ( .A(n5957), .Y(n5796) );
  CLKBUFX3 U8225 ( .A(n5955), .Y(n5817) );
  CLKBUFX3 U8226 ( .A(n5955), .Y(n5818) );
  CLKBUFX3 U8227 ( .A(n5955), .Y(n5819) );
  CLKBUFX3 U8228 ( .A(n5955), .Y(n5820) );
  CLKBUFX3 U8229 ( .A(n5955), .Y(n5821) );
  CLKBUFX3 U8230 ( .A(n5955), .Y(n5822) );
  CLKBUFX3 U8231 ( .A(n5955), .Y(n5823) );
  CLKBUFX3 U8232 ( .A(n5955), .Y(n5824) );
  CLKBUFX3 U8233 ( .A(n5955), .Y(n5825) );
  CLKBUFX3 U8234 ( .A(n5956), .Y(n5806) );
  CLKBUFX3 U8235 ( .A(n5956), .Y(n5807) );
  CLKBUFX3 U8236 ( .A(n5956), .Y(n5808) );
  CLKBUFX3 U8237 ( .A(n5956), .Y(n5809) );
  CLKBUFX3 U8238 ( .A(n5956), .Y(n5810) );
  CLKBUFX3 U8239 ( .A(n5956), .Y(n5811) );
  CLKBUFX3 U8240 ( .A(n5956), .Y(n5812) );
  CLKBUFX3 U8241 ( .A(n5956), .Y(n5813) );
  CLKBUFX3 U8242 ( .A(n5956), .Y(n5814) );
  CLKBUFX3 U8243 ( .A(n5955), .Y(n5815) );
  CLKBUFX3 U8244 ( .A(n5955), .Y(n5816) );
  CLKBUFX3 U8245 ( .A(n5955), .Y(n5826) );
  CLKBUFX3 U8246 ( .A(n5948), .Y(n5917) );
  CLKBUFX3 U8247 ( .A(n5948), .Y(n5918) );
  CLKBUFX3 U8248 ( .A(n5948), .Y(n5919) );
  CLKBUFX3 U8249 ( .A(n5948), .Y(n5920) );
  CLKBUFX3 U8250 ( .A(n5948), .Y(n5921) );
  CLKBUFX3 U8251 ( .A(n5948), .Y(n5922) );
  CLKBUFX3 U8252 ( .A(n5947), .Y(n5923) );
  CLKBUFX3 U8253 ( .A(n5947), .Y(n5924) );
  CLKBUFX3 U8254 ( .A(n5947), .Y(n5925) );
  CLKBUFX3 U8255 ( .A(n5971), .Y(n5907) );
  CLKBUFX3 U8256 ( .A(n5961), .Y(n5908) );
  CLKBUFX3 U8257 ( .A(n5947), .Y(n5909) );
  CLKBUFX3 U8258 ( .A(n5966), .Y(n5910) );
  CLKBUFX3 U8259 ( .A(n5948), .Y(n5911) );
  CLKBUFX3 U8260 ( .A(n5948), .Y(n5912) );
  CLKBUFX3 U8261 ( .A(n5948), .Y(n5913) );
  CLKBUFX3 U8262 ( .A(n5948), .Y(n5914) );
  CLKBUFX3 U8263 ( .A(n5948), .Y(n5915) );
  CLKBUFX3 U8264 ( .A(n5948), .Y(n5916) );
  CLKBUFX3 U8265 ( .A(n5946), .Y(n5937) );
  CLKBUFX3 U8266 ( .A(n5946), .Y(n5938) );
  CLKBUFX3 U8267 ( .A(n5968), .Y(n5659) );
  CLKBUFX3 U8268 ( .A(n5968), .Y(n5660) );
  CLKBUFX3 U8269 ( .A(n5968), .Y(n5661) );
  CLKBUFX3 U8270 ( .A(n5968), .Y(n5662) );
  CLKBUFX3 U8271 ( .A(n5968), .Y(n5663) );
  CLKBUFX3 U8272 ( .A(n5968), .Y(n5664) );
  CLKBUFX3 U8273 ( .A(n5968), .Y(n5665) );
  CLKBUFX3 U8274 ( .A(n5968), .Y(n5666) );
  CLKBUFX3 U8275 ( .A(n5960), .Y(n5757) );
  CLKBUFX3 U8276 ( .A(n5960), .Y(n5758) );
  CLKBUFX3 U8277 ( .A(n5960), .Y(n5759) );
  CLKBUFX3 U8278 ( .A(n5960), .Y(n5760) );
  CLKBUFX3 U8279 ( .A(n5960), .Y(n5761) );
  CLKBUFX3 U8280 ( .A(n5960), .Y(n5762) );
  CLKBUFX3 U8281 ( .A(n5960), .Y(n5763) );
  CLKBUFX3 U8282 ( .A(n5960), .Y(n5764) );
  CLKBUFX3 U8283 ( .A(n5960), .Y(n5765) );
  CLKBUFX3 U8284 ( .A(n5961), .Y(n5747) );
  CLKBUFX3 U8285 ( .A(n5961), .Y(n5748) );
  CLKBUFX3 U8286 ( .A(n5961), .Y(n5749) );
  CLKBUFX3 U8287 ( .A(n5961), .Y(n5750) );
  CLKBUFX3 U8288 ( .A(n5961), .Y(n5751) );
  CLKBUFX3 U8289 ( .A(n5961), .Y(n5752) );
  CLKBUFX3 U8290 ( .A(n5961), .Y(n5753) );
  CLKBUFX3 U8291 ( .A(n5961), .Y(n5754) );
  CLKBUFX3 U8292 ( .A(n5960), .Y(n5755) );
  CLKBUFX3 U8293 ( .A(n5960), .Y(n5756) );
  CLKBUFX3 U8294 ( .A(n5959), .Y(n5777) );
  CLKBUFX3 U8295 ( .A(n5959), .Y(n5778) );
  CLKBUFX3 U8296 ( .A(n5958), .Y(n5779) );
  CLKBUFX3 U8297 ( .A(n5958), .Y(n5780) );
  CLKBUFX3 U8298 ( .A(n5958), .Y(n5781) );
  CLKBUFX3 U8299 ( .A(n5958), .Y(n5782) );
  CLKBUFX3 U8300 ( .A(n5958), .Y(n5783) );
  CLKBUFX3 U8301 ( .A(n5958), .Y(n5784) );
  CLKBUFX3 U8302 ( .A(n5958), .Y(n5785) );
  CLKBUFX3 U8303 ( .A(n5960), .Y(n5766) );
  CLKBUFX3 U8304 ( .A(n5959), .Y(n5767) );
  CLKBUFX3 U8305 ( .A(n5959), .Y(n5768) );
  CLKBUFX3 U8306 ( .A(n5959), .Y(n5769) );
  CLKBUFX3 U8307 ( .A(n5959), .Y(n5770) );
  CLKBUFX3 U8308 ( .A(n5959), .Y(n5771) );
  CLKBUFX3 U8309 ( .A(n5959), .Y(n5772) );
  CLKBUFX3 U8310 ( .A(n5959), .Y(n5773) );
  CLKBUFX3 U8311 ( .A(n5959), .Y(n5774) );
  CLKBUFX3 U8312 ( .A(n5959), .Y(n5775) );
  CLKBUFX3 U8313 ( .A(n5959), .Y(n5776) );
  CLKBUFX3 U8314 ( .A(n5964), .Y(n5717) );
  CLKBUFX3 U8315 ( .A(n5964), .Y(n5718) );
  CLKBUFX3 U8316 ( .A(n5963), .Y(n5719) );
  CLKBUFX3 U8317 ( .A(n5963), .Y(n5720) );
  CLKBUFX3 U8318 ( .A(n5963), .Y(n5721) );
  CLKBUFX3 U8319 ( .A(n5963), .Y(n5722) );
  CLKBUFX3 U8320 ( .A(n5963), .Y(n5723) );
  CLKBUFX3 U8321 ( .A(n5963), .Y(n5724) );
  CLKBUFX3 U8322 ( .A(n5963), .Y(n5725) );
  CLKBUFX3 U8323 ( .A(n5964), .Y(n5707) );
  CLKBUFX3 U8324 ( .A(n5964), .Y(n5708) );
  CLKBUFX3 U8325 ( .A(n5964), .Y(n5709) );
  CLKBUFX3 U8326 ( .A(n5964), .Y(n5710) );
  CLKBUFX3 U8327 ( .A(n5964), .Y(n5711) );
  CLKBUFX3 U8328 ( .A(n5964), .Y(n5712) );
  CLKBUFX3 U8329 ( .A(n5946), .Y(n5939) );
  CLKBUFX3 U8330 ( .A(n5946), .Y(n5940) );
  CLKBUFX3 U8331 ( .A(n5946), .Y(n5941) );
  CLKBUFX3 U8332 ( .A(n5946), .Y(n5942) );
  CLKBUFX3 U8333 ( .A(n5946), .Y(n5943) );
  CLKBUFX3 U8334 ( .A(n5946), .Y(n5944) );
  CLKBUFX3 U8335 ( .A(n5946), .Y(n5945) );
  CLKBUFX3 U8336 ( .A(n5947), .Y(n5926) );
  CLKBUFX3 U8337 ( .A(n5947), .Y(n5927) );
  CLKBUFX3 U8338 ( .A(n5947), .Y(n5928) );
  CLKBUFX3 U8339 ( .A(n5947), .Y(n5929) );
  CLKBUFX3 U8340 ( .A(n5947), .Y(n5930) );
  CLKBUFX3 U8341 ( .A(n5947), .Y(n5931) );
  CLKBUFX3 U8342 ( .A(n5947), .Y(n5932) );
  CLKBUFX3 U8343 ( .A(n5947), .Y(n5933) );
  CLKBUFX3 U8344 ( .A(n5947), .Y(n5934) );
  CLKBUFX3 U8345 ( .A(n5946), .Y(n5935) );
  CLKBUFX3 U8346 ( .A(n5946), .Y(n5936) );
  CLKBUFX3 U8347 ( .A(n5950), .Y(n5877) );
  CLKBUFX3 U8348 ( .A(n5950), .Y(n5878) );
  CLKBUFX3 U8349 ( .A(n5950), .Y(n5879) );
  CLKBUFX3 U8350 ( .A(n5950), .Y(n5880) );
  CLKBUFX3 U8351 ( .A(n5950), .Y(n5881) );
  CLKBUFX3 U8352 ( .A(n5950), .Y(n5882) );
  CLKBUFX3 U8353 ( .A(n5950), .Y(n5883) );
  CLKBUFX3 U8354 ( .A(n5950), .Y(n5884) );
  CLKBUFX3 U8355 ( .A(n5950), .Y(n5885) );
  CLKBUFX3 U8356 ( .A(n5951), .Y(n5866) );
  CLKBUFX3 U8357 ( .A(n5951), .Y(n5867) );
  CLKBUFX3 U8358 ( .A(n5951), .Y(n5868) );
  CLKBUFX3 U8359 ( .A(n5951), .Y(n5869) );
  CLKBUFX3 U8360 ( .A(n5951), .Y(n5870) );
  CLKBUFX3 U8361 ( .A(n5951), .Y(n5871) );
  CLKBUFX3 U8362 ( .A(n5951), .Y(n5872) );
  CLKBUFX3 U8363 ( .A(n5951), .Y(n5873) );
  CLKBUFX3 U8364 ( .A(n5951), .Y(n5874) );
  CLKBUFX3 U8365 ( .A(n5950), .Y(n5875) );
  CLKBUFX3 U8366 ( .A(n5950), .Y(n5876) );
  CLKBUFX3 U8367 ( .A(n5949), .Y(n5897) );
  CLKBUFX3 U8368 ( .A(n5949), .Y(n5898) );
  CLKBUFX3 U8369 ( .A(n5959), .Y(n5899) );
  CLKBUFX3 U8370 ( .A(n5969), .Y(n5900) );
  CLKBUFX3 U8371 ( .A(n5960), .Y(n5901) );
  CLKBUFX3 U8372 ( .A(n5958), .Y(n5902) );
  CLKBUFX3 U8373 ( .A(n5962), .Y(n5903) );
  CLKBUFX3 U8374 ( .A(n5970), .Y(n5904) );
  CLKBUFX3 U8375 ( .A(n5956), .Y(n5905) );
  CLKBUFX3 U8376 ( .A(n5950), .Y(n5886) );
  CLKBUFX3 U8377 ( .A(n5949), .Y(n5887) );
  CLKBUFX3 U8378 ( .A(n5949), .Y(n5888) );
  CLKBUFX3 U8379 ( .A(n5949), .Y(n5889) );
  CLKBUFX3 U8380 ( .A(n5949), .Y(n5890) );
  CLKBUFX3 U8381 ( .A(n5949), .Y(n5891) );
  CLKBUFX3 U8382 ( .A(n5949), .Y(n5892) );
  CLKBUFX3 U8383 ( .A(n5949), .Y(n5893) );
  CLKBUFX3 U8384 ( .A(n5949), .Y(n5894) );
  CLKBUFX3 U8385 ( .A(n5949), .Y(n5895) );
  CLKBUFX3 U8386 ( .A(n5949), .Y(n5896) );
  CLKBUFX3 U8387 ( .A(n5953), .Y(n5906) );
  CLKBUFX3 U8388 ( .A(n5967), .Y(n5677) );
  CLKBUFX3 U8389 ( .A(n5967), .Y(n5678) );
  CLKBUFX3 U8390 ( .A(n5967), .Y(n5679) );
  CLKBUFX3 U8391 ( .A(n5967), .Y(n5680) );
  CLKBUFX3 U8392 ( .A(n5967), .Y(n5681) );
  CLKBUFX3 U8393 ( .A(n5967), .Y(n5682) );
  CLKBUFX3 U8394 ( .A(n5966), .Y(n5683) );
  CLKBUFX3 U8395 ( .A(n5966), .Y(n5684) );
  CLKBUFX3 U8396 ( .A(n5966), .Y(n5685) );
  CLKBUFX3 U8397 ( .A(n5968), .Y(n5667) );
  CLKBUFX3 U8398 ( .A(n5968), .Y(n5668) );
  CLKBUFX3 U8399 ( .A(n5968), .Y(n5669) );
  CLKBUFX3 U8400 ( .A(n5968), .Y(n5670) );
  CLKBUFX3 U8401 ( .A(n5967), .Y(n5671) );
  CLKBUFX3 U8402 ( .A(n5967), .Y(n5672) );
  CLKBUFX3 U8403 ( .A(n5967), .Y(n5673) );
  CLKBUFX3 U8404 ( .A(n5967), .Y(n5674) );
  CLKBUFX3 U8405 ( .A(n5967), .Y(n5675) );
  CLKBUFX3 U8406 ( .A(n5967), .Y(n5676) );
  CLKBUFX3 U8407 ( .A(n5965), .Y(n5697) );
  CLKBUFX3 U8408 ( .A(n5965), .Y(n5698) );
  CLKBUFX3 U8409 ( .A(n5965), .Y(n5699) );
  CLKBUFX3 U8410 ( .A(n5965), .Y(n5700) );
  CLKBUFX3 U8411 ( .A(n5965), .Y(n5701) );
  CLKBUFX3 U8412 ( .A(n5965), .Y(n5702) );
  CLKBUFX3 U8413 ( .A(n5965), .Y(n5703) );
  CLKBUFX3 U8414 ( .A(n5965), .Y(n5704) );
  CLKBUFX3 U8415 ( .A(n5965), .Y(n5705) );
  CLKBUFX3 U8416 ( .A(n5965), .Y(n5706) );
  CLKBUFX3 U8417 ( .A(n5966), .Y(n5686) );
  CLKBUFX3 U8418 ( .A(n5966), .Y(n5687) );
  CLKBUFX3 U8419 ( .A(n5966), .Y(n5688) );
  CLKBUFX3 U8420 ( .A(n5966), .Y(n5689) );
  CLKBUFX3 U8421 ( .A(n5966), .Y(n5690) );
  CLKBUFX3 U8422 ( .A(n5966), .Y(n5691) );
  CLKBUFX3 U8423 ( .A(n5966), .Y(n5692) );
  CLKBUFX3 U8424 ( .A(n5966), .Y(n5693) );
  CLKBUFX3 U8425 ( .A(n5966), .Y(n5694) );
  CLKBUFX3 U8426 ( .A(n5965), .Y(n5695) );
  CLKBUFX3 U8427 ( .A(n5965), .Y(n5696) );
  CLKBUFX3 U8428 ( .A(n5964), .Y(n5713) );
  CLKBUFX3 U8429 ( .A(n5964), .Y(n5714) );
  CLKBUFX3 U8430 ( .A(n5964), .Y(n5715) );
  CLKBUFX3 U8431 ( .A(n5964), .Y(n5716) );
  CLKBUFX3 U8432 ( .A(n5962), .Y(n5737) );
  CLKBUFX3 U8433 ( .A(n5962), .Y(n5738) );
  CLKBUFX3 U8434 ( .A(n5962), .Y(n5739) );
  CLKBUFX3 U8435 ( .A(n5962), .Y(n5740) );
  CLKBUFX3 U8436 ( .A(n5962), .Y(n5741) );
  CLKBUFX3 U8437 ( .A(n5962), .Y(n5742) );
  CLKBUFX3 U8438 ( .A(n5963), .Y(n5726) );
  CLKBUFX3 U8439 ( .A(n5963), .Y(n5727) );
  CLKBUFX3 U8440 ( .A(n5963), .Y(n5728) );
  CLKBUFX3 U8441 ( .A(n5963), .Y(n5729) );
  CLKBUFX3 U8442 ( .A(n5963), .Y(n5730) );
  CLKBUFX3 U8443 ( .A(n5962), .Y(n5731) );
  CLKBUFX3 U8444 ( .A(n5962), .Y(n5732) );
  CLKBUFX3 U8445 ( .A(n5962), .Y(n5733) );
  CLKBUFX3 U8446 ( .A(n5962), .Y(n5734) );
  CLKBUFX3 U8447 ( .A(n5962), .Y(n5735) );
  CLKBUFX3 U8448 ( .A(n5962), .Y(n5736) );
  CLKBUFX3 U8449 ( .A(n5958), .Y(n5786) );
  CLKBUFX3 U8450 ( .A(n5961), .Y(n5743) );
  CLKBUFX3 U8451 ( .A(n5961), .Y(n5746) );
  CLKBUFX3 U8452 ( .A(n5961), .Y(n5744) );
  CLKBUFX3 U8453 ( .A(n5961), .Y(n5745) );
  INVX12 U8454 ( .A(n4622), .Y(mem_wdata_D[45]) );
  INVX12 U8455 ( .A(n4606), .Y(mem_wdata_D[106]) );
  INVX12 U8456 ( .A(n4609), .Y(mem_wdata_D[109]) );
  INVX12 U8457 ( .A(n4604), .Y(mem_wdata_D[110]) );
  INVX12 U8458 ( .A(n4607), .Y(mem_wdata_D[113]) );
  INVX12 U8459 ( .A(n4605), .Y(mem_wdata_D[117]) );
  INVX12 U8460 ( .A(n4603), .Y(mem_wdata_D[103]) );
  INVX12 U8461 ( .A(n4600), .Y(mem_wdata_D[107]) );
  INVX12 U8462 ( .A(n4602), .Y(mem_wdata_D[114]) );
  OA22X1 U8463 ( .A0(n10769), .A1(n4245), .B0(n10772), .B1(n4246), .Y(n7853)
         );
  CLKINVX1 U8464 ( .A(n8151), .Y(n8178) );
  OA22X1 U8465 ( .A0(n10713), .A1(n4245), .B0(n10716), .B1(n4246), .Y(n7280)
         );
  AND2XL U8466 ( .A(n11089), .B(n11088), .Y(n4387) );
  OA22X1 U8467 ( .A0(n10294), .A1(n4245), .B0(n10297), .B1(n4246), .Y(n8108)
         );
  OA22X1 U8468 ( .A0(n10145), .A1(n4245), .B0(n10148), .B1(n4246), .Y(n6438)
         );
  CLKBUFX3 U8469 ( .A(net97418), .Y(net108190) );
  CLKBUFX3 U8470 ( .A(net97418), .Y(net108194) );
  CLKBUFX3 U8471 ( .A(n5309), .Y(n5284) );
  CLKBUFX3 U8472 ( .A(n5311), .Y(n5279) );
  CLKBUFX3 U8473 ( .A(n5311), .Y(n5280) );
  CLKBUFX3 U8474 ( .A(n5311), .Y(n5278) );
  CLKBUFX3 U8475 ( .A(n5310), .Y(n5281) );
  CLKINVX1 U8476 ( .A(n10346), .Y(n6296) );
  INVX3 U8477 ( .A(n4478), .Y(n4693) );
  CLKBUFX3 U8478 ( .A(n5308), .Y(n5287) );
  CLKBUFX3 U8479 ( .A(n5307), .Y(n5296) );
  CLKBUFX3 U8480 ( .A(n5305), .Y(n5301) );
  CLKBUFX3 U8481 ( .A(n5306), .Y(n5297) );
  CLKBUFX3 U8482 ( .A(n5307), .Y(n5293) );
  CLKBUFX3 U8483 ( .A(n5307), .Y(n5290) );
  CLKBUFX3 U8484 ( .A(n5295), .Y(n5291) );
  CLKBUFX3 U8485 ( .A(n5295), .Y(n5289) );
  CLKBUFX3 U8486 ( .A(n5305), .Y(n5299) );
  CLKBUFX3 U8487 ( .A(n5307), .Y(n5292) );
  INVX3 U8488 ( .A(n4478), .Y(n4694) );
  INVX3 U8489 ( .A(n5409), .Y(n5407) );
  INVX3 U8490 ( .A(n5409), .Y(n5408) );
  CLKBUFX3 U8491 ( .A(net112084), .Y(net112076) );
  CLKBUFX3 U8492 ( .A(n9533), .Y(n4720) );
  CLKBUFX3 U8493 ( .A(net100601), .Y(net112050) );
  INVX3 U8494 ( .A(n5481), .Y(n5479) );
  CLKBUFX3 U8495 ( .A(n1979), .Y(n5481) );
  INVX3 U8496 ( .A(n5481), .Y(n5480) );
  INVX3 U8497 ( .A(n4777), .Y(n4775) );
  CLKBUFX3 U8498 ( .A(n2000), .Y(n4777) );
  INVX3 U8499 ( .A(n4777), .Y(n4776) );
  INVX3 U8500 ( .A(n1998), .Y(n5469) );
  INVX3 U8501 ( .A(n1993), .Y(n5440) );
  INVX3 U8502 ( .A(n5415), .Y(n5413) );
  CLKBUFX3 U8503 ( .A(n1999), .Y(n5415) );
  INVX3 U8504 ( .A(n1987), .Y(n5460) );
  INVX3 U8505 ( .A(n5439), .Y(n5437) );
  CLKBUFX3 U8506 ( .A(n1985), .Y(n5439) );
  INVX3 U8507 ( .A(n1996), .Y(n5455) );
  INVX3 U8508 ( .A(n4437), .Y(n5453) );
  INVX3 U8509 ( .A(n5447), .Y(n5445) );
  CLKBUFX3 U8510 ( .A(n1989), .Y(n5447) );
  INVX3 U8511 ( .A(n5421), .Y(n5419) );
  CLKBUFX3 U8512 ( .A(n1990), .Y(n5421) );
  INVX3 U8513 ( .A(n5444), .Y(n5442) );
  INVX3 U8514 ( .A(n1997), .Y(n5474) );
  INVX3 U8515 ( .A(n5044), .Y(n5042) );
  CLKBUFX3 U8516 ( .A(n4391), .Y(n5044) );
  INVX3 U8517 ( .A(n5492), .Y(n5490) );
  CLKBUFX3 U8518 ( .A(n301), .Y(n5492) );
  INVX3 U8519 ( .A(n5489), .Y(n5487) );
  CLKBUFX3 U8520 ( .A(n1986), .Y(n5489) );
  INVX3 U8521 ( .A(n1998), .Y(n5470) );
  INVX3 U8522 ( .A(n1993), .Y(n5441) );
  INVX3 U8523 ( .A(n5415), .Y(n5414) );
  INVX3 U8524 ( .A(n1987), .Y(n5461) );
  INVX3 U8525 ( .A(n5439), .Y(n5438) );
  INVX3 U8526 ( .A(n1996), .Y(n5456) );
  INVX3 U8527 ( .A(n4437), .Y(n5454) );
  INVX3 U8528 ( .A(n5447), .Y(n5446) );
  INVX3 U8529 ( .A(n5421), .Y(n5420) );
  INVX3 U8530 ( .A(n5444), .Y(n5443) );
  CLKBUFX3 U8531 ( .A(n1991), .Y(n5444) );
  INVX3 U8532 ( .A(n1997), .Y(n5475) );
  INVX3 U8533 ( .A(n5492), .Y(n5491) );
  INVX3 U8534 ( .A(n5489), .Y(n5488) );
  INVX3 U8535 ( .A(net112158), .Y(net112148) );
  INVX3 U8536 ( .A(n5424), .Y(n5422) );
  CLKBUFX3 U8537 ( .A(n4411), .Y(n5424) );
  INVX3 U8538 ( .A(n5424), .Y(n5423) );
  CLKBUFX3 U8539 ( .A(n5240), .Y(n5267) );
  NAND2X1 U8540 ( .A(n5468), .B(n5559), .Y(n10864) );
  INVX3 U8541 ( .A(n4488), .Y(n5558) );
  INVX3 U8542 ( .A(n4488), .Y(n5559) );
  CLKBUFX3 U8543 ( .A(n5970), .Y(n5645) );
  CLKBUFX3 U8544 ( .A(n5971), .Y(n5628) );
  CLKBUFX3 U8545 ( .A(n5971), .Y(n5629) );
  CLKBUFX3 U8546 ( .A(n5971), .Y(n5630) );
  CLKBUFX3 U8547 ( .A(n5971), .Y(n5631) );
  CLKBUFX3 U8548 ( .A(n5971), .Y(n5632) );
  CLKBUFX3 U8549 ( .A(n5971), .Y(n5633) );
  CLKBUFX3 U8550 ( .A(n5971), .Y(n5634) );
  CLKBUFX3 U8551 ( .A(n5970), .Y(n5635) );
  CLKBUFX3 U8552 ( .A(n5970), .Y(n5636) );
  CLKBUFX3 U8553 ( .A(n5969), .Y(n5657) );
  CLKBUFX3 U8554 ( .A(n5969), .Y(n5658) );
  CLKBUFX3 U8555 ( .A(n5969), .Y(n5647) );
  CLKBUFX3 U8556 ( .A(n5969), .Y(n5648) );
  CLKBUFX3 U8557 ( .A(n5969), .Y(n5649) );
  CLKBUFX3 U8558 ( .A(n5969), .Y(n5650) );
  CLKBUFX3 U8559 ( .A(n5969), .Y(n5651) );
  CLKBUFX3 U8560 ( .A(n5969), .Y(n5652) );
  CLKBUFX3 U8561 ( .A(n5969), .Y(n5653) );
  CLKBUFX3 U8562 ( .A(n5969), .Y(n5654) );
  CLKBUFX3 U8563 ( .A(n5969), .Y(n5655) );
  CLKBUFX3 U8564 ( .A(n5969), .Y(n5656) );
  CLKBUFX3 U8565 ( .A(n5970), .Y(n5646) );
  CLKBUFX3 U8566 ( .A(n5970), .Y(n5637) );
  CLKBUFX3 U8567 ( .A(n5970), .Y(n5638) );
  CLKBUFX3 U8568 ( .A(n5970), .Y(n5639) );
  CLKBUFX3 U8569 ( .A(n5970), .Y(n5640) );
  CLKBUFX3 U8570 ( .A(n5970), .Y(n5641) );
  CLKBUFX3 U8571 ( .A(n5970), .Y(n5642) );
  CLKBUFX3 U8572 ( .A(n5970), .Y(n5643) );
  CLKBUFX3 U8573 ( .A(n5970), .Y(n5644) );
  CLKBUFX3 U8574 ( .A(n5971), .Y(n5627) );
  CLKBUFX3 U8575 ( .A(rst_n), .Y(n5954) );
  CLKBUFX3 U8576 ( .A(n5972), .Y(n5953) );
  CLKBUFX3 U8577 ( .A(n5972), .Y(n5952) );
  CLKBUFX3 U8578 ( .A(n5972), .Y(n5957) );
  CLKBUFX3 U8579 ( .A(n5972), .Y(n5956) );
  CLKBUFX3 U8580 ( .A(rst_n), .Y(n5955) );
  CLKBUFX3 U8581 ( .A(n5972), .Y(n5948) );
  CLKBUFX3 U8582 ( .A(n5948), .Y(n5960) );
  CLKBUFX3 U8583 ( .A(n5968), .Y(n5959) );
  CLKBUFX3 U8584 ( .A(n5972), .Y(n5947) );
  CLKBUFX3 U8585 ( .A(n5972), .Y(n5946) );
  CLKBUFX3 U8586 ( .A(n5971), .Y(n5951) );
  CLKBUFX3 U8587 ( .A(rst_n), .Y(n5950) );
  CLKBUFX3 U8588 ( .A(rst_n), .Y(n5949) );
  CLKBUFX3 U8589 ( .A(n5972), .Y(n5968) );
  CLKBUFX3 U8590 ( .A(rst_n), .Y(n5967) );
  CLKBUFX3 U8591 ( .A(n5972), .Y(n5966) );
  CLKBUFX3 U8592 ( .A(n5972), .Y(n5965) );
  CLKBUFX3 U8593 ( .A(n5972), .Y(n5964) );
  CLKBUFX3 U8594 ( .A(n5971), .Y(n5963) );
  CLKBUFX3 U8595 ( .A(n5946), .Y(n5962) );
  CLKBUFX3 U8596 ( .A(n5972), .Y(n5961) );
  CLKBUFX3 U8597 ( .A(n5946), .Y(n5958) );
  CLKINVX1 U8598 ( .A(n8871), .Y(n8872) );
  INVX12 U8599 ( .A(n1956), .Y(mem_wdata_D[43]) );
  INVX12 U8600 ( .A(n1958), .Y(mem_wdata_D[91]) );
  INVX12 U8601 ( .A(n1959), .Y(mem_wdata_D[94]) );
  INVX12 U8602 ( .A(n1960), .Y(mem_wdata_D[97]) );
  INVX12 U8603 ( .A(n1962), .Y(mem_wdata_D[104]) );
  INVX12 U8604 ( .A(n1964), .Y(mem_wdata_D[116]) );
  CLKINVX1 U8605 ( .A(n8238), .Y(n8247) );
  INVX12 U8606 ( .A(n1961), .Y(mem_wdata_D[100]) );
  INVX12 U8607 ( .A(n1963), .Y(mem_wdata_D[112]) );
  INVX12 U8608 ( .A(n1965), .Y(mem_wdata_D[118]) );
  INVX12 U8609 ( .A(n1966), .Y(mem_wdata_D[119]) );
  INVX12 U8610 ( .A(n1967), .Y(mem_wdata_D[121]) );
  INVX12 U8611 ( .A(n1968), .Y(mem_wdata_D[124]) );
  INVX12 U8612 ( .A(n1969), .Y(mem_wdata_D[127]) );
  NAND2BX1 U8613 ( .AN(n5429), .B(n11228), .Y(n10060) );
  CLKINVX1 U8614 ( .A(n8075), .Y(n8083) );
  CLKMX2X2 U8615 ( .A(net100573), .B(net112438), .S0(n8079), .Y(n8080) );
  NAND2BX1 U8616 ( .AN(n5429), .B(n11227), .Y(n10036) );
  NAND2BX1 U8617 ( .AN(n5425), .B(n11278), .Y(n6294) );
  NAND2BX1 U8618 ( .AN(n5425), .B(n11277), .Y(n6258) );
  NAND2BX1 U8619 ( .AN(n5429), .B(n11245), .Y(n6256) );
  NAND2X2 U8620 ( .A(n10650), .B(n4571), .Y(n10324) );
  NAND2XL U8621 ( .A(n3416), .B(n10580), .Y(n10692) );
  CLKINVX1 U8622 ( .A(n9348), .Y(n9338) );
  INVXL U8623 ( .A(net101401), .Y(net104248) );
  XOR3XL U8624 ( .A(n11108), .B(n11107), .C(n11106), .Y(n11111) );
  INVXL U8625 ( .A(n10609), .Y(n10610) );
  INVXL U8626 ( .A(n10404), .Y(n10405) );
  INVXL U8627 ( .A(n10389), .Y(n10390) );
  CLKINVX1 U8628 ( .A(n10382), .Y(n10391) );
  AOI2BB1X1 U8629 ( .A0N(n4466), .A1N(n4390), .B0(n10811), .Y(n10813) );
  INVXL U8630 ( .A(n10810), .Y(n10811) );
  AOI2BB1X1 U8631 ( .A0N(n4475), .A1N(n10801), .B0(n10367), .Y(n10369) );
  CLKINVX1 U8632 ( .A(n10366), .Y(n10367) );
  AOI2BB1X1 U8633 ( .A0N(n4387), .A1N(n4435), .B0(n11091), .Y(n11093) );
  INVXL U8634 ( .A(n11090), .Y(n11091) );
  AOI2BB1XL U8635 ( .A0N(n3838), .A1N(net101906), .B0(n8260), .Y(n7466) );
  XOR3XL U8636 ( .A(n11077), .B(n4456), .C(n11076), .Y(n11079) );
  CLKINVX1 U8637 ( .A(n11373), .Y(n10946) );
  CLKINVX1 U8638 ( .A(n11452), .Y(n10067) );
  CLKINVX1 U8639 ( .A(n11362), .Y(n10725) );
  CLKINVX1 U8640 ( .A(n11375), .Y(n10497) );
  CLKINVX1 U8641 ( .A(n11368), .Y(n10514) );
  CLKINVX1 U8642 ( .A(n11384), .Y(n10937) );
  INVXL U8643 ( .A(n8750), .Y(n8754) );
  CLKINVX1 U8644 ( .A(n11469), .Y(n10940) );
  NAND2BX1 U8645 ( .AN(n5425), .B(n11281), .Y(n6282) );
  NAND2BX1 U8646 ( .AN(n5429), .B(n11249), .Y(n6280) );
  NAND2BX1 U8647 ( .AN(n5425), .B(n11276), .Y(n6278) );
  NAND2BX1 U8648 ( .AN(n5429), .B(n11244), .Y(n6276) );
  NAND2BX1 U8649 ( .AN(n4247), .B(n11308), .Y(n6279) );
  NAND2BX1 U8650 ( .AN(n5425), .B(n11279), .Y(n6290) );
  NAND2BXL U8651 ( .AN(n4247), .B(n11311), .Y(n6291) );
  INVXL U8652 ( .A(n260), .Y(n7043) );
  AOI2BB1XL U8653 ( .A0N(n9275), .A1N(n9273), .B0(n9272), .Y(n9278) );
  AND2XL U8654 ( .A(n6), .B(n10285), .Y(n4397) );
  AND2XL U8655 ( .A(n3418), .B(net98550), .Y(n4401) );
  AND2XL U8656 ( .A(net98216), .B(net98217), .Y(n4402) );
  AND2XL U8657 ( .A(n3324), .B(n10926), .Y(n4409) );
  INVXL U8658 ( .A(n10636), .Y(n11007) );
  AND2XL U8659 ( .A(n3423), .B(n10455), .Y(n4410) );
  OA22X1 U8660 ( .A0(n10209), .A1(n4676), .B0(n10212), .B1(n4250), .Y(n9514)
         );
  INVXL U8661 ( .A(n3846), .Y(n10796) );
  AND2XL U8662 ( .A(n10356), .B(n10355), .Y(n4414) );
  CLKINVX1 U8663 ( .A(net104866), .Y(net104230) );
  CLKINVX1 U8664 ( .A(n10173), .Y(n10174) );
  CLKINVX1 U8665 ( .A(n10365), .Y(n10801) );
  NAND2BX1 U8666 ( .AN(n10364), .B(n10363), .Y(n10365) );
  AOI2BB1X1 U8667 ( .A0N(n10362), .A1N(n10361), .B0(n10360), .Y(n10364) );
  CLKINVX1 U8668 ( .A(n8260), .Y(n8263) );
  CLKINVX1 U8669 ( .A(n9354), .Y(n9352) );
  AND2XL U8670 ( .A(n3417), .B(n10548), .Y(n4426) );
  AND2XL U8671 ( .A(n10679), .B(n10678), .Y(n4427) );
  AND2XL U8672 ( .A(n3663), .B(n10530), .Y(n4428) );
  AND2X2 U8673 ( .A(n3321), .B(net98514), .Y(n4429) );
  AND2XL U8674 ( .A(n3414), .B(net98598), .Y(n4431) );
  CLKINVX1 U8675 ( .A(n8745), .Y(n8760) );
  CLKINVX1 U8676 ( .A(n8237), .Y(n6568) );
  CLKINVX1 U8677 ( .A(n9263), .Y(n9253) );
  INVXL U8678 ( .A(n7975), .Y(n7974) );
  CLKINVX1 U8679 ( .A(n8175), .Y(n8162) );
  CLKINVX1 U8680 ( .A(n8726), .Y(n8728) );
  CLKINVX1 U8681 ( .A(n9492), .Y(n9490) );
  CLKINVX1 U8682 ( .A(n8560), .Y(n8562) );
  CLKINVX1 U8683 ( .A(n9067), .Y(n9045) );
  CLKBUFX3 U8684 ( .A(net128159), .Y(net112158) );
  CLKBUFX3 U8685 ( .A(net128155), .Y(net112246) );
  CLKBUFX3 U8686 ( .A(net128154), .Y(net112228) );
  CLKINVX1 U8687 ( .A(n7522), .Y(n7516) );
  CLKBUFX3 U8688 ( .A(net128155), .Y(net112250) );
  CLKBUFX3 U8689 ( .A(net128158), .Y(net112178) );
  CLKBUFX3 U8690 ( .A(net128154), .Y(net112232) );
  CLKBUFX3 U8691 ( .A(net128160), .Y(net112196) );
  CLKBUFX3 U8692 ( .A(net128159), .Y(net112160) );
  AND2X2 U8693 ( .A(n4448), .B(n4445), .Y(n4440) );
  CLKINVX1 U8694 ( .A(n9252), .Y(n9256) );
  CLKINVX1 U8695 ( .A(n9251), .Y(n9257) );
  CLKMX2X2 U8696 ( .A(net100573), .B(net112438), .S0(n9253), .Y(n9254) );
  CLKINVX1 U8697 ( .A(n8181), .Y(n8182) );
  CLKINVX1 U8698 ( .A(n9167), .Y(n9169) );
  CLKINVX1 U8699 ( .A(n7463), .Y(n7467) );
  CLKINVX1 U8700 ( .A(n8959), .Y(n8732) );
  CLKINVX1 U8701 ( .A(n9051), .Y(n7826) );
  AO22X1 U8702 ( .A0(n6760), .A1(net137952), .B0(net112296), .B1(n6759), .Y(
        n6762) );
  AND2XL U8703 ( .A(net111994), .B(n6695), .Y(n6703) );
  CLKINVX1 U8704 ( .A(n7889), .Y(n7879) );
  AND2X2 U8705 ( .A(n8452), .B(n8451), .Y(n8460) );
  INVX1 U8706 ( .A(n8450), .Y(n8452) );
  CLKINVX1 U8707 ( .A(n9476), .Y(n9465) );
  INVX3 U8708 ( .A(n1978), .Y(n5482) );
  INVX3 U8709 ( .A(n1978), .Y(n5483) );
  INVX3 U8710 ( .A(n5418), .Y(n5416) );
  INVX3 U8711 ( .A(n5418), .Y(n5417) );
  INVX3 U8712 ( .A(n5436), .Y(n5434) );
  CLKBUFX3 U8713 ( .A(n1980), .Y(n5436) );
  INVX3 U8714 ( .A(n5459), .Y(n5457) );
  INVX3 U8715 ( .A(n4479), .Y(n5451) );
  INVX3 U8716 ( .A(n5450), .Y(n5448) );
  INVX3 U8717 ( .A(n5436), .Y(n5435) );
  INVX3 U8718 ( .A(n5459), .Y(n5458) );
  CLKBUFX3 U8719 ( .A(n1988), .Y(n5459) );
  INVX3 U8720 ( .A(n4479), .Y(n5452) );
  INVX3 U8721 ( .A(n5450), .Y(n5449) );
  INVX3 U8722 ( .A(n2211), .Y(n5402) );
  INVX3 U8723 ( .A(n2211), .Y(n5403) );
  INVX3 U8724 ( .A(n5433), .Y(n5431) );
  CLKBUFX3 U8725 ( .A(n4458), .Y(n5433) );
  INVX3 U8726 ( .A(n5433), .Y(n5432) );
  INVX3 U8727 ( .A(n5412), .Y(n5410) );
  CLKBUFX3 U8728 ( .A(n1995), .Y(n5412) );
  INVX3 U8729 ( .A(n5406), .Y(n5404) );
  CLKBUFX3 U8730 ( .A(n4442), .Y(n5406) );
  INVX3 U8731 ( .A(n5473), .Y(n5471) );
  CLKBUFX3 U8732 ( .A(n1992), .Y(n5473) );
  INVX3 U8733 ( .A(n5478), .Y(n5476) );
  CLKBUFX3 U8734 ( .A(n302), .Y(n5478) );
  INVX3 U8735 ( .A(n5486), .Y(n5484) );
  CLKBUFX3 U8736 ( .A(n1994), .Y(n5486) );
  INVX3 U8737 ( .A(n5412), .Y(n5411) );
  INVX3 U8738 ( .A(n5406), .Y(n5405) );
  INVX3 U8739 ( .A(n5473), .Y(n5472) );
  INVX3 U8740 ( .A(n5478), .Y(n5477) );
  INVX3 U8741 ( .A(n5486), .Y(n5485) );
  CLKBUFX3 U8742 ( .A(n11002), .Y(n5509) );
  CLKBUFX3 U8743 ( .A(n11171), .Y(n5533) );
  CLKBUFX3 U8744 ( .A(n11171), .Y(n5532) );
  CLKBUFX3 U8745 ( .A(n11002), .Y(n5508) );
  CLKBUFX3 U8746 ( .A(n9527), .Y(n4689) );
  CLKBUFX3 U8747 ( .A(n5090), .Y(n5132) );
  CLKBUFX3 U8748 ( .A(n5534), .Y(n5529) );
  CLKBUFX3 U8749 ( .A(n11171), .Y(n5534) );
  CLKBUFX3 U8750 ( .A(net133468), .Y(net112104) );
  CLKBUFX3 U8751 ( .A(n4349), .Y(n4685) );
  CLKINVX1 U8752 ( .A(net111910), .Y(net111906) );
  NAND4X1 U8753 ( .A(n9638), .B(n9637), .C(n9636), .D(n9635), .Y(n10550) );
  NAND2BXL U8754 ( .AN(n4247), .B(n11302), .Y(n9638) );
  NAND4X1 U8755 ( .A(n9590), .B(n9589), .C(n9588), .D(n9587), .Y(n11124) );
  NAND2BXL U8756 ( .AN(n4247), .B(n11301), .Y(n9590) );
  NAND4X1 U8757 ( .A(n9687), .B(n9686), .C(n9685), .D(n9684), .Y(n10532) );
  NAND2BXL U8758 ( .AN(n4247), .B(n11300), .Y(n9687) );
  NAND4X1 U8759 ( .A(n10644), .B(n10643), .C(n10642), .D(n10641), .Y(n11175)
         );
  NAND2BXL U8760 ( .AN(n4247), .B(n11299), .Y(n10644) );
  NAND4X1 U8761 ( .A(n9736), .B(n9735), .C(n9734), .D(n9733), .Y(n10628) );
  NAND2BXL U8762 ( .AN(n4247), .B(n11298), .Y(n9736) );
  NAND4X1 U8763 ( .A(n9825), .B(n9824), .C(n9823), .D(n9822), .Y(n10840) );
  NAND2BXL U8764 ( .AN(n4247), .B(n11307), .Y(n9825) );
  NAND4X1 U8765 ( .A(n9805), .B(n9804), .C(n9803), .D(n9802), .Y(n10829) );
  NAND2BXL U8766 ( .AN(n4247), .B(n11306), .Y(n9805) );
  NAND4X1 U8767 ( .A(n9845), .B(n9844), .C(n9843), .D(n9842), .Y(n10469) );
  NAND2BXL U8768 ( .AN(n4247), .B(n11305), .Y(n9845) );
  NAND4X1 U8769 ( .A(n9881), .B(n9880), .C(n9879), .D(n9878), .Y(n10457) );
  NAND2BXL U8770 ( .AN(n4247), .B(n11304), .Y(n9881) );
  NAND2BXL U8771 ( .AN(n4247), .B(n11303), .Y(net99633) );
  NAND2BXL U8772 ( .AN(n5428), .B(n11211), .Y(n9823) );
  NAND2BXL U8773 ( .AN(n5428), .B(n11210), .Y(n9803) );
  NAND2BXL U8774 ( .AN(n5428), .B(n11209), .Y(n9843) );
  NAND2BXL U8775 ( .AN(n5427), .B(n11208), .Y(n9879) );
  NAND2BXL U8776 ( .AN(n5427), .B(n11207), .Y(net99635) );
  NAND2BXL U8777 ( .AN(n5428), .B(n11206), .Y(n9636) );
  NAND2BXL U8778 ( .AN(n5428), .B(n11205), .Y(n9588) );
  NAND2BXL U8779 ( .AN(n5428), .B(n11204), .Y(n9685) );
  NAND2BXL U8780 ( .AN(n5428), .B(n11203), .Y(n10642) );
  NAND2BXL U8781 ( .AN(n5428), .B(n11202), .Y(n9734) );
  CLKBUFX3 U8782 ( .A(\i_MIPS/Register/n147 ), .Y(n5621) );
  CLKBUFX3 U8783 ( .A(\i_MIPS/Register/n147 ), .Y(n5620) );
  CLKBUFX3 U8784 ( .A(\i_MIPS/Register/n146 ), .Y(n5618) );
  CLKBUFX3 U8785 ( .A(\i_MIPS/Register/n146 ), .Y(n5619) );
  CLKBUFX3 U8786 ( .A(\i_MIPS/Register/n145 ), .Y(n5616) );
  CLKBUFX3 U8787 ( .A(\i_MIPS/Register/n145 ), .Y(n5617) );
  CLKBUFX3 U8788 ( .A(\i_MIPS/Register/n144 ), .Y(n5614) );
  CLKBUFX3 U8789 ( .A(\i_MIPS/Register/n144 ), .Y(n5615) );
  CLKBUFX3 U8790 ( .A(\i_MIPS/Register/n143 ), .Y(n5612) );
  CLKBUFX3 U8791 ( .A(\i_MIPS/Register/n143 ), .Y(n5613) );
  CLKBUFX3 U8792 ( .A(\i_MIPS/Register/n142 ), .Y(n5610) );
  CLKBUFX3 U8793 ( .A(\i_MIPS/Register/n142 ), .Y(n5611) );
  CLKBUFX3 U8794 ( .A(\i_MIPS/Register/n141 ), .Y(n5608) );
  CLKBUFX3 U8795 ( .A(\i_MIPS/Register/n141 ), .Y(n5609) );
  CLKBUFX3 U8796 ( .A(\i_MIPS/Register/n139 ), .Y(n5606) );
  CLKBUFX3 U8797 ( .A(\i_MIPS/Register/n139 ), .Y(n5607) );
  CLKBUFX3 U8798 ( .A(\i_MIPS/Register/n138 ), .Y(n5604) );
  CLKBUFX3 U8799 ( .A(\i_MIPS/Register/n138 ), .Y(n5605) );
  CLKBUFX3 U8800 ( .A(\i_MIPS/Register/n137 ), .Y(n5602) );
  CLKBUFX3 U8801 ( .A(\i_MIPS/Register/n137 ), .Y(n5603) );
  CLKBUFX3 U8802 ( .A(\i_MIPS/Register/n136 ), .Y(n5600) );
  CLKBUFX3 U8803 ( .A(\i_MIPS/Register/n136 ), .Y(n5601) );
  CLKBUFX3 U8804 ( .A(\i_MIPS/Register/n135 ), .Y(n5598) );
  CLKBUFX3 U8805 ( .A(\i_MIPS/Register/n135 ), .Y(n5599) );
  CLKBUFX3 U8806 ( .A(\i_MIPS/Register/n134 ), .Y(n5596) );
  CLKBUFX3 U8807 ( .A(\i_MIPS/Register/n134 ), .Y(n5597) );
  CLKBUFX3 U8808 ( .A(\i_MIPS/Register/n133 ), .Y(n5594) );
  CLKBUFX3 U8809 ( .A(\i_MIPS/Register/n133 ), .Y(n5595) );
  CLKBUFX3 U8810 ( .A(\i_MIPS/Register/n132 ), .Y(n5592) );
  CLKBUFX3 U8811 ( .A(\i_MIPS/Register/n132 ), .Y(n5593) );
  CLKBUFX3 U8812 ( .A(\i_MIPS/Register/n130 ), .Y(n5590) );
  CLKBUFX3 U8813 ( .A(\i_MIPS/Register/n130 ), .Y(n5591) );
  CLKBUFX3 U8814 ( .A(\i_MIPS/Register/n129 ), .Y(n5588) );
  CLKBUFX3 U8815 ( .A(\i_MIPS/Register/n129 ), .Y(n5589) );
  CLKBUFX3 U8816 ( .A(\i_MIPS/Register/n128 ), .Y(n5586) );
  CLKBUFX3 U8817 ( .A(\i_MIPS/Register/n128 ), .Y(n5587) );
  CLKBUFX3 U8818 ( .A(\i_MIPS/Register/n127 ), .Y(n5584) );
  CLKBUFX3 U8819 ( .A(\i_MIPS/Register/n127 ), .Y(n5585) );
  CLKBUFX3 U8820 ( .A(\i_MIPS/Register/n126 ), .Y(n5582) );
  CLKBUFX3 U8821 ( .A(\i_MIPS/Register/n126 ), .Y(n5583) );
  CLKBUFX3 U8822 ( .A(\i_MIPS/Register/n125 ), .Y(n5580) );
  CLKBUFX3 U8823 ( .A(\i_MIPS/Register/n125 ), .Y(n5581) );
  CLKBUFX3 U8824 ( .A(\i_MIPS/Register/n124 ), .Y(n5578) );
  CLKBUFX3 U8825 ( .A(\i_MIPS/Register/n124 ), .Y(n5579) );
  CLKBUFX3 U8826 ( .A(\i_MIPS/Register/n123 ), .Y(n5576) );
  CLKBUFX3 U8827 ( .A(\i_MIPS/Register/n123 ), .Y(n5577) );
  CLKBUFX3 U8828 ( .A(\i_MIPS/Register/n121 ), .Y(n5574) );
  CLKBUFX3 U8829 ( .A(\i_MIPS/Register/n121 ), .Y(n5575) );
  CLKBUFX3 U8830 ( .A(\i_MIPS/Register/n112 ), .Y(n5566) );
  CLKBUFX3 U8831 ( .A(\i_MIPS/Register/n112 ), .Y(n5567) );
  CLKBUFX3 U8832 ( .A(\i_MIPS/Register/n108 ), .Y(n5562) );
  CLKBUFX3 U8833 ( .A(\i_MIPS/Register/n108 ), .Y(n5563) );
  CLKBUFX3 U8834 ( .A(\i_MIPS/Register/n106 ), .Y(n5560) );
  CLKBUFX3 U8835 ( .A(\i_MIPS/Register/n106 ), .Y(n5561) );
  CLKBUFX3 U8836 ( .A(\i_MIPS/Register/n116 ), .Y(n5570) );
  CLKBUFX3 U8837 ( .A(\i_MIPS/Register/n116 ), .Y(n5571) );
  CLKBUFX3 U8838 ( .A(\i_MIPS/Register/n114 ), .Y(n5568) );
  CLKBUFX3 U8839 ( .A(\i_MIPS/Register/n114 ), .Y(n5569) );
  CLKBUFX3 U8840 ( .A(\i_MIPS/Register/n110 ), .Y(n5564) );
  CLKBUFX3 U8841 ( .A(\i_MIPS/Register/n110 ), .Y(n5565) );
  CLKBUFX3 U8842 ( .A(n10865), .Y(n5467) );
  CLKBUFX3 U8843 ( .A(n10865), .Y(n5468) );
  CLKBUFX3 U8844 ( .A(\i_MIPS/Register/n118 ), .Y(n5572) );
  CLKBUFX3 U8845 ( .A(\i_MIPS/Register/n118 ), .Y(n5573) );
  CLKBUFX3 U8846 ( .A(n5957), .Y(n5969) );
  CLKBUFX3 U8847 ( .A(n5972), .Y(n5970) );
  CLKBUFX3 U8848 ( .A(rst_n), .Y(n5971) );
  AND2XL U8849 ( .A(n7694), .B(n3684), .Y(n7717) );
  AND2X2 U8850 ( .A(n7693), .B(n7692), .Y(n7714) );
  INVX12 U8851 ( .A(n4648), .Y(mem_addr_D[31]) );
  CLKINVX1 U8852 ( .A(n11507), .Y(n4650) );
  CLKINVX1 U8853 ( .A(n8440), .Y(n8441) );
  INVX12 U8854 ( .A(n4636), .Y(mem_addr_D[15]) );
  XOR2X1 U8855 ( .A(n10223), .B(n3783), .Y(n11110) );
  CLKMX2X2 U8856 ( .A(n6836), .B(n6835), .S0(net107812), .Y(net105194) );
  CLKMX2X2 U8857 ( .A(n7776), .B(n7775), .S0(net107812), .Y(net103416) );
  CLKMX2X2 U8858 ( .A(n8224), .B(n8223), .S0(net107810), .Y(n8226) );
  AOI2BB1X1 U8859 ( .A0N(net112332), .A1N(\i_MIPS/n355 ), .B0(n4526), .Y(n6853) );
  AOI2BB2X1 U8860 ( .B0(net111960), .B1(n9381), .A0N(net111906), .A1N(n10313), 
        .Y(n9400) );
  OA22X2 U8861 ( .A0(n4757), .A1(n656), .B0(n4793), .B1(n2237), .Y(n7197) );
  OA22X1 U8862 ( .A0(n4819), .A1(n1087), .B0(n4865), .B1(n2682), .Y(n8589) );
  CLKINVX1 U8863 ( .A(n7891), .Y(n7894) );
  INVX1 U8864 ( .A(net103060), .Y(net103224) );
  NAND2X1 U8865 ( .A(n4662), .B(\i_MIPS/n340 ), .Y(n8648) );
  OA22X1 U8866 ( .A0(n4817), .A1(n1232), .B0(n4863), .B1(n2773), .Y(n8981) );
  OA22X2 U8867 ( .A0(n4975), .A1(n795), .B0(n5020), .B1(n2358), .Y(n8188) );
  OA22X1 U8868 ( .A0(n4822), .A1(n1233), .B0(n4868), .B1(n2774), .Y(n8190) );
  OA22X1 U8869 ( .A0(n5101), .A1(n1234), .B0(n5066), .B1(n2775), .Y(n6007) );
  OA22X1 U8870 ( .A0(n5221), .A1(n1235), .B0(n5152), .B1(n2776), .Y(n6006) );
  OA22X1 U8871 ( .A0(n5221), .A1(n1236), .B0(n5178), .B1(n2777), .Y(n6002) );
  OA22X1 U8872 ( .A0(n5282), .A1(n1237), .B0(n5260), .B1(n2778), .Y(n6001) );
  OA22X1 U8873 ( .A0(n5194), .A1(n1239), .B0(n5153), .B1(n2780), .Y(n6046) );
  OA22X1 U8874 ( .A0(n5129), .A1(n1240), .B0(n5088), .B1(n2781), .Y(n6019) );
  OA22X1 U8875 ( .A0(n5211), .A1(n1241), .B0(n5147), .B1(n2782), .Y(n6018) );
  OA22X1 U8876 ( .A0(n5221), .A1(n1242), .B0(n5148), .B1(n2783), .Y(n6022) );
  OA22X1 U8877 ( .A0(n5212), .A1(n1243), .B0(n5170), .B1(n2784), .Y(n6098) );
  OA22X2 U8878 ( .A0(n5212), .A1(n1482), .B0(n5169), .B1(n3056), .Y(n10034) );
  OA22X2 U8879 ( .A0(n5386), .A1(n1483), .B0(n5346), .B1(n3057), .Y(n10032) );
  OA22X1 U8880 ( .A0(n5288), .A1(n1656), .B0(n5241), .B1(n3240), .Y(n6153) );
  OA22X1 U8881 ( .A0(n5196), .A1(n1657), .B0(n5152), .B1(n3241), .Y(n6154) );
  OA22X1 U8882 ( .A0(n5196), .A1(n1659), .B0(n5153), .B1(n3243), .Y(n6144) );
  OA22XL U8883 ( .A0(n5104), .A1(n1709), .B0(n5082), .B1(n3306), .Y(n6135) );
  OA22X1 U8884 ( .A0(n5288), .A1(n1661), .B0(n5241), .B1(n3245), .Y(n6148) );
  OA22X1 U8885 ( .A0(n5196), .A1(n1662), .B0(n5168), .B1(n3246), .Y(n6149) );
  OA22X1 U8886 ( .A0(n5120), .A1(n1663), .B0(n5062), .B1(n3247), .Y(n9961) );
  OA22X1 U8887 ( .A0(n5304), .A1(n1664), .B0(n5260), .B1(n3248), .Y(n10197) );
  OA22X1 U8888 ( .A0(n5222), .A1(n1665), .B0(n5172), .B1(n3249), .Y(n10198) );
  OA22X1 U8889 ( .A0(n230), .A1(n1666), .B0(n5260), .B1(n3250), .Y(n10184) );
  OA22X1 U8890 ( .A0(n5213), .A1(n1667), .B0(n5172), .B1(n3251), .Y(n10185) );
  OA22X1 U8891 ( .A0(n5304), .A1(n1668), .B0(n5260), .B1(n3252), .Y(n10180) );
  OA22X1 U8892 ( .A0(n5213), .A1(n1669), .B0(n5172), .B1(n3253), .Y(n10181) );
  OA22X1 U8893 ( .A0(n5205), .A1(n1088), .B0(n5161), .B1(n2731), .Y(n9754) );
  OA22X1 U8894 ( .A0(n5114), .A1(n1089), .B0(n5054), .B1(n2732), .Y(n9755) );
  OA22X1 U8895 ( .A0(n5369), .A1(n1090), .B0(n5340), .B1(n2733), .Y(n9752) );
  NAND4X1 U8896 ( .A(n10048), .B(n10047), .C(n10046), .D(n10045), .Y(n11260)
         );
  OA22X1 U8897 ( .A0(n5212), .A1(n1492), .B0(n5169), .B1(n3210), .Y(n10047) );
  OA22X1 U8898 ( .A0(n5121), .A1(n1493), .B0(n5075), .B1(n3211), .Y(n10048) );
  OA22X1 U8899 ( .A0(n5389), .A1(n1494), .B0(n5346), .B1(n3212), .Y(n10045) );
  OA22X1 U8900 ( .A0(n5201), .A1(n3061), .B0(n5157), .B1(n1170), .Y(n9607) );
  OA22X1 U8901 ( .A0(n5110), .A1(n3062), .B0(n5085), .B1(n1171), .Y(n9608) );
  OA22X1 U8902 ( .A0(n5399), .A1(n3063), .B0(n5337), .B1(n1172), .Y(n9605) );
  OA22X1 U8903 ( .A0(n5212), .A1(n1670), .B0(n5169), .B1(n3254), .Y(n10042) );
  OA22X1 U8904 ( .A0(n5121), .A1(n1495), .B0(n5078), .B1(n3255), .Y(n10043) );
  OA22X1 U8905 ( .A0(n5376), .A1(n1671), .B0(n5346), .B1(n3256), .Y(n10040) );
  OA22X1 U8906 ( .A0(n5212), .A1(n1496), .B0(n5169), .B1(n3257), .Y(n10052) );
  OA22X1 U8907 ( .A0(n5121), .A1(n1497), .B0(n5064), .B1(n3258), .Y(n10053) );
  OA22X1 U8908 ( .A0(n5377), .A1(n1498), .B0(n5346), .B1(n3259), .Y(n10050) );
  OA22X1 U8909 ( .A0(n5205), .A1(n1091), .B0(n5161), .B1(n2683), .Y(n9744) );
  OA22X1 U8910 ( .A0(n5114), .A1(n1092), .B0(n5087), .B1(n2684), .Y(n9745) );
  OA22X1 U8911 ( .A0(n5387), .A1(n1093), .B0(n5340), .B1(n2734), .Y(n9742) );
  OA22X1 U8912 ( .A0(n5201), .A1(n3064), .B0(n5157), .B1(n1173), .Y(n9597) );
  OA22X1 U8913 ( .A0(n5110), .A1(n1499), .B0(n5059), .B1(n3079), .Y(n9598) );
  OA22X1 U8914 ( .A0(n5206), .A1(n1094), .B0(n5162), .B1(n2685), .Y(n9777) );
  OA22X1 U8915 ( .A0(n5400), .A1(n1095), .B0(n5341), .B1(n2686), .Y(n9775) );
  OA22X1 U8916 ( .A0(n5374), .A1(n1096), .B0(n5340), .B1(n2735), .Y(n9738) );
  OA22X1 U8917 ( .A0(n5120), .A1(n1500), .B0(n5086), .B1(n3080), .Y(n9928) );
  OA22XL U8918 ( .A0(n5301), .A1(n1609), .B0(n5256), .B1(n3186), .Y(n9926) );
  OA22XL U8919 ( .A0(n5210), .A1(n1610), .B0(n5167), .B1(n3187), .Y(n9927) );
  OA22XL U8920 ( .A0(n5301), .A1(n1612), .B0(n5267), .B1(n3189), .Y(n9943) );
  OA22X1 U8921 ( .A0(n5205), .A1(n3065), .B0(n5161), .B1(n1277), .Y(n9749) );
  OA22X1 U8922 ( .A0(n5114), .A1(n3066), .B0(n5058), .B1(n1174), .Y(n9750) );
  OA22X1 U8923 ( .A0(n5392), .A1(n1097), .B0(n5340), .B1(n2736), .Y(n9747) );
  OA22X1 U8924 ( .A0(n5201), .A1(n1501), .B0(n5157), .B1(n3081), .Y(n9602) );
  OA22X1 U8925 ( .A0(n5110), .A1(n1502), .B0(n5084), .B1(n3082), .Y(n9603) );
  OA22X1 U8926 ( .A0(n237), .A1(n1503), .B0(n5337), .B1(n3083), .Y(n9600) );
  OA22X1 U8927 ( .A0(n5201), .A1(n1504), .B0(n5157), .B1(n3084), .Y(n9593) );
  OA22X1 U8928 ( .A0(n5377), .A1(n1505), .B0(n5337), .B1(n3085), .Y(n9591) );
  OA22X1 U8929 ( .A0(n5206), .A1(n1098), .B0(n5162), .B1(n2687), .Y(n9772) );
  OA22X1 U8930 ( .A0(n5115), .A1(n1099), .B0(n5068), .B1(n2688), .Y(n9773) );
  OA22X1 U8931 ( .A0(n5383), .A1(n1100), .B0(n5341), .B1(n2689), .Y(n9770) );
  OA22XL U8932 ( .A0(n5301), .A1(n1615), .B0(n5247), .B1(n3192), .Y(n9935) );
  OA22X1 U8933 ( .A0(n5209), .A1(n1506), .B0(n5166), .B1(n3086), .Y(n9917) );
  OA22X1 U8934 ( .A0(n5206), .A1(n1101), .B0(n5162), .B1(n2690), .Y(n9767) );
  OA22X1 U8935 ( .A0(n5115), .A1(n1102), .B0(n5085), .B1(n2691), .Y(n9768) );
  OA22X1 U8936 ( .A0(n5397), .A1(n1103), .B0(n5341), .B1(n2692), .Y(n9765) );
  OA22XL U8937 ( .A0(n5104), .A1(n1617), .B0(n5057), .B1(n3194), .Y(n6126) );
  OA22X1 U8938 ( .A0(n5300), .A1(n1507), .B0(n5255), .B1(n3087), .Y(n9911) );
  OA22X1 U8939 ( .A0(n5209), .A1(n1508), .B0(n5166), .B1(n3088), .Y(n9912) );
  OA22X1 U8940 ( .A0(n5300), .A1(n1672), .B0(n5255), .B1(n3260), .Y(n9903) );
  OA22X1 U8941 ( .A0(n5209), .A1(n1673), .B0(n5166), .B1(n3261), .Y(n9904) );
  OA22X1 U8942 ( .A0(n5373), .A1(n3067), .B0(n5341), .B1(n1175), .Y(n9761) );
  OA22X1 U8943 ( .A0(n5300), .A1(n1674), .B0(n5255), .B1(n3262), .Y(n9895) );
  OA22X1 U8944 ( .A0(n5209), .A1(n1675), .B0(n5166), .B1(n3263), .Y(n9896) );
  OA22X1 U8945 ( .A0(n5300), .A1(n1509), .B0(n5255), .B1(n3089), .Y(n9921) );
  OA22X1 U8946 ( .A0(n5209), .A1(n1510), .B0(n5166), .B1(n3090), .Y(n9922) );
  OA22XL U8947 ( .A0(n5104), .A1(n1710), .B0(n5087), .B1(n3307), .Y(n6130) );
  OA22X1 U8948 ( .A0(n5199), .A1(n1511), .B0(n5156), .B1(n3091), .Y(n6229) );
  OA22X1 U8949 ( .A0(n5108), .A1(n1512), .B0(n5055), .B1(n3092), .Y(n6230) );
  OA22X1 U8950 ( .A0(n5367), .A1(n1513), .B0(n5335), .B1(n3093), .Y(n6227) );
  OA22X1 U8951 ( .A0(n5198), .A1(n1514), .B0(n5155), .B1(n3094), .Y(n6219) );
  OA22X1 U8952 ( .A0(n5107), .A1(n1515), .B0(n5066), .B1(n3095), .Y(n6220) );
  OA22X1 U8953 ( .A0(n5380), .A1(n1516), .B0(n5334), .B1(n3096), .Y(n6217) );
  OA22X1 U8954 ( .A0(n5199), .A1(n1517), .B0(n5156), .B1(n3097), .Y(n6234) );
  OA22X1 U8955 ( .A0(n5108), .A1(n1518), .B0(n5077), .B1(n3098), .Y(n6235) );
  OA22X1 U8956 ( .A0(n5383), .A1(n1519), .B0(n5335), .B1(n3099), .Y(n6232) );
  NAND4X1 U8957 ( .A(n6225), .B(n6224), .C(n6223), .D(n6222), .Y(n11279) );
  OA22X1 U8958 ( .A0(n5198), .A1(n1520), .B0(n5155), .B1(n3100), .Y(n6224) );
  OA22X1 U8959 ( .A0(n5107), .A1(n1521), .B0(n5057), .B1(n3101), .Y(n6225) );
  OA22X1 U8960 ( .A0(n5381), .A1(n1522), .B0(n5334), .B1(n3102), .Y(n6222) );
  OA22X1 U8961 ( .A0(n5198), .A1(n1523), .B0(n5155), .B1(n3103), .Y(n6209) );
  OA22X1 U8962 ( .A0(n5107), .A1(n1524), .B0(n5081), .B1(n3104), .Y(n6210) );
  OA22X1 U8963 ( .A0(n5382), .A1(n1525), .B0(n5334), .B1(n3105), .Y(n6207) );
  OA22X1 U8964 ( .A0(n5107), .A1(n1526), .B0(n181), .B1(n3106), .Y(n6200) );
  OA22X1 U8965 ( .A0(n5390), .A1(n1527), .B0(n5334), .B1(n3107), .Y(n6197) );
  OA22X1 U8966 ( .A0(n5107), .A1(n1528), .B0(n5065), .B1(n3108), .Y(n6215) );
  NAND4X1 U8967 ( .A(n6205), .B(n6204), .C(n6203), .D(n6202), .Y(n11280) );
  OA22X1 U8968 ( .A0(n5107), .A1(n1530), .B0(n5074), .B1(n3110), .Y(n6205) );
  OA22X1 U8969 ( .A0(n5378), .A1(n1531), .B0(n5334), .B1(n3111), .Y(n6202) );
  OA22X1 U8970 ( .A0(n5289), .A1(n1104), .B0(n5242), .B1(n2693), .Y(n6168) );
  OA22X1 U8971 ( .A0(n5197), .A1(n1105), .B0(n5154), .B1(n2694), .Y(n6169) );
  NAND4X1 U8972 ( .A(n6160), .B(n6159), .C(n6158), .D(n6157), .Y(n11310) );
  OA22XL U8973 ( .A0(n5288), .A1(n1619), .B0(n5241), .B1(n3196), .Y(n6158) );
  OA22XL U8974 ( .A0(n5196), .A1(n1620), .B0(n5149), .B1(n3197), .Y(n6159) );
  OA22X1 U8975 ( .A0(n5106), .A1(n1106), .B0(n5068), .B1(n2695), .Y(n6175) );
  OA22X1 U8976 ( .A0(n5289), .A1(n1107), .B0(n5242), .B1(n2696), .Y(n6173) );
  OA22X1 U8977 ( .A0(n5197), .A1(n1108), .B0(n5154), .B1(n2697), .Y(n6174) );
  NAND4X1 U8978 ( .A(n6165), .B(n6164), .C(n6163), .D(n6162), .Y(n11278) );
  OA22XL U8979 ( .A0(n5288), .A1(n3112), .B0(n5241), .B1(n1202), .Y(n6163) );
  OA22XL U8980 ( .A0(n5196), .A1(n3113), .B0(n5165), .B1(n1203), .Y(n6164) );
  OA22X1 U8981 ( .A0(n5199), .A1(n1532), .B0(n5156), .B1(n3114), .Y(n6250) );
  OA22X1 U8982 ( .A0(n5108), .A1(n1533), .B0(n5071), .B1(n3115), .Y(n6251) );
  OA22X1 U8983 ( .A0(n5393), .A1(n1534), .B0(n5335), .B1(n3116), .Y(n6248) );
  NAND4X1 U8984 ( .A(n6243), .B(n6242), .C(n6241), .D(n6240), .Y(n11309) );
  OA22X1 U8985 ( .A0(n5199), .A1(n1535), .B0(n5156), .B1(n3117), .Y(n6242) );
  OA22X1 U8986 ( .A0(n5108), .A1(n1536), .B0(n5063), .B1(n3118), .Y(n6243) );
  NAND4X1 U8987 ( .A(n6255), .B(n6254), .C(n6253), .D(n6252), .Y(n11245) );
  OA22X1 U8988 ( .A0(n5199), .A1(n1538), .B0(n5156), .B1(n3120), .Y(n6254) );
  OA22X1 U8989 ( .A0(n5108), .A1(n1539), .B0(n5076), .B1(n3121), .Y(n6255) );
  OA22X1 U8990 ( .A0(n269), .A1(n1540), .B0(n5335), .B1(n3122), .Y(n6252) );
  NAND4X1 U8991 ( .A(n6247), .B(n6246), .C(n6245), .D(n6244), .Y(n11277) );
  OA22X1 U8992 ( .A0(n5199), .A1(n1541), .B0(n5156), .B1(n3123), .Y(n6246) );
  OA22X1 U8993 ( .A0(n5108), .A1(n1542), .B0(n5058), .B1(n3124), .Y(n6247) );
  OA22X1 U8994 ( .A0(n5394), .A1(n1543), .B0(n5335), .B1(n3125), .Y(n6244) );
  NAND4X1 U8995 ( .A(n6190), .B(n6189), .C(n6188), .D(n6187), .Y(n11217) );
  OA22X1 U8996 ( .A0(n5197), .A1(n1544), .B0(n5154), .B1(n3126), .Y(n6189) );
  OA22X1 U8997 ( .A0(n5106), .A1(n1545), .B0(n5086), .B1(n3127), .Y(n6190) );
  OA22X1 U8998 ( .A0(n5374), .A1(n1546), .B0(n5333), .B1(n3128), .Y(n6187) );
  OA22X1 U8999 ( .A0(n5197), .A1(n1547), .B0(n5154), .B1(n3129), .Y(n6179) );
  OA22X1 U9000 ( .A0(n5106), .A1(n1548), .B0(n5058), .B1(n3130), .Y(n6180) );
  OA22X1 U9001 ( .A0(n5369), .A1(n1549), .B0(n5333), .B1(n3131), .Y(n6177) );
  OA22X1 U9002 ( .A0(n5197), .A1(n1550), .B0(n5154), .B1(n3132), .Y(n6194) );
  OA22X1 U9003 ( .A0(n5106), .A1(n1551), .B0(n5062), .B1(n3133), .Y(n6195) );
  OA22X1 U9004 ( .A0(n5375), .A1(n1552), .B0(n5333), .B1(n3134), .Y(n6192) );
  NAND4X1 U9005 ( .A(n6185), .B(n6184), .C(n6183), .D(n6182), .Y(n11281) );
  OA22X1 U9006 ( .A0(n5197), .A1(n1553), .B0(n5154), .B1(n3135), .Y(n6184) );
  OA22X1 U9007 ( .A0(n5106), .A1(n1554), .B0(n5084), .B1(n3136), .Y(n6185) );
  OA22X1 U9008 ( .A0(n5401), .A1(n1555), .B0(n5333), .B1(n3137), .Y(n6182) );
  NAND4X1 U9009 ( .A(n6271), .B(n6270), .C(n6269), .D(n6268), .Y(n11212) );
  OA22X1 U9010 ( .A0(n5200), .A1(n1556), .B0(n5155), .B1(n3138), .Y(n6270) );
  OA22X1 U9011 ( .A0(n5109), .A1(n1557), .B0(n5070), .B1(n3139), .Y(n6271) );
  OA22X1 U9012 ( .A0(n5388), .A1(n1558), .B0(n5336), .B1(n3140), .Y(n6268) );
  NAND4X1 U9013 ( .A(n6263), .B(n6262), .C(n6261), .D(n6260), .Y(n11308) );
  OA22X1 U9014 ( .A0(n5200), .A1(n1455), .B0(n5154), .B1(n3141), .Y(n6262) );
  OA22X1 U9015 ( .A0(n5109), .A1(n1559), .B0(n5055), .B1(n3142), .Y(n6263) );
  OA22X1 U9016 ( .A0(n5379), .A1(n1560), .B0(n5336), .B1(n3143), .Y(n6260) );
  NAND4X1 U9017 ( .A(n6275), .B(n6274), .C(n6273), .D(n6272), .Y(n11244) );
  OA22X1 U9018 ( .A0(n5200), .A1(n1561), .B0(n5145), .B1(n3144), .Y(n6274) );
  OA22X1 U9019 ( .A0(n5109), .A1(n1562), .B0(n5060), .B1(n3145), .Y(n6275) );
  OA22X1 U9020 ( .A0(n5391), .A1(n1563), .B0(n5336), .B1(n3146), .Y(n6272) );
  NAND4X1 U9021 ( .A(n6267), .B(n6266), .C(n6265), .D(n6264), .Y(n11276) );
  OA22X1 U9022 ( .A0(n5200), .A1(n1564), .B0(n5155), .B1(n3147), .Y(n6266) );
  OA22X1 U9023 ( .A0(n5109), .A1(n1565), .B0(n5082), .B1(n3148), .Y(n6267) );
  OA22X1 U9024 ( .A0(n5371), .A1(n1566), .B0(n5336), .B1(n3149), .Y(n6264) );
  OA22X1 U9025 ( .A0(n5299), .A1(n1794), .B0(n5252), .B1(n3450), .Y(n9815) );
  OA22X1 U9026 ( .A0(n5207), .A1(n1795), .B0(n5163), .B1(n3451), .Y(n9816) );
  OA22X1 U9027 ( .A0(n5299), .A1(n1796), .B0(n5252), .B1(n3452), .Y(n9807) );
  OA22X1 U9028 ( .A0(n5207), .A1(n1797), .B0(n5163), .B1(n3453), .Y(n9808) );
  OA22X1 U9029 ( .A0(n5299), .A1(n1798), .B0(n5252), .B1(n3454), .Y(n9819) );
  OA22X1 U9030 ( .A0(n5207), .A1(n1799), .B0(n5163), .B1(n3455), .Y(n9820) );
  OA22X1 U9031 ( .A0(n5299), .A1(n1800), .B0(n5252), .B1(n3456), .Y(n9811) );
  OA22X1 U9032 ( .A0(n5207), .A1(n1801), .B0(n5163), .B1(n3457), .Y(n9812) );
  OA22X1 U9033 ( .A0(n5299), .A1(n1802), .B0(n5252), .B1(n3458), .Y(n9795) );
  OA22X1 U9034 ( .A0(n5207), .A1(n1803), .B0(n5163), .B1(n3459), .Y(n9796) );
  NAND4X1 U9035 ( .A(n9787), .B(n9786), .C(n9785), .D(n9784), .Y(n11306) );
  OA22XL U9036 ( .A0(n5115), .A1(n1871), .B0(n5056), .B1(n3527), .Y(n9787) );
  OA22XL U9037 ( .A0(n5206), .A1(n1872), .B0(n5162), .B1(n3528), .Y(n9786) );
  OA22X1 U9038 ( .A0(n5299), .A1(n1804), .B0(n5252), .B1(n3460), .Y(n9799) );
  OA22X1 U9039 ( .A0(n5207), .A1(n1805), .B0(n5163), .B1(n3461), .Y(n9800) );
  NAND4X1 U9040 ( .A(n9792), .B(n9791), .C(n9790), .D(n9789), .Y(n11274) );
  OA22XL U9041 ( .A0(n5115), .A1(n1873), .B0(n167), .B1(n3529), .Y(n9792) );
  OA22XL U9042 ( .A0(n5206), .A1(n1874), .B0(n5162), .B1(n3530), .Y(n9791) );
  OA22X1 U9043 ( .A0(n5299), .A1(n1806), .B0(n5253), .B1(n3462), .Y(n9835) );
  OA22X1 U9044 ( .A0(n5208), .A1(n1807), .B0(n5164), .B1(n3463), .Y(n9836) );
  OA22X1 U9045 ( .A0(n5299), .A1(n1808), .B0(n5253), .B1(n3464), .Y(n9827) );
  OA22X1 U9046 ( .A0(n5208), .A1(n1809), .B0(n5164), .B1(n3465), .Y(n9828) );
  OA22X1 U9047 ( .A0(n5299), .A1(n1810), .B0(n5253), .B1(n3466), .Y(n9839) );
  OA22X1 U9048 ( .A0(n5208), .A1(n1811), .B0(n5164), .B1(n3467), .Y(n9840) );
  OA22X1 U9049 ( .A0(n5299), .A1(n1812), .B0(n5253), .B1(n3468), .Y(n9831) );
  OA22X1 U9050 ( .A0(n5208), .A1(n1813), .B0(n5164), .B1(n3469), .Y(n9832) );
  OA22X1 U9051 ( .A0(n5299), .A1(n1814), .B0(n5254), .B1(n3470), .Y(n9871) );
  OA22X1 U9052 ( .A0(n5207), .A1(n3589), .B0(n5165), .B1(n1875), .Y(n9872) );
  OA22X1 U9053 ( .A0(n5299), .A1(n1935), .B0(n5254), .B1(n3591), .Y(n9863) );
  OA22X1 U9054 ( .A0(n5208), .A1(n1936), .B0(n5165), .B1(n3592), .Y(n9864) );
  OA22X1 U9055 ( .A0(n5299), .A1(n1815), .B0(n5254), .B1(n3471), .Y(n9875) );
  OA22X1 U9056 ( .A0(n5207), .A1(n1816), .B0(n5165), .B1(n3472), .Y(n9876) );
  OA22X1 U9057 ( .A0(n5299), .A1(n1817), .B0(n5254), .B1(n3473), .Y(n9867) );
  OA22X1 U9058 ( .A0(n5207), .A1(n1818), .B0(n5165), .B1(n3474), .Y(n9868) );
  OA22X1 U9059 ( .A0(n5299), .A1(n1819), .B0(n5254), .B1(n3475), .Y(n9855) );
  OA22X1 U9060 ( .A0(n5208), .A1(n1820), .B0(n5165), .B1(n3476), .Y(n9856) );
  OA22X1 U9061 ( .A0(n5299), .A1(n1821), .B0(n5253), .B1(n3477), .Y(n9847) );
  OA22X1 U9062 ( .A0(n5208), .A1(n1822), .B0(n5164), .B1(n3478), .Y(n9848) );
  OA22X1 U9063 ( .A0(n5299), .A1(n1823), .B0(n5254), .B1(n3479), .Y(n9859) );
  OA22X1 U9064 ( .A0(n5208), .A1(n1824), .B0(n5165), .B1(n3480), .Y(n9860) );
  OA22X1 U9065 ( .A0(n5299), .A1(n1825), .B0(n5253), .B1(n3481), .Y(n9851) );
  OA22X1 U9066 ( .A0(n5208), .A1(n1826), .B0(n5164), .B1(n3482), .Y(n9852) );
  NAND4X1 U9067 ( .A(n9628), .B(n9627), .C(n9626), .D(n9625), .Y(n11206) );
  OA22XL U9068 ( .A0(n5111), .A1(n1876), .B0(n5087), .B1(n3531), .Y(n9628) );
  OA22XL U9069 ( .A0(n230), .A1(n1877), .B0(n5247), .B1(n3532), .Y(n9626) );
  OA22XL U9070 ( .A0(n5202), .A1(n1878), .B0(n183), .B1(n3533), .Y(n9627) );
  NAND4X1 U9071 ( .A(n9618), .B(n9617), .C(n9616), .D(n9615), .Y(n11302) );
  OA22XL U9072 ( .A0(n5111), .A1(n1879), .B0(n5089), .B1(n3534), .Y(n9618) );
  OA22XL U9073 ( .A0(n230), .A1(n1880), .B0(n5247), .B1(n3535), .Y(n9616) );
  OA22XL U9074 ( .A0(n5202), .A1(n1881), .B0(n183), .B1(n3536), .Y(n9617) );
  NAND4X1 U9075 ( .A(n9633), .B(n9632), .C(n9631), .D(n9630), .Y(n11238) );
  OA22XL U9076 ( .A0(n5111), .A1(n1882), .B0(n5063), .B1(n3537), .Y(n9633) );
  OA22XL U9077 ( .A0(n230), .A1(n1883), .B0(n5247), .B1(n3538), .Y(n9631) );
  OA22XL U9078 ( .A0(n5202), .A1(n1884), .B0(n183), .B1(n3539), .Y(n9632) );
  NAND4X1 U9079 ( .A(n9623), .B(n9622), .C(n9621), .D(n9620), .Y(n11270) );
  OA22XL U9080 ( .A0(n5111), .A1(n1885), .B0(n5073), .B1(n3540), .Y(n9623) );
  OA22XL U9081 ( .A0(n230), .A1(n1886), .B0(n5247), .B1(n3541), .Y(n9621) );
  OA22XL U9082 ( .A0(n5202), .A1(n1887), .B0(n183), .B1(n3542), .Y(n9622) );
  NAND4X1 U9083 ( .A(n9582), .B(n9581), .C(n9580), .D(n9579), .Y(n11205) );
  OA22XL U9084 ( .A0(n5110), .A1(n1888), .B0(n5077), .B1(n3543), .Y(n9582) );
  OA22XL U9085 ( .A0(n5201), .A1(n1889), .B0(n5157), .B1(n3544), .Y(n9581) );
  NAND4X1 U9086 ( .A(n9574), .B(n9573), .C(n9572), .D(n9571), .Y(n11301) );
  NAND4X1 U9087 ( .A(n9586), .B(n9585), .C(n9584), .D(n9583), .Y(n11237) );
  OA22XL U9088 ( .A0(n5110), .A1(n1890), .B0(n5059), .B1(n3545), .Y(n9586) );
  OA22XL U9089 ( .A0(n5201), .A1(n1891), .B0(n5157), .B1(n3546), .Y(n9585) );
  NAND4X1 U9090 ( .A(n9578), .B(n9577), .C(n9576), .D(n9575), .Y(n11269) );
  NAND4X1 U9091 ( .A(n9677), .B(n9676), .C(n9675), .D(n9674), .Y(n11204) );
  OA22XL U9092 ( .A0(n5112), .A1(n1892), .B0(n5079), .B1(n3547), .Y(n9677) );
  NAND4X1 U9093 ( .A(n9667), .B(n9666), .C(n9665), .D(n9664), .Y(n11300) );
  OA22XL U9094 ( .A0(n5112), .A1(n1893), .B0(n5080), .B1(n3548), .Y(n9667) );
  NAND4X1 U9095 ( .A(n9682), .B(n9681), .C(n9680), .D(n9679), .Y(n11236) );
  OA22XL U9096 ( .A0(n5112), .A1(n1894), .B0(n5061), .B1(n3549), .Y(n9682) );
  NAND4X1 U9097 ( .A(n9672), .B(n9671), .C(n9670), .D(n9669), .Y(n11268) );
  OA22XL U9098 ( .A0(n5112), .A1(n1895), .B0(n5086), .B1(n3550), .Y(n9672) );
  OA22X1 U9099 ( .A0(n5203), .A1(n1827), .B0(n5159), .B1(n3483), .Y(n9671) );
  NAND4X1 U9100 ( .A(n10166), .B(n10165), .C(n10164), .D(n10163), .Y(n11203)
         );
  OA22XL U9101 ( .A0(n5123), .A1(n1896), .B0(n5068), .B1(n3551), .Y(n10166) );
  OA22X1 U9102 ( .A0(n5304), .A1(n1828), .B0(n5259), .B1(n3484), .Y(n10164) );
  OA22XL U9103 ( .A0(n5214), .A1(n1897), .B0(n5171), .B1(n3552), .Y(n10165) );
  NAND4X1 U9104 ( .A(n10156), .B(n10155), .C(n10154), .D(n10153), .Y(n11299)
         );
  OA22XL U9105 ( .A0(n5123), .A1(n1898), .B0(n5089), .B1(n3553), .Y(n10156) );
  OA22X1 U9106 ( .A0(n5304), .A1(n1829), .B0(n5259), .B1(n3485), .Y(n10154) );
  OA22XL U9107 ( .A0(n5214), .A1(n1899), .B0(n5171), .B1(n3554), .Y(n10155) );
  NAND4X1 U9108 ( .A(n10171), .B(n10170), .C(n10169), .D(n10168), .Y(n11235)
         );
  OA22XL U9109 ( .A0(n5124), .A1(n1900), .B0(n167), .B1(n3555), .Y(n10171) );
  OA22XL U9110 ( .A0(n5299), .A1(n1901), .B0(n5260), .B1(n3556), .Y(n10169) );
  OA22XL U9111 ( .A0(n5207), .A1(n1902), .B0(n5172), .B1(n3557), .Y(n10170) );
  NAND4X1 U9112 ( .A(n10161), .B(n10160), .C(n10159), .D(n10158), .Y(n11267)
         );
  OA22XL U9113 ( .A0(n5123), .A1(n1903), .B0(n5085), .B1(n3558), .Y(n10161) );
  OA22X1 U9114 ( .A0(n5304), .A1(n1830), .B0(n5259), .B1(n3486), .Y(n10159) );
  OA22XL U9115 ( .A0(n5214), .A1(n1904), .B0(n5171), .B1(n3559), .Y(n10160) );
  NAND4X1 U9116 ( .A(n9726), .B(n9725), .C(n9724), .D(n9723), .Y(n11202) );
  OA22XL U9117 ( .A0(n5114), .A1(n1905), .B0(n5057), .B1(n3560), .Y(n9726) );
  OA22XL U9118 ( .A0(n5205), .A1(n1906), .B0(n5161), .B1(n3561), .Y(n9725) );
  NAND4X1 U9119 ( .A(n9716), .B(n9715), .C(n9714), .D(n9713), .Y(n11298) );
  OA22XL U9120 ( .A0(n5113), .A1(n1907), .B0(n5088), .B1(n3562), .Y(n9716) );
  OA22XL U9121 ( .A0(n5204), .A1(n1908), .B0(n5160), .B1(n3563), .Y(n9715) );
  NAND4X1 U9122 ( .A(n9731), .B(n9730), .C(n9729), .D(n9728), .Y(n11234) );
  OA22XL U9123 ( .A0(n5114), .A1(n1909), .B0(n5062), .B1(n3564), .Y(n9731) );
  OA22XL U9124 ( .A0(n5205), .A1(n1910), .B0(n5161), .B1(n3565), .Y(n9730) );
  NAND4X1 U9125 ( .A(n9721), .B(n9720), .C(n9719), .D(n9718), .Y(n11266) );
  OA22XL U9126 ( .A0(n5113), .A1(n1911), .B0(n5088), .B1(n3566), .Y(n9721) );
  OA22XL U9127 ( .A0(n5204), .A1(n1912), .B0(n5160), .B1(n3567), .Y(n9720) );
  OA22XL U9128 ( .A0(n4986), .A1(n1391), .B0(n5032), .B1(n2921), .Y(n6432) );
  OA22XL U9129 ( .A0(n4761), .A1(n3265), .B0(n4795), .B1(n1425), .Y(n6435) );
  OA22XL U9130 ( .A0(n4986), .A1(n1392), .B0(n5032), .B1(n2922), .Y(n6428) );
  OA22X2 U9131 ( .A0(n4975), .A1(n799), .B0(n5020), .B1(n2362), .Y(n8104) );
  OA22X2 U9132 ( .A0(n4973), .A1(n703), .B0(n5011), .B1(n2271), .Y(n9390) );
  OA22X2 U9133 ( .A0(n4982), .A1(n667), .B0(n5028), .B1(n2238), .Y(n7016) );
  OA22X2 U9134 ( .A0(n4758), .A1(n2292), .B0(n4794), .B1(n675), .Y(n7019) );
  OA22X2 U9135 ( .A0(n4979), .A1(n802), .B0(n5024), .B1(n2365), .Y(n7657) );
  OA22X2 U9136 ( .A0(n4826), .A1(n803), .B0(n4871), .B1(n2366), .Y(n7659) );
  OA22X2 U9137 ( .A0(n4753), .A1(n657), .B0(n4792), .B1(n2240), .Y(n7660) );
  OA22XL U9138 ( .A0(n4837), .A1(n1176), .B0(n4883), .B1(n2726), .Y(n6323) );
  OA22XL U9139 ( .A0(n4765), .A1(n2785), .B0(n4796), .B1(n1126), .Y(n6324) );
  OA22X2 U9140 ( .A0(n4971), .A1(n705), .B0(n5013), .B1(n2273), .Y(n9299) );
  OA22X2 U9141 ( .A0(n4813), .A1(n669), .B0(n4863), .B1(n2241), .Y(n9301) );
  OA22X2 U9142 ( .A0(n4976), .A1(n804), .B0(n185), .B1(n2367), .Y(n8021) );
  OA22X2 U9143 ( .A0(n4974), .A1(n670), .B0(n5019), .B1(n2242), .Y(n8309) );
  OA22X2 U9144 ( .A0(n4821), .A1(n671), .B0(n4867), .B1(n2243), .Y(n8311) );
  OA22X2 U9145 ( .A0(n4748), .A1(n658), .B0(n4790), .B1(n2244), .Y(n8312) );
  OA22X2 U9146 ( .A0(n4978), .A1(n806), .B0(n5025), .B1(n2369), .Y(n7437) );
  OA22X2 U9147 ( .A0(n4755), .A1(n659), .B0(n4793), .B1(n2245), .Y(n7440) );
  OA22X2 U9148 ( .A0(n4830), .A1(n672), .B0(n4861), .B1(n2246), .Y(n9090) );
  OA22X2 U9149 ( .A0(n4743), .A1(n2293), .B0(n4789), .B1(n676), .Y(n9091) );
  OA22X2 U9150 ( .A0(n4973), .A1(n811), .B0(n5018), .B1(n2374), .Y(n8400) );
  OA22X2 U9151 ( .A0(n4820), .A1(n812), .B0(n4866), .B1(n2375), .Y(n8402) );
  OA22X2 U9152 ( .A0(n4748), .A1(n813), .B0(n4790), .B1(n2376), .Y(n8403) );
  OA22X2 U9153 ( .A0(n4833), .A1(n673), .B0(n4878), .B1(n2247), .Y(n6655) );
  OA22XL U9154 ( .A0(n4761), .A1(n2737), .B0(n4795), .B1(n1138), .Y(n6656) );
  OA22X2 U9155 ( .A0(n4983), .A1(n814), .B0(n5029), .B1(n2377), .Y(n7008) );
  OA22X2 U9156 ( .A0(n4758), .A1(n816), .B0(n4794), .B1(n2379), .Y(n7011) );
  OA22X2 U9157 ( .A0(n4746), .A1(n2413), .B0(n4790), .B1(n677), .Y(n8602) );
  OA22X2 U9158 ( .A0(n4995), .A1(n706), .B0(n5018), .B1(n2274), .Y(n9295) );
  OA22X2 U9159 ( .A0(n4814), .A1(n707), .B0(n4859), .B1(n2275), .Y(n9297) );
  OA22XL U9160 ( .A0(n4837), .A1(n1177), .B0(n4883), .B1(n2727), .Y(n6319) );
  OA22XL U9161 ( .A0(n4765), .A1(n2976), .B0(n4796), .B1(n1204), .Y(n6320) );
  OA22X2 U9162 ( .A0(n4749), .A1(n817), .B0(n4791), .B1(n2380), .Y(n8304) );
  OA22X2 U9163 ( .A0(n4743), .A1(n2415), .B0(n4789), .B1(n729), .Y(n9083) );
  OA22X2 U9164 ( .A0(n4997), .A1(n818), .B0(n5029), .B1(n2381), .Y(n9510) );
  OA22X2 U9165 ( .A0(n4810), .A1(n819), .B0(n4856), .B1(n2382), .Y(n9512) );
  OA22X2 U9166 ( .A0(n4985), .A1(n710), .B0(n5031), .B1(n2278), .Y(n6645) );
  OA22X2 U9167 ( .A0(n4833), .A1(n711), .B0(n4878), .B1(n2279), .Y(n6647) );
  OA22XL U9168 ( .A0(n4761), .A1(n2977), .B0(n4795), .B1(n1205), .Y(n6648) );
  OA22X1 U9169 ( .A0(n4819), .A1(n1244), .B0(n4865), .B1(n2786), .Y(n8597) );
  OA22X1 U9170 ( .A0(n4832), .A1(n1245), .B0(n4877), .B1(n2787), .Y(n6890) );
  OA22X1 U9171 ( .A0(n4833), .A1(n1246), .B0(n4878), .B1(n2788), .Y(n6651) );
  OA22XL U9172 ( .A0(n4761), .A1(n1393), .B0(n4795), .B1(n2923), .Y(n6652) );
  OA22X2 U9173 ( .A0(n4975), .A1(n824), .B0(n5020), .B1(n2387), .Y(n8195) );
  OA22X1 U9174 ( .A0(n4822), .A1(n1247), .B0(n4868), .B1(n2789), .Y(n8197) );
  OA22X2 U9175 ( .A0(n4977), .A1(n826), .B0(n5022), .B1(n2389), .Y(n7845) );
  OA22X2 U9176 ( .A0(n4752), .A1(n827), .B0(n4792), .B1(n2390), .Y(n7848) );
  OA22X1 U9177 ( .A0(n4819), .A1(n1110), .B0(n4865), .B1(n2699), .Y(n8593) );
  OA22X2 U9178 ( .A0(n4747), .A1(n851), .B0(n4790), .B1(n2421), .Y(n8594) );
  OA22X1 U9179 ( .A0(n4832), .A1(n1249), .B0(n4877), .B1(n2791), .Y(n6809) );
  OA22XL U9180 ( .A0(n4760), .A1(n1178), .B0(n4795), .B1(n2925), .Y(n6810) );
  OA22X2 U9181 ( .A0(n4985), .A1(n829), .B0(n5031), .B1(n2392), .Y(n6799) );
  OA22X1 U9182 ( .A0(n4833), .A1(n1250), .B0(n4878), .B1(n2792), .Y(n6801) );
  OA22XL U9183 ( .A0(n4760), .A1(n3266), .B0(n4795), .B1(n1426), .Y(n6802) );
  OA22XL U9184 ( .A0(n5212), .A1(n1395), .B0(n5150), .B1(n2926), .Y(n6070) );
  OA22XL U9185 ( .A0(n5287), .A1(n1396), .B0(n5255), .B1(n2927), .Y(n6069) );
  OA22XL U9186 ( .A0(n5102), .A1(n1397), .B0(n5076), .B1(n2928), .Y(n6067) );
  OA22XL U9187 ( .A0(n5194), .A1(n1398), .B0(n5150), .B1(n2929), .Y(n6066) );
  OA22XL U9188 ( .A0(n5286), .A1(n1399), .B0(n5239), .B1(n2930), .Y(n6065) );
  OA22XL U9189 ( .A0(n5102), .A1(n1400), .B0(n167), .B1(n2931), .Y(n6039) );
  OA22XL U9190 ( .A0(n5194), .A1(n1401), .B0(n5150), .B1(n2932), .Y(n6038) );
  OA22XL U9191 ( .A0(n5286), .A1(n1402), .B0(n5239), .B1(n2933), .Y(n6037) );
  OA22X1 U9192 ( .A0(n5221), .A1(n1252), .B0(n5150), .B1(n2794), .Y(n6034) );
  OA22XL U9193 ( .A0(n5102), .A1(n1403), .B0(n5057), .B1(n2934), .Y(n6059) );
  OA22XL U9194 ( .A0(n5194), .A1(n1404), .B0(n5148), .B1(n2935), .Y(n6058) );
  OA22XL U9195 ( .A0(n5286), .A1(n1405), .B0(n5239), .B1(n2936), .Y(n6057) );
  OA22XL U9196 ( .A0(n5102), .A1(n1406), .B0(n5071), .B1(n2937), .Y(n6055) );
  OA22XL U9197 ( .A0(n5194), .A1(n1407), .B0(n5169), .B1(n2938), .Y(n6054) );
  OA22XL U9198 ( .A0(n5286), .A1(n1408), .B0(n5239), .B1(n2939), .Y(n6053) );
  OA22XL U9199 ( .A0(n5194), .A1(n1410), .B0(n5151), .B1(n2941), .Y(n6050) );
  OA22XL U9200 ( .A0(n5286), .A1(n1411), .B0(n5239), .B1(n2942), .Y(n6049) );
  OA22X1 U9201 ( .A0(n5122), .A1(n1253), .B0(n5056), .B1(n2795), .Y(n6027) );
  OA22X1 U9202 ( .A0(n5221), .A1(n1254), .B0(n5149), .B1(n2796), .Y(n6026) );
  OA22X1 U9203 ( .A0(n5309), .A1(n1255), .B0(n5266), .B1(n2797), .Y(n6025) );
  OA22XL U9204 ( .A0(n5103), .A1(n1135), .B0(n5075), .B1(n2671), .Y(n6091) );
  OA22XL U9205 ( .A0(n5220), .A1(n1136), .B0(n5153), .B1(n2672), .Y(n6090) );
  OA22XL U9206 ( .A0(n5220), .A1(n1412), .B0(n5170), .B1(n2943), .Y(n6086) );
  OA22XL U9207 ( .A0(n5103), .A1(n1413), .B0(n167), .B1(n2944), .Y(n6083) );
  OA22XL U9208 ( .A0(n5220), .A1(n1414), .B0(n5151), .B1(n2945), .Y(n6082) );
  OA22XL U9209 ( .A0(n5103), .A1(n1415), .B0(n5068), .B1(n2946), .Y(n6079) );
  OA22XL U9210 ( .A0(n5220), .A1(n1416), .B0(n5168), .B1(n2947), .Y(n6078) );
  OA22XL U9211 ( .A0(n5104), .A1(n1417), .B0(n5075), .B1(n2948), .Y(n6102) );
  OAI222XL U9212 ( .A0(n5467), .A1(n266), .B0(n5424), .B1(n5466), .C0(n5558), 
        .C1(\i_MIPS/n205 ), .Y(n11523) );
  OAI222XL U9213 ( .A0(n5467), .A1(n272), .B0(n5433), .B1(n5464), .C0(n5558), 
        .C1(\i_MIPS/n202 ), .Y(n11526) );
  OAI222XL U9214 ( .A0(n5467), .A1(n282), .B0(n2211), .B1(n5465), .C0(n5559), 
        .C1(\i_MIPS/n199 ), .Y(n11529) );
  OAI222XL U9215 ( .A0(n5468), .A1(n267), .B0(n5406), .B1(n5465), .C0(n5559), 
        .C1(\i_MIPS/n209 ), .Y(n11519) );
  OAI222XL U9216 ( .A0(n5467), .A1(n304), .B0(n1999), .B1(n5465), .C0(n5559), 
        .C1(\i_MIPS/n208 ), .Y(n11520) );
  OAI222XL U9217 ( .A0(n5467), .A1(n271), .B0(n1987), .B1(n5464), .C0(n5558), 
        .C1(\i_MIPS/n207 ), .Y(n11521) );
  OAI222XL U9218 ( .A0(n5467), .A1(n308), .B0(n1978), .B1(n5466), .C0(n5558), 
        .C1(\i_MIPS/n206 ), .Y(n11522) );
  OAI222XL U9219 ( .A0(n5467), .A1(n311), .B0(n1985), .B1(n5464), .C0(n5558), 
        .C1(\i_MIPS/n204 ), .Y(n11524) );
  OAI222XL U9220 ( .A0(n5467), .A1(n305), .B0(n1980), .B1(n5464), .C0(n5558), 
        .C1(\i_MIPS/n203 ), .Y(n11525) );
  OAI222XL U9221 ( .A0(n5467), .A1(n418), .B0(n5418), .B1(n5466), .C0(n5559), 
        .C1(\i_MIPS/n201 ), .Y(n11527) );
  OAI222XL U9222 ( .A0(n5467), .A1(n279), .B0(n1988), .B1(n5466), .C0(n5558), 
        .C1(\i_MIPS/n200 ), .Y(n11528) );
  OAI222XL U9223 ( .A0(n5467), .A1(n312), .B0(n1996), .B1(n5466), .C0(n5559), 
        .C1(\i_MIPS/n198 ), .Y(n11530) );
  OAI222XL U9224 ( .A0(n5467), .A1(n273), .B0(n4437), .B1(n5466), .C0(n5559), 
        .C1(\i_MIPS/n197 ), .Y(n11531) );
  OAI222XL U9225 ( .A0(n5467), .A1(n283), .B0(n4479), .B1(n5466), .C0(n5559), 
        .C1(\i_MIPS/n196 ), .Y(n11532) );
  OAI222XL U9226 ( .A0(n5467), .A1(n419), .B0(n5450), .B1(n5466), .C0(n5559), 
        .C1(\i_MIPS/n195 ), .Y(n11533) );
  OAI222XL U9227 ( .A0(n5468), .A1(n313), .B0(n1989), .B1(n5465), .C0(n5559), 
        .C1(\i_MIPS/n194 ), .Y(n11534) );
  OAI222XL U9228 ( .A0(n5468), .A1(n314), .B0(n1990), .B1(n5465), .C0(n5559), 
        .C1(\i_MIPS/n193 ), .Y(n11535) );
  OAI222XL U9229 ( .A0(n5467), .A1(n276), .B0(n1991), .B1(n5464), .C0(n5558), 
        .C1(\i_MIPS/n192 ), .Y(n11536) );
  OAI222XL U9230 ( .A0(n5467), .A1(n309), .B0(n1997), .B1(n5466), .C0(n5559), 
        .C1(\i_MIPS/n191 ), .Y(n11537) );
  OAI222XL U9231 ( .A0(n5467), .A1(n280), .B0(n1992), .B1(n5466), .C0(n5558), 
        .C1(\i_MIPS/n190 ), .Y(n11538) );
  OAI222XL U9232 ( .A0(n5468), .A1(n317), .B0(n5044), .B1(n5465), .C0(n5558), 
        .C1(\i_MIPS/n189 ), .Y(n11539) );
  OAI222XL U9233 ( .A0(n5468), .A1(n277), .B0(n5492), .B1(n5465), .C0(n5559), 
        .C1(\i_MIPS/n188 ), .Y(n11540) );
  OAI222XL U9234 ( .A0(n5468), .A1(n310), .B0(n1986), .B1(n5465), .C0(n5558), 
        .C1(\i_MIPS/n187 ), .Y(n11541) );
  OAI222XL U9235 ( .A0(n5468), .A1(n268), .B0(n2000), .B1(n5465), .C0(n5558), 
        .C1(\i_MIPS/n186 ), .Y(n11542) );
  OAI222XL U9236 ( .A0(n5468), .A1(n316), .B0(n1979), .B1(n5465), .C0(n5559), 
        .C1(\i_MIPS/n185 ), .Y(n11543) );
  OAI222XL U9237 ( .A0(n5468), .A1(n281), .B0(n5478), .B1(n5466), .C0(n5558), 
        .C1(\i_MIPS/n184 ), .Y(n11544) );
  OAI222XL U9238 ( .A0(n5468), .A1(n315), .B0(n1994), .B1(n5466), .C0(n5558), 
        .C1(\i_MIPS/n183 ), .Y(n11545) );
  OA22X2 U9239 ( .A0(n4811), .A1(n715), .B0(n263), .B1(n2283), .Y(n9388) );
  OA22X2 U9240 ( .A0(n4742), .A1(n2418), .B0(n4788), .B1(n733), .Y(n9389) );
  OA22X2 U9241 ( .A0(n4968), .A1(n830), .B0(n5014), .B1(n2393), .Y(n9382) );
  OA22X2 U9242 ( .A0(n4812), .A1(n831), .B0(n4858), .B1(n2394), .Y(n9384) );
  OA22X2 U9243 ( .A0(n4754), .A1(n832), .B0(n4788), .B1(n2395), .Y(n9385) );
  OA22XL U9244 ( .A0(n4837), .A1(n1179), .B0(n4883), .B1(n2728), .Y(n6315) );
  OA22XL U9245 ( .A0(n4765), .A1(n2978), .B0(n4796), .B1(n1206), .Y(n6316) );
  OA22X2 U9246 ( .A0(n4979), .A1(n716), .B0(n5025), .B1(n2284), .Y(n6299) );
  OA22X2 U9247 ( .A0(n4817), .A1(n717), .B0(n4875), .B1(n2285), .Y(n6301) );
  OA22X1 U9248 ( .A0(n4751), .A1(n2956), .B0(n4788), .B1(n1180), .Y(n6302) );
  OA22X2 U9249 ( .A0(n4976), .A1(n833), .B0(n185), .B1(n2396), .Y(n8009) );
  OA22X2 U9250 ( .A0(n4974), .A1(n835), .B0(n5019), .B1(n2398), .Y(n8297) );
  OA22X1 U9251 ( .A0(n4821), .A1(n1256), .B0(n4867), .B1(n2798), .Y(n8299) );
  OA22X2 U9252 ( .A0(n4749), .A1(n836), .B0(n4791), .B1(n2399), .Y(n8300) );
  OA22X2 U9253 ( .A0(n4980), .A1(n837), .B0(n5025), .B1(n2400), .Y(n7425) );
  OA22X2 U9254 ( .A0(n4755), .A1(n838), .B0(n4793), .B1(n2401), .Y(n7428) );
  OA22X2 U9255 ( .A0(n4758), .A1(n2419), .B0(n4794), .B1(n734), .Y(n7092) );
  OA22X1 U9256 ( .A0(n4819), .A1(n1258), .B0(n4865), .B1(n2800), .Y(n8686) );
  OA22X2 U9257 ( .A0(n4981), .A1(n841), .B0(n5027), .B1(n2404), .Y(n7182) );
  OA22X1 U9258 ( .A0(n4829), .A1(n1259), .B0(n4874), .B1(n2801), .Y(n7184) );
  OA22X2 U9259 ( .A0(n4757), .A1(n842), .B0(n4793), .B1(n2405), .Y(n7185) );
  OA22X2 U9260 ( .A0(n4985), .A1(n720), .B0(n5031), .B1(n2288), .Y(n6641) );
  OA22XL U9261 ( .A0(n4761), .A1(n2979), .B0(n4795), .B1(n1207), .Y(n6644) );
  OA22X2 U9262 ( .A0(n4981), .A1(n843), .B0(n5010), .B1(n2406), .Y(n9500) );
  OA22X1 U9263 ( .A0(n4825), .A1(n1260), .B0(n4861), .B1(n2802), .Y(n9502) );
  NAND2X1 U9264 ( .A(n11180), .B(\i_MIPS/n341 ), .Y(n6705) );
  OA22X1 U9265 ( .A0(n5288), .A1(n1678), .B0(n5241), .B1(n3268), .Y(n6138) );
  OA22X1 U9266 ( .A0(n5196), .A1(n1679), .B0(n5152), .B1(n3269), .Y(n6139) );
  OA22X2 U9267 ( .A0(n5111), .A1(n1484), .B0(n5079), .B1(n3058), .Y(n9642) );
  OA22X2 U9268 ( .A0(n5202), .A1(n3031), .B0(n183), .B1(n1447), .Y(n9641) );
  AO22X2 U9269 ( .A0(n5528), .A1(DCACHE_addr[29]), .B0(n5526), .B1(n11507), 
        .Y(n11018) );
  AO22X2 U9270 ( .A0(n5528), .A1(DCACHE_addr[19]), .B0(n5527), .B1(n11497), 
        .Y(n11040) );
  AO22X2 U9271 ( .A0(n5528), .A1(DCACHE_addr[6]), .B0(n5527), .B1(n11484), .Y(
        n11038) );
  AO22X2 U9272 ( .A0(n5528), .A1(DCACHE_addr[9]), .B0(n5527), .B1(n11487), .Y(
        n11027) );
  AO22X2 U9273 ( .A0(n5528), .A1(DCACHE_addr[25]), .B0(n5526), .B1(n11503), 
        .Y(n11026) );
  AO22X2 U9274 ( .A0(n5528), .A1(DCACHE_addr[22]), .B0(n5527), .B1(n11500), 
        .Y(n11028) );
  OA22XL U9275 ( .A0(n5104), .A1(n1729), .B0(n5081), .B1(n3336), .Y(n6118) );
  NOR4X1 U9276 ( .A(n6472), .B(n6471), .C(n6470), .D(n6469), .Y(n6473) );
  NOR4X1 U9277 ( .A(n6463), .B(n6462), .C(n6461), .D(n6460), .Y(n6464) );
  NOR4X1 U9278 ( .A(n6617), .B(n6616), .C(n6615), .D(n6614), .Y(n6618) );
  NOR4X1 U9279 ( .A(n9098), .B(n9097), .C(n9096), .D(n9095), .Y(n9099) );
  NOR4X1 U9280 ( .A(n8571), .B(n8570), .C(n8569), .D(n8568), .Y(n8572) );
  NOR4X1 U9281 ( .A(n9539), .B(n9538), .C(n9537), .D(n9536), .Y(n9540) );
  NOR4X1 U9282 ( .A(n9519), .B(n9518), .C(n9517), .D(n9516), .Y(n9520) );
  AO22X1 U9283 ( .A0(n9531), .A1(n994), .B0(n4714), .B1(n2518), .Y(n9316) );
  AO22X1 U9284 ( .A0(n4713), .A1(n281), .B0(n4707), .B1(n2519), .Y(n8040) );
  AO22X1 U9285 ( .A0(n9531), .A1(n995), .B0(n4717), .B1(n2520), .Y(n8039) );
  AO22X1 U9286 ( .A0(n4722), .A1(n996), .B0(n4719), .B1(n2521), .Y(n8038) );
  AO22X1 U9287 ( .A0(n4713), .A1(n947), .B0(n4710), .B1(n2459), .Y(n9308) );
  AO22X1 U9288 ( .A0(n9531), .A1(n997), .B0(n4715), .B1(n2522), .Y(n9307) );
  NOR4X1 U9289 ( .A(n8123), .B(n8122), .C(n8121), .D(n8120), .Y(n8124) );
  AO22X1 U9290 ( .A0(n4711), .A1(n282), .B0(n4708), .B1(n2523), .Y(n8123) );
  AO22X1 U9291 ( .A0(n9531), .A1(n998), .B0(n4717), .B1(n2524), .Y(n8122) );
  AO22X1 U9292 ( .A0(n4711), .A1(n999), .B0(n4708), .B1(n2525), .Y(n8031) );
  AO22X1 U9293 ( .A0(n9531), .A1(n1000), .B0(n4717), .B1(n2526), .Y(n8030) );
  AO22X1 U9294 ( .A0(n4722), .A1(n1001), .B0(n4719), .B1(n2527), .Y(n8029) );
  AO22X1 U9295 ( .A0(n9531), .A1(n393), .B0(n4716), .B1(n1042), .Y(n7675) );
  AO22X1 U9296 ( .A0(n4712), .A1(n283), .B0(n4708), .B1(n2460), .Y(n7770) );
  AO22X1 U9297 ( .A0(n9531), .A1(n1002), .B0(n4717), .B1(n2528), .Y(n7769) );
  NOR4X1 U9298 ( .A(n8114), .B(n8113), .C(n8112), .D(n8111), .Y(n8115) );
  AO22X1 U9299 ( .A0(n4713), .A1(n1003), .B0(n4708), .B1(n2529), .Y(n8114) );
  AO22X1 U9300 ( .A0(n9531), .A1(n1004), .B0(n4717), .B1(n2530), .Y(n8113) );
  AO22X1 U9301 ( .A0(n4712), .A1(n436), .B0(n4708), .B1(n2461), .Y(n7667) );
  NOR4X1 U9302 ( .A(n6955), .B(n6954), .C(n6953), .D(n6952), .Y(n6956) );
  AO22X1 U9303 ( .A0(n4711), .A1(n316), .B0(n4707), .B1(n2462), .Y(n6955) );
  AO22X1 U9304 ( .A0(n9531), .A1(n1005), .B0(n4715), .B1(n2531), .Y(n6954) );
  AO22X1 U9305 ( .A0(n4721), .A1(n948), .B0(n4719), .B1(n2463), .Y(n6953) );
  AO22X1 U9306 ( .A0(n4711), .A1(n949), .B0(n4709), .B1(n2464), .Y(n7761) );
  AO22X1 U9307 ( .A0(n9531), .A1(n1006), .B0(n4717), .B1(n2532), .Y(n7760) );
  AO22X1 U9308 ( .A0(n4711), .A1(n317), .B0(n4707), .B1(n2465), .Y(n7035) );
  AO22X1 U9309 ( .A0(n9531), .A1(n950), .B0(n4715), .B1(n2466), .Y(n7034) );
  AO22X1 U9310 ( .A0(n4721), .A1(n951), .B0(n4719), .B1(n2467), .Y(n7033) );
  NOR4X1 U9311 ( .A(n6946), .B(n6945), .C(n6944), .D(n6943), .Y(n6947) );
  AO22X1 U9312 ( .A0(n4711), .A1(n952), .B0(n4707), .B1(n2468), .Y(n6946) );
  AO22X1 U9313 ( .A0(n9531), .A1(n1007), .B0(n4715), .B1(n2533), .Y(n6945) );
  AO22X1 U9314 ( .A0(n4721), .A1(n953), .B0(n4719), .B1(n2469), .Y(n6944) );
  AO22X1 U9315 ( .A0(n4711), .A1(n954), .B0(n4707), .B1(n2470), .Y(n7026) );
  AO22X1 U9316 ( .A0(n9531), .A1(n955), .B0(n4715), .B1(n2471), .Y(n7025) );
  AO22X1 U9317 ( .A0(n4721), .A1(n956), .B0(n4719), .B1(n2472), .Y(n7024) );
  NOR4X1 U9318 ( .A(n8509), .B(n8508), .C(n8507), .D(n8506), .Y(n8510) );
  NOR4X1 U9319 ( .A(n7447), .B(n7446), .C(n7445), .D(n7444), .Y(n7448) );
  NOR4X1 U9320 ( .A(n8319), .B(n8318), .C(n8317), .D(n8316), .Y(n8320) );
  NOR4X1 U9321 ( .A(n8909), .B(n8908), .C(n8907), .D(n8906), .Y(n8910) );
  AO22X1 U9322 ( .A0(n4713), .A1(n272), .B0(n4709), .B1(n2004), .Y(n8620) );
  AO22X1 U9323 ( .A0(n9531), .A1(n318), .B0(n4714), .B1(n2005), .Y(n8619) );
  NOR4X1 U9324 ( .A(n8611), .B(n8610), .C(n8609), .D(n8608), .Y(n8612) );
  AO22X1 U9325 ( .A0(n4712), .A1(n425), .B0(n4709), .B1(n2006), .Y(n8611) );
  AO22X1 U9326 ( .A0(n9531), .A1(n319), .B0(n4714), .B1(n2007), .Y(n8610) );
  NOR4X1 U9327 ( .A(n7286), .B(n7285), .C(n7284), .D(n7283), .Y(n7287) );
  NOR4X1 U9328 ( .A(n6830), .B(n6829), .C(n6828), .D(n6827), .Y(n6831) );
  NOR4X1 U9329 ( .A(n6821), .B(n6820), .C(n6819), .D(n6818), .Y(n6822) );
  NOR4X1 U9330 ( .A(n8715), .B(n8714), .C(n8713), .D(n8712), .Y(n8716) );
  NOR4X1 U9331 ( .A(n7375), .B(n7374), .C(n7373), .D(n7372), .Y(n7376) );
  NOR4X1 U9332 ( .A(n7213), .B(n7212), .C(n7211), .D(n7210), .Y(n7214) );
  NOR4X1 U9333 ( .A(n9010), .B(n9009), .C(n9008), .D(n9007), .Y(n9011) );
  NOR4X1 U9334 ( .A(n6911), .B(n6910), .C(n6909), .D(n6908), .Y(n6912) );
  NOR4X1 U9335 ( .A(n7366), .B(n7365), .C(n7364), .D(n7363), .Y(n7367) );
  NOR4X1 U9336 ( .A(n7204), .B(n7203), .C(n7202), .D(n7201), .Y(n7205) );
  NOR4X1 U9337 ( .A(n9001), .B(n9000), .C(n8999), .D(n8998), .Y(n9002) );
  NOR4X1 U9338 ( .A(n6902), .B(n6901), .C(n6900), .D(n6899), .Y(n6903) );
  NOR4X1 U9339 ( .A(n8808), .B(n8807), .C(n8806), .D(n8805), .Y(n8809) );
  NAND2XL U9340 ( .A(n7688), .B(n7523), .Y(n7417) );
  NAND2XL U9341 ( .A(n7610), .B(n7609), .Y(n7614) );
  NAND2XL U9342 ( .A(n7803), .B(n7617), .Y(n7611) );
  NAND2XL U9343 ( .A(n8341), .B(n8360), .Y(n8342) );
  CLKINVX1 U9344 ( .A(n8236), .Y(n7491) );
  NAND2X1 U9345 ( .A(n8970), .B(n9347), .Y(n8179) );
  NOR4X1 U9346 ( .A(n9409), .B(n9408), .C(n9407), .D(n9406), .Y(n9428) );
  NAND4X1 U9347 ( .A(n9404), .B(n9403), .C(n9402), .D(n9401), .Y(n9409) );
  AO22X1 U9348 ( .A0(n4696), .A1(n285), .B0(n4477), .B1(n430), .Y(n9407) );
  AO22X1 U9349 ( .A0(n4482), .A1(n274), .B0(n4705), .B1(n306), .Y(n9406) );
  NOR4X1 U9350 ( .A(n9426), .B(n9425), .C(n9424), .D(n9423), .Y(n9427) );
  NAND4X1 U9351 ( .A(n9421), .B(n9420), .C(n9419), .D(n9418), .Y(n9426) );
  AO22X1 U9352 ( .A0(n4696), .A1(n286), .B0(n4477), .B1(n431), .Y(n9424) );
  AO22X1 U9353 ( .A0(n4482), .A1(n275), .B0(n4705), .B1(n307), .Y(n9423) );
  NAND2X1 U9354 ( .A(DCACHE_addr[23]), .B(n4674), .Y(n10489) );
  OAI211X1 U9355 ( .A0(n9334), .A1(n8555), .B0(n8554), .C0(n4658), .Y(n8556)
         );
  NAND2XL U9356 ( .A(n6598), .B(\i_MIPS/n341 ), .Y(n6708) );
  NAND2X1 U9357 ( .A(DCACHE_addr[2]), .B(n4673), .Y(net99164) );
  INVXL U9358 ( .A(n10542), .Y(n10543) );
  INVXL U9359 ( .A(n10449), .Y(n10450) );
  NAND2X1 U9360 ( .A(DCACHE_addr[20]), .B(n4674), .Y(n10222) );
  INVX1 U9361 ( .A(n7880), .Y(n7517) );
  NAND2X2 U9362 ( .A(n4662), .B(net107808), .Y(n8353) );
  NAND2X1 U9363 ( .A(DCACHE_addr[25]), .B(n4674), .Y(n10313) );
  AOI2BB1XL U9364 ( .A0N(n7475), .A1N(\i_MIPS/n371 ), .B0(n4298), .Y(n7476) );
  CLKINVX1 U9365 ( .A(n10627), .Y(n10505) );
  NAND2XL U9366 ( .A(n7881), .B(n7880), .Y(n7888) );
  OA22XL U9367 ( .A0(net112368), .A1(\i_MIPS/n355 ), .B0(net112350), .B1(
        \i_MIPS/n356 ), .Y(n6765) );
  NAND2X1 U9368 ( .A(n6707), .B(n6705), .Y(n6599) );
  AND3X2 U9369 ( .A(n3907), .B(n7481), .C(n6708), .Y(n6602) );
  NAND2XL U9370 ( .A(n8849), .B(n8848), .Y(n8857) );
  NAND2X1 U9371 ( .A(DCACHE_addr[1]), .B(n2651), .Y(n10078) );
  CLKINVX1 U9372 ( .A(n11180), .Y(n6598) );
  NAND2XL U9373 ( .A(n9487), .B(n9152), .Y(n9150) );
  NAND2XL U9374 ( .A(n9476), .B(n9475), .Y(n9494) );
  NAND2XL U9375 ( .A(n9348), .B(n9347), .Y(n9356) );
  NAND2XL U9376 ( .A(n9263), .B(n9262), .Y(n9283) );
  CLKMX2X2 U9377 ( .A(net100573), .B(net112438), .S0(n7974), .Y(n7987) );
  NAND2XL U9378 ( .A(net112376), .B(\i_MIPS/n357 ), .Y(n7824) );
  NAND2XL U9379 ( .A(n8072), .B(n8071), .Y(n8075) );
  NAND2XL U9380 ( .A(n8553), .B(n8546), .Y(n8544) );
  NAND2XL U9381 ( .A(n9043), .B(n9042), .Y(n9069) );
  NAND2XL U9382 ( .A(n8750), .B(n8752), .Y(n7808) );
  CLKINVX1 U9383 ( .A(n8848), .Y(n8861) );
  NAND2X1 U9384 ( .A(n8444), .B(n8432), .Y(n8451) );
  INVXL U9385 ( .A(n10823), .Y(n10824) );
  INVXL U9386 ( .A(n10622), .Y(n10623) );
  NAND2X1 U9387 ( .A(n9159), .B(n8864), .Y(n8869) );
  NAND2XL U9388 ( .A(n11012), .B(n11011), .Y(n11499) );
  NAND2XL U9389 ( .A(n11015), .B(n11014), .Y(n11494) );
  NOR2X1 U9390 ( .A(n6719), .B(n6718), .Y(n6730) );
  NAND2XL U9391 ( .A(n4064), .B(n3359), .Y(n11495) );
  INVXL U9392 ( .A(n8947), .Y(n9064) );
  AND2X2 U9393 ( .A(n10374), .B(n10375), .Y(n4453) );
  OA22X2 U9394 ( .A0(n4978), .A1(n844), .B0(n5023), .B1(n2407), .Y(n7751) );
  OA22X1 U9395 ( .A0(n4825), .A1(n1261), .B0(n4870), .B1(n2803), .Y(n7753) );
  OA22X1 U9396 ( .A0(n4825), .A1(n1262), .B0(n4870), .B1(n2804), .Y(n7741) );
  OA22X1 U9397 ( .A0(n4753), .A1(n2957), .B0(n4792), .B1(n1278), .Y(n7742) );
  OA22X1 U9398 ( .A0(n4979), .A1(n1263), .B0(n5024), .B1(n2805), .Y(n7646) );
  OA22X1 U9399 ( .A0(n4826), .A1(n1264), .B0(n4871), .B1(n2806), .Y(n7648) );
  OA22X1 U9400 ( .A0(n4754), .A1(n2958), .B0(n4792), .B1(n1181), .Y(n7649) );
  OA22X1 U9401 ( .A0(n4981), .A1(n1265), .B0(n5027), .B1(n2807), .Y(n7264) );
  OA22X1 U9402 ( .A0(n4829), .A1(n1266), .B0(n4874), .B1(n2808), .Y(n7266) );
  OA22X1 U9403 ( .A0(n4756), .A1(n1077), .B0(n4793), .B1(n2809), .Y(n7267) );
  OA22X1 U9404 ( .A0(n4830), .A1(n1112), .B0(n4861), .B1(n2701), .Y(n9183) );
  OA22X1 U9405 ( .A0(n4824), .A1(n1267), .B0(n4869), .B1(n2810), .Y(n7933) );
  OA22X1 U9406 ( .A0(n4752), .A1(n1268), .B0(n4792), .B1(n2811), .Y(n7934) );
  OA22X1 U9407 ( .A0(n4971), .A1(n1269), .B0(n5016), .B1(n2812), .Y(n8786) );
  OA22X1 U9408 ( .A0(n4818), .A1(n1270), .B0(n263), .B1(n2813), .Y(n8788) );
  OA22X1 U9409 ( .A0(n4980), .A1(n1271), .B0(n5026), .B1(n2814), .Y(n7344) );
  OA22X1 U9410 ( .A0(n4828), .A1(n1272), .B0(n4873), .B1(n2815), .Y(n7346) );
  OA22XL U9411 ( .A0(n4825), .A1(n1418), .B0(n4870), .B1(n2949), .Y(n7839) );
  OA22XL U9412 ( .A0(n4752), .A1(n1182), .B0(n4792), .B1(n2950), .Y(n7840) );
  INVXL U9413 ( .A(n9152), .Y(n9486) );
  NAND2XL U9414 ( .A(n3685), .B(n6844), .Y(n6845) );
  INVXL U9415 ( .A(n8546), .Y(n9276) );
  CLKMX2X2 U9416 ( .A(n9452), .B(n9451), .S0(\i_MIPS/IR_ID[25] ), .Y(n9499) );
  NOR4X1 U9417 ( .A(n9441), .B(n9440), .C(n9439), .D(n9438), .Y(n9452) );
  CLKMX2X2 U9418 ( .A(n8149), .B(n8148), .S0(\i_MIPS/IR_ID[25] ), .Y(n8187) );
  NOR4X1 U9419 ( .A(n8138), .B(n8137), .C(n8136), .D(n8135), .Y(n8149) );
  NOR4X1 U9420 ( .A(n9125), .B(n9124), .C(n9123), .D(n9122), .Y(n9136) );
  CLKMX2X2 U9421 ( .A(n8386), .B(n8385), .S0(\i_MIPS/IR_ID[25] ), .Y(n8387) );
  NOR4X1 U9422 ( .A(n8375), .B(n8374), .C(n8373), .D(n8372), .Y(n8386) );
  CLKMX2X2 U9423 ( .A(n8484), .B(n8483), .S0(\i_MIPS/IR_ID[25] ), .Y(n8485) );
  NOR4X1 U9424 ( .A(n8473), .B(n8472), .C(n8471), .D(n8470), .Y(n8484) );
  NOR4X1 U9425 ( .A(n7388), .B(n7387), .C(n7386), .D(n7385), .Y(n7399) );
  NOR4X1 U9426 ( .A(n7076), .B(n7075), .C(n7074), .D(n7073), .Y(n7087) );
  NOR4X1 U9427 ( .A(n8055), .B(n8054), .C(n8053), .D(n8052), .Y(n8066) );
  CLKMX2X2 U9428 ( .A(n9039), .B(n9038), .S0(\i_MIPS/IR_ID[25] ), .Y(n9074) );
  NOR4X1 U9429 ( .A(n9028), .B(n9027), .C(n9026), .D(n9025), .Y(n9039) );
  NOR4X1 U9430 ( .A(n7135), .B(n7134), .C(n7133), .D(n7132), .Y(n7146) );
  NOR4X1 U9431 ( .A(n7560), .B(n7559), .C(n7558), .D(n7557), .Y(n7571) );
  NOR4X1 U9432 ( .A(n7785), .B(n7784), .C(n7783), .D(n7782), .Y(n7796) );
  CLKMX2X2 U9433 ( .A(n8682), .B(n8681), .S0(\i_MIPS/IR_ID[25] ), .Y(n8683) );
  CLKMX2X2 U9434 ( .A(n7003), .B(n7002), .S0(net107816), .Y(n7004) );
  NOR4X1 U9435 ( .A(n6992), .B(n6991), .C(n6990), .D(n6989), .Y(n7003) );
  CLKMX2X2 U9436 ( .A(n6878), .B(n6877), .S0(\i_MIPS/IR_ID[25] ), .Y(n6879) );
  NOR4X1 U9437 ( .A(n6867), .B(n6866), .C(n6865), .D(n6864), .Y(n6878) );
  CLKMX2X2 U9438 ( .A(n8784), .B(n8783), .S0(net107816), .Y(n8785) );
  NOR4X1 U9439 ( .A(n8773), .B(n8772), .C(n8771), .D(n8770), .Y(n8784) );
  CLKMX2X2 U9440 ( .A(n6797), .B(n6796), .S0(\i_MIPS/IR_ID[25] ), .Y(n6798) );
  NOR4X1 U9441 ( .A(n6786), .B(n6785), .C(n6784), .D(n6783), .Y(n6797) );
  NOR4X1 U9442 ( .A(n8836), .B(n8835), .C(n8834), .D(n8833), .Y(n8847) );
  NAND2XL U9443 ( .A(n7891), .B(n7902), .Y(n7885) );
  NAND2XL U9444 ( .A(n8636), .B(n8635), .Y(n7057) );
  CLKINVX1 U9445 ( .A(n11183), .Y(n7482) );
  AND2X2 U9446 ( .A(n9041), .B(n8955), .Y(n6522) );
  NAND2XL U9447 ( .A(n7492), .B(n7496), .Y(n7312) );
  NAND2BX1 U9448 ( .AN(n8239), .B(n8854), .Y(n8246) );
  INVXL U9449 ( .A(n10324), .Y(n10253) );
  CLKINVX1 U9450 ( .A(n9329), .Y(n7480) );
  NAND2XL U9451 ( .A(n4), .B(n7975), .Y(n7979) );
  NAND2XL U9452 ( .A(n6964), .B(n6966), .Y(n6761) );
  NAND2XL U9453 ( .A(n7877), .B(n7876), .Y(n6972) );
  NAND2XL U9454 ( .A(n7502), .B(n4381), .Y(n6764) );
  NAND2X1 U9455 ( .A(DCACHE_addr[19]), .B(n4674), .Y(n10563) );
  CLKINVX1 U9456 ( .A(n6605), .Y(n9886) );
  MX2XL U9457 ( .A(\i_MIPS/n366 ), .B(n7696), .S0(\i_MIPS/ID_EX[79] ), .Y(
        n8358) );
  NAND2XL U9458 ( .A(n4305), .B(n7406), .Y(n7309) );
  NOR4X1 U9459 ( .A(n8927), .B(n8926), .C(n8925), .D(n8924), .Y(n8938) );
  AO21X2 U9460 ( .A0(n10322), .A1(n4610), .B0(net111902), .Y(n10355) );
  CLKMX2X2 U9461 ( .A(n7061), .B(n7042), .S0(net107796), .Y(n7420) );
  INVXL U9462 ( .A(n8752), .Y(n7819) );
  MXI2X1 U9463 ( .A(n8549), .B(n8548), .S0(net107794), .Y(n4471) );
  MX2XL U9464 ( .A(n3358), .B(n7149), .S0(\i_MIPS/ID_EX[79] ), .Y(n8156) );
  MX2XL U9465 ( .A(n7149), .B(\i_MIPS/n344 ), .S0(\i_MIPS/ID_EX[79] ), .Y(
        n8440) );
  MX2XL U9466 ( .A(\i_MIPS/n368 ), .B(\i_MIPS/n367 ), .S0(\i_MIPS/ID_EX[79] ), 
        .Y(n8357) );
  AND2X2 U9467 ( .A(n10806), .B(n10804), .Y(n4475) );
  NAND4BX1 U9468 ( .AN(n8615), .B(n8614), .C(n8613), .D(n8612), .Y(n8626) );
  INVXL U9469 ( .A(n8751), .Y(n8748) );
  CLKINVX1 U9470 ( .A(n6707), .Y(n6710) );
  CLKMX2X2 U9471 ( .A(n9545), .B(n9544), .S0(net107810), .Y(n9548) );
  CLKMX2X2 U9472 ( .A(n8425), .B(n8424), .S0(net107810), .Y(n8428) );
  CLKMX2X2 U9473 ( .A(n8295), .B(n8294), .S0(\i_MIPS/IR_ID[25] ), .Y(n8296) );
  NOR4X1 U9474 ( .A(n8284), .B(n8283), .C(n8282), .D(n8281), .Y(n8295) );
  CLKBUFX3 U9475 ( .A(net107808), .Y(net107802) );
  NAND3BX2 U9476 ( .AN(n8856), .B(n9457), .C(n8855), .Y(n8860) );
  CLKINVX1 U9477 ( .A(n9059), .Y(n8652) );
  CLKINVX1 U9478 ( .A(net103914), .Y(net103911) );
  AND2X2 U9479 ( .A(n4501), .B(n4448), .Y(n4478) );
  CLKINVX1 U9480 ( .A(n10506), .Y(n5418) );
  NAND2XL U9481 ( .A(n10504), .B(n10503), .Y(n10506) );
  NOR2BX1 U9482 ( .AN(net98375), .B(n4480), .Y(n4479) );
  INVXL U9483 ( .A(n10521), .Y(n4480) );
  CLKINVX1 U9484 ( .A(n10718), .Y(n5450) );
  MX2XL U9485 ( .A(net101082), .B(net112415), .S0(n4481), .Y(n7465) );
  NAND2XL U9486 ( .A(n7464), .B(\i_MIPS/n371 ), .Y(n4481) );
  INVX1 U9487 ( .A(n8727), .Y(n8540) );
  NAND4XL U9488 ( .A(n9457), .B(n9268), .C(n9243), .D(n8071), .Y(n7530) );
  MX2XL U9489 ( .A(DCACHE_addr[19]), .B(n10665), .S0(n210), .Y(\i_MIPS/n448 )
         );
  MX2XL U9490 ( .A(DCACHE_addr[1]), .B(n10965), .S0(n213), .Y(\i_MIPS/n466 )
         );
  MX2XL U9491 ( .A(DCACHE_addr[28]), .B(n258), .S0(n217), .Y(\i_MIPS/n439 ) );
  AO22X1 U9492 ( .A0(n145), .A1(n321), .B0(n227), .B1(n429), .Y(n8568) );
  AO22X1 U9493 ( .A0(n145), .A1(n426), .B0(n229), .B1(n2008), .Y(n6469) );
  AO22X1 U9494 ( .A0(n145), .A1(n427), .B0(n228), .B1(n2009), .Y(n6460) );
  AO22X1 U9495 ( .A0(n4729), .A1(n320), .B0(n4725), .B1(n428), .Y(n8617) );
  AO22X1 U9496 ( .A0(n4729), .A1(n321), .B0(n4727), .B1(n429), .Y(n8608) );
  INVXL U9497 ( .A(n9475), .Y(n9458) );
  MX2XL U9498 ( .A(n4664), .B(net97703), .S0(n207), .Y(\i_MIPS/n464 ) );
  MX2XL U9499 ( .A(DCACHE_addr[4]), .B(net97684), .S0(n216), .Y(\i_MIPS/n463 )
         );
  MX2XL U9500 ( .A(DCACHE_addr[2]), .B(net97770), .S0(n211), .Y(\i_MIPS/n465 )
         );
  INVX1 U9501 ( .A(n9459), .Y(n9155) );
  INVXL U9502 ( .A(n9262), .Y(n9244) );
  CLKMX2X2 U9503 ( .A(\i_MIPS/PHT_2/history_state[1] ), .B(
        \i_MIPS/PHT_2/history_state[0] ), .S0(n11045), .Y(\i_MIPS/PHT_2/n53 )
         );
  MX2XL U9504 ( .A(DCACHE_addr[7]), .B(n10693), .S0(n217), .Y(\i_MIPS/n460 )
         );
  MX2XL U9505 ( .A(DCACHE_addr[20]), .B(n20), .S0(n204), .Y(\i_MIPS/n447 ) );
  MX2XL U9506 ( .A(DCACHE_addr[13]), .B(net98012), .S0(n223), .Y(\i_MIPS/n454 ) );
  AND2X2 U9507 ( .A(n7510), .B(n4381), .Y(n7512) );
  INVXL U9508 ( .A(n7509), .Y(n7510) );
  NAND2XL U9509 ( .A(n6531), .B(\i_MIPS/n364 ), .Y(n4483) );
  MX2XL U9510 ( .A(DCACHE_addr[25]), .B(n3689), .S0(n207), .Y(\i_MIPS/n442 )
         );
  MX2XL U9511 ( .A(DCACHE_addr[8]), .B(net98393), .S0(n214), .Y(\i_MIPS/n459 )
         );
  MX2XL U9512 ( .A(DCACHE_addr[27]), .B(n3830), .S0(n205), .Y(\i_MIPS/n440 )
         );
  AND2XL U9513 ( .A(net103910), .B(n9329), .Y(n7547) );
  NOR4X1 U9514 ( .A(n7252), .B(n7251), .C(n7250), .D(n7249), .Y(n7263) );
  INVXL U9515 ( .A(\i_MIPS/forward_unit/n10 ), .Y(n6633) );
  CLKBUFX3 U9516 ( .A(n10195), .Y(n5312) );
  NAND3BX1 U9517 ( .AN(n9567), .B(n9887), .C(\i_MIPS/n324 ), .Y(
        \i_MIPS/Control_ID/n10 ) );
  NAND2X1 U9518 ( .A(\i_MIPS/n322 ), .B(\i_MIPS/n332 ), .Y(n9891) );
  CLKINVX1 U9519 ( .A(n4651), .Y(n11314) );
  NOR2BX1 U9520 ( .AN(n4544), .B(n9567), .Y(n4487) );
  AND2X2 U9521 ( .A(n4487), .B(\i_MIPS/n332 ), .Y(n4488) );
  CLKINVX1 U9522 ( .A(n11046), .Y(n11065) );
  CLKBUFX3 U9523 ( .A(n5967), .Y(n5972) );
  MXI2X2 U9524 ( .A(n10875), .B(n10874), .S0(n5520), .Y(n10876) );
  AOI222XL U9525 ( .A0(n5504), .A1(n11380), .B0(mem_rdata_D[30]), .B1(n232), 
        .C0(n12957), .C1(n5501), .Y(n10146) );
  MXI2X2 U9526 ( .A(n10688), .B(n10687), .S0(n5517), .Y(n10689) );
  MXI2X2 U9527 ( .A(n10308), .B(n10307), .S0(n5514), .Y(n10309) );
  MXI2X2 U9528 ( .A(n10276), .B(n10275), .S0(n5514), .Y(n10277) );
  MXI2X2 U9529 ( .A(n10498), .B(n10497), .S0(n5514), .Y(n10499) );
  MXI2X2 U9530 ( .A(n10783), .B(n10782), .S0(n5519), .Y(n10784) );
  MXI2X2 U9531 ( .A(n10661), .B(n10660), .S0(n5516), .Y(n10662) );
  MXI2X2 U9532 ( .A(n10515), .B(n10514), .S0(n5516), .Y(n10516) );
  AOI222XL U9533 ( .A0(n5504), .A1(n11368), .B0(mem_rdata_D[18]), .B1(n233), 
        .C0(n12969), .C1(n5501), .Y(n10515) );
  MXI2X2 U9534 ( .A(n10770), .B(n10769), .S0(n5519), .Y(n10771) );
  AOI222XL U9535 ( .A0(n5504), .A1(n11366), .B0(mem_rdata_D[16]), .B1(n233), 
        .C0(n12971), .C1(n5501), .Y(n10295) );
  MXI2X2 U9536 ( .A(n10759), .B(n10758), .S0(n5519), .Y(n10760) );
  AOI222XL U9537 ( .A0(n5505), .A1(n11362), .B0(mem_rdata_D[12]), .B1(n234), 
        .C0(n12975), .C1(n5502), .Y(n10726) );
  AOI222XL U9538 ( .A0(n5505), .A1(n11361), .B0(mem_rdata_D[11]), .B1(n235), 
        .C0(n12976), .C1(n5502), .Y(n10714) );
  MXI2X2 U9539 ( .A(n10080), .B(n10079), .S0(n5513), .Y(n10081) );
  AOI222XL U9540 ( .A0(n5503), .A1(n11373), .B0(mem_rdata_D[23]), .B1(n236), 
        .C0(n12964), .C1(n5502), .Y(n10947) );
  MXI2X2 U9541 ( .A(n10973), .B(n10972), .S0(n5522), .Y(n10974) );
  MXI2X2 U9542 ( .A(n10935), .B(n10934), .S0(n5521), .Y(n10936) );
  NAND2XL U9543 ( .A(n12931), .B(\i_MIPS/n336 ), .Y(n10322) );
  NAND2XL U9544 ( .A(n12933), .B(n4674), .Y(n10282) );
  NAND2XL U9545 ( .A(n12952), .B(n4674), .Y(net98335) );
  AOI222XL U9546 ( .A0(n5499), .A1(n11445), .B0(mem_rdata_D[95]), .B1(n232), 
        .C0(n12956), .C1(n5497), .Y(n10872) );
  AOI222XL U9547 ( .A0(n5498), .A1(n11441), .B0(mem_rdata_D[91]), .B1(n232), 
        .C0(n12960), .C1(n4385), .Y(n10305) );
  MXI2X2 U9548 ( .A(n10495), .B(n10494), .S0(n5514), .Y(n10496) );
  MXI2X2 U9549 ( .A(n10780), .B(n10779), .S0(n5519), .Y(n10781) );
  MXI2X2 U9550 ( .A(n10213), .B(n10212), .S0(n5513), .Y(n10214) );
  MXI2X2 U9551 ( .A(n10658), .B(n10657), .S0(n5516), .Y(n10659) );
  AOI222XL U9552 ( .A0(n5498), .A1(n11430), .B0(mem_rdata_D[80]), .B1(n235), 
        .C0(n12971), .C1(n4385), .Y(n10292) );
  AOI222XL U9553 ( .A0(n5499), .A1(n11428), .B0(mem_rdata_D[78]), .B1(n236), 
        .C0(n12973), .C1(n5497), .Y(n10745) );
  AOI222XL U9554 ( .A0(n5499), .A1(n11426), .B0(mem_rdata_D[76]), .B1(n233), 
        .C0(n12975), .C1(n5497), .Y(n10723) );
  AOI222XL U9555 ( .A0(n5499), .A1(n11425), .B0(mem_rdata_D[75]), .B1(n234), 
        .C0(n12976), .C1(n5497), .Y(n10711) );
  MXI2X2 U9556 ( .A(n10074), .B(n10073), .S0(n5513), .Y(n10075) );
  AOI222XL U9557 ( .A0(n5496), .A1(n11477), .B0(mem_rdata_D[127]), .B1(n234), 
        .C0(n12956), .C1(n5493), .Y(n10869) );
  MXI2X2 U9558 ( .A(n10140), .B(n10139), .S0(n5513), .Y(n10141) );
  AOI222XL U9559 ( .A0(n5495), .A1(n11474), .B0(mem_rdata_D[124]), .B1(n236), 
        .C0(n12959), .C1(n5494), .Y(n10476) );
  AOI222XL U9560 ( .A0(n5496), .A1(n11467), .B0(mem_rdata_D[117]), .B1(n233), 
        .C0(n12966), .C1(n5493), .Y(n10668) );
  MXI2X2 U9561 ( .A(n10720), .B(n10719), .S0(n5518), .Y(n10721) );
  AOI222XL U9562 ( .A0(n5511), .A1(n11413), .B0(mem_rdata_D[63]), .B1(n235), 
        .C0(n12956), .C1(n5507), .Y(n10878) );
  AOI222XL U9563 ( .A0(n5511), .A1(n11411), .B0(mem_rdata_D[61]), .B1(n235), 
        .C0(n12958), .C1(n5507), .Y(n10691) );
  MXI2X2 U9564 ( .A(n10485), .B(n10484), .S0(n5514), .Y(n10486) );
  MXI2X2 U9565 ( .A(n10311), .B(n10310), .S0(n5514), .Y(n10312) );
  MXI2X2 U9566 ( .A(n10279), .B(n10278), .S0(n5514), .Y(n10280) );
  AOI222XL U9567 ( .A0(n5511), .A1(n11399), .B0(mem_rdata_D[49]), .B1(n236), 
        .C0(n12970), .C1(n5507), .Y(n10773) );
  MXI2X2 U9568 ( .A(n10298), .B(n10297), .S0(n5514), .Y(n10299) );
  AOI222XL U9569 ( .A0(n5511), .A1(n11397), .B0(mem_rdata_D[47]), .B1(n232), 
        .C0(n12972), .C1(n5507), .Y(n10762) );
  AOI222XL U9570 ( .A0(n5511), .A1(n11396), .B0(mem_rdata_D[46]), .B1(n236), 
        .C0(n12973), .C1(n5507), .Y(n10751) );
  MXI2X2 U9571 ( .A(n10705), .B(n10704), .S0(n5517), .Y(n10706) );
  MXI2X2 U9572 ( .A(n10944), .B(n10943), .S0(n5522), .Y(n10945) );
  MXI2X2 U9573 ( .A(n10982), .B(n10981), .S0(n5523), .Y(n10983) );
  MXI2X2 U9574 ( .A(n10970), .B(n10969), .S0(n5522), .Y(n10971) );
  AOI222XL U9575 ( .A0(n5500), .A1(n11414), .B0(mem_rdata_D[64]), .B1(n233), 
        .C0(n12987), .C1(n4385), .Y(n10957) );
  MXI2X2 U9576 ( .A(n10941), .B(n10940), .S0(n5522), .Y(n10942) );
  AOI222XL U9577 ( .A0(n5495), .A1(n11454), .B0(mem_rdata_D[104]), .B1(n233), 
        .C0(n12979), .C1(n5494), .Y(n10894) );
  MXI2X2 U9578 ( .A(n10979), .B(n10978), .S0(n5523), .Y(n10980) );
  MXI2X2 U9579 ( .A(n10967), .B(n10966), .S0(n5522), .Y(n10968) );
  AOI222XL U9580 ( .A0(n5495), .A1(n11446), .B0(mem_rdata_D[96]), .B1(n236), 
        .C0(n12987), .C1(n5494), .Y(n10954) );
  AOI222XL U9581 ( .A0(n5512), .A1(n11405), .B0(mem_rdata_D[55]), .B1(n235), 
        .C0(n12964), .C1(n4421), .Y(n10950) );
  MXI2X2 U9582 ( .A(n10976), .B(n10975), .S0(n5522), .Y(n10977) );
  MXI2X2 U9583 ( .A(n10924), .B(n10923), .S0(n5521), .Y(n10925) );
  MXI2X2 U9584 ( .A(n10938), .B(n10937), .S0(n5521), .Y(n10939) );
  MXI2X2 U9585 ( .A(n10992), .B(n10991), .S0(n5523), .Y(n10993) );
  MXI2X2 U9586 ( .A(n11000), .B(n10999), .S0(n5523), .Y(n11001) );
  XOR2X1 U9587 ( .A(n10176), .B(ICACHE_addr[1]), .Y(n11078) );
  AOI21X2 U9588 ( .A0(n9976), .A1(n9983), .B0(n9975), .Y(n10927) );
  NOR2XL U9589 ( .A(n11349), .B(n11346), .Y(n9975) );
  OAI21XL U9590 ( .A0(n3854), .A1(n11479), .B0(n11349), .Y(n9976) );
  XOR2X1 U9591 ( .A(n10173), .B(ICACHE_addr[5]), .Y(n10804) );
  XOR2X1 U9592 ( .A(n10232), .B(ICACHE_addr[9]), .Y(n10595) );
  XOR2X1 U9593 ( .A(n10235), .B(ICACHE_addr[11]), .Y(n10604) );
  XOR2X1 U9594 ( .A(n10241), .B(ICACHE_addr[13]), .Y(n10425) );
  NAND2XL U9595 ( .A(n10138), .B(n4661), .Y(n10066) );
  NAND2XL U9596 ( .A(n10174), .B(ICACHE_addr[5]), .Y(n10175) );
  XOR2X1 U9597 ( .A(n10243), .B(ICACHE_addr[12]), .Y(n10410) );
  NAND2X1 U9598 ( .A(n10242), .B(ICACHE_addr[11]), .Y(n10243) );
  OA22XL U9599 ( .A0(\i_MIPS/ALUin1[7] ), .A1(n4670), .B0(\i_MIPS/ALUin1[6] ), 
        .B1(n3828), .Y(net105043) );
  OA22XL U9600 ( .A0(\i_MIPS/ALUin1[5] ), .A1(n4669), .B0(\i_MIPS/ALUin1[4] ), 
        .B1(n3828), .Y(n6851) );
  OA22XL U9601 ( .A0(\i_MIPS/ALUin1[24] ), .A1(n4670), .B0(\i_MIPS/ALUin1[25] ), .B1(n3828), .Y(n8164) );
  NAND2X1 U9602 ( .A(\i_MIPS/ALUin1[25] ), .B(n6586), .Y(n9040) );
  OAI222XL U9603 ( .A0(n5468), .A1(n1938), .B0(n5409), .B1(n5465), .C0(n5559), 
        .C1(\i_MIPS/n210 ), .Y(n11518) );
  OAI222XL U9604 ( .A0(n5467), .A1(n1937), .B0(n1998), .B1(n5464), .C0(n5558), 
        .C1(\i_MIPS/n214 ), .Y(n11514) );
  OAI222XL U9605 ( .A0(n5467), .A1(n265), .B0(n4439), .B1(n5464), .C0(n5558), 
        .C1(\i_MIPS/n213 ), .Y(n11515) );
  OAI222XL U9606 ( .A0(n5467), .A1(n284), .B0(n1993), .B1(n5464), .C0(n5558), 
        .C1(\i_MIPS/n212 ), .Y(n11516) );
  OAI222XL U9607 ( .A0(n10865), .A1(n278), .B0(n1995), .B1(n5465), .C0(n5559), 
        .C1(\i_MIPS/n211 ), .Y(n11517) );
  AO22X2 U9608 ( .A0(n5528), .A1(n12931), .B0(n5526), .B1(n11504), .Y(n11023)
         );
  AO22X2 U9609 ( .A0(n5528), .A1(n12933), .B0(n5526), .B1(n11502), .Y(n11022)
         );
  AO22X2 U9610 ( .A0(n5528), .A1(n12942), .B0(n5527), .B1(n11493), .Y(n11032)
         );
  AO22X2 U9611 ( .A0(n5528), .A1(n12946), .B0(n5527), .B1(n11489), .Y(n11030)
         );
  AO22X2 U9612 ( .A0(n5528), .A1(n12947), .B0(n5527), .B1(n11488), .Y(n11031)
         );
  AO22X2 U9613 ( .A0(n5544), .A1(ICACHE_addr[5]), .B0(n239), .B1(n11320), .Y(
        n11151) );
  AO22X2 U9614 ( .A0(mem_rdata_I[23]), .A1(n5538), .B0(n252), .B1(n11209), .Y(
        n9837) );
  AO22X2 U9615 ( .A0(mem_rdata_I[22]), .A1(n5538), .B0(n250), .B1(n11208), .Y(
        n9873) );
  AO22X2 U9616 ( .A0(mem_rdata_I[21]), .A1(n5538), .B0(n250), .B1(n11207), .Y(
        n9857) );
  AO22X2 U9617 ( .A0(mem_rdata_I[19]), .A1(n5535), .B0(n249), .B1(n11205), .Y(
        n11118) );
  AO22X2 U9618 ( .A0(mem_rdata_I[55]), .A1(n5538), .B0(n251), .B1(n11241), .Y(
        n9841) );
  AO22X2 U9619 ( .A0(mem_rdata_I[53]), .A1(n5538), .B0(n249), .B1(n11239), .Y(
        n9861) );
  AO22X2 U9620 ( .A0(mem_rdata_I[92]), .A1(n5543), .B0(n250), .B1(n11278), .Y(
        n6166) );
  AO22X2 U9621 ( .A0(mem_rdata_I[87]), .A1(n5538), .B0(n250), .B1(n11273), .Y(
        n9833) );
  AO22X2 U9622 ( .A0(mem_rdata_I[86]), .A1(n5538), .B0(n250), .B1(n11272), .Y(
        n9869) );
  AO22X2 U9623 ( .A0(mem_rdata_I[85]), .A1(n5538), .B0(n249), .B1(n11271), .Y(
        n9853) );
  AO22X2 U9624 ( .A0(mem_rdata_I[83]), .A1(n5535), .B0(n250), .B1(n11269), .Y(
        n11117) );
  AO22X2 U9625 ( .A0(mem_rdata_I[124]), .A1(n5543), .B0(n251), .B1(n11310), 
        .Y(n6161) );
  AO22X2 U9626 ( .A0(mem_rdata_I[115]), .A1(n5535), .B0(n252), .B1(n11301), 
        .Y(n11116) );
  AO22X2 U9627 ( .A0(mem_rdata_I[113]), .A1(n5544), .B0(n249), .B1(n11299), 
        .Y(n10157) );
  AO22X2 U9628 ( .A0(mem_rdata_I[108]), .A1(n5539), .B0(n249), .B1(n11294), 
        .Y(n9764) );
  AO22X2 U9629 ( .A0(mem_rdata_I[101]), .A1(n5538), .B0(n250), .B1(n11287), 
        .Y(n9914) );
  AO22X2 U9630 ( .A0(n5544), .A1(ICACHE_addr[17]), .B0(n239), .B1(n11332), .Y(
        n11156) );
  OAI221XL U9631 ( .A0(\i_MIPS/Register/register[2][24] ), .A1(net112076), 
        .B0(\i_MIPS/Register/register[10][24] ), .B1(net112096), .C0(n8280), 
        .Y(n8283) );
  OAI221XL U9632 ( .A0(\i_MIPS/Register/register[2][21] ), .A1(net112078), 
        .B0(\i_MIPS/Register/register[10][21] ), .B1(net112098), .C0(n9121), 
        .Y(n9124) );
  OAI221XL U9633 ( .A0(\i_MIPS/Register/register[2][28] ), .A1(net112078), 
        .B0(\i_MIPS/Register/register[10][28] ), .B1(net112096), .C0(n8469), 
        .Y(n8472) );
  OAI221XL U9634 ( .A0(\i_MIPS/Register/register[2][20] ), .A1(net112078), 
        .B0(\i_MIPS/Register/register[10][20] ), .B1(net112098), .C0(n9226), 
        .Y(n9229) );
  OA22X1 U9635 ( .A0(\i_MIPS/Register/register[6][20] ), .A1(net112116), .B0(
        \i_MIPS/Register/register[14][20] ), .B1(net112142), .Y(n9226) );
  OAI221XL U9636 ( .A0(\i_MIPS/Register/register[2][14] ), .A1(net112072), 
        .B0(\i_MIPS/Register/register[10][14] ), .B1(net112090), .C0(n7629), 
        .Y(n7632) );
  OAI221XL U9637 ( .A0(\i_MIPS/Register/register[2][16] ), .A1(net112076), 
        .B0(\i_MIPS/Register/register[10][16] ), .B1(net112090), .C0(n8051), 
        .Y(n8054) );
  OAI221XL U9638 ( .A0(\i_MIPS/Register/register[2][6] ), .A1(net112072), .B0(
        \i_MIPS/Register/register[10][6] ), .B1(net112090), .C0(n6988), .Y(
        n6991) );
  OA22X1 U9639 ( .A0(\i_MIPS/Register/register[6][6] ), .A1(net112110), .B0(
        \i_MIPS/Register/register[14][6] ), .B1(net112128), .Y(n6988) );
  OAI221XL U9640 ( .A0(\i_MIPS/Register/register[2][4] ), .A1(net112072), .B0(
        \i_MIPS/Register/register[10][4] ), .B1(net112090), .C0(n6863), .Y(
        n6866) );
  OAI221XL U9641 ( .A0(\i_MIPS/Register/register[2][7] ), .A1(net112076), .B0(
        \i_MIPS/Register/register[10][7] ), .B1(net112090), .C0(n7914), .Y(
        n7917) );
  OAI221XL U9642 ( .A0(\i_MIPS/Register/register[2][0] ), .A1(net112072), .B0(
        \i_MIPS/Register/register[10][0] ), .B1(net112098), .C0(n7556), .Y(
        n7559) );
  OAI221XL U9643 ( .A0(\i_MIPS/Register/register[2][23] ), .A1(net112078), 
        .B0(\i_MIPS/Register/register[10][23] ), .B1(net112098), .C0(n8832), 
        .Y(n8835) );
  OAI221XL U9644 ( .A0(\i_MIPS/Register/register[2][18] ), .A1(net112078), 
        .B0(\i_MIPS/Register/register[10][18] ), .B1(net112098), .C0(n8769), 
        .Y(n8772) );
  OA22X1 U9645 ( .A0(\i_MIPS/Register/register[6][18] ), .A1(net112116), .B0(
        \i_MIPS/Register/register[14][18] ), .B1(net112134), .Y(n8769) );
  OAI221XL U9646 ( .A0(\i_MIPS/Register/register[2][5] ), .A1(net112072), .B0(
        \i_MIPS/Register/register[10][5] ), .B1(net112090), .C0(n6782), .Y(
        n6785) );
  OAI221XL U9647 ( .A0(\i_MIPS/Register/register[2][11] ), .A1(net112072), 
        .B0(\i_MIPS/Register/register[10][11] ), .B1(net112098), .C0(n7248), 
        .Y(n7251) );
  OAI221XL U9648 ( .A0(\i_MIPS/Register/register[2][25] ), .A1(net112078), 
        .B0(\i_MIPS/Register/register[10][25] ), .B1(net112098), .C0(n9024), 
        .Y(n9027) );
  OAI221XL U9649 ( .A0(\i_MIPS/Register/register[2][26] ), .A1(net112078), 
        .B0(\i_MIPS/Register/register[10][26] ), .B1(net112098), .C0(n8923), 
        .Y(n8926) );
  OAI221XL U9650 ( .A0(\i_MIPS/Register/register[2][29] ), .A1(net112076), 
        .B0(\i_MIPS/Register/register[10][29] ), .B1(net112096), .C0(n8134), 
        .Y(n8137) );
  OAI221XL U9651 ( .A0(\i_MIPS/Register/register[2][22] ), .A1(net112078), 
        .B0(\i_MIPS/Register/register[10][22] ), .B1(net112100), .C0(n9437), 
        .Y(n9440) );
  OAI221XL U9652 ( .A0(\i_MIPS/Register/register[2][31] ), .A1(net112072), 
        .B0(\i_MIPS/Register/register[10][31] ), .B1(net112090), .C0(n6663), 
        .Y(n6666) );
  OAI221XL U9653 ( .A0(\i_MIPS/Register/register[2][27] ), .A1(n4690), .B0(
        \i_MIPS/Register/register[10][27] ), .B1(n4686), .C0(n9405), .Y(n9408)
         );
  OAI31XL U9654 ( .A0(n9892), .A1(\i_MIPS/IR_ID[30] ), .A2(\i_MIPS/IR_ID[27] ), 
        .B0(\i_MIPS/Control_ID/n15 ), .Y(n9893) );
  CLKINVX1 U9655 ( .A(\i_MIPS/n251 ), .Y(n10680) );
  OA22XL U9656 ( .A0(n4626), .A1(n3804), .B0(n4649), .B1(n4625), .Y(n4624) );
  NOR4X1 U9657 ( .A(n9369), .B(n9368), .C(n9367), .D(n9366), .Y(n9380) );
  NAND4X1 U9658 ( .A(n9364), .B(n9363), .C(n9362), .D(n9361), .Y(n9369) );
  AO22X1 U9659 ( .A0(net112050), .A1(n285), .B0(net100603), .B1(n430), .Y(
        n9367) );
  NOR4X1 U9660 ( .A(n6676), .B(n6675), .C(n6674), .D(n6673), .Y(n6677) );
  OAI221XL U9661 ( .A0(\i_MIPS/Register/register[18][31] ), .A1(net112072), 
        .B0(\i_MIPS/Register/register[26][31] ), .B1(net112090), .C0(n6672), 
        .Y(n6675) );
  NAND4X1 U9662 ( .A(n6671), .B(n6670), .C(n6669), .D(n6668), .Y(n6676) );
  AO22X1 U9663 ( .A0(net112036), .A1(n434), .B0(net100603), .B1(n2014), .Y(
        n6674) );
  NOR4X1 U9664 ( .A(n9450), .B(n9449), .C(n9448), .D(n9447), .Y(n9451) );
  OAI221XL U9665 ( .A0(\i_MIPS/Register/register[18][22] ), .A1(net112078), 
        .B0(\i_MIPS/Register/register[26][22] ), .B1(net112100), .C0(n9446), 
        .Y(n9449) );
  NAND4X1 U9666 ( .A(n9445), .B(n9444), .C(n9443), .D(n9442), .Y(n9450) );
  AO22X1 U9667 ( .A0(net112050), .A1(n957), .B0(net100603), .B1(n2473), .Y(
        n9448) );
  NOR4X1 U9668 ( .A(n9378), .B(n9377), .C(n9376), .D(n9375), .Y(n9379) );
  NAND4X1 U9669 ( .A(n9373), .B(n9372), .C(n9371), .D(n9370), .Y(n9378) );
  AO22X1 U9670 ( .A0(net112050), .A1(n286), .B0(net100603), .B1(n431), .Y(
        n9376) );
  NOR4X1 U9671 ( .A(n7340), .B(n7339), .C(n7338), .D(n7337), .Y(n7341) );
  NAND4X1 U9672 ( .A(n7335), .B(n7334), .C(n7333), .D(n7332), .Y(n7340) );
  AO22X1 U9673 ( .A0(net112038), .A1(n394), .B0(net100603), .B1(n1043), .Y(
        n7338) );
  NOR4X1 U9674 ( .A(n8782), .B(n8781), .C(n8780), .D(n8779), .Y(n8783) );
  NAND4X1 U9675 ( .A(n8777), .B(n8776), .C(n8775), .D(n8774), .Y(n8782) );
  AO22X1 U9676 ( .A0(net112038), .A1(n1008), .B0(net100603), .B1(n2534), .Y(
        n8780) );
  NAND4X1 U9677 ( .A(n8001), .B(n8000), .C(n7999), .D(n7998), .Y(n8006) );
  AO22X1 U9678 ( .A0(net112036), .A1(n1009), .B0(net100603), .B1(n2535), .Y(
        n8004) );
  NAND4X1 U9679 ( .A(n7730), .B(n7729), .C(n7728), .D(n7727), .Y(n7735) );
  NOR4X1 U9680 ( .A(n9239), .B(n9238), .C(n9237), .D(n9236), .Y(n9240) );
  NAND4X1 U9681 ( .A(n9234), .B(n9233), .C(n9232), .D(n9231), .Y(n9239) );
  AO22X1 U9682 ( .A0(net112050), .A1(n958), .B0(net100603), .B1(n2474), .Y(
        n9237) );
  NAND4X1 U9683 ( .A(n7637), .B(n7636), .C(n7635), .D(n7634), .Y(n7642) );
  AO22X1 U9684 ( .A0(net112038), .A1(n395), .B0(net100603), .B1(n1044), .Y(
        n7640) );
  NOR4X1 U9685 ( .A(n9134), .B(n9133), .C(n9132), .D(n9131), .Y(n9135) );
  OAI221XL U9686 ( .A0(\i_MIPS/Register/register[18][21] ), .A1(net112078), 
        .B0(\i_MIPS/Register/register[26][21] ), .B1(net112098), .C0(n9130), 
        .Y(n9133) );
  NAND4X1 U9687 ( .A(n9129), .B(n9128), .C(n9127), .D(n9126), .Y(n9134) );
  AO22X1 U9688 ( .A0(net112050), .A1(n1010), .B0(net100603), .B1(n2536), .Y(
        n9132) );
  NOR4X1 U9689 ( .A(n7001), .B(n7000), .C(n6999), .D(n6998), .Y(n7002) );
  NAND4X1 U9690 ( .A(n6996), .B(n6995), .C(n6994), .D(n6993), .Y(n7001) );
  NOR4X1 U9691 ( .A(n8064), .B(n8063), .C(n8062), .D(n8061), .Y(n8065) );
  NAND4X1 U9692 ( .A(n8059), .B(n8058), .C(n8057), .D(n8056), .Y(n8064) );
  NOR4X1 U9693 ( .A(n8845), .B(n8844), .C(n8843), .D(n8842), .Y(n8846) );
  OAI221XL U9694 ( .A0(\i_MIPS/Register/register[18][23] ), .A1(net112078), 
        .B0(\i_MIPS/Register/register[26][23] ), .B1(net112098), .C0(n8841), 
        .Y(n8844) );
  NAND4X1 U9695 ( .A(n8840), .B(n8839), .C(n8838), .D(n8837), .Y(n8845) );
  AO22X1 U9696 ( .A0(net112038), .A1(n1011), .B0(net100603), .B1(n2537), .Y(
        n8843) );
  NOR4X1 U9697 ( .A(n8482), .B(n8481), .C(n8480), .D(n8479), .Y(n8483) );
  NAND4X1 U9698 ( .A(n8477), .B(n8476), .C(n8475), .D(n8474), .Y(n8482) );
  AO22X1 U9699 ( .A0(net112038), .A1(n959), .B0(net100603), .B1(n2475), .Y(
        n8480) );
  NOR4X1 U9700 ( .A(n8384), .B(n8383), .C(n8382), .D(n8381), .Y(n8385) );
  OAI221XL U9701 ( .A0(\i_MIPS/Register/register[18][3] ), .A1(net112078), 
        .B0(\i_MIPS/Register/register[26][3] ), .B1(net112096), .C0(n8380), 
        .Y(n8383) );
  NAND4X1 U9702 ( .A(n8379), .B(n8378), .C(n8377), .D(n8376), .Y(n8384) );
  AO22X1 U9703 ( .A0(net112038), .A1(n1012), .B0(net100603), .B1(n2538), .Y(
        n8382) );
  NOR4X1 U9704 ( .A(n8680), .B(n8679), .C(n8678), .D(n8677), .Y(n8681) );
  OAI221XL U9705 ( .A0(\i_MIPS/Register/register[18][9] ), .A1(net112078), 
        .B0(\i_MIPS/Register/register[26][9] ), .B1(net112096), .C0(n8676), 
        .Y(n8679) );
  NAND4X1 U9706 ( .A(n8675), .B(n8674), .C(n8673), .D(n8672), .Y(n8680) );
  AO22X1 U9707 ( .A0(net112038), .A1(n1013), .B0(net100603), .B1(n2539), .Y(
        n8678) );
  OAI221XL U9708 ( .A0(\i_MIPS/Register/register[18][7] ), .A1(net112076), 
        .B0(\i_MIPS/Register/register[26][7] ), .B1(net112090), .C0(n7923), 
        .Y(n7926) );
  NAND4X1 U9709 ( .A(n7564), .B(n7563), .C(n7562), .D(n7561), .Y(n7569) );
  AO22X1 U9710 ( .A0(net112038), .A1(n396), .B0(net100603), .B1(n1045), .Y(
        n7567) );
  NOR4X1 U9711 ( .A(n9037), .B(n9036), .C(n9035), .D(n9034), .Y(n9038) );
  OAI221XL U9712 ( .A0(\i_MIPS/Register/register[18][25] ), .A1(net112078), 
        .B0(\i_MIPS/Register/register[26][25] ), .B1(net112098), .C0(n9033), 
        .Y(n9036) );
  NAND4X1 U9713 ( .A(n9032), .B(n9031), .C(n9030), .D(n9029), .Y(n9037) );
  AO22X1 U9714 ( .A0(net112050), .A1(n1014), .B0(net100603), .B1(n2540), .Y(
        n9035) );
  NOR4X1 U9715 ( .A(n6876), .B(n6875), .C(n6874), .D(n6873), .Y(n6877) );
  OAI221XL U9716 ( .A0(\i_MIPS/Register/register[18][4] ), .A1(net112072), 
        .B0(\i_MIPS/Register/register[26][4] ), .B1(net112090), .C0(n6872), 
        .Y(n6875) );
  NAND4X1 U9717 ( .A(n6871), .B(n6870), .C(n6869), .D(n6868), .Y(n6876) );
  AO22X1 U9718 ( .A0(net112036), .A1(n1015), .B0(net100603), .B1(n2541), .Y(
        n6874) );
  NOR4X1 U9719 ( .A(n8936), .B(n8935), .C(n8934), .D(n8933), .Y(n8937) );
  OAI221XL U9720 ( .A0(\i_MIPS/Register/register[18][26] ), .A1(net112078), 
        .B0(\i_MIPS/Register/register[26][26] ), .B1(net112098), .C0(n8932), 
        .Y(n8935) );
  NAND4X1 U9721 ( .A(n8931), .B(n8930), .C(n8929), .D(n8928), .Y(n8936) );
  AO22X1 U9722 ( .A0(net112050), .A1(n960), .B0(net100603), .B1(n2476), .Y(
        n8934) );
  NOR4X1 U9723 ( .A(n8293), .B(n8292), .C(n8291), .D(n8290), .Y(n8294) );
  OAI221XL U9724 ( .A0(\i_MIPS/Register/register[18][24] ), .A1(net112078), 
        .B0(\i_MIPS/Register/register[26][24] ), .B1(net112096), .C0(n8289), 
        .Y(n8292) );
  NAND4X1 U9725 ( .A(n8288), .B(n8287), .C(n8286), .D(n8285), .Y(n8293) );
  AO22X1 U9726 ( .A0(net112038), .A1(n1016), .B0(net100603), .B1(n2542), .Y(
        n8291) );
  NOR4X1 U9727 ( .A(n7144), .B(n7143), .C(n7142), .D(n7141), .Y(n7145) );
  NAND4X1 U9728 ( .A(n7139), .B(n7138), .C(n7137), .D(n7136), .Y(n7144) );
  AO22X1 U9729 ( .A0(net112038), .A1(n397), .B0(net100603), .B1(n1046), .Y(
        n7142) );
  NOR4X1 U9730 ( .A(n7085), .B(n7084), .C(n7083), .D(n7082), .Y(n7086) );
  NAND4X1 U9731 ( .A(n7080), .B(n7079), .C(n7078), .D(n7077), .Y(n7085) );
  AO22X1 U9732 ( .A0(net112036), .A1(n961), .B0(net100603), .B1(n2477), .Y(
        n7083) );
  NOR4X1 U9733 ( .A(n7261), .B(n7260), .C(n7259), .D(n7258), .Y(n7262) );
  OAI221XL U9734 ( .A0(\i_MIPS/Register/register[18][11] ), .A1(net112072), 
        .B0(\i_MIPS/Register/register[26][11] ), .B1(net112098), .C0(n7257), 
        .Y(n7260) );
  NAND4X1 U9735 ( .A(n7256), .B(n7255), .C(n7254), .D(n7253), .Y(n7261) );
  AO22X1 U9736 ( .A0(net112038), .A1(n398), .B0(net100603), .B1(n1047), .Y(
        n7259) );
  NOR4X1 U9737 ( .A(n6795), .B(n6794), .C(n6793), .D(n6792), .Y(n6796) );
  OAI221XL U9738 ( .A0(\i_MIPS/Register/register[18][5] ), .A1(net112072), 
        .B0(\i_MIPS/Register/register[26][5] ), .B1(net112090), .C0(n6791), 
        .Y(n6794) );
  NAND4X1 U9739 ( .A(n6790), .B(n6789), .C(n6788), .D(n6787), .Y(n6795) );
  AO22X1 U9740 ( .A0(net112036), .A1(n1017), .B0(net100603), .B1(n2543), .Y(
        n6793) );
  NOR4X1 U9741 ( .A(n7397), .B(n7396), .C(n7395), .D(n7394), .Y(n7398) );
  NAND4X1 U9742 ( .A(n7392), .B(n7391), .C(n7390), .D(n7389), .Y(n7397) );
  AO22X1 U9743 ( .A0(net112038), .A1(n399), .B0(net100603), .B1(n1048), .Y(
        n7395) );
  NOR4X1 U9744 ( .A(n8147), .B(n8146), .C(n8145), .D(n8144), .Y(n8148) );
  OAI221XL U9745 ( .A0(\i_MIPS/Register/register[18][29] ), .A1(net112076), 
        .B0(\i_MIPS/Register/register[26][29] ), .B1(net112096), .C0(n8143), 
        .Y(n8146) );
  NAND4X1 U9746 ( .A(n8142), .B(n8141), .C(n8140), .D(n8139), .Y(n8147) );
  NOR4X1 U9747 ( .A(n7794), .B(n7793), .C(n7792), .D(n7791), .Y(n7795) );
  NAND4X1 U9748 ( .A(n7789), .B(n7788), .C(n7787), .D(n7786), .Y(n7794) );
  AO22X1 U9749 ( .A0(net112036), .A1(n1018), .B0(net100603), .B1(n2544), .Y(
        n7792) );
  MXI2X1 U9750 ( .A(\i_MIPS/ID_EX[70] ), .B(\i_MIPS/ID_EX[102] ), .S0(n5622), 
        .Y(n6594) );
  OA22X1 U9751 ( .A0(\i_MIPS/Register/register[6][23] ), .A1(n4683), .B0(
        \i_MIPS/Register/register[14][23] ), .B1(n4678), .Y(n8896) );
  OAI221XL U9752 ( .A0(\i_MIPS/Register/register[2][30] ), .A1(n4690), .B0(
        \i_MIPS/Register/register[10][30] ), .B1(n4686), .C0(n6613), .Y(n6621)
         );
  OAI221XL U9753 ( .A0(\i_MIPS/Register/register[2][4] ), .A1(n4692), .B0(
        \i_MIPS/Register/register[10][4] ), .B1(n4688), .C0(n6898), .Y(n6906)
         );
  OA22X1 U9754 ( .A0(\i_MIPS/Register/register[6][4] ), .A1(n4684), .B0(
        \i_MIPS/Register/register[14][4] ), .B1(n4680), .Y(n6898) );
  OAI221XL U9755 ( .A0(\i_MIPS/Register/register[18][7] ), .A1(n4692), .B0(
        \i_MIPS/Register/register[26][7] ), .B1(n4687), .C0(n7958), .Y(n7966)
         );
  OAI221XL U9756 ( .A0(\i_MIPS/Register/register[2][7] ), .A1(n4692), .B0(
        \i_MIPS/Register/register[10][7] ), .B1(n4687), .C0(n7949), .Y(n7957)
         );
  OAI221XL U9757 ( .A0(\i_MIPS/Register/register[2][17] ), .A1(n4692), .B0(
        \i_MIPS/Register/register[10][17] ), .B1(n4687), .C0(n7855), .Y(n7863)
         );
  OAI221XL U9758 ( .A0(\i_MIPS/Register/register[18][0] ), .A1(n4692), .B0(
        \i_MIPS/Register/register[26][0] ), .B1(n4687), .C0(n7600), .Y(n7608)
         );
  OAI221XL U9759 ( .A0(\i_MIPS/Register/register[18][11] ), .A1(n4691), .B0(
        \i_MIPS/Register/register[26][11] ), .B1(n4688), .C0(n7291), .Y(n7299)
         );
  OAI221XL U9760 ( .A0(\i_MIPS/Register/register[2][11] ), .A1(n4690), .B0(
        \i_MIPS/Register/register[10][11] ), .B1(n4688), .C0(n7282), .Y(n7290)
         );
  OAI221XL U9761 ( .A0(\i_MIPS/Register/register[18][10] ), .A1(n4692), .B0(
        \i_MIPS/Register/register[26][10] ), .B1(n4688), .C0(n7371), .Y(n7379)
         );
  OAI221XL U9762 ( .A0(\i_MIPS/Register/register[2][10] ), .A1(n4691), .B0(
        \i_MIPS/Register/register[10][10] ), .B1(n4688), .C0(n7362), .Y(n7370)
         );
  OAI221XL U9763 ( .A0(\i_MIPS/Register/register[18][15] ), .A1(n4690), .B0(
        \i_MIPS/Register/register[26][15] ), .B1(n4688), .C0(n7209), .Y(n7217)
         );
  OAI221XL U9764 ( .A0(\i_MIPS/Register/register[2][15] ), .A1(n4690), .B0(
        \i_MIPS/Register/register[10][15] ), .B1(n4688), .C0(n7200), .Y(n7208)
         );
  OAI221XL U9765 ( .A0(\i_MIPS/Register/register[18][9] ), .A1(n4691), .B0(
        \i_MIPS/Register/register[26][9] ), .B1(n4688), .C0(n8711), .Y(n8719)
         );
  OA22X1 U9766 ( .A0(\i_MIPS/Register/register[22][9] ), .A1(n4682), .B0(
        \i_MIPS/Register/register[30][9] ), .B1(n4679), .Y(n8711) );
  OAI221XL U9767 ( .A0(\i_MIPS/Register/register[2][9] ), .A1(n4691), .B0(
        \i_MIPS/Register/register[10][9] ), .B1(n4687), .C0(n8702), .Y(n8710)
         );
  OA22X1 U9768 ( .A0(\i_MIPS/Register/register[6][9] ), .A1(n4682), .B0(
        \i_MIPS/Register/register[14][9] ), .B1(n4679), .Y(n8702) );
  OAI221XL U9769 ( .A0(\i_MIPS/Register/register[18][18] ), .A1(n4691), .B0(
        \i_MIPS/Register/register[26][18] ), .B1(n4688), .C0(n8813), .Y(n8821)
         );
  OA22X1 U9770 ( .A0(\i_MIPS/Register/register[22][18] ), .A1(n4684), .B0(
        \i_MIPS/Register/register[30][18] ), .B1(n4678), .Y(n8813) );
  OAI221XL U9771 ( .A0(\i_MIPS/Register/register[2][18] ), .A1(n4691), .B0(
        \i_MIPS/Register/register[10][18] ), .B1(n4686), .C0(n8804), .Y(n8812)
         );
  OA22X1 U9772 ( .A0(\i_MIPS/Register/register[6][18] ), .A1(n4683), .B0(
        \i_MIPS/Register/register[14][18] ), .B1(n4678), .Y(n8804) );
  OAI221XL U9773 ( .A0(\i_MIPS/Register/register[2][19] ), .A1(n4691), .B0(
        \i_MIPS/Register/register[10][19] ), .B1(n4687), .C0(n8607), .Y(n8615)
         );
  OA22X1 U9774 ( .A0(\i_MIPS/Register/register[6][19] ), .A1(n4682), .B0(
        \i_MIPS/Register/register[14][19] ), .B1(n4679), .Y(n8607) );
  OAI221XL U9775 ( .A0(\i_MIPS/Register/register[2][19] ), .A1(net112078), 
        .B0(\i_MIPS/Register/register[10][19] ), .B1(net112096), .C0(n8567), 
        .Y(n8575) );
  OAI221XL U9776 ( .A0(\i_MIPS/Register/register[18][25] ), .A1(n4690), .B0(
        \i_MIPS/Register/register[26][25] ), .B1(n4686), .C0(n9103), .Y(n9111)
         );
  OAI221XL U9777 ( .A0(\i_MIPS/Register/register[2][25] ), .A1(n4690), .B0(
        \i_MIPS/Register/register[10][25] ), .B1(n4686), .C0(n9094), .Y(n9102)
         );
  OAI221XL U9778 ( .A0(\i_MIPS/Register/register[18][30] ), .A1(net112072), 
        .B0(\i_MIPS/Register/register[26][30] ), .B1(net112090), .C0(n6468), 
        .Y(n6476) );
  OAI221XL U9779 ( .A0(\i_MIPS/Register/register[2][30] ), .A1(net112072), 
        .B0(\i_MIPS/Register/register[10][30] ), .B1(net112090), .C0(n6459), 
        .Y(n6467) );
  AND3XL U9780 ( .A(net108200), .B(\i_MIPS/n326 ), .C(\i_MIPS/n330 ), .Y(n9570) );
  XNOR2XL U9781 ( .A(\i_MIPS/IR_ID[16] ), .B(\i_MIPS/Reg_W[0] ), .Y(n6634) );
  XNOR2XL U9782 ( .A(\i_MIPS/IR_ID[17] ), .B(\i_MIPS/Reg_W[1] ), .Y(n6635) );
  XNOR2XL U9783 ( .A(\i_MIPS/IR_ID[18] ), .B(\i_MIPS/Reg_W[2] ), .Y(n6636) );
  XOR2X1 U9784 ( .A(\i_MIPS/PHT_2/counter ), .B(n11042), .Y(\i_MIPS/PHT_2/n54 ) );
  OAI22XL U9785 ( .A0(\i_MIPS/Register/register[9][31] ), .A1(n9410), .B0(
        \i_MIPS/Register/register[1][31] ), .B1(n9411), .Y(n6718) );
  NOR2X1 U9786 ( .A(n6734), .B(n6733), .Y(n6742) );
  OAI22XL U9787 ( .A0(\i_MIPS/Register/register[31][31] ), .A1(n9416), .B0(
        \i_MIPS/Register/register[23][31] ), .B1(n9417), .Y(n6734) );
  OAI22XL U9788 ( .A0(\i_MIPS/Register/register[27][31] ), .A1(n9414), .B0(
        \i_MIPS/Register/register[19][31] ), .B1(n9415), .Y(n6733) );
  NOR2X1 U9789 ( .A(n6732), .B(n6731), .Y(n6743) );
  OAI22XL U9790 ( .A0(\i_MIPS/Register/register[29][31] ), .A1(n9412), .B0(
        \i_MIPS/Register/register[21][31] ), .B1(n187), .Y(n6732) );
  OAI22XL U9791 ( .A0(\i_MIPS/Register/register[25][31] ), .A1(n9410), .B0(
        \i_MIPS/Register/register[17][31] ), .B1(n9411), .Y(n6731) );
  NOR2X1 U9792 ( .A(n6721), .B(n6720), .Y(n6729) );
  OAI22XL U9793 ( .A0(\i_MIPS/Register/register[15][31] ), .A1(n9416), .B0(
        \i_MIPS/Register/register[7][31] ), .B1(n9417), .Y(n6721) );
  OAI22XL U9794 ( .A0(\i_MIPS/Register/register[11][31] ), .A1(n9414), .B0(
        \i_MIPS/Register/register[3][31] ), .B1(n9415), .Y(n6720) );
  OAI22XL U9795 ( .A0(\i_MIPS/Register/register[13][31] ), .A1(n9412), .B0(
        \i_MIPS/Register/register[5][31] ), .B1(n189), .Y(n6719) );
  XNOR2XL U9796 ( .A(\i_MIPS/Reg_W[2] ), .B(\i_MIPS/IR_ID[23] ), .Y(n6440) );
  XNOR2XL U9797 ( .A(\i_MIPS/Reg_W[3] ), .B(\i_MIPS/IR_ID[24] ), .Y(n6442) );
  NAND3BX1 U9798 ( .AN(n4472), .B(n8153), .C(n7151), .Y(n7230) );
  XOR2X1 U9799 ( .A(n11335), .B(ICACHE_addr[20]), .Y(n5991) );
  XNOR2XL U9800 ( .A(\i_MIPS/Reg_W[3] ), .B(\i_MIPS/IR_ID[19] ), .Y(n6637) );
  OAI22XL U9801 ( .A0(n4681), .A1(\i_MIPS/Register/register[22][31] ), .B0(
        n4678), .B1(\i_MIPS/Register/register[30][31] ), .Y(n6738) );
  OAI22XL U9802 ( .A0(\i_MIPS/Register/register[18][31] ), .A1(n4690), .B0(
        \i_MIPS/Register/register[26][31] ), .B1(n4686), .Y(n6737) );
  OAI22XL U9803 ( .A0(n4697), .A1(\i_MIPS/Register/register[20][31] ), .B0(
        n4693), .B1(\i_MIPS/Register/register[28][31] ), .Y(n6739) );
  OAI22XL U9804 ( .A0(n4681), .A1(\i_MIPS/Register/register[6][31] ), .B0(
        n4678), .B1(\i_MIPS/Register/register[14][31] ), .Y(n6725) );
  OAI22XL U9805 ( .A0(\i_MIPS/Register/register[2][31] ), .A1(n4690), .B0(
        \i_MIPS/Register/register[10][31] ), .B1(n4686), .Y(n6724) );
  OAI22XL U9806 ( .A0(n4697), .A1(\i_MIPS/Register/register[4][31] ), .B0(
        n4693), .B1(\i_MIPS/Register/register[12][31] ), .Y(n6726) );
  OAI2BB2XL U9807 ( .B0(\i_MIPS/n224 ), .B1(net108198), .A0N(n5545), .A1N(
        n10591), .Y(\i_MIPS/N67 ) );
  OAI2BB2XL U9808 ( .B0(\i_MIPS/n223 ), .B1(net108198), .A0N(n4073), .A1N(
        n10812), .Y(\i_MIPS/N66 ) );
  OAI2BB2XL U9809 ( .B0(\i_MIPS/n185 ), .B1(net108198), .A0N(n4072), .A1N(
        n10176), .Y(\i_MIPS/N28 ) );
  OAI2BB2XL U9810 ( .B0(\i_MIPS/n245 ), .B1(net108198), .A0N(n5545), .A1N(
        n10371), .Y(\i_MIPS/N99 ) );
  OAI2BB2XL U9811 ( .B0(\i_MIPS/n165 ), .B1(net108194), .A0N(n4072), .A1N(
        n10409), .Y(\i_MIPS/N105 ) );
  OAI2BB2XL U9812 ( .B0(\i_MIPS/n166 ), .B1(net108194), .A0N(n4073), .A1N(
        n10424), .Y(\i_MIPS/N106 ) );
  CLKINVX1 U9813 ( .A(n10440), .Y(n10438) );
  OAI2BB2XL U9814 ( .B0(\i_MIPS/n174 ), .B1(net108194), .A0N(n4073), .A1N(
        net98501), .Y(\i_MIPS/N114 ) );
  OAI2BB2XL U9815 ( .B0(\i_MIPS/n228 ), .B1(net108200), .A0N(n4072), .A1N(
        n10422), .Y(\i_MIPS/N71 ) );
  OAI2BB2XL U9816 ( .B0(\i_MIPS/n227 ), .B1(net108200), .A0N(n4073), .A1N(
        n10406), .Y(\i_MIPS/N70 ) );
  OAI2BB2XL U9817 ( .B0(\i_MIPS/n226 ), .B1(net108200), .A0N(n4315), .A1N(
        n10601), .Y(\i_MIPS/N69 ) );
  OAI2BB2XL U9818 ( .B0(\i_MIPS/n240 ), .B1(net108190), .A0N(n5545), .A1N(
        n11079), .Y(\i_MIPS/N94 ) );
  CLKINVX1 U9819 ( .A(n11111), .Y(n11109) );
  OAI2BB2XL U9820 ( .B0(\i_MIPS/n243 ), .B1(net108190), .A0N(n4072), .A1N(
        n11095), .Y(\i_MIPS/N97 ) );
  CLKINVX1 U9821 ( .A(n11097), .Y(n11095) );
  OAI2BB2XL U9822 ( .B0(\i_MIPS/n244 ), .B1(net108192), .A0N(n4073), .A1N(
        n10803), .Y(\i_MIPS/N98 ) );
  OAI2BB2XL U9823 ( .B0(\i_MIPS/n161 ), .B1(net108190), .A0N(n4073), .A1N(
        n10815), .Y(\i_MIPS/N101 ) );
  OAI2BB2XL U9824 ( .B0(\i_MIPS/n170 ), .B1(net108192), .A0N(n4072), .A1N(
        n10635), .Y(\i_MIPS/N110 ) );
  OAI2BB2XL U9825 ( .B0(\i_MIPS/n220 ), .B1(net108198), .A0N(n4072), .A1N(
        n10800), .Y(\i_MIPS/N63 ) );
  OAI2BB2XL U9826 ( .B0(\i_MIPS/n217 ), .B1(net108198), .A0N(n5545), .A1N(
        n11106), .Y(\i_MIPS/N60 ) );
  OAI2BB2XL U9827 ( .B0(\i_MIPS/n186 ), .B1(net108198), .A0N(n4073), .A1N(
        n11077), .Y(\i_MIPS/N29 ) );
  OAI2BB2XL U9828 ( .B0(\i_MIPS/n162 ), .B1(net108192), .A0N(n4072), .A1N(
        n10594), .Y(\i_MIPS/N102 ) );
  CLKINVX1 U9829 ( .A(n10596), .Y(n10594) );
  OAI2BB2XL U9830 ( .B0(\i_MIPS/n164 ), .B1(net108192), .A0N(n5545), .A1N(n637), .Y(\i_MIPS/N104 ) );
  OAI2BB2XL U9831 ( .B0(\i_MIPS/n180 ), .B1(net108192), .A0N(n5545), .A1N(
        n4424), .Y(\i_MIPS/N120 ) );
  OAI2BB2XL U9832 ( .B0(\i_MIPS/n189 ), .B1(net108198), .A0N(n11094), .A1N(
        n4073), .Y(\i_MIPS/N32 ) );
  OAI2BB2XL U9833 ( .B0(\i_MIPS/n190 ), .B1(net108198), .A0N(n10802), .A1N(
        n4073), .Y(\i_MIPS/N33 ) );
  OAI2BB2XL U9834 ( .B0(\i_MIPS/n191 ), .B1(net108198), .A0N(n10370), .A1N(
        n5545), .Y(\i_MIPS/N34 ) );
  OAI2BB2XL U9835 ( .B0(\i_MIPS/n192 ), .B1(net108198), .A0N(n10227), .A1N(
        n4073), .Y(\i_MIPS/N35 ) );
  OAI2BB2XL U9836 ( .B0(\i_MIPS/n194 ), .B1(net108198), .A0N(n10593), .A1N(
        n4072), .Y(\i_MIPS/N37 ) );
  OAI2BB2XL U9837 ( .B0(\i_MIPS/n195 ), .B1(net108198), .A0N(n409), .A1N(n4072), .Y(\i_MIPS/N38 ) );
  OAI2BB2XL U9838 ( .B0(\i_MIPS/n197 ), .B1(net108194), .A0N(n10408), .A1N(
        n4072), .Y(\i_MIPS/N40 ) );
  OAI2BB2XL U9839 ( .B0(\i_MIPS/n198 ), .B1(net108194), .A0N(n10423), .A1N(
        n4072), .Y(\i_MIPS/N41 ) );
  OAI2BB2XL U9840 ( .B0(\i_MIPS/n199 ), .B1(net108198), .A0N(n10613), .A1N(
        n4072), .Y(\i_MIPS/N42 ) );
  OAI2BB2XL U9841 ( .B0(\i_MIPS/n209 ), .B1(net108198), .A0N(n10340), .A1N(
        n5545), .Y(\i_MIPS/N52 ) );
  OAI2BB2XL U9842 ( .B0(\i_MIPS/n210 ), .B1(net108198), .A0N(n10836), .A1N(
        n4073), .Y(\i_MIPS/N53 ) );
  OAI2BB2XL U9843 ( .B0(\i_MIPS/n212 ), .B1(net108192), .A0N(n10791), .A1N(
        n4072), .Y(\i_MIPS/N55 ) );
  OAI2BB2XL U9844 ( .B0(\i_MIPS/n206 ), .B1(net108194), .A0N(net98502), .A1N(
        n4073), .Y(\i_MIPS/N49 ) );
  OAI2BB2XL U9845 ( .B0(\i_MIPS/n207 ), .B1(net108194), .A0N(n10448), .A1N(
        n5545), .Y(\i_MIPS/N50 ) );
  OAI2BB2XL U9846 ( .B0(\i_MIPS/n208 ), .B1(net108194), .A0N(n10465), .A1N(
        n5545), .Y(\i_MIPS/N51 ) );
  OAI2BB2XL U9847 ( .B0(\i_MIPS/n211 ), .B1(net108194), .A0N(n10579), .A1N(
        n4072), .Y(\i_MIPS/N54 ) );
  OAI2BB2XL U9848 ( .B0(\i_MIPS/n239 ), .B1(net108190), .A0N(n11066), .A1N(
        n4073), .Y(\i_MIPS/N93 ) );
  CLKINVX1 U9849 ( .A(n11068), .Y(n11066) );
  OAI2BB2XL U9850 ( .B0(\i_MIPS/n214 ), .B1(net108190), .A0N(n10863), .A1N(
        n5545), .Y(\i_MIPS/N57 ) );
  OAI2BB2XL U9851 ( .B0(\i_MIPS/n230 ), .B1(net108200), .A0N(n5545), .A1N(
        n3865), .Y(\i_MIPS/N73 ) );
  OAI2BB2XL U9852 ( .B0(\i_MIPS/n229 ), .B1(net108200), .A0N(n4072), .A1N(
        n10611), .Y(\i_MIPS/N72 ) );
  OAI2BB2XL U9853 ( .B0(\i_MIPS/n242 ), .B1(net108190), .A0N(n5545), .A1N(
        n2016), .Y(\i_MIPS/N96 ) );
  AOI221X2 U9854 ( .A0(n4507), .A1(\D_cache/cache[0][140] ), .B0(n4508), .B1(
        \D_cache/cache[1][140] ), .C0(n3403), .Y(n4506) );
  NAND2XL U9855 ( .A(net112415), .B(\i_MIPS/ALU/N303 ), .Y(n6698) );
  NAND2XL U9856 ( .A(net112415), .B(n6694), .Y(n6697) );
  AOI2BB1XL U9857 ( .A0N(n9164), .A1N(n3838), .B0(n7887), .Y(n6699) );
  NAND4X1 U9858 ( .A(n8922), .B(n8921), .C(n8920), .D(n8919), .Y(n8927) );
  NAND4X1 U9859 ( .A(n7071), .B(n7070), .C(n7069), .D(n7068), .Y(n7076) );
  NAND4X1 U9860 ( .A(n8133), .B(n8132), .C(n8131), .D(n8130), .Y(n8138) );
  NAND4X1 U9861 ( .A(n8279), .B(n8278), .C(n8277), .D(n8276), .Y(n8284) );
  OA22X1 U9862 ( .A0(\i_MIPS/Register/register[5][24] ), .A1(net112222), .B0(
        \i_MIPS/Register/register[13][24] ), .B1(net112236), .Y(n8278) );
  OA22X1 U9863 ( .A0(\i_MIPS/Register/register[1][24] ), .A1(net112254), .B0(
        \i_MIPS/Register/register[9][24] ), .B1(n151), .Y(n8279) );
  OA22X1 U9864 ( .A0(\i_MIPS/Register/register[7][24] ), .A1(net112150), .B0(
        \i_MIPS/Register/register[15][24] ), .B1(net112170), .Y(n8276) );
  NAND4X1 U9865 ( .A(n9120), .B(n9119), .C(n9118), .D(n9117), .Y(n9125) );
  OA22X1 U9866 ( .A0(\i_MIPS/Register/register[1][21] ), .A1(net112260), .B0(
        \i_MIPS/Register/register[9][21] ), .B1(n147), .Y(n9120) );
  OA22X1 U9867 ( .A0(\i_MIPS/Register/register[7][21] ), .A1(net112152), .B0(
        \i_MIPS/Register/register[15][21] ), .B1(net112172), .Y(n9117) );
  NAND4X1 U9868 ( .A(n8370), .B(n8369), .C(n8368), .D(n8367), .Y(n8375) );
  OA22X1 U9869 ( .A0(\i_MIPS/Register/register[5][3] ), .A1(net112222), .B0(
        \i_MIPS/Register/register[13][3] ), .B1(net112236), .Y(n8369) );
  OA22X1 U9870 ( .A0(\i_MIPS/Register/register[1][3] ), .A1(net112258), .B0(
        \i_MIPS/Register/register[9][3] ), .B1(n151), .Y(n8370) );
  OA22X1 U9871 ( .A0(\i_MIPS/Register/register[7][3] ), .A1(net112150), .B0(
        \i_MIPS/Register/register[15][3] ), .B1(net112170), .Y(n8367) );
  NAND4X1 U9872 ( .A(n8468), .B(n8467), .C(n8466), .D(n8465), .Y(n8473) );
  OA22X1 U9873 ( .A0(\i_MIPS/Register/register[5][28] ), .A1(net112224), .B0(
        \i_MIPS/Register/register[13][28] ), .B1(net112244), .Y(n8467) );
  OA22X1 U9874 ( .A0(\i_MIPS/Register/register[1][28] ), .A1(net112260), .B0(
        \i_MIPS/Register/register[9][28] ), .B1(n148), .Y(n8468) );
  OA22X1 U9875 ( .A0(\i_MIPS/Register/register[7][28] ), .A1(net112152), .B0(
        \i_MIPS/Register/register[15][28] ), .B1(net112170), .Y(n8465) );
  NAND4X1 U9876 ( .A(n7383), .B(n7382), .C(n7381), .D(n7380), .Y(n7388) );
  NAND4X1 U9877 ( .A(n9225), .B(n9224), .C(n9223), .D(n9222), .Y(n9230) );
  OA22X1 U9878 ( .A0(\i_MIPS/Register/register[1][20] ), .A1(net112254), .B0(
        \i_MIPS/Register/register[9][20] ), .B1(n148), .Y(n9225) );
  OA22X1 U9879 ( .A0(\i_MIPS/Register/register[7][20] ), .A1(net112152), .B0(
        \i_MIPS/Register/register[15][20] ), .B1(net112172), .Y(n9222) );
  NAND4X1 U9880 ( .A(n7628), .B(n7627), .C(n7626), .D(n7625), .Y(n7633) );
  OA22X1 U9881 ( .A0(\i_MIPS/Register/register[5][14] ), .A1(net112222), .B0(
        \i_MIPS/Register/register[13][14] ), .B1(net112244), .Y(n7627) );
  OA22X1 U9882 ( .A0(\i_MIPS/Register/register[1][14] ), .A1(net112254), .B0(
        \i_MIPS/Register/register[9][14] ), .B1(n147), .Y(n7628) );
  OA22X1 U9883 ( .A0(\i_MIPS/Register/register[7][14] ), .A1(net112148), .B0(
        \i_MIPS/Register/register[15][14] ), .B1(net112166), .Y(n7625) );
  NAND4X1 U9884 ( .A(n9023), .B(n9022), .C(n9021), .D(n9020), .Y(n9028) );
  OA22X1 U9885 ( .A0(\i_MIPS/Register/register[5][25] ), .A1(net112224), .B0(
        \i_MIPS/Register/register[13][25] ), .B1(net112236), .Y(n9022) );
  OA22X1 U9886 ( .A0(\i_MIPS/Register/register[1][25] ), .A1(net112258), .B0(
        \i_MIPS/Register/register[9][25] ), .B1(n150), .Y(n9023) );
  OA22X1 U9887 ( .A0(\i_MIPS/Register/register[7][25] ), .A1(net112152), .B0(
        \i_MIPS/Register/register[15][25] ), .B1(net112170), .Y(n9020) );
  NAND4X1 U9888 ( .A(n7721), .B(n7720), .C(n7719), .D(n7718), .Y(n7726) );
  OA22X1 U9889 ( .A0(\i_MIPS/Register/register[5][13] ), .A1(net112222), .B0(
        \i_MIPS/Register/register[13][13] ), .B1(net112242), .Y(n7720) );
  OA22X1 U9890 ( .A0(\i_MIPS/Register/register[7][13] ), .A1(net112148), .B0(
        \i_MIPS/Register/register[15][13] ), .B1(net112166), .Y(n7718) );
  NAND4X1 U9891 ( .A(n7992), .B(n7991), .C(n7990), .D(n7989), .Y(n7997) );
  NAND4X1 U9892 ( .A(n8050), .B(n8049), .C(n8048), .D(n8047), .Y(n8055) );
  NAND4X1 U9893 ( .A(n7130), .B(n7129), .C(n7128), .D(n7127), .Y(n7135) );
  NAND4X1 U9894 ( .A(n7247), .B(n7246), .C(n7245), .D(n7244), .Y(n7252) );
  OA22X1 U9895 ( .A0(\i_MIPS/Register/register[5][11] ), .A1(net112222), .B0(
        \i_MIPS/Register/register[13][11] ), .B1(net112240), .Y(n7246) );
  OA22X1 U9896 ( .A0(\i_MIPS/Register/register[1][11] ), .A1(net112260), .B0(
        \i_MIPS/Register/register[9][11] ), .B1(n150), .Y(n7247) );
  OA22X1 U9897 ( .A0(\i_MIPS/Register/register[7][11] ), .A1(net112148), .B0(
        \i_MIPS/Register/register[15][11] ), .B1(net112166), .Y(n7244) );
  NAND4X1 U9898 ( .A(n6987), .B(n6986), .C(n6985), .D(n6984), .Y(n6992) );
  OA22X1 U9899 ( .A0(\i_MIPS/Register/register[5][6] ), .A1(n192), .B0(
        \i_MIPS/Register/register[13][6] ), .B1(net112236), .Y(n6986) );
  OA22X1 U9900 ( .A0(\i_MIPS/Register/register[1][6] ), .A1(net112260), .B0(
        \i_MIPS/Register/register[9][6] ), .B1(n148), .Y(n6987) );
  OA22X1 U9901 ( .A0(\i_MIPS/Register/register[7][6] ), .A1(net112152), .B0(
        \i_MIPS/Register/register[15][6] ), .B1(net112164), .Y(n6984) );
  NAND4X1 U9902 ( .A(n6781), .B(n6780), .C(n6779), .D(n6778), .Y(n6786) );
  OA22X1 U9903 ( .A0(\i_MIPS/Register/register[5][5] ), .A1(n192), .B0(
        \i_MIPS/Register/register[13][5] ), .B1(net112242), .Y(n6780) );
  OA22X1 U9904 ( .A0(\i_MIPS/Register/register[1][5] ), .A1(net112258), .B0(
        \i_MIPS/Register/register[9][5] ), .B1(n150), .Y(n6781) );
  OA22X1 U9905 ( .A0(\i_MIPS/Register/register[7][5] ), .A1(net112152), .B0(
        \i_MIPS/Register/register[15][5] ), .B1(net112164), .Y(n6778) );
  NAND4X1 U9906 ( .A(n6862), .B(n6861), .C(n6860), .D(n6859), .Y(n6867) );
  OA22X1 U9907 ( .A0(\i_MIPS/Register/register[5][4] ), .A1(n192), .B0(
        \i_MIPS/Register/register[13][4] ), .B1(net112236), .Y(n6861) );
  OA22X1 U9908 ( .A0(\i_MIPS/Register/register[1][4] ), .A1(net112260), .B0(
        \i_MIPS/Register/register[9][4] ), .B1(n151), .Y(n6862) );
  OA22X1 U9909 ( .A0(\i_MIPS/Register/register[7][4] ), .A1(net112148), .B0(
        \i_MIPS/Register/register[15][4] ), .B1(net112164), .Y(n6859) );
  NAND4X1 U9910 ( .A(n7913), .B(n7912), .C(n7911), .D(n7910), .Y(n7918) );
  NAND4X1 U9911 ( .A(n7780), .B(n7779), .C(n7778), .D(n7777), .Y(n7785) );
  NAND4X1 U9912 ( .A(n7555), .B(n7554), .C(n7553), .D(n7552), .Y(n7560) );
  OA22X1 U9913 ( .A0(\i_MIPS/Register/register[5][0] ), .A1(net112222), .B0(
        \i_MIPS/Register/register[13][0] ), .B1(net112240), .Y(n7554) );
  OA22X1 U9914 ( .A0(\i_MIPS/Register/register[1][0] ), .A1(net112260), .B0(
        \i_MIPS/Register/register[9][0] ), .B1(n151), .Y(n7555) );
  OA22X1 U9915 ( .A0(\i_MIPS/Register/register[7][0] ), .A1(net112148), .B0(
        \i_MIPS/Register/register[15][0] ), .B1(net112166), .Y(n7552) );
  OA22X1 U9916 ( .A0(\i_MIPS/Register/register[5][10] ), .A1(net112222), .B0(
        \i_MIPS/Register/register[13][10] ), .B1(net112236), .Y(n7325) );
  OA22X1 U9917 ( .A0(\i_MIPS/Register/register[7][10] ), .A1(net112148), .B0(
        \i_MIPS/Register/register[15][10] ), .B1(net112166), .Y(n7323) );
  OA22X1 U9918 ( .A0(\i_MIPS/Register/register[5][9] ), .A1(net112224), .B0(
        \i_MIPS/Register/register[13][9] ), .B1(net112236), .Y(n8665) );
  OA22X1 U9919 ( .A0(\i_MIPS/Register/register[1][9] ), .A1(net112254), .B0(
        \i_MIPS/Register/register[9][9] ), .B1(n147), .Y(n8666) );
  OA22X1 U9920 ( .A0(\i_MIPS/Register/register[7][9] ), .A1(net112152), .B0(
        \i_MIPS/Register/register[15][9] ), .B1(net112170), .Y(n8663) );
  NAND4X1 U9921 ( .A(n8831), .B(n8830), .C(n8829), .D(n8828), .Y(n8836) );
  OA22X1 U9922 ( .A0(\i_MIPS/Register/register[5][23] ), .A1(net112224), .B0(
        \i_MIPS/Register/register[13][23] ), .B1(net112240), .Y(n8830) );
  OA22X1 U9923 ( .A0(\i_MIPS/Register/register[1][23] ), .A1(net112260), .B0(
        \i_MIPS/Register/register[9][23] ), .B1(n147), .Y(n8831) );
  OA22X1 U9924 ( .A0(\i_MIPS/Register/register[7][23] ), .A1(net112152), .B0(
        \i_MIPS/Register/register[15][23] ), .B1(net112170), .Y(n8828) );
  NAND4X1 U9925 ( .A(n8768), .B(n8767), .C(n8766), .D(n8765), .Y(n8773) );
  OA22X1 U9926 ( .A0(\i_MIPS/Register/register[5][18] ), .A1(net112224), .B0(
        \i_MIPS/Register/register[13][18] ), .B1(net112236), .Y(n8767) );
  OA22X1 U9927 ( .A0(\i_MIPS/Register/register[1][18] ), .A1(net112258), .B0(
        \i_MIPS/Register/register[9][18] ), .B1(n151), .Y(n8768) );
  OA22X1 U9928 ( .A0(\i_MIPS/Register/register[7][18] ), .A1(net112152), .B0(
        \i_MIPS/Register/register[15][18] ), .B1(net112170), .Y(n8765) );
  NAND4X1 U9929 ( .A(n9436), .B(n9435), .C(n9434), .D(n9433), .Y(n9441) );
  NAND4X1 U9930 ( .A(n6662), .B(n6661), .C(n6660), .D(n6659), .Y(n6667) );
  OA22X1 U9931 ( .A0(\i_MIPS/Register/register[0][20] ), .A1(n4702), .B0(
        \i_MIPS/Register/register[8][20] ), .B1(n4700), .Y(n9310) );
  OA22X1 U9932 ( .A0(\i_MIPS/Register/register[4][20] ), .A1(n4697), .B0(
        \i_MIPS/Register/register[12][20] ), .B1(n4693), .Y(n9311) );
  OAI221XL U9933 ( .A0(\i_MIPS/Register/register[2][20] ), .A1(n4690), .B0(
        \i_MIPS/Register/register[10][20] ), .B1(n4686), .C0(n9304), .Y(n9312)
         );
  OA22X1 U9934 ( .A0(\i_MIPS/Register/register[4][1] ), .A1(n4698), .B0(
        \i_MIPS/Register/register[12][1] ), .B1(n4694), .Y(n8034) );
  OA22X1 U9935 ( .A0(\i_MIPS/Register/register[0][1] ), .A1(n4703), .B0(
        \i_MIPS/Register/register[8][1] ), .B1(n4701), .Y(n8033) );
  NAND4BX1 U9936 ( .AN(n7765), .B(n7764), .C(n7763), .D(n7762), .Y(n7776) );
  OA22X1 U9937 ( .A0(\i_MIPS/Register/register[4][13] ), .A1(n4699), .B0(
        \i_MIPS/Register/register[12][13] ), .B1(n4695), .Y(n7764) );
  OA22X1 U9938 ( .A0(\i_MIPS/Register/register[0][13] ), .A1(n4703), .B0(
        \i_MIPS/Register/register[8][13] ), .B1(n4701), .Y(n7763) );
  OAI221XL U9939 ( .A0(\i_MIPS/Register/register[2][13] ), .A1(n4692), .B0(
        \i_MIPS/Register/register[10][13] ), .B1(n4687), .C0(n7757), .Y(n7765)
         );
  OAI221XL U9940 ( .A0(\i_MIPS/Register/register[2][21] ), .A1(n4690), .B0(
        \i_MIPS/Register/register[10][21] ), .B1(n4686), .C0(n9198), .Y(n9206)
         );
  NAND4BX1 U9941 ( .AN(n9523), .B(n9522), .C(n9521), .D(n9520), .Y(n9545) );
  OAI221XL U9942 ( .A0(\i_MIPS/Register/register[2][22] ), .A1(n4690), .B0(
        \i_MIPS/Register/register[10][22] ), .B1(n4686), .C0(n9515), .Y(n9523)
         );
  NAND4BX1 U9943 ( .AN(n7671), .B(n7670), .C(n7669), .D(n7668), .Y(n7682) );
  OA22X1 U9944 ( .A0(\i_MIPS/Register/register[4][14] ), .A1(n4699), .B0(
        \i_MIPS/Register/register[12][14] ), .B1(n4695), .Y(n7670) );
  OA22X1 U9945 ( .A0(\i_MIPS/Register/register[0][14] ), .A1(n4703), .B0(
        \i_MIPS/Register/register[8][14] ), .B1(n4701), .Y(n7669) );
  OAI221XL U9946 ( .A0(\i_MIPS/Register/register[2][14] ), .A1(n4692), .B0(
        \i_MIPS/Register/register[10][14] ), .B1(n4687), .C0(n7663), .Y(n7671)
         );
  NAND4BX1 U9947 ( .AN(n8118), .B(n8117), .C(n8116), .D(n8115), .Y(n8129) );
  OA22X1 U9948 ( .A0(\i_MIPS/Register/register[4][16] ), .A1(n4698), .B0(
        \i_MIPS/Register/register[12][16] ), .B1(n4694), .Y(n8117) );
  OA22X1 U9949 ( .A0(\i_MIPS/Register/register[0][16] ), .A1(n4703), .B0(
        \i_MIPS/Register/register[8][16] ), .B1(n4701), .Y(n8116) );
  OAI221XL U9950 ( .A0(\i_MIPS/Register/register[2][16] ), .A1(n4691), .B0(
        \i_MIPS/Register/register[10][16] ), .B1(n4687), .C0(n8110), .Y(n8118)
         );
  NAND4BX1 U9951 ( .AN(n6950), .B(n6949), .C(n6948), .D(n6947), .Y(n6961) );
  OA22X1 U9952 ( .A0(\i_MIPS/Register/register[4][2] ), .A1(n4698), .B0(
        \i_MIPS/Register/register[12][2] ), .B1(n4695), .Y(n6949) );
  OA22X1 U9953 ( .A0(\i_MIPS/Register/register[0][2] ), .A1(n4704), .B0(
        \i_MIPS/Register/register[8][2] ), .B1(n4700), .Y(n6948) );
  NAND4BX1 U9954 ( .AN(n8213), .B(n8212), .C(n8211), .D(n8210), .Y(n8224) );
  OA22X1 U9955 ( .A0(\i_MIPS/Register/register[4][29] ), .A1(n4698), .B0(
        \i_MIPS/Register/register[12][29] ), .B1(n4694), .Y(n8212) );
  OA22X1 U9956 ( .A0(\i_MIPS/Register/register[0][29] ), .A1(n4703), .B0(
        \i_MIPS/Register/register[8][29] ), .B1(n4701), .Y(n8211) );
  OAI221XL U9957 ( .A0(\i_MIPS/Register/register[2][29] ), .A1(n4691), .B0(
        \i_MIPS/Register/register[10][29] ), .B1(n4688), .C0(n8205), .Y(n8213)
         );
  OA22X1 U9958 ( .A0(\i_MIPS/Register/register[4][6] ), .A1(n4699), .B0(
        \i_MIPS/Register/register[12][6] ), .B1(n4695), .Y(n7029) );
  OA22X1 U9959 ( .A0(\i_MIPS/Register/register[0][6] ), .A1(n4704), .B0(
        \i_MIPS/Register/register[8][6] ), .B1(n4700), .Y(n7028) );
  OAI221XL U9960 ( .A0(\i_MIPS/Register/register[2][6] ), .A1(n4692), .B0(
        \i_MIPS/Register/register[10][6] ), .B1(n4688), .C0(n7022), .Y(n7030)
         );
  OA22X1 U9961 ( .A0(\i_MIPS/Register/register[4][28] ), .A1(n4698), .B0(
        \i_MIPS/Register/register[12][28] ), .B1(n4694), .Y(n8512) );
  OA22X1 U9962 ( .A0(\i_MIPS/Register/register[0][28] ), .A1(n4703), .B0(
        \i_MIPS/Register/register[8][28] ), .B1(n4701), .Y(n8511) );
  OAI221XL U9963 ( .A0(\i_MIPS/Register/register[2][28] ), .A1(n4691), .B0(
        \i_MIPS/Register/register[10][28] ), .B1(n4688), .C0(n8505), .Y(n8513)
         );
  NAND4BX1 U9964 ( .AN(n8414), .B(n8413), .C(n8412), .D(n8411), .Y(n8425) );
  OA22X1 U9965 ( .A0(\i_MIPS/Register/register[4][3] ), .A1(n4698), .B0(
        \i_MIPS/Register/register[12][3] ), .B1(n4694), .Y(n8413) );
  OA22X1 U9966 ( .A0(\i_MIPS/Register/register[0][3] ), .A1(n4703), .B0(
        \i_MIPS/Register/register[8][3] ), .B1(n4701), .Y(n8412) );
  OAI221XL U9967 ( .A0(\i_MIPS/Register/register[2][3] ), .A1(n4691), .B0(
        \i_MIPS/Register/register[10][3] ), .B1(n4688), .C0(n8406), .Y(n8414)
         );
  OAI221XL U9968 ( .A0(\i_MIPS/Register/register[2][8] ), .A1(n4692), .B0(
        \i_MIPS/Register/register[10][8] ), .B1(n4688), .C0(n7107), .Y(n7115)
         );
  NAND4BX1 U9969 ( .AN(n7451), .B(n7450), .C(n7449), .D(n7448), .Y(n7462) );
  OA22X1 U9970 ( .A0(\i_MIPS/Register/register[4][12] ), .A1(n4699), .B0(
        \i_MIPS/Register/register[12][12] ), .B1(n4695), .Y(n7450) );
  OA22X1 U9971 ( .A0(\i_MIPS/Register/register[0][12] ), .A1(n4704), .B0(
        \i_MIPS/Register/register[8][12] ), .B1(n4700), .Y(n7449) );
  NAND4BX1 U9972 ( .AN(n8323), .B(n8322), .C(n8321), .D(n8320), .Y(n8334) );
  OA22X1 U9973 ( .A0(\i_MIPS/Register/register[4][24] ), .A1(n4698), .B0(
        \i_MIPS/Register/register[12][24] ), .B1(n4694), .Y(n8322) );
  OA22X1 U9974 ( .A0(\i_MIPS/Register/register[0][24] ), .A1(n4703), .B0(
        \i_MIPS/Register/register[8][24] ), .B1(n4701), .Y(n8321) );
  OAI221XL U9975 ( .A0(\i_MIPS/Register/register[2][24] ), .A1(n4691), .B0(
        \i_MIPS/Register/register[10][24] ), .B1(n4687), .C0(n8315), .Y(n8323)
         );
  NAND4BX1 U9976 ( .AN(n6825), .B(n6824), .C(n6823), .D(n6822), .Y(n6836) );
  OA22X1 U9977 ( .A0(\i_MIPS/Register/register[4][5] ), .A1(n4698), .B0(
        \i_MIPS/Register/register[12][5] ), .B1(n4695), .Y(n6824) );
  OA22X1 U9978 ( .A0(\i_MIPS/Register/register[0][5] ), .A1(n4704), .B0(
        \i_MIPS/Register/register[8][5] ), .B1(n4700), .Y(n6823) );
  OAI221XL U9979 ( .A0(\i_MIPS/Register/register[2][5] ), .A1(n4690), .B0(
        \i_MIPS/Register/register[10][5] ), .B1(n4688), .C0(n6817), .Y(n6825)
         );
  NAND4BX1 U9980 ( .AN(n9005), .B(n9004), .C(n9003), .D(n9002), .Y(n9016) );
  OA22X1 U9981 ( .A0(\i_MIPS/Register/register[0][26] ), .A1(n4702), .B0(
        \i_MIPS/Register/register[8][26] ), .B1(n4700), .Y(n9003) );
  OA22X1 U9982 ( .A0(\i_MIPS/Register/register[4][26] ), .A1(n4697), .B0(
        \i_MIPS/Register/register[12][26] ), .B1(n4693), .Y(n9004) );
  NAND4BX1 U9983 ( .AN(n6630), .B(n6629), .C(n6628), .D(n6627), .Y(n6631) );
  NAND4BX1 U9984 ( .AN(n9321), .B(n9320), .C(n9319), .D(n9318), .Y(n9322) );
  OA22X1 U9985 ( .A0(\i_MIPS/Register/register[16][20] ), .A1(n4702), .B0(
        \i_MIPS/Register/register[24][20] ), .B1(n4700), .Y(n9319) );
  OA22X1 U9986 ( .A0(\i_MIPS/Register/register[20][20] ), .A1(n4697), .B0(
        \i_MIPS/Register/register[28][20] ), .B1(n4693), .Y(n9320) );
  OAI221XL U9987 ( .A0(\i_MIPS/Register/register[18][20] ), .A1(n4690), .B0(
        \i_MIPS/Register/register[26][20] ), .B1(n4686), .C0(n9313), .Y(n9321)
         );
  OAI221XL U9988 ( .A0(\i_MIPS/Register/register[18][1] ), .A1(n4692), .B0(
        \i_MIPS/Register/register[26][1] ), .B1(n4687), .C0(n8036), .Y(n8044)
         );
  OA22XL U9989 ( .A0(\i_MIPS/Register/register[20][19] ), .A1(net102050), .B0(
        \i_MIPS/Register/register[28][19] ), .B1(net102051), .Y(n8583) );
  OA22XL U9990 ( .A0(\i_MIPS/Register/register[16][19] ), .A1(net102048), .B0(
        \i_MIPS/Register/register[24][19] ), .B1(net102049), .Y(n8582) );
  NAND4BX1 U9991 ( .AN(n9215), .B(n9214), .C(n9213), .D(n9212), .Y(n9216) );
  OAI221XL U9992 ( .A0(\i_MIPS/Register/register[18][21] ), .A1(n4690), .B0(
        \i_MIPS/Register/register[26][21] ), .B1(n4686), .C0(n9207), .Y(n9215)
         );
  NAND4BX1 U9993 ( .AN(n7774), .B(n7773), .C(n7772), .D(n7771), .Y(n7775) );
  OAI221XL U9994 ( .A0(\i_MIPS/Register/register[18][13] ), .A1(n4692), .B0(
        \i_MIPS/Register/register[26][13] ), .B1(n4687), .C0(n7766), .Y(n7774)
         );
  NAND4BX1 U9995 ( .AN(n9543), .B(n9542), .C(n9541), .D(n9540), .Y(n9544) );
  OA22X1 U9996 ( .A0(\i_MIPS/Register/register[20][22] ), .A1(n4698), .B0(
        \i_MIPS/Register/register[28][22] ), .B1(n4694), .Y(n9542) );
  OA22X1 U9997 ( .A0(\i_MIPS/Register/register[16][22] ), .A1(n4703), .B0(
        \i_MIPS/Register/register[24][22] ), .B1(n4701), .Y(n9541) );
  OAI221XL U9998 ( .A0(\i_MIPS/Register/register[18][22] ), .A1(n4692), .B0(
        \i_MIPS/Register/register[26][22] ), .B1(n4687), .C0(n9526), .Y(n9543)
         );
  NAND4BX1 U9999 ( .AN(n7680), .B(n7679), .C(n7678), .D(n7677), .Y(n7681) );
  OAI221XL U10000 ( .A0(\i_MIPS/Register/register[18][14] ), .A1(n4692), .B0(
        \i_MIPS/Register/register[26][14] ), .B1(n4687), .C0(n7672), .Y(n7680)
         );
  NAND4BX1 U10001 ( .AN(n8127), .B(n8126), .C(n8125), .D(n8124), .Y(n8128) );
  OAI221XL U10002 ( .A0(\i_MIPS/Register/register[18][16] ), .A1(n4691), .B0(
        \i_MIPS/Register/register[26][16] ), .B1(n4687), .C0(n8119), .Y(n8127)
         );
  OA22X1 U10003 ( .A0(\i_MIPS/Register/register[20][2] ), .A1(n4699), .B0(
        \i_MIPS/Register/register[28][2] ), .B1(n4695), .Y(n6958) );
  OA22X1 U10004 ( .A0(\i_MIPS/Register/register[16][2] ), .A1(n4704), .B0(
        \i_MIPS/Register/register[24][2] ), .B1(n4700), .Y(n6957) );
  NAND4BX1 U10005 ( .AN(n8222), .B(n8221), .C(n8220), .D(n8219), .Y(n8223) );
  OAI221XL U10006 ( .A0(\i_MIPS/Register/register[18][29] ), .A1(n4691), .B0(
        \i_MIPS/Register/register[26][29] ), .B1(n4688), .C0(n8214), .Y(n8222)
         );
  OA22X1 U10007 ( .A0(\i_MIPS/Register/register[20][6] ), .A1(n4699), .B0(
        \i_MIPS/Register/register[28][6] ), .B1(n4695), .Y(n7038) );
  OA22X1 U10008 ( .A0(\i_MIPS/Register/register[16][6] ), .A1(n4704), .B0(
        \i_MIPS/Register/register[24][6] ), .B1(n4700), .Y(n7037) );
  OAI221XL U10009 ( .A0(\i_MIPS/Register/register[18][6] ), .A1(n4691), .B0(
        \i_MIPS/Register/register[26][6] ), .B1(n4688), .C0(n7031), .Y(n7039)
         );
  NAND4BX1 U10010 ( .AN(n8522), .B(n8521), .C(n8520), .D(n8519), .Y(n8523) );
  OA22X1 U10011 ( .A0(\i_MIPS/Register/register[20][28] ), .A1(n4698), .B0(
        \i_MIPS/Register/register[28][28] ), .B1(n4694), .Y(n8521) );
  OA22X1 U10012 ( .A0(\i_MIPS/Register/register[16][28] ), .A1(n4703), .B0(
        \i_MIPS/Register/register[24][28] ), .B1(n4701), .Y(n8520) );
  NAND4BX1 U10013 ( .AN(n8423), .B(n8422), .C(n8421), .D(n8420), .Y(n8424) );
  OAI221XL U10014 ( .A0(\i_MIPS/Register/register[18][3] ), .A1(n4691), .B0(
        \i_MIPS/Register/register[26][3] ), .B1(n4687), .C0(n8415), .Y(n8423)
         );
  NAND4BX1 U10015 ( .AN(n7460), .B(n7459), .C(n7458), .D(n7457), .Y(n7461) );
  OAI221XL U10016 ( .A0(\i_MIPS/Register/register[18][12] ), .A1(n4692), .B0(
        \i_MIPS/Register/register[26][12] ), .B1(n4687), .C0(n7452), .Y(n7460)
         );
  NAND4BX1 U10017 ( .AN(n8332), .B(n8331), .C(n8330), .D(n8329), .Y(n8333) );
  OAI221XL U10018 ( .A0(\i_MIPS/Register/register[18][24] ), .A1(n4691), .B0(
        \i_MIPS/Register/register[26][24] ), .B1(n4688), .C0(n8324), .Y(n8332)
         );
  NAND4BX1 U10019 ( .AN(n8624), .B(n8623), .C(n8622), .D(n8621), .Y(n8625) );
  OA22X1 U10020 ( .A0(\i_MIPS/Register/register[20][19] ), .A1(n4698), .B0(
        \i_MIPS/Register/register[28][19] ), .B1(n4694), .Y(n8623) );
  OAI221XL U10021 ( .A0(\i_MIPS/Register/register[18][19] ), .A1(n4691), .B0(
        \i_MIPS/Register/register[26][19] ), .B1(n4688), .C0(n8616), .Y(n8624)
         );
  NAND4BX1 U10022 ( .AN(n6834), .B(n6833), .C(n6832), .D(n6831), .Y(n6835) );
  OAI221XL U10023 ( .A0(\i_MIPS/Register/register[18][5] ), .A1(n4692), .B0(
        \i_MIPS/Register/register[26][5] ), .B1(n4688), .C0(n6826), .Y(n6834)
         );
  OA22X1 U10024 ( .A0(\i_MIPS/Register/register[16][26] ), .A1(n4702), .B0(
        \i_MIPS/Register/register[24][26] ), .B1(n4700), .Y(n9012) );
  OA22X1 U10025 ( .A0(\i_MIPS/Register/register[20][26] ), .A1(n4697), .B0(
        \i_MIPS/Register/register[28][26] ), .B1(n4693), .Y(n9013) );
  OAI221XL U10026 ( .A0(\i_MIPS/Register/register[18][26] ), .A1(n4690), .B0(
        \i_MIPS/Register/register[26][26] ), .B1(n4686), .C0(n9006), .Y(n9014)
         );
  INVX1 U10027 ( .A(n6483), .Y(n8960) );
  MXI2XL U10028 ( .A(\i_MIPS/n361 ), .B(n4430), .S0(n205), .Y(\i_MIPS/n552 )
         );
  OA22X1 U10029 ( .A0(\i_MIPS/PHT_2/n3 ), .A1(n11047), .B0(\i_MIPS/PHT_2/n7 ), 
        .B1(n11046), .Y(n10352) );
  AOI32X1 U10030 ( .A0(n406), .A1(\i_MIPS/PHT_2/history_state[0] ), .A2(
        \i_MIPS/PHT_2/history_state[1] ), .B0(n270), .B1(
        \i_MIPS/PHT_2/current_state_2[1] ), .Y(n10353) );
  MXI2XL U10031 ( .A(\i_MIPS/n344 ), .B(n10838), .S0(n216), .Y(\i_MIPS/n535 )
         );
  MXI2X1 U10032 ( .A(\i_MIPS/n355 ), .B(net128955), .S0(n223), .Y(
        \i_MIPS/n546 ) );
  MXI2X1 U10033 ( .A(\i_MIPS/n360 ), .B(n4396), .S0(n220), .Y(\i_MIPS/n551 )
         );
  MXI2X1 U10034 ( .A(\i_MIPS/n367 ), .B(n4408), .S0(n216), .Y(\i_MIPS/n558 )
         );
  MXI2X1 U10035 ( .A(\i_MIPS/n366 ), .B(n4407), .S0(n210), .Y(\i_MIPS/n557 )
         );
  MXI2X1 U10036 ( .A(\i_MIPS/n365 ), .B(n4406), .S0(n207), .Y(\i_MIPS/n556 )
         );
  MXI2X1 U10037 ( .A(\i_MIPS/n364 ), .B(n4405), .S0(n208), .Y(\i_MIPS/n555 )
         );
  MXI2X1 U10038 ( .A(\i_MIPS/n363 ), .B(n4431), .S0(n205), .Y(\i_MIPS/n554 )
         );
  MXI2X1 U10039 ( .A(\i_MIPS/n362 ), .B(n4404), .S0(n219), .Y(\i_MIPS/n553 )
         );
  MXI2X1 U10040 ( .A(\i_MIPS/n359 ), .B(n4403), .S0(n222), .Y(\i_MIPS/n550 )
         );
  MXI2XL U10041 ( .A(\i_MIPS/n358 ), .B(n4402), .S0(n223), .Y(\i_MIPS/n549 )
         );
  MXI2XL U10042 ( .A(\i_MIPS/n357 ), .B(n4401), .S0(n204), .Y(\i_MIPS/n548 )
         );
  MXI2X1 U10043 ( .A(\i_MIPS/n356 ), .B(n4400), .S0(n220), .Y(\i_MIPS/n547 )
         );
  MXI2XL U10044 ( .A(\i_MIPS/n354 ), .B(n4429), .S0(n223), .Y(\i_MIPS/n545 )
         );
  MXI2XL U10045 ( .A(\i_MIPS/n353 ), .B(n4399), .S0(n217), .Y(\i_MIPS/n544 )
         );
  MXI2X1 U10046 ( .A(\i_MIPS/n350 ), .B(n4427), .S0(n207), .Y(\i_MIPS/n541 )
         );
  MXI2X1 U10047 ( .A(\i_MIPS/n352 ), .B(n11007), .S0(n208), .Y(\i_MIPS/n543 )
         );
  MXI2XL U10048 ( .A(\i_MIPS/n341 ), .B(n10796), .S0(n220), .Y(\i_MIPS/n532 )
         );
  MXI2XL U10049 ( .A(\i_MIPS/n343 ), .B(n4414), .S0(n207), .Y(\i_MIPS/n534 )
         );
  MXI2XL U10050 ( .A(\i_MIPS/n371 ), .B(n4432), .S0(n210), .Y(\i_MIPS/n562 )
         );
  MXI2XL U10051 ( .A(\i_MIPS/n294 ), .B(\i_MIPS/n295 ), .S0(n211), .Y(
        \i_MIPS/n422 ) );
  MXI2X1 U10052 ( .A(\i_MIPS/PHT_2/n2 ), .B(n11049), .S0(n11048), .Y(
        \i_MIPS/PHT_2/n45 ) );
  MXI2XL U10053 ( .A(\i_MIPS/n313 ), .B(\i_MIPS/n312 ), .S0(n210), .Y(
        \i_MIPS/n513 ) );
  MXI2X1 U10054 ( .A(\i_MIPS/n296 ), .B(\i_MIPS/n297 ), .S0(n220), .Y(
        \i_MIPS/n424 ) );
  MXI2X1 U10055 ( .A(\i_MIPS/n264 ), .B(\i_MIPS/n265 ), .S0(n222), .Y(
        \i_MIPS/n392 ) );
  MXI2XL U10056 ( .A(\i_MIPS/n334 ), .B(\i_MIPS/n335 ), .S0(n213), .Y(
        \i_MIPS/n524 ) );
  MXI2XL U10057 ( .A(\i_MIPS/n325 ), .B(\i_MIPS/n324 ), .S0(n219), .Y(
        \i_MIPS/n519 ) );
  MXI2X1 U10058 ( .A(\i_MIPS/n308 ), .B(\i_MIPS/n309 ), .S0(n223), .Y(
        \i_MIPS/n436 ) );
  MXI2X1 U10059 ( .A(\i_MIPS/n306 ), .B(\i_MIPS/n307 ), .S0(n210), .Y(
        \i_MIPS/n434 ) );
  MXI2X1 U10060 ( .A(\i_MIPS/n304 ), .B(\i_MIPS/n305 ), .S0(n204), .Y(
        \i_MIPS/n432 ) );
  MXI2X1 U10061 ( .A(\i_MIPS/n292 ), .B(\i_MIPS/n293 ), .S0(n211), .Y(
        \i_MIPS/n420 ) );
  MXI2X1 U10062 ( .A(\i_MIPS/n290 ), .B(\i_MIPS/n291 ), .S0(n213), .Y(
        \i_MIPS/n418 ) );
  MXI2X1 U10063 ( .A(\i_MIPS/n262 ), .B(\i_MIPS/n263 ), .S0(n216), .Y(
        \i_MIPS/n390 ) );
  MXI2X1 U10064 ( .A(\i_MIPS/n256 ), .B(\i_MIPS/n257 ), .S0(n217), .Y(
        \i_MIPS/n384 ) );
  MXI2XL U10065 ( .A(\i_MIPS/n373 ), .B(\i_MIPS/n372 ), .S0(n204), .Y(
        \i_MIPS/n563 ) );
  MXI2XL U10066 ( .A(\i_MIPS/n338 ), .B(\i_MIPS/n339 ), .S0(n222), .Y(
        \i_MIPS/n529 ) );
  MXI2XL U10067 ( .A(\i_MIPS/n336 ), .B(\i_MIPS/n337 ), .S0(n214), .Y(
        \i_MIPS/n526 ) );
  MXI2XL U10068 ( .A(\i_MIPS/n319 ), .B(\i_MIPS/n318 ), .S0(n220), .Y(
        \i_MIPS/n516 ) );
  MXI2XL U10069 ( .A(\i_MIPS/n254 ), .B(\i_MIPS/n255 ), .S0(n207), .Y(
        \i_MIPS/n382 ) );
  MXI2XL U10070 ( .A(\i_MIPS/n252 ), .B(\i_MIPS/n253 ), .S0(n208), .Y(
        \i_MIPS/n380 ) );
  CLKINVX1 U10071 ( .A(n6768), .Y(n7984) );
  XNOR2X1 U10072 ( .A(\i_MIPS/IR_ID[25] ), .B(\i_MIPS/Reg_W[4] ), .Y(n6453) );
  NOR3X1 U10073 ( .A(\i_MIPS/Hazard_detection/n8 ), .B(
        \i_MIPS/Hazard_detection/n9 ), .C(\i_MIPS/Hazard_detection/n10 ), .Y(
        \i_MIPS/Hazard_detection/n7 ) );
  XOR2XL U10074 ( .A(\i_MIPS/IR_ID[24] ), .B(\i_MIPS/ID_EX[114] ), .Y(
        \i_MIPS/Hazard_detection/n8 ) );
  XOR2XL U10075 ( .A(\i_MIPS/IR_ID[22] ), .B(\i_MIPS/ID_EX[112] ), .Y(
        \i_MIPS/Hazard_detection/n9 ) );
  XOR2XL U10076 ( .A(\i_MIPS/IR_ID[25] ), .B(\i_MIPS/ID_EX[115] ), .Y(
        \i_MIPS/Hazard_detection/n10 ) );
  NOR3X1 U10077 ( .A(\i_MIPS/Hazard_detection/n11 ), .B(
        \i_MIPS/Hazard_detection/n12 ), .C(\i_MIPS/Hazard_detection/n13 ), .Y(
        \i_MIPS/Hazard_detection/n4 ) );
  XOR2XL U10078 ( .A(\i_MIPS/IR_ID[19] ), .B(\i_MIPS/ID_EX[114] ), .Y(
        \i_MIPS/Hazard_detection/n11 ) );
  XOR2XL U10079 ( .A(\i_MIPS/IR_ID[17] ), .B(\i_MIPS/ID_EX[112] ), .Y(
        \i_MIPS/Hazard_detection/n12 ) );
  XOR2XL U10080 ( .A(net107812), .B(\i_MIPS/ID_EX[115] ), .Y(
        \i_MIPS/Hazard_detection/n13 ) );
  INVX1 U10081 ( .A(n11043), .Y(n11045) );
  NAND3BXL U10082 ( .AN(\i_MIPS/n567 ), .B(\i_MIPS/PHT_2/counter ), .C(
        net108200), .Y(n11043) );
  AND2XL U10083 ( .A(\i_MIPS/ALU/N303 ), .B(n6694), .Y(n4509) );
  NAND2X1 U10084 ( .A(n10283), .B(ICACHE_addr[17]), .Y(n10225) );
  XOR2X1 U10085 ( .A(n10240), .B(ICACHE_addr[14]), .Y(n10615) );
  NAND2XL U10086 ( .A(n10239), .B(ICACHE_addr[13]), .Y(n10240) );
  NAND2X1 U10087 ( .A(n11056), .B(n11055), .Y(\i_MIPS/PHT_2/n46 ) );
  CLKMX2X2 U10088 ( .A(\i_MIPS/PHT_2/n5 ), .B(n11054), .S0(n4461), .Y(n11055)
         );
  NAND2XL U10089 ( .A(net112691), .B(\i_MIPS/PHT_2/current_state_2[0] ), .Y(
        n11054) );
  NAND4BX1 U10090 ( .AN(n9111), .B(n9110), .C(n9109), .D(n9108), .Y(n9112) );
  NAND4BX1 U10091 ( .AN(n7299), .B(n7298), .C(n7297), .D(n7296), .Y(net104255)
         );
  NAND4BX1 U10092 ( .AN(n7957), .B(n7956), .C(n7955), .D(n7954), .Y(net103092)
         );
  NAND4BX1 U10093 ( .AN(n7599), .B(n7598), .C(n7597), .D(n7596), .Y(net103721)
         );
  NAND4BX1 U10094 ( .AN(n7608), .B(n7607), .C(n7606), .D(n7605), .Y(net103722)
         );
  NAND4BX1 U10095 ( .AN(n7208), .B(n7207), .C(n7206), .D(n7205), .Y(net104410)
         );
  NAND4BX1 U10096 ( .AN(n7370), .B(n7369), .C(n7368), .D(n7367), .Y(net104108)
         );
  CLKMX2X2 U10097 ( .A(n8721), .B(n8720), .S0(net107810), .Y(n8724) );
  NAND4BX1 U10098 ( .AN(n8710), .B(n8709), .C(n8708), .D(n8707), .Y(n8721) );
  NAND4BX1 U10099 ( .AN(n8719), .B(n8718), .C(n8717), .D(n8716), .Y(n8720) );
  OA22X1 U10100 ( .A0(\i_MIPS/Register/register[0][9] ), .A1(n4702), .B0(
        \i_MIPS/Register/register[8][9] ), .B1(n4700), .Y(n8708) );
  NAND4BX1 U10101 ( .AN(n8821), .B(n8820), .C(n8819), .D(n8818), .Y(n8822) );
  NAND2X1 U10102 ( .A(n10847), .B(ICACHE_addr[28]), .Y(n10848) );
  NOR2X1 U10103 ( .A(n6736), .B(n6735), .Y(n6741) );
  NOR2X1 U10104 ( .A(n6723), .B(n6722), .Y(n6728) );
  NAND2X2 U10105 ( .A(n6104), .B(n6103), .Y(n6105) );
  XOR2X4 U10106 ( .A(n4528), .B(\i_MIPS/n236 ), .Y(n9559) );
  OA22XL U10107 ( .A0(n4908), .A1(n1622), .B0(n4947), .B1(n3199), .Y(n9182) );
  OA22XL U10108 ( .A0(n4912), .A1(n1711), .B0(n4947), .B1(n3308), .Y(n8787) );
  OA22XL U10109 ( .A0(n4917), .A1(n1712), .B0(n4948), .B1(n3309), .Y(n7838) );
  MX2XL U10110 ( .A(n12931), .B(n3914), .S0(n210), .Y(\i_MIPS/n441 ) );
  NAND2BX1 U10111 ( .AN(n9556), .B(\i_MIPS/ID_EX_3 ), .Y(n9558) );
  AOI33X1 U10112 ( .A0(\i_MIPS/Hazard_detection/n7 ), .A1(n9555), .A2(n9554), 
        .B0(\i_MIPS/Hazard_detection/n4 ), .B1(n9553), .B2(n9552), .Y(n9556)
         );
  MX2XL U10113 ( .A(\D_cache/cache[7][137] ), .B(n11025), .S0(n5006), .Y(
        \D_cache/n693 ) );
  MX2XL U10114 ( .A(\D_cache/cache[6][137] ), .B(n11025), .S0(n4962), .Y(
        \D_cache/n694 ) );
  MX2XL U10115 ( .A(\D_cache/cache[5][137] ), .B(n11025), .S0(n4940), .Y(
        \D_cache/n695 ) );
  MX2XL U10116 ( .A(\D_cache/cache[4][137] ), .B(n11025), .S0(n4898), .Y(
        \D_cache/n696 ) );
  MX2XL U10117 ( .A(\D_cache/cache[3][137] ), .B(n11025), .S0(n4852), .Y(
        \D_cache/n697 ) );
  MX2XL U10118 ( .A(\D_cache/cache[2][137] ), .B(n11025), .S0(n4805), .Y(
        \D_cache/n698 ) );
  MX2XL U10119 ( .A(\D_cache/cache[1][137] ), .B(n11025), .S0(n4785), .Y(
        \D_cache/n699 ) );
  MX2XL U10120 ( .A(\D_cache/cache[0][137] ), .B(n11025), .S0(n4732), .Y(
        \D_cache/n700 ) );
  MX2XL U10121 ( .A(\D_cache/cache[7][150] ), .B(n11029), .S0(n5007), .Y(
        \D_cache/n589 ) );
  MX2XL U10122 ( .A(\D_cache/cache[6][150] ), .B(n11029), .S0(n4963), .Y(
        \D_cache/n590 ) );
  MX2XL U10123 ( .A(\D_cache/cache[5][150] ), .B(n11029), .S0(n4944), .Y(
        \D_cache/n591 ) );
  MX2XL U10124 ( .A(\D_cache/cache[4][150] ), .B(n11029), .S0(n4899), .Y(
        \D_cache/n592 ) );
  MX2XL U10125 ( .A(\D_cache/cache[3][150] ), .B(n11029), .S0(n4853), .Y(
        \D_cache/n593 ) );
  MX2XL U10126 ( .A(\D_cache/cache[2][150] ), .B(n11029), .S0(n4808), .Y(
        \D_cache/n594 ) );
  MX2XL U10127 ( .A(\D_cache/cache[1][150] ), .B(n11029), .S0(n4786), .Y(
        \D_cache/n595 ) );
  MX2XL U10128 ( .A(\D_cache/cache[0][150] ), .B(n11029), .S0(n4740), .Y(
        \D_cache/n596 ) );
  MX2XL U10129 ( .A(\D_cache/cache[7][144] ), .B(n11013), .S0(n5006), .Y(
        \D_cache/n637 ) );
  MX2XL U10130 ( .A(\D_cache/cache[6][144] ), .B(n11013), .S0(n4962), .Y(
        \D_cache/n638 ) );
  MX2XL U10131 ( .A(\D_cache/cache[5][144] ), .B(n11013), .S0(n4942), .Y(
        \D_cache/n639 ) );
  MX2XL U10132 ( .A(\D_cache/cache[4][144] ), .B(n11013), .S0(n4898), .Y(
        \D_cache/n640 ) );
  MX2XL U10133 ( .A(\D_cache/cache[3][144] ), .B(n11013), .S0(n4852), .Y(
        \D_cache/n641 ) );
  MX2XL U10134 ( .A(\D_cache/cache[2][144] ), .B(n11013), .S0(n4806), .Y(
        \D_cache/n642 ) );
  MX2XL U10135 ( .A(\D_cache/cache[1][144] ), .B(n11013), .S0(n4784), .Y(
        \D_cache/n643 ) );
  MX2XL U10136 ( .A(\D_cache/cache[0][144] ), .B(n11013), .S0(n4735), .Y(
        \D_cache/n644 ) );
  MX2XL U10137 ( .A(\D_cache/cache[7][140] ), .B(n11010), .S0(n5006), .Y(
        \D_cache/n669 ) );
  MX2XL U10138 ( .A(\D_cache/cache[6][140] ), .B(n11010), .S0(n4962), .Y(
        \D_cache/n670 ) );
  MX2XL U10139 ( .A(\D_cache/cache[5][140] ), .B(n11010), .S0(n4941), .Y(
        \D_cache/n671 ) );
  MX2XL U10140 ( .A(\D_cache/cache[4][140] ), .B(n11010), .S0(n4898), .Y(
        \D_cache/n672 ) );
  MX2XL U10141 ( .A(\D_cache/cache[3][140] ), .B(n11010), .S0(n4852), .Y(
        \D_cache/n673 ) );
  MX2XL U10142 ( .A(\D_cache/cache[2][140] ), .B(n11010), .S0(n4801), .Y(
        \D_cache/n674 ) );
  MX2XL U10143 ( .A(\D_cache/cache[1][140] ), .B(n11010), .S0(n4785), .Y(
        \D_cache/n675 ) );
  MX2XL U10144 ( .A(\D_cache/cache[0][140] ), .B(n11010), .S0(n4738), .Y(
        \D_cache/n676 ) );
  MX2XL U10145 ( .A(\D_cache/cache[1][139] ), .B(n11016), .S0(n4784), .Y(
        \D_cache/n683 ) );
  MX2XL U10146 ( .A(\D_cache/cache[0][139] ), .B(n11016), .S0(n4736), .Y(
        \D_cache/n684 ) );
  OA22XL U10147 ( .A0(\i_MIPS/Register/register[23][27] ), .A1(n9417), .B0(
        \i_MIPS/Register/register[31][27] ), .B1(n9416), .Y(n9418) );
  OA22XL U10148 ( .A0(\i_MIPS/Register/register[7][27] ), .A1(n9417), .B0(
        \i_MIPS/Register/register[15][27] ), .B1(n9416), .Y(n9401) );
  OA22X1 U10149 ( .A0(\i_MIPS/Register/register[23][6] ), .A1(net112152), .B0(
        \i_MIPS/Register/register[31][6] ), .B1(net112164), .Y(n6993) );
  OA22X1 U10150 ( .A0(\i_MIPS/Register/register[23][13] ), .A1(net112148), 
        .B0(\i_MIPS/Register/register[31][13] ), .B1(net112166), .Y(n7727) );
  OA22X1 U10151 ( .A0(\i_MIPS/Register/register[23][10] ), .A1(net112148), 
        .B0(\i_MIPS/Register/register[31][10] ), .B1(net112166), .Y(n7332) );
  OA22X1 U10152 ( .A0(\i_MIPS/Register/register[23][23] ), .A1(net112152), 
        .B0(\i_MIPS/Register/register[31][23] ), .B1(net112170), .Y(n8837) );
  OA22X1 U10153 ( .A0(\i_MIPS/Register/register[23][18] ), .A1(net112152), 
        .B0(\i_MIPS/Register/register[31][18] ), .B1(net112170), .Y(n8774) );
  OA22X1 U10154 ( .A0(\i_MIPS/Register/register[23][20] ), .A1(net112150), 
        .B0(\i_MIPS/Register/register[31][20] ), .B1(net112172), .Y(n9231) );
  OA22X1 U10155 ( .A0(\i_MIPS/Register/register[23][25] ), .A1(net112152), 
        .B0(\i_MIPS/Register/register[31][25] ), .B1(net112170), .Y(n9029) );
  OA22X1 U10156 ( .A0(\i_MIPS/Register/register[23][21] ), .A1(net112150), 
        .B0(\i_MIPS/Register/register[31][21] ), .B1(net112172), .Y(n9126) );
  OA22X1 U10157 ( .A0(\i_MIPS/Register/register[23][24] ), .A1(net112150), 
        .B0(\i_MIPS/Register/register[31][24] ), .B1(net112170), .Y(n8285) );
  OA22XL U10158 ( .A0(n5395), .A1(n1634), .B0(n5331), .B1(n3214), .Y(n6115) );
  OA22X1 U10159 ( .A0(n5400), .A1(n1079), .B0(n5330), .B1(n2657), .Y(n6088) );
  OA22X1 U10160 ( .A0(n5373), .A1(n1273), .B0(n5330), .B1(n2816), .Y(n6084) );
  OA22X1 U10161 ( .A0(n5376), .A1(n1274), .B0(n5330), .B1(n2817), .Y(n6080) );
  OA22X1 U10162 ( .A0(n5395), .A1(n1275), .B0(n5329), .B1(n2818), .Y(n6044) );
  OA22X1 U10163 ( .A0(n5401), .A1(n1276), .B0(n5330), .B1(n2819), .Y(n6076) );
  OA22XL U10164 ( .A0(n5391), .A1(n1623), .B0(n5344), .B1(n3200), .Y(n9925) );
  OA22XL U10165 ( .A0(n5380), .A1(n1624), .B0(n5344), .B1(n3201), .Y(n9934) );
  OA22XL U10166 ( .A0(n5388), .A1(n1625), .B0(n5331), .B1(n3311), .Y(n6123) );
  OA22XL U10167 ( .A0(n5389), .A1(n1626), .B0(n5332), .B1(n3202), .Y(n6157) );
  OA22XL U10168 ( .A0(n5397), .A1(n1627), .B0(n5332), .B1(n3203), .Y(n6162) );
  OA22X1 U10169 ( .A0(n5376), .A1(n1831), .B0(n5342), .B1(n3487), .Y(n9814) );
  OA22X1 U10170 ( .A0(n5399), .A1(n1832), .B0(n5342), .B1(n3488), .Y(n9806) );
  OA22X1 U10171 ( .A0(n5381), .A1(n1833), .B0(n5342), .B1(n3489), .Y(n9818) );
  OA22X1 U10172 ( .A0(n5373), .A1(n1834), .B0(n5342), .B1(n3490), .Y(n9810) );
  OA22X1 U10173 ( .A0(n5372), .A1(n1835), .B0(n5342), .B1(n3491), .Y(n9794) );
  OA22XL U10174 ( .A0(n5400), .A1(n1913), .B0(n5341), .B1(n3568), .Y(n9784) );
  OA22X1 U10175 ( .A0(n5377), .A1(n1836), .B0(n5342), .B1(n3492), .Y(n9798) );
  OA22XL U10176 ( .A0(n5391), .A1(n1914), .B0(n5341), .B1(n3569), .Y(n9789) );
  OA22X1 U10177 ( .A0(n5387), .A1(n1837), .B0(n5343), .B1(n3493), .Y(n9834) );
  OA22X1 U10178 ( .A0(n5399), .A1(n1838), .B0(n5343), .B1(n3494), .Y(n9826) );
  OA22X1 U10179 ( .A0(n5379), .A1(n1839), .B0(n5343), .B1(n3495), .Y(n9838) );
  OA22X1 U10180 ( .A0(n269), .A1(n1840), .B0(n5343), .B1(n3496), .Y(n9830) );
  OA22X1 U10181 ( .A0(n5385), .A1(n1841), .B0(n5342), .B1(n3497), .Y(n9870) );
  OA22X1 U10182 ( .A0(n5398), .A1(n3590), .B0(n5343), .B1(n1915), .Y(n9862) );
  OA22X1 U10183 ( .A0(n5389), .A1(n1842), .B0(n5342), .B1(n3498), .Y(n9874) );
  OA22X1 U10184 ( .A0(n5397), .A1(n1843), .B0(n5342), .B1(n3499), .Y(n9866) );
  OA22X1 U10185 ( .A0(n5386), .A1(n1844), .B0(n5343), .B1(n3500), .Y(n9854) );
  OA22X1 U10186 ( .A0(n5394), .A1(n1845), .B0(n5343), .B1(n3501), .Y(n9846) );
  OA22X1 U10187 ( .A0(n5398), .A1(n1846), .B0(n5343), .B1(n3502), .Y(n9858) );
  OA22X1 U10188 ( .A0(n5384), .A1(n1847), .B0(n5343), .B1(n3503), .Y(n9850) );
  OA22XL U10189 ( .A0(n5371), .A1(n1916), .B0(n5338), .B1(n3570), .Y(n9625) );
  OA22XL U10190 ( .A0(n5383), .A1(n1917), .B0(n5338), .B1(n3571), .Y(n9615) );
  OA22XL U10191 ( .A0(n5378), .A1(n1918), .B0(n5338), .B1(n3572), .Y(n9630) );
  OA22XL U10192 ( .A0(n5370), .A1(n1919), .B0(n5338), .B1(n3573), .Y(n9620) );
  OA22XL U10193 ( .A0(n5367), .A1(n1920), .B0(n5337), .B1(n3574), .Y(n9579) );
  OA22XL U10194 ( .A0(n5375), .A1(n1921), .B0(n5337), .B1(n3575), .Y(n9583) );
  OA22XL U10195 ( .A0(n5390), .A1(n1922), .B0(n5343), .B1(n3576), .Y(n9674) );
  OA22XL U10196 ( .A0(n5401), .A1(n1923), .B0(n5343), .B1(n3577), .Y(n9664) );
  OA22XL U10197 ( .A0(n5369), .A1(n1924), .B0(n5342), .B1(n3578), .Y(n9679) );
  OA22XL U10198 ( .A0(n5397), .A1(n1925), .B0(n5342), .B1(n3579), .Y(n9669) );
  OA22XL U10199 ( .A0(n5382), .A1(n1926), .B0(n5347), .B1(n3580), .Y(n10163)
         );
  OA22XL U10200 ( .A0(n237), .A1(n1927), .B0(n5347), .B1(n3581), .Y(n10153) );
  OA22XL U10201 ( .A0(n5388), .A1(n1928), .B0(n5348), .B1(n3582), .Y(n10168)
         );
  OA22XL U10202 ( .A0(n5374), .A1(n1929), .B0(n5347), .B1(n3583), .Y(n10158)
         );
  OA22XL U10203 ( .A0(n5395), .A1(n1930), .B0(n5340), .B1(n3584), .Y(n9723) );
  OA22XL U10204 ( .A0(n5393), .A1(n1931), .B0(n5339), .B1(n3585), .Y(n9713) );
  OA22XL U10205 ( .A0(n5380), .A1(n1932), .B0(n5340), .B1(n3586), .Y(n9728) );
  OA22XL U10206 ( .A0(n5368), .A1(n1933), .B0(n5339), .B1(n3587), .Y(n9718) );
  OA22XL U10207 ( .A0(\i_MIPS/Register/register[19][27] ), .A1(n9415), .B0(
        \i_MIPS/Register/register[27][27] ), .B1(n9414), .Y(n9419) );
  OA22XL U10208 ( .A0(\i_MIPS/Register/register[3][27] ), .A1(n9415), .B0(
        \i_MIPS/Register/register[11][27] ), .B1(n9414), .Y(n9402) );
  OA22XL U10209 ( .A0(\i_MIPS/Register/register[0][19] ), .A1(net102048), .B0(
        \i_MIPS/Register/register[8][19] ), .B1(net102049), .Y(n8573) );
  OA22XL U10210 ( .A0(\i_MIPS/Register/register[16][30] ), .A1(net102048), 
        .B0(\i_MIPS/Register/register[24][30] ), .B1(net102049), .Y(n6474) );
  OA22XL U10211 ( .A0(\i_MIPS/Register/register[0][30] ), .A1(net102048), .B0(
        \i_MIPS/Register/register[8][30] ), .B1(net102049), .Y(n6465) );
  MX2XL U10212 ( .A(\D_cache/cache[6][146] ), .B(n11033), .S0(n4963), .Y(
        \D_cache/n622 ) );
  MX2XL U10213 ( .A(\D_cache/cache[5][146] ), .B(n11033), .S0(n4944), .Y(
        \D_cache/n623 ) );
  MX2XL U10214 ( .A(\D_cache/cache[4][146] ), .B(n11033), .S0(n4899), .Y(
        \D_cache/n624 ) );
  MX2XL U10215 ( .A(\D_cache/cache[3][146] ), .B(n11033), .S0(n4853), .Y(
        \D_cache/n625 ) );
  MX2XL U10216 ( .A(\D_cache/cache[2][146] ), .B(n11033), .S0(n4808), .Y(
        \D_cache/n626 ) );
  MX2XL U10217 ( .A(\D_cache/cache[1][146] ), .B(n11033), .S0(n4783), .Y(
        \D_cache/n627 ) );
  MX2XL U10218 ( .A(\D_cache/cache[0][146] ), .B(n11033), .S0(n4740), .Y(
        \D_cache/n628 ) );
  MX2XL U10219 ( .A(\D_cache/cache[6][135] ), .B(n11024), .S0(n4962), .Y(
        \D_cache/n710 ) );
  MX2XL U10220 ( .A(\D_cache/cache[5][135] ), .B(n11024), .S0(n4942), .Y(
        \D_cache/n711 ) );
  MX2XL U10221 ( .A(\D_cache/cache[4][135] ), .B(n11024), .S0(n4898), .Y(
        \D_cache/n712 ) );
  MX2XL U10222 ( .A(\D_cache/cache[3][135] ), .B(n11024), .S0(n4852), .Y(
        \D_cache/n713 ) );
  MX2XL U10223 ( .A(\D_cache/cache[2][135] ), .B(n11024), .S0(n4802), .Y(
        \D_cache/n714 ) );
  MX2XL U10224 ( .A(\D_cache/cache[1][135] ), .B(n11024), .S0(n4785), .Y(
        \D_cache/n715 ) );
  MX2XL U10225 ( .A(\D_cache/cache[0][135] ), .B(n11024), .S0(n4732), .Y(
        \D_cache/n716 ) );
  OA22X1 U10226 ( .A0(\i_MIPS/Register/register[19][6] ), .A1(net112182), .B0(
        \i_MIPS/Register/register[27][6] ), .B1(n198), .Y(n6994) );
  OA22X1 U10227 ( .A0(\i_MIPS/Register/register[3][6] ), .A1(net112182), .B0(
        \i_MIPS/Register/register[11][6] ), .B1(n199), .Y(n6985) );
  OA22X1 U10228 ( .A0(\i_MIPS/Register/register[19][10] ), .A1(net112188), 
        .B0(\i_MIPS/Register/register[27][10] ), .B1(n200), .Y(n7333) );
  OA22X1 U10229 ( .A0(\i_MIPS/Register/register[3][10] ), .A1(net112188), .B0(
        \i_MIPS/Register/register[11][10] ), .B1(n200), .Y(n7324) );
  OA22X1 U10230 ( .A0(\i_MIPS/Register/register[19][18] ), .A1(net112188), 
        .B0(\i_MIPS/Register/register[27][18] ), .B1(n200), .Y(n8775) );
  OA22X1 U10231 ( .A0(\i_MIPS/Register/register[3][18] ), .A1(net112188), .B0(
        \i_MIPS/Register/register[11][18] ), .B1(n199), .Y(n8766) );
  OA22X1 U10232 ( .A0(\i_MIPS/Register/register[19][24] ), .A1(net112182), 
        .B0(\i_MIPS/Register/register[27][24] ), .B1(n197), .Y(n8286) );
  OA22X1 U10233 ( .A0(\i_MIPS/Register/register[3][24] ), .A1(net112188), .B0(
        \i_MIPS/Register/register[11][24] ), .B1(n199), .Y(n8277) );
  OA22X2 U10234 ( .A0(n4910), .A1(n1452), .B0(n4947), .B1(n3022), .Y(n8984) );
  OA22X2 U10235 ( .A0(n4917), .A1(n1454), .B0(n4948), .B1(n3025), .Y(n7842) );
  OA22XL U10236 ( .A0(n4905), .A1(n1628), .B0(n4947), .B1(n3204), .Y(n6300) );
  OA22XL U10237 ( .A0(n4915), .A1(n1715), .B0(n4947), .B1(n3313), .Y(n9189) );
  OA22XL U10238 ( .A0(n4909), .A1(n3270), .B0(n4947), .B1(n1635), .Y(n9289) );
  OA22XL U10239 ( .A0(n4910), .A1(n1716), .B0(n4947), .B1(n3314), .Y(n9511) );
  OA22XL U10240 ( .A0(n4912), .A1(n1457), .B0(n4950), .B1(n3027), .Y(n6654) );
  OA22XL U10241 ( .A0(n4923), .A1(n1717), .B0(n4950), .B1(n3315), .Y(n6808) );
  OA22XL U10242 ( .A0(n4907), .A1(n1629), .B0(n4947), .B1(n3205), .Y(n9508) );
  OA22XL U10243 ( .A0(n4906), .A1(n1718), .B0(n4947), .B1(n3316), .Y(n9501) );
  OA22XL U10244 ( .A0(n4923), .A1(n1719), .B0(n4950), .B1(n3317), .Y(n6800) );
  OA22XL U10245 ( .A0(n4912), .A1(n1630), .B0(n4950), .B1(n3206), .Y(n6646) );
  OA22XL U10246 ( .A0(n4907), .A1(n1720), .B0(n4950), .B1(n3318), .Y(n6650) );
  OA22XL U10247 ( .A0(n4912), .A1(n1631), .B0(n4950), .B1(n3207), .Y(n6642) );
  OA22XL U10248 ( .A0(n4927), .A1(n1632), .B0(n4950), .B1(n3208), .Y(n6318) );
  AO22X1 U10249 ( .A0(n4729), .A1(n375), .B0(n4727), .B1(n1029), .Y(n9314) );
  AO22X1 U10250 ( .A0(n4729), .A1(n376), .B0(n4727), .B1(n1030), .Y(n9305) );
  AO22X1 U10251 ( .A0(n4730), .A1(n854), .B0(n4725), .B1(n2422), .Y(n8120) );
  AO22X1 U10252 ( .A0(n4731), .A1(n377), .B0(n4724), .B1(n2478), .Y(n7673) );
  AO22X1 U10253 ( .A0(n4728), .A1(n962), .B0(n4725), .B1(n2479), .Y(n7767) );
  AO22X1 U10254 ( .A0(n4728), .A1(n855), .B0(n4725), .B1(n2423), .Y(n8111) );
  AO22X1 U10255 ( .A0(n4731), .A1(n378), .B0(n4724), .B1(n2480), .Y(n7664) );
  AO22X1 U10256 ( .A0(n4730), .A1(n963), .B0(n4726), .B1(n2481), .Y(n6952) );
  AO22X1 U10257 ( .A0(n4730), .A1(n964), .B0(n4726), .B1(n2482), .Y(n7032) );
  AO22X1 U10258 ( .A0(n4730), .A1(n965), .B0(n4726), .B1(n2483), .Y(n6943) );
  AO22X1 U10259 ( .A0(n4730), .A1(n966), .B0(n4726), .B1(n2484), .Y(n7023) );
  AO22X1 U10260 ( .A0(net112002), .A1(n856), .B0(net112020), .B1(n2424), .Y(
        n7328) );
  AO22X1 U10261 ( .A0(net112006), .A1(n857), .B0(net112020), .B1(n2425), .Y(
        n8779) );
  AO22X1 U10262 ( .A0(net112006), .A1(n858), .B0(net112020), .B1(n2426), .Y(
        n8770) );
  AO22X1 U10263 ( .A0(net112008), .A1(n967), .B0(net112026), .B1(n2485), .Y(
        n9227) );
  AO22X1 U10264 ( .A0(net112004), .A1(n379), .B0(net112030), .B1(n1031), .Y(
        n8135) );
  AO22X1 U10265 ( .A0(net112004), .A1(n400), .B0(net112030), .B1(n1049), .Y(
        n8144) );
  OA22X1 U10266 ( .A0(n5303), .A1(n3216), .B0(n5258), .B1(n1419), .Y(n10089)
         );
  OA22XL U10267 ( .A0(n5303), .A1(n1633), .B0(n5258), .B1(n3319), .Y(n10056)
         );
  OA22X1 U10268 ( .A0(n5297), .A1(n1567), .B0(n5250), .B1(n3213), .Y(n9739) );
  OA22X1 U10269 ( .A0(n5293), .A1(n1568), .B0(n5246), .B1(n3150), .Y(n9592) );
  OA22X1 U10270 ( .A0(n5298), .A1(n1569), .B0(n5251), .B1(n3151), .Y(n9762) );
  OA22X1 U10271 ( .A0(n5292), .A1(n1570), .B0(n5245), .B1(n3152), .Y(n6269) );
  OA22X1 U10272 ( .A0(n5292), .A1(n1571), .B0(n5245), .B1(n3153), .Y(n6261) );
  OA22X1 U10273 ( .A0(n5292), .A1(n1572), .B0(n5245), .B1(n3154), .Y(n6273) );
  OA22X1 U10274 ( .A0(n5292), .A1(n1573), .B0(n5245), .B1(n3155), .Y(n6265) );
  OA22XL U10275 ( .A0(\i_MIPS/Register/register[21][27] ), .A1(n188), .B0(
        \i_MIPS/Register/register[29][27] ), .B1(n9412), .Y(n9420) );
  OA22XL U10276 ( .A0(\i_MIPS/Register/register[5][27] ), .A1(n186), .B0(
        \i_MIPS/Register/register[13][27] ), .B1(n9412), .Y(n9403) );
  OAI221XL U10277 ( .A0(\i_MIPS/ALUin1[24] ), .A1(net112364), .B0(
        \i_MIPS/ALUin1[25] ), .B1(net112346), .C0(n6681), .Y(n9335) );
  OA22XL U10278 ( .A0(\i_MIPS/Register/register[4][19] ), .A1(net102050), .B0(
        \i_MIPS/Register/register[12][19] ), .B1(net102051), .Y(n8574) );
  OA22XL U10279 ( .A0(\i_MIPS/Register/register[20][30] ), .A1(net102050), 
        .B0(\i_MIPS/Register/register[28][30] ), .B1(net102051), .Y(n6475) );
  OA22XL U10280 ( .A0(\i_MIPS/Register/register[4][30] ), .A1(net102050), .B0(
        \i_MIPS/Register/register[12][30] ), .B1(net102051), .Y(n6466) );
  OA22X1 U10281 ( .A0(\i_MIPS/Register/register[22][6] ), .A1(net112110), .B0(
        \i_MIPS/Register/register[30][6] ), .B1(net112128), .Y(n6997) );
  OA22X1 U10282 ( .A0(\i_MIPS/Register/register[22][18] ), .A1(net112116), 
        .B0(\i_MIPS/Register/register[30][18] ), .B1(net112134), .Y(n8778) );
  OA22X1 U10283 ( .A0(\i_MIPS/Register/register[22][20] ), .A1(net112112), 
        .B0(\i_MIPS/Register/register[30][20] ), .B1(net112142), .Y(n9235) );
  OA22X1 U10284 ( .A0(\i_MIPS/Register/register[22][26] ), .A1(n4684), .B0(
        \i_MIPS/Register/register[30][26] ), .B1(n4678), .Y(n9006) );
  OA22X1 U10285 ( .A0(\i_MIPS/Register/register[6][26] ), .A1(n4684), .B0(
        \i_MIPS/Register/register[14][26] ), .B1(n4678), .Y(n8997) );
  OA22X1 U10286 ( .A0(\i_MIPS/Register/register[6][6] ), .A1(n4684), .B0(
        \i_MIPS/Register/register[14][6] ), .B1(n4680), .Y(n7022) );
  OA22X1 U10287 ( .A0(\i_MIPS/Register/register[22][22] ), .A1(n4682), .B0(
        \i_MIPS/Register/register[30][22] ), .B1(n4679), .Y(n9526) );
  OAI221XL U10288 ( .A0(\i_MIPS/Register/register[18][27] ), .A1(n4690), .B0(
        \i_MIPS/Register/register[26][27] ), .B1(n4686), .C0(n9422), .Y(n9425)
         );
  MX2XL U10289 ( .A(n12941), .B(n10502), .S0(n211), .Y(\i_MIPS/n451 ) );
  OA22XL U10290 ( .A0(\i_MIPS/Register/register[17][27] ), .A1(n9411), .B0(
        \i_MIPS/Register/register[25][27] ), .B1(n9410), .Y(n9421) );
  OA22XL U10291 ( .A0(\i_MIPS/Register/register[1][27] ), .A1(n9411), .B0(
        \i_MIPS/Register/register[9][27] ), .B1(n9410), .Y(n9404) );
  OA22X1 U10292 ( .A0(\i_MIPS/Register/register[4][19] ), .A1(n4698), .B0(
        \i_MIPS/Register/register[12][19] ), .B1(n4694), .Y(n8614) );
  OA22X1 U10293 ( .A0(\i_MIPS/Register/register[21][6] ), .A1(n192), .B0(
        \i_MIPS/Register/register[29][6] ), .B1(net112236), .Y(n6995) );
  OA22X1 U10294 ( .A0(\i_MIPS/Register/register[21][4] ), .A1(n192), .B0(
        \i_MIPS/Register/register[29][4] ), .B1(net112242), .Y(n6870) );
  OA22X1 U10295 ( .A0(\i_MIPS/Register/register[21][13] ), .A1(net112222), 
        .B0(\i_MIPS/Register/register[29][13] ), .B1(net112236), .Y(n7729) );
  OA22X1 U10296 ( .A0(\i_MIPS/Register/register[21][14] ), .A1(net112222), 
        .B0(\i_MIPS/Register/register[29][14] ), .B1(net112242), .Y(n7636) );
  OA22X1 U10297 ( .A0(\i_MIPS/Register/register[21][11] ), .A1(net112222), 
        .B0(\i_MIPS/Register/register[29][11] ), .B1(net112236), .Y(n7255) );
  OA22X1 U10298 ( .A0(\i_MIPS/Register/register[21][10] ), .A1(net112222), 
        .B0(\i_MIPS/Register/register[29][10] ), .B1(net112236), .Y(n7334) );
  OA22X1 U10299 ( .A0(\i_MIPS/Register/register[21][9] ), .A1(net112224), .B0(
        \i_MIPS/Register/register[29][9] ), .B1(net112236), .Y(n8674) );
  OA22X1 U10300 ( .A0(\i_MIPS/Register/register[21][23] ), .A1(net112224), 
        .B0(\i_MIPS/Register/register[29][23] ), .B1(net112242), .Y(n8839) );
  OA22X1 U10301 ( .A0(\i_MIPS/Register/register[21][18] ), .A1(net112224), 
        .B0(\i_MIPS/Register/register[29][18] ), .B1(net112244), .Y(n8776) );
  OA22X1 U10302 ( .A0(\i_MIPS/Register/register[21][25] ), .A1(net112224), 
        .B0(\i_MIPS/Register/register[29][25] ), .B1(net112236), .Y(n9031) );
  OA22X1 U10303 ( .A0(\i_MIPS/Register/register[21][24] ), .A1(net112222), 
        .B0(\i_MIPS/Register/register[29][24] ), .B1(net112236), .Y(n8287) );
  AO22X1 U10304 ( .A0(net112038), .A1(n380), .B0(net100603), .B1(n1032), .Y(
        n7386) );
  AO22X1 U10305 ( .A0(net112050), .A1(n1019), .B0(net100603), .B1(n2545), .Y(
        n9439) );
  AO22X1 U10306 ( .A0(net112036), .A1(n968), .B0(net100603), .B1(n2486), .Y(
        n6784) );
  AO22X1 U10307 ( .A0(net112036), .A1(n859), .B0(net100603), .B1(n2427), .Y(
        n7783) );
  AO22X1 U10308 ( .A0(net112038), .A1(n334), .B0(net100603), .B1(n978), .Y(
        n7329) );
  AO22X1 U10309 ( .A0(net112038), .A1(n860), .B0(net100603), .B1(n2428), .Y(
        n8771) );
  AO22X1 U10310 ( .A0(net112036), .A1(n969), .B0(net100603), .B1(n2487), .Y(
        n7995) );
  AO22X1 U10311 ( .A0(net112036), .A1(n970), .B0(net100603), .B1(n2488), .Y(
        n7724) );
  AO22X1 U10312 ( .A0(net112050), .A1(n971), .B0(net100603), .B1(n2489), .Y(
        n9228) );
  AO22X1 U10313 ( .A0(net112038), .A1(n381), .B0(net100603), .B1(n1033), .Y(
        n7631) );
  AO22X1 U10314 ( .A0(net112036), .A1(n972), .B0(net100603), .B1(n2490), .Y(
        n6990) );
  AO22X1 U10315 ( .A0(net112036), .A1(n973), .B0(net100603), .B1(n2491), .Y(
        n8053) );
  AO22X1 U10316 ( .A0(net112050), .A1(n1020), .B0(net100603), .B1(n2546), .Y(
        n9123) );
  AO22X1 U10317 ( .A0(net112038), .A1(n861), .B0(net100603), .B1(n2429), .Y(
        n8834) );
  AO22X1 U10318 ( .A0(net112038), .A1(n974), .B0(net100603), .B1(n2492), .Y(
        n8471) );
  AO22X1 U10319 ( .A0(net112038), .A1(n862), .B0(net100603), .B1(n2430), .Y(
        n8669) );
  AO22X1 U10320 ( .A0(net112038), .A1(n975), .B0(net100603), .B1(n2493), .Y(
        n8373) );
  AO22X1 U10321 ( .A0(net112036), .A1(n863), .B0(net100603), .B1(n2431), .Y(
        n7916) );
  AO22X1 U10322 ( .A0(net112038), .A1(n335), .B0(net100603), .B1(n979), .Y(
        n7558) );
  AO22X1 U10323 ( .A0(net112050), .A1(n864), .B0(net100603), .B1(n2432), .Y(
        n9026) );
  AO22X1 U10324 ( .A0(net112036), .A1(n865), .B0(net100603), .B1(n2433), .Y(
        n6865) );
  AO22X1 U10325 ( .A0(net112038), .A1(n401), .B0(net100603), .B1(n1050), .Y(
        n7133) );
  AO22X1 U10326 ( .A0(net112050), .A1(n976), .B0(net100603), .B1(n2494), .Y(
        n8925) );
  AO22X1 U10327 ( .A0(net112038), .A1(n977), .B0(net100603), .B1(n2495), .Y(
        n8282) );
  AO22X1 U10328 ( .A0(net112036), .A1(n1021), .B0(net100603), .B1(n2547), .Y(
        n7074) );
  AO22X1 U10329 ( .A0(net112038), .A1(n336), .B0(net100603), .B1(n980), .Y(
        n7250) );
  AO22X1 U10330 ( .A0(net112036), .A1(n435), .B0(net100603), .B1(n2015), .Y(
        n6665) );
  MX2XL U10331 ( .A(\D_cache/cache[6][115] ), .B(n11001), .S0(n4964), .Y(
        \D_cache/n870 ) );
  MX2XL U10332 ( .A(\D_cache/cache[5][115] ), .B(n11001), .S0(n4943), .Y(
        \D_cache/n871 ) );
  MX2XL U10333 ( .A(\D_cache/cache[4][115] ), .B(n11001), .S0(n4900), .Y(
        \D_cache/n872 ) );
  MX2XL U10334 ( .A(\D_cache/cache[3][115] ), .B(n11001), .S0(n4854), .Y(
        \D_cache/n873 ) );
  MX2XL U10335 ( .A(\D_cache/cache[2][115] ), .B(n11001), .S0(n4809), .Y(
        \D_cache/n874 ) );
  MX2XL U10336 ( .A(\D_cache/cache[1][115] ), .B(n11001), .S0(n4786), .Y(
        \D_cache/n875 ) );
  MX2XL U10337 ( .A(\D_cache/cache[0][115] ), .B(n11001), .S0(n4741), .Y(
        \D_cache/n876 ) );
  MX2XL U10338 ( .A(\D_cache/cache[5][61] ), .B(n10686), .S0(n4937), .Y(
        \D_cache/n1303 ) );
  MX2XL U10339 ( .A(\D_cache/cache[4][61] ), .B(n10686), .S0(n4893), .Y(
        \D_cache/n1304 ) );
  MX2XL U10340 ( .A(\D_cache/cache[3][61] ), .B(n10686), .S0(n4847), .Y(
        \D_cache/n1305 ) );
  MX2XL U10341 ( .A(\D_cache/cache[2][61] ), .B(n10686), .S0(n4802), .Y(
        \D_cache/n1306 ) );
  MX2XL U10342 ( .A(\D_cache/cache[1][61] ), .B(n10686), .S0(n4779), .Y(
        \D_cache/n1307 ) );
  MX2XL U10343 ( .A(\D_cache/cache[0][61] ), .B(n10686), .S0(n4738), .Y(
        \D_cache/n1308 ) );
  MX2XL U10344 ( .A(\D_cache/cache[6][60] ), .B(n10480), .S0(n4956), .Y(
        \D_cache/n1310 ) );
  MX2XL U10345 ( .A(\D_cache/cache[5][60] ), .B(n10480), .S0(n4937), .Y(
        \D_cache/n1311 ) );
  MX2XL U10346 ( .A(\D_cache/cache[4][60] ), .B(n10480), .S0(n4892), .Y(
        \D_cache/n1312 ) );
  MX2XL U10347 ( .A(\D_cache/cache[3][60] ), .B(n10480), .S0(n4846), .Y(
        \D_cache/n1313 ) );
  MX2XL U10348 ( .A(\D_cache/cache[2][60] ), .B(n10480), .S0(n4801), .Y(
        \D_cache/n1314 ) );
  MX2XL U10349 ( .A(\D_cache/cache[1][60] ), .B(n10480), .S0(n4778), .Y(
        \D_cache/n1315 ) );
  MX2XL U10350 ( .A(\D_cache/cache[0][60] ), .B(n10480), .S0(n4732), .Y(
        \D_cache/n1316 ) );
  MX2XL U10351 ( .A(\D_cache/cache[6][56] ), .B(n10781), .S0(n4959), .Y(
        \D_cache/n1342 ) );
  MX2XL U10352 ( .A(\D_cache/cache[5][56] ), .B(n10781), .S0(n4939), .Y(
        \D_cache/n1343 ) );
  MX2XL U10353 ( .A(\D_cache/cache[4][56] ), .B(n10781), .S0(n4894), .Y(
        \D_cache/n1344 ) );
  MX2XL U10354 ( .A(\D_cache/cache[3][56] ), .B(n10781), .S0(n4849), .Y(
        \D_cache/n1345 ) );
  MX2XL U10355 ( .A(\D_cache/cache[2][56] ), .B(n10781), .S0(n4805), .Y(
        \D_cache/n1346 ) );
  MX2XL U10356 ( .A(\D_cache/cache[1][56] ), .B(n10781), .S0(n4782), .Y(
        \D_cache/n1347 ) );
  MX2XL U10357 ( .A(\D_cache/cache[0][56] ), .B(n10781), .S0(n4736), .Y(
        \D_cache/n1348 ) );
  MX2XL U10358 ( .A(\D_cache/cache[6][54] ), .B(n10214), .S0(n4957), .Y(
        \D_cache/n1358 ) );
  MX2XL U10359 ( .A(\D_cache/cache[5][54] ), .B(n10214), .S0(n4937), .Y(
        \D_cache/n1359 ) );
  MX2XL U10360 ( .A(\D_cache/cache[4][54] ), .B(n10214), .S0(n4894), .Y(
        \D_cache/n1360 ) );
  MX2XL U10361 ( .A(\D_cache/cache[3][54] ), .B(n10214), .S0(n4846), .Y(
        \D_cache/n1361 ) );
  MX2XL U10362 ( .A(\D_cache/cache[2][54] ), .B(n10214), .S0(n4803), .Y(
        \D_cache/n1362 ) );
  MX2XL U10363 ( .A(\D_cache/cache[1][54] ), .B(n10214), .S0(n4780), .Y(
        \D_cache/n1363 ) );
  MX2XL U10364 ( .A(\D_cache/cache[0][54] ), .B(n10214), .S0(n4734), .Y(
        \D_cache/n1364 ) );
  MX2XL U10365 ( .A(\D_cache/cache[6][53] ), .B(n10672), .S0(n4957), .Y(
        \D_cache/n1366 ) );
  MX2XL U10366 ( .A(\D_cache/cache[5][53] ), .B(n10672), .S0(n4937), .Y(
        \D_cache/n1367 ) );
  MX2XL U10367 ( .A(\D_cache/cache[4][53] ), .B(n10672), .S0(n4893), .Y(
        \D_cache/n1368 ) );
  MX2XL U10368 ( .A(\D_cache/cache[3][53] ), .B(n10672), .S0(n4847), .Y(
        \D_cache/n1369 ) );
  MX2XL U10369 ( .A(\D_cache/cache[2][53] ), .B(n10672), .S0(n4802), .Y(
        \D_cache/n1370 ) );
  MX2XL U10370 ( .A(\D_cache/cache[1][53] ), .B(n10672), .S0(n4779), .Y(
        \D_cache/n1371 ) );
  MX2XL U10371 ( .A(\D_cache/cache[0][53] ), .B(n10672), .S0(n4733), .Y(
        \D_cache/n1372 ) );
  MX2XL U10372 ( .A(\D_cache/cache[6][52] ), .B(n10659), .S0(n4957), .Y(
        \D_cache/n1374 ) );
  MX2XL U10373 ( .A(\D_cache/cache[5][52] ), .B(n10659), .S0(n4937), .Y(
        \D_cache/n1375 ) );
  MX2XL U10374 ( .A(\D_cache/cache[4][52] ), .B(n10659), .S0(n4893), .Y(
        \D_cache/n1376 ) );
  MX2XL U10375 ( .A(\D_cache/cache[3][52] ), .B(n10659), .S0(n4847), .Y(
        \D_cache/n1377 ) );
  MX2XL U10376 ( .A(\D_cache/cache[2][52] ), .B(n10659), .S0(n4802), .Y(
        \D_cache/n1378 ) );
  MX2XL U10377 ( .A(\D_cache/cache[1][52] ), .B(n10659), .S0(n4779), .Y(
        \D_cache/n1379 ) );
  MX2XL U10378 ( .A(\D_cache/cache[0][52] ), .B(n10659), .S0(n4733), .Y(
        \D_cache/n1380 ) );
  MX2XL U10379 ( .A(\D_cache/cache[0][49] ), .B(n10768), .S0(n4736), .Y(
        \D_cache/n1404 ) );
  MX2XL U10380 ( .A(\D_cache/cache[6][47] ), .B(n10757), .S0(n4961), .Y(
        \D_cache/n1414 ) );
  MX2XL U10381 ( .A(\D_cache/cache[5][47] ), .B(n10757), .S0(n4941), .Y(
        \D_cache/n1415 ) );
  MX2XL U10382 ( .A(\D_cache/cache[4][47] ), .B(n10757), .S0(n4897), .Y(
        \D_cache/n1416 ) );
  MX2XL U10383 ( .A(\D_cache/cache[3][47] ), .B(n10757), .S0(n4851), .Y(
        \D_cache/n1417 ) );
  MX2XL U10384 ( .A(\D_cache/cache[2][47] ), .B(n10757), .S0(n4807), .Y(
        \D_cache/n1418 ) );
  MX2XL U10385 ( .A(\D_cache/cache[1][47] ), .B(n10757), .S0(n4784), .Y(
        \D_cache/n1419 ) );
  MX2XL U10386 ( .A(\D_cache/cache[6][43] ), .B(n10712), .S0(n4960), .Y(
        \D_cache/n1446 ) );
  MX2XL U10387 ( .A(\D_cache/cache[5][43] ), .B(n10712), .S0(n4942), .Y(
        \D_cache/n1447 ) );
  MX2XL U10388 ( .A(\D_cache/cache[4][43] ), .B(n10712), .S0(n4896), .Y(
        \D_cache/n1448 ) );
  MX2XL U10389 ( .A(\D_cache/cache[3][43] ), .B(n10712), .S0(n4850), .Y(
        \D_cache/n1449 ) );
  MX2XL U10390 ( .A(\D_cache/cache[2][43] ), .B(n10712), .S0(n4806), .Y(
        \D_cache/n1450 ) );
  MX2XL U10391 ( .A(\D_cache/cache[1][43] ), .B(n10712), .S0(n4780), .Y(
        \D_cache/n1451 ) );
  MX2XL U10392 ( .A(\D_cache/cache[0][43] ), .B(n10712), .S0(n4738), .Y(
        \D_cache/n1452 ) );
  MX2XL U10393 ( .A(\D_cache/cache[6][42] ), .B(n10262), .S0(n4958), .Y(
        \D_cache/n1454 ) );
  MX2XL U10394 ( .A(\D_cache/cache[5][42] ), .B(n10262), .S0(n4939), .Y(
        \D_cache/n1455 ) );
  MX2XL U10395 ( .A(\D_cache/cache[4][42] ), .B(n10262), .S0(n4895), .Y(
        \D_cache/n1456 ) );
  MX2XL U10396 ( .A(\D_cache/cache[3][42] ), .B(n10262), .S0(n4848), .Y(
        \D_cache/n1457 ) );
  MX2XL U10397 ( .A(\D_cache/cache[2][42] ), .B(n10262), .S0(n4804), .Y(
        \D_cache/n1458 ) );
  MX2XL U10398 ( .A(\D_cache/cache[1][42] ), .B(n10262), .S0(n4782), .Y(
        \D_cache/n1459 ) );
  MX2XL U10399 ( .A(\D_cache/cache[0][42] ), .B(n10262), .S0(n4735), .Y(
        \D_cache/n1460 ) );
  MX2XL U10400 ( .A(\D_cache/cache[6][41] ), .B(n10700), .S0(n4960), .Y(
        \D_cache/n1462 ) );
  MX2XL U10401 ( .A(\D_cache/cache[5][41] ), .B(n10700), .S0(n4938), .Y(
        \D_cache/n1463 ) );
  MX2XL U10402 ( .A(\D_cache/cache[4][41] ), .B(n10700), .S0(n4896), .Y(
        \D_cache/n1464 ) );
  MX2XL U10403 ( .A(\D_cache/cache[3][41] ), .B(n10700), .S0(n4850), .Y(
        \D_cache/n1465 ) );
  MX2XL U10404 ( .A(\D_cache/cache[2][41] ), .B(n10700), .S0(n4806), .Y(
        \D_cache/n1466 ) );
  MX2XL U10405 ( .A(\D_cache/cache[1][41] ), .B(n10700), .S0(n4780), .Y(
        \D_cache/n1467 ) );
  MX2XL U10406 ( .A(\D_cache/cache[0][41] ), .B(n10700), .S0(n4738), .Y(
        \D_cache/n1468 ) );
  MX2XL U10407 ( .A(\D_cache/cache[6][40] ), .B(n10898), .S0(n4958), .Y(
        \D_cache/n1470 ) );
  MX2XL U10408 ( .A(\D_cache/cache[5][40] ), .B(n10898), .S0(n4940), .Y(
        \D_cache/n1471 ) );
  MX2XL U10409 ( .A(\D_cache/cache[4][40] ), .B(n10898), .S0(n4893), .Y(
        \D_cache/n1472 ) );
  MX2XL U10410 ( .A(\D_cache/cache[3][40] ), .B(n10898), .S0(n4849), .Y(
        \D_cache/n1473 ) );
  MX2XL U10411 ( .A(\D_cache/cache[2][40] ), .B(n10898), .S0(n4801), .Y(
        \D_cache/n1474 ) );
  MX2XL U10412 ( .A(\D_cache/cache[1][40] ), .B(n10898), .S0(n4781), .Y(
        \D_cache/n1475 ) );
  MX2XL U10413 ( .A(\D_cache/cache[0][40] ), .B(n10898), .S0(n4737), .Y(
        \D_cache/n1476 ) );
  MX2XL U10414 ( .A(\D_cache/cache[6][39] ), .B(n10886), .S0(n4956), .Y(
        \D_cache/n1478 ) );
  MX2XL U10415 ( .A(\D_cache/cache[5][39] ), .B(n10886), .S0(n4938), .Y(
        \D_cache/n1479 ) );
  MX2XL U10416 ( .A(\D_cache/cache[4][39] ), .B(n10886), .S0(n4894), .Y(
        \D_cache/n1480 ) );
  MX2XL U10417 ( .A(\D_cache/cache[3][39] ), .B(n10886), .S0(n4848), .Y(
        \D_cache/n1481 ) );
  MX2XL U10418 ( .A(\D_cache/cache[2][39] ), .B(n10886), .S0(n4802), .Y(
        \D_cache/n1482 ) );
  MX2XL U10419 ( .A(\D_cache/cache[1][39] ), .B(n10886), .S0(n4783), .Y(
        \D_cache/n1483 ) );
  MX2XL U10420 ( .A(\D_cache/cache[6][38] ), .B(n10075), .S0(n4956), .Y(
        \D_cache/n1486 ) );
  MX2XL U10421 ( .A(\D_cache/cache[5][38] ), .B(n10075), .S0(n4937), .Y(
        \D_cache/n1487 ) );
  MX2XL U10422 ( .A(\D_cache/cache[4][38] ), .B(n10075), .S0(n4894), .Y(
        \D_cache/n1488 ) );
  MX2XL U10423 ( .A(\D_cache/cache[3][38] ), .B(n10075), .S0(n4847), .Y(
        \D_cache/n1489 ) );
  MX2XL U10424 ( .A(\D_cache/cache[2][38] ), .B(n10075), .S0(n4803), .Y(
        \D_cache/n1490 ) );
  MX2XL U10425 ( .A(\D_cache/cache[1][38] ), .B(n10075), .S0(n4780), .Y(
        \D_cache/n1491 ) );
  MX2XL U10426 ( .A(\D_cache/cache[0][38] ), .B(n10075), .S0(n4734), .Y(
        \D_cache/n1492 ) );
  MX2XL U10427 ( .A(\D_cache/cache[6][29] ), .B(n10683), .S0(n4957), .Y(
        \D_cache/n1558 ) );
  MX2XL U10428 ( .A(\D_cache/cache[5][29] ), .B(n10683), .S0(n4937), .Y(
        \D_cache/n1559 ) );
  MX2XL U10429 ( .A(\D_cache/cache[4][29] ), .B(n10683), .S0(n4893), .Y(
        \D_cache/n1560 ) );
  MX2XL U10430 ( .A(\D_cache/cache[3][29] ), .B(n10683), .S0(n4847), .Y(
        \D_cache/n1561 ) );
  MX2XL U10431 ( .A(\D_cache/cache[2][29] ), .B(n10683), .S0(n4802), .Y(
        \D_cache/n1562 ) );
  MX2XL U10432 ( .A(\D_cache/cache[1][29] ), .B(n10683), .S0(n4779), .Y(
        \D_cache/n1563 ) );
  MX2XL U10433 ( .A(\D_cache/cache[0][29] ), .B(n10683), .S0(n4733), .Y(
        \D_cache/n1564 ) );
  MX2XL U10434 ( .A(\D_cache/cache[6][27] ), .B(n10303), .S0(n4956), .Y(
        \D_cache/n1574 ) );
  MX2XL U10435 ( .A(\D_cache/cache[5][27] ), .B(n10303), .S0(n4937), .Y(
        \D_cache/n1575 ) );
  MX2XL U10436 ( .A(\D_cache/cache[4][27] ), .B(n10303), .S0(n4892), .Y(
        \D_cache/n1576 ) );
  MX2XL U10437 ( .A(\D_cache/cache[3][27] ), .B(n10303), .S0(n4846), .Y(
        \D_cache/n1577 ) );
  MX2XL U10438 ( .A(\D_cache/cache[2][27] ), .B(n10303), .S0(n4801), .Y(
        \D_cache/n1578 ) );
  MX2XL U10439 ( .A(\D_cache/cache[1][27] ), .B(n10303), .S0(n4778), .Y(
        \D_cache/n1579 ) );
  MX2XL U10440 ( .A(\D_cache/cache[0][27] ), .B(n10303), .S0(n4732), .Y(
        \D_cache/n1580 ) );
  MX2XL U10441 ( .A(\D_cache/cache[6][26] ), .B(n10271), .S0(n4958), .Y(
        \D_cache/n1582 ) );
  MX2XL U10442 ( .A(\D_cache/cache[5][26] ), .B(n10271), .S0(n4939), .Y(
        \D_cache/n1583 ) );
  MX2XL U10443 ( .A(\D_cache/cache[4][26] ), .B(n10271), .S0(n4895), .Y(
        \D_cache/n1584 ) );
  MX2XL U10444 ( .A(\D_cache/cache[3][26] ), .B(n10271), .S0(n4848), .Y(
        \D_cache/n1585 ) );
  MX2XL U10445 ( .A(\D_cache/cache[2][26] ), .B(n10271), .S0(n4804), .Y(
        \D_cache/n1586 ) );
  MX2XL U10446 ( .A(\D_cache/cache[1][26] ), .B(n10271), .S0(n4782), .Y(
        \D_cache/n1587 ) );
  MX2XL U10447 ( .A(\D_cache/cache[6][25] ), .B(n10493), .S0(n4956), .Y(
        \D_cache/n1590 ) );
  MX2XL U10448 ( .A(\D_cache/cache[5][25] ), .B(n10493), .S0(n4937), .Y(
        \D_cache/n1591 ) );
  MX2XL U10449 ( .A(\D_cache/cache[4][25] ), .B(n10493), .S0(n4892), .Y(
        \D_cache/n1592 ) );
  MX2XL U10450 ( .A(\D_cache/cache[3][25] ), .B(n10493), .S0(n4846), .Y(
        \D_cache/n1593 ) );
  MX2XL U10451 ( .A(\D_cache/cache[2][25] ), .B(n10493), .S0(n4801), .Y(
        \D_cache/n1594 ) );
  MX2XL U10452 ( .A(\D_cache/cache[1][25] ), .B(n10493), .S0(n4778), .Y(
        \D_cache/n1595 ) );
  MX2XL U10453 ( .A(\D_cache/cache[0][25] ), .B(n10493), .S0(n4732), .Y(
        \D_cache/n1596 ) );
  MX2XL U10454 ( .A(\D_cache/cache[6][24] ), .B(n10778), .S0(n4959), .Y(
        \D_cache/n1598 ) );
  MX2XL U10455 ( .A(\D_cache/cache[5][24] ), .B(n10778), .S0(n4939), .Y(
        \D_cache/n1599 ) );
  MX2XL U10456 ( .A(\D_cache/cache[4][24] ), .B(n10778), .S0(n4900), .Y(
        \D_cache/n1600 ) );
  MX2XL U10457 ( .A(\D_cache/cache[3][24] ), .B(n10778), .S0(n4849), .Y(
        \D_cache/n1601 ) );
  MX2XL U10458 ( .A(\D_cache/cache[2][24] ), .B(n10778), .S0(n4805), .Y(
        \D_cache/n1602 ) );
  MX2XL U10459 ( .A(\D_cache/cache[1][24] ), .B(n10778), .S0(n4782), .Y(
        \D_cache/n1603 ) );
  MX2XL U10460 ( .A(\D_cache/cache[0][24] ), .B(n10778), .S0(n4736), .Y(
        \D_cache/n1604 ) );
  MX2XL U10461 ( .A(\D_cache/cache[6][22] ), .B(n10211), .S0(n4960), .Y(
        \D_cache/n1614 ) );
  MX2XL U10462 ( .A(\D_cache/cache[5][22] ), .B(n10211), .S0(n4937), .Y(
        \D_cache/n1615 ) );
  MX2XL U10463 ( .A(\D_cache/cache[4][22] ), .B(n10211), .S0(n4894), .Y(
        \D_cache/n1616 ) );
  MX2XL U10464 ( .A(\D_cache/cache[3][22] ), .B(n10211), .S0(n4850), .Y(
        \D_cache/n1617 ) );
  MX2XL U10465 ( .A(\D_cache/cache[2][22] ), .B(n10211), .S0(n4803), .Y(
        \D_cache/n1618 ) );
  MX2XL U10466 ( .A(\D_cache/cache[1][22] ), .B(n10211), .S0(n4780), .Y(
        \D_cache/n1619 ) );
  MX2XL U10467 ( .A(\D_cache/cache[0][22] ), .B(n10211), .S0(n4734), .Y(
        \D_cache/n1620 ) );
  MX2XL U10468 ( .A(\D_cache/cache[4][20] ), .B(n10656), .S0(n4893), .Y(
        \D_cache/n1632 ) );
  MX2XL U10469 ( .A(\D_cache/cache[3][20] ), .B(n10656), .S0(n4847), .Y(
        \D_cache/n1633 ) );
  MX2XL U10470 ( .A(\D_cache/cache[2][20] ), .B(n10656), .S0(n4802), .Y(
        \D_cache/n1634 ) );
  MX2XL U10471 ( .A(\D_cache/cache[1][20] ), .B(n10656), .S0(n4779), .Y(
        \D_cache/n1635 ) );
  MX2XL U10472 ( .A(\D_cache/cache[0][20] ), .B(n10656), .S0(n4733), .Y(
        \D_cache/n1636 ) );
  MX2XL U10473 ( .A(\D_cache/cache[6][18] ), .B(n10510), .S0(n4964), .Y(
        \D_cache/n1646 ) );
  MX2XL U10474 ( .A(\D_cache/cache[5][18] ), .B(n10510), .S0(n4940), .Y(
        \D_cache/n1647 ) );
  MX2XL U10475 ( .A(\D_cache/cache[4][18] ), .B(n10510), .S0(n4898), .Y(
        \D_cache/n1648 ) );
  MX2XL U10476 ( .A(\D_cache/cache[3][18] ), .B(n10510), .S0(n4854), .Y(
        \D_cache/n1649 ) );
  MX2XL U10477 ( .A(\D_cache/cache[2][18] ), .B(n10510), .S0(n4803), .Y(
        \D_cache/n1650 ) );
  MX2XL U10478 ( .A(\D_cache/cache[1][18] ), .B(n10510), .S0(n4781), .Y(
        \D_cache/n1651 ) );
  MX2XL U10479 ( .A(\D_cache/cache[0][18] ), .B(n10510), .S0(n4733), .Y(
        \D_cache/n1652 ) );
  MX2XL U10480 ( .A(\D_cache/cache[6][17] ), .B(n10765), .S0(n4959), .Y(
        \D_cache/n1654 ) );
  MX2XL U10481 ( .A(\D_cache/cache[5][17] ), .B(n10765), .S0(n4939), .Y(
        \D_cache/n1655 ) );
  MX2XL U10482 ( .A(\D_cache/cache[4][17] ), .B(n10765), .S0(n4893), .Y(
        \D_cache/n1656 ) );
  MX2XL U10483 ( .A(\D_cache/cache[3][17] ), .B(n10765), .S0(n4849), .Y(
        \D_cache/n1657 ) );
  MX2XL U10484 ( .A(\D_cache/cache[2][17] ), .B(n10765), .S0(n4805), .Y(
        \D_cache/n1658 ) );
  MX2XL U10485 ( .A(\D_cache/cache[1][17] ), .B(n10765), .S0(n4782), .Y(
        \D_cache/n1659 ) );
  MX2XL U10486 ( .A(\D_cache/cache[6][16] ), .B(n10290), .S0(n4958), .Y(
        \D_cache/n1662 ) );
  MX2XL U10487 ( .A(\D_cache/cache[5][16] ), .B(n10290), .S0(n4939), .Y(
        \D_cache/n1663 ) );
  MX2XL U10488 ( .A(\D_cache/cache[4][16] ), .B(n10290), .S0(n4895), .Y(
        \D_cache/n1664 ) );
  MX2XL U10489 ( .A(\D_cache/cache[3][16] ), .B(n10290), .S0(n4848), .Y(
        \D_cache/n1665 ) );
  MX2XL U10490 ( .A(\D_cache/cache[2][16] ), .B(n10290), .S0(n4804), .Y(
        \D_cache/n1666 ) );
  MX2XL U10491 ( .A(\D_cache/cache[1][16] ), .B(n10290), .S0(n4782), .Y(
        \D_cache/n1667 ) );
  MX2XL U10492 ( .A(\D_cache/cache[6][15] ), .B(n10754), .S0(n4961), .Y(
        \D_cache/n1670 ) );
  MX2XL U10493 ( .A(\D_cache/cache[5][15] ), .B(n10754), .S0(n4938), .Y(
        \D_cache/n1671 ) );
  MX2XL U10494 ( .A(\D_cache/cache[4][15] ), .B(n10754), .S0(n4897), .Y(
        \D_cache/n1672 ) );
  MX2XL U10495 ( .A(\D_cache/cache[3][15] ), .B(n10754), .S0(n4851), .Y(
        \D_cache/n1673 ) );
  MX2XL U10496 ( .A(\D_cache/cache[2][15] ), .B(n10754), .S0(n4807), .Y(
        \D_cache/n1674 ) );
  MX2XL U10497 ( .A(\D_cache/cache[1][15] ), .B(n10754), .S0(n4781), .Y(
        \D_cache/n1675 ) );
  MX2XL U10498 ( .A(\D_cache/cache[0][15] ), .B(n10754), .S0(n4739), .Y(
        \D_cache/n1676 ) );
  MX2XL U10499 ( .A(\D_cache/cache[0][13] ), .B(n10732), .S0(n4739), .Y(
        \D_cache/n1692 ) );
  MX2XL U10500 ( .A(\D_cache/cache[6][12] ), .B(n10721), .S0(n4960), .Y(
        \D_cache/n1694 ) );
  MX2XL U10501 ( .A(\D_cache/cache[5][12] ), .B(n10721), .S0(n4941), .Y(
        \D_cache/n1695 ) );
  MX2XL U10502 ( .A(\D_cache/cache[4][12] ), .B(n10721), .S0(n4896), .Y(
        \D_cache/n1696 ) );
  MX2XL U10503 ( .A(\D_cache/cache[3][12] ), .B(n10721), .S0(n4850), .Y(
        \D_cache/n1697 ) );
  MX2XL U10504 ( .A(\D_cache/cache[2][12] ), .B(n10721), .S0(n4806), .Y(
        \D_cache/n1698 ) );
  MX2XL U10505 ( .A(\D_cache/cache[1][12] ), .B(n10721), .S0(n4784), .Y(
        \D_cache/n1699 ) );
  MX2XL U10506 ( .A(\D_cache/cache[0][12] ), .B(n10721), .S0(n4738), .Y(
        \D_cache/n1700 ) );
  MX2XL U10507 ( .A(\D_cache/cache[6][11] ), .B(n10709), .S0(n4960), .Y(
        \D_cache/n1702 ) );
  MX2XL U10508 ( .A(\D_cache/cache[5][11] ), .B(n10709), .S0(n4937), .Y(
        \D_cache/n1703 ) );
  MX2XL U10509 ( .A(\D_cache/cache[4][11] ), .B(n10709), .S0(n4896), .Y(
        \D_cache/n1704 ) );
  MX2XL U10510 ( .A(\D_cache/cache[3][11] ), .B(n10709), .S0(n4850), .Y(
        \D_cache/n1705 ) );
  MX2XL U10511 ( .A(\D_cache/cache[2][11] ), .B(n10709), .S0(n4806), .Y(
        \D_cache/n1706 ) );
  MX2XL U10512 ( .A(\D_cache/cache[1][11] ), .B(n10709), .S0(n4779), .Y(
        \D_cache/n1707 ) );
  MX2XL U10513 ( .A(\D_cache/cache[6][10] ), .B(n10259), .S0(n4958), .Y(
        \D_cache/n1710 ) );
  MX2XL U10514 ( .A(\D_cache/cache[5][10] ), .B(n10259), .S0(n4939), .Y(
        \D_cache/n1711 ) );
  MX2XL U10515 ( .A(\D_cache/cache[4][10] ), .B(n10259), .S0(n4895), .Y(
        \D_cache/n1712 ) );
  MX2XL U10516 ( .A(\D_cache/cache[3][10] ), .B(n10259), .S0(n4848), .Y(
        \D_cache/n1713 ) );
  MX2XL U10517 ( .A(\D_cache/cache[2][10] ), .B(n10259), .S0(n4804), .Y(
        \D_cache/n1714 ) );
  MX2XL U10518 ( .A(\D_cache/cache[1][10] ), .B(n10259), .S0(n4782), .Y(
        \D_cache/n1715 ) );
  MX2XL U10519 ( .A(\D_cache/cache[0][10] ), .B(n10259), .S0(n4735), .Y(
        \D_cache/n1716 ) );
  MX2XL U10520 ( .A(\D_cache/cache[6][9] ), .B(n10697), .S0(n4960), .Y(
        \D_cache/n1718 ) );
  MX2XL U10521 ( .A(\D_cache/cache[5][9] ), .B(n10697), .S0(n4936), .Y(
        \D_cache/n1719 ) );
  MX2XL U10522 ( .A(\D_cache/cache[4][9] ), .B(n10697), .S0(n4896), .Y(
        \D_cache/n1720 ) );
  MX2XL U10523 ( .A(\D_cache/cache[3][9] ), .B(n10697), .S0(n4850), .Y(
        \D_cache/n1721 ) );
  MX2XL U10524 ( .A(\D_cache/cache[2][9] ), .B(n10697), .S0(n4806), .Y(
        \D_cache/n1722 ) );
  MX2XL U10525 ( .A(\D_cache/cache[1][9] ), .B(n10697), .S0(n4785), .Y(
        \D_cache/n1723 ) );
  MX2XL U10526 ( .A(\D_cache/cache[0][9] ), .B(n10697), .S0(n4738), .Y(
        \D_cache/n1724 ) );
  MX2XL U10527 ( .A(\D_cache/cache[6][7] ), .B(n10883), .S0(n4958), .Y(
        \D_cache/n1734 ) );
  MX2XL U10528 ( .A(\D_cache/cache[5][7] ), .B(n10883), .S0(n4938), .Y(
        \D_cache/n1735 ) );
  MX2XL U10529 ( .A(\D_cache/cache[4][7] ), .B(n10883), .S0(n4892), .Y(
        \D_cache/n1736 ) );
  MX2XL U10530 ( .A(\D_cache/cache[3][7] ), .B(n10883), .S0(n4850), .Y(
        \D_cache/n1737 ) );
  MX2XL U10531 ( .A(\D_cache/cache[2][7] ), .B(n10883), .S0(n4804), .Y(
        \D_cache/n1738 ) );
  MX2XL U10532 ( .A(\D_cache/cache[1][7] ), .B(n10883), .S0(n4783), .Y(
        \D_cache/n1739 ) );
  MX2XL U10533 ( .A(\D_cache/cache[0][7] ), .B(n10883), .S0(n4737), .Y(
        \D_cache/n1740 ) );
  MX2XL U10534 ( .A(\D_cache/cache[6][6] ), .B(n10069), .S0(n4964), .Y(
        \D_cache/n1742 ) );
  MX2XL U10535 ( .A(\D_cache/cache[5][6] ), .B(n10069), .S0(n4937), .Y(
        \D_cache/n1743 ) );
  MX2XL U10536 ( .A(\D_cache/cache[4][6] ), .B(n10069), .S0(n4894), .Y(
        \D_cache/n1744 ) );
  MX2XL U10537 ( .A(\D_cache/cache[3][6] ), .B(n10069), .S0(n4849), .Y(
        \D_cache/n1745 ) );
  MX2XL U10538 ( .A(\D_cache/cache[2][6] ), .B(n10069), .S0(n4803), .Y(
        \D_cache/n1746 ) );
  MX2XL U10539 ( .A(\D_cache/cache[1][6] ), .B(n10069), .S0(n4780), .Y(
        \D_cache/n1747 ) );
  MX2XL U10540 ( .A(\D_cache/cache[6][3] ), .B(n9992), .S0(n4962), .Y(
        \D_cache/n1766 ) );
  MX2XL U10541 ( .A(\D_cache/cache[5][3] ), .B(n9992), .S0(n4941), .Y(
        \D_cache/n1767 ) );
  MX2XL U10542 ( .A(\D_cache/cache[4][3] ), .B(n9992), .S0(n4898), .Y(
        \D_cache/n1768 ) );
  MX2XL U10543 ( .A(\D_cache/cache[3][3] ), .B(n9992), .S0(n4852), .Y(
        \D_cache/n1769 ) );
  MX2XL U10544 ( .A(\D_cache/cache[2][3] ), .B(n9992), .S0(n4808), .Y(
        \D_cache/n1770 ) );
  MX2XL U10545 ( .A(\D_cache/cache[1][3] ), .B(n9992), .S0(n4784), .Y(
        \D_cache/n1771 ) );
  MX2XL U10546 ( .A(\D_cache/cache[6][127] ), .B(n10876), .S0(n4958), .Y(
        \D_cache/n774 ) );
  MX2XL U10547 ( .A(\D_cache/cache[5][127] ), .B(n10876), .S0(n4939), .Y(
        \D_cache/n775 ) );
  MX2XL U10548 ( .A(\D_cache/cache[4][127] ), .B(n10876), .S0(n4895), .Y(
        \D_cache/n776 ) );
  MX2XL U10549 ( .A(\D_cache/cache[3][127] ), .B(n10876), .S0(n4848), .Y(
        \D_cache/n777 ) );
  MX2XL U10550 ( .A(\D_cache/cache[2][127] ), .B(n10876), .S0(n4804), .Y(
        \D_cache/n778 ) );
  MX2XL U10551 ( .A(\D_cache/cache[1][127] ), .B(n10876), .S0(n4782), .Y(
        \D_cache/n779 ) );
  MX2XL U10552 ( .A(\D_cache/cache[0][127] ), .B(n10876), .S0(n4735), .Y(
        \D_cache/n780 ) );
  MX2XL U10553 ( .A(\D_cache/cache[6][125] ), .B(n10689), .S0(n4960), .Y(
        \D_cache/n790 ) );
  MX2XL U10554 ( .A(\D_cache/cache[5][125] ), .B(n10689), .S0(n4942), .Y(
        \D_cache/n791 ) );
  MX2XL U10555 ( .A(\D_cache/cache[4][125] ), .B(n10689), .S0(n4896), .Y(
        \D_cache/n792 ) );
  MX2XL U10556 ( .A(\D_cache/cache[3][125] ), .B(n10689), .S0(n4850), .Y(
        \D_cache/n793 ) );
  MX2XL U10557 ( .A(\D_cache/cache[2][125] ), .B(n10689), .S0(n4806), .Y(
        \D_cache/n794 ) );
  MX2XL U10558 ( .A(\D_cache/cache[1][125] ), .B(n10689), .S0(n4781), .Y(
        \D_cache/n795 ) );
  MX2XL U10559 ( .A(\D_cache/cache[0][125] ), .B(n10689), .S0(n4738), .Y(
        \D_cache/n796 ) );
  MX2XL U10560 ( .A(\D_cache/cache[5][124] ), .B(n10483), .S0(n4937), .Y(
        \D_cache/n799 ) );
  MX2XL U10561 ( .A(\D_cache/cache[4][124] ), .B(n10483), .S0(n4892), .Y(
        \D_cache/n800 ) );
  MX2XL U10562 ( .A(\D_cache/cache[3][124] ), .B(n10483), .S0(n4846), .Y(
        \D_cache/n801 ) );
  MX2XL U10563 ( .A(\D_cache/cache[2][124] ), .B(n10483), .S0(n4801), .Y(
        \D_cache/n802 ) );
  MX2XL U10564 ( .A(\D_cache/cache[1][124] ), .B(n10483), .S0(n4778), .Y(
        \D_cache/n803 ) );
  MX2XL U10565 ( .A(\D_cache/cache[0][124] ), .B(n10483), .S0(n4732), .Y(
        \D_cache/n804 ) );
  MX2XL U10566 ( .A(\D_cache/cache[6][120] ), .B(n10784), .S0(n4959), .Y(
        \D_cache/n830 ) );
  MX2XL U10567 ( .A(\D_cache/cache[5][120] ), .B(n10784), .S0(n4939), .Y(
        \D_cache/n831 ) );
  MX2XL U10568 ( .A(\D_cache/cache[4][120] ), .B(n10784), .S0(n4895), .Y(
        \D_cache/n832 ) );
  MX2XL U10569 ( .A(\D_cache/cache[3][120] ), .B(n10784), .S0(n4849), .Y(
        \D_cache/n833 ) );
  MX2XL U10570 ( .A(\D_cache/cache[2][120] ), .B(n10784), .S0(n4805), .Y(
        \D_cache/n834 ) );
  MX2XL U10571 ( .A(\D_cache/cache[1][120] ), .B(n10784), .S0(n4782), .Y(
        \D_cache/n835 ) );
  MX2XL U10572 ( .A(\D_cache/cache[0][120] ), .B(n10784), .S0(n4736), .Y(
        \D_cache/n836 ) );
  MX2XL U10573 ( .A(\D_cache/cache[5][117] ), .B(n10675), .S0(n4937), .Y(
        \D_cache/n855 ) );
  MX2XL U10574 ( .A(\D_cache/cache[4][117] ), .B(n10675), .S0(n4893), .Y(
        \D_cache/n856 ) );
  MX2XL U10575 ( .A(\D_cache/cache[3][117] ), .B(n10675), .S0(n4847), .Y(
        \D_cache/n857 ) );
  MX2XL U10576 ( .A(\D_cache/cache[2][117] ), .B(n10675), .S0(n4802), .Y(
        \D_cache/n858 ) );
  MX2XL U10577 ( .A(\D_cache/cache[1][117] ), .B(n10675), .S0(n4779), .Y(
        \D_cache/n859 ) );
  MX2XL U10578 ( .A(\D_cache/cache[0][117] ), .B(n10675), .S0(n4733), .Y(
        \D_cache/n860 ) );
  MX2XL U10579 ( .A(\D_cache/cache[6][113] ), .B(n10771), .S0(n4959), .Y(
        \D_cache/n886 ) );
  MX2XL U10580 ( .A(\D_cache/cache[5][113] ), .B(n10771), .S0(n4939), .Y(
        \D_cache/n887 ) );
  MX2XL U10581 ( .A(\D_cache/cache[4][113] ), .B(n10771), .S0(n4898), .Y(
        \D_cache/n888 ) );
  MX2XL U10582 ( .A(\D_cache/cache[3][113] ), .B(n10771), .S0(n4849), .Y(
        \D_cache/n889 ) );
  MX2XL U10583 ( .A(\D_cache/cache[2][113] ), .B(n10771), .S0(n4805), .Y(
        \D_cache/n890 ) );
  MX2XL U10584 ( .A(\D_cache/cache[1][113] ), .B(n10771), .S0(n4782), .Y(
        \D_cache/n891 ) );
  MX2XL U10585 ( .A(\D_cache/cache[0][113] ), .B(n10771), .S0(n4736), .Y(
        \D_cache/n892 ) );
  MX2XL U10586 ( .A(\D_cache/cache[6][111] ), .B(n10760), .S0(n4961), .Y(
        \D_cache/n902 ) );
  MX2XL U10587 ( .A(\D_cache/cache[5][111] ), .B(n10760), .S0(n4936), .Y(
        \D_cache/n903 ) );
  MX2XL U10588 ( .A(\D_cache/cache[4][111] ), .B(n10760), .S0(n4897), .Y(
        \D_cache/n904 ) );
  MX2XL U10589 ( .A(\D_cache/cache[3][111] ), .B(n10760), .S0(n4851), .Y(
        \D_cache/n905 ) );
  MX2XL U10590 ( .A(\D_cache/cache[2][111] ), .B(n10760), .S0(n4807), .Y(
        \D_cache/n906 ) );
  MX2XL U10591 ( .A(\D_cache/cache[1][111] ), .B(n10760), .S0(n4784), .Y(
        \D_cache/n907 ) );
  MX2XL U10592 ( .A(\D_cache/cache[0][111] ), .B(n10760), .S0(n4738), .Y(
        \D_cache/n908 ) );
  MX2XL U10593 ( .A(\D_cache/cache[6][110] ), .B(n10749), .S0(n4961), .Y(
        \D_cache/n910 ) );
  MX2XL U10594 ( .A(\D_cache/cache[5][110] ), .B(n10749), .S0(n4938), .Y(
        \D_cache/n911 ) );
  MX2XL U10595 ( .A(\D_cache/cache[4][110] ), .B(n10749), .S0(n4897), .Y(
        \D_cache/n912 ) );
  MX2XL U10596 ( .A(\D_cache/cache[3][110] ), .B(n10749), .S0(n4851), .Y(
        \D_cache/n913 ) );
  MX2XL U10597 ( .A(\D_cache/cache[2][110] ), .B(n10749), .S0(n4807), .Y(
        \D_cache/n914 ) );
  MX2XL U10598 ( .A(\D_cache/cache[1][110] ), .B(n10749), .S0(n4784), .Y(
        \D_cache/n915 ) );
  MX2XL U10599 ( .A(\D_cache/cache[0][110] ), .B(n10749), .S0(n4739), .Y(
        \D_cache/n916 ) );
  MX2XL U10600 ( .A(\D_cache/cache[6][109] ), .B(n10738), .S0(n4961), .Y(
        \D_cache/n918 ) );
  MX2XL U10601 ( .A(\D_cache/cache[5][109] ), .B(n10738), .S0(n4940), .Y(
        \D_cache/n919 ) );
  MX2XL U10602 ( .A(\D_cache/cache[4][109] ), .B(n10738), .S0(n4897), .Y(
        \D_cache/n920 ) );
  MX2XL U10603 ( .A(\D_cache/cache[3][109] ), .B(n10738), .S0(n4851), .Y(
        \D_cache/n921 ) );
  MX2XL U10604 ( .A(\D_cache/cache[2][109] ), .B(n10738), .S0(n4807), .Y(
        \D_cache/n922 ) );
  MX2XL U10605 ( .A(\D_cache/cache[1][109] ), .B(n10738), .S0(n4785), .Y(
        \D_cache/n923 ) );
  MX2XL U10606 ( .A(\D_cache/cache[0][109] ), .B(n10738), .S0(n4739), .Y(
        \D_cache/n924 ) );
  MX2XL U10607 ( .A(\D_cache/cache[0][108] ), .B(n10727), .S0(n4739), .Y(
        \D_cache/n932 ) );
  MX2XL U10608 ( .A(\D_cache/cache[6][106] ), .B(n10265), .S0(n4958), .Y(
        \D_cache/n942 ) );
  MX2XL U10609 ( .A(\D_cache/cache[5][106] ), .B(n10265), .S0(n4938), .Y(
        \D_cache/n943 ) );
  MX2XL U10610 ( .A(\D_cache/cache[4][106] ), .B(n10265), .S0(n4895), .Y(
        \D_cache/n944 ) );
  MX2XL U10611 ( .A(\D_cache/cache[3][106] ), .B(n10265), .S0(n4848), .Y(
        \D_cache/n945 ) );
  MX2XL U10612 ( .A(\D_cache/cache[2][106] ), .B(n10265), .S0(n4804), .Y(
        \D_cache/n946 ) );
  MX2XL U10613 ( .A(\D_cache/cache[1][106] ), .B(n10265), .S0(n4781), .Y(
        \D_cache/n947 ) );
  MX2XL U10614 ( .A(\D_cache/cache[0][106] ), .B(n10265), .S0(n4735), .Y(
        \D_cache/n948 ) );
  MX2XL U10615 ( .A(\D_cache/cache[3][105] ), .B(n10703), .S0(n4850), .Y(
        \D_cache/n953 ) );
  MX2XL U10616 ( .A(\D_cache/cache[2][105] ), .B(n10703), .S0(n4806), .Y(
        \D_cache/n954 ) );
  MX2XL U10617 ( .A(\D_cache/cache[1][105] ), .B(n10703), .S0(n4778), .Y(
        \D_cache/n955 ) );
  MX2XL U10618 ( .A(\D_cache/cache[0][105] ), .B(n10703), .S0(n4738), .Y(
        \D_cache/n956 ) );
  MX2XL U10619 ( .A(\D_cache/cache[6][104] ), .B(n10901), .S0(n4957), .Y(
        \D_cache/n958 ) );
  MX2XL U10620 ( .A(\D_cache/cache[5][104] ), .B(n10901), .S0(n4940), .Y(
        \D_cache/n959 ) );
  MX2XL U10621 ( .A(\D_cache/cache[4][104] ), .B(n10901), .S0(n4893), .Y(
        \D_cache/n960 ) );
  MX2XL U10622 ( .A(\D_cache/cache[3][104] ), .B(n10901), .S0(n4846), .Y(
        \D_cache/n961 ) );
  MX2XL U10623 ( .A(\D_cache/cache[2][104] ), .B(n10901), .S0(n4805), .Y(
        \D_cache/n962 ) );
  MX2XL U10624 ( .A(\D_cache/cache[1][104] ), .B(n10901), .S0(n4781), .Y(
        \D_cache/n963 ) );
  MX2XL U10625 ( .A(\D_cache/cache[0][104] ), .B(n10901), .S0(n4737), .Y(
        \D_cache/n964 ) );
  MX2XL U10626 ( .A(\D_cache/cache[6][103] ), .B(n10889), .S0(n4957), .Y(
        \D_cache/n966 ) );
  MX2XL U10627 ( .A(\D_cache/cache[5][103] ), .B(n10889), .S0(n4938), .Y(
        \D_cache/n967 ) );
  MX2XL U10628 ( .A(\D_cache/cache[4][103] ), .B(n10889), .S0(n4895), .Y(
        \D_cache/n968 ) );
  MX2XL U10629 ( .A(\D_cache/cache[3][103] ), .B(n10889), .S0(n4849), .Y(
        \D_cache/n969 ) );
  MX2XL U10630 ( .A(\D_cache/cache[2][103] ), .B(n10889), .S0(n4806), .Y(
        \D_cache/n970 ) );
  MX2XL U10631 ( .A(\D_cache/cache[1][103] ), .B(n10889), .S0(n4783), .Y(
        \D_cache/n971 ) );
  MX2XL U10632 ( .A(\D_cache/cache[0][103] ), .B(n10889), .S0(n4737), .Y(
        \D_cache/n972 ) );
  MX2XL U10633 ( .A(\D_cache/cache[6][92] ), .B(n10486), .S0(n4956), .Y(
        \D_cache/n1054 ) );
  MX2XL U10634 ( .A(\D_cache/cache[5][92] ), .B(n10486), .S0(n4936), .Y(
        \D_cache/n1055 ) );
  MX2XL U10635 ( .A(\D_cache/cache[4][92] ), .B(n10486), .S0(n4892), .Y(
        \D_cache/n1056 ) );
  MX2XL U10636 ( .A(\D_cache/cache[3][92] ), .B(n10486), .S0(n4846), .Y(
        \D_cache/n1057 ) );
  MX2XL U10637 ( .A(\D_cache/cache[2][92] ), .B(n10486), .S0(n4801), .Y(
        \D_cache/n1058 ) );
  MX2XL U10638 ( .A(\D_cache/cache[1][92] ), .B(n10486), .S0(n4778), .Y(
        \D_cache/n1059 ) );
  MX2XL U10639 ( .A(\D_cache/cache[0][92] ), .B(n10486), .S0(n4732), .Y(
        \D_cache/n1060 ) );
  MX2XL U10640 ( .A(\D_cache/cache[6][91] ), .B(n10312), .S0(n4956), .Y(
        \D_cache/n1062 ) );
  MX2XL U10641 ( .A(\D_cache/cache[5][91] ), .B(n10312), .S0(n4940), .Y(
        \D_cache/n1063 ) );
  MX2XL U10642 ( .A(\D_cache/cache[4][91] ), .B(n10312), .S0(n4892), .Y(
        \D_cache/n1064 ) );
  MX2XL U10643 ( .A(\D_cache/cache[3][91] ), .B(n10312), .S0(n4846), .Y(
        \D_cache/n1065 ) );
  MX2XL U10644 ( .A(\D_cache/cache[2][91] ), .B(n10312), .S0(n4801), .Y(
        \D_cache/n1066 ) );
  MX2XL U10645 ( .A(\D_cache/cache[1][91] ), .B(n10312), .S0(n4778), .Y(
        \D_cache/n1067 ) );
  MX2XL U10646 ( .A(\D_cache/cache[0][91] ), .B(n10312), .S0(n4732), .Y(
        \D_cache/n1068 ) );
  MX2XL U10647 ( .A(\D_cache/cache[6][90] ), .B(n10280), .S0(n4958), .Y(
        \D_cache/n1070 ) );
  MX2XL U10648 ( .A(\D_cache/cache[5][90] ), .B(n10280), .S0(n4940), .Y(
        \D_cache/n1071 ) );
  MX2XL U10649 ( .A(\D_cache/cache[4][90] ), .B(n10280), .S0(n4895), .Y(
        \D_cache/n1072 ) );
  MX2XL U10650 ( .A(\D_cache/cache[3][90] ), .B(n10280), .S0(n4848), .Y(
        \D_cache/n1073 ) );
  MX2XL U10651 ( .A(\D_cache/cache[2][90] ), .B(n10280), .S0(n4804), .Y(
        \D_cache/n1074 ) );
  MX2XL U10652 ( .A(\D_cache/cache[1][90] ), .B(n10280), .S0(n4783), .Y(
        \D_cache/n1075 ) );
  MX2XL U10653 ( .A(\D_cache/cache[0][90] ), .B(n10280), .S0(n4735), .Y(
        \D_cache/n1076 ) );
  MX2XL U10654 ( .A(\D_cache/cache[6][86] ), .B(n10220), .S0(n4958), .Y(
        \D_cache/n1102 ) );
  MX2XL U10655 ( .A(\D_cache/cache[5][86] ), .B(n10220), .S0(n4938), .Y(
        \D_cache/n1103 ) );
  MX2XL U10656 ( .A(\D_cache/cache[4][86] ), .B(n10220), .S0(n4895), .Y(
        \D_cache/n1104 ) );
  MX2XL U10657 ( .A(\D_cache/cache[3][86] ), .B(n10220), .S0(n4848), .Y(
        \D_cache/n1105 ) );
  MX2XL U10658 ( .A(\D_cache/cache[2][86] ), .B(n10220), .S0(n4804), .Y(
        \D_cache/n1106 ) );
  MX2XL U10659 ( .A(\D_cache/cache[1][86] ), .B(n10220), .S0(n4781), .Y(
        \D_cache/n1107 ) );
  MX2XL U10660 ( .A(\D_cache/cache[0][86] ), .B(n10220), .S0(n4735), .Y(
        \D_cache/n1108 ) );
  MX2XL U10661 ( .A(\D_cache/cache[6][80] ), .B(n10299), .S0(n4956), .Y(
        \D_cache/n1150 ) );
  MX2XL U10662 ( .A(\D_cache/cache[5][80] ), .B(n10299), .S0(n4937), .Y(
        \D_cache/n1151 ) );
  MX2XL U10663 ( .A(\D_cache/cache[4][80] ), .B(n10299), .S0(n4894), .Y(
        \D_cache/n1152 ) );
  MX2XL U10664 ( .A(\D_cache/cache[3][80] ), .B(n10299), .S0(n4850), .Y(
        \D_cache/n1153 ) );
  MX2XL U10665 ( .A(\D_cache/cache[2][80] ), .B(n10299), .S0(n4803), .Y(
        \D_cache/n1154 ) );
  MX2XL U10666 ( .A(\D_cache/cache[1][80] ), .B(n10299), .S0(n4780), .Y(
        \D_cache/n1155 ) );
  MX2XL U10667 ( .A(\D_cache/cache[0][80] ), .B(n10299), .S0(n4732), .Y(
        \D_cache/n1156 ) );
  MX2XL U10668 ( .A(\D_cache/cache[6][74] ), .B(n10268), .S0(n4958), .Y(
        \D_cache/n1198 ) );
  MX2XL U10669 ( .A(\D_cache/cache[5][74] ), .B(n10268), .S0(n4940), .Y(
        \D_cache/n1199 ) );
  MX2XL U10670 ( .A(\D_cache/cache[4][74] ), .B(n10268), .S0(n4895), .Y(
        \D_cache/n1200 ) );
  MX2XL U10671 ( .A(\D_cache/cache[3][74] ), .B(n10268), .S0(n4848), .Y(
        \D_cache/n1201 ) );
  MX2XL U10672 ( .A(\D_cache/cache[2][74] ), .B(n10268), .S0(n4804), .Y(
        \D_cache/n1202 ) );
  MX2XL U10673 ( .A(\D_cache/cache[1][74] ), .B(n10268), .S0(n4783), .Y(
        \D_cache/n1203 ) );
  MX2XL U10674 ( .A(\D_cache/cache[0][74] ), .B(n10268), .S0(n4735), .Y(
        \D_cache/n1204 ) );
  MX2XL U10675 ( .A(\D_cache/cache[6][73] ), .B(n10706), .S0(n4960), .Y(
        \D_cache/n1206 ) );
  MX2XL U10676 ( .A(\D_cache/cache[5][73] ), .B(n10706), .S0(n4937), .Y(
        \D_cache/n1207 ) );
  MX2XL U10677 ( .A(\D_cache/cache[4][73] ), .B(n10706), .S0(n4896), .Y(
        \D_cache/n1208 ) );
  MX2XL U10678 ( .A(\D_cache/cache[3][73] ), .B(n10706), .S0(n4850), .Y(
        \D_cache/n1209 ) );
  MX2XL U10679 ( .A(\D_cache/cache[2][73] ), .B(n10706), .S0(n4806), .Y(
        \D_cache/n1210 ) );
  MX2XL U10680 ( .A(\D_cache/cache[1][73] ), .B(n10706), .S0(n4779), .Y(
        \D_cache/n1211 ) );
  MX2XL U10681 ( .A(\D_cache/cache[0][73] ), .B(n10706), .S0(n4738), .Y(
        \D_cache/n1212 ) );
  MX2XL U10682 ( .A(\D_cache/cache[6][72] ), .B(n4244), .S0(n4956), .Y(
        \D_cache/n1214 ) );
  MX2XL U10683 ( .A(\D_cache/cache[5][72] ), .B(n4244), .S0(n4938), .Y(
        \D_cache/n1215 ) );
  MX2XL U10684 ( .A(\D_cache/cache[4][72] ), .B(n4244), .S0(n4895), .Y(
        \D_cache/n1216 ) );
  MX2XL U10685 ( .A(\D_cache/cache[3][72] ), .B(n4244), .S0(n4847), .Y(
        \D_cache/n1217 ) );
  MX2XL U10686 ( .A(\D_cache/cache[2][72] ), .B(n4244), .S0(n4801), .Y(
        \D_cache/n1218 ) );
  MX2XL U10687 ( .A(\D_cache/cache[1][72] ), .B(n4244), .S0(n4781), .Y(
        \D_cache/n1219 ) );
  MX2XL U10688 ( .A(\D_cache/cache[0][72] ), .B(n4244), .S0(n4737), .Y(
        \D_cache/n1220 ) );
  MX2XL U10689 ( .A(\D_cache/cache[6][71] ), .B(n10892), .S0(n4959), .Y(
        \D_cache/n1222 ) );
  MX2XL U10690 ( .A(\D_cache/cache[5][71] ), .B(n10892), .S0(n4940), .Y(
        \D_cache/n1223 ) );
  MX2XL U10691 ( .A(\D_cache/cache[4][71] ), .B(n10892), .S0(n4894), .Y(
        \D_cache/n1224 ) );
  MX2XL U10692 ( .A(\D_cache/cache[3][71] ), .B(n10892), .S0(n4848), .Y(
        \D_cache/n1225 ) );
  MX2XL U10693 ( .A(\D_cache/cache[2][71] ), .B(n10892), .S0(n4802), .Y(
        \D_cache/n1226 ) );
  MX2XL U10694 ( .A(\D_cache/cache[1][71] ), .B(n10892), .S0(n4783), .Y(
        \D_cache/n1227 ) );
  MX2XL U10695 ( .A(\D_cache/cache[0][71] ), .B(n10892), .S0(n4737), .Y(
        \D_cache/n1228 ) );
  MX2XL U10696 ( .A(\D_cache/cache[6][37] ), .B(n10983), .S0(n4965), .Y(
        \D_cache/n1494 ) );
  MX2XL U10697 ( .A(\D_cache/cache[5][37] ), .B(n10983), .S0(n4944), .Y(
        \D_cache/n1495 ) );
  MX2XL U10698 ( .A(\D_cache/cache[4][37] ), .B(n10983), .S0(n4901), .Y(
        \D_cache/n1496 ) );
  MX2XL U10699 ( .A(\D_cache/cache[3][37] ), .B(n10983), .S0(n4855), .Y(
        \D_cache/n1497 ) );
  MX2XL U10700 ( .A(\D_cache/cache[2][37] ), .B(n10983), .S0(n4805), .Y(
        \D_cache/n1498 ) );
  MX2XL U10701 ( .A(\D_cache/cache[1][37] ), .B(n10983), .S0(n4786), .Y(
        \D_cache/n1499 ) );
  MX2XL U10702 ( .A(\D_cache/cache[0][37] ), .B(n10983), .S0(n4739), .Y(
        \D_cache/n1500 ) );
  MX2XL U10703 ( .A(\D_cache/cache[6][36] ), .B(n10971), .S0(n4965), .Y(
        \D_cache/n1502 ) );
  MX2XL U10704 ( .A(\D_cache/cache[5][36] ), .B(n10971), .S0(n4944), .Y(
        \D_cache/n1503 ) );
  MX2XL U10705 ( .A(\D_cache/cache[4][36] ), .B(n10971), .S0(n4901), .Y(
        \D_cache/n1504 ) );
  MX2XL U10706 ( .A(\D_cache/cache[3][36] ), .B(n10971), .S0(n4855), .Y(
        \D_cache/n1505 ) );
  MX2XL U10707 ( .A(\D_cache/cache[2][36] ), .B(n10971), .S0(n4806), .Y(
        \D_cache/n1506 ) );
  MX2XL U10708 ( .A(\D_cache/cache[1][36] ), .B(n10971), .S0(n4786), .Y(
        \D_cache/n1507 ) );
  MX2XL U10709 ( .A(\D_cache/cache[0][36] ), .B(n10971), .S0(n4732), .Y(
        \D_cache/n1508 ) );
  MX2XL U10710 ( .A(\D_cache/cache[6][35] ), .B(n10919), .S0(n4959), .Y(
        \D_cache/n1510 ) );
  MX2XL U10711 ( .A(\D_cache/cache[5][35] ), .B(n10919), .S0(n4939), .Y(
        \D_cache/n1511 ) );
  MX2XL U10712 ( .A(\D_cache/cache[4][35] ), .B(n10919), .S0(n4900), .Y(
        \D_cache/n1512 ) );
  MX2XL U10713 ( .A(\D_cache/cache[3][35] ), .B(n10919), .S0(n4849), .Y(
        \D_cache/n1513 ) );
  MX2XL U10714 ( .A(\D_cache/cache[2][35] ), .B(n10919), .S0(n4805), .Y(
        \D_cache/n1514 ) );
  MX2XL U10715 ( .A(\D_cache/cache[1][35] ), .B(n10919), .S0(n4782), .Y(
        \D_cache/n1515 ) );
  MX2XL U10716 ( .A(\D_cache/cache[0][35] ), .B(n10919), .S0(n4741), .Y(
        \D_cache/n1516 ) );
  MX2XL U10717 ( .A(\D_cache/cache[6][34] ), .B(n10933), .S0(n4964), .Y(
        \D_cache/n1518 ) );
  MX2XL U10718 ( .A(\D_cache/cache[5][34] ), .B(n10933), .S0(n4943), .Y(
        \D_cache/n1519 ) );
  MX2XL U10719 ( .A(\D_cache/cache[4][34] ), .B(n10933), .S0(n4900), .Y(
        \D_cache/n1520 ) );
  MX2XL U10720 ( .A(\D_cache/cache[3][34] ), .B(n10933), .S0(n4854), .Y(
        \D_cache/n1521 ) );
  MX2XL U10721 ( .A(\D_cache/cache[2][34] ), .B(n10933), .S0(n4809), .Y(
        \D_cache/n1522 ) );
  MX2XL U10722 ( .A(\D_cache/cache[1][34] ), .B(n10933), .S0(n4783), .Y(
        \D_cache/n1523 ) );
  MX2XL U10723 ( .A(\D_cache/cache[0][34] ), .B(n10933), .S0(n4741), .Y(
        \D_cache/n1524 ) );
  MX2XL U10724 ( .A(\D_cache/cache[6][33] ), .B(n10910), .S0(n4958), .Y(
        \D_cache/n1526 ) );
  MX2XL U10725 ( .A(\D_cache/cache[5][33] ), .B(n10910), .S0(n4938), .Y(
        \D_cache/n1527 ) );
  MX2XL U10726 ( .A(\D_cache/cache[4][33] ), .B(n10910), .S0(n4895), .Y(
        \D_cache/n1528 ) );
  MX2XL U10727 ( .A(\D_cache/cache[3][33] ), .B(n10910), .S0(n4849), .Y(
        \D_cache/n1529 ) );
  MX2XL U10728 ( .A(\D_cache/cache[2][33] ), .B(n10910), .S0(n4804), .Y(
        \D_cache/n1530 ) );
  MX2XL U10729 ( .A(\D_cache/cache[1][33] ), .B(n10910), .S0(n4781), .Y(
        \D_cache/n1531 ) );
  MX2XL U10730 ( .A(\D_cache/cache[0][33] ), .B(n10910), .S0(n4737), .Y(
        \D_cache/n1532 ) );
  MX2XL U10731 ( .A(\D_cache/cache[0][8] ), .B(n169), .S0(n4737), .Y(
        \D_cache/n1732 ) );
  MX2XL U10732 ( .A(\D_cache/cache[6][5] ), .B(n10980), .S0(n4965), .Y(
        \D_cache/n1750 ) );
  MX2XL U10733 ( .A(\D_cache/cache[5][5] ), .B(n10980), .S0(n4944), .Y(
        \D_cache/n1751 ) );
  MX2XL U10734 ( .A(\D_cache/cache[4][5] ), .B(n10980), .S0(n4901), .Y(
        \D_cache/n1752 ) );
  MX2XL U10735 ( .A(\D_cache/cache[3][5] ), .B(n10980), .S0(n4855), .Y(
        \D_cache/n1753 ) );
  MX2XL U10736 ( .A(\D_cache/cache[2][5] ), .B(n10980), .S0(n4804), .Y(
        \D_cache/n1754 ) );
  MX2XL U10737 ( .A(\D_cache/cache[1][5] ), .B(n10980), .S0(n4786), .Y(
        \D_cache/n1755 ) );
  MX2XL U10738 ( .A(\D_cache/cache[0][5] ), .B(n10980), .S0(n4736), .Y(
        \D_cache/n1756 ) );
  MX2XL U10739 ( .A(\D_cache/cache[6][2] ), .B(n10930), .S0(n4964), .Y(
        \D_cache/n1774 ) );
  MX2XL U10740 ( .A(\D_cache/cache[5][2] ), .B(n10930), .S0(n4943), .Y(
        \D_cache/n1775 ) );
  MX2XL U10741 ( .A(\D_cache/cache[4][2] ), .B(n10930), .S0(n4900), .Y(
        \D_cache/n1776 ) );
  MX2XL U10742 ( .A(\D_cache/cache[3][2] ), .B(n10930), .S0(n4854), .Y(
        \D_cache/n1777 ) );
  MX2XL U10743 ( .A(\D_cache/cache[2][2] ), .B(n10930), .S0(n4809), .Y(
        \D_cache/n1778 ) );
  MX2XL U10744 ( .A(\D_cache/cache[1][2] ), .B(n10930), .S0(n4786), .Y(
        \D_cache/n1779 ) );
  MX2XL U10745 ( .A(\D_cache/cache[0][2] ), .B(n10930), .S0(n4741), .Y(
        \D_cache/n1780 ) );
  MX2XL U10746 ( .A(\D_cache/cache[6][1] ), .B(n10907), .S0(n4956), .Y(
        \D_cache/n1782 ) );
  MX2XL U10747 ( .A(\D_cache/cache[5][1] ), .B(n10907), .S0(n4940), .Y(
        \D_cache/n1783 ) );
  MX2XL U10748 ( .A(\D_cache/cache[4][1] ), .B(n10907), .S0(n4898), .Y(
        \D_cache/n1784 ) );
  MX2XL U10749 ( .A(\D_cache/cache[3][1] ), .B(n10907), .S0(n4854), .Y(
        \D_cache/n1785 ) );
  MX2XL U10750 ( .A(\D_cache/cache[2][1] ), .B(n10907), .S0(n4805), .Y(
        \D_cache/n1786 ) );
  MX2XL U10751 ( .A(\D_cache/cache[1][1] ), .B(n10907), .S0(n4783), .Y(
        \D_cache/n1787 ) );
  MX2XL U10752 ( .A(\D_cache/cache[0][1] ), .B(n10907), .S0(n4737), .Y(
        \D_cache/n1788 ) );
  MX2XL U10753 ( .A(\D_cache/cache[6][68] ), .B(n10977), .S0(n4965), .Y(
        \D_cache/n1246 ) );
  MX2XL U10754 ( .A(\D_cache/cache[5][68] ), .B(n10977), .S0(n4944), .Y(
        \D_cache/n1247 ) );
  MX2XL U10755 ( .A(\D_cache/cache[4][68] ), .B(n10977), .S0(n4901), .Y(
        \D_cache/n1248 ) );
  MX2XL U10756 ( .A(\D_cache/cache[3][68] ), .B(n10977), .S0(n4855), .Y(
        \D_cache/n1249 ) );
  MX2XL U10757 ( .A(\D_cache/cache[2][68] ), .B(n10977), .S0(n4801), .Y(
        \D_cache/n1250 ) );
  MX2XL U10758 ( .A(\D_cache/cache[1][68] ), .B(n10977), .S0(n4786), .Y(
        \D_cache/n1251 ) );
  MX2XL U10759 ( .A(\D_cache/cache[0][68] ), .B(n10977), .S0(n4735), .Y(
        \D_cache/n1252 ) );
  MX2XL U10760 ( .A(\D_cache/cache[6][67] ), .B(n10925), .S0(n4964), .Y(
        \D_cache/n1254 ) );
  MX2XL U10761 ( .A(\D_cache/cache[5][67] ), .B(n10925), .S0(n4943), .Y(
        \D_cache/n1255 ) );
  MX2XL U10762 ( .A(\D_cache/cache[4][67] ), .B(n10925), .S0(n4900), .Y(
        \D_cache/n1256 ) );
  MX2XL U10763 ( .A(\D_cache/cache[3][67] ), .B(n10925), .S0(n4854), .Y(
        \D_cache/n1257 ) );
  MX2XL U10764 ( .A(\D_cache/cache[2][67] ), .B(n10925), .S0(n4809), .Y(
        \D_cache/n1258 ) );
  MX2XL U10765 ( .A(\D_cache/cache[1][67] ), .B(n10925), .S0(n4778), .Y(
        \D_cache/n1259 ) );
  MX2XL U10766 ( .A(\D_cache/cache[0][67] ), .B(n10925), .S0(n4741), .Y(
        \D_cache/n1260 ) );
  MX2XL U10767 ( .A(\D_cache/cache[6][66] ), .B(n10939), .S0(n4964), .Y(
        \D_cache/n1262 ) );
  MX2XL U10768 ( .A(\D_cache/cache[5][66] ), .B(n10939), .S0(n4943), .Y(
        \D_cache/n1263 ) );
  MX2XL U10769 ( .A(\D_cache/cache[4][66] ), .B(n10939), .S0(n4900), .Y(
        \D_cache/n1264 ) );
  MX2XL U10770 ( .A(\D_cache/cache[3][66] ), .B(n10939), .S0(n4854), .Y(
        \D_cache/n1265 ) );
  MX2XL U10771 ( .A(\D_cache/cache[2][66] ), .B(n10939), .S0(n4809), .Y(
        \D_cache/n1266 ) );
  MX2XL U10772 ( .A(\D_cache/cache[1][66] ), .B(n10939), .S0(n4779), .Y(
        \D_cache/n1267 ) );
  MX2XL U10773 ( .A(\D_cache/cache[0][66] ), .B(n10939), .S0(n4741), .Y(
        \D_cache/n1268 ) );
  MX2XL U10774 ( .A(\D_cache/cache[6][65] ), .B(n10916), .S0(n4959), .Y(
        \D_cache/n1270 ) );
  MX2XL U10775 ( .A(\D_cache/cache[5][65] ), .B(n10916), .S0(n4939), .Y(
        \D_cache/n1271 ) );
  MX2XL U10776 ( .A(\D_cache/cache[4][65] ), .B(n10916), .S0(n4893), .Y(
        \D_cache/n1272 ) );
  MX2XL U10777 ( .A(\D_cache/cache[3][65] ), .B(n10916), .S0(n4849), .Y(
        \D_cache/n1273 ) );
  MX2XL U10778 ( .A(\D_cache/cache[2][65] ), .B(n10916), .S0(n4805), .Y(
        \D_cache/n1274 ) );
  MX2XL U10779 ( .A(\D_cache/cache[1][65] ), .B(n10916), .S0(n4782), .Y(
        \D_cache/n1275 ) );
  MX2XL U10780 ( .A(\D_cache/cache[0][65] ), .B(n10916), .S0(n4736), .Y(
        \D_cache/n1276 ) );
  MX2XL U10781 ( .A(\D_cache/cache[3][64] ), .B(n10964), .S0(n4855), .Y(
        \D_cache/n1281 ) );
  MX2XL U10782 ( .A(\D_cache/cache[2][64] ), .B(n10964), .S0(n4802), .Y(
        \D_cache/n1282 ) );
  MX2XL U10783 ( .A(\D_cache/cache[1][64] ), .B(n10964), .S0(n4786), .Y(
        \D_cache/n1283 ) );
  MX2XL U10784 ( .A(\D_cache/cache[0][64] ), .B(n10964), .S0(n4736), .Y(
        \D_cache/n1284 ) );
  MX2XL U10785 ( .A(\D_cache/cache[6][101] ), .B(n10986), .S0(n4965), .Y(
        \D_cache/n982 ) );
  MX2XL U10786 ( .A(\D_cache/cache[5][101] ), .B(n10986), .S0(n4944), .Y(
        \D_cache/n983 ) );
  MX2XL U10787 ( .A(\D_cache/cache[4][101] ), .B(n10986), .S0(n4901), .Y(
        \D_cache/n984 ) );
  MX2XL U10788 ( .A(\D_cache/cache[3][101] ), .B(n10986), .S0(n4855), .Y(
        \D_cache/n985 ) );
  MX2XL U10789 ( .A(\D_cache/cache[2][101] ), .B(n10986), .S0(n4803), .Y(
        \D_cache/n986 ) );
  MX2XL U10790 ( .A(\D_cache/cache[1][101] ), .B(n10986), .S0(n4786), .Y(
        \D_cache/n987 ) );
  MX2XL U10791 ( .A(\D_cache/cache[6][100] ), .B(n10974), .S0(n4965), .Y(
        \D_cache/n990 ) );
  MX2XL U10792 ( .A(\D_cache/cache[5][100] ), .B(n10974), .S0(n4944), .Y(
        \D_cache/n991 ) );
  MX2XL U10793 ( .A(\D_cache/cache[4][100] ), .B(n10974), .S0(n4901), .Y(
        \D_cache/n992 ) );
  MX2XL U10794 ( .A(\D_cache/cache[3][100] ), .B(n10974), .S0(n4855), .Y(
        \D_cache/n993 ) );
  MX2XL U10795 ( .A(\D_cache/cache[2][100] ), .B(n10974), .S0(n4803), .Y(
        \D_cache/n994 ) );
  MX2XL U10796 ( .A(\D_cache/cache[1][100] ), .B(n10974), .S0(n4786), .Y(
        \D_cache/n995 ) );
  MX2XL U10797 ( .A(\D_cache/cache[0][100] ), .B(n10974), .S0(n4738), .Y(
        \D_cache/n996 ) );
  MX2XL U10798 ( .A(\D_cache/cache[6][99] ), .B(n10922), .S0(n4964), .Y(
        \D_cache/n998 ) );
  MX2XL U10799 ( .A(\D_cache/cache[5][99] ), .B(n10922), .S0(n4943), .Y(
        \D_cache/n999 ) );
  MX2XL U10800 ( .A(\D_cache/cache[4][99] ), .B(n10922), .S0(n4900), .Y(
        \D_cache/n1000 ) );
  MX2XL U10801 ( .A(\D_cache/cache[3][99] ), .B(n10922), .S0(n4854), .Y(
        \D_cache/n1001 ) );
  MX2XL U10802 ( .A(\D_cache/cache[2][99] ), .B(n10922), .S0(n4809), .Y(
        \D_cache/n1002 ) );
  MX2XL U10803 ( .A(\D_cache/cache[1][99] ), .B(n10922), .S0(n4780), .Y(
        \D_cache/n1003 ) );
  MX2XL U10804 ( .A(\D_cache/cache[0][99] ), .B(n10922), .S0(n4741), .Y(
        \D_cache/n1004 ) );
  MX2XL U10805 ( .A(\D_cache/cache[6][98] ), .B(n10936), .S0(n4964), .Y(
        \D_cache/n1006 ) );
  MX2XL U10806 ( .A(\D_cache/cache[5][98] ), .B(n10936), .S0(n4943), .Y(
        \D_cache/n1007 ) );
  MX2XL U10807 ( .A(\D_cache/cache[4][98] ), .B(n10936), .S0(n4900), .Y(
        \D_cache/n1008 ) );
  MX2XL U10808 ( .A(\D_cache/cache[3][98] ), .B(n10936), .S0(n4854), .Y(
        \D_cache/n1009 ) );
  MX2XL U10809 ( .A(\D_cache/cache[2][98] ), .B(n10936), .S0(n4809), .Y(
        \D_cache/n1010 ) );
  MX2XL U10810 ( .A(\D_cache/cache[1][98] ), .B(n10936), .S0(n4783), .Y(
        \D_cache/n1011 ) );
  MX2XL U10811 ( .A(\D_cache/cache[0][98] ), .B(n10936), .S0(n4741), .Y(
        \D_cache/n1012 ) );
  MX2XL U10812 ( .A(\D_cache/cache[6][97] ), .B(n190), .S0(n4958), .Y(
        \D_cache/n1014 ) );
  MX2XL U10813 ( .A(\D_cache/cache[5][97] ), .B(n190), .S0(n4938), .Y(
        \D_cache/n1015 ) );
  MX2XL U10814 ( .A(\D_cache/cache[4][97] ), .B(n190), .S0(n4892), .Y(
        \D_cache/n1016 ) );
  MX2XL U10815 ( .A(\D_cache/cache[3][97] ), .B(n190), .S0(n4850), .Y(
        \D_cache/n1017 ) );
  MX2XL U10816 ( .A(\D_cache/cache[2][97] ), .B(n190), .S0(n4806), .Y(
        \D_cache/n1018 ) );
  MX2XL U10817 ( .A(\D_cache/cache[1][97] ), .B(n190), .S0(n4781), .Y(
        \D_cache/n1019 ) );
  MX2XL U10818 ( .A(\D_cache/cache[0][97] ), .B(n190), .S0(n4736), .Y(
        \D_cache/n1020 ) );
  MX2XL U10819 ( .A(\D_cache/cache[6][96] ), .B(n10961), .S0(n4956), .Y(
        \D_cache/n1022 ) );
  MX2XL U10820 ( .A(\D_cache/cache[5][96] ), .B(n10961), .S0(n4936), .Y(
        \D_cache/n1023 ) );
  MX2XL U10821 ( .A(\D_cache/cache[4][96] ), .B(n10961), .S0(n4892), .Y(
        \D_cache/n1024 ) );
  MX2XL U10822 ( .A(\D_cache/cache[3][96] ), .B(n10961), .S0(n4846), .Y(
        \D_cache/n1025 ) );
  MX2XL U10823 ( .A(\D_cache/cache[2][96] ), .B(n10961), .S0(n4801), .Y(
        \D_cache/n1026 ) );
  MX2XL U10824 ( .A(\D_cache/cache[1][96] ), .B(n10961), .S0(n4778), .Y(
        \D_cache/n1027 ) );
  MX2XL U10825 ( .A(\D_cache/cache[0][96] ), .B(n10961), .S0(n4732), .Y(
        \D_cache/n1028 ) );
  OA22X1 U10826 ( .A0(\i_MIPS/Register/register[17][6] ), .A1(net112254), .B0(
        \i_MIPS/Register/register[25][6] ), .B1(n147), .Y(n6996) );
  OA22X1 U10827 ( .A0(\i_MIPS/Register/register[17][4] ), .A1(net112258), .B0(
        \i_MIPS/Register/register[25][4] ), .B1(n148), .Y(n6871) );
  OA22X1 U10828 ( .A0(\i_MIPS/Register/register[17][13] ), .A1(net112260), 
        .B0(\i_MIPS/Register/register[25][13] ), .B1(n147), .Y(n7730) );
  OA22X1 U10829 ( .A0(\i_MIPS/Register/register[17][14] ), .A1(net112260), 
        .B0(\i_MIPS/Register/register[25][14] ), .B1(n150), .Y(n7637) );
  OA22X1 U10830 ( .A0(\i_MIPS/Register/register[17][11] ), .A1(net112258), 
        .B0(\i_MIPS/Register/register[25][11] ), .B1(n148), .Y(n7256) );
  OA22X1 U10831 ( .A0(\i_MIPS/Register/register[17][9] ), .A1(net112260), .B0(
        \i_MIPS/Register/register[25][9] ), .B1(n148), .Y(n8675) );
  OA22X1 U10832 ( .A0(\i_MIPS/Register/register[17][23] ), .A1(net112260), 
        .B0(\i_MIPS/Register/register[25][23] ), .B1(n151), .Y(n8840) );
  OA22X1 U10833 ( .A0(\i_MIPS/Register/register[17][18] ), .A1(net112260), 
        .B0(\i_MIPS/Register/register[25][18] ), .B1(n150), .Y(n8777) );
  OA22X1 U10834 ( .A0(\i_MIPS/Register/register[17][20] ), .A1(net112260), 
        .B0(\i_MIPS/Register/register[25][20] ), .B1(n151), .Y(n9234) );
  OA22X1 U10835 ( .A0(\i_MIPS/Register/register[17][25] ), .A1(net112254), 
        .B0(\i_MIPS/Register/register[25][25] ), .B1(n148), .Y(n9032) );
  OA22X1 U10836 ( .A0(\i_MIPS/Register/register[17][21] ), .A1(net112260), 
        .B0(\i_MIPS/Register/register[25][21] ), .B1(n150), .Y(n9129) );
  OA22X1 U10837 ( .A0(\i_MIPS/Register/register[17][24] ), .A1(net112260), 
        .B0(\i_MIPS/Register/register[25][24] ), .B1(n150), .Y(n8288) );
  MXI2X1 U10838 ( .A(\i_MIPS/PHT_2/n8 ), .B(\i_MIPS/PHT_2/n7 ), .S0(n4529), 
        .Y(\i_MIPS/PHT_2/n48 ) );
  MX2XL U10839 ( .A(\i_MIPS/EX_MEM[5] ), .B(n3875), .S0(n223), .Y(
        \i_MIPS/n469 ) );
  MX2XL U10840 ( .A(\i_MIPS/ID_EX[66] ), .B(n4615), .S0(n211), .Y(
        \i_MIPS/n387 ) );
  CLKINVX1 U10841 ( .A(\i_MIPS/n309 ), .Y(n10952) );
  CLKMX2X2 U10842 ( .A(\D_cache/cache[7][153] ), .B(n10927), .S0(n5008), .Y(
        \D_cache/n565 ) );
  CLKMX2X2 U10843 ( .A(\D_cache/cache[6][153] ), .B(n10927), .S0(n4964), .Y(
        \D_cache/n566 ) );
  CLKMX2X2 U10844 ( .A(\D_cache/cache[5][153] ), .B(n10927), .S0(n4943), .Y(
        \D_cache/n567 ) );
  CLKMX2X2 U10845 ( .A(\D_cache/cache[4][153] ), .B(n10927), .S0(n4900), .Y(
        \D_cache/n568 ) );
  CLKMX2X2 U10846 ( .A(\D_cache/cache[3][153] ), .B(n10927), .S0(n4854), .Y(
        \D_cache/n569 ) );
  CLKMX2X2 U10847 ( .A(\D_cache/cache[2][153] ), .B(n10927), .S0(n4809), .Y(
        \D_cache/n570 ) );
  CLKMX2X2 U10848 ( .A(\D_cache/cache[1][153] ), .B(n10927), .S0(n4780), .Y(
        \D_cache/n571 ) );
  CLKMX2X2 U10849 ( .A(\D_cache/cache[0][153] ), .B(n10927), .S0(n4735), .Y(
        \D_cache/n572 ) );
  MX2XL U10850 ( .A(\i_MIPS/ID_EX[68] ), .B(n10318), .S0(n204), .Y(
        \i_MIPS/n383 ) );
  MXI2XL U10851 ( .A(n4534), .B(n9885), .S0(n217), .Y(\i_MIPS/n475 ) );
  MXI2XL U10852 ( .A(n4542), .B(n259), .S0(n217), .Y(\i_MIPS/n473 ) );
  MX2XL U10853 ( .A(\i_MIPS/Reg_W[1] ), .B(n9884), .S0(n210), .Y(\i_MIPS/n476 ) );
  MX2XL U10854 ( .A(n3603), .B(n3918), .S0(n222), .Y(\i_MIPS/n427 ) );
  MX2XL U10855 ( .A(\i_MIPS/ID_EX[42] ), .B(n3780), .S0(n213), .Y(
        \i_MIPS/n435 ) );
  MX2XL U10856 ( .A(\i_MIPS/Reg_W[0] ), .B(n9886), .S0(n205), .Y(\i_MIPS/n477 ) );
  MX2XL U10857 ( .A(\D_cache/cache[6][149] ), .B(n11023), .S0(n4962), .Y(
        \D_cache/n598 ) );
  MX2XL U10858 ( .A(\D_cache/cache[5][149] ), .B(n11023), .S0(n4942), .Y(
        \D_cache/n599 ) );
  MX2XL U10859 ( .A(\D_cache/cache[4][149] ), .B(n11023), .S0(n4898), .Y(
        \D_cache/n600 ) );
  MX2XL U10860 ( .A(\D_cache/cache[3][149] ), .B(n11023), .S0(n4852), .Y(
        \D_cache/n601 ) );
  MX2XL U10861 ( .A(\D_cache/cache[2][149] ), .B(n11023), .S0(n4803), .Y(
        \D_cache/n602 ) );
  MX2XL U10862 ( .A(\D_cache/cache[1][149] ), .B(n11023), .S0(n4785), .Y(
        \D_cache/n603 ) );
  MX2XL U10863 ( .A(\D_cache/cache[0][149] ), .B(n11023), .S0(n4739), .Y(
        \D_cache/n604 ) );
  MX2XL U10864 ( .A(\D_cache/cache[6][147] ), .B(n11022), .S0(n4962), .Y(
        \D_cache/n614 ) );
  MX2XL U10865 ( .A(\D_cache/cache[5][147] ), .B(n11022), .S0(n4941), .Y(
        \D_cache/n615 ) );
  MX2XL U10866 ( .A(\D_cache/cache[4][147] ), .B(n11022), .S0(n4898), .Y(
        \D_cache/n616 ) );
  MX2XL U10867 ( .A(\D_cache/cache[3][147] ), .B(n11022), .S0(n4852), .Y(
        \D_cache/n617 ) );
  MX2XL U10868 ( .A(\D_cache/cache[2][147] ), .B(n11022), .S0(n4805), .Y(
        \D_cache/n618 ) );
  MX2XL U10869 ( .A(\D_cache/cache[1][147] ), .B(n11022), .S0(n4784), .Y(
        \D_cache/n619 ) );
  MX2XL U10870 ( .A(\D_cache/cache[0][147] ), .B(n11022), .S0(n4735), .Y(
        \D_cache/n620 ) );
  MX2XL U10871 ( .A(\D_cache/cache[6][128] ), .B(n11019), .S0(n4962), .Y(
        \D_cache/n766 ) );
  MX2XL U10872 ( .A(\D_cache/cache[5][128] ), .B(n11019), .S0(n4942), .Y(
        \D_cache/n767 ) );
  MX2XL U10873 ( .A(\D_cache/cache[4][128] ), .B(n11019), .S0(n4898), .Y(
        \D_cache/n768 ) );
  MX2XL U10874 ( .A(\D_cache/cache[3][128] ), .B(n11019), .S0(n4852), .Y(
        \D_cache/n769 ) );
  MX2XL U10875 ( .A(\D_cache/cache[2][128] ), .B(n11019), .S0(n4806), .Y(
        \D_cache/n770 ) );
  MX2XL U10876 ( .A(\D_cache/cache[1][128] ), .B(n11019), .S0(n4785), .Y(
        \D_cache/n771 ) );
  MX2XL U10877 ( .A(\D_cache/cache[0][128] ), .B(n11019), .S0(n4738), .Y(
        \D_cache/n772 ) );
  MX2XL U10878 ( .A(\i_MIPS/Reg_W[3] ), .B(n9883), .S0(n219), .Y(\i_MIPS/n474 ) );
  MX2XL U10879 ( .A(\D_cache/cache[6][143] ), .B(n11034), .S0(n4963), .Y(
        \D_cache/n646 ) );
  MX2XL U10880 ( .A(\D_cache/cache[5][143] ), .B(n11034), .S0(n4943), .Y(
        \D_cache/n647 ) );
  MX2XL U10881 ( .A(\D_cache/cache[4][143] ), .B(n11034), .S0(n4899), .Y(
        \D_cache/n648 ) );
  MX2XL U10882 ( .A(\D_cache/cache[3][143] ), .B(n11034), .S0(n4853), .Y(
        \D_cache/n649 ) );
  MX2XL U10883 ( .A(\D_cache/cache[2][143] ), .B(n11034), .S0(n4808), .Y(
        \D_cache/n650 ) );
  MX2XL U10884 ( .A(\D_cache/cache[1][143] ), .B(n11034), .S0(n4781), .Y(
        \D_cache/n651 ) );
  MX2XL U10885 ( .A(\D_cache/cache[0][143] ), .B(n11034), .S0(n4740), .Y(
        \D_cache/n652 ) );
  MX2XL U10886 ( .A(\D_cache/cache[6][145] ), .B(n11028), .S0(n4963), .Y(
        \D_cache/n630 ) );
  MX2XL U10887 ( .A(\D_cache/cache[5][145] ), .B(n11028), .S0(n4944), .Y(
        \D_cache/n631 ) );
  MX2XL U10888 ( .A(\D_cache/cache[4][145] ), .B(n11028), .S0(n4899), .Y(
        \D_cache/n632 ) );
  MX2XL U10889 ( .A(\D_cache/cache[3][145] ), .B(n11028), .S0(n4853), .Y(
        \D_cache/n633 ) );
  MX2XL U10890 ( .A(\D_cache/cache[2][145] ), .B(n11028), .S0(n4808), .Y(
        \D_cache/n634 ) );
  MX2XL U10891 ( .A(\D_cache/cache[1][145] ), .B(n11028), .S0(n4778), .Y(
        \D_cache/n635 ) );
  MX2XL U10892 ( .A(\D_cache/cache[0][145] ), .B(n11028), .S0(n4740), .Y(
        \D_cache/n636 ) );
  MX2XL U10893 ( .A(\D_cache/cache[6][130] ), .B(n3834), .S0(n4963), .Y(
        \D_cache/n750 ) );
  MX2XL U10894 ( .A(\D_cache/cache[5][130] ), .B(n3834), .S0(n4940), .Y(
        \D_cache/n751 ) );
  MX2XL U10895 ( .A(\D_cache/cache[4][130] ), .B(n3834), .S0(n4899), .Y(
        \D_cache/n752 ) );
  MX2XL U10896 ( .A(\D_cache/cache[3][130] ), .B(n3834), .S0(n4853), .Y(
        \D_cache/n753 ) );
  MX2XL U10897 ( .A(\D_cache/cache[1][130] ), .B(n3834), .S0(n4786), .Y(
        \D_cache/n755 ) );
  MX2XL U10898 ( .A(\D_cache/cache[0][130] ), .B(n3834), .S0(n4740), .Y(
        \D_cache/n756 ) );
  MX2XL U10899 ( .A(\D_cache/cache[6][136] ), .B(n11020), .S0(n4962), .Y(
        \D_cache/n702 ) );
  MX2XL U10900 ( .A(\D_cache/cache[5][136] ), .B(n11020), .S0(n4941), .Y(
        \D_cache/n703 ) );
  MX2XL U10901 ( .A(\D_cache/cache[4][136] ), .B(n11020), .S0(n4898), .Y(
        \D_cache/n704 ) );
  MX2XL U10902 ( .A(\D_cache/cache[3][136] ), .B(n11020), .S0(n4852), .Y(
        \D_cache/n705 ) );
  MX2XL U10903 ( .A(\D_cache/cache[2][136] ), .B(n11020), .S0(n4804), .Y(
        \D_cache/n706 ) );
  MX2XL U10904 ( .A(\D_cache/cache[1][136] ), .B(n11020), .S0(n4784), .Y(
        \D_cache/n707 ) );
  MX2XL U10905 ( .A(\D_cache/cache[0][136] ), .B(n11020), .S0(n4736), .Y(
        \D_cache/n708 ) );
  MX2XL U10906 ( .A(\D_cache/cache[5][142] ), .B(n11040), .S0(n4939), .Y(
        \D_cache/n655 ) );
  MX2XL U10907 ( .A(\D_cache/cache[4][142] ), .B(n11040), .S0(n4892), .Y(
        \D_cache/n656 ) );
  MX2XL U10908 ( .A(\D_cache/cache[6][129] ), .B(n11038), .S0(n4963), .Y(
        \D_cache/n758 ) );
  MX2XL U10909 ( .A(\D_cache/cache[5][129] ), .B(n11038), .S0(n4938), .Y(
        \D_cache/n759 ) );
  MX2XL U10910 ( .A(\D_cache/cache[4][129] ), .B(n11038), .S0(n4899), .Y(
        \D_cache/n760 ) );
  MX2XL U10911 ( .A(\D_cache/cache[3][129] ), .B(n11038), .S0(n4853), .Y(
        \D_cache/n761 ) );
  MX2XL U10912 ( .A(\D_cache/cache[2][129] ), .B(n11038), .S0(n4808), .Y(
        \D_cache/n762 ) );
  MX2XL U10913 ( .A(\D_cache/cache[1][129] ), .B(n11038), .S0(n4778), .Y(
        \D_cache/n763 ) );
  MX2XL U10914 ( .A(\D_cache/cache[0][129] ), .B(n11038), .S0(n4740), .Y(
        \D_cache/n764 ) );
  MX2XL U10915 ( .A(\D_cache/cache[6][132] ), .B(n11027), .S0(n4963), .Y(
        \D_cache/n734 ) );
  MX2XL U10916 ( .A(\D_cache/cache[5][132] ), .B(n11027), .S0(n4943), .Y(
        \D_cache/n735 ) );
  MX2XL U10917 ( .A(\D_cache/cache[4][132] ), .B(n11027), .S0(n4899), .Y(
        \D_cache/n736 ) );
  MX2XL U10918 ( .A(\D_cache/cache[3][132] ), .B(n11027), .S0(n4853), .Y(
        \D_cache/n737 ) );
  MX2XL U10919 ( .A(\D_cache/cache[2][132] ), .B(n11027), .S0(n4808), .Y(
        \D_cache/n738 ) );
  MX2XL U10920 ( .A(\D_cache/cache[1][132] ), .B(n11027), .S0(n4783), .Y(
        \D_cache/n739 ) );
  MX2XL U10921 ( .A(\D_cache/cache[0][132] ), .B(n11027), .S0(n4740), .Y(
        \D_cache/n740 ) );
  MX2XL U10922 ( .A(\D_cache/cache[6][141] ), .B(n11035), .S0(n4963), .Y(
        \D_cache/n662 ) );
  MX2XL U10923 ( .A(\D_cache/cache[5][141] ), .B(n11035), .S0(n4944), .Y(
        \D_cache/n663 ) );
  MX2XL U10924 ( .A(\D_cache/cache[4][141] ), .B(n11035), .S0(n4899), .Y(
        \D_cache/n664 ) );
  MX2XL U10925 ( .A(\D_cache/cache[3][141] ), .B(n11035), .S0(n4853), .Y(
        \D_cache/n665 ) );
  MX2XL U10926 ( .A(\D_cache/cache[1][141] ), .B(n11035), .S0(n4781), .Y(
        \D_cache/n667 ) );
  MX2XL U10927 ( .A(\D_cache/cache[0][141] ), .B(n11035), .S0(n4740), .Y(
        \D_cache/n668 ) );
  MX2XL U10928 ( .A(\D_cache/cache[6][138] ), .B(n11032), .S0(n4963), .Y(
        \D_cache/n686 ) );
  MX2XL U10929 ( .A(\D_cache/cache[5][138] ), .B(n11032), .S0(n4940), .Y(
        \D_cache/n687 ) );
  MX2XL U10930 ( .A(\D_cache/cache[4][138] ), .B(n11032), .S0(n4899), .Y(
        \D_cache/n688 ) );
  MX2XL U10931 ( .A(\D_cache/cache[3][138] ), .B(n11032), .S0(n4853), .Y(
        \D_cache/n689 ) );
  MX2XL U10932 ( .A(\D_cache/cache[2][138] ), .B(n11032), .S0(n4808), .Y(
        \D_cache/n690 ) );
  MX2XL U10933 ( .A(\D_cache/cache[1][138] ), .B(n11032), .S0(n4779), .Y(
        \D_cache/n691 ) );
  MX2XL U10934 ( .A(\D_cache/cache[0][138] ), .B(n11032), .S0(n4740), .Y(
        \D_cache/n692 ) );
  MX2XL U10935 ( .A(\D_cache/cache[6][134] ), .B(n11030), .S0(n4963), .Y(
        \D_cache/n718 ) );
  MX2XL U10936 ( .A(\D_cache/cache[5][134] ), .B(n11030), .S0(n4938), .Y(
        \D_cache/n719 ) );
  MX2XL U10937 ( .A(\D_cache/cache[4][134] ), .B(n11030), .S0(n4899), .Y(
        \D_cache/n720 ) );
  MX2XL U10938 ( .A(\D_cache/cache[3][134] ), .B(n11030), .S0(n4853), .Y(
        \D_cache/n721 ) );
  MX2XL U10939 ( .A(\D_cache/cache[2][134] ), .B(n11030), .S0(n4808), .Y(
        \D_cache/n722 ) );
  MX2XL U10940 ( .A(\D_cache/cache[1][134] ), .B(n11030), .S0(n4786), .Y(
        \D_cache/n723 ) );
  MX2XL U10941 ( .A(\D_cache/cache[0][134] ), .B(n11030), .S0(n4740), .Y(
        \D_cache/n724 ) );
  MX2XL U10942 ( .A(\D_cache/cache[6][133] ), .B(n11031), .S0(n4963), .Y(
        \D_cache/n726 ) );
  MX2XL U10943 ( .A(\D_cache/cache[5][133] ), .B(n11031), .S0(n4943), .Y(
        \D_cache/n727 ) );
  MX2XL U10944 ( .A(\D_cache/cache[4][133] ), .B(n11031), .S0(n4899), .Y(
        \D_cache/n728 ) );
  MX2XL U10945 ( .A(\D_cache/cache[3][133] ), .B(n11031), .S0(n4853), .Y(
        \D_cache/n729 ) );
  MX2XL U10946 ( .A(\D_cache/cache[2][133] ), .B(n11031), .S0(n4808), .Y(
        \D_cache/n730 ) );
  MX2XL U10947 ( .A(\D_cache/cache[1][133] ), .B(n11031), .S0(n4780), .Y(
        \D_cache/n731 ) );
  MX2XL U10948 ( .A(\D_cache/cache[0][133] ), .B(n11031), .S0(n4740), .Y(
        \D_cache/n732 ) );
  MX2XL U10949 ( .A(\D_cache/cache[6][131] ), .B(n11037), .S0(n4963), .Y(
        \D_cache/n742 ) );
  MX2XL U10950 ( .A(\D_cache/cache[5][131] ), .B(n11037), .S0(n4937), .Y(
        \D_cache/n743 ) );
  MX2XL U10951 ( .A(\D_cache/cache[4][131] ), .B(n11037), .S0(n4899), .Y(
        \D_cache/n744 ) );
  MX2XL U10952 ( .A(\D_cache/cache[3][131] ), .B(n11037), .S0(n4853), .Y(
        \D_cache/n745 ) );
  MX2XL U10953 ( .A(\D_cache/cache[2][131] ), .B(n11037), .S0(n4808), .Y(
        \D_cache/n746 ) );
  MX2XL U10954 ( .A(\D_cache/cache[1][131] ), .B(n11037), .S0(n4781), .Y(
        \D_cache/n747 ) );
  MX2XL U10955 ( .A(\D_cache/cache[0][131] ), .B(n11037), .S0(n4740), .Y(
        \D_cache/n748 ) );
  MX2XL U10956 ( .A(\D_cache/cache[7][152] ), .B(n11018), .S0(n5006), .Y(
        \D_cache/n573 ) );
  MX2XL U10957 ( .A(\D_cache/cache[6][152] ), .B(n11018), .S0(n4962), .Y(
        \D_cache/n574 ) );
  MX2XL U10958 ( .A(\D_cache/cache[5][152] ), .B(n11018), .S0(n4942), .Y(
        \D_cache/n575 ) );
  MX2XL U10959 ( .A(\D_cache/cache[4][152] ), .B(n11018), .S0(n4898), .Y(
        \D_cache/n576 ) );
  MX2XL U10960 ( .A(\D_cache/cache[3][152] ), .B(n11018), .S0(n4852), .Y(
        \D_cache/n577 ) );
  MX2XL U10961 ( .A(\D_cache/cache[2][152] ), .B(n11018), .S0(n4809), .Y(
        \D_cache/n578 ) );
  MX2XL U10962 ( .A(\D_cache/cache[1][152] ), .B(n11018), .S0(n4785), .Y(
        \D_cache/n579 ) );
  MX2XL U10963 ( .A(\D_cache/cache[0][152] ), .B(n11018), .S0(n4732), .Y(
        \D_cache/n580 ) );
  MX2XL U10964 ( .A(\D_cache/cache[6][151] ), .B(n11021), .S0(n4962), .Y(
        \D_cache/n582 ) );
  MX2XL U10965 ( .A(\D_cache/cache[5][151] ), .B(n11021), .S0(n4942), .Y(
        \D_cache/n583 ) );
  MX2XL U10966 ( .A(\D_cache/cache[4][151] ), .B(n11021), .S0(n4898), .Y(
        \D_cache/n584 ) );
  MX2XL U10967 ( .A(\D_cache/cache[3][151] ), .B(n11021), .S0(n4852), .Y(
        \D_cache/n585 ) );
  MX2XL U10968 ( .A(\D_cache/cache[2][151] ), .B(n11021), .S0(n4801), .Y(
        \D_cache/n586 ) );
  MX2XL U10969 ( .A(\D_cache/cache[1][151] ), .B(n11021), .S0(n4784), .Y(
        \D_cache/n587 ) );
  MX2XL U10970 ( .A(\D_cache/cache[0][151] ), .B(n11021), .S0(n4739), .Y(
        \D_cache/n588 ) );
  MX2XL U10971 ( .A(\D_cache/cache[6][148] ), .B(n11026), .S0(n4961), .Y(
        \D_cache/n606 ) );
  MX2XL U10972 ( .A(\D_cache/cache[5][148] ), .B(n11026), .S0(n4941), .Y(
        \D_cache/n607 ) );
  MX2XL U10973 ( .A(\D_cache/cache[4][148] ), .B(n11026), .S0(n4897), .Y(
        \D_cache/n608 ) );
  MX2XL U10974 ( .A(\D_cache/cache[3][148] ), .B(n11026), .S0(n4851), .Y(
        \D_cache/n609 ) );
  MX2XL U10975 ( .A(\D_cache/cache[2][148] ), .B(n11026), .S0(n4807), .Y(
        \D_cache/n610 ) );
  MX2XL U10976 ( .A(\D_cache/cache[1][148] ), .B(n11026), .S0(n4785), .Y(
        \D_cache/n611 ) );
  MX2XL U10977 ( .A(\D_cache/cache[0][148] ), .B(n11026), .S0(n4739), .Y(
        \D_cache/n612 ) );
  MX2XL U10978 ( .A(\I_cache/cache[7][128] ), .B(n11151), .S0(n5321), .Y(
        n11756) );
  MX2XL U10979 ( .A(\I_cache/cache[7][151] ), .B(n11150), .S0(n5316), .Y(
        n11572) );
  MX2XL U10980 ( .A(\I_cache/cache[6][151] ), .B(n11150), .S0(n5363), .Y(
        n11573) );
  MX2XL U10981 ( .A(\I_cache/cache[7][150] ), .B(n11138), .S0(n5320), .Y(
        n11580) );
  MX2XL U10982 ( .A(\I_cache/cache[6][150] ), .B(n11138), .S0(n5365), .Y(
        n11581) );
  MX2XL U10983 ( .A(\I_cache/cache[7][149] ), .B(n11144), .S0(n5320), .Y(
        n11588) );
  MX2XL U10984 ( .A(\I_cache/cache[6][149] ), .B(n11144), .S0(n5363), .Y(
        n11589) );
  MX2XL U10985 ( .A(\I_cache/cache[7][148] ), .B(n11146), .S0(n5320), .Y(
        n11596) );
  MX2XL U10986 ( .A(\I_cache/cache[6][148] ), .B(n11146), .S0(n5358), .Y(
        n11597) );
  MX2XL U10987 ( .A(\I_cache/cache[7][147] ), .B(n11145), .S0(n5320), .Y(
        n11604) );
  MX2XL U10988 ( .A(\I_cache/cache[6][147] ), .B(n11145), .S0(n5365), .Y(
        n11605) );
  MX2XL U10989 ( .A(\I_cache/cache[7][146] ), .B(n11137), .S0(n5322), .Y(
        n11612) );
  MX2XL U10990 ( .A(\I_cache/cache[6][146] ), .B(n11137), .S0(n5365), .Y(
        n11613) );
  MX2XL U10991 ( .A(\I_cache/cache[7][145] ), .B(n11139), .S0(n5320), .Y(
        n11620) );
  MX2XL U10992 ( .A(\I_cache/cache[6][145] ), .B(n11139), .S0(n5366), .Y(
        n11621) );
  MX2XL U10993 ( .A(\I_cache/cache[7][144] ), .B(n11154), .S0(n5321), .Y(
        n11628) );
  MX2XL U10994 ( .A(\I_cache/cache[6][144] ), .B(n11154), .S0(n5365), .Y(
        n11629) );
  MX2XL U10995 ( .A(\I_cache/cache[7][143] ), .B(n11133), .S0(n5315), .Y(
        n11636) );
  MX2XL U10996 ( .A(\I_cache/cache[6][143] ), .B(n11133), .S0(n5364), .Y(
        n11637) );
  MX2XL U10997 ( .A(\I_cache/cache[7][142] ), .B(n11131), .S0(n5316), .Y(
        n11644) );
  MX2XL U10998 ( .A(\I_cache/cache[6][142] ), .B(n11131), .S0(n5362), .Y(
        n11645) );
  MX2XL U10999 ( .A(\I_cache/cache[7][141] ), .B(n11132), .S0(n5314), .Y(
        n11652) );
  MX2XL U11000 ( .A(\I_cache/cache[6][141] ), .B(n11132), .S0(n5361), .Y(
        n11653) );
  MX2XL U11001 ( .A(\I_cache/cache[7][140] ), .B(n11156), .S0(n5321), .Y(
        n11660) );
  MX2XL U11002 ( .A(\I_cache/cache[6][140] ), .B(n11156), .S0(n5363), .Y(
        n11661) );
  MX2XL U11003 ( .A(\I_cache/cache[7][139] ), .B(n11153), .S0(n5321), .Y(
        n11668) );
  MX2XL U11004 ( .A(\I_cache/cache[6][139] ), .B(n11153), .S0(n5360), .Y(
        n11669) );
  MX2XL U11005 ( .A(\I_cache/cache[7][138] ), .B(n11140), .S0(n5320), .Y(
        n11676) );
  MX2XL U11006 ( .A(\I_cache/cache[6][138] ), .B(n11140), .S0(n5358), .Y(
        n11677) );
  MX2XL U11007 ( .A(\I_cache/cache[7][137] ), .B(n11147), .S0(n5320), .Y(
        n11684) );
  MX2XL U11008 ( .A(\I_cache/cache[6][137] ), .B(n11147), .S0(n5358), .Y(
        n11685) );
  MX2XL U11009 ( .A(\I_cache/cache[7][136] ), .B(n11149), .S0(n5320), .Y(
        n11692) );
  MX2XL U11010 ( .A(\I_cache/cache[6][136] ), .B(n11149), .S0(n5364), .Y(
        n11693) );
  MX2XL U11011 ( .A(\I_cache/cache[7][135] ), .B(n11148), .S0(n5320), .Y(
        n11700) );
  MX2XL U11012 ( .A(\I_cache/cache[6][135] ), .B(n11148), .S0(n5360), .Y(
        n11701) );
  MX2XL U11013 ( .A(\I_cache/cache[7][134] ), .B(n11142), .S0(n5320), .Y(
        n11708) );
  MX2XL U11014 ( .A(\I_cache/cache[6][134] ), .B(n11142), .S0(n5364), .Y(
        n11709) );
  MX2XL U11015 ( .A(\I_cache/cache[7][133] ), .B(n11141), .S0(n5320), .Y(
        n11716) );
  MX2XL U11016 ( .A(\I_cache/cache[6][133] ), .B(n11141), .S0(n5361), .Y(
        n11717) );
  MX2XL U11017 ( .A(\I_cache/cache[7][132] ), .B(n11143), .S0(n5320), .Y(
        n11724) );
  MX2XL U11018 ( .A(\I_cache/cache[6][132] ), .B(n11143), .S0(n5358), .Y(
        n11725) );
  MX2XL U11019 ( .A(\I_cache/cache[7][131] ), .B(n11135), .S0(n5317), .Y(
        n11732) );
  MX2XL U11020 ( .A(\I_cache/cache[6][131] ), .B(n11135), .S0(n5364), .Y(
        n11733) );
  MX2XL U11021 ( .A(\I_cache/cache[7][130] ), .B(n11136), .S0(n5320), .Y(
        n11740) );
  MX2XL U11022 ( .A(\I_cache/cache[6][130] ), .B(n11136), .S0(n5359), .Y(
        n11741) );
  MX2XL U11023 ( .A(\I_cache/cache[7][129] ), .B(n11134), .S0(n5315), .Y(
        n11748) );
  MX2XL U11024 ( .A(\I_cache/cache[6][129] ), .B(n11134), .S0(n5361), .Y(
        n11749) );
  MX2XL U11025 ( .A(\I_cache/cache[6][128] ), .B(n11151), .S0(n5362), .Y(
        n11757) );
  CLKMX2X2 U11026 ( .A(\I_cache/cache[7][127] ), .B(n164), .S0(n5317), .Y(
        n11764) );
  CLKMX2X2 U11027 ( .A(\I_cache/cache[6][127] ), .B(n164), .S0(n5364), .Y(
        n11765) );
  CLKMX2X2 U11028 ( .A(\I_cache/cache[5][127] ), .B(n164), .S0(n5231), .Y(
        n11766) );
  CLKMX2X2 U11029 ( .A(\I_cache/cache[4][127] ), .B(n164), .S0(n5271), .Y(
        n11767) );
  CLKMX2X2 U11030 ( .A(\I_cache/cache[3][127] ), .B(n164), .S0(n5138), .Y(
        n11768) );
  CLKMX2X2 U11031 ( .A(\I_cache/cache[2][127] ), .B(n164), .S0(n5184), .Y(
        n11769) );
  CLKMX2X2 U11032 ( .A(\I_cache/cache[1][127] ), .B(n164), .S0(n5053), .Y(
        n11770) );
  CLKMX2X2 U11033 ( .A(\I_cache/cache[0][127] ), .B(n164), .S0(n5094), .Y(
        n11771) );
  CLKMX2X2 U11034 ( .A(\I_cache/cache[6][126] ), .B(n6211), .S0(n5363), .Y(
        n11773) );
  CLKMX2X2 U11035 ( .A(\I_cache/cache[5][126] ), .B(n6211), .S0(n5225), .Y(
        n11774) );
  CLKMX2X2 U11036 ( .A(\I_cache/cache[4][126] ), .B(n6211), .S0(n5271), .Y(
        n11775) );
  CLKMX2X2 U11037 ( .A(\I_cache/cache[3][126] ), .B(n6211), .S0(n5138), .Y(
        n11776) );
  CLKMX2X2 U11038 ( .A(\I_cache/cache[1][126] ), .B(n6211), .S0(n5051), .Y(
        n11778) );
  CLKMX2X2 U11039 ( .A(\I_cache/cache[0][126] ), .B(n6211), .S0(n5094), .Y(
        n11779) );
  CLKMX2X2 U11040 ( .A(\I_cache/cache[7][125] ), .B(n6231), .S0(n5317), .Y(
        n11780) );
  CLKMX2X2 U11041 ( .A(\I_cache/cache[6][125] ), .B(n6231), .S0(n5365), .Y(
        n11781) );
  CLKMX2X2 U11042 ( .A(\I_cache/cache[5][125] ), .B(n6231), .S0(n5228), .Y(
        n11782) );
  CLKMX2X2 U11043 ( .A(\I_cache/cache[4][125] ), .B(n6231), .S0(n5271), .Y(
        n11783) );
  CLKMX2X2 U11044 ( .A(\I_cache/cache[3][125] ), .B(n6231), .S0(n5138), .Y(
        n11784) );
  CLKMX2X2 U11045 ( .A(\I_cache/cache[2][125] ), .B(n6231), .S0(n5184), .Y(
        n11785) );
  CLKMX2X2 U11046 ( .A(\I_cache/cache[1][125] ), .B(n6231), .S0(n5046), .Y(
        n11786) );
  CLKMX2X2 U11047 ( .A(\I_cache/cache[0][125] ), .B(n6231), .S0(n5094), .Y(
        n11787) );
  CLKMX2X2 U11048 ( .A(\I_cache/cache[7][124] ), .B(n157), .S0(n5316), .Y(
        n11788) );
  CLKMX2X2 U11049 ( .A(\I_cache/cache[6][124] ), .B(n157), .S0(n5364), .Y(
        n11789) );
  CLKMX2X2 U11050 ( .A(\I_cache/cache[5][124] ), .B(n157), .S0(n5227), .Y(
        n11790) );
  CLKMX2X2 U11051 ( .A(\I_cache/cache[4][124] ), .B(n157), .S0(n5270), .Y(
        n11791) );
  CLKMX2X2 U11052 ( .A(\I_cache/cache[3][124] ), .B(n157), .S0(n5137), .Y(
        n11792) );
  CLKMX2X2 U11053 ( .A(\I_cache/cache[2][124] ), .B(n157), .S0(n5183), .Y(
        n11793) );
  CLKMX2X2 U11054 ( .A(\I_cache/cache[1][124] ), .B(n157), .S0(n5050), .Y(
        n11794) );
  CLKMX2X2 U11055 ( .A(\I_cache/cache[0][124] ), .B(n157), .S0(n5093), .Y(
        n11795) );
  CLKMX2X2 U11056 ( .A(\I_cache/cache[7][123] ), .B(n11159), .S0(n5321), .Y(
        n11796) );
  CLKMX2X2 U11057 ( .A(\I_cache/cache[6][123] ), .B(n11159), .S0(n5362), .Y(
        n11797) );
  CLKMX2X2 U11058 ( .A(\I_cache/cache[5][123] ), .B(n11159), .S0(n5233), .Y(
        n11798) );
  CLKMX2X2 U11059 ( .A(\I_cache/cache[4][123] ), .B(n11159), .S0(n5276), .Y(
        n11799) );
  CLKMX2X2 U11060 ( .A(\I_cache/cache[3][123] ), .B(n11159), .S0(n5143), .Y(
        n11800) );
  CLKMX2X2 U11061 ( .A(\I_cache/cache[2][123] ), .B(n11159), .S0(n5189), .Y(
        n11801) );
  CLKMX2X2 U11062 ( .A(\I_cache/cache[1][123] ), .B(n11159), .S0(n5046), .Y(
        n11802) );
  CLKMX2X2 U11063 ( .A(\I_cache/cache[0][123] ), .B(n11159), .S0(n5098), .Y(
        n11803) );
  CLKMX2X2 U11064 ( .A(\I_cache/cache[7][122] ), .B(n9563), .S0(n5316), .Y(
        n11804) );
  CLKMX2X2 U11065 ( .A(\I_cache/cache[6][122] ), .B(n9563), .S0(n5366), .Y(
        n11805) );
  CLKMX2X2 U11066 ( .A(\I_cache/cache[5][122] ), .B(n9563), .S0(n5227), .Y(
        n11806) );
  CLKMX2X2 U11067 ( .A(\I_cache/cache[4][122] ), .B(n9563), .S0(n5270), .Y(
        n11807) );
  CLKMX2X2 U11068 ( .A(\I_cache/cache[3][122] ), .B(n9563), .S0(n5137), .Y(
        n11808) );
  CLKMX2X2 U11069 ( .A(\I_cache/cache[2][122] ), .B(n9563), .S0(n5183), .Y(
        n11809) );
  CLKMX2X2 U11070 ( .A(\I_cache/cache[1][122] ), .B(n9563), .S0(n5048), .Y(
        n11810) );
  CLKMX2X2 U11071 ( .A(\I_cache/cache[0][122] ), .B(n9563), .S0(n5091), .Y(
        n11811) );
  CLKMX2X2 U11072 ( .A(\I_cache/cache[7][121] ), .B(n9817), .S0(n5322), .Y(
        n11812) );
  CLKMX2X2 U11073 ( .A(\I_cache/cache[6][121] ), .B(n9817), .S0(n5361), .Y(
        n11813) );
  CLKMX2X2 U11074 ( .A(\I_cache/cache[5][121] ), .B(n9817), .S0(n5231), .Y(
        n11814) );
  CLKMX2X2 U11075 ( .A(\I_cache/cache[4][121] ), .B(n9817), .S0(n5274), .Y(
        n11815) );
  CLKMX2X2 U11076 ( .A(\I_cache/cache[3][121] ), .B(n9817), .S0(n5142), .Y(
        n11816) );
  CLKMX2X2 U11077 ( .A(\I_cache/cache[2][121] ), .B(n9817), .S0(n5188), .Y(
        n11817) );
  CLKMX2X2 U11078 ( .A(\I_cache/cache[1][121] ), .B(n9817), .S0(n5049), .Y(
        n11818) );
  CLKMX2X2 U11079 ( .A(\I_cache/cache[0][121] ), .B(n9817), .S0(n5096), .Y(
        n11819) );
  CLKMX2X2 U11080 ( .A(\I_cache/cache[7][120] ), .B(n9797), .S0(n5319), .Y(
        n11820) );
  CLKMX2X2 U11081 ( .A(\I_cache/cache[6][120] ), .B(n9797), .S0(n5366), .Y(
        n11821) );
  CLKMX2X2 U11082 ( .A(\I_cache/cache[5][120] ), .B(n9797), .S0(n5230), .Y(
        n11822) );
  CLKMX2X2 U11083 ( .A(\I_cache/cache[4][120] ), .B(n9797), .S0(n5273), .Y(
        n11823) );
  CLKMX2X2 U11084 ( .A(\I_cache/cache[3][120] ), .B(n9797), .S0(n5141), .Y(
        n11824) );
  CLKMX2X2 U11085 ( .A(\I_cache/cache[2][120] ), .B(n9797), .S0(n5187), .Y(
        n11825) );
  CLKMX2X2 U11086 ( .A(\I_cache/cache[1][120] ), .B(n9797), .S0(n5048), .Y(
        n11826) );
  CLKMX2X2 U11087 ( .A(\I_cache/cache[0][120] ), .B(n9797), .S0(n5095), .Y(
        n11827) );
  CLKMX2X2 U11088 ( .A(\I_cache/cache[7][119] ), .B(n9837), .S0(n5320), .Y(
        n11828) );
  CLKMX2X2 U11089 ( .A(\I_cache/cache[6][119] ), .B(n9837), .S0(n5361), .Y(
        n11829) );
  CLKMX2X2 U11090 ( .A(\I_cache/cache[5][119] ), .B(n9837), .S0(n5231), .Y(
        n11830) );
  CLKMX2X2 U11091 ( .A(\I_cache/cache[4][119] ), .B(n9837), .S0(n5274), .Y(
        n11831) );
  CLKMX2X2 U11092 ( .A(\I_cache/cache[3][119] ), .B(n9837), .S0(n5142), .Y(
        n11832) );
  CLKMX2X2 U11093 ( .A(\I_cache/cache[2][119] ), .B(n9837), .S0(n5188), .Y(
        n11833) );
  CLKMX2X2 U11094 ( .A(\I_cache/cache[1][119] ), .B(n9837), .S0(n5048), .Y(
        n11834) );
  CLKMX2X2 U11095 ( .A(\I_cache/cache[0][119] ), .B(n9837), .S0(n5096), .Y(
        n11835) );
  CLKMX2X2 U11096 ( .A(\I_cache/cache[7][118] ), .B(n9873), .S0(n5319), .Y(
        n11836) );
  CLKMX2X2 U11097 ( .A(\I_cache/cache[6][118] ), .B(n9873), .S0(n5360), .Y(
        n11837) );
  CLKMX2X2 U11098 ( .A(\I_cache/cache[5][118] ), .B(n9873), .S0(n5230), .Y(
        n11838) );
  CLKMX2X2 U11099 ( .A(\I_cache/cache[4][118] ), .B(n9873), .S0(n5273), .Y(
        n11839) );
  CLKMX2X2 U11100 ( .A(\I_cache/cache[3][118] ), .B(n9873), .S0(n5141), .Y(
        n11840) );
  CLKMX2X2 U11101 ( .A(\I_cache/cache[1][118] ), .B(n9873), .S0(n5051), .Y(
        n11842) );
  CLKMX2X2 U11102 ( .A(\I_cache/cache[0][118] ), .B(n9873), .S0(n5097), .Y(
        n11843) );
  CLKMX2X2 U11103 ( .A(\I_cache/cache[7][117] ), .B(n9857), .S0(n5314), .Y(
        n11844) );
  CLKMX2X2 U11104 ( .A(\I_cache/cache[6][117] ), .B(n9857), .S0(n5366), .Y(
        n11845) );
  CLKMX2X2 U11105 ( .A(\I_cache/cache[5][117] ), .B(n9857), .S0(n5231), .Y(
        n11846) );
  CLKMX2X2 U11106 ( .A(\I_cache/cache[4][117] ), .B(n9857), .S0(n5274), .Y(
        n11847) );
  CLKMX2X2 U11107 ( .A(\I_cache/cache[3][117] ), .B(n9857), .S0(n5142), .Y(
        n11848) );
  CLKMX2X2 U11108 ( .A(\I_cache/cache[2][117] ), .B(n9857), .S0(n5188), .Y(
        n11849) );
  CLKMX2X2 U11109 ( .A(\I_cache/cache[1][117] ), .B(n9857), .S0(n5050), .Y(
        n11850) );
  CLKMX2X2 U11110 ( .A(\I_cache/cache[0][117] ), .B(n9857), .S0(n5096), .Y(
        n11851) );
  CLKMX2X2 U11111 ( .A(\I_cache/cache[7][116] ), .B(n158), .S0(n5314), .Y(
        n11852) );
  CLKMX2X2 U11112 ( .A(\I_cache/cache[6][116] ), .B(n158), .S0(n5366), .Y(
        n11853) );
  CLKMX2X2 U11113 ( .A(\I_cache/cache[5][116] ), .B(n158), .S0(n5225), .Y(
        n11854) );
  CLKMX2X2 U11114 ( .A(\I_cache/cache[4][116] ), .B(n158), .S0(n5273), .Y(
        n11855) );
  CLKMX2X2 U11115 ( .A(\I_cache/cache[3][116] ), .B(n158), .S0(n5135), .Y(
        n11856) );
  CLKMX2X2 U11116 ( .A(\I_cache/cache[2][116] ), .B(n158), .S0(n5181), .Y(
        n11857) );
  CLKMX2X2 U11117 ( .A(\I_cache/cache[1][116] ), .B(n158), .S0(n5052), .Y(
        n11858) );
  CLKMX2X2 U11118 ( .A(\I_cache/cache[0][116] ), .B(n158), .S0(n5091), .Y(
        n11859) );
  CLKMX2X2 U11119 ( .A(\I_cache/cache[7][115] ), .B(n11118), .S0(n5316), .Y(
        n11860) );
  CLKMX2X2 U11120 ( .A(\I_cache/cache[6][115] ), .B(n11118), .S0(n5359), .Y(
        n11861) );
  CLKMX2X2 U11121 ( .A(\I_cache/cache[5][115] ), .B(n11118), .S0(n5233), .Y(
        n11862) );
  CLKMX2X2 U11122 ( .A(\I_cache/cache[4][115] ), .B(n11118), .S0(n5273), .Y(
        n11863) );
  CLKMX2X2 U11123 ( .A(\I_cache/cache[3][115] ), .B(n11118), .S0(n5140), .Y(
        n11864) );
  CLKMX2X2 U11124 ( .A(\I_cache/cache[2][115] ), .B(n11118), .S0(n5187), .Y(
        n11865) );
  CLKMX2X2 U11125 ( .A(\I_cache/cache[1][115] ), .B(n11118), .S0(n5049), .Y(
        n11866) );
  CLKMX2X2 U11126 ( .A(\I_cache/cache[0][115] ), .B(n11118), .S0(n5093), .Y(
        n11867) );
  CLKMX2X2 U11127 ( .A(\I_cache/cache[7][114] ), .B(n153), .S0(n5315), .Y(
        n11868) );
  CLKMX2X2 U11128 ( .A(\I_cache/cache[6][114] ), .B(n153), .S0(n5358), .Y(
        n11869) );
  CLKMX2X2 U11129 ( .A(\I_cache/cache[5][114] ), .B(n153), .S0(n5226), .Y(
        n11870) );
  CLKMX2X2 U11130 ( .A(\I_cache/cache[4][114] ), .B(n153), .S0(n5269), .Y(
        n11871) );
  CLKMX2X2 U11131 ( .A(\I_cache/cache[3][114] ), .B(n153), .S0(n5136), .Y(
        n11872) );
  CLKMX2X2 U11132 ( .A(\I_cache/cache[2][114] ), .B(n153), .S0(n5182), .Y(
        n11873) );
  CLKMX2X2 U11133 ( .A(\I_cache/cache[1][114] ), .B(n153), .S0(n5046), .Y(
        n11874) );
  CLKMX2X2 U11134 ( .A(\I_cache/cache[0][114] ), .B(n153), .S0(n5092), .Y(
        n11875) );
  CLKMX2X2 U11135 ( .A(\I_cache/cache[7][113] ), .B(n10167), .S0(n5322), .Y(
        n11876) );
  CLKMX2X2 U11136 ( .A(\I_cache/cache[6][113] ), .B(n10167), .S0(n5360), .Y(
        n11877) );
  CLKMX2X2 U11137 ( .A(\I_cache/cache[5][113] ), .B(n10167), .S0(n5233), .Y(
        n11878) );
  CLKMX2X2 U11138 ( .A(\I_cache/cache[4][113] ), .B(n10167), .S0(n5277), .Y(
        n11879) );
  CLKMX2X2 U11139 ( .A(\I_cache/cache[3][113] ), .B(n10167), .S0(n5135), .Y(
        n11880) );
  CLKMX2X2 U11140 ( .A(\I_cache/cache[2][113] ), .B(n10167), .S0(n5183), .Y(
        n11881) );
  CLKMX2X2 U11141 ( .A(\I_cache/cache[1][113] ), .B(n10167), .S0(n5051), .Y(
        n11882) );
  CLKMX2X2 U11142 ( .A(\I_cache/cache[0][113] ), .B(n10167), .S0(n5099), .Y(
        n11883) );
  CLKMX2X2 U11143 ( .A(\I_cache/cache[7][112] ), .B(n9727), .S0(n5315), .Y(
        n11884) );
  CLKMX2X2 U11144 ( .A(\I_cache/cache[6][112] ), .B(n9727), .S0(n5360), .Y(
        n11885) );
  CLKMX2X2 U11145 ( .A(\I_cache/cache[5][112] ), .B(n9727), .S0(n5226), .Y(
        n11886) );
  CLKMX2X2 U11146 ( .A(\I_cache/cache[4][112] ), .B(n9727), .S0(n5269), .Y(
        n11887) );
  CLKMX2X2 U11147 ( .A(\I_cache/cache[3][112] ), .B(n9727), .S0(n5136), .Y(
        n11888) );
  CLKMX2X2 U11148 ( .A(\I_cache/cache[2][112] ), .B(n9727), .S0(n5182), .Y(
        n11889) );
  CLKMX2X2 U11149 ( .A(\I_cache/cache[1][112] ), .B(n9727), .S0(n5053), .Y(
        n11890) );
  CLKMX2X2 U11150 ( .A(\I_cache/cache[0][112] ), .B(n9727), .S0(n5092), .Y(
        n11891) );
  MX2XL U11151 ( .A(\I_cache/cache[5][111] ), .B(n9648), .S0(n5225), .Y(n11894) );
  MX2XL U11152 ( .A(\I_cache/cache[4][111] ), .B(n9648), .S0(n5270), .Y(n11895) );
  CLKMX2X2 U11153 ( .A(\I_cache/cache[7][110] ), .B(n9604), .S0(n5314), .Y(
        n11900) );
  CLKMX2X2 U11154 ( .A(\I_cache/cache[6][110] ), .B(n9604), .S0(n5366), .Y(
        n11901) );
  CLKMX2X2 U11155 ( .A(\I_cache/cache[5][110] ), .B(n9604), .S0(n5225), .Y(
        n11902) );
  CLKMX2X2 U11156 ( .A(\I_cache/cache[4][110] ), .B(n9604), .S0(n5274), .Y(
        n11903) );
  CLKMX2X2 U11157 ( .A(\I_cache/cache[3][110] ), .B(n9604), .S0(n5135), .Y(
        n11904) );
  CLKMX2X2 U11158 ( .A(\I_cache/cache[2][110] ), .B(n9604), .S0(n5181), .Y(
        n11905) );
  CLKMX2X2 U11159 ( .A(\I_cache/cache[1][110] ), .B(n9604), .S0(n5050), .Y(
        n11906) );
  CLKMX2X2 U11160 ( .A(\I_cache/cache[0][110] ), .B(n9604), .S0(n5091), .Y(
        n11907) );
  CLKMX2X2 U11161 ( .A(\I_cache/cache[6][109] ), .B(n9698), .S0(n5361), .Y(
        n11909) );
  CLKMX2X2 U11162 ( .A(\I_cache/cache[2][109] ), .B(n9698), .S0(n5182), .Y(
        n11913) );
  CLKMX2X2 U11163 ( .A(\I_cache/cache[1][109] ), .B(n9698), .S0(n5046), .Y(
        n11914) );
  CLKMX2X2 U11164 ( .A(\I_cache/cache[0][109] ), .B(n9698), .S0(n5092), .Y(
        n11915) );
  CLKMX2X2 U11165 ( .A(\I_cache/cache[6][107] ), .B(n9751), .S0(n5358), .Y(
        n11925) );
  CLKMX2X2 U11166 ( .A(\I_cache/cache[4][107] ), .B(n9751), .S0(n5273), .Y(
        n11927) );
  CLKMX2X2 U11167 ( .A(\I_cache/cache[2][107] ), .B(n9751), .S0(n5187), .Y(
        n11929) );
  CLKMX2X2 U11168 ( .A(\I_cache/cache[1][107] ), .B(n9751), .S0(n5048), .Y(
        n11930) );
  CLKMX2X2 U11169 ( .A(\I_cache/cache[0][107] ), .B(n9751), .S0(n5095), .Y(
        n11931) );
  CLKMX2X2 U11170 ( .A(\I_cache/cache[6][106] ), .B(n10054), .S0(n5359), .Y(
        n11933) );
  CLKMX2X2 U11171 ( .A(\I_cache/cache[2][106] ), .B(n10054), .S0(n5186), .Y(
        n11937) );
  CLKMX2X2 U11172 ( .A(\I_cache/cache[0][106] ), .B(n10054), .S0(n5095), .Y(
        n11939) );
  CLKMX2X2 U11173 ( .A(\I_cache/cache[7][101] ), .B(n9924), .S0(n5319), .Y(
        n11972) );
  CLKMX2X2 U11174 ( .A(\I_cache/cache[6][101] ), .B(n9924), .S0(n5359), .Y(
        n11973) );
  CLKMX2X2 U11175 ( .A(\I_cache/cache[5][101] ), .B(n9924), .S0(n5228), .Y(
        n11974) );
  CLKMX2X2 U11176 ( .A(\I_cache/cache[4][101] ), .B(n9924), .S0(n5274), .Y(
        n11975) );
  CLKMX2X2 U11177 ( .A(\I_cache/cache[3][101] ), .B(n9924), .S0(n5139), .Y(
        n11976) );
  CLKMX2X2 U11178 ( .A(\I_cache/cache[2][101] ), .B(n9924), .S0(n5185), .Y(
        n11977) );
  CLKMX2X2 U11179 ( .A(\I_cache/cache[1][101] ), .B(n9924), .S0(n5053), .Y(
        n11978) );
  CLKMX2X2 U11180 ( .A(\I_cache/cache[0][101] ), .B(n9924), .S0(n5092), .Y(
        n11979) );
  CLKMX2X2 U11181 ( .A(\I_cache/cache[7][98] ), .B(n11104), .S0(n5321), .Y(
        n11996) );
  CLKMX2X2 U11182 ( .A(\I_cache/cache[6][98] ), .B(n11104), .S0(n5358), .Y(
        n11997) );
  CLKMX2X2 U11183 ( .A(\I_cache/cache[5][98] ), .B(n11104), .S0(n5233), .Y(
        n11998) );
  CLKMX2X2 U11184 ( .A(\I_cache/cache[4][98] ), .B(n11104), .S0(n5276), .Y(
        n11999) );
  CLKMX2X2 U11185 ( .A(\I_cache/cache[3][98] ), .B(n11104), .S0(n5143), .Y(
        n12000) );
  CLKMX2X2 U11186 ( .A(\I_cache/cache[2][98] ), .B(n11104), .S0(n5189), .Y(
        n12001) );
  CLKMX2X2 U11187 ( .A(\I_cache/cache[1][98] ), .B(n11104), .S0(n5052), .Y(
        n12002) );
  CLKMX2X2 U11188 ( .A(\I_cache/cache[0][98] ), .B(n11104), .S0(n5091), .Y(
        n12003) );
  CLKMX2X2 U11189 ( .A(\I_cache/cache[7][95] ), .B(n154), .S0(n5317), .Y(
        n12020) );
  CLKMX2X2 U11190 ( .A(\I_cache/cache[6][95] ), .B(n154), .S0(n5364), .Y(
        n12021) );
  CLKMX2X2 U11191 ( .A(\I_cache/cache[5][95] ), .B(n154), .S0(n5233), .Y(
        n12022) );
  CLKMX2X2 U11192 ( .A(\I_cache/cache[4][95] ), .B(n154), .S0(n5271), .Y(
        n12023) );
  CLKMX2X2 U11193 ( .A(\I_cache/cache[3][95] ), .B(n154), .S0(n5138), .Y(
        n12024) );
  CLKMX2X2 U11194 ( .A(\I_cache/cache[2][95] ), .B(n154), .S0(n5184), .Y(
        n12025) );
  CLKMX2X2 U11195 ( .A(\I_cache/cache[1][95] ), .B(n154), .S0(n5047), .Y(
        n12026) );
  CLKMX2X2 U11196 ( .A(\I_cache/cache[0][95] ), .B(n154), .S0(n5094), .Y(
        n12027) );
  CLKMX2X2 U11197 ( .A(\I_cache/cache[7][94] ), .B(n6216), .S0(n5317), .Y(
        n12028) );
  CLKMX2X2 U11198 ( .A(\I_cache/cache[5][94] ), .B(n6216), .S0(n5226), .Y(
        n12030) );
  CLKMX2X2 U11199 ( .A(\I_cache/cache[4][94] ), .B(n6216), .S0(n5271), .Y(
        n12031) );
  CLKMX2X2 U11200 ( .A(\I_cache/cache[3][94] ), .B(n6216), .S0(n5138), .Y(
        n12032) );
  CLKMX2X2 U11201 ( .A(\I_cache/cache[2][94] ), .B(n6216), .S0(n5184), .Y(
        n12033) );
  CLKMX2X2 U11202 ( .A(\I_cache/cache[0][94] ), .B(n6216), .S0(n5094), .Y(
        n12035) );
  CLKMX2X2 U11203 ( .A(\I_cache/cache[7][93] ), .B(n6236), .S0(n5317), .Y(
        n12036) );
  CLKMX2X2 U11204 ( .A(\I_cache/cache[6][93] ), .B(n6236), .S0(n5359), .Y(
        n12037) );
  CLKMX2X2 U11205 ( .A(\I_cache/cache[5][93] ), .B(n6236), .S0(n5232), .Y(
        n12038) );
  CLKMX2X2 U11206 ( .A(\I_cache/cache[4][93] ), .B(n6236), .S0(n5271), .Y(
        n12039) );
  CLKMX2X2 U11207 ( .A(\I_cache/cache[3][93] ), .B(n6236), .S0(n5138), .Y(
        n12040) );
  CLKMX2X2 U11208 ( .A(\I_cache/cache[2][93] ), .B(n6236), .S0(n5184), .Y(
        n12041) );
  CLKMX2X2 U11209 ( .A(\I_cache/cache[1][93] ), .B(n6236), .S0(n5051), .Y(
        n12042) );
  CLKMX2X2 U11210 ( .A(\I_cache/cache[0][93] ), .B(n6236), .S0(n5093), .Y(
        n12043) );
  CLKMX2X2 U11211 ( .A(\I_cache/cache[7][92] ), .B(n6176), .S0(n5316), .Y(
        n12044) );
  CLKMX2X2 U11212 ( .A(\I_cache/cache[5][92] ), .B(n6176), .S0(n5227), .Y(
        n12046) );
  CLKMX2X2 U11213 ( .A(\I_cache/cache[4][92] ), .B(n6176), .S0(n5270), .Y(
        n12047) );
  CLKMX2X2 U11214 ( .A(\I_cache/cache[3][92] ), .B(n6176), .S0(n5137), .Y(
        n12048) );
  CLKMX2X2 U11215 ( .A(\I_cache/cache[2][92] ), .B(n6176), .S0(n5183), .Y(
        n12049) );
  CLKMX2X2 U11216 ( .A(\I_cache/cache[0][92] ), .B(n6176), .S0(n5093), .Y(
        n12051) );
  CLKMX2X2 U11217 ( .A(\I_cache/cache[7][91] ), .B(n11160), .S0(n5321), .Y(
        n12052) );
  CLKMX2X2 U11218 ( .A(\I_cache/cache[6][91] ), .B(n11160), .S0(n5363), .Y(
        n12053) );
  CLKMX2X2 U11219 ( .A(\I_cache/cache[5][91] ), .B(n11160), .S0(n5233), .Y(
        n12054) );
  CLKMX2X2 U11220 ( .A(\I_cache/cache[4][91] ), .B(n11160), .S0(n5276), .Y(
        n12055) );
  CLKMX2X2 U11221 ( .A(\I_cache/cache[3][91] ), .B(n11160), .S0(n5143), .Y(
        n12056) );
  CLKMX2X2 U11222 ( .A(\I_cache/cache[2][91] ), .B(n11160), .S0(n5189), .Y(
        n12057) );
  CLKMX2X2 U11223 ( .A(\I_cache/cache[1][91] ), .B(n11160), .S0(n5046), .Y(
        n12058) );
  CLKMX2X2 U11224 ( .A(\I_cache/cache[0][91] ), .B(n11160), .S0(n5098), .Y(
        n12059) );
  CLKMX2X2 U11225 ( .A(\I_cache/cache[7][90] ), .B(n9564), .S0(n5314), .Y(
        n12060) );
  CLKMX2X2 U11226 ( .A(\I_cache/cache[6][90] ), .B(n9564), .S0(n5358), .Y(
        n12061) );
  CLKMX2X2 U11227 ( .A(\I_cache/cache[5][90] ), .B(n9564), .S0(n5225), .Y(
        n12062) );
  CLKMX2X2 U11228 ( .A(\I_cache/cache[4][90] ), .B(n9564), .S0(n5276), .Y(
        n12063) );
  CLKMX2X2 U11229 ( .A(\I_cache/cache[3][90] ), .B(n9564), .S0(n5135), .Y(
        n12064) );
  CLKMX2X2 U11230 ( .A(\I_cache/cache[2][90] ), .B(n9564), .S0(n5181), .Y(
        n12065) );
  CLKMX2X2 U11231 ( .A(\I_cache/cache[1][90] ), .B(n9564), .S0(n5045), .Y(
        n12066) );
  CLKMX2X2 U11232 ( .A(\I_cache/cache[0][90] ), .B(n9564), .S0(n5091), .Y(
        n12067) );
  CLKMX2X2 U11233 ( .A(\I_cache/cache[7][89] ), .B(n9821), .S0(n5317), .Y(
        n12068) );
  CLKMX2X2 U11234 ( .A(\I_cache/cache[6][89] ), .B(n9821), .S0(n5358), .Y(
        n12069) );
  CLKMX2X2 U11235 ( .A(\I_cache/cache[5][89] ), .B(n9821), .S0(n5231), .Y(
        n12070) );
  CLKMX2X2 U11236 ( .A(\I_cache/cache[4][89] ), .B(n9821), .S0(n5274), .Y(
        n12071) );
  CLKMX2X2 U11237 ( .A(\I_cache/cache[3][89] ), .B(n9821), .S0(n5142), .Y(
        n12072) );
  CLKMX2X2 U11238 ( .A(\I_cache/cache[2][89] ), .B(n9821), .S0(n5188), .Y(
        n12073) );
  CLKMX2X2 U11239 ( .A(\I_cache/cache[1][89] ), .B(n9821), .S0(n5051), .Y(
        n12074) );
  CLKMX2X2 U11240 ( .A(\I_cache/cache[0][89] ), .B(n9821), .S0(n5096), .Y(
        n12075) );
  CLKMX2X2 U11241 ( .A(\I_cache/cache[7][88] ), .B(n9801), .S0(n5319), .Y(
        n12076) );
  CLKMX2X2 U11242 ( .A(\I_cache/cache[6][88] ), .B(n9801), .S0(n5365), .Y(
        n12077) );
  CLKMX2X2 U11243 ( .A(\I_cache/cache[5][88] ), .B(n9801), .S0(n5230), .Y(
        n12078) );
  CLKMX2X2 U11244 ( .A(\I_cache/cache[4][88] ), .B(n9801), .S0(n5273), .Y(
        n12079) );
  CLKMX2X2 U11245 ( .A(\I_cache/cache[3][88] ), .B(n9801), .S0(n5141), .Y(
        n12080) );
  CLKMX2X2 U11246 ( .A(\I_cache/cache[2][88] ), .B(n9801), .S0(n5187), .Y(
        n12081) );
  CLKMX2X2 U11247 ( .A(\I_cache/cache[1][88] ), .B(n9801), .S0(n5051), .Y(
        n12082) );
  CLKMX2X2 U11248 ( .A(\I_cache/cache[0][88] ), .B(n9801), .S0(n5098), .Y(
        n12083) );
  CLKMX2X2 U11249 ( .A(\I_cache/cache[7][87] ), .B(n9841), .S0(n5321), .Y(
        n12084) );
  CLKMX2X2 U11250 ( .A(\I_cache/cache[6][87] ), .B(n9841), .S0(n5366), .Y(
        n12085) );
  CLKMX2X2 U11251 ( .A(\I_cache/cache[5][87] ), .B(n9841), .S0(n5231), .Y(
        n12086) );
  CLKMX2X2 U11252 ( .A(\I_cache/cache[4][87] ), .B(n9841), .S0(n5274), .Y(
        n12087) );
  CLKMX2X2 U11253 ( .A(\I_cache/cache[3][87] ), .B(n9841), .S0(n5142), .Y(
        n12088) );
  CLKMX2X2 U11254 ( .A(\I_cache/cache[2][87] ), .B(n9841), .S0(n5188), .Y(
        n12089) );
  CLKMX2X2 U11255 ( .A(\I_cache/cache[1][87] ), .B(n9841), .S0(n5053), .Y(
        n12090) );
  CLKMX2X2 U11256 ( .A(\I_cache/cache[0][87] ), .B(n9841), .S0(n5096), .Y(
        n12091) );
  CLKMX2X2 U11257 ( .A(\I_cache/cache[7][86] ), .B(n9877), .S0(n5321), .Y(
        n12092) );
  CLKMX2X2 U11258 ( .A(\I_cache/cache[6][86] ), .B(n9877), .S0(n5358), .Y(
        n12093) );
  CLKMX2X2 U11259 ( .A(\I_cache/cache[5][86] ), .B(n9877), .S0(n5228), .Y(
        n12094) );
  CLKMX2X2 U11260 ( .A(\I_cache/cache[4][86] ), .B(n9877), .S0(n5277), .Y(
        n12095) );
  CLKMX2X2 U11261 ( .A(\I_cache/cache[3][86] ), .B(n9877), .S0(n5139), .Y(
        n12096) );
  CLKMX2X2 U11262 ( .A(\I_cache/cache[2][86] ), .B(n9877), .S0(n5185), .Y(
        n12097) );
  CLKMX2X2 U11263 ( .A(\I_cache/cache[1][86] ), .B(n9877), .S0(n5051), .Y(
        n12098) );
  CLKMX2X2 U11264 ( .A(\I_cache/cache[0][86] ), .B(n9877), .S0(n5094), .Y(
        n12099) );
  CLKMX2X2 U11265 ( .A(\I_cache/cache[7][85] ), .B(n9861), .S0(n5316), .Y(
        n12100) );
  CLKMX2X2 U11266 ( .A(\I_cache/cache[6][85] ), .B(n9861), .S0(n5366), .Y(
        n12101) );
  CLKMX2X2 U11267 ( .A(\I_cache/cache[5][85] ), .B(n9861), .S0(n5231), .Y(
        n12102) );
  CLKMX2X2 U11268 ( .A(\I_cache/cache[4][85] ), .B(n9861), .S0(n5274), .Y(
        n12103) );
  CLKMX2X2 U11269 ( .A(\I_cache/cache[3][85] ), .B(n9861), .S0(n5142), .Y(
        n12104) );
  CLKMX2X2 U11270 ( .A(\I_cache/cache[2][85] ), .B(n9861), .S0(n5188), .Y(
        n12105) );
  CLKMX2X2 U11271 ( .A(\I_cache/cache[1][85] ), .B(n9861), .S0(n5047), .Y(
        n12106) );
  CLKMX2X2 U11272 ( .A(\I_cache/cache[0][85] ), .B(n9861), .S0(n5096), .Y(
        n12107) );
  CLKMX2X2 U11273 ( .A(\I_cache/cache[7][84] ), .B(n141), .S0(n5314), .Y(
        n12108) );
  CLKMX2X2 U11274 ( .A(\I_cache/cache[6][84] ), .B(n141), .S0(n5358), .Y(
        n12109) );
  CLKMX2X2 U11275 ( .A(\I_cache/cache[5][84] ), .B(n141), .S0(n5225), .Y(
        n12110) );
  CLKMX2X2 U11276 ( .A(\I_cache/cache[4][84] ), .B(n141), .S0(n5277), .Y(
        n12111) );
  CLKMX2X2 U11277 ( .A(\I_cache/cache[3][84] ), .B(n141), .S0(n5135), .Y(
        n12112) );
  CLKMX2X2 U11278 ( .A(\I_cache/cache[2][84] ), .B(n141), .S0(n5181), .Y(
        n12113) );
  CLKMX2X2 U11279 ( .A(\I_cache/cache[1][84] ), .B(n141), .S0(n5050), .Y(
        n12114) );
  CLKMX2X2 U11280 ( .A(\I_cache/cache[0][84] ), .B(n141), .S0(n5091), .Y(
        n12115) );
  CLKMX2X2 U11281 ( .A(\I_cache/cache[7][83] ), .B(n11119), .S0(n5314), .Y(
        n12116) );
  CLKMX2X2 U11282 ( .A(\I_cache/cache[6][83] ), .B(n11119), .S0(n5362), .Y(
        n12117) );
  CLKMX2X2 U11283 ( .A(\I_cache/cache[5][83] ), .B(n11119), .S0(n5232), .Y(
        n12118) );
  CLKMX2X2 U11284 ( .A(\I_cache/cache[4][83] ), .B(n11119), .S0(n5272), .Y(
        n12119) );
  CLKMX2X2 U11285 ( .A(\I_cache/cache[3][83] ), .B(n11119), .S0(n5139), .Y(
        n12120) );
  CLKMX2X2 U11286 ( .A(\I_cache/cache[2][83] ), .B(n11119), .S0(n5183), .Y(
        n12121) );
  CLKMX2X2 U11287 ( .A(\I_cache/cache[1][83] ), .B(n11119), .S0(n5045), .Y(
        n12122) );
  CLKMX2X2 U11288 ( .A(\I_cache/cache[0][83] ), .B(n11119), .S0(n5099), .Y(
        n12123) );
  CLKMX2X2 U11289 ( .A(\I_cache/cache[7][82] ), .B(n162), .S0(n5315), .Y(
        n12124) );
  CLKMX2X2 U11290 ( .A(\I_cache/cache[6][82] ), .B(n162), .S0(n5359), .Y(
        n12125) );
  CLKMX2X2 U11291 ( .A(\I_cache/cache[5][82] ), .B(n162), .S0(n5226), .Y(
        n12126) );
  CLKMX2X2 U11292 ( .A(\I_cache/cache[4][82] ), .B(n162), .S0(n5269), .Y(
        n12127) );
  CLKMX2X2 U11293 ( .A(\I_cache/cache[3][82] ), .B(n162), .S0(n5136), .Y(
        n12128) );
  CLKMX2X2 U11294 ( .A(\I_cache/cache[2][82] ), .B(n162), .S0(n5182), .Y(
        n12129) );
  CLKMX2X2 U11295 ( .A(\I_cache/cache[1][82] ), .B(n162), .S0(n5050), .Y(
        n12130) );
  CLKMX2X2 U11296 ( .A(\I_cache/cache[0][82] ), .B(n162), .S0(n5092), .Y(
        n12131) );
  CLKMX2X2 U11297 ( .A(\I_cache/cache[7][81] ), .B(n10172), .S0(n5322), .Y(
        n12132) );
  CLKMX2X2 U11298 ( .A(\I_cache/cache[6][81] ), .B(n10172), .S0(n5363), .Y(
        n12133) );
  CLKMX2X2 U11299 ( .A(\I_cache/cache[5][81] ), .B(n10172), .S0(n5227), .Y(
        n12134) );
  CLKMX2X2 U11300 ( .A(\I_cache/cache[4][81] ), .B(n10172), .S0(n5277), .Y(
        n12135) );
  CLKMX2X2 U11301 ( .A(\I_cache/cache[3][81] ), .B(n10172), .S0(n5138), .Y(
        n12136) );
  CLKMX2X2 U11302 ( .A(\I_cache/cache[2][81] ), .B(n10172), .S0(n5186), .Y(
        n12137) );
  CLKMX2X2 U11303 ( .A(\I_cache/cache[1][81] ), .B(n10172), .S0(n5053), .Y(
        n12138) );
  CLKMX2X2 U11304 ( .A(\I_cache/cache[0][81] ), .B(n10172), .S0(n5099), .Y(
        n12139) );
  CLKMX2X2 U11305 ( .A(\I_cache/cache[7][80] ), .B(n9732), .S0(n5315), .Y(
        n12140) );
  CLKMX2X2 U11306 ( .A(\I_cache/cache[6][80] ), .B(n9732), .S0(n5360), .Y(
        n12141) );
  CLKMX2X2 U11307 ( .A(\I_cache/cache[5][80] ), .B(n9732), .S0(n5226), .Y(
        n12142) );
  CLKMX2X2 U11308 ( .A(\I_cache/cache[4][80] ), .B(n9732), .S0(n5269), .Y(
        n12143) );
  CLKMX2X2 U11309 ( .A(\I_cache/cache[3][80] ), .B(n9732), .S0(n5136), .Y(
        n12144) );
  CLKMX2X2 U11310 ( .A(\I_cache/cache[2][80] ), .B(n9732), .S0(n5182), .Y(
        n12145) );
  CLKMX2X2 U11311 ( .A(\I_cache/cache[1][80] ), .B(n9732), .S0(n5052), .Y(
        n12146) );
  CLKMX2X2 U11312 ( .A(\I_cache/cache[0][80] ), .B(n9732), .S0(n5095), .Y(
        n12147) );
  CLKMX2X2 U11313 ( .A(\I_cache/cache[7][78] ), .B(n9609), .S0(n5314), .Y(
        n12156) );
  CLKMX2X2 U11314 ( .A(\I_cache/cache[6][78] ), .B(n9609), .S0(n5361), .Y(
        n12157) );
  CLKMX2X2 U11315 ( .A(\I_cache/cache[5][78] ), .B(n9609), .S0(n5225), .Y(
        n12158) );
  CLKMX2X2 U11316 ( .A(\I_cache/cache[4][78] ), .B(n9609), .S0(n5272), .Y(
        n12159) );
  CLKMX2X2 U11317 ( .A(\I_cache/cache[3][78] ), .B(n9609), .S0(n5135), .Y(
        n12160) );
  CLKMX2X2 U11318 ( .A(\I_cache/cache[2][78] ), .B(n9609), .S0(n5181), .Y(
        n12161) );
  CLKMX2X2 U11319 ( .A(\I_cache/cache[1][78] ), .B(n9609), .S0(n5045), .Y(
        n12162) );
  CLKMX2X2 U11320 ( .A(\I_cache/cache[0][78] ), .B(n9609), .S0(n5091), .Y(
        n12163) );
  CLKMX2X2 U11321 ( .A(\I_cache/cache[2][77] ), .B(n9708), .S0(n5182), .Y(
        n12169) );
  CLKMX2X2 U11322 ( .A(\I_cache/cache[0][77] ), .B(n9708), .S0(n5092), .Y(
        n12171) );
  CLKMX2X2 U11323 ( .A(\I_cache/cache[7][76] ), .B(n9779), .S0(n5319), .Y(
        n12172) );
  CLKMX2X2 U11324 ( .A(\I_cache/cache[6][76] ), .B(n9779), .S0(n5363), .Y(
        n12173) );
  CLKMX2X2 U11325 ( .A(\I_cache/cache[5][76] ), .B(n9779), .S0(n5230), .Y(
        n12174) );
  CLKMX2X2 U11326 ( .A(\I_cache/cache[4][76] ), .B(n9779), .S0(n5273), .Y(
        n12175) );
  CLKMX2X2 U11327 ( .A(\I_cache/cache[3][76] ), .B(n9779), .S0(n5141), .Y(
        n12176) );
  CLKMX2X2 U11328 ( .A(\I_cache/cache[2][76] ), .B(n9779), .S0(n5187), .Y(
        n12177) );
  CLKMX2X2 U11329 ( .A(\I_cache/cache[1][76] ), .B(n9779), .S0(n5049), .Y(
        n12178) );
  CLKMX2X2 U11330 ( .A(\I_cache/cache[0][76] ), .B(n9779), .S0(n5095), .Y(
        n12179) );
  CLKMX2X2 U11331 ( .A(\I_cache/cache[6][75] ), .B(n9756), .S0(n5362), .Y(
        n12181) );
  CLKMX2X2 U11332 ( .A(\I_cache/cache[4][75] ), .B(n9756), .S0(n5273), .Y(
        n12183) );
  CLKMX2X2 U11333 ( .A(\I_cache/cache[2][75] ), .B(n9756), .S0(n5187), .Y(
        n12185) );
  CLKMX2X2 U11334 ( .A(\I_cache/cache[0][75] ), .B(n9756), .S0(n5095), .Y(
        n12187) );
  CLKMX2X2 U11335 ( .A(\I_cache/cache[7][74] ), .B(n10059), .S0(n5318), .Y(
        n12188) );
  CLKMX2X2 U11336 ( .A(\I_cache/cache[6][74] ), .B(n10059), .S0(n5364), .Y(
        n12189) );
  CLKMX2X2 U11337 ( .A(\I_cache/cache[3][74] ), .B(n10059), .S0(n5140), .Y(
        n12192) );
  CLKMX2X2 U11338 ( .A(\I_cache/cache[2][74] ), .B(n10059), .S0(n5186), .Y(
        n12193) );
  CLKMX2X2 U11339 ( .A(\I_cache/cache[1][74] ), .B(n10059), .S0(n5049), .Y(
        n12194) );
  CLKMX2X2 U11340 ( .A(\I_cache/cache[0][74] ), .B(n10059), .S0(n5093), .Y(
        n12195) );
  CLKMX2X2 U11341 ( .A(\I_cache/cache[7][69] ), .B(n9929), .S0(n5317), .Y(
        n12228) );
  CLKMX2X2 U11342 ( .A(\I_cache/cache[6][69] ), .B(n9929), .S0(n5362), .Y(
        n12229) );
  CLKMX2X2 U11343 ( .A(\I_cache/cache[5][69] ), .B(n9929), .S0(n5228), .Y(
        n12230) );
  CLKMX2X2 U11344 ( .A(\I_cache/cache[4][69] ), .B(n9929), .S0(n5272), .Y(
        n12231) );
  CLKMX2X2 U11345 ( .A(\I_cache/cache[3][69] ), .B(n9929), .S0(n5139), .Y(
        n12232) );
  CLKMX2X2 U11346 ( .A(\I_cache/cache[2][69] ), .B(n9929), .S0(n5185), .Y(
        n12233) );
  CLKMX2X2 U11347 ( .A(\I_cache/cache[1][69] ), .B(n9929), .S0(n5048), .Y(
        n12234) );
  CLKMX2X2 U11348 ( .A(\I_cache/cache[0][69] ), .B(n9929), .S0(n5091), .Y(
        n12235) );
  CLKMX2X2 U11349 ( .A(\I_cache/cache[7][66] ), .B(n11105), .S0(n5314), .Y(
        n12252) );
  CLKMX2X2 U11350 ( .A(\I_cache/cache[6][66] ), .B(n11105), .S0(n5363), .Y(
        n12253) );
  CLKMX2X2 U11351 ( .A(\I_cache/cache[5][66] ), .B(n11105), .S0(n5225), .Y(
        n12254) );
  CLKMX2X2 U11352 ( .A(\I_cache/cache[4][66] ), .B(n11105), .S0(n5275), .Y(
        n12255) );
  CLKMX2X2 U11353 ( .A(\I_cache/cache[3][66] ), .B(n11105), .S0(n5135), .Y(
        n12256) );
  CLKMX2X2 U11354 ( .A(\I_cache/cache[2][66] ), .B(n11105), .S0(n5181), .Y(
        n12257) );
  CLKMX2X2 U11355 ( .A(\I_cache/cache[1][66] ), .B(n11105), .S0(n5046), .Y(
        n12258) );
  CLKMX2X2 U11356 ( .A(\I_cache/cache[0][66] ), .B(n11105), .S0(n5097), .Y(
        n12259) );
  CLKMX2X2 U11357 ( .A(\I_cache/cache[7][63] ), .B(n165), .S0(n5316), .Y(
        n12276) );
  CLKMX2X2 U11358 ( .A(\I_cache/cache[6][63] ), .B(n165), .S0(n5362), .Y(
        n12277) );
  CLKMX2X2 U11359 ( .A(\I_cache/cache[5][63] ), .B(n165), .S0(n5227), .Y(
        n12278) );
  CLKMX2X2 U11360 ( .A(\I_cache/cache[4][63] ), .B(n165), .S0(n5270), .Y(
        n12279) );
  CLKMX2X2 U11361 ( .A(\I_cache/cache[3][63] ), .B(n165), .S0(n5137), .Y(
        n12280) );
  CLKMX2X2 U11362 ( .A(\I_cache/cache[2][63] ), .B(n165), .S0(n5183), .Y(
        n12281) );
  CLKMX2X2 U11363 ( .A(\I_cache/cache[1][63] ), .B(n165), .S0(n5053), .Y(
        n12282) );
  CLKMX2X2 U11364 ( .A(\I_cache/cache[0][63] ), .B(n165), .S0(n5094), .Y(
        n12283) );
  CLKMX2X2 U11365 ( .A(\I_cache/cache[7][62] ), .B(n161), .S0(n5317), .Y(
        n12284) );
  CLKMX2X2 U11366 ( .A(\I_cache/cache[6][62] ), .B(n161), .S0(n5360), .Y(
        n12285) );
  CLKMX2X2 U11367 ( .A(\I_cache/cache[5][62] ), .B(n161), .S0(n5227), .Y(
        n12286) );
  CLKMX2X2 U11368 ( .A(\I_cache/cache[4][62] ), .B(n161), .S0(n5271), .Y(
        n12287) );
  CLKMX2X2 U11369 ( .A(\I_cache/cache[3][62] ), .B(n161), .S0(n5138), .Y(
        n12288) );
  CLKMX2X2 U11370 ( .A(\I_cache/cache[2][62] ), .B(n161), .S0(n5184), .Y(
        n12289) );
  CLKMX2X2 U11371 ( .A(\I_cache/cache[1][62] ), .B(n161), .S0(n5047), .Y(
        n12290) );
  CLKMX2X2 U11372 ( .A(\I_cache/cache[0][62] ), .B(n161), .S0(n5094), .Y(
        n12291) );
  CLKMX2X2 U11373 ( .A(\I_cache/cache[7][61] ), .B(n152), .S0(n5317), .Y(
        n12292) );
  CLKMX2X2 U11374 ( .A(\I_cache/cache[6][61] ), .B(n152), .S0(n5364), .Y(
        n12293) );
  CLKMX2X2 U11375 ( .A(\I_cache/cache[5][61] ), .B(n152), .S0(n5231), .Y(
        n12294) );
  CLKMX2X2 U11376 ( .A(\I_cache/cache[4][61] ), .B(n152), .S0(n5271), .Y(
        n12295) );
  CLKMX2X2 U11377 ( .A(\I_cache/cache[3][61] ), .B(n152), .S0(n5138), .Y(
        n12296) );
  CLKMX2X2 U11378 ( .A(\I_cache/cache[2][61] ), .B(n152), .S0(n5184), .Y(
        n12297) );
  CLKMX2X2 U11379 ( .A(\I_cache/cache[1][61] ), .B(n152), .S0(n5050), .Y(
        n12298) );
  CLKMX2X2 U11380 ( .A(\I_cache/cache[0][61] ), .B(n152), .S0(n5094), .Y(
        n12299) );
  CLKMX2X2 U11381 ( .A(\I_cache/cache[7][60] ), .B(n6166), .S0(n5316), .Y(
        n12300) );
  CLKMX2X2 U11382 ( .A(\I_cache/cache[6][60] ), .B(n6166), .S0(n5358), .Y(
        n12301) );
  CLKMX2X2 U11383 ( .A(\I_cache/cache[5][60] ), .B(n6166), .S0(n5227), .Y(
        n12302) );
  CLKMX2X2 U11384 ( .A(\I_cache/cache[4][60] ), .B(n6166), .S0(n5270), .Y(
        n12303) );
  CLKMX2X2 U11385 ( .A(\I_cache/cache[3][60] ), .B(n6166), .S0(n5137), .Y(
        n12304) );
  CLKMX2X2 U11386 ( .A(\I_cache/cache[2][60] ), .B(n6166), .S0(n5183), .Y(
        n12305) );
  CLKMX2X2 U11387 ( .A(\I_cache/cache[1][60] ), .B(n6166), .S0(n5051), .Y(
        n12306) );
  CLKMX2X2 U11388 ( .A(\I_cache/cache[0][60] ), .B(n6166), .S0(n5093), .Y(
        n12307) );
  CLKMX2X2 U11389 ( .A(\I_cache/cache[7][59] ), .B(n11158), .S0(n5321), .Y(
        n12308) );
  CLKMX2X2 U11390 ( .A(\I_cache/cache[6][59] ), .B(n11158), .S0(n5366), .Y(
        n12309) );
  CLKMX2X2 U11391 ( .A(\I_cache/cache[5][59] ), .B(n11158), .S0(n5233), .Y(
        n12310) );
  CLKMX2X2 U11392 ( .A(\I_cache/cache[4][59] ), .B(n11158), .S0(n5276), .Y(
        n12311) );
  CLKMX2X2 U11393 ( .A(\I_cache/cache[3][59] ), .B(n11158), .S0(n5143), .Y(
        n12312) );
  CLKMX2X2 U11394 ( .A(\I_cache/cache[2][59] ), .B(n11158), .S0(n5189), .Y(
        n12313) );
  CLKMX2X2 U11395 ( .A(\I_cache/cache[1][59] ), .B(n11158), .S0(n5052), .Y(
        n12314) );
  CLKMX2X2 U11396 ( .A(\I_cache/cache[0][59] ), .B(n11158), .S0(n5098), .Y(
        n12315) );
  CLKMX2X2 U11397 ( .A(\I_cache/cache[7][58] ), .B(n9562), .S0(n5316), .Y(
        n12316) );
  CLKMX2X2 U11398 ( .A(\I_cache/cache[6][58] ), .B(n9562), .S0(n5366), .Y(
        n12317) );
  CLKMX2X2 U11399 ( .A(\I_cache/cache[5][58] ), .B(n9562), .S0(n5227), .Y(
        n12318) );
  CLKMX2X2 U11400 ( .A(\I_cache/cache[4][58] ), .B(n9562), .S0(n5270), .Y(
        n12319) );
  CLKMX2X2 U11401 ( .A(\I_cache/cache[3][58] ), .B(n9562), .S0(n5137), .Y(
        n12320) );
  CLKMX2X2 U11402 ( .A(\I_cache/cache[2][58] ), .B(n9562), .S0(n5183), .Y(
        n12321) );
  CLKMX2X2 U11403 ( .A(\I_cache/cache[1][58] ), .B(n9562), .S0(n5050), .Y(
        n12322) );
  CLKMX2X2 U11404 ( .A(\I_cache/cache[0][58] ), .B(n9562), .S0(n5091), .Y(
        n12323) );
  CLKMX2X2 U11405 ( .A(\I_cache/cache[7][57] ), .B(n156), .S0(n5318), .Y(
        n12324) );
  CLKMX2X2 U11406 ( .A(\I_cache/cache[6][57] ), .B(n156), .S0(n5361), .Y(
        n12325) );
  CLKMX2X2 U11407 ( .A(\I_cache/cache[5][57] ), .B(n156), .S0(n5229), .Y(
        n12326) );
  CLKMX2X2 U11408 ( .A(\I_cache/cache[4][57] ), .B(n156), .S0(n5272), .Y(
        n12327) );
  CLKMX2X2 U11409 ( .A(\I_cache/cache[3][57] ), .B(n156), .S0(n5140), .Y(
        n12328) );
  CLKMX2X2 U11410 ( .A(\I_cache/cache[2][57] ), .B(n156), .S0(n5186), .Y(
        n12329) );
  CLKMX2X2 U11411 ( .A(\I_cache/cache[1][57] ), .B(n156), .S0(n5045), .Y(
        n12330) );
  CLKMX2X2 U11412 ( .A(\I_cache/cache[0][57] ), .B(n156), .S0(n5096), .Y(
        n12331) );
  CLKMX2X2 U11413 ( .A(\I_cache/cache[7][56] ), .B(n9793), .S0(n5319), .Y(
        n12332) );
  CLKMX2X2 U11414 ( .A(\I_cache/cache[6][56] ), .B(n9793), .S0(n5363), .Y(
        n12333) );
  CLKMX2X2 U11415 ( .A(\I_cache/cache[5][56] ), .B(n9793), .S0(n5230), .Y(
        n12334) );
  CLKMX2X2 U11416 ( .A(\I_cache/cache[4][56] ), .B(n9793), .S0(n5273), .Y(
        n12335) );
  CLKMX2X2 U11417 ( .A(\I_cache/cache[3][56] ), .B(n9793), .S0(n5141), .Y(
        n12336) );
  CLKMX2X2 U11418 ( .A(\I_cache/cache[2][56] ), .B(n9793), .S0(n5187), .Y(
        n12337) );
  CLKMX2X2 U11419 ( .A(\I_cache/cache[1][56] ), .B(n9793), .S0(n5052), .Y(
        n12338) );
  CLKMX2X2 U11420 ( .A(\I_cache/cache[0][56] ), .B(n9793), .S0(n5095), .Y(
        n12339) );
  CLKMX2X2 U11421 ( .A(\I_cache/cache[7][55] ), .B(n9833), .S0(n5318), .Y(
        n12340) );
  CLKMX2X2 U11422 ( .A(\I_cache/cache[6][55] ), .B(n9833), .S0(n5363), .Y(
        n12341) );
  CLKMX2X2 U11423 ( .A(\I_cache/cache[5][55] ), .B(n9833), .S0(n5231), .Y(
        n12342) );
  CLKMX2X2 U11424 ( .A(\I_cache/cache[4][55] ), .B(n9833), .S0(n5274), .Y(
        n12343) );
  CLKMX2X2 U11425 ( .A(\I_cache/cache[3][55] ), .B(n9833), .S0(n5142), .Y(
        n12344) );
  CLKMX2X2 U11426 ( .A(\I_cache/cache[2][55] ), .B(n9833), .S0(n5188), .Y(
        n12345) );
  CLKMX2X2 U11427 ( .A(\I_cache/cache[1][55] ), .B(n9833), .S0(n5048), .Y(
        n12346) );
  CLKMX2X2 U11428 ( .A(\I_cache/cache[0][55] ), .B(n9833), .S0(n5096), .Y(
        n12347) );
  CLKMX2X2 U11429 ( .A(\I_cache/cache[7][54] ), .B(n9869), .S0(n5319), .Y(
        n12348) );
  CLKMX2X2 U11430 ( .A(\I_cache/cache[6][54] ), .B(n9869), .S0(n5358), .Y(
        n12349) );
  CLKMX2X2 U11431 ( .A(\I_cache/cache[5][54] ), .B(n9869), .S0(n5231), .Y(
        n12350) );
  CLKMX2X2 U11432 ( .A(\I_cache/cache[4][54] ), .B(n9869), .S0(n5274), .Y(
        n12351) );
  CLKMX2X2 U11433 ( .A(\I_cache/cache[3][54] ), .B(n9869), .S0(n5142), .Y(
        n12352) );
  CLKMX2X2 U11434 ( .A(\I_cache/cache[2][54] ), .B(n9869), .S0(n5188), .Y(
        n12353) );
  CLKMX2X2 U11435 ( .A(\I_cache/cache[1][54] ), .B(n9869), .S0(n5047), .Y(
        n12354) );
  CLKMX2X2 U11436 ( .A(\I_cache/cache[0][54] ), .B(n9869), .S0(n5093), .Y(
        n12355) );
  CLKMX2X2 U11437 ( .A(\I_cache/cache[7][53] ), .B(n9853), .S0(n5322), .Y(
        n12356) );
  CLKMX2X2 U11438 ( .A(\I_cache/cache[6][53] ), .B(n9853), .S0(n5362), .Y(
        n12357) );
  CLKMX2X2 U11439 ( .A(\I_cache/cache[5][53] ), .B(n9853), .S0(n5231), .Y(
        n12358) );
  CLKMX2X2 U11440 ( .A(\I_cache/cache[4][53] ), .B(n9853), .S0(n5274), .Y(
        n12359) );
  CLKMX2X2 U11441 ( .A(\I_cache/cache[3][53] ), .B(n9853), .S0(n5142), .Y(
        n12360) );
  CLKMX2X2 U11442 ( .A(\I_cache/cache[2][53] ), .B(n9853), .S0(n5188), .Y(
        n12361) );
  CLKMX2X2 U11443 ( .A(\I_cache/cache[1][53] ), .B(n9853), .S0(n5045), .Y(
        n12362) );
  CLKMX2X2 U11444 ( .A(\I_cache/cache[0][53] ), .B(n9853), .S0(n5096), .Y(
        n12363) );
  CLKMX2X2 U11445 ( .A(\I_cache/cache[7][52] ), .B(n9624), .S0(n5314), .Y(
        n12364) );
  CLKMX2X2 U11446 ( .A(\I_cache/cache[6][52] ), .B(n9624), .S0(n5366), .Y(
        n12365) );
  CLKMX2X2 U11447 ( .A(\I_cache/cache[5][52] ), .B(n9624), .S0(n5225), .Y(
        n12366) );
  CLKMX2X2 U11448 ( .A(\I_cache/cache[4][52] ), .B(n9624), .S0(n5269), .Y(
        n12367) );
  CLKMX2X2 U11449 ( .A(\I_cache/cache[3][52] ), .B(n9624), .S0(n5135), .Y(
        n12368) );
  CLKMX2X2 U11450 ( .A(\I_cache/cache[2][52] ), .B(n9624), .S0(n5181), .Y(
        n12369) );
  CLKMX2X2 U11451 ( .A(\I_cache/cache[1][52] ), .B(n9624), .S0(n5048), .Y(
        n12370) );
  CLKMX2X2 U11452 ( .A(\I_cache/cache[0][52] ), .B(n9624), .S0(n5091), .Y(
        n12371) );
  CLKMX2X2 U11453 ( .A(\I_cache/cache[7][51] ), .B(n11117), .S0(n5318), .Y(
        n12372) );
  CLKMX2X2 U11454 ( .A(\I_cache/cache[6][51] ), .B(n11117), .S0(n5365), .Y(
        n12373) );
  CLKMX2X2 U11455 ( .A(\I_cache/cache[5][51] ), .B(n11117), .S0(n5228), .Y(
        n12374) );
  CLKMX2X2 U11456 ( .A(\I_cache/cache[4][51] ), .B(n11117), .S0(n5276), .Y(
        n12375) );
  CLKMX2X2 U11457 ( .A(\I_cache/cache[3][51] ), .B(n11117), .S0(n5136), .Y(
        n12376) );
  CLKMX2X2 U11458 ( .A(\I_cache/cache[2][51] ), .B(n11117), .S0(n5182), .Y(
        n12377) );
  CLKMX2X2 U11459 ( .A(\I_cache/cache[1][51] ), .B(n11117), .S0(n5050), .Y(
        n12378) );
  CLKMX2X2 U11460 ( .A(\I_cache/cache[0][51] ), .B(n11117), .S0(n5095), .Y(
        n12379) );
  CLKMX2X2 U11461 ( .A(\I_cache/cache[7][50] ), .B(n155), .S0(n5315), .Y(
        n12380) );
  CLKMX2X2 U11462 ( .A(\I_cache/cache[6][50] ), .B(n155), .S0(n5365), .Y(
        n12381) );
  CLKMX2X2 U11463 ( .A(\I_cache/cache[5][50] ), .B(n155), .S0(n5226), .Y(
        n12382) );
  CLKMX2X2 U11464 ( .A(\I_cache/cache[4][50] ), .B(n155), .S0(n5269), .Y(
        n12383) );
  CLKMX2X2 U11465 ( .A(\I_cache/cache[3][50] ), .B(n155), .S0(n5136), .Y(
        n12384) );
  CLKMX2X2 U11466 ( .A(\I_cache/cache[2][50] ), .B(n155), .S0(n5182), .Y(
        n12385) );
  CLKMX2X2 U11467 ( .A(\I_cache/cache[1][50] ), .B(n155), .S0(n5050), .Y(
        n12386) );
  CLKMX2X2 U11468 ( .A(\I_cache/cache[0][50] ), .B(n155), .S0(n5092), .Y(
        n12387) );
  CLKMX2X2 U11469 ( .A(\I_cache/cache[7][49] ), .B(n10162), .S0(n5322), .Y(
        n12388) );
  CLKMX2X2 U11470 ( .A(\I_cache/cache[6][49] ), .B(n10162), .S0(n5364), .Y(
        n12389) );
  CLKMX2X2 U11471 ( .A(\I_cache/cache[5][49] ), .B(n10162), .S0(n5225), .Y(
        n12390) );
  CLKMX2X2 U11472 ( .A(\I_cache/cache[4][49] ), .B(n10162), .S0(n5277), .Y(
        n12391) );
  CLKMX2X2 U11473 ( .A(\I_cache/cache[3][49] ), .B(n10162), .S0(n5143), .Y(
        n12392) );
  CLKMX2X2 U11474 ( .A(\I_cache/cache[2][49] ), .B(n10162), .S0(n5188), .Y(
        n12393) );
  CLKMX2X2 U11475 ( .A(\I_cache/cache[1][49] ), .B(n10162), .S0(n5045), .Y(
        n12394) );
  CLKMX2X2 U11476 ( .A(\I_cache/cache[0][49] ), .B(n10162), .S0(n5099), .Y(
        n12395) );
  CLKMX2X2 U11477 ( .A(\I_cache/cache[7][48] ), .B(n9722), .S0(n5315), .Y(
        n12396) );
  CLKMX2X2 U11478 ( .A(\I_cache/cache[6][48] ), .B(n9722), .S0(n5361), .Y(
        n12397) );
  CLKMX2X2 U11479 ( .A(\I_cache/cache[5][48] ), .B(n9722), .S0(n5226), .Y(
        n12398) );
  CLKMX2X2 U11480 ( .A(\I_cache/cache[4][48] ), .B(n9722), .S0(n5269), .Y(
        n12399) );
  CLKMX2X2 U11481 ( .A(\I_cache/cache[3][48] ), .B(n9722), .S0(n5136), .Y(
        n12400) );
  CLKMX2X2 U11482 ( .A(\I_cache/cache[2][48] ), .B(n9722), .S0(n5182), .Y(
        n12401) );
  CLKMX2X2 U11483 ( .A(\I_cache/cache[1][48] ), .B(n9722), .S0(n5050), .Y(
        n12402) );
  CLKMX2X2 U11484 ( .A(\I_cache/cache[0][48] ), .B(n9722), .S0(n5092), .Y(
        n12403) );
  MX2XL U11485 ( .A(\I_cache/cache[7][47] ), .B(n9653), .S0(n5314), .Y(n12404)
         );
  MX2XL U11486 ( .A(\I_cache/cache[6][47] ), .B(n9653), .S0(n5359), .Y(n12405)
         );
  CLKMX2X2 U11487 ( .A(\I_cache/cache[7][46] ), .B(n9599), .S0(n5314), .Y(
        n12412) );
  CLKMX2X2 U11488 ( .A(\I_cache/cache[6][46] ), .B(n9599), .S0(n5365), .Y(
        n12413) );
  CLKMX2X2 U11489 ( .A(\I_cache/cache[5][46] ), .B(n9599), .S0(n5225), .Y(
        n12414) );
  CLKMX2X2 U11490 ( .A(\I_cache/cache[4][46] ), .B(n9599), .S0(n5271), .Y(
        n12415) );
  CLKMX2X2 U11491 ( .A(\I_cache/cache[3][46] ), .B(n9599), .S0(n5135), .Y(
        n12416) );
  CLKMX2X2 U11492 ( .A(\I_cache/cache[2][46] ), .B(n9599), .S0(n5181), .Y(
        n12417) );
  CLKMX2X2 U11493 ( .A(\I_cache/cache[1][46] ), .B(n9599), .S0(n5046), .Y(
        n12418) );
  CLKMX2X2 U11494 ( .A(\I_cache/cache[0][46] ), .B(n9599), .S0(n5091), .Y(
        n12419) );
  CLKMX2X2 U11495 ( .A(\I_cache/cache[2][45] ), .B(n9703), .S0(n5182), .Y(
        n12425) );
  CLKMX2X2 U11496 ( .A(\I_cache/cache[0][45] ), .B(n9703), .S0(n5092), .Y(
        n12427) );
  CLKMX2X2 U11497 ( .A(\I_cache/cache[7][44] ), .B(n9769), .S0(n5319), .Y(
        n12428) );
  CLKMX2X2 U11498 ( .A(\I_cache/cache[6][44] ), .B(n9769), .S0(n5361), .Y(
        n12429) );
  CLKMX2X2 U11499 ( .A(\I_cache/cache[5][44] ), .B(n9769), .S0(n5230), .Y(
        n12430) );
  CLKMX2X2 U11500 ( .A(\I_cache/cache[4][44] ), .B(n9769), .S0(n5273), .Y(
        n12431) );
  CLKMX2X2 U11501 ( .A(\I_cache/cache[3][44] ), .B(n9769), .S0(n5141), .Y(
        n12432) );
  CLKMX2X2 U11502 ( .A(\I_cache/cache[2][44] ), .B(n9769), .S0(n5187), .Y(
        n12433) );
  CLKMX2X2 U11503 ( .A(\I_cache/cache[1][44] ), .B(n9769), .S0(n5046), .Y(
        n12434) );
  CLKMX2X2 U11504 ( .A(\I_cache/cache[0][44] ), .B(n9769), .S0(n5095), .Y(
        n12435) );
  CLKMX2X2 U11505 ( .A(\I_cache/cache[6][43] ), .B(n9746), .S0(n5362), .Y(
        n12437) );
  CLKMX2X2 U11506 ( .A(\I_cache/cache[4][43] ), .B(n9746), .S0(n5273), .Y(
        n12439) );
  CLKMX2X2 U11507 ( .A(\I_cache/cache[3][43] ), .B(n9746), .S0(n5141), .Y(
        n12440) );
  CLKMX2X2 U11508 ( .A(\I_cache/cache[2][43] ), .B(n9746), .S0(n5187), .Y(
        n12441) );
  CLKMX2X2 U11509 ( .A(\I_cache/cache[1][43] ), .B(n9746), .S0(n5050), .Y(
        n12442) );
  CLKMX2X2 U11510 ( .A(\I_cache/cache[0][43] ), .B(n9746), .S0(n5095), .Y(
        n12443) );
  CLKMX2X2 U11511 ( .A(\I_cache/cache[6][42] ), .B(n10049), .S0(n5363), .Y(
        n12445) );
  CLKMX2X2 U11512 ( .A(\I_cache/cache[4][42] ), .B(n10049), .S0(n5272), .Y(
        n12447) );
  CLKMX2X2 U11513 ( .A(\I_cache/cache[2][42] ), .B(n10049), .S0(n5186), .Y(
        n12449) );
  CLKMX2X2 U11514 ( .A(\I_cache/cache[0][42] ), .B(n10049), .S0(n5097), .Y(
        n12451) );
  CLKMX2X2 U11515 ( .A(\I_cache/cache[7][37] ), .B(n180), .S0(n5319), .Y(
        n12484) );
  CLKMX2X2 U11516 ( .A(\I_cache/cache[6][37] ), .B(n180), .S0(n5360), .Y(
        n12485) );
  CLKMX2X2 U11517 ( .A(\I_cache/cache[5][37] ), .B(n180), .S0(n5228), .Y(
        n12486) );
  CLKMX2X2 U11518 ( .A(\I_cache/cache[4][37] ), .B(n180), .S0(n5271), .Y(
        n12487) );
  CLKMX2X2 U11519 ( .A(\I_cache/cache[3][37] ), .B(n180), .S0(n5139), .Y(
        n12488) );
  CLKMX2X2 U11520 ( .A(\I_cache/cache[2][37] ), .B(n180), .S0(n5185), .Y(
        n12489) );
  CLKMX2X2 U11521 ( .A(\I_cache/cache[1][37] ), .B(n180), .S0(n5053), .Y(
        n12490) );
  CLKMX2X2 U11522 ( .A(\I_cache/cache[0][37] ), .B(n180), .S0(n5096), .Y(
        n12491) );
  CLKMX2X2 U11523 ( .A(\I_cache/cache[7][34] ), .B(n11103), .S0(n5322), .Y(
        n12508) );
  CLKMX2X2 U11524 ( .A(\I_cache/cache[6][34] ), .B(n11103), .S0(n5365), .Y(
        n12509) );
  CLKMX2X2 U11525 ( .A(\I_cache/cache[5][34] ), .B(n11103), .S0(n5232), .Y(
        n12510) );
  CLKMX2X2 U11526 ( .A(\I_cache/cache[4][34] ), .B(n11103), .S0(n5277), .Y(
        n12511) );
  CLKMX2X2 U11527 ( .A(\I_cache/cache[3][34] ), .B(n11103), .S0(n5136), .Y(
        n12512) );
  CLKMX2X2 U11528 ( .A(\I_cache/cache[2][34] ), .B(n11103), .S0(n5185), .Y(
        n12513) );
  CLKMX2X2 U11529 ( .A(\I_cache/cache[1][34] ), .B(n11103), .S0(n5052), .Y(
        n12514) );
  CLKMX2X2 U11530 ( .A(\I_cache/cache[0][34] ), .B(n11103), .S0(n5098), .Y(
        n12515) );
  CLKMX2X2 U11531 ( .A(\I_cache/cache[7][31] ), .B(n159), .S0(n5316), .Y(
        n12532) );
  CLKMX2X2 U11532 ( .A(\I_cache/cache[6][31] ), .B(n159), .S0(n5364), .Y(
        n12533) );
  CLKMX2X2 U11533 ( .A(\I_cache/cache[5][31] ), .B(n159), .S0(n5227), .Y(
        n12534) );
  CLKMX2X2 U11534 ( .A(\I_cache/cache[4][31] ), .B(n159), .S0(n5270), .Y(
        n12535) );
  CLKMX2X2 U11535 ( .A(\I_cache/cache[3][31] ), .B(n159), .S0(n5137), .Y(
        n12536) );
  CLKMX2X2 U11536 ( .A(\I_cache/cache[2][31] ), .B(n159), .S0(n5183), .Y(
        n12537) );
  CLKMX2X2 U11537 ( .A(\I_cache/cache[1][31] ), .B(n159), .S0(n5053), .Y(
        n12538) );
  CLKMX2X2 U11538 ( .A(\I_cache/cache[0][31] ), .B(n159), .S0(n5094), .Y(
        n12539) );
  CLKMX2X2 U11539 ( .A(\I_cache/cache[7][30] ), .B(n140), .S0(n5317), .Y(
        n12540) );
  CLKMX2X2 U11540 ( .A(\I_cache/cache[6][30] ), .B(n140), .S0(n5362), .Y(
        n12541) );
  CLKMX2X2 U11541 ( .A(\I_cache/cache[5][30] ), .B(n140), .S0(n5225), .Y(
        n12542) );
  CLKMX2X2 U11542 ( .A(\I_cache/cache[4][30] ), .B(n140), .S0(n5271), .Y(
        n12543) );
  CLKMX2X2 U11543 ( .A(\I_cache/cache[3][30] ), .B(n140), .S0(n5138), .Y(
        n12544) );
  CLKMX2X2 U11544 ( .A(\I_cache/cache[2][30] ), .B(n140), .S0(n5184), .Y(
        n12545) );
  CLKMX2X2 U11545 ( .A(\I_cache/cache[1][30] ), .B(n140), .S0(n5047), .Y(
        n12546) );
  CLKMX2X2 U11546 ( .A(\I_cache/cache[0][30] ), .B(n140), .S0(n5094), .Y(
        n12547) );
  CLKMX2X2 U11547 ( .A(\I_cache/cache[6][29] ), .B(n6221), .S0(n5365), .Y(
        n12549) );
  CLKMX2X2 U11548 ( .A(\I_cache/cache[5][29] ), .B(n6221), .S0(n5228), .Y(
        n12550) );
  CLKMX2X2 U11549 ( .A(\I_cache/cache[4][29] ), .B(n6221), .S0(n5271), .Y(
        n12551) );
  CLKMX2X2 U11550 ( .A(\I_cache/cache[3][29] ), .B(n6221), .S0(n5138), .Y(
        n12552) );
  CLKMX2X2 U11551 ( .A(\I_cache/cache[2][29] ), .B(n6221), .S0(n5184), .Y(
        n12553) );
  CLKMX2X2 U11552 ( .A(\I_cache/cache[1][29] ), .B(n6221), .S0(n5049), .Y(
        n12554) );
  CLKMX2X2 U11553 ( .A(\I_cache/cache[7][28] ), .B(n6161), .S0(n5316), .Y(
        n12556) );
  CLKMX2X2 U11554 ( .A(\I_cache/cache[6][28] ), .B(n6161), .S0(n5359), .Y(
        n12557) );
  CLKMX2X2 U11555 ( .A(\I_cache/cache[5][28] ), .B(n6161), .S0(n5227), .Y(
        n12558) );
  CLKMX2X2 U11556 ( .A(\I_cache/cache[4][28] ), .B(n6161), .S0(n5270), .Y(
        n12559) );
  CLKMX2X2 U11557 ( .A(\I_cache/cache[3][28] ), .B(n6161), .S0(n5137), .Y(
        n12560) );
  CLKMX2X2 U11558 ( .A(\I_cache/cache[2][28] ), .B(n6161), .S0(n5183), .Y(
        n12561) );
  CLKMX2X2 U11559 ( .A(\I_cache/cache[1][28] ), .B(n6161), .S0(n5047), .Y(
        n12562) );
  CLKMX2X2 U11560 ( .A(\I_cache/cache[0][28] ), .B(n6161), .S0(n5093), .Y(
        n12563) );
  CLKMX2X2 U11561 ( .A(\I_cache/cache[7][27] ), .B(n11157), .S0(n5321), .Y(
        n12564) );
  CLKMX2X2 U11562 ( .A(\I_cache/cache[6][27] ), .B(n11157), .S0(n5364), .Y(
        n12565) );
  CLKMX2X2 U11563 ( .A(\I_cache/cache[5][27] ), .B(n11157), .S0(n5233), .Y(
        n12566) );
  CLKMX2X2 U11564 ( .A(\I_cache/cache[4][27] ), .B(n11157), .S0(n5276), .Y(
        n12567) );
  CLKMX2X2 U11565 ( .A(\I_cache/cache[3][27] ), .B(n11157), .S0(n5143), .Y(
        n12568) );
  CLKMX2X2 U11566 ( .A(\I_cache/cache[2][27] ), .B(n11157), .S0(n5189), .Y(
        n12569) );
  CLKMX2X2 U11567 ( .A(\I_cache/cache[1][27] ), .B(n11157), .S0(n5045), .Y(
        n12570) );
  CLKMX2X2 U11568 ( .A(\I_cache/cache[0][27] ), .B(n11157), .S0(n5098), .Y(
        n12571) );
  CLKMX2X2 U11569 ( .A(\I_cache/cache[7][26] ), .B(n9561), .S0(n5317), .Y(
        n12572) );
  CLKMX2X2 U11570 ( .A(\I_cache/cache[6][26] ), .B(n9561), .S0(n5359), .Y(
        n12573) );
  CLKMX2X2 U11571 ( .A(\I_cache/cache[5][26] ), .B(n9561), .S0(n5232), .Y(
        n12574) );
  CLKMX2X2 U11572 ( .A(\I_cache/cache[4][26] ), .B(n9561), .S0(n5271), .Y(
        n12575) );
  CLKMX2X2 U11573 ( .A(\I_cache/cache[3][26] ), .B(n9561), .S0(n5138), .Y(
        n12576) );
  CLKMX2X2 U11574 ( .A(\I_cache/cache[1][26] ), .B(n9561), .S0(n5050), .Y(
        n12578) );
  CLKMX2X2 U11575 ( .A(\I_cache/cache[0][26] ), .B(n9561), .S0(n5093), .Y(
        n12579) );
  CLKMX2X2 U11576 ( .A(\I_cache/cache[7][25] ), .B(n9809), .S0(n5319), .Y(
        n12580) );
  CLKMX2X2 U11577 ( .A(\I_cache/cache[6][25] ), .B(n9809), .S0(n5362), .Y(
        n12581) );
  CLKMX2X2 U11578 ( .A(\I_cache/cache[5][25] ), .B(n9809), .S0(n5230), .Y(
        n12582) );
  CLKMX2X2 U11579 ( .A(\I_cache/cache[4][25] ), .B(n9809), .S0(n5273), .Y(
        n12583) );
  CLKMX2X2 U11580 ( .A(\I_cache/cache[3][25] ), .B(n9809), .S0(n5141), .Y(
        n12584) );
  CLKMX2X2 U11581 ( .A(\I_cache/cache[2][25] ), .B(n9809), .S0(n5187), .Y(
        n12585) );
  CLKMX2X2 U11582 ( .A(\I_cache/cache[1][25] ), .B(n9809), .S0(n5048), .Y(
        n12586) );
  CLKMX2X2 U11583 ( .A(\I_cache/cache[0][25] ), .B(n9809), .S0(n5096), .Y(
        n12587) );
  CLKMX2X2 U11584 ( .A(\I_cache/cache[7][24] ), .B(n160), .S0(n5319), .Y(
        n12588) );
  CLKMX2X2 U11585 ( .A(\I_cache/cache[6][24] ), .B(n160), .S0(n5360), .Y(
        n12589) );
  CLKMX2X2 U11586 ( .A(\I_cache/cache[5][24] ), .B(n160), .S0(n5230), .Y(
        n12590) );
  CLKMX2X2 U11587 ( .A(\I_cache/cache[4][24] ), .B(n160), .S0(n5273), .Y(
        n12591) );
  CLKMX2X2 U11588 ( .A(\I_cache/cache[3][24] ), .B(n160), .S0(n5141), .Y(
        n12592) );
  CLKMX2X2 U11589 ( .A(\I_cache/cache[2][24] ), .B(n160), .S0(n5187), .Y(
        n12593) );
  CLKMX2X2 U11590 ( .A(\I_cache/cache[1][24] ), .B(n160), .S0(n5052), .Y(
        n12594) );
  CLKMX2X2 U11591 ( .A(\I_cache/cache[0][24] ), .B(n160), .S0(n5095), .Y(
        n12595) );
  CLKMX2X2 U11592 ( .A(\I_cache/cache[7][23] ), .B(n9829), .S0(n5320), .Y(
        n12596) );
  CLKMX2X2 U11593 ( .A(\I_cache/cache[6][23] ), .B(n9829), .S0(n5361), .Y(
        n12597) );
  CLKMX2X2 U11594 ( .A(\I_cache/cache[5][23] ), .B(n9829), .S0(n5231), .Y(
        n12598) );
  CLKMX2X2 U11595 ( .A(\I_cache/cache[4][23] ), .B(n9829), .S0(n5274), .Y(
        n12599) );
  CLKMX2X2 U11596 ( .A(\I_cache/cache[3][23] ), .B(n9829), .S0(n5142), .Y(
        n12600) );
  CLKMX2X2 U11597 ( .A(\I_cache/cache[2][23] ), .B(n9829), .S0(n5188), .Y(
        n12601) );
  CLKMX2X2 U11598 ( .A(\I_cache/cache[1][23] ), .B(n9829), .S0(n5048), .Y(
        n12602) );
  CLKMX2X2 U11599 ( .A(\I_cache/cache[0][23] ), .B(n9829), .S0(n5096), .Y(
        n12603) );
  CLKMX2X2 U11600 ( .A(\I_cache/cache[7][22] ), .B(n9865), .S0(n5318), .Y(
        n12604) );
  CLKMX2X2 U11601 ( .A(\I_cache/cache[6][22] ), .B(n9865), .S0(n5365), .Y(
        n12605) );
  CLKMX2X2 U11602 ( .A(\I_cache/cache[5][22] ), .B(n9865), .S0(n5231), .Y(
        n12606) );
  CLKMX2X2 U11603 ( .A(\I_cache/cache[4][22] ), .B(n9865), .S0(n5274), .Y(
        n12607) );
  CLKMX2X2 U11604 ( .A(\I_cache/cache[3][22] ), .B(n9865), .S0(n5142), .Y(
        n12608) );
  CLKMX2X2 U11605 ( .A(\I_cache/cache[2][22] ), .B(n9865), .S0(n5188), .Y(
        n12609) );
  CLKMX2X2 U11606 ( .A(\I_cache/cache[1][22] ), .B(n9865), .S0(n5052), .Y(
        n12610) );
  CLKMX2X2 U11607 ( .A(\I_cache/cache[0][22] ), .B(n9865), .S0(n5095), .Y(
        n12611) );
  CLKMX2X2 U11608 ( .A(\I_cache/cache[7][21] ), .B(n9849), .S0(n5321), .Y(
        n12612) );
  CLKMX2X2 U11609 ( .A(\I_cache/cache[6][21] ), .B(n9849), .S0(n5361), .Y(
        n12613) );
  CLKMX2X2 U11610 ( .A(\I_cache/cache[5][21] ), .B(n9849), .S0(n5231), .Y(
        n12614) );
  CLKMX2X2 U11611 ( .A(\I_cache/cache[4][21] ), .B(n9849), .S0(n5274), .Y(
        n12615) );
  CLKMX2X2 U11612 ( .A(\I_cache/cache[3][21] ), .B(n9849), .S0(n5142), .Y(
        n12616) );
  CLKMX2X2 U11613 ( .A(\I_cache/cache[2][21] ), .B(n9849), .S0(n5188), .Y(
        n12617) );
  CLKMX2X2 U11614 ( .A(\I_cache/cache[1][21] ), .B(n9849), .S0(n5052), .Y(
        n12618) );
  CLKMX2X2 U11615 ( .A(\I_cache/cache[0][21] ), .B(n9849), .S0(n5096), .Y(
        n12619) );
  CLKMX2X2 U11616 ( .A(\I_cache/cache[7][20] ), .B(n9619), .S0(n5314), .Y(
        n12620) );
  CLKMX2X2 U11617 ( .A(\I_cache/cache[6][20] ), .B(n9619), .S0(n5360), .Y(
        n12621) );
  CLKMX2X2 U11618 ( .A(\I_cache/cache[5][20] ), .B(n9619), .S0(n5225), .Y(
        n12622) );
  CLKMX2X2 U11619 ( .A(\I_cache/cache[4][20] ), .B(n9619), .S0(n5270), .Y(
        n12623) );
  CLKMX2X2 U11620 ( .A(\I_cache/cache[3][20] ), .B(n9619), .S0(n5135), .Y(
        n12624) );
  CLKMX2X2 U11621 ( .A(\I_cache/cache[2][20] ), .B(n9619), .S0(n5181), .Y(
        n12625) );
  CLKMX2X2 U11622 ( .A(\I_cache/cache[1][20] ), .B(n9619), .S0(n5045), .Y(
        n12626) );
  CLKMX2X2 U11623 ( .A(\I_cache/cache[0][20] ), .B(n9619), .S0(n5091), .Y(
        n12627) );
  CLKMX2X2 U11624 ( .A(\I_cache/cache[7][19] ), .B(n11116), .S0(n5317), .Y(
        n12628) );
  CLKMX2X2 U11625 ( .A(\I_cache/cache[6][19] ), .B(n11116), .S0(n5362), .Y(
        n12629) );
  CLKMX2X2 U11626 ( .A(\I_cache/cache[5][19] ), .B(n11116), .S0(n5230), .Y(
        n12630) );
  CLKMX2X2 U11627 ( .A(\I_cache/cache[4][19] ), .B(n11116), .S0(n5275), .Y(
        n12631) );
  CLKMX2X2 U11628 ( .A(\I_cache/cache[3][19] ), .B(n11116), .S0(n5143), .Y(
        n12632) );
  CLKMX2X2 U11629 ( .A(\I_cache/cache[2][19] ), .B(n11116), .S0(n5186), .Y(
        n12633) );
  CLKMX2X2 U11630 ( .A(\I_cache/cache[1][19] ), .B(n11116), .S0(n5047), .Y(
        n12634) );
  CLKMX2X2 U11631 ( .A(\I_cache/cache[0][19] ), .B(n11116), .S0(n5094), .Y(
        n12635) );
  CLKMX2X2 U11632 ( .A(\I_cache/cache[7][18] ), .B(n163), .S0(n5315), .Y(
        n12636) );
  CLKMX2X2 U11633 ( .A(\I_cache/cache[6][18] ), .B(n163), .S0(n5364), .Y(
        n12637) );
  CLKMX2X2 U11634 ( .A(\I_cache/cache[5][18] ), .B(n163), .S0(n5226), .Y(
        n12638) );
  CLKMX2X2 U11635 ( .A(\I_cache/cache[4][18] ), .B(n163), .S0(n5269), .Y(
        n12639) );
  CLKMX2X2 U11636 ( .A(\I_cache/cache[3][18] ), .B(n163), .S0(n5136), .Y(
        n12640) );
  CLKMX2X2 U11637 ( .A(\I_cache/cache[2][18] ), .B(n163), .S0(n5182), .Y(
        n12641) );
  CLKMX2X2 U11638 ( .A(\I_cache/cache[1][18] ), .B(n163), .S0(n5053), .Y(
        n12642) );
  CLKMX2X2 U11639 ( .A(\I_cache/cache[0][18] ), .B(n163), .S0(n5092), .Y(
        n12643) );
  CLKMX2X2 U11640 ( .A(\I_cache/cache[7][17] ), .B(n10157), .S0(n5322), .Y(
        n12644) );
  CLKMX2X2 U11641 ( .A(\I_cache/cache[6][17] ), .B(n10157), .S0(n5358), .Y(
        n12645) );
  CLKMX2X2 U11642 ( .A(\I_cache/cache[5][17] ), .B(n10157), .S0(n5229), .Y(
        n12646) );
  CLKMX2X2 U11643 ( .A(\I_cache/cache[4][17] ), .B(n10157), .S0(n5277), .Y(
        n12647) );
  CLKMX2X2 U11644 ( .A(\I_cache/cache[3][17] ), .B(n10157), .S0(n5142), .Y(
        n12648) );
  CLKMX2X2 U11645 ( .A(\I_cache/cache[2][17] ), .B(n10157), .S0(n5189), .Y(
        n12649) );
  CLKMX2X2 U11646 ( .A(\I_cache/cache[1][17] ), .B(n10157), .S0(n5049), .Y(
        n12650) );
  CLKMX2X2 U11647 ( .A(\I_cache/cache[0][17] ), .B(n10157), .S0(n5099), .Y(
        n12651) );
  CLKMX2X2 U11648 ( .A(\I_cache/cache[7][16] ), .B(n9717), .S0(n5315), .Y(
        n12652) );
  CLKMX2X2 U11649 ( .A(\I_cache/cache[6][16] ), .B(n9717), .S0(n5366), .Y(
        n12653) );
  CLKMX2X2 U11650 ( .A(\I_cache/cache[5][16] ), .B(n9717), .S0(n5226), .Y(
        n12654) );
  CLKMX2X2 U11651 ( .A(\I_cache/cache[4][16] ), .B(n9717), .S0(n5269), .Y(
        n12655) );
  CLKMX2X2 U11652 ( .A(\I_cache/cache[3][16] ), .B(n9717), .S0(n5136), .Y(
        n12656) );
  CLKMX2X2 U11653 ( .A(\I_cache/cache[2][16] ), .B(n9717), .S0(n5182), .Y(
        n12657) );
  CLKMX2X2 U11654 ( .A(\I_cache/cache[1][16] ), .B(n9717), .S0(n5047), .Y(
        n12658) );
  CLKMX2X2 U11655 ( .A(\I_cache/cache[0][16] ), .B(n9717), .S0(n5092), .Y(
        n12659) );
  MX2XL U11656 ( .A(\I_cache/cache[7][15] ), .B(n9643), .S0(n5314), .Y(n12660)
         );
  CLKMX2X2 U11657 ( .A(\I_cache/cache[6][14] ), .B(n9594), .S0(n5361), .Y(
        n12669) );
  CLKMX2X2 U11658 ( .A(\I_cache/cache[5][14] ), .B(n9594), .S0(n5225), .Y(
        n12670) );
  CLKMX2X2 U11659 ( .A(\I_cache/cache[4][14] ), .B(n9594), .S0(n5274), .Y(
        n12671) );
  CLKMX2X2 U11660 ( .A(\I_cache/cache[3][14] ), .B(n9594), .S0(n5135), .Y(
        n12672) );
  CLKMX2X2 U11661 ( .A(\I_cache/cache[2][14] ), .B(n9594), .S0(n5181), .Y(
        n12673) );
  CLKMX2X2 U11662 ( .A(\I_cache/cache[1][14] ), .B(n9594), .S0(n5046), .Y(
        n12674) );
  CLKMX2X2 U11663 ( .A(\I_cache/cache[0][14] ), .B(n9594), .S0(n5091), .Y(
        n12675) );
  CLKMX2X2 U11664 ( .A(\I_cache/cache[6][13] ), .B(n9693), .S0(n5365), .Y(
        n12677) );
  CLKMX2X2 U11665 ( .A(\I_cache/cache[3][13] ), .B(n9693), .S0(n5136), .Y(
        n12680) );
  CLKMX2X2 U11666 ( .A(\I_cache/cache[2][13] ), .B(n9693), .S0(n5182), .Y(
        n12681) );
  CLKMX2X2 U11667 ( .A(\I_cache/cache[1][13] ), .B(n9693), .S0(n5050), .Y(
        n12682) );
  CLKMX2X2 U11668 ( .A(\I_cache/cache[0][13] ), .B(n9693), .S0(n5092), .Y(
        n12683) );
  CLKMX2X2 U11669 ( .A(\I_cache/cache[6][12] ), .B(n9764), .S0(n5360), .Y(
        n12685) );
  CLKMX2X2 U11670 ( .A(\I_cache/cache[5][12] ), .B(n9764), .S0(n5230), .Y(
        n12686) );
  CLKMX2X2 U11671 ( .A(\I_cache/cache[4][12] ), .B(n9764), .S0(n5273), .Y(
        n12687) );
  CLKMX2X2 U11672 ( .A(\I_cache/cache[3][12] ), .B(n9764), .S0(n5141), .Y(
        n12688) );
  CLKMX2X2 U11673 ( .A(\I_cache/cache[2][12] ), .B(n9764), .S0(n5187), .Y(
        n12689) );
  CLKMX2X2 U11674 ( .A(\I_cache/cache[1][12] ), .B(n9764), .S0(n5049), .Y(
        n12690) );
  CLKMX2X2 U11675 ( .A(\I_cache/cache[0][12] ), .B(n9764), .S0(n5095), .Y(
        n12691) );
  CLKMX2X2 U11676 ( .A(\I_cache/cache[6][11] ), .B(n9741), .S0(n5365), .Y(
        n12693) );
  CLKMX2X2 U11677 ( .A(\I_cache/cache[4][11] ), .B(n9741), .S0(n5269), .Y(
        n12695) );
  CLKMX2X2 U11678 ( .A(\I_cache/cache[2][11] ), .B(n9741), .S0(n5182), .Y(
        n12697) );
  CLKMX2X2 U11679 ( .A(\I_cache/cache[0][11] ), .B(n9741), .S0(n5095), .Y(
        n12699) );
  CLKMX2X2 U11680 ( .A(\I_cache/cache[0][10] ), .B(n10044), .S0(n5091), .Y(
        n12707) );
  CLKMX2X2 U11681 ( .A(\I_cache/cache[7][5] ), .B(n9914), .S0(n5315), .Y(
        n12740) );
  CLKMX2X2 U11682 ( .A(\I_cache/cache[6][5] ), .B(n9914), .S0(n5363), .Y(
        n12741) );
  CLKMX2X2 U11683 ( .A(\I_cache/cache[5][5] ), .B(n9914), .S0(n5228), .Y(
        n12742) );
  CLKMX2X2 U11684 ( .A(\I_cache/cache[4][5] ), .B(n9914), .S0(n5275), .Y(
        n12743) );
  CLKMX2X2 U11685 ( .A(\I_cache/cache[3][5] ), .B(n9914), .S0(n5139), .Y(
        n12744) );
  CLKMX2X2 U11686 ( .A(\I_cache/cache[2][5] ), .B(n9914), .S0(n5185), .Y(
        n12745) );
  CLKMX2X2 U11687 ( .A(\I_cache/cache[1][5] ), .B(n9914), .S0(n5052), .Y(
        n12746) );
  CLKMX2X2 U11688 ( .A(\I_cache/cache[0][5] ), .B(n9914), .S0(n5096), .Y(
        n12747) );
  CLKMX2X2 U11689 ( .A(\I_cache/cache[6][2] ), .B(n11102), .S0(n5360), .Y(
        n12765) );
  CLKMX2X2 U11690 ( .A(\I_cache/cache[4][2] ), .B(n11102), .S0(n5277), .Y(
        n12767) );
  CLKMX2X2 U11691 ( .A(\I_cache/cache[3][2] ), .B(n11102), .S0(n5140), .Y(
        n12768) );
  CLKMX2X2 U11692 ( .A(\I_cache/cache[2][2] ), .B(n11102), .S0(n5186), .Y(
        n12769) );
  CLKMX2X2 U11693 ( .A(\I_cache/cache[1][2] ), .B(n11102), .S0(n5046), .Y(
        n12770) );
  CLKMX2X2 U11694 ( .A(\I_cache/cache[0][2] ), .B(n11102), .S0(n5093), .Y(
        n12771) );
  MXI2X1 U11695 ( .A(net112764), .B(\i_MIPS/n222 ), .S0(n213), .Y(
        \i_MIPS/n505 ) );
  MXI2XL U11696 ( .A(\i_MIPS/n303 ), .B(n8429), .S0(n210), .Y(\i_MIPS/n431 )
         );
  CLKMX2X2 U11697 ( .A(n5482), .B(\i_MIPS/Register/register[0][23] ), .S0(
        n5621), .Y(\i_MIPS/Register/n1131 ) );
  CLKMX2X2 U11698 ( .A(n5491), .B(\i_MIPS/Register/register[0][5] ), .S0(n5620), .Y(\i_MIPS/Register/n1113 ) );
  CLKMX2X2 U11699 ( .A(n5487), .B(\i_MIPS/Register/register[0][4] ), .S0(n5621), .Y(\i_MIPS/Register/n1112 ) );
  CLKMX2X2 U11700 ( .A(n5479), .B(\i_MIPS/Register/register[0][2] ), .S0(n5620), .Y(\i_MIPS/Register/n1110 ) );
  CLKMX2X2 U11701 ( .A(n5477), .B(\i_MIPS/Register/register[0][1] ), .S0(
        \i_MIPS/Register/n147 ), .Y(\i_MIPS/Register/n1109 ) );
  CLKMX2X2 U11702 ( .A(n5484), .B(\i_MIPS/Register/register[0][0] ), .S0(
        \i_MIPS/Register/n147 ), .Y(\i_MIPS/Register/n1108 ) );
  CLKMX2X2 U11703 ( .A(n5462), .B(\i_MIPS/Register/register[1][30] ), .S0(
        n5618), .Y(\i_MIPS/Register/n1106 ) );
  CLKMX2X2 U11704 ( .A(n5440), .B(\i_MIPS/Register/register[1][29] ), .S0(
        n5619), .Y(\i_MIPS/Register/n1105 ) );
  CLKMX2X2 U11705 ( .A(n5460), .B(\i_MIPS/Register/register[1][24] ), .S0(
        n5618), .Y(\i_MIPS/Register/n1100 ) );
  CLKMX2X2 U11706 ( .A(n5437), .B(\i_MIPS/Register/register[1][21] ), .S0(
        n5619), .Y(\i_MIPS/Register/n1097 ) );
  CLKMX2X2 U11707 ( .A(n5434), .B(\i_MIPS/Register/register[1][20] ), .S0(
        \i_MIPS/Register/n146 ), .Y(\i_MIPS/Register/n1096 ) );
  CLKMX2X2 U11708 ( .A(n5442), .B(\i_MIPS/Register/register[1][9] ), .S0(
        \i_MIPS/Register/n146 ), .Y(\i_MIPS/Register/n1085 ) );
  CLKMX2X2 U11709 ( .A(n5462), .B(\i_MIPS/Register/register[2][30] ), .S0(
        n5616), .Y(\i_MIPS/Register/n1074 ) );
  CLKMX2X2 U11710 ( .A(n5440), .B(\i_MIPS/Register/register[2][29] ), .S0(
        n5617), .Y(\i_MIPS/Register/n1073 ) );
  CLKMX2X2 U11711 ( .A(n5460), .B(\i_MIPS/Register/register[2][24] ), .S0(
        n5616), .Y(\i_MIPS/Register/n1068 ) );
  CLKMX2X2 U11712 ( .A(n5437), .B(\i_MIPS/Register/register[2][21] ), .S0(
        n5617), .Y(\i_MIPS/Register/n1065 ) );
  CLKMX2X2 U11713 ( .A(n5434), .B(\i_MIPS/Register/register[2][20] ), .S0(
        \i_MIPS/Register/n145 ), .Y(\i_MIPS/Register/n1064 ) );
  CLKMX2X2 U11714 ( .A(n5442), .B(\i_MIPS/Register/register[2][9] ), .S0(
        \i_MIPS/Register/n145 ), .Y(\i_MIPS/Register/n1053 ) );
  CLKMX2X2 U11715 ( .A(n5462), .B(\i_MIPS/Register/register[3][30] ), .S0(
        n5614), .Y(\i_MIPS/Register/n1042 ) );
  CLKMX2X2 U11716 ( .A(n5440), .B(\i_MIPS/Register/register[3][29] ), .S0(
        n5615), .Y(\i_MIPS/Register/n1041 ) );
  CLKMX2X2 U11717 ( .A(n5460), .B(\i_MIPS/Register/register[3][24] ), .S0(
        n5614), .Y(\i_MIPS/Register/n1036 ) );
  CLKMX2X2 U11718 ( .A(n5437), .B(\i_MIPS/Register/register[3][21] ), .S0(
        n5615), .Y(\i_MIPS/Register/n1033 ) );
  CLKMX2X2 U11719 ( .A(n5434), .B(\i_MIPS/Register/register[3][20] ), .S0(
        \i_MIPS/Register/n144 ), .Y(\i_MIPS/Register/n1032 ) );
  CLKMX2X2 U11720 ( .A(n5442), .B(\i_MIPS/Register/register[3][9] ), .S0(
        \i_MIPS/Register/n144 ), .Y(\i_MIPS/Register/n1021 ) );
  CLKMX2X2 U11721 ( .A(n5462), .B(\i_MIPS/Register/register[4][30] ), .S0(
        n5612), .Y(\i_MIPS/Register/n1010 ) );
  CLKMX2X2 U11722 ( .A(n5440), .B(\i_MIPS/Register/register[4][29] ), .S0(
        n5613), .Y(\i_MIPS/Register/n1009 ) );
  CLKMX2X2 U11723 ( .A(n5460), .B(\i_MIPS/Register/register[4][24] ), .S0(
        n5612), .Y(\i_MIPS/Register/n1004 ) );
  CLKMX2X2 U11724 ( .A(n5437), .B(\i_MIPS/Register/register[4][21] ), .S0(
        n5613), .Y(\i_MIPS/Register/n1001 ) );
  CLKMX2X2 U11725 ( .A(n5434), .B(\i_MIPS/Register/register[4][20] ), .S0(
        \i_MIPS/Register/n143 ), .Y(\i_MIPS/Register/n1000 ) );
  CLKMX2X2 U11726 ( .A(n5442), .B(\i_MIPS/Register/register[4][9] ), .S0(
        \i_MIPS/Register/n143 ), .Y(\i_MIPS/Register/n989 ) );
  CLKMX2X2 U11727 ( .A(n5462), .B(\i_MIPS/Register/register[5][30] ), .S0(
        n5610), .Y(\i_MIPS/Register/n978 ) );
  CLKMX2X2 U11728 ( .A(n5440), .B(\i_MIPS/Register/register[5][29] ), .S0(
        n5611), .Y(\i_MIPS/Register/n977 ) );
  CLKMX2X2 U11729 ( .A(n5460), .B(\i_MIPS/Register/register[5][24] ), .S0(
        n5610), .Y(\i_MIPS/Register/n972 ) );
  CLKMX2X2 U11730 ( .A(n5437), .B(\i_MIPS/Register/register[5][21] ), .S0(
        n5611), .Y(\i_MIPS/Register/n969 ) );
  CLKMX2X2 U11731 ( .A(n5434), .B(\i_MIPS/Register/register[5][20] ), .S0(
        \i_MIPS/Register/n142 ), .Y(\i_MIPS/Register/n968 ) );
  CLKMX2X2 U11732 ( .A(n5442), .B(\i_MIPS/Register/register[5][9] ), .S0(
        \i_MIPS/Register/n142 ), .Y(\i_MIPS/Register/n957 ) );
  CLKMX2X2 U11733 ( .A(n5462), .B(\i_MIPS/Register/register[6][30] ), .S0(
        n5608), .Y(\i_MIPS/Register/n946 ) );
  CLKMX2X2 U11734 ( .A(n5440), .B(\i_MIPS/Register/register[6][29] ), .S0(
        n5609), .Y(\i_MIPS/Register/n945 ) );
  CLKMX2X2 U11735 ( .A(n5460), .B(\i_MIPS/Register/register[6][24] ), .S0(
        n5608), .Y(\i_MIPS/Register/n940 ) );
  CLKMX2X2 U11736 ( .A(n5437), .B(\i_MIPS/Register/register[6][21] ), .S0(
        n5609), .Y(\i_MIPS/Register/n937 ) );
  CLKMX2X2 U11737 ( .A(n5434), .B(\i_MIPS/Register/register[6][20] ), .S0(
        \i_MIPS/Register/n141 ), .Y(\i_MIPS/Register/n936 ) );
  CLKMX2X2 U11738 ( .A(n5442), .B(\i_MIPS/Register/register[6][9] ), .S0(
        \i_MIPS/Register/n141 ), .Y(\i_MIPS/Register/n925 ) );
  CLKMX2X2 U11739 ( .A(n5463), .B(\i_MIPS/Register/register[7][30] ), .S0(
        n5606), .Y(\i_MIPS/Register/n914 ) );
  CLKMX2X2 U11740 ( .A(n5441), .B(\i_MIPS/Register/register[7][29] ), .S0(
        n5607), .Y(\i_MIPS/Register/n913 ) );
  CLKMX2X2 U11741 ( .A(n5461), .B(\i_MIPS/Register/register[7][24] ), .S0(
        n5606), .Y(\i_MIPS/Register/n908 ) );
  CLKMX2X2 U11742 ( .A(n5438), .B(\i_MIPS/Register/register[7][21] ), .S0(
        n5607), .Y(\i_MIPS/Register/n905 ) );
  CLKMX2X2 U11743 ( .A(n5435), .B(\i_MIPS/Register/register[7][20] ), .S0(
        \i_MIPS/Register/n139 ), .Y(\i_MIPS/Register/n904 ) );
  CLKMX2X2 U11744 ( .A(n5443), .B(\i_MIPS/Register/register[7][9] ), .S0(
        \i_MIPS/Register/n139 ), .Y(\i_MIPS/Register/n893 ) );
  CLKMX2X2 U11745 ( .A(n5462), .B(\i_MIPS/Register/register[8][30] ), .S0(
        n5604), .Y(\i_MIPS/Register/n882 ) );
  CLKMX2X2 U11746 ( .A(n5440), .B(\i_MIPS/Register/register[8][29] ), .S0(
        n5605), .Y(\i_MIPS/Register/n881 ) );
  CLKMX2X2 U11747 ( .A(n5460), .B(\i_MIPS/Register/register[8][24] ), .S0(
        n5604), .Y(\i_MIPS/Register/n876 ) );
  CLKMX2X2 U11748 ( .A(n5437), .B(\i_MIPS/Register/register[8][21] ), .S0(
        n5605), .Y(\i_MIPS/Register/n873 ) );
  CLKMX2X2 U11749 ( .A(n5434), .B(\i_MIPS/Register/register[8][20] ), .S0(
        \i_MIPS/Register/n138 ), .Y(\i_MIPS/Register/n872 ) );
  CLKMX2X2 U11750 ( .A(n5442), .B(\i_MIPS/Register/register[8][9] ), .S0(
        \i_MIPS/Register/n138 ), .Y(\i_MIPS/Register/n861 ) );
  CLKMX2X2 U11751 ( .A(n5462), .B(\i_MIPS/Register/register[9][30] ), .S0(
        n5602), .Y(\i_MIPS/Register/n850 ) );
  CLKMX2X2 U11752 ( .A(n5440), .B(\i_MIPS/Register/register[9][29] ), .S0(
        n5603), .Y(\i_MIPS/Register/n849 ) );
  CLKMX2X2 U11753 ( .A(n5460), .B(\i_MIPS/Register/register[9][24] ), .S0(
        n5602), .Y(\i_MIPS/Register/n844 ) );
  CLKMX2X2 U11754 ( .A(n5437), .B(\i_MIPS/Register/register[9][21] ), .S0(
        n5603), .Y(\i_MIPS/Register/n841 ) );
  CLKMX2X2 U11755 ( .A(n5434), .B(\i_MIPS/Register/register[9][20] ), .S0(
        \i_MIPS/Register/n137 ), .Y(\i_MIPS/Register/n840 ) );
  CLKMX2X2 U11756 ( .A(n5442), .B(\i_MIPS/Register/register[9][9] ), .S0(
        \i_MIPS/Register/n137 ), .Y(\i_MIPS/Register/n829 ) );
  CLKMX2X2 U11757 ( .A(n5462), .B(\i_MIPS/Register/register[10][30] ), .S0(
        n5600), .Y(\i_MIPS/Register/n818 ) );
  CLKMX2X2 U11758 ( .A(n5440), .B(\i_MIPS/Register/register[10][29] ), .S0(
        n5601), .Y(\i_MIPS/Register/n817 ) );
  CLKMX2X2 U11759 ( .A(n5460), .B(\i_MIPS/Register/register[10][24] ), .S0(
        n5600), .Y(\i_MIPS/Register/n812 ) );
  CLKMX2X2 U11760 ( .A(n5437), .B(\i_MIPS/Register/register[10][21] ), .S0(
        n5601), .Y(\i_MIPS/Register/n809 ) );
  CLKMX2X2 U11761 ( .A(n5434), .B(\i_MIPS/Register/register[10][20] ), .S0(
        \i_MIPS/Register/n136 ), .Y(\i_MIPS/Register/n808 ) );
  CLKMX2X2 U11762 ( .A(n5442), .B(\i_MIPS/Register/register[10][9] ), .S0(
        \i_MIPS/Register/n136 ), .Y(\i_MIPS/Register/n797 ) );
  CLKMX2X2 U11763 ( .A(n5463), .B(\i_MIPS/Register/register[11][30] ), .S0(
        n5598), .Y(\i_MIPS/Register/n786 ) );
  CLKMX2X2 U11764 ( .A(n5440), .B(\i_MIPS/Register/register[11][29] ), .S0(
        n5599), .Y(\i_MIPS/Register/n785 ) );
  CLKMX2X2 U11765 ( .A(n5460), .B(\i_MIPS/Register/register[11][24] ), .S0(
        n5598), .Y(\i_MIPS/Register/n780 ) );
  CLKMX2X2 U11766 ( .A(n5437), .B(\i_MIPS/Register/register[11][21] ), .S0(
        n5599), .Y(\i_MIPS/Register/n777 ) );
  CLKMX2X2 U11767 ( .A(n5434), .B(\i_MIPS/Register/register[11][20] ), .S0(
        \i_MIPS/Register/n135 ), .Y(\i_MIPS/Register/n776 ) );
  CLKMX2X2 U11768 ( .A(n5442), .B(\i_MIPS/Register/register[11][9] ), .S0(
        \i_MIPS/Register/n135 ), .Y(\i_MIPS/Register/n765 ) );
  CLKMX2X2 U11769 ( .A(n5462), .B(\i_MIPS/Register/register[12][30] ), .S0(
        n5596), .Y(\i_MIPS/Register/n754 ) );
  CLKMX2X2 U11770 ( .A(n5440), .B(\i_MIPS/Register/register[12][29] ), .S0(
        n5597), .Y(\i_MIPS/Register/n753 ) );
  CLKMX2X2 U11771 ( .A(n5460), .B(\i_MIPS/Register/register[12][24] ), .S0(
        n5596), .Y(\i_MIPS/Register/n748 ) );
  CLKMX2X2 U11772 ( .A(n5437), .B(\i_MIPS/Register/register[12][21] ), .S0(
        n5597), .Y(\i_MIPS/Register/n745 ) );
  CLKMX2X2 U11773 ( .A(n5434), .B(\i_MIPS/Register/register[12][20] ), .S0(
        \i_MIPS/Register/n134 ), .Y(\i_MIPS/Register/n744 ) );
  CLKMX2X2 U11774 ( .A(n5442), .B(\i_MIPS/Register/register[12][9] ), .S0(
        \i_MIPS/Register/n134 ), .Y(\i_MIPS/Register/n733 ) );
  CLKMX2X2 U11775 ( .A(n5462), .B(\i_MIPS/Register/register[13][30] ), .S0(
        n5594), .Y(\i_MIPS/Register/n722 ) );
  CLKMX2X2 U11776 ( .A(n5440), .B(\i_MIPS/Register/register[13][29] ), .S0(
        n5595), .Y(\i_MIPS/Register/n721 ) );
  CLKMX2X2 U11777 ( .A(n5460), .B(\i_MIPS/Register/register[13][24] ), .S0(
        n5594), .Y(\i_MIPS/Register/n716 ) );
  CLKMX2X2 U11778 ( .A(n5437), .B(\i_MIPS/Register/register[13][21] ), .S0(
        n5595), .Y(\i_MIPS/Register/n713 ) );
  CLKMX2X2 U11779 ( .A(n5434), .B(\i_MIPS/Register/register[13][20] ), .S0(
        \i_MIPS/Register/n133 ), .Y(\i_MIPS/Register/n712 ) );
  CLKMX2X2 U11780 ( .A(n5442), .B(\i_MIPS/Register/register[13][9] ), .S0(
        \i_MIPS/Register/n133 ), .Y(\i_MIPS/Register/n701 ) );
  CLKMX2X2 U11781 ( .A(n5462), .B(\i_MIPS/Register/register[14][30] ), .S0(
        n5592), .Y(\i_MIPS/Register/n690 ) );
  CLKMX2X2 U11782 ( .A(n5440), .B(\i_MIPS/Register/register[14][29] ), .S0(
        n5593), .Y(\i_MIPS/Register/n689 ) );
  CLKMX2X2 U11783 ( .A(n5460), .B(\i_MIPS/Register/register[14][24] ), .S0(
        n5592), .Y(\i_MIPS/Register/n684 ) );
  CLKMX2X2 U11784 ( .A(n5437), .B(\i_MIPS/Register/register[14][21] ), .S0(
        n5593), .Y(\i_MIPS/Register/n681 ) );
  CLKMX2X2 U11785 ( .A(n5434), .B(\i_MIPS/Register/register[14][20] ), .S0(
        \i_MIPS/Register/n132 ), .Y(\i_MIPS/Register/n680 ) );
  CLKMX2X2 U11786 ( .A(n5442), .B(\i_MIPS/Register/register[14][9] ), .S0(
        \i_MIPS/Register/n132 ), .Y(\i_MIPS/Register/n669 ) );
  CLKMX2X2 U11787 ( .A(n5463), .B(\i_MIPS/Register/register[15][30] ), .S0(
        n5590), .Y(\i_MIPS/Register/n658 ) );
  CLKMX2X2 U11788 ( .A(n5441), .B(\i_MIPS/Register/register[15][29] ), .S0(
        n5591), .Y(\i_MIPS/Register/n657 ) );
  CLKMX2X2 U11789 ( .A(n5461), .B(\i_MIPS/Register/register[15][24] ), .S0(
        n5590), .Y(\i_MIPS/Register/n652 ) );
  CLKMX2X2 U11790 ( .A(n5438), .B(\i_MIPS/Register/register[15][21] ), .S0(
        n5591), .Y(\i_MIPS/Register/n649 ) );
  CLKMX2X2 U11791 ( .A(n5435), .B(\i_MIPS/Register/register[15][20] ), .S0(
        \i_MIPS/Register/n130 ), .Y(\i_MIPS/Register/n648 ) );
  CLKMX2X2 U11792 ( .A(n5443), .B(\i_MIPS/Register/register[15][9] ), .S0(
        \i_MIPS/Register/n130 ), .Y(\i_MIPS/Register/n637 ) );
  CLKMX2X2 U11793 ( .A(n5463), .B(\i_MIPS/Register/register[16][30] ), .S0(
        n5588), .Y(\i_MIPS/Register/n626 ) );
  CLKMX2X2 U11794 ( .A(n5441), .B(\i_MIPS/Register/register[16][29] ), .S0(
        n5589), .Y(\i_MIPS/Register/n625 ) );
  CLKMX2X2 U11795 ( .A(n5461), .B(\i_MIPS/Register/register[16][24] ), .S0(
        n5588), .Y(\i_MIPS/Register/n620 ) );
  CLKMX2X2 U11796 ( .A(n5438), .B(\i_MIPS/Register/register[16][21] ), .S0(
        n5589), .Y(\i_MIPS/Register/n617 ) );
  CLKMX2X2 U11797 ( .A(n5435), .B(\i_MIPS/Register/register[16][20] ), .S0(
        \i_MIPS/Register/n129 ), .Y(\i_MIPS/Register/n616 ) );
  CLKMX2X2 U11798 ( .A(n5443), .B(\i_MIPS/Register/register[16][9] ), .S0(
        \i_MIPS/Register/n129 ), .Y(\i_MIPS/Register/n605 ) );
  CLKMX2X2 U11799 ( .A(n5463), .B(\i_MIPS/Register/register[17][30] ), .S0(
        n5586), .Y(\i_MIPS/Register/n594 ) );
  CLKMX2X2 U11800 ( .A(n5441), .B(\i_MIPS/Register/register[17][29] ), .S0(
        n5587), .Y(\i_MIPS/Register/n593 ) );
  CLKMX2X2 U11801 ( .A(n5461), .B(\i_MIPS/Register/register[17][24] ), .S0(
        n5586), .Y(\i_MIPS/Register/n588 ) );
  CLKMX2X2 U11802 ( .A(n5438), .B(\i_MIPS/Register/register[17][21] ), .S0(
        n5587), .Y(\i_MIPS/Register/n585 ) );
  CLKMX2X2 U11803 ( .A(n5435), .B(\i_MIPS/Register/register[17][20] ), .S0(
        \i_MIPS/Register/n128 ), .Y(\i_MIPS/Register/n584 ) );
  CLKMX2X2 U11804 ( .A(n5443), .B(\i_MIPS/Register/register[17][9] ), .S0(
        \i_MIPS/Register/n128 ), .Y(\i_MIPS/Register/n573 ) );
  CLKMX2X2 U11805 ( .A(n5463), .B(\i_MIPS/Register/register[18][30] ), .S0(
        n5584), .Y(\i_MIPS/Register/n562 ) );
  CLKMX2X2 U11806 ( .A(n5441), .B(\i_MIPS/Register/register[18][29] ), .S0(
        n5585), .Y(\i_MIPS/Register/n561 ) );
  CLKMX2X2 U11807 ( .A(n5461), .B(\i_MIPS/Register/register[18][24] ), .S0(
        n5584), .Y(\i_MIPS/Register/n556 ) );
  CLKMX2X2 U11808 ( .A(n5438), .B(\i_MIPS/Register/register[18][21] ), .S0(
        n5585), .Y(\i_MIPS/Register/n553 ) );
  CLKMX2X2 U11809 ( .A(n5435), .B(\i_MIPS/Register/register[18][20] ), .S0(
        \i_MIPS/Register/n127 ), .Y(\i_MIPS/Register/n552 ) );
  CLKMX2X2 U11810 ( .A(n5443), .B(\i_MIPS/Register/register[18][9] ), .S0(
        \i_MIPS/Register/n127 ), .Y(\i_MIPS/Register/n541 ) );
  CLKMX2X2 U11811 ( .A(n5462), .B(\i_MIPS/Register/register[19][30] ), .S0(
        \i_MIPS/Register/n126 ), .Y(\i_MIPS/Register/n530 ) );
  CLKMX2X2 U11812 ( .A(n5440), .B(\i_MIPS/Register/register[19][29] ), .S0(
        n5582), .Y(\i_MIPS/Register/n529 ) );
  CLKMX2X2 U11813 ( .A(n5460), .B(\i_MIPS/Register/register[19][24] ), .S0(
        n5583), .Y(\i_MIPS/Register/n524 ) );
  CLKMX2X2 U11814 ( .A(n5437), .B(\i_MIPS/Register/register[19][21] ), .S0(
        n5582), .Y(\i_MIPS/Register/n521 ) );
  CLKMX2X2 U11815 ( .A(n5434), .B(\i_MIPS/Register/register[19][20] ), .S0(
        n5583), .Y(\i_MIPS/Register/n520 ) );
  CLKMX2X2 U11816 ( .A(n5442), .B(\i_MIPS/Register/register[19][9] ), .S0(
        \i_MIPS/Register/n126 ), .Y(\i_MIPS/Register/n509 ) );
  CLKMX2X2 U11817 ( .A(n5463), .B(\i_MIPS/Register/register[20][30] ), .S0(
        n5580), .Y(\i_MIPS/Register/n498 ) );
  CLKMX2X2 U11818 ( .A(n5441), .B(\i_MIPS/Register/register[20][29] ), .S0(
        n5581), .Y(\i_MIPS/Register/n497 ) );
  CLKMX2X2 U11819 ( .A(n5461), .B(\i_MIPS/Register/register[20][24] ), .S0(
        n5580), .Y(\i_MIPS/Register/n492 ) );
  CLKMX2X2 U11820 ( .A(n5438), .B(\i_MIPS/Register/register[20][21] ), .S0(
        n5581), .Y(\i_MIPS/Register/n489 ) );
  CLKMX2X2 U11821 ( .A(n5435), .B(\i_MIPS/Register/register[20][20] ), .S0(
        \i_MIPS/Register/n125 ), .Y(\i_MIPS/Register/n488 ) );
  CLKMX2X2 U11822 ( .A(n5443), .B(\i_MIPS/Register/register[20][9] ), .S0(
        \i_MIPS/Register/n125 ), .Y(\i_MIPS/Register/n477 ) );
  CLKMX2X2 U11823 ( .A(n5463), .B(\i_MIPS/Register/register[21][30] ), .S0(
        \i_MIPS/Register/n124 ), .Y(\i_MIPS/Register/n466 ) );
  CLKMX2X2 U11824 ( .A(n5441), .B(\i_MIPS/Register/register[21][29] ), .S0(
        n5578), .Y(\i_MIPS/Register/n465 ) );
  CLKMX2X2 U11825 ( .A(n5461), .B(\i_MIPS/Register/register[21][24] ), .S0(
        n5579), .Y(\i_MIPS/Register/n460 ) );
  CLKMX2X2 U11826 ( .A(n5438), .B(\i_MIPS/Register/register[21][21] ), .S0(
        n5578), .Y(\i_MIPS/Register/n457 ) );
  CLKMX2X2 U11827 ( .A(n5435), .B(\i_MIPS/Register/register[21][20] ), .S0(
        n5579), .Y(\i_MIPS/Register/n456 ) );
  CLKMX2X2 U11828 ( .A(n5443), .B(\i_MIPS/Register/register[21][9] ), .S0(
        \i_MIPS/Register/n124 ), .Y(\i_MIPS/Register/n445 ) );
  CLKMX2X2 U11829 ( .A(n5463), .B(\i_MIPS/Register/register[22][30] ), .S0(
        n5576), .Y(\i_MIPS/Register/n434 ) );
  CLKMX2X2 U11830 ( .A(n5441), .B(\i_MIPS/Register/register[22][29] ), .S0(
        n5577), .Y(\i_MIPS/Register/n433 ) );
  CLKMX2X2 U11831 ( .A(n5461), .B(\i_MIPS/Register/register[22][24] ), .S0(
        n5576), .Y(\i_MIPS/Register/n428 ) );
  CLKMX2X2 U11832 ( .A(n5438), .B(\i_MIPS/Register/register[22][21] ), .S0(
        n5577), .Y(\i_MIPS/Register/n425 ) );
  CLKMX2X2 U11833 ( .A(n5435), .B(\i_MIPS/Register/register[22][20] ), .S0(
        \i_MIPS/Register/n123 ), .Y(\i_MIPS/Register/n424 ) );
  CLKMX2X2 U11834 ( .A(n5443), .B(\i_MIPS/Register/register[22][9] ), .S0(
        \i_MIPS/Register/n123 ), .Y(\i_MIPS/Register/n413 ) );
  CLKMX2X2 U11835 ( .A(n5463), .B(\i_MIPS/Register/register[23][30] ), .S0(
        \i_MIPS/Register/n121 ), .Y(\i_MIPS/Register/n402 ) );
  CLKMX2X2 U11836 ( .A(n5441), .B(\i_MIPS/Register/register[23][29] ), .S0(
        n5574), .Y(\i_MIPS/Register/n401 ) );
  CLKMX2X2 U11837 ( .A(n5461), .B(\i_MIPS/Register/register[23][24] ), .S0(
        n5575), .Y(\i_MIPS/Register/n396 ) );
  CLKMX2X2 U11838 ( .A(n5438), .B(\i_MIPS/Register/register[23][21] ), .S0(
        n5574), .Y(\i_MIPS/Register/n393 ) );
  CLKMX2X2 U11839 ( .A(n5435), .B(\i_MIPS/Register/register[23][20] ), .S0(
        n5575), .Y(\i_MIPS/Register/n392 ) );
  CLKMX2X2 U11840 ( .A(n5443), .B(\i_MIPS/Register/register[23][9] ), .S0(
        \i_MIPS/Register/n121 ), .Y(\i_MIPS/Register/n381 ) );
  CLKMX2X2 U11841 ( .A(n5463), .B(\i_MIPS/Register/register[24][30] ), .S0(
        n5572), .Y(\i_MIPS/Register/n370 ) );
  CLKMX2X2 U11842 ( .A(n5441), .B(\i_MIPS/Register/register[24][29] ), .S0(
        n5573), .Y(\i_MIPS/Register/n369 ) );
  CLKMX2X2 U11843 ( .A(n5461), .B(\i_MIPS/Register/register[24][24] ), .S0(
        n5572), .Y(\i_MIPS/Register/n364 ) );
  CLKMX2X2 U11844 ( .A(n5438), .B(\i_MIPS/Register/register[24][21] ), .S0(
        n5573), .Y(\i_MIPS/Register/n361 ) );
  CLKMX2X2 U11845 ( .A(n5435), .B(\i_MIPS/Register/register[24][20] ), .S0(
        \i_MIPS/Register/n118 ), .Y(\i_MIPS/Register/n360 ) );
  CLKMX2X2 U11846 ( .A(n5443), .B(\i_MIPS/Register/register[24][9] ), .S0(
        \i_MIPS/Register/n118 ), .Y(\i_MIPS/Register/n349 ) );
  CLKMX2X2 U11847 ( .A(n5463), .B(\i_MIPS/Register/register[25][30] ), .S0(
        n5570), .Y(\i_MIPS/Register/n338 ) );
  CLKMX2X2 U11848 ( .A(n5441), .B(\i_MIPS/Register/register[25][29] ), .S0(
        n5571), .Y(\i_MIPS/Register/n337 ) );
  CLKMX2X2 U11849 ( .A(n5461), .B(\i_MIPS/Register/register[25][24] ), .S0(
        n5570), .Y(\i_MIPS/Register/n332 ) );
  CLKMX2X2 U11850 ( .A(n5438), .B(\i_MIPS/Register/register[25][21] ), .S0(
        n5571), .Y(\i_MIPS/Register/n329 ) );
  CLKMX2X2 U11851 ( .A(n5435), .B(\i_MIPS/Register/register[25][20] ), .S0(
        \i_MIPS/Register/n116 ), .Y(\i_MIPS/Register/n328 ) );
  CLKMX2X2 U11852 ( .A(n5443), .B(\i_MIPS/Register/register[25][9] ), .S0(
        \i_MIPS/Register/n116 ), .Y(\i_MIPS/Register/n317 ) );
  CLKMX2X2 U11853 ( .A(n5463), .B(\i_MIPS/Register/register[26][30] ), .S0(
        n5568), .Y(\i_MIPS/Register/n306 ) );
  CLKMX2X2 U11854 ( .A(n5441), .B(\i_MIPS/Register/register[26][29] ), .S0(
        n5569), .Y(\i_MIPS/Register/n305 ) );
  CLKMX2X2 U11855 ( .A(n5461), .B(\i_MIPS/Register/register[26][24] ), .S0(
        n5568), .Y(\i_MIPS/Register/n300 ) );
  CLKMX2X2 U11856 ( .A(n5438), .B(\i_MIPS/Register/register[26][21] ), .S0(
        n5569), .Y(\i_MIPS/Register/n297 ) );
  CLKMX2X2 U11857 ( .A(n5435), .B(\i_MIPS/Register/register[26][20] ), .S0(
        \i_MIPS/Register/n114 ), .Y(\i_MIPS/Register/n296 ) );
  CLKMX2X2 U11858 ( .A(n5443), .B(\i_MIPS/Register/register[26][9] ), .S0(
        \i_MIPS/Register/n114 ), .Y(\i_MIPS/Register/n285 ) );
  CLKMX2X2 U11859 ( .A(n5462), .B(\i_MIPS/Register/register[27][30] ), .S0(
        \i_MIPS/Register/n112 ), .Y(\i_MIPS/Register/n274 ) );
  CLKMX2X2 U11860 ( .A(n5440), .B(\i_MIPS/Register/register[27][29] ), .S0(
        n5566), .Y(\i_MIPS/Register/n273 ) );
  CLKMX2X2 U11861 ( .A(n5460), .B(\i_MIPS/Register/register[27][24] ), .S0(
        n5567), .Y(\i_MIPS/Register/n268 ) );
  CLKMX2X2 U11862 ( .A(n5437), .B(\i_MIPS/Register/register[27][21] ), .S0(
        n5566), .Y(\i_MIPS/Register/n265 ) );
  CLKMX2X2 U11863 ( .A(n5434), .B(\i_MIPS/Register/register[27][20] ), .S0(
        n5567), .Y(\i_MIPS/Register/n264 ) );
  CLKMX2X2 U11864 ( .A(n5442), .B(\i_MIPS/Register/register[27][9] ), .S0(
        \i_MIPS/Register/n112 ), .Y(\i_MIPS/Register/n253 ) );
  CLKMX2X2 U11865 ( .A(n5463), .B(\i_MIPS/Register/register[28][30] ), .S0(
        n5564), .Y(\i_MIPS/Register/n242 ) );
  CLKMX2X2 U11866 ( .A(n5441), .B(\i_MIPS/Register/register[28][29] ), .S0(
        n5565), .Y(\i_MIPS/Register/n241 ) );
  CLKMX2X2 U11867 ( .A(n5461), .B(\i_MIPS/Register/register[28][24] ), .S0(
        n5564), .Y(\i_MIPS/Register/n236 ) );
  CLKMX2X2 U11868 ( .A(n5438), .B(\i_MIPS/Register/register[28][21] ), .S0(
        n5565), .Y(\i_MIPS/Register/n233 ) );
  CLKMX2X2 U11869 ( .A(n5435), .B(\i_MIPS/Register/register[28][20] ), .S0(
        \i_MIPS/Register/n110 ), .Y(\i_MIPS/Register/n232 ) );
  CLKMX2X2 U11870 ( .A(n5443), .B(\i_MIPS/Register/register[28][9] ), .S0(
        \i_MIPS/Register/n110 ), .Y(\i_MIPS/Register/n221 ) );
  CLKMX2X2 U11871 ( .A(n5463), .B(\i_MIPS/Register/register[29][30] ), .S0(
        \i_MIPS/Register/n108 ), .Y(\i_MIPS/Register/n210 ) );
  CLKMX2X2 U11872 ( .A(n5441), .B(\i_MIPS/Register/register[29][29] ), .S0(
        n5562), .Y(\i_MIPS/Register/n209 ) );
  CLKMX2X2 U11873 ( .A(n5461), .B(\i_MIPS/Register/register[29][24] ), .S0(
        n5563), .Y(\i_MIPS/Register/n204 ) );
  CLKMX2X2 U11874 ( .A(n5438), .B(\i_MIPS/Register/register[29][21] ), .S0(
        n5562), .Y(\i_MIPS/Register/n201 ) );
  CLKMX2X2 U11875 ( .A(n5435), .B(\i_MIPS/Register/register[29][20] ), .S0(
        n5563), .Y(\i_MIPS/Register/n200 ) );
  CLKMX2X2 U11876 ( .A(n5443), .B(\i_MIPS/Register/register[29][9] ), .S0(
        \i_MIPS/Register/n108 ), .Y(\i_MIPS/Register/n189 ) );
  CLKMX2X2 U11877 ( .A(n5463), .B(\i_MIPS/Register/register[30][30] ), .S0(
        n5560), .Y(\i_MIPS/Register/n178 ) );
  CLKMX2X2 U11878 ( .A(n5441), .B(\i_MIPS/Register/register[30][29] ), .S0(
        n5561), .Y(\i_MIPS/Register/n177 ) );
  CLKMX2X2 U11879 ( .A(n5461), .B(\i_MIPS/Register/register[30][24] ), .S0(
        n5560), .Y(\i_MIPS/Register/n172 ) );
  CLKMX2X2 U11880 ( .A(n5438), .B(\i_MIPS/Register/register[30][21] ), .S0(
        n5561), .Y(\i_MIPS/Register/n169 ) );
  CLKMX2X2 U11881 ( .A(n5435), .B(\i_MIPS/Register/register[30][20] ), .S0(
        \i_MIPS/Register/n106 ), .Y(\i_MIPS/Register/n168 ) );
  CLKMX2X2 U11882 ( .A(n5443), .B(\i_MIPS/Register/register[30][9] ), .S0(
        \i_MIPS/Register/n106 ), .Y(\i_MIPS/Register/n157 ) );
  CLKMX2X2 U11883 ( .A(n5402), .B(\i_MIPS/Register/register[0][16] ), .S0(
        n5620), .Y(\i_MIPS/Register/n1124 ) );
  CLKMX2X2 U11884 ( .A(n5402), .B(\i_MIPS/Register/register[1][16] ), .S0(
        n5618), .Y(\i_MIPS/Register/n1092 ) );
  CLKMX2X2 U11885 ( .A(n5402), .B(\i_MIPS/Register/register[2][16] ), .S0(
        n5616), .Y(\i_MIPS/Register/n1060 ) );
  CLKMX2X2 U11886 ( .A(n5402), .B(\i_MIPS/Register/register[3][16] ), .S0(
        n5614), .Y(\i_MIPS/Register/n1028 ) );
  CLKMX2X2 U11887 ( .A(n5402), .B(\i_MIPS/Register/register[4][16] ), .S0(
        n5612), .Y(\i_MIPS/Register/n996 ) );
  CLKMX2X2 U11888 ( .A(n5402), .B(\i_MIPS/Register/register[5][16] ), .S0(
        n5610), .Y(\i_MIPS/Register/n964 ) );
  CLKMX2X2 U11889 ( .A(n5402), .B(\i_MIPS/Register/register[6][16] ), .S0(
        n5608), .Y(\i_MIPS/Register/n932 ) );
  CLKMX2X2 U11890 ( .A(n5403), .B(\i_MIPS/Register/register[7][16] ), .S0(
        n5606), .Y(\i_MIPS/Register/n900 ) );
  CLKMX2X2 U11891 ( .A(n5402), .B(\i_MIPS/Register/register[8][16] ), .S0(
        n5604), .Y(\i_MIPS/Register/n868 ) );
  CLKMX2X2 U11892 ( .A(n5402), .B(\i_MIPS/Register/register[9][16] ), .S0(
        n5602), .Y(\i_MIPS/Register/n836 ) );
  CLKMX2X2 U11893 ( .A(n5402), .B(\i_MIPS/Register/register[10][16] ), .S0(
        n5600), .Y(\i_MIPS/Register/n804 ) );
  CLKMX2X2 U11894 ( .A(n5403), .B(\i_MIPS/Register/register[11][16] ), .S0(
        n5598), .Y(\i_MIPS/Register/n772 ) );
  CLKMX2X2 U11895 ( .A(n5402), .B(\i_MIPS/Register/register[12][16] ), .S0(
        n5596), .Y(\i_MIPS/Register/n740 ) );
  CLKMX2X2 U11896 ( .A(n5402), .B(\i_MIPS/Register/register[13][16] ), .S0(
        n5594), .Y(\i_MIPS/Register/n708 ) );
  CLKMX2X2 U11897 ( .A(n5402), .B(\i_MIPS/Register/register[14][16] ), .S0(
        n5592), .Y(\i_MIPS/Register/n676 ) );
  CLKMX2X2 U11898 ( .A(n5403), .B(\i_MIPS/Register/register[15][16] ), .S0(
        n5590), .Y(\i_MIPS/Register/n644 ) );
  CLKMX2X2 U11899 ( .A(n5403), .B(\i_MIPS/Register/register[16][16] ), .S0(
        n5588), .Y(\i_MIPS/Register/n612 ) );
  CLKMX2X2 U11900 ( .A(n5403), .B(\i_MIPS/Register/register[17][16] ), .S0(
        n5586), .Y(\i_MIPS/Register/n580 ) );
  CLKMX2X2 U11901 ( .A(n5403), .B(\i_MIPS/Register/register[18][16] ), .S0(
        n5584), .Y(\i_MIPS/Register/n548 ) );
  CLKMX2X2 U11902 ( .A(n5402), .B(\i_MIPS/Register/register[19][16] ), .S0(
        n5582), .Y(\i_MIPS/Register/n516 ) );
  CLKMX2X2 U11903 ( .A(n5403), .B(\i_MIPS/Register/register[20][16] ), .S0(
        n5580), .Y(\i_MIPS/Register/n484 ) );
  CLKMX2X2 U11904 ( .A(n5403), .B(\i_MIPS/Register/register[21][16] ), .S0(
        n5578), .Y(\i_MIPS/Register/n452 ) );
  CLKMX2X2 U11905 ( .A(n5403), .B(\i_MIPS/Register/register[22][16] ), .S0(
        n5576), .Y(\i_MIPS/Register/n420 ) );
  CLKMX2X2 U11906 ( .A(n5402), .B(\i_MIPS/Register/register[23][16] ), .S0(
        n5574), .Y(\i_MIPS/Register/n388 ) );
  CLKMX2X2 U11907 ( .A(n5403), .B(\i_MIPS/Register/register[24][16] ), .S0(
        n5572), .Y(\i_MIPS/Register/n356 ) );
  CLKMX2X2 U11908 ( .A(n5403), .B(\i_MIPS/Register/register[25][16] ), .S0(
        n5570), .Y(\i_MIPS/Register/n324 ) );
  CLKMX2X2 U11909 ( .A(n5403), .B(\i_MIPS/Register/register[26][16] ), .S0(
        n5568), .Y(\i_MIPS/Register/n292 ) );
  CLKMX2X2 U11910 ( .A(n5403), .B(\i_MIPS/Register/register[27][16] ), .S0(
        n5566), .Y(\i_MIPS/Register/n260 ) );
  CLKMX2X2 U11911 ( .A(n5403), .B(\i_MIPS/Register/register[28][16] ), .S0(
        n5564), .Y(\i_MIPS/Register/n228 ) );
  CLKMX2X2 U11912 ( .A(n5402), .B(\i_MIPS/Register/register[29][16] ), .S0(
        n5562), .Y(\i_MIPS/Register/n196 ) );
  CLKMX2X2 U11913 ( .A(n5403), .B(\i_MIPS/Register/register[30][16] ), .S0(
        n5560), .Y(\i_MIPS/Register/n164 ) );
  CLKMX2X2 U11914 ( .A(n5469), .B(\i_MIPS/Register/register[0][31] ), .S0(
        n5621), .Y(\i_MIPS/Register/n1139 ) );
  CLKMX2X2 U11915 ( .A(n5462), .B(\i_MIPS/Register/register[0][30] ), .S0(
        n5621), .Y(\i_MIPS/Register/n1138 ) );
  CLKMX2X2 U11916 ( .A(n5440), .B(\i_MIPS/Register/register[0][29] ), .S0(
        n5621), .Y(\i_MIPS/Register/n1137 ) );
  CLKMX2X2 U11917 ( .A(n5410), .B(\i_MIPS/Register/register[0][28] ), .S0(
        n5620), .Y(\i_MIPS/Register/n1136 ) );
  CLKMX2X2 U11918 ( .A(n5407), .B(\i_MIPS/Register/register[0][27] ), .S0(
        n5620), .Y(\i_MIPS/Register/n1135 ) );
  CLKMX2X2 U11919 ( .A(n5404), .B(\i_MIPS/Register/register[0][26] ), .S0(
        n5620), .Y(\i_MIPS/Register/n1134 ) );
  CLKMX2X2 U11920 ( .A(n5413), .B(\i_MIPS/Register/register[0][25] ), .S0(
        n5620), .Y(\i_MIPS/Register/n1133 ) );
  CLKMX2X2 U11921 ( .A(n5460), .B(\i_MIPS/Register/register[0][24] ), .S0(
        n5621), .Y(\i_MIPS/Register/n1132 ) );
  CLKMX2X2 U11922 ( .A(n5422), .B(\i_MIPS/Register/register[0][22] ), .S0(
        n5620), .Y(\i_MIPS/Register/n1130 ) );
  CLKMX2X2 U11923 ( .A(n5437), .B(\i_MIPS/Register/register[0][21] ), .S0(
        n5620), .Y(\i_MIPS/Register/n1129 ) );
  CLKMX2X2 U11924 ( .A(n5434), .B(\i_MIPS/Register/register[0][20] ), .S0(
        n5620), .Y(\i_MIPS/Register/n1128 ) );
  CLKMX2X2 U11925 ( .A(n5431), .B(\i_MIPS/Register/register[0][19] ), .S0(
        n5620), .Y(\i_MIPS/Register/n1127 ) );
  CLKMX2X2 U11926 ( .A(n5416), .B(\i_MIPS/Register/register[0][18] ), .S0(
        n5620), .Y(\i_MIPS/Register/n1126 ) );
  CLKMX2X2 U11927 ( .A(n5457), .B(\i_MIPS/Register/register[0][17] ), .S0(
        n5621), .Y(\i_MIPS/Register/n1125 ) );
  CLKMX2X2 U11928 ( .A(n5455), .B(\i_MIPS/Register/register[0][15] ), .S0(
        n5621), .Y(\i_MIPS/Register/n1123 ) );
  CLKMX2X2 U11929 ( .A(n5453), .B(\i_MIPS/Register/register[0][14] ), .S0(
        n5621), .Y(\i_MIPS/Register/n1122 ) );
  CLKMX2X2 U11930 ( .A(n5451), .B(\i_MIPS/Register/register[0][13] ), .S0(
        n5621), .Y(\i_MIPS/Register/n1121 ) );
  CLKMX2X2 U11931 ( .A(n5449), .B(\i_MIPS/Register/register[0][12] ), .S0(
        n5621), .Y(\i_MIPS/Register/n1120 ) );
  CLKMX2X2 U11932 ( .A(n5445), .B(\i_MIPS/Register/register[0][11] ), .S0(
        n5621), .Y(\i_MIPS/Register/n1119 ) );
  CLKMX2X2 U11933 ( .A(n5419), .B(\i_MIPS/Register/register[0][10] ), .S0(
        n5620), .Y(\i_MIPS/Register/n1118 ) );
  CLKMX2X2 U11934 ( .A(n5443), .B(\i_MIPS/Register/register[0][9] ), .S0(n5621), .Y(\i_MIPS/Register/n1117 ) );
  CLKMX2X2 U11935 ( .A(n5474), .B(\i_MIPS/Register/register[0][8] ), .S0(n5621), .Y(\i_MIPS/Register/n1116 ) );
  CLKMX2X2 U11936 ( .A(n5471), .B(\i_MIPS/Register/register[0][7] ), .S0(n5621), .Y(\i_MIPS/Register/n1115 ) );
  CLKMX2X2 U11937 ( .A(n5042), .B(\i_MIPS/Register/register[0][6] ), .S0(n5620), .Y(\i_MIPS/Register/n1114 ) );
  CLKMX2X2 U11938 ( .A(n4775), .B(\i_MIPS/Register/register[0][3] ), .S0(n5620), .Y(\i_MIPS/Register/n1111 ) );
  CLKMX2X2 U11939 ( .A(n5469), .B(\i_MIPS/Register/register[1][31] ), .S0(
        n5618), .Y(\i_MIPS/Register/n1107 ) );
  CLKMX2X2 U11940 ( .A(n5410), .B(\i_MIPS/Register/register[1][28] ), .S0(
        n5619), .Y(\i_MIPS/Register/n1104 ) );
  CLKMX2X2 U11941 ( .A(n5407), .B(\i_MIPS/Register/register[1][27] ), .S0(
        n5618), .Y(\i_MIPS/Register/n1103 ) );
  CLKMX2X2 U11942 ( .A(n5404), .B(\i_MIPS/Register/register[1][26] ), .S0(
        n5618), .Y(\i_MIPS/Register/n1102 ) );
  CLKMX2X2 U11943 ( .A(n5413), .B(\i_MIPS/Register/register[1][25] ), .S0(
        n5619), .Y(\i_MIPS/Register/n1101 ) );
  CLKMX2X2 U11944 ( .A(n5482), .B(\i_MIPS/Register/register[1][23] ), .S0(
        n5619), .Y(\i_MIPS/Register/n1099 ) );
  CLKMX2X2 U11945 ( .A(n5422), .B(\i_MIPS/Register/register[1][22] ), .S0(
        n5618), .Y(\i_MIPS/Register/n1098 ) );
  CLKMX2X2 U11946 ( .A(n5431), .B(\i_MIPS/Register/register[1][19] ), .S0(
        n5618), .Y(\i_MIPS/Register/n1095 ) );
  CLKMX2X2 U11947 ( .A(n5416), .B(\i_MIPS/Register/register[1][18] ), .S0(
        n5619), .Y(\i_MIPS/Register/n1094 ) );
  CLKMX2X2 U11948 ( .A(n5457), .B(\i_MIPS/Register/register[1][17] ), .S0(
        n5619), .Y(\i_MIPS/Register/n1093 ) );
  CLKMX2X2 U11949 ( .A(n5455), .B(\i_MIPS/Register/register[1][15] ), .S0(
        n5619), .Y(\i_MIPS/Register/n1091 ) );
  CLKMX2X2 U11950 ( .A(n5453), .B(\i_MIPS/Register/register[1][14] ), .S0(
        n5619), .Y(\i_MIPS/Register/n1090 ) );
  CLKMX2X2 U11951 ( .A(n5451), .B(\i_MIPS/Register/register[1][13] ), .S0(
        n5619), .Y(\i_MIPS/Register/n1089 ) );
  CLKMX2X2 U11952 ( .A(n5448), .B(\i_MIPS/Register/register[1][12] ), .S0(
        n5619), .Y(\i_MIPS/Register/n1088 ) );
  CLKMX2X2 U11953 ( .A(n5445), .B(\i_MIPS/Register/register[1][11] ), .S0(
        n5618), .Y(\i_MIPS/Register/n1087 ) );
  CLKMX2X2 U11954 ( .A(n5419), .B(\i_MIPS/Register/register[1][10] ), .S0(
        n5618), .Y(\i_MIPS/Register/n1086 ) );
  CLKMX2X2 U11955 ( .A(n5474), .B(\i_MIPS/Register/register[1][8] ), .S0(n5619), .Y(\i_MIPS/Register/n1084 ) );
  CLKMX2X2 U11956 ( .A(n5471), .B(\i_MIPS/Register/register[1][7] ), .S0(n5619), .Y(\i_MIPS/Register/n1083 ) );
  CLKMX2X2 U11957 ( .A(n5042), .B(\i_MIPS/Register/register[1][6] ), .S0(n5618), .Y(\i_MIPS/Register/n1082 ) );
  CLKMX2X2 U11958 ( .A(n5490), .B(\i_MIPS/Register/register[1][5] ), .S0(n5618), .Y(\i_MIPS/Register/n1081 ) );
  CLKMX2X2 U11959 ( .A(n5487), .B(\i_MIPS/Register/register[1][4] ), .S0(n5618), .Y(\i_MIPS/Register/n1080 ) );
  CLKMX2X2 U11960 ( .A(n4775), .B(\i_MIPS/Register/register[1][3] ), .S0(n5618), .Y(\i_MIPS/Register/n1079 ) );
  CLKMX2X2 U11961 ( .A(n5479), .B(\i_MIPS/Register/register[1][2] ), .S0(n5618), .Y(\i_MIPS/Register/n1078 ) );
  CLKMX2X2 U11962 ( .A(n5476), .B(\i_MIPS/Register/register[1][1] ), .S0(n5619), .Y(\i_MIPS/Register/n1077 ) );
  CLKMX2X2 U11963 ( .A(n5484), .B(\i_MIPS/Register/register[1][0] ), .S0(n5619), .Y(\i_MIPS/Register/n1076 ) );
  CLKMX2X2 U11964 ( .A(n5469), .B(\i_MIPS/Register/register[2][31] ), .S0(
        n5616), .Y(\i_MIPS/Register/n1075 ) );
  CLKMX2X2 U11965 ( .A(n5410), .B(\i_MIPS/Register/register[2][28] ), .S0(
        n5617), .Y(\i_MIPS/Register/n1072 ) );
  CLKMX2X2 U11966 ( .A(n5407), .B(\i_MIPS/Register/register[2][27] ), .S0(
        n5616), .Y(\i_MIPS/Register/n1071 ) );
  CLKMX2X2 U11967 ( .A(n5404), .B(\i_MIPS/Register/register[2][26] ), .S0(
        n5616), .Y(\i_MIPS/Register/n1070 ) );
  CLKMX2X2 U11968 ( .A(n5413), .B(\i_MIPS/Register/register[2][25] ), .S0(
        n5617), .Y(\i_MIPS/Register/n1069 ) );
  CLKMX2X2 U11969 ( .A(n5482), .B(\i_MIPS/Register/register[2][23] ), .S0(
        n5617), .Y(\i_MIPS/Register/n1067 ) );
  CLKMX2X2 U11970 ( .A(n5422), .B(\i_MIPS/Register/register[2][22] ), .S0(
        n5616), .Y(\i_MIPS/Register/n1066 ) );
  CLKMX2X2 U11971 ( .A(n5431), .B(\i_MIPS/Register/register[2][19] ), .S0(
        n5616), .Y(\i_MIPS/Register/n1063 ) );
  CLKMX2X2 U11972 ( .A(n5416), .B(\i_MIPS/Register/register[2][18] ), .S0(
        n5617), .Y(\i_MIPS/Register/n1062 ) );
  CLKMX2X2 U11973 ( .A(n5457), .B(\i_MIPS/Register/register[2][17] ), .S0(
        n5617), .Y(\i_MIPS/Register/n1061 ) );
  CLKMX2X2 U11974 ( .A(n5455), .B(\i_MIPS/Register/register[2][15] ), .S0(
        n5617), .Y(\i_MIPS/Register/n1059 ) );
  CLKMX2X2 U11975 ( .A(n5453), .B(\i_MIPS/Register/register[2][14] ), .S0(
        n5617), .Y(\i_MIPS/Register/n1058 ) );
  CLKMX2X2 U11976 ( .A(n5451), .B(\i_MIPS/Register/register[2][13] ), .S0(
        n5617), .Y(\i_MIPS/Register/n1057 ) );
  CLKMX2X2 U11977 ( .A(n5448), .B(\i_MIPS/Register/register[2][12] ), .S0(
        n5617), .Y(\i_MIPS/Register/n1056 ) );
  CLKMX2X2 U11978 ( .A(n5445), .B(\i_MIPS/Register/register[2][11] ), .S0(
        n5616), .Y(\i_MIPS/Register/n1055 ) );
  CLKMX2X2 U11979 ( .A(n5419), .B(\i_MIPS/Register/register[2][10] ), .S0(
        n5616), .Y(\i_MIPS/Register/n1054 ) );
  CLKMX2X2 U11980 ( .A(n5474), .B(\i_MIPS/Register/register[2][8] ), .S0(n5617), .Y(\i_MIPS/Register/n1052 ) );
  CLKMX2X2 U11981 ( .A(n5471), .B(\i_MIPS/Register/register[2][7] ), .S0(n5617), .Y(\i_MIPS/Register/n1051 ) );
  CLKMX2X2 U11982 ( .A(n5042), .B(\i_MIPS/Register/register[2][6] ), .S0(n5616), .Y(\i_MIPS/Register/n1050 ) );
  CLKMX2X2 U11983 ( .A(n5490), .B(\i_MIPS/Register/register[2][5] ), .S0(n5616), .Y(\i_MIPS/Register/n1049 ) );
  CLKMX2X2 U11984 ( .A(n5487), .B(\i_MIPS/Register/register[2][4] ), .S0(n5616), .Y(\i_MIPS/Register/n1048 ) );
  CLKMX2X2 U11985 ( .A(n4775), .B(\i_MIPS/Register/register[2][3] ), .S0(n5616), .Y(\i_MIPS/Register/n1047 ) );
  CLKMX2X2 U11986 ( .A(n5479), .B(\i_MIPS/Register/register[2][2] ), .S0(n5616), .Y(\i_MIPS/Register/n1046 ) );
  CLKMX2X2 U11987 ( .A(n5476), .B(\i_MIPS/Register/register[2][1] ), .S0(n5617), .Y(\i_MIPS/Register/n1045 ) );
  CLKMX2X2 U11988 ( .A(n5484), .B(\i_MIPS/Register/register[2][0] ), .S0(n5617), .Y(\i_MIPS/Register/n1044 ) );
  CLKMX2X2 U11989 ( .A(n5469), .B(\i_MIPS/Register/register[3][31] ), .S0(
        n5614), .Y(\i_MIPS/Register/n1043 ) );
  CLKMX2X2 U11990 ( .A(n5410), .B(\i_MIPS/Register/register[3][28] ), .S0(
        n5615), .Y(\i_MIPS/Register/n1040 ) );
  CLKMX2X2 U11991 ( .A(n5407), .B(\i_MIPS/Register/register[3][27] ), .S0(
        n5614), .Y(\i_MIPS/Register/n1039 ) );
  CLKMX2X2 U11992 ( .A(n5404), .B(\i_MIPS/Register/register[3][26] ), .S0(
        n5614), .Y(\i_MIPS/Register/n1038 ) );
  CLKMX2X2 U11993 ( .A(n5413), .B(\i_MIPS/Register/register[3][25] ), .S0(
        n5615), .Y(\i_MIPS/Register/n1037 ) );
  CLKMX2X2 U11994 ( .A(n5482), .B(\i_MIPS/Register/register[3][23] ), .S0(
        n5615), .Y(\i_MIPS/Register/n1035 ) );
  CLKMX2X2 U11995 ( .A(n5422), .B(\i_MIPS/Register/register[3][22] ), .S0(
        n5614), .Y(\i_MIPS/Register/n1034 ) );
  CLKMX2X2 U11996 ( .A(n5431), .B(\i_MIPS/Register/register[3][19] ), .S0(
        n5614), .Y(\i_MIPS/Register/n1031 ) );
  CLKMX2X2 U11997 ( .A(n5416), .B(\i_MIPS/Register/register[3][18] ), .S0(
        n5615), .Y(\i_MIPS/Register/n1030 ) );
  CLKMX2X2 U11998 ( .A(n5457), .B(\i_MIPS/Register/register[3][17] ), .S0(
        n5615), .Y(\i_MIPS/Register/n1029 ) );
  CLKMX2X2 U11999 ( .A(n5455), .B(\i_MIPS/Register/register[3][15] ), .S0(
        n5615), .Y(\i_MIPS/Register/n1027 ) );
  CLKMX2X2 U12000 ( .A(n5453), .B(\i_MIPS/Register/register[3][14] ), .S0(
        n5615), .Y(\i_MIPS/Register/n1026 ) );
  CLKMX2X2 U12001 ( .A(n5451), .B(\i_MIPS/Register/register[3][13] ), .S0(
        n5615), .Y(\i_MIPS/Register/n1025 ) );
  CLKMX2X2 U12002 ( .A(n5448), .B(\i_MIPS/Register/register[3][12] ), .S0(
        n5615), .Y(\i_MIPS/Register/n1024 ) );
  CLKMX2X2 U12003 ( .A(n5445), .B(\i_MIPS/Register/register[3][11] ), .S0(
        n5614), .Y(\i_MIPS/Register/n1023 ) );
  CLKMX2X2 U12004 ( .A(n5419), .B(\i_MIPS/Register/register[3][10] ), .S0(
        n5614), .Y(\i_MIPS/Register/n1022 ) );
  CLKMX2X2 U12005 ( .A(n5474), .B(\i_MIPS/Register/register[3][8] ), .S0(n5615), .Y(\i_MIPS/Register/n1020 ) );
  CLKMX2X2 U12006 ( .A(n5471), .B(\i_MIPS/Register/register[3][7] ), .S0(n5615), .Y(\i_MIPS/Register/n1019 ) );
  CLKMX2X2 U12007 ( .A(n5042), .B(\i_MIPS/Register/register[3][6] ), .S0(n5614), .Y(\i_MIPS/Register/n1018 ) );
  CLKMX2X2 U12008 ( .A(n5490), .B(\i_MIPS/Register/register[3][5] ), .S0(n5614), .Y(\i_MIPS/Register/n1017 ) );
  CLKMX2X2 U12009 ( .A(n5487), .B(\i_MIPS/Register/register[3][4] ), .S0(n5614), .Y(\i_MIPS/Register/n1016 ) );
  CLKMX2X2 U12010 ( .A(n4775), .B(\i_MIPS/Register/register[3][3] ), .S0(n5614), .Y(\i_MIPS/Register/n1015 ) );
  CLKMX2X2 U12011 ( .A(n5479), .B(\i_MIPS/Register/register[3][2] ), .S0(n5614), .Y(\i_MIPS/Register/n1014 ) );
  CLKMX2X2 U12012 ( .A(n5476), .B(\i_MIPS/Register/register[3][1] ), .S0(n5615), .Y(\i_MIPS/Register/n1013 ) );
  CLKMX2X2 U12013 ( .A(n5484), .B(\i_MIPS/Register/register[3][0] ), .S0(n5615), .Y(\i_MIPS/Register/n1012 ) );
  CLKMX2X2 U12014 ( .A(n5469), .B(\i_MIPS/Register/register[4][31] ), .S0(
        n5612), .Y(\i_MIPS/Register/n1011 ) );
  CLKMX2X2 U12015 ( .A(n5410), .B(\i_MIPS/Register/register[4][28] ), .S0(
        n5613), .Y(\i_MIPS/Register/n1008 ) );
  CLKMX2X2 U12016 ( .A(n5407), .B(\i_MIPS/Register/register[4][27] ), .S0(
        n5612), .Y(\i_MIPS/Register/n1007 ) );
  CLKMX2X2 U12017 ( .A(n5404), .B(\i_MIPS/Register/register[4][26] ), .S0(
        n5612), .Y(\i_MIPS/Register/n1006 ) );
  CLKMX2X2 U12018 ( .A(n5413), .B(\i_MIPS/Register/register[4][25] ), .S0(
        n5613), .Y(\i_MIPS/Register/n1005 ) );
  CLKMX2X2 U12019 ( .A(n5482), .B(\i_MIPS/Register/register[4][23] ), .S0(
        n5613), .Y(\i_MIPS/Register/n1003 ) );
  CLKMX2X2 U12020 ( .A(n5422), .B(\i_MIPS/Register/register[4][22] ), .S0(
        n5612), .Y(\i_MIPS/Register/n1002 ) );
  CLKMX2X2 U12021 ( .A(n5431), .B(\i_MIPS/Register/register[4][19] ), .S0(
        n5612), .Y(\i_MIPS/Register/n999 ) );
  CLKMX2X2 U12022 ( .A(n5416), .B(\i_MIPS/Register/register[4][18] ), .S0(
        n5613), .Y(\i_MIPS/Register/n998 ) );
  CLKMX2X2 U12023 ( .A(n5457), .B(\i_MIPS/Register/register[4][17] ), .S0(
        n5613), .Y(\i_MIPS/Register/n997 ) );
  CLKMX2X2 U12024 ( .A(n5455), .B(\i_MIPS/Register/register[4][15] ), .S0(
        n5613), .Y(\i_MIPS/Register/n995 ) );
  CLKMX2X2 U12025 ( .A(n5453), .B(\i_MIPS/Register/register[4][14] ), .S0(
        n5613), .Y(\i_MIPS/Register/n994 ) );
  CLKMX2X2 U12026 ( .A(n5451), .B(\i_MIPS/Register/register[4][13] ), .S0(
        n5613), .Y(\i_MIPS/Register/n993 ) );
  CLKMX2X2 U12027 ( .A(n5448), .B(\i_MIPS/Register/register[4][12] ), .S0(
        n5613), .Y(\i_MIPS/Register/n992 ) );
  CLKMX2X2 U12028 ( .A(n5445), .B(\i_MIPS/Register/register[4][11] ), .S0(
        n5612), .Y(\i_MIPS/Register/n991 ) );
  CLKMX2X2 U12029 ( .A(n5419), .B(\i_MIPS/Register/register[4][10] ), .S0(
        n5612), .Y(\i_MIPS/Register/n990 ) );
  CLKMX2X2 U12030 ( .A(n5474), .B(\i_MIPS/Register/register[4][8] ), .S0(n5613), .Y(\i_MIPS/Register/n988 ) );
  CLKMX2X2 U12031 ( .A(n5471), .B(\i_MIPS/Register/register[4][7] ), .S0(n5613), .Y(\i_MIPS/Register/n987 ) );
  CLKMX2X2 U12032 ( .A(n5042), .B(\i_MIPS/Register/register[4][6] ), .S0(n5612), .Y(\i_MIPS/Register/n986 ) );
  CLKMX2X2 U12033 ( .A(n5490), .B(\i_MIPS/Register/register[4][5] ), .S0(n5612), .Y(\i_MIPS/Register/n985 ) );
  CLKMX2X2 U12034 ( .A(n5487), .B(\i_MIPS/Register/register[4][4] ), .S0(n5612), .Y(\i_MIPS/Register/n984 ) );
  CLKMX2X2 U12035 ( .A(n4775), .B(\i_MIPS/Register/register[4][3] ), .S0(n5612), .Y(\i_MIPS/Register/n983 ) );
  CLKMX2X2 U12036 ( .A(n5479), .B(\i_MIPS/Register/register[4][2] ), .S0(n5612), .Y(\i_MIPS/Register/n982 ) );
  CLKMX2X2 U12037 ( .A(n5476), .B(\i_MIPS/Register/register[4][1] ), .S0(n5613), .Y(\i_MIPS/Register/n981 ) );
  CLKMX2X2 U12038 ( .A(n5484), .B(\i_MIPS/Register/register[4][0] ), .S0(n5613), .Y(\i_MIPS/Register/n980 ) );
  CLKMX2X2 U12039 ( .A(n5469), .B(\i_MIPS/Register/register[5][31] ), .S0(
        n5610), .Y(\i_MIPS/Register/n979 ) );
  CLKMX2X2 U12040 ( .A(n5410), .B(\i_MIPS/Register/register[5][28] ), .S0(
        n5611), .Y(\i_MIPS/Register/n976 ) );
  CLKMX2X2 U12041 ( .A(n5407), .B(\i_MIPS/Register/register[5][27] ), .S0(
        n5610), .Y(\i_MIPS/Register/n975 ) );
  CLKMX2X2 U12042 ( .A(n5404), .B(\i_MIPS/Register/register[5][26] ), .S0(
        n5610), .Y(\i_MIPS/Register/n974 ) );
  CLKMX2X2 U12043 ( .A(n5413), .B(\i_MIPS/Register/register[5][25] ), .S0(
        n5611), .Y(\i_MIPS/Register/n973 ) );
  CLKMX2X2 U12044 ( .A(n5482), .B(\i_MIPS/Register/register[5][23] ), .S0(
        n5611), .Y(\i_MIPS/Register/n971 ) );
  CLKMX2X2 U12045 ( .A(n5422), .B(\i_MIPS/Register/register[5][22] ), .S0(
        n5610), .Y(\i_MIPS/Register/n970 ) );
  CLKMX2X2 U12046 ( .A(n5431), .B(\i_MIPS/Register/register[5][19] ), .S0(
        n5610), .Y(\i_MIPS/Register/n967 ) );
  CLKMX2X2 U12047 ( .A(n5416), .B(\i_MIPS/Register/register[5][18] ), .S0(
        n5611), .Y(\i_MIPS/Register/n966 ) );
  CLKMX2X2 U12048 ( .A(n5457), .B(\i_MIPS/Register/register[5][17] ), .S0(
        n5611), .Y(\i_MIPS/Register/n965 ) );
  CLKMX2X2 U12049 ( .A(n5455), .B(\i_MIPS/Register/register[5][15] ), .S0(
        n5611), .Y(\i_MIPS/Register/n963 ) );
  CLKMX2X2 U12050 ( .A(n5453), .B(\i_MIPS/Register/register[5][14] ), .S0(
        n5611), .Y(\i_MIPS/Register/n962 ) );
  CLKMX2X2 U12051 ( .A(n5451), .B(\i_MIPS/Register/register[5][13] ), .S0(
        n5611), .Y(\i_MIPS/Register/n961 ) );
  CLKMX2X2 U12052 ( .A(n5448), .B(\i_MIPS/Register/register[5][12] ), .S0(
        n5611), .Y(\i_MIPS/Register/n960 ) );
  CLKMX2X2 U12053 ( .A(n5445), .B(\i_MIPS/Register/register[5][11] ), .S0(
        n5610), .Y(\i_MIPS/Register/n959 ) );
  CLKMX2X2 U12054 ( .A(n5419), .B(\i_MIPS/Register/register[5][10] ), .S0(
        n5610), .Y(\i_MIPS/Register/n958 ) );
  CLKMX2X2 U12055 ( .A(n5474), .B(\i_MIPS/Register/register[5][8] ), .S0(n5611), .Y(\i_MIPS/Register/n956 ) );
  CLKMX2X2 U12056 ( .A(n5471), .B(\i_MIPS/Register/register[5][7] ), .S0(n5611), .Y(\i_MIPS/Register/n955 ) );
  CLKMX2X2 U12057 ( .A(n5042), .B(\i_MIPS/Register/register[5][6] ), .S0(n5610), .Y(\i_MIPS/Register/n954 ) );
  CLKMX2X2 U12058 ( .A(n5490), .B(\i_MIPS/Register/register[5][5] ), .S0(n5610), .Y(\i_MIPS/Register/n953 ) );
  CLKMX2X2 U12059 ( .A(n5487), .B(\i_MIPS/Register/register[5][4] ), .S0(n5610), .Y(\i_MIPS/Register/n952 ) );
  CLKMX2X2 U12060 ( .A(n4775), .B(\i_MIPS/Register/register[5][3] ), .S0(n5610), .Y(\i_MIPS/Register/n951 ) );
  CLKMX2X2 U12061 ( .A(n5479), .B(\i_MIPS/Register/register[5][2] ), .S0(n5610), .Y(\i_MIPS/Register/n950 ) );
  CLKMX2X2 U12062 ( .A(n5476), .B(\i_MIPS/Register/register[5][1] ), .S0(n5611), .Y(\i_MIPS/Register/n949 ) );
  CLKMX2X2 U12063 ( .A(n5484), .B(\i_MIPS/Register/register[5][0] ), .S0(n5611), .Y(\i_MIPS/Register/n948 ) );
  CLKMX2X2 U12064 ( .A(n5469), .B(\i_MIPS/Register/register[6][31] ), .S0(
        n5608), .Y(\i_MIPS/Register/n947 ) );
  CLKMX2X2 U12065 ( .A(n5410), .B(\i_MIPS/Register/register[6][28] ), .S0(
        n5609), .Y(\i_MIPS/Register/n944 ) );
  CLKMX2X2 U12066 ( .A(n5407), .B(\i_MIPS/Register/register[6][27] ), .S0(
        n5608), .Y(\i_MIPS/Register/n943 ) );
  CLKMX2X2 U12067 ( .A(n5404), .B(\i_MIPS/Register/register[6][26] ), .S0(
        n5608), .Y(\i_MIPS/Register/n942 ) );
  CLKMX2X2 U12068 ( .A(n5413), .B(\i_MIPS/Register/register[6][25] ), .S0(
        n5609), .Y(\i_MIPS/Register/n941 ) );
  CLKMX2X2 U12069 ( .A(n5482), .B(\i_MIPS/Register/register[6][23] ), .S0(
        n5609), .Y(\i_MIPS/Register/n939 ) );
  CLKMX2X2 U12070 ( .A(n5422), .B(\i_MIPS/Register/register[6][22] ), .S0(
        n5608), .Y(\i_MIPS/Register/n938 ) );
  CLKMX2X2 U12071 ( .A(n5431), .B(\i_MIPS/Register/register[6][19] ), .S0(
        n5608), .Y(\i_MIPS/Register/n935 ) );
  CLKMX2X2 U12072 ( .A(n5416), .B(\i_MIPS/Register/register[6][18] ), .S0(
        n5609), .Y(\i_MIPS/Register/n934 ) );
  CLKMX2X2 U12073 ( .A(n5457), .B(\i_MIPS/Register/register[6][17] ), .S0(
        n5609), .Y(\i_MIPS/Register/n933 ) );
  CLKMX2X2 U12074 ( .A(n5455), .B(\i_MIPS/Register/register[6][15] ), .S0(
        n5609), .Y(\i_MIPS/Register/n931 ) );
  CLKMX2X2 U12075 ( .A(n5453), .B(\i_MIPS/Register/register[6][14] ), .S0(
        n5609), .Y(\i_MIPS/Register/n930 ) );
  CLKMX2X2 U12076 ( .A(n5451), .B(\i_MIPS/Register/register[6][13] ), .S0(
        n5609), .Y(\i_MIPS/Register/n929 ) );
  CLKMX2X2 U12077 ( .A(n5448), .B(\i_MIPS/Register/register[6][12] ), .S0(
        n5609), .Y(\i_MIPS/Register/n928 ) );
  CLKMX2X2 U12078 ( .A(n5445), .B(\i_MIPS/Register/register[6][11] ), .S0(
        n5608), .Y(\i_MIPS/Register/n927 ) );
  CLKMX2X2 U12079 ( .A(n5419), .B(\i_MIPS/Register/register[6][10] ), .S0(
        n5608), .Y(\i_MIPS/Register/n926 ) );
  CLKMX2X2 U12080 ( .A(n5474), .B(\i_MIPS/Register/register[6][8] ), .S0(n5609), .Y(\i_MIPS/Register/n924 ) );
  CLKMX2X2 U12081 ( .A(n5471), .B(\i_MIPS/Register/register[6][7] ), .S0(n5609), .Y(\i_MIPS/Register/n923 ) );
  CLKMX2X2 U12082 ( .A(n5042), .B(\i_MIPS/Register/register[6][6] ), .S0(n5608), .Y(\i_MIPS/Register/n922 ) );
  CLKMX2X2 U12083 ( .A(n5490), .B(\i_MIPS/Register/register[6][5] ), .S0(n5608), .Y(\i_MIPS/Register/n921 ) );
  CLKMX2X2 U12084 ( .A(n5487), .B(\i_MIPS/Register/register[6][4] ), .S0(n5608), .Y(\i_MIPS/Register/n920 ) );
  CLKMX2X2 U12085 ( .A(n4775), .B(\i_MIPS/Register/register[6][3] ), .S0(n5608), .Y(\i_MIPS/Register/n919 ) );
  CLKMX2X2 U12086 ( .A(n5479), .B(\i_MIPS/Register/register[6][2] ), .S0(n5608), .Y(\i_MIPS/Register/n918 ) );
  CLKMX2X2 U12087 ( .A(n5476), .B(\i_MIPS/Register/register[6][1] ), .S0(n5609), .Y(\i_MIPS/Register/n917 ) );
  CLKMX2X2 U12088 ( .A(n5484), .B(\i_MIPS/Register/register[6][0] ), .S0(n5609), .Y(\i_MIPS/Register/n916 ) );
  CLKMX2X2 U12089 ( .A(n5470), .B(\i_MIPS/Register/register[7][31] ), .S0(
        n5606), .Y(\i_MIPS/Register/n915 ) );
  CLKMX2X2 U12090 ( .A(n5411), .B(\i_MIPS/Register/register[7][28] ), .S0(
        n5607), .Y(\i_MIPS/Register/n912 ) );
  CLKMX2X2 U12091 ( .A(n5408), .B(\i_MIPS/Register/register[7][27] ), .S0(
        n5606), .Y(\i_MIPS/Register/n911 ) );
  CLKMX2X2 U12092 ( .A(n5405), .B(\i_MIPS/Register/register[7][26] ), .S0(
        n5606), .Y(\i_MIPS/Register/n910 ) );
  CLKMX2X2 U12093 ( .A(n5414), .B(\i_MIPS/Register/register[7][25] ), .S0(
        n5607), .Y(\i_MIPS/Register/n909 ) );
  CLKMX2X2 U12094 ( .A(n5483), .B(\i_MIPS/Register/register[7][23] ), .S0(
        n5607), .Y(\i_MIPS/Register/n907 ) );
  CLKMX2X2 U12095 ( .A(n5423), .B(\i_MIPS/Register/register[7][22] ), .S0(
        n5606), .Y(\i_MIPS/Register/n906 ) );
  CLKMX2X2 U12096 ( .A(n5432), .B(\i_MIPS/Register/register[7][19] ), .S0(
        n5606), .Y(\i_MIPS/Register/n903 ) );
  CLKMX2X2 U12097 ( .A(n5417), .B(\i_MIPS/Register/register[7][18] ), .S0(
        n5607), .Y(\i_MIPS/Register/n902 ) );
  CLKMX2X2 U12098 ( .A(n5458), .B(\i_MIPS/Register/register[7][17] ), .S0(
        n5607), .Y(\i_MIPS/Register/n901 ) );
  CLKMX2X2 U12099 ( .A(n5456), .B(\i_MIPS/Register/register[7][15] ), .S0(
        n5607), .Y(\i_MIPS/Register/n899 ) );
  CLKMX2X2 U12100 ( .A(n5454), .B(\i_MIPS/Register/register[7][14] ), .S0(
        n5607), .Y(\i_MIPS/Register/n898 ) );
  CLKMX2X2 U12101 ( .A(n5452), .B(\i_MIPS/Register/register[7][13] ), .S0(
        n5607), .Y(\i_MIPS/Register/n897 ) );
  CLKMX2X2 U12102 ( .A(n5449), .B(\i_MIPS/Register/register[7][12] ), .S0(
        n5607), .Y(\i_MIPS/Register/n896 ) );
  CLKMX2X2 U12103 ( .A(n5446), .B(\i_MIPS/Register/register[7][11] ), .S0(
        n5606), .Y(\i_MIPS/Register/n895 ) );
  CLKMX2X2 U12104 ( .A(n5420), .B(\i_MIPS/Register/register[7][10] ), .S0(
        n5606), .Y(\i_MIPS/Register/n894 ) );
  CLKMX2X2 U12105 ( .A(n5475), .B(\i_MIPS/Register/register[7][8] ), .S0(n5607), .Y(\i_MIPS/Register/n892 ) );
  CLKMX2X2 U12106 ( .A(n5472), .B(\i_MIPS/Register/register[7][7] ), .S0(n5607), .Y(\i_MIPS/Register/n891 ) );
  CLKMX2X2 U12107 ( .A(n5043), .B(\i_MIPS/Register/register[7][6] ), .S0(n5606), .Y(\i_MIPS/Register/n890 ) );
  CLKMX2X2 U12108 ( .A(n5491), .B(\i_MIPS/Register/register[7][5] ), .S0(n5606), .Y(\i_MIPS/Register/n889 ) );
  CLKMX2X2 U12109 ( .A(n5488), .B(\i_MIPS/Register/register[7][4] ), .S0(n5606), .Y(\i_MIPS/Register/n888 ) );
  CLKMX2X2 U12110 ( .A(n4776), .B(\i_MIPS/Register/register[7][3] ), .S0(n5606), .Y(\i_MIPS/Register/n887 ) );
  CLKMX2X2 U12111 ( .A(n5480), .B(\i_MIPS/Register/register[7][2] ), .S0(n5606), .Y(\i_MIPS/Register/n886 ) );
  CLKMX2X2 U12112 ( .A(n5477), .B(\i_MIPS/Register/register[7][1] ), .S0(n5607), .Y(\i_MIPS/Register/n885 ) );
  CLKMX2X2 U12113 ( .A(n5485), .B(\i_MIPS/Register/register[7][0] ), .S0(n5607), .Y(\i_MIPS/Register/n884 ) );
  CLKMX2X2 U12114 ( .A(n5469), .B(\i_MIPS/Register/register[8][31] ), .S0(
        n5604), .Y(\i_MIPS/Register/n883 ) );
  CLKMX2X2 U12115 ( .A(n5410), .B(\i_MIPS/Register/register[8][28] ), .S0(
        n5605), .Y(\i_MIPS/Register/n880 ) );
  CLKMX2X2 U12116 ( .A(n5407), .B(\i_MIPS/Register/register[8][27] ), .S0(
        n5604), .Y(\i_MIPS/Register/n879 ) );
  CLKMX2X2 U12117 ( .A(n5404), .B(\i_MIPS/Register/register[8][26] ), .S0(
        n5604), .Y(\i_MIPS/Register/n878 ) );
  CLKMX2X2 U12118 ( .A(n5413), .B(\i_MIPS/Register/register[8][25] ), .S0(
        n5605), .Y(\i_MIPS/Register/n877 ) );
  CLKMX2X2 U12119 ( .A(n5482), .B(\i_MIPS/Register/register[8][23] ), .S0(
        n5605), .Y(\i_MIPS/Register/n875 ) );
  CLKMX2X2 U12120 ( .A(n5422), .B(\i_MIPS/Register/register[8][22] ), .S0(
        n5604), .Y(\i_MIPS/Register/n874 ) );
  CLKMX2X2 U12121 ( .A(n5431), .B(\i_MIPS/Register/register[8][19] ), .S0(
        n5604), .Y(\i_MIPS/Register/n871 ) );
  CLKMX2X2 U12122 ( .A(n5416), .B(\i_MIPS/Register/register[8][18] ), .S0(
        n5605), .Y(\i_MIPS/Register/n870 ) );
  CLKMX2X2 U12123 ( .A(n5457), .B(\i_MIPS/Register/register[8][17] ), .S0(
        n5605), .Y(\i_MIPS/Register/n869 ) );
  CLKMX2X2 U12124 ( .A(n5455), .B(\i_MIPS/Register/register[8][15] ), .S0(
        n5605), .Y(\i_MIPS/Register/n867 ) );
  CLKMX2X2 U12125 ( .A(n5453), .B(\i_MIPS/Register/register[8][14] ), .S0(
        n5605), .Y(\i_MIPS/Register/n866 ) );
  CLKMX2X2 U12126 ( .A(n5451), .B(\i_MIPS/Register/register[8][13] ), .S0(
        n5605), .Y(\i_MIPS/Register/n865 ) );
  CLKMX2X2 U12127 ( .A(n5448), .B(\i_MIPS/Register/register[8][12] ), .S0(
        n5605), .Y(\i_MIPS/Register/n864 ) );
  CLKMX2X2 U12128 ( .A(n5445), .B(\i_MIPS/Register/register[8][11] ), .S0(
        n5604), .Y(\i_MIPS/Register/n863 ) );
  CLKMX2X2 U12129 ( .A(n5419), .B(\i_MIPS/Register/register[8][10] ), .S0(
        n5604), .Y(\i_MIPS/Register/n862 ) );
  CLKMX2X2 U12130 ( .A(n5474), .B(\i_MIPS/Register/register[8][8] ), .S0(n5605), .Y(\i_MIPS/Register/n860 ) );
  CLKMX2X2 U12131 ( .A(n5471), .B(\i_MIPS/Register/register[8][7] ), .S0(n5605), .Y(\i_MIPS/Register/n859 ) );
  CLKMX2X2 U12132 ( .A(n5042), .B(\i_MIPS/Register/register[8][6] ), .S0(n5604), .Y(\i_MIPS/Register/n858 ) );
  CLKMX2X2 U12133 ( .A(n5490), .B(\i_MIPS/Register/register[8][5] ), .S0(n5604), .Y(\i_MIPS/Register/n857 ) );
  CLKMX2X2 U12134 ( .A(n5487), .B(\i_MIPS/Register/register[8][4] ), .S0(n5604), .Y(\i_MIPS/Register/n856 ) );
  CLKMX2X2 U12135 ( .A(n4775), .B(\i_MIPS/Register/register[8][3] ), .S0(n5604), .Y(\i_MIPS/Register/n855 ) );
  CLKMX2X2 U12136 ( .A(n5479), .B(\i_MIPS/Register/register[8][2] ), .S0(n5604), .Y(\i_MIPS/Register/n854 ) );
  CLKMX2X2 U12137 ( .A(n5476), .B(\i_MIPS/Register/register[8][1] ), .S0(n5605), .Y(\i_MIPS/Register/n853 ) );
  CLKMX2X2 U12138 ( .A(n5484), .B(\i_MIPS/Register/register[8][0] ), .S0(n5605), .Y(\i_MIPS/Register/n852 ) );
  CLKMX2X2 U12139 ( .A(n5469), .B(\i_MIPS/Register/register[9][31] ), .S0(
        n5602), .Y(\i_MIPS/Register/n851 ) );
  CLKMX2X2 U12140 ( .A(n5410), .B(\i_MIPS/Register/register[9][28] ), .S0(
        n5603), .Y(\i_MIPS/Register/n848 ) );
  CLKMX2X2 U12141 ( .A(n5407), .B(\i_MIPS/Register/register[9][27] ), .S0(
        n5602), .Y(\i_MIPS/Register/n847 ) );
  CLKMX2X2 U12142 ( .A(n5404), .B(\i_MIPS/Register/register[9][26] ), .S0(
        n5602), .Y(\i_MIPS/Register/n846 ) );
  CLKMX2X2 U12143 ( .A(n5413), .B(\i_MIPS/Register/register[9][25] ), .S0(
        n5603), .Y(\i_MIPS/Register/n845 ) );
  CLKMX2X2 U12144 ( .A(n5482), .B(\i_MIPS/Register/register[9][23] ), .S0(
        n5603), .Y(\i_MIPS/Register/n843 ) );
  CLKMX2X2 U12145 ( .A(n5422), .B(\i_MIPS/Register/register[9][22] ), .S0(
        n5602), .Y(\i_MIPS/Register/n842 ) );
  CLKMX2X2 U12146 ( .A(n5431), .B(\i_MIPS/Register/register[9][19] ), .S0(
        n5602), .Y(\i_MIPS/Register/n839 ) );
  CLKMX2X2 U12147 ( .A(n5416), .B(\i_MIPS/Register/register[9][18] ), .S0(
        n5603), .Y(\i_MIPS/Register/n838 ) );
  CLKMX2X2 U12148 ( .A(n5457), .B(\i_MIPS/Register/register[9][17] ), .S0(
        n5603), .Y(\i_MIPS/Register/n837 ) );
  CLKMX2X2 U12149 ( .A(n5455), .B(\i_MIPS/Register/register[9][15] ), .S0(
        n5603), .Y(\i_MIPS/Register/n835 ) );
  CLKMX2X2 U12150 ( .A(n5453), .B(\i_MIPS/Register/register[9][14] ), .S0(
        n5603), .Y(\i_MIPS/Register/n834 ) );
  CLKMX2X2 U12151 ( .A(n5451), .B(\i_MIPS/Register/register[9][13] ), .S0(
        n5603), .Y(\i_MIPS/Register/n833 ) );
  CLKMX2X2 U12152 ( .A(n5448), .B(\i_MIPS/Register/register[9][12] ), .S0(
        n5603), .Y(\i_MIPS/Register/n832 ) );
  CLKMX2X2 U12153 ( .A(n5445), .B(\i_MIPS/Register/register[9][11] ), .S0(
        n5602), .Y(\i_MIPS/Register/n831 ) );
  CLKMX2X2 U12154 ( .A(n5419), .B(\i_MIPS/Register/register[9][10] ), .S0(
        n5602), .Y(\i_MIPS/Register/n830 ) );
  CLKMX2X2 U12155 ( .A(n5474), .B(\i_MIPS/Register/register[9][8] ), .S0(n5603), .Y(\i_MIPS/Register/n828 ) );
  CLKMX2X2 U12156 ( .A(n5471), .B(\i_MIPS/Register/register[9][7] ), .S0(n5603), .Y(\i_MIPS/Register/n827 ) );
  CLKMX2X2 U12157 ( .A(n5042), .B(\i_MIPS/Register/register[9][6] ), .S0(n5602), .Y(\i_MIPS/Register/n826 ) );
  CLKMX2X2 U12158 ( .A(n5490), .B(\i_MIPS/Register/register[9][5] ), .S0(n5602), .Y(\i_MIPS/Register/n825 ) );
  CLKMX2X2 U12159 ( .A(n5487), .B(\i_MIPS/Register/register[9][4] ), .S0(n5602), .Y(\i_MIPS/Register/n824 ) );
  CLKMX2X2 U12160 ( .A(n4775), .B(\i_MIPS/Register/register[9][3] ), .S0(n5602), .Y(\i_MIPS/Register/n823 ) );
  CLKMX2X2 U12161 ( .A(n5479), .B(\i_MIPS/Register/register[9][2] ), .S0(n5602), .Y(\i_MIPS/Register/n822 ) );
  CLKMX2X2 U12162 ( .A(n5476), .B(\i_MIPS/Register/register[9][1] ), .S0(n5603), .Y(\i_MIPS/Register/n821 ) );
  CLKMX2X2 U12163 ( .A(n5484), .B(\i_MIPS/Register/register[9][0] ), .S0(n5603), .Y(\i_MIPS/Register/n820 ) );
  CLKMX2X2 U12164 ( .A(n5469), .B(\i_MIPS/Register/register[10][31] ), .S0(
        n5600), .Y(\i_MIPS/Register/n819 ) );
  CLKMX2X2 U12165 ( .A(n5410), .B(\i_MIPS/Register/register[10][28] ), .S0(
        n5601), .Y(\i_MIPS/Register/n816 ) );
  CLKMX2X2 U12166 ( .A(n5407), .B(\i_MIPS/Register/register[10][27] ), .S0(
        n5600), .Y(\i_MIPS/Register/n815 ) );
  CLKMX2X2 U12167 ( .A(n5404), .B(\i_MIPS/Register/register[10][26] ), .S0(
        n5600), .Y(\i_MIPS/Register/n814 ) );
  CLKMX2X2 U12168 ( .A(n5413), .B(\i_MIPS/Register/register[10][25] ), .S0(
        n5601), .Y(\i_MIPS/Register/n813 ) );
  CLKMX2X2 U12169 ( .A(n5482), .B(\i_MIPS/Register/register[10][23] ), .S0(
        n5601), .Y(\i_MIPS/Register/n811 ) );
  CLKMX2X2 U12170 ( .A(n5422), .B(\i_MIPS/Register/register[10][22] ), .S0(
        n5600), .Y(\i_MIPS/Register/n810 ) );
  CLKMX2X2 U12171 ( .A(n5431), .B(\i_MIPS/Register/register[10][19] ), .S0(
        n5600), .Y(\i_MIPS/Register/n807 ) );
  CLKMX2X2 U12172 ( .A(n5416), .B(\i_MIPS/Register/register[10][18] ), .S0(
        n5601), .Y(\i_MIPS/Register/n806 ) );
  CLKMX2X2 U12173 ( .A(n5457), .B(\i_MIPS/Register/register[10][17] ), .S0(
        n5601), .Y(\i_MIPS/Register/n805 ) );
  CLKMX2X2 U12174 ( .A(n5455), .B(\i_MIPS/Register/register[10][15] ), .S0(
        n5601), .Y(\i_MIPS/Register/n803 ) );
  CLKMX2X2 U12175 ( .A(n5453), .B(\i_MIPS/Register/register[10][14] ), .S0(
        n5601), .Y(\i_MIPS/Register/n802 ) );
  CLKMX2X2 U12176 ( .A(n5451), .B(\i_MIPS/Register/register[10][13] ), .S0(
        n5601), .Y(\i_MIPS/Register/n801 ) );
  CLKMX2X2 U12177 ( .A(n5448), .B(\i_MIPS/Register/register[10][12] ), .S0(
        n5601), .Y(\i_MIPS/Register/n800 ) );
  CLKMX2X2 U12178 ( .A(n5445), .B(\i_MIPS/Register/register[10][11] ), .S0(
        n5600), .Y(\i_MIPS/Register/n799 ) );
  CLKMX2X2 U12179 ( .A(n5419), .B(\i_MIPS/Register/register[10][10] ), .S0(
        n5600), .Y(\i_MIPS/Register/n798 ) );
  CLKMX2X2 U12180 ( .A(n5474), .B(\i_MIPS/Register/register[10][8] ), .S0(
        n5601), .Y(\i_MIPS/Register/n796 ) );
  CLKMX2X2 U12181 ( .A(n5471), .B(\i_MIPS/Register/register[10][7] ), .S0(
        n5601), .Y(\i_MIPS/Register/n795 ) );
  CLKMX2X2 U12182 ( .A(n5042), .B(\i_MIPS/Register/register[10][6] ), .S0(
        n5600), .Y(\i_MIPS/Register/n794 ) );
  CLKMX2X2 U12183 ( .A(n5490), .B(\i_MIPS/Register/register[10][5] ), .S0(
        n5600), .Y(\i_MIPS/Register/n793 ) );
  CLKMX2X2 U12184 ( .A(n5487), .B(\i_MIPS/Register/register[10][4] ), .S0(
        n5600), .Y(\i_MIPS/Register/n792 ) );
  CLKMX2X2 U12185 ( .A(n4775), .B(\i_MIPS/Register/register[10][3] ), .S0(
        n5600), .Y(\i_MIPS/Register/n791 ) );
  CLKMX2X2 U12186 ( .A(n5479), .B(\i_MIPS/Register/register[10][2] ), .S0(
        n5600), .Y(\i_MIPS/Register/n790 ) );
  CLKMX2X2 U12187 ( .A(n5476), .B(\i_MIPS/Register/register[10][1] ), .S0(
        n5601), .Y(\i_MIPS/Register/n789 ) );
  CLKMX2X2 U12188 ( .A(n5484), .B(\i_MIPS/Register/register[10][0] ), .S0(
        n5601), .Y(\i_MIPS/Register/n788 ) );
  CLKMX2X2 U12189 ( .A(n5469), .B(\i_MIPS/Register/register[11][31] ), .S0(
        n5598), .Y(\i_MIPS/Register/n787 ) );
  CLKMX2X2 U12190 ( .A(n5411), .B(\i_MIPS/Register/register[11][28] ), .S0(
        n5599), .Y(\i_MIPS/Register/n784 ) );
  CLKMX2X2 U12191 ( .A(n5408), .B(\i_MIPS/Register/register[11][27] ), .S0(
        n5598), .Y(\i_MIPS/Register/n783 ) );
  CLKMX2X2 U12192 ( .A(n5404), .B(\i_MIPS/Register/register[11][26] ), .S0(
        n5598), .Y(\i_MIPS/Register/n782 ) );
  CLKMX2X2 U12193 ( .A(n5414), .B(\i_MIPS/Register/register[11][25] ), .S0(
        n5599), .Y(\i_MIPS/Register/n781 ) );
  CLKMX2X2 U12194 ( .A(n5482), .B(\i_MIPS/Register/register[11][23] ), .S0(
        n5599), .Y(\i_MIPS/Register/n779 ) );
  CLKMX2X2 U12195 ( .A(n5422), .B(\i_MIPS/Register/register[11][22] ), .S0(
        n5598), .Y(\i_MIPS/Register/n778 ) );
  CLKMX2X2 U12196 ( .A(n5432), .B(\i_MIPS/Register/register[11][19] ), .S0(
        n5598), .Y(\i_MIPS/Register/n775 ) );
  CLKMX2X2 U12197 ( .A(n5417), .B(\i_MIPS/Register/register[11][18] ), .S0(
        n5599), .Y(\i_MIPS/Register/n774 ) );
  CLKMX2X2 U12198 ( .A(n5457), .B(\i_MIPS/Register/register[11][17] ), .S0(
        n5599), .Y(\i_MIPS/Register/n773 ) );
  CLKMX2X2 U12199 ( .A(n5455), .B(\i_MIPS/Register/register[11][15] ), .S0(
        n5599), .Y(\i_MIPS/Register/n771 ) );
  CLKMX2X2 U12200 ( .A(n5453), .B(\i_MIPS/Register/register[11][14] ), .S0(
        n5599), .Y(\i_MIPS/Register/n770 ) );
  CLKMX2X2 U12201 ( .A(n5451), .B(\i_MIPS/Register/register[11][13] ), .S0(
        n5599), .Y(\i_MIPS/Register/n769 ) );
  CLKMX2X2 U12202 ( .A(n5448), .B(\i_MIPS/Register/register[11][12] ), .S0(
        n5599), .Y(\i_MIPS/Register/n768 ) );
  CLKMX2X2 U12203 ( .A(n5445), .B(\i_MIPS/Register/register[11][11] ), .S0(
        n5598), .Y(\i_MIPS/Register/n767 ) );
  CLKMX2X2 U12204 ( .A(n5419), .B(\i_MIPS/Register/register[11][10] ), .S0(
        n5598), .Y(\i_MIPS/Register/n766 ) );
  CLKMX2X2 U12205 ( .A(n5474), .B(\i_MIPS/Register/register[11][8] ), .S0(
        n5599), .Y(\i_MIPS/Register/n764 ) );
  CLKMX2X2 U12206 ( .A(n5471), .B(\i_MIPS/Register/register[11][7] ), .S0(
        n5599), .Y(\i_MIPS/Register/n763 ) );
  CLKMX2X2 U12207 ( .A(n5043), .B(\i_MIPS/Register/register[11][6] ), .S0(
        n5598), .Y(\i_MIPS/Register/n762 ) );
  CLKMX2X2 U12208 ( .A(n5490), .B(\i_MIPS/Register/register[11][5] ), .S0(
        n5598), .Y(\i_MIPS/Register/n761 ) );
  CLKMX2X2 U12209 ( .A(n5487), .B(\i_MIPS/Register/register[11][4] ), .S0(
        n5598), .Y(\i_MIPS/Register/n760 ) );
  CLKMX2X2 U12210 ( .A(n4776), .B(\i_MIPS/Register/register[11][3] ), .S0(
        n5598), .Y(\i_MIPS/Register/n759 ) );
  CLKMX2X2 U12211 ( .A(n5479), .B(\i_MIPS/Register/register[11][2] ), .S0(
        n5598), .Y(\i_MIPS/Register/n758 ) );
  CLKMX2X2 U12212 ( .A(n5476), .B(\i_MIPS/Register/register[11][1] ), .S0(
        n5599), .Y(\i_MIPS/Register/n757 ) );
  CLKMX2X2 U12213 ( .A(n5484), .B(\i_MIPS/Register/register[11][0] ), .S0(
        n5599), .Y(\i_MIPS/Register/n756 ) );
  CLKMX2X2 U12214 ( .A(n5469), .B(\i_MIPS/Register/register[12][31] ), .S0(
        n5596), .Y(\i_MIPS/Register/n755 ) );
  CLKMX2X2 U12215 ( .A(n5410), .B(\i_MIPS/Register/register[12][28] ), .S0(
        n5597), .Y(\i_MIPS/Register/n752 ) );
  CLKMX2X2 U12216 ( .A(n5407), .B(\i_MIPS/Register/register[12][27] ), .S0(
        n5596), .Y(\i_MIPS/Register/n751 ) );
  CLKMX2X2 U12217 ( .A(n5404), .B(\i_MIPS/Register/register[12][26] ), .S0(
        n5596), .Y(\i_MIPS/Register/n750 ) );
  CLKMX2X2 U12218 ( .A(n5413), .B(\i_MIPS/Register/register[12][25] ), .S0(
        n5597), .Y(\i_MIPS/Register/n749 ) );
  CLKMX2X2 U12219 ( .A(n5482), .B(\i_MIPS/Register/register[12][23] ), .S0(
        n5597), .Y(\i_MIPS/Register/n747 ) );
  CLKMX2X2 U12220 ( .A(n5422), .B(\i_MIPS/Register/register[12][22] ), .S0(
        n5596), .Y(\i_MIPS/Register/n746 ) );
  CLKMX2X2 U12221 ( .A(n5431), .B(\i_MIPS/Register/register[12][19] ), .S0(
        n5596), .Y(\i_MIPS/Register/n743 ) );
  CLKMX2X2 U12222 ( .A(n5416), .B(\i_MIPS/Register/register[12][18] ), .S0(
        n5597), .Y(\i_MIPS/Register/n742 ) );
  CLKMX2X2 U12223 ( .A(n5457), .B(\i_MIPS/Register/register[12][17] ), .S0(
        n5597), .Y(\i_MIPS/Register/n741 ) );
  CLKMX2X2 U12224 ( .A(n5455), .B(\i_MIPS/Register/register[12][15] ), .S0(
        n5597), .Y(\i_MIPS/Register/n739 ) );
  CLKMX2X2 U12225 ( .A(n5453), .B(\i_MIPS/Register/register[12][14] ), .S0(
        n5597), .Y(\i_MIPS/Register/n738 ) );
  CLKMX2X2 U12226 ( .A(n5451), .B(\i_MIPS/Register/register[12][13] ), .S0(
        n5597), .Y(\i_MIPS/Register/n737 ) );
  CLKMX2X2 U12227 ( .A(n5448), .B(\i_MIPS/Register/register[12][12] ), .S0(
        n5597), .Y(\i_MIPS/Register/n736 ) );
  CLKMX2X2 U12228 ( .A(n5445), .B(\i_MIPS/Register/register[12][11] ), .S0(
        n5596), .Y(\i_MIPS/Register/n735 ) );
  CLKMX2X2 U12229 ( .A(n5419), .B(\i_MIPS/Register/register[12][10] ), .S0(
        n5596), .Y(\i_MIPS/Register/n734 ) );
  CLKMX2X2 U12230 ( .A(n5474), .B(\i_MIPS/Register/register[12][8] ), .S0(
        n5597), .Y(\i_MIPS/Register/n732 ) );
  CLKMX2X2 U12231 ( .A(n5471), .B(\i_MIPS/Register/register[12][7] ), .S0(
        n5597), .Y(\i_MIPS/Register/n731 ) );
  CLKMX2X2 U12232 ( .A(n5042), .B(\i_MIPS/Register/register[12][6] ), .S0(
        n5596), .Y(\i_MIPS/Register/n730 ) );
  CLKMX2X2 U12233 ( .A(n5490), .B(\i_MIPS/Register/register[12][5] ), .S0(
        n5596), .Y(\i_MIPS/Register/n729 ) );
  CLKMX2X2 U12234 ( .A(n5487), .B(\i_MIPS/Register/register[12][4] ), .S0(
        n5596), .Y(\i_MIPS/Register/n728 ) );
  CLKMX2X2 U12235 ( .A(n4775), .B(\i_MIPS/Register/register[12][3] ), .S0(
        n5596), .Y(\i_MIPS/Register/n727 ) );
  CLKMX2X2 U12236 ( .A(n5479), .B(\i_MIPS/Register/register[12][2] ), .S0(
        n5596), .Y(\i_MIPS/Register/n726 ) );
  CLKMX2X2 U12237 ( .A(n5476), .B(\i_MIPS/Register/register[12][1] ), .S0(
        n5597), .Y(\i_MIPS/Register/n725 ) );
  CLKMX2X2 U12238 ( .A(n5484), .B(\i_MIPS/Register/register[12][0] ), .S0(
        n5597), .Y(\i_MIPS/Register/n724 ) );
  CLKMX2X2 U12239 ( .A(n5469), .B(\i_MIPS/Register/register[13][31] ), .S0(
        n5594), .Y(\i_MIPS/Register/n723 ) );
  CLKMX2X2 U12240 ( .A(n5410), .B(\i_MIPS/Register/register[13][28] ), .S0(
        n5595), .Y(\i_MIPS/Register/n720 ) );
  CLKMX2X2 U12241 ( .A(n5407), .B(\i_MIPS/Register/register[13][27] ), .S0(
        n5594), .Y(\i_MIPS/Register/n719 ) );
  CLKMX2X2 U12242 ( .A(n5404), .B(\i_MIPS/Register/register[13][26] ), .S0(
        n5594), .Y(\i_MIPS/Register/n718 ) );
  CLKMX2X2 U12243 ( .A(n5413), .B(\i_MIPS/Register/register[13][25] ), .S0(
        n5595), .Y(\i_MIPS/Register/n717 ) );
  CLKMX2X2 U12244 ( .A(n5482), .B(\i_MIPS/Register/register[13][23] ), .S0(
        n5595), .Y(\i_MIPS/Register/n715 ) );
  CLKMX2X2 U12245 ( .A(n5422), .B(\i_MIPS/Register/register[13][22] ), .S0(
        n5594), .Y(\i_MIPS/Register/n714 ) );
  CLKMX2X2 U12246 ( .A(n5431), .B(\i_MIPS/Register/register[13][19] ), .S0(
        n5594), .Y(\i_MIPS/Register/n711 ) );
  CLKMX2X2 U12247 ( .A(n5416), .B(\i_MIPS/Register/register[13][18] ), .S0(
        n5595), .Y(\i_MIPS/Register/n710 ) );
  CLKMX2X2 U12248 ( .A(n5457), .B(\i_MIPS/Register/register[13][17] ), .S0(
        n5595), .Y(\i_MIPS/Register/n709 ) );
  CLKMX2X2 U12249 ( .A(n5455), .B(\i_MIPS/Register/register[13][15] ), .S0(
        n5595), .Y(\i_MIPS/Register/n707 ) );
  CLKMX2X2 U12250 ( .A(n5453), .B(\i_MIPS/Register/register[13][14] ), .S0(
        n5595), .Y(\i_MIPS/Register/n706 ) );
  CLKMX2X2 U12251 ( .A(n5451), .B(\i_MIPS/Register/register[13][13] ), .S0(
        n5595), .Y(\i_MIPS/Register/n705 ) );
  CLKMX2X2 U12252 ( .A(n5448), .B(\i_MIPS/Register/register[13][12] ), .S0(
        n5595), .Y(\i_MIPS/Register/n704 ) );
  CLKMX2X2 U12253 ( .A(n5445), .B(\i_MIPS/Register/register[13][11] ), .S0(
        n5594), .Y(\i_MIPS/Register/n703 ) );
  CLKMX2X2 U12254 ( .A(n5419), .B(\i_MIPS/Register/register[13][10] ), .S0(
        n5594), .Y(\i_MIPS/Register/n702 ) );
  CLKMX2X2 U12255 ( .A(n5474), .B(\i_MIPS/Register/register[13][8] ), .S0(
        n5595), .Y(\i_MIPS/Register/n700 ) );
  CLKMX2X2 U12256 ( .A(n5471), .B(\i_MIPS/Register/register[13][7] ), .S0(
        n5595), .Y(\i_MIPS/Register/n699 ) );
  CLKMX2X2 U12257 ( .A(n5042), .B(\i_MIPS/Register/register[13][6] ), .S0(
        n5594), .Y(\i_MIPS/Register/n698 ) );
  CLKMX2X2 U12258 ( .A(n5490), .B(\i_MIPS/Register/register[13][5] ), .S0(
        n5594), .Y(\i_MIPS/Register/n697 ) );
  CLKMX2X2 U12259 ( .A(n5487), .B(\i_MIPS/Register/register[13][4] ), .S0(
        n5594), .Y(\i_MIPS/Register/n696 ) );
  CLKMX2X2 U12260 ( .A(n4775), .B(\i_MIPS/Register/register[13][3] ), .S0(
        n5594), .Y(\i_MIPS/Register/n695 ) );
  CLKMX2X2 U12261 ( .A(n5479), .B(\i_MIPS/Register/register[13][2] ), .S0(
        n5594), .Y(\i_MIPS/Register/n694 ) );
  CLKMX2X2 U12262 ( .A(n5476), .B(\i_MIPS/Register/register[13][1] ), .S0(
        n5595), .Y(\i_MIPS/Register/n693 ) );
  CLKMX2X2 U12263 ( .A(n5484), .B(\i_MIPS/Register/register[13][0] ), .S0(
        n5595), .Y(\i_MIPS/Register/n692 ) );
  CLKMX2X2 U12264 ( .A(n5469), .B(\i_MIPS/Register/register[14][31] ), .S0(
        n5592), .Y(\i_MIPS/Register/n691 ) );
  CLKMX2X2 U12265 ( .A(n5410), .B(\i_MIPS/Register/register[14][28] ), .S0(
        n5593), .Y(\i_MIPS/Register/n688 ) );
  CLKMX2X2 U12266 ( .A(n5407), .B(\i_MIPS/Register/register[14][27] ), .S0(
        n5592), .Y(\i_MIPS/Register/n687 ) );
  CLKMX2X2 U12267 ( .A(n5404), .B(\i_MIPS/Register/register[14][26] ), .S0(
        n5592), .Y(\i_MIPS/Register/n686 ) );
  CLKMX2X2 U12268 ( .A(n5413), .B(\i_MIPS/Register/register[14][25] ), .S0(
        n5593), .Y(\i_MIPS/Register/n685 ) );
  CLKMX2X2 U12269 ( .A(n5482), .B(\i_MIPS/Register/register[14][23] ), .S0(
        n5593), .Y(\i_MIPS/Register/n683 ) );
  CLKMX2X2 U12270 ( .A(n5422), .B(\i_MIPS/Register/register[14][22] ), .S0(
        n5592), .Y(\i_MIPS/Register/n682 ) );
  CLKMX2X2 U12271 ( .A(n5431), .B(\i_MIPS/Register/register[14][19] ), .S0(
        n5592), .Y(\i_MIPS/Register/n679 ) );
  CLKMX2X2 U12272 ( .A(n5416), .B(\i_MIPS/Register/register[14][18] ), .S0(
        n5593), .Y(\i_MIPS/Register/n678 ) );
  CLKMX2X2 U12273 ( .A(n5457), .B(\i_MIPS/Register/register[14][17] ), .S0(
        n5593), .Y(\i_MIPS/Register/n677 ) );
  CLKMX2X2 U12274 ( .A(n5455), .B(\i_MIPS/Register/register[14][15] ), .S0(
        n5593), .Y(\i_MIPS/Register/n675 ) );
  CLKMX2X2 U12275 ( .A(n5453), .B(\i_MIPS/Register/register[14][14] ), .S0(
        n5593), .Y(\i_MIPS/Register/n674 ) );
  CLKMX2X2 U12276 ( .A(n5451), .B(\i_MIPS/Register/register[14][13] ), .S0(
        n5593), .Y(\i_MIPS/Register/n673 ) );
  CLKMX2X2 U12277 ( .A(n5448), .B(\i_MIPS/Register/register[14][12] ), .S0(
        n5593), .Y(\i_MIPS/Register/n672 ) );
  CLKMX2X2 U12278 ( .A(n5445), .B(\i_MIPS/Register/register[14][11] ), .S0(
        n5592), .Y(\i_MIPS/Register/n671 ) );
  CLKMX2X2 U12279 ( .A(n5419), .B(\i_MIPS/Register/register[14][10] ), .S0(
        n5592), .Y(\i_MIPS/Register/n670 ) );
  CLKMX2X2 U12280 ( .A(n5474), .B(\i_MIPS/Register/register[14][8] ), .S0(
        n5593), .Y(\i_MIPS/Register/n668 ) );
  CLKMX2X2 U12281 ( .A(n5471), .B(\i_MIPS/Register/register[14][7] ), .S0(
        n5593), .Y(\i_MIPS/Register/n667 ) );
  CLKMX2X2 U12282 ( .A(n5042), .B(\i_MIPS/Register/register[14][6] ), .S0(
        n5592), .Y(\i_MIPS/Register/n666 ) );
  CLKMX2X2 U12283 ( .A(n5490), .B(\i_MIPS/Register/register[14][5] ), .S0(
        n5592), .Y(\i_MIPS/Register/n665 ) );
  CLKMX2X2 U12284 ( .A(n5487), .B(\i_MIPS/Register/register[14][4] ), .S0(
        n5592), .Y(\i_MIPS/Register/n664 ) );
  CLKMX2X2 U12285 ( .A(n4775), .B(\i_MIPS/Register/register[14][3] ), .S0(
        n5592), .Y(\i_MIPS/Register/n663 ) );
  CLKMX2X2 U12286 ( .A(n5479), .B(\i_MIPS/Register/register[14][2] ), .S0(
        n5592), .Y(\i_MIPS/Register/n662 ) );
  CLKMX2X2 U12287 ( .A(n5476), .B(\i_MIPS/Register/register[14][1] ), .S0(
        n5593), .Y(\i_MIPS/Register/n661 ) );
  CLKMX2X2 U12288 ( .A(n5484), .B(\i_MIPS/Register/register[14][0] ), .S0(
        n5593), .Y(\i_MIPS/Register/n660 ) );
  CLKMX2X2 U12289 ( .A(n5470), .B(\i_MIPS/Register/register[15][31] ), .S0(
        n5590), .Y(\i_MIPS/Register/n659 ) );
  CLKMX2X2 U12290 ( .A(n5411), .B(\i_MIPS/Register/register[15][28] ), .S0(
        n5591), .Y(\i_MIPS/Register/n656 ) );
  CLKMX2X2 U12291 ( .A(n5408), .B(\i_MIPS/Register/register[15][27] ), .S0(
        n5590), .Y(\i_MIPS/Register/n655 ) );
  CLKMX2X2 U12292 ( .A(n5405), .B(\i_MIPS/Register/register[15][26] ), .S0(
        n5590), .Y(\i_MIPS/Register/n654 ) );
  CLKMX2X2 U12293 ( .A(n5414), .B(\i_MIPS/Register/register[15][25] ), .S0(
        n5591), .Y(\i_MIPS/Register/n653 ) );
  CLKMX2X2 U12294 ( .A(n5483), .B(\i_MIPS/Register/register[15][23] ), .S0(
        n5591), .Y(\i_MIPS/Register/n651 ) );
  CLKMX2X2 U12295 ( .A(n5423), .B(\i_MIPS/Register/register[15][22] ), .S0(
        n5590), .Y(\i_MIPS/Register/n650 ) );
  CLKMX2X2 U12296 ( .A(n5432), .B(\i_MIPS/Register/register[15][19] ), .S0(
        n5590), .Y(\i_MIPS/Register/n647 ) );
  CLKMX2X2 U12297 ( .A(n5417), .B(\i_MIPS/Register/register[15][18] ), .S0(
        n5591), .Y(\i_MIPS/Register/n646 ) );
  CLKMX2X2 U12298 ( .A(n5458), .B(\i_MIPS/Register/register[15][17] ), .S0(
        n5591), .Y(\i_MIPS/Register/n645 ) );
  CLKMX2X2 U12299 ( .A(n5456), .B(\i_MIPS/Register/register[15][15] ), .S0(
        n5591), .Y(\i_MIPS/Register/n643 ) );
  CLKMX2X2 U12300 ( .A(n5454), .B(\i_MIPS/Register/register[15][14] ), .S0(
        n5591), .Y(\i_MIPS/Register/n642 ) );
  CLKMX2X2 U12301 ( .A(n5452), .B(\i_MIPS/Register/register[15][13] ), .S0(
        n5591), .Y(\i_MIPS/Register/n641 ) );
  CLKMX2X2 U12302 ( .A(n5449), .B(\i_MIPS/Register/register[15][12] ), .S0(
        n5591), .Y(\i_MIPS/Register/n640 ) );
  CLKMX2X2 U12303 ( .A(n5446), .B(\i_MIPS/Register/register[15][11] ), .S0(
        n5590), .Y(\i_MIPS/Register/n639 ) );
  CLKMX2X2 U12304 ( .A(n5420), .B(\i_MIPS/Register/register[15][10] ), .S0(
        n5590), .Y(\i_MIPS/Register/n638 ) );
  CLKMX2X2 U12305 ( .A(n5475), .B(\i_MIPS/Register/register[15][8] ), .S0(
        n5591), .Y(\i_MIPS/Register/n636 ) );
  CLKMX2X2 U12306 ( .A(n5472), .B(\i_MIPS/Register/register[15][7] ), .S0(
        n5591), .Y(\i_MIPS/Register/n635 ) );
  CLKMX2X2 U12307 ( .A(n5043), .B(\i_MIPS/Register/register[15][6] ), .S0(
        n5590), .Y(\i_MIPS/Register/n634 ) );
  CLKMX2X2 U12308 ( .A(n5491), .B(\i_MIPS/Register/register[15][5] ), .S0(
        n5590), .Y(\i_MIPS/Register/n633 ) );
  CLKMX2X2 U12309 ( .A(n5488), .B(\i_MIPS/Register/register[15][4] ), .S0(
        n5590), .Y(\i_MIPS/Register/n632 ) );
  CLKMX2X2 U12310 ( .A(n4776), .B(\i_MIPS/Register/register[15][3] ), .S0(
        n5590), .Y(\i_MIPS/Register/n631 ) );
  CLKMX2X2 U12311 ( .A(n5480), .B(\i_MIPS/Register/register[15][2] ), .S0(
        n5590), .Y(\i_MIPS/Register/n630 ) );
  CLKMX2X2 U12312 ( .A(n5477), .B(\i_MIPS/Register/register[15][1] ), .S0(
        n5591), .Y(\i_MIPS/Register/n629 ) );
  CLKMX2X2 U12313 ( .A(n5485), .B(\i_MIPS/Register/register[15][0] ), .S0(
        n5591), .Y(\i_MIPS/Register/n628 ) );
  CLKMX2X2 U12314 ( .A(n5470), .B(\i_MIPS/Register/register[16][31] ), .S0(
        n5588), .Y(\i_MIPS/Register/n627 ) );
  CLKMX2X2 U12315 ( .A(n5411), .B(\i_MIPS/Register/register[16][28] ), .S0(
        n5589), .Y(\i_MIPS/Register/n624 ) );
  CLKMX2X2 U12316 ( .A(n5408), .B(\i_MIPS/Register/register[16][27] ), .S0(
        n5588), .Y(\i_MIPS/Register/n623 ) );
  CLKMX2X2 U12317 ( .A(n5405), .B(\i_MIPS/Register/register[16][26] ), .S0(
        n5588), .Y(\i_MIPS/Register/n622 ) );
  CLKMX2X2 U12318 ( .A(n5414), .B(\i_MIPS/Register/register[16][25] ), .S0(
        n5589), .Y(\i_MIPS/Register/n621 ) );
  CLKMX2X2 U12319 ( .A(n5483), .B(\i_MIPS/Register/register[16][23] ), .S0(
        n5589), .Y(\i_MIPS/Register/n619 ) );
  CLKMX2X2 U12320 ( .A(n5423), .B(\i_MIPS/Register/register[16][22] ), .S0(
        n5588), .Y(\i_MIPS/Register/n618 ) );
  CLKMX2X2 U12321 ( .A(n5432), .B(\i_MIPS/Register/register[16][19] ), .S0(
        n5588), .Y(\i_MIPS/Register/n615 ) );
  CLKMX2X2 U12322 ( .A(n5417), .B(\i_MIPS/Register/register[16][18] ), .S0(
        n5589), .Y(\i_MIPS/Register/n614 ) );
  CLKMX2X2 U12323 ( .A(n5458), .B(\i_MIPS/Register/register[16][17] ), .S0(
        n5589), .Y(\i_MIPS/Register/n613 ) );
  CLKMX2X2 U12324 ( .A(n5456), .B(\i_MIPS/Register/register[16][15] ), .S0(
        n5589), .Y(\i_MIPS/Register/n611 ) );
  CLKMX2X2 U12325 ( .A(n5454), .B(\i_MIPS/Register/register[16][14] ), .S0(
        n5589), .Y(\i_MIPS/Register/n610 ) );
  CLKMX2X2 U12326 ( .A(n5452), .B(\i_MIPS/Register/register[16][13] ), .S0(
        n5589), .Y(\i_MIPS/Register/n609 ) );
  CLKMX2X2 U12327 ( .A(n5449), .B(\i_MIPS/Register/register[16][12] ), .S0(
        n5589), .Y(\i_MIPS/Register/n608 ) );
  CLKMX2X2 U12328 ( .A(n5446), .B(\i_MIPS/Register/register[16][11] ), .S0(
        n5588), .Y(\i_MIPS/Register/n607 ) );
  CLKMX2X2 U12329 ( .A(n5420), .B(\i_MIPS/Register/register[16][10] ), .S0(
        n5588), .Y(\i_MIPS/Register/n606 ) );
  CLKMX2X2 U12330 ( .A(n5475), .B(\i_MIPS/Register/register[16][8] ), .S0(
        n5589), .Y(\i_MIPS/Register/n604 ) );
  CLKMX2X2 U12331 ( .A(n5472), .B(\i_MIPS/Register/register[16][7] ), .S0(
        n5589), .Y(\i_MIPS/Register/n603 ) );
  CLKMX2X2 U12332 ( .A(n5043), .B(\i_MIPS/Register/register[16][6] ), .S0(
        n5588), .Y(\i_MIPS/Register/n602 ) );
  CLKMX2X2 U12333 ( .A(n5491), .B(\i_MIPS/Register/register[16][5] ), .S0(
        n5588), .Y(\i_MIPS/Register/n601 ) );
  CLKMX2X2 U12334 ( .A(n5488), .B(\i_MIPS/Register/register[16][4] ), .S0(
        n5588), .Y(\i_MIPS/Register/n600 ) );
  CLKMX2X2 U12335 ( .A(n4776), .B(\i_MIPS/Register/register[16][3] ), .S0(
        n5588), .Y(\i_MIPS/Register/n599 ) );
  CLKMX2X2 U12336 ( .A(n5480), .B(\i_MIPS/Register/register[16][2] ), .S0(
        n5588), .Y(\i_MIPS/Register/n598 ) );
  CLKMX2X2 U12337 ( .A(n5477), .B(\i_MIPS/Register/register[16][1] ), .S0(
        n5589), .Y(\i_MIPS/Register/n597 ) );
  CLKMX2X2 U12338 ( .A(n5485), .B(\i_MIPS/Register/register[16][0] ), .S0(
        n5589), .Y(\i_MIPS/Register/n596 ) );
  CLKMX2X2 U12339 ( .A(n5470), .B(\i_MIPS/Register/register[17][31] ), .S0(
        n5586), .Y(\i_MIPS/Register/n595 ) );
  CLKMX2X2 U12340 ( .A(n5411), .B(\i_MIPS/Register/register[17][28] ), .S0(
        n5587), .Y(\i_MIPS/Register/n592 ) );
  CLKMX2X2 U12341 ( .A(n5408), .B(\i_MIPS/Register/register[17][27] ), .S0(
        n5586), .Y(\i_MIPS/Register/n591 ) );
  CLKMX2X2 U12342 ( .A(n5405), .B(\i_MIPS/Register/register[17][26] ), .S0(
        n5586), .Y(\i_MIPS/Register/n590 ) );
  CLKMX2X2 U12343 ( .A(n5414), .B(\i_MIPS/Register/register[17][25] ), .S0(
        n5587), .Y(\i_MIPS/Register/n589 ) );
  CLKMX2X2 U12344 ( .A(n5483), .B(\i_MIPS/Register/register[17][23] ), .S0(
        n5587), .Y(\i_MIPS/Register/n587 ) );
  CLKMX2X2 U12345 ( .A(n5423), .B(\i_MIPS/Register/register[17][22] ), .S0(
        n5586), .Y(\i_MIPS/Register/n586 ) );
  CLKMX2X2 U12346 ( .A(n5432), .B(\i_MIPS/Register/register[17][19] ), .S0(
        n5586), .Y(\i_MIPS/Register/n583 ) );
  CLKMX2X2 U12347 ( .A(n5417), .B(\i_MIPS/Register/register[17][18] ), .S0(
        n5587), .Y(\i_MIPS/Register/n582 ) );
  CLKMX2X2 U12348 ( .A(n5458), .B(\i_MIPS/Register/register[17][17] ), .S0(
        n5587), .Y(\i_MIPS/Register/n581 ) );
  CLKMX2X2 U12349 ( .A(n5456), .B(\i_MIPS/Register/register[17][15] ), .S0(
        n5587), .Y(\i_MIPS/Register/n579 ) );
  CLKMX2X2 U12350 ( .A(n5454), .B(\i_MIPS/Register/register[17][14] ), .S0(
        n5587), .Y(\i_MIPS/Register/n578 ) );
  CLKMX2X2 U12351 ( .A(n5452), .B(\i_MIPS/Register/register[17][13] ), .S0(
        n5587), .Y(\i_MIPS/Register/n577 ) );
  CLKMX2X2 U12352 ( .A(n5449), .B(\i_MIPS/Register/register[17][12] ), .S0(
        n5587), .Y(\i_MIPS/Register/n576 ) );
  CLKMX2X2 U12353 ( .A(n5446), .B(\i_MIPS/Register/register[17][11] ), .S0(
        n5586), .Y(\i_MIPS/Register/n575 ) );
  CLKMX2X2 U12354 ( .A(n5420), .B(\i_MIPS/Register/register[17][10] ), .S0(
        n5586), .Y(\i_MIPS/Register/n574 ) );
  CLKMX2X2 U12355 ( .A(n5475), .B(\i_MIPS/Register/register[17][8] ), .S0(
        n5587), .Y(\i_MIPS/Register/n572 ) );
  CLKMX2X2 U12356 ( .A(n5472), .B(\i_MIPS/Register/register[17][7] ), .S0(
        n5587), .Y(\i_MIPS/Register/n571 ) );
  CLKMX2X2 U12357 ( .A(n5043), .B(\i_MIPS/Register/register[17][6] ), .S0(
        n5586), .Y(\i_MIPS/Register/n570 ) );
  CLKMX2X2 U12358 ( .A(n5491), .B(\i_MIPS/Register/register[17][5] ), .S0(
        n5586), .Y(\i_MIPS/Register/n569 ) );
  CLKMX2X2 U12359 ( .A(n5488), .B(\i_MIPS/Register/register[17][4] ), .S0(
        n5586), .Y(\i_MIPS/Register/n568 ) );
  CLKMX2X2 U12360 ( .A(n4776), .B(\i_MIPS/Register/register[17][3] ), .S0(
        n5586), .Y(\i_MIPS/Register/n567 ) );
  CLKMX2X2 U12361 ( .A(n5480), .B(\i_MIPS/Register/register[17][2] ), .S0(
        n5586), .Y(\i_MIPS/Register/n566 ) );
  CLKMX2X2 U12362 ( .A(n5477), .B(\i_MIPS/Register/register[17][1] ), .S0(
        n5587), .Y(\i_MIPS/Register/n565 ) );
  CLKMX2X2 U12363 ( .A(n5485), .B(\i_MIPS/Register/register[17][0] ), .S0(
        n5587), .Y(\i_MIPS/Register/n564 ) );
  CLKMX2X2 U12364 ( .A(n5470), .B(\i_MIPS/Register/register[18][31] ), .S0(
        n5584), .Y(\i_MIPS/Register/n563 ) );
  CLKMX2X2 U12365 ( .A(n5411), .B(\i_MIPS/Register/register[18][28] ), .S0(
        n5585), .Y(\i_MIPS/Register/n560 ) );
  CLKMX2X2 U12366 ( .A(n5408), .B(\i_MIPS/Register/register[18][27] ), .S0(
        n5584), .Y(\i_MIPS/Register/n559 ) );
  CLKMX2X2 U12367 ( .A(n5405), .B(\i_MIPS/Register/register[18][26] ), .S0(
        n5584), .Y(\i_MIPS/Register/n558 ) );
  CLKMX2X2 U12368 ( .A(n5414), .B(\i_MIPS/Register/register[18][25] ), .S0(
        n5585), .Y(\i_MIPS/Register/n557 ) );
  CLKMX2X2 U12369 ( .A(n5483), .B(\i_MIPS/Register/register[18][23] ), .S0(
        n5585), .Y(\i_MIPS/Register/n555 ) );
  CLKMX2X2 U12370 ( .A(n5423), .B(\i_MIPS/Register/register[18][22] ), .S0(
        n5584), .Y(\i_MIPS/Register/n554 ) );
  CLKMX2X2 U12371 ( .A(n5432), .B(\i_MIPS/Register/register[18][19] ), .S0(
        n5584), .Y(\i_MIPS/Register/n551 ) );
  CLKMX2X2 U12372 ( .A(n5417), .B(\i_MIPS/Register/register[18][18] ), .S0(
        n5585), .Y(\i_MIPS/Register/n550 ) );
  CLKMX2X2 U12373 ( .A(n5458), .B(\i_MIPS/Register/register[18][17] ), .S0(
        n5585), .Y(\i_MIPS/Register/n549 ) );
  CLKMX2X2 U12374 ( .A(n5456), .B(\i_MIPS/Register/register[18][15] ), .S0(
        n5585), .Y(\i_MIPS/Register/n547 ) );
  CLKMX2X2 U12375 ( .A(n5454), .B(\i_MIPS/Register/register[18][14] ), .S0(
        n5585), .Y(\i_MIPS/Register/n546 ) );
  CLKMX2X2 U12376 ( .A(n5452), .B(\i_MIPS/Register/register[18][13] ), .S0(
        n5585), .Y(\i_MIPS/Register/n545 ) );
  CLKMX2X2 U12377 ( .A(n5449), .B(\i_MIPS/Register/register[18][12] ), .S0(
        n5585), .Y(\i_MIPS/Register/n544 ) );
  CLKMX2X2 U12378 ( .A(n5446), .B(\i_MIPS/Register/register[18][11] ), .S0(
        n5584), .Y(\i_MIPS/Register/n543 ) );
  CLKMX2X2 U12379 ( .A(n5420), .B(\i_MIPS/Register/register[18][10] ), .S0(
        n5584), .Y(\i_MIPS/Register/n542 ) );
  CLKMX2X2 U12380 ( .A(n5475), .B(\i_MIPS/Register/register[18][8] ), .S0(
        n5585), .Y(\i_MIPS/Register/n540 ) );
  CLKMX2X2 U12381 ( .A(n5472), .B(\i_MIPS/Register/register[18][7] ), .S0(
        n5585), .Y(\i_MIPS/Register/n539 ) );
  CLKMX2X2 U12382 ( .A(n5043), .B(\i_MIPS/Register/register[18][6] ), .S0(
        n5584), .Y(\i_MIPS/Register/n538 ) );
  CLKMX2X2 U12383 ( .A(n5491), .B(\i_MIPS/Register/register[18][5] ), .S0(
        n5584), .Y(\i_MIPS/Register/n537 ) );
  CLKMX2X2 U12384 ( .A(n5488), .B(\i_MIPS/Register/register[18][4] ), .S0(
        n5584), .Y(\i_MIPS/Register/n536 ) );
  CLKMX2X2 U12385 ( .A(n4776), .B(\i_MIPS/Register/register[18][3] ), .S0(
        n5584), .Y(\i_MIPS/Register/n535 ) );
  CLKMX2X2 U12386 ( .A(n5480), .B(\i_MIPS/Register/register[18][2] ), .S0(
        n5584), .Y(\i_MIPS/Register/n534 ) );
  CLKMX2X2 U12387 ( .A(n5477), .B(\i_MIPS/Register/register[18][1] ), .S0(
        n5585), .Y(\i_MIPS/Register/n533 ) );
  CLKMX2X2 U12388 ( .A(n5485), .B(\i_MIPS/Register/register[18][0] ), .S0(
        n5585), .Y(\i_MIPS/Register/n532 ) );
  CLKMX2X2 U12389 ( .A(n5470), .B(\i_MIPS/Register/register[19][31] ), .S0(
        n5582), .Y(\i_MIPS/Register/n531 ) );
  CLKMX2X2 U12390 ( .A(n5410), .B(\i_MIPS/Register/register[19][28] ), .S0(
        n5583), .Y(\i_MIPS/Register/n528 ) );
  CLKMX2X2 U12391 ( .A(n5407), .B(\i_MIPS/Register/register[19][27] ), .S0(
        n5582), .Y(\i_MIPS/Register/n527 ) );
  CLKMX2X2 U12392 ( .A(n5405), .B(\i_MIPS/Register/register[19][26] ), .S0(
        n5582), .Y(\i_MIPS/Register/n526 ) );
  CLKMX2X2 U12393 ( .A(n5413), .B(\i_MIPS/Register/register[19][25] ), .S0(
        n5583), .Y(\i_MIPS/Register/n525 ) );
  CLKMX2X2 U12394 ( .A(n5483), .B(\i_MIPS/Register/register[19][23] ), .S0(
        n5583), .Y(\i_MIPS/Register/n523 ) );
  CLKMX2X2 U12395 ( .A(n5423), .B(\i_MIPS/Register/register[19][22] ), .S0(
        n5582), .Y(\i_MIPS/Register/n522 ) );
  CLKMX2X2 U12396 ( .A(n5431), .B(\i_MIPS/Register/register[19][19] ), .S0(
        n5582), .Y(\i_MIPS/Register/n519 ) );
  CLKMX2X2 U12397 ( .A(n5417), .B(\i_MIPS/Register/register[19][18] ), .S0(
        n5583), .Y(\i_MIPS/Register/n518 ) );
  CLKMX2X2 U12398 ( .A(n5458), .B(\i_MIPS/Register/register[19][17] ), .S0(
        n5583), .Y(\i_MIPS/Register/n517 ) );
  CLKMX2X2 U12399 ( .A(n5456), .B(\i_MIPS/Register/register[19][15] ), .S0(
        n5583), .Y(\i_MIPS/Register/n515 ) );
  CLKMX2X2 U12400 ( .A(n5454), .B(\i_MIPS/Register/register[19][14] ), .S0(
        n5583), .Y(\i_MIPS/Register/n514 ) );
  CLKMX2X2 U12401 ( .A(n5452), .B(\i_MIPS/Register/register[19][13] ), .S0(
        n5583), .Y(\i_MIPS/Register/n513 ) );
  CLKMX2X2 U12402 ( .A(n5448), .B(\i_MIPS/Register/register[19][12] ), .S0(
        n5583), .Y(\i_MIPS/Register/n512 ) );
  CLKMX2X2 U12403 ( .A(n5446), .B(\i_MIPS/Register/register[19][11] ), .S0(
        n5582), .Y(\i_MIPS/Register/n511 ) );
  CLKMX2X2 U12404 ( .A(n5420), .B(\i_MIPS/Register/register[19][10] ), .S0(
        n5582), .Y(\i_MIPS/Register/n510 ) );
  CLKMX2X2 U12405 ( .A(n5475), .B(\i_MIPS/Register/register[19][8] ), .S0(
        n5583), .Y(\i_MIPS/Register/n508 ) );
  CLKMX2X2 U12406 ( .A(n5472), .B(\i_MIPS/Register/register[19][7] ), .S0(
        n5583), .Y(\i_MIPS/Register/n507 ) );
  CLKMX2X2 U12407 ( .A(n5043), .B(\i_MIPS/Register/register[19][6] ), .S0(
        n5582), .Y(\i_MIPS/Register/n506 ) );
  CLKMX2X2 U12408 ( .A(n5490), .B(\i_MIPS/Register/register[19][5] ), .S0(
        n5582), .Y(\i_MIPS/Register/n505 ) );
  CLKMX2X2 U12409 ( .A(n5488), .B(\i_MIPS/Register/register[19][4] ), .S0(
        n5582), .Y(\i_MIPS/Register/n504 ) );
  CLKMX2X2 U12410 ( .A(n4775), .B(\i_MIPS/Register/register[19][3] ), .S0(
        n5582), .Y(\i_MIPS/Register/n503 ) );
  CLKMX2X2 U12411 ( .A(n5480), .B(\i_MIPS/Register/register[19][2] ), .S0(
        n5582), .Y(\i_MIPS/Register/n502 ) );
  CLKMX2X2 U12412 ( .A(n5477), .B(\i_MIPS/Register/register[19][1] ), .S0(
        n5583), .Y(\i_MIPS/Register/n501 ) );
  CLKMX2X2 U12413 ( .A(n5484), .B(\i_MIPS/Register/register[19][0] ), .S0(
        n5583), .Y(\i_MIPS/Register/n500 ) );
  CLKMX2X2 U12414 ( .A(n5470), .B(\i_MIPS/Register/register[20][31] ), .S0(
        n5580), .Y(\i_MIPS/Register/n499 ) );
  CLKMX2X2 U12415 ( .A(n5411), .B(\i_MIPS/Register/register[20][28] ), .S0(
        n5581), .Y(\i_MIPS/Register/n496 ) );
  CLKMX2X2 U12416 ( .A(n5408), .B(\i_MIPS/Register/register[20][27] ), .S0(
        n5580), .Y(\i_MIPS/Register/n495 ) );
  CLKMX2X2 U12417 ( .A(n5405), .B(\i_MIPS/Register/register[20][26] ), .S0(
        n5580), .Y(\i_MIPS/Register/n494 ) );
  CLKMX2X2 U12418 ( .A(n5414), .B(\i_MIPS/Register/register[20][25] ), .S0(
        n5581), .Y(\i_MIPS/Register/n493 ) );
  CLKMX2X2 U12419 ( .A(n5483), .B(\i_MIPS/Register/register[20][23] ), .S0(
        n5581), .Y(\i_MIPS/Register/n491 ) );
  CLKMX2X2 U12420 ( .A(n5423), .B(\i_MIPS/Register/register[20][22] ), .S0(
        n5580), .Y(\i_MIPS/Register/n490 ) );
  CLKMX2X2 U12421 ( .A(n5432), .B(\i_MIPS/Register/register[20][19] ), .S0(
        n5580), .Y(\i_MIPS/Register/n487 ) );
  CLKMX2X2 U12422 ( .A(n5417), .B(\i_MIPS/Register/register[20][18] ), .S0(
        n5581), .Y(\i_MIPS/Register/n486 ) );
  CLKMX2X2 U12423 ( .A(n5458), .B(\i_MIPS/Register/register[20][17] ), .S0(
        n5581), .Y(\i_MIPS/Register/n485 ) );
  CLKMX2X2 U12424 ( .A(n5456), .B(\i_MIPS/Register/register[20][15] ), .S0(
        n5581), .Y(\i_MIPS/Register/n483 ) );
  CLKMX2X2 U12425 ( .A(n5454), .B(\i_MIPS/Register/register[20][14] ), .S0(
        n5581), .Y(\i_MIPS/Register/n482 ) );
  CLKMX2X2 U12426 ( .A(n5452), .B(\i_MIPS/Register/register[20][13] ), .S0(
        n5581), .Y(\i_MIPS/Register/n481 ) );
  CLKMX2X2 U12427 ( .A(n5449), .B(\i_MIPS/Register/register[20][12] ), .S0(
        n5581), .Y(\i_MIPS/Register/n480 ) );
  CLKMX2X2 U12428 ( .A(n5446), .B(\i_MIPS/Register/register[20][11] ), .S0(
        n5580), .Y(\i_MIPS/Register/n479 ) );
  CLKMX2X2 U12429 ( .A(n5420), .B(\i_MIPS/Register/register[20][10] ), .S0(
        n5580), .Y(\i_MIPS/Register/n478 ) );
  CLKMX2X2 U12430 ( .A(n5475), .B(\i_MIPS/Register/register[20][8] ), .S0(
        n5581), .Y(\i_MIPS/Register/n476 ) );
  CLKMX2X2 U12431 ( .A(n5472), .B(\i_MIPS/Register/register[20][7] ), .S0(
        n5581), .Y(\i_MIPS/Register/n475 ) );
  CLKMX2X2 U12432 ( .A(n5043), .B(\i_MIPS/Register/register[20][6] ), .S0(
        n5580), .Y(\i_MIPS/Register/n474 ) );
  CLKMX2X2 U12433 ( .A(n5491), .B(\i_MIPS/Register/register[20][5] ), .S0(
        n5580), .Y(\i_MIPS/Register/n473 ) );
  CLKMX2X2 U12434 ( .A(n5488), .B(\i_MIPS/Register/register[20][4] ), .S0(
        n5580), .Y(\i_MIPS/Register/n472 ) );
  CLKMX2X2 U12435 ( .A(n4776), .B(\i_MIPS/Register/register[20][3] ), .S0(
        n5580), .Y(\i_MIPS/Register/n471 ) );
  CLKMX2X2 U12436 ( .A(n5480), .B(\i_MIPS/Register/register[20][2] ), .S0(
        n5580), .Y(\i_MIPS/Register/n470 ) );
  CLKMX2X2 U12437 ( .A(n5477), .B(\i_MIPS/Register/register[20][1] ), .S0(
        n5581), .Y(\i_MIPS/Register/n469 ) );
  CLKMX2X2 U12438 ( .A(n5485), .B(\i_MIPS/Register/register[20][0] ), .S0(
        n5581), .Y(\i_MIPS/Register/n468 ) );
  CLKMX2X2 U12439 ( .A(n5470), .B(\i_MIPS/Register/register[21][31] ), .S0(
        n5578), .Y(\i_MIPS/Register/n467 ) );
  CLKMX2X2 U12440 ( .A(n5411), .B(\i_MIPS/Register/register[21][28] ), .S0(
        n5579), .Y(\i_MIPS/Register/n464 ) );
  CLKMX2X2 U12441 ( .A(n5408), .B(\i_MIPS/Register/register[21][27] ), .S0(
        n5578), .Y(\i_MIPS/Register/n463 ) );
  CLKMX2X2 U12442 ( .A(n5405), .B(\i_MIPS/Register/register[21][26] ), .S0(
        n5578), .Y(\i_MIPS/Register/n462 ) );
  CLKMX2X2 U12443 ( .A(n5414), .B(\i_MIPS/Register/register[21][25] ), .S0(
        n5579), .Y(\i_MIPS/Register/n461 ) );
  CLKMX2X2 U12444 ( .A(n5483), .B(\i_MIPS/Register/register[21][23] ), .S0(
        n5579), .Y(\i_MIPS/Register/n459 ) );
  CLKMX2X2 U12445 ( .A(n5423), .B(\i_MIPS/Register/register[21][22] ), .S0(
        n5578), .Y(\i_MIPS/Register/n458 ) );
  CLKMX2X2 U12446 ( .A(n5432), .B(\i_MIPS/Register/register[21][19] ), .S0(
        n5578), .Y(\i_MIPS/Register/n455 ) );
  CLKMX2X2 U12447 ( .A(n5416), .B(\i_MIPS/Register/register[21][18] ), .S0(
        n5579), .Y(\i_MIPS/Register/n454 ) );
  CLKMX2X2 U12448 ( .A(n5458), .B(\i_MIPS/Register/register[21][17] ), .S0(
        n5579), .Y(\i_MIPS/Register/n453 ) );
  CLKMX2X2 U12449 ( .A(n5456), .B(\i_MIPS/Register/register[21][15] ), .S0(
        n5579), .Y(\i_MIPS/Register/n451 ) );
  CLKMX2X2 U12450 ( .A(n5454), .B(\i_MIPS/Register/register[21][14] ), .S0(
        n5579), .Y(\i_MIPS/Register/n450 ) );
  CLKMX2X2 U12451 ( .A(n5452), .B(\i_MIPS/Register/register[21][13] ), .S0(
        n5579), .Y(\i_MIPS/Register/n449 ) );
  CLKMX2X2 U12452 ( .A(n5449), .B(\i_MIPS/Register/register[21][12] ), .S0(
        n5579), .Y(\i_MIPS/Register/n448 ) );
  CLKMX2X2 U12453 ( .A(n5446), .B(\i_MIPS/Register/register[21][11] ), .S0(
        n5578), .Y(\i_MIPS/Register/n447 ) );
  CLKMX2X2 U12454 ( .A(n5420), .B(\i_MIPS/Register/register[21][10] ), .S0(
        n5578), .Y(\i_MIPS/Register/n446 ) );
  CLKMX2X2 U12455 ( .A(n5475), .B(\i_MIPS/Register/register[21][8] ), .S0(
        n5579), .Y(\i_MIPS/Register/n444 ) );
  CLKMX2X2 U12456 ( .A(n5472), .B(\i_MIPS/Register/register[21][7] ), .S0(
        n5579), .Y(\i_MIPS/Register/n443 ) );
  CLKMX2X2 U12457 ( .A(n5043), .B(\i_MIPS/Register/register[21][6] ), .S0(
        n5578), .Y(\i_MIPS/Register/n442 ) );
  CLKMX2X2 U12458 ( .A(n5491), .B(\i_MIPS/Register/register[21][5] ), .S0(
        n5578), .Y(\i_MIPS/Register/n441 ) );
  CLKMX2X2 U12459 ( .A(n5488), .B(\i_MIPS/Register/register[21][4] ), .S0(
        n5578), .Y(\i_MIPS/Register/n440 ) );
  CLKMX2X2 U12460 ( .A(n4776), .B(\i_MIPS/Register/register[21][3] ), .S0(
        n5578), .Y(\i_MIPS/Register/n439 ) );
  CLKMX2X2 U12461 ( .A(n5480), .B(\i_MIPS/Register/register[21][2] ), .S0(
        n5578), .Y(\i_MIPS/Register/n438 ) );
  CLKMX2X2 U12462 ( .A(n5477), .B(\i_MIPS/Register/register[21][1] ), .S0(
        n5579), .Y(\i_MIPS/Register/n437 ) );
  CLKMX2X2 U12463 ( .A(n5485), .B(\i_MIPS/Register/register[21][0] ), .S0(
        n5579), .Y(\i_MIPS/Register/n436 ) );
  CLKMX2X2 U12464 ( .A(n5470), .B(\i_MIPS/Register/register[22][31] ), .S0(
        n5576), .Y(\i_MIPS/Register/n435 ) );
  CLKMX2X2 U12465 ( .A(n5411), .B(\i_MIPS/Register/register[22][28] ), .S0(
        n5577), .Y(\i_MIPS/Register/n432 ) );
  CLKMX2X2 U12466 ( .A(n5408), .B(\i_MIPS/Register/register[22][27] ), .S0(
        n5576), .Y(\i_MIPS/Register/n431 ) );
  CLKMX2X2 U12467 ( .A(n5405), .B(\i_MIPS/Register/register[22][26] ), .S0(
        n5576), .Y(\i_MIPS/Register/n430 ) );
  CLKMX2X2 U12468 ( .A(n5414), .B(\i_MIPS/Register/register[22][25] ), .S0(
        n5577), .Y(\i_MIPS/Register/n429 ) );
  CLKMX2X2 U12469 ( .A(n5483), .B(\i_MIPS/Register/register[22][23] ), .S0(
        n5577), .Y(\i_MIPS/Register/n427 ) );
  CLKMX2X2 U12470 ( .A(n5423), .B(\i_MIPS/Register/register[22][22] ), .S0(
        n5576), .Y(\i_MIPS/Register/n426 ) );
  CLKMX2X2 U12471 ( .A(n5432), .B(\i_MIPS/Register/register[22][19] ), .S0(
        n5576), .Y(\i_MIPS/Register/n423 ) );
  CLKMX2X2 U12472 ( .A(n5417), .B(\i_MIPS/Register/register[22][18] ), .S0(
        n5577), .Y(\i_MIPS/Register/n422 ) );
  CLKMX2X2 U12473 ( .A(n5458), .B(\i_MIPS/Register/register[22][17] ), .S0(
        n5577), .Y(\i_MIPS/Register/n421 ) );
  CLKMX2X2 U12474 ( .A(n5456), .B(\i_MIPS/Register/register[22][15] ), .S0(
        n5577), .Y(\i_MIPS/Register/n419 ) );
  CLKMX2X2 U12475 ( .A(n5454), .B(\i_MIPS/Register/register[22][14] ), .S0(
        n5577), .Y(\i_MIPS/Register/n418 ) );
  CLKMX2X2 U12476 ( .A(n5452), .B(\i_MIPS/Register/register[22][13] ), .S0(
        n5577), .Y(\i_MIPS/Register/n417 ) );
  CLKMX2X2 U12477 ( .A(n5449), .B(\i_MIPS/Register/register[22][12] ), .S0(
        n5577), .Y(\i_MIPS/Register/n416 ) );
  CLKMX2X2 U12478 ( .A(n5446), .B(\i_MIPS/Register/register[22][11] ), .S0(
        n5576), .Y(\i_MIPS/Register/n415 ) );
  CLKMX2X2 U12479 ( .A(n5420), .B(\i_MIPS/Register/register[22][10] ), .S0(
        n5576), .Y(\i_MIPS/Register/n414 ) );
  CLKMX2X2 U12480 ( .A(n5475), .B(\i_MIPS/Register/register[22][8] ), .S0(
        n5577), .Y(\i_MIPS/Register/n412 ) );
  CLKMX2X2 U12481 ( .A(n5472), .B(\i_MIPS/Register/register[22][7] ), .S0(
        n5577), .Y(\i_MIPS/Register/n411 ) );
  CLKMX2X2 U12482 ( .A(n5042), .B(\i_MIPS/Register/register[22][6] ), .S0(
        n5576), .Y(\i_MIPS/Register/n410 ) );
  CLKMX2X2 U12483 ( .A(n5491), .B(\i_MIPS/Register/register[22][5] ), .S0(
        n5576), .Y(\i_MIPS/Register/n409 ) );
  CLKMX2X2 U12484 ( .A(n5488), .B(\i_MIPS/Register/register[22][4] ), .S0(
        n5576), .Y(\i_MIPS/Register/n408 ) );
  CLKMX2X2 U12485 ( .A(n4776), .B(\i_MIPS/Register/register[22][3] ), .S0(
        n5576), .Y(\i_MIPS/Register/n407 ) );
  CLKMX2X2 U12486 ( .A(n5480), .B(\i_MIPS/Register/register[22][2] ), .S0(
        n5576), .Y(\i_MIPS/Register/n406 ) );
  CLKMX2X2 U12487 ( .A(n5477), .B(\i_MIPS/Register/register[22][1] ), .S0(
        n5577), .Y(\i_MIPS/Register/n405 ) );
  CLKMX2X2 U12488 ( .A(n5485), .B(\i_MIPS/Register/register[22][0] ), .S0(
        n5577), .Y(\i_MIPS/Register/n404 ) );
  CLKMX2X2 U12489 ( .A(n5469), .B(\i_MIPS/Register/register[23][31] ), .S0(
        n5574), .Y(\i_MIPS/Register/n403 ) );
  CLKMX2X2 U12490 ( .A(n5410), .B(\i_MIPS/Register/register[23][28] ), .S0(
        n5575), .Y(\i_MIPS/Register/n400 ) );
  CLKMX2X2 U12491 ( .A(n5407), .B(\i_MIPS/Register/register[23][27] ), .S0(
        n5574), .Y(\i_MIPS/Register/n399 ) );
  CLKMX2X2 U12492 ( .A(n5404), .B(\i_MIPS/Register/register[23][26] ), .S0(
        n5574), .Y(\i_MIPS/Register/n398 ) );
  CLKMX2X2 U12493 ( .A(n5413), .B(\i_MIPS/Register/register[23][25] ), .S0(
        n5575), .Y(\i_MIPS/Register/n397 ) );
  CLKMX2X2 U12494 ( .A(n5482), .B(\i_MIPS/Register/register[23][23] ), .S0(
        n5575), .Y(\i_MIPS/Register/n395 ) );
  CLKMX2X2 U12495 ( .A(n5422), .B(\i_MIPS/Register/register[23][22] ), .S0(
        n5574), .Y(\i_MIPS/Register/n394 ) );
  CLKMX2X2 U12496 ( .A(n5431), .B(\i_MIPS/Register/register[23][19] ), .S0(
        n5574), .Y(\i_MIPS/Register/n391 ) );
  CLKMX2X2 U12497 ( .A(n5417), .B(\i_MIPS/Register/register[23][18] ), .S0(
        n5575), .Y(\i_MIPS/Register/n390 ) );
  CLKMX2X2 U12498 ( .A(n5457), .B(\i_MIPS/Register/register[23][17] ), .S0(
        n5575), .Y(\i_MIPS/Register/n389 ) );
  CLKMX2X2 U12499 ( .A(n5455), .B(\i_MIPS/Register/register[23][15] ), .S0(
        n5575), .Y(\i_MIPS/Register/n387 ) );
  CLKMX2X2 U12500 ( .A(n5453), .B(\i_MIPS/Register/register[23][14] ), .S0(
        n5575), .Y(\i_MIPS/Register/n386 ) );
  CLKMX2X2 U12501 ( .A(n5451), .B(\i_MIPS/Register/register[23][13] ), .S0(
        n5575), .Y(\i_MIPS/Register/n385 ) );
  CLKMX2X2 U12502 ( .A(n5449), .B(\i_MIPS/Register/register[23][12] ), .S0(
        n5575), .Y(\i_MIPS/Register/n384 ) );
  CLKMX2X2 U12503 ( .A(n5445), .B(\i_MIPS/Register/register[23][11] ), .S0(
        n5574), .Y(\i_MIPS/Register/n383 ) );
  CLKMX2X2 U12504 ( .A(n5419), .B(\i_MIPS/Register/register[23][10] ), .S0(
        n5574), .Y(\i_MIPS/Register/n382 ) );
  CLKMX2X2 U12505 ( .A(n5474), .B(\i_MIPS/Register/register[23][8] ), .S0(
        n5575), .Y(\i_MIPS/Register/n380 ) );
  CLKMX2X2 U12506 ( .A(n5471), .B(\i_MIPS/Register/register[23][7] ), .S0(
        n5575), .Y(\i_MIPS/Register/n379 ) );
  CLKMX2X2 U12507 ( .A(n5043), .B(\i_MIPS/Register/register[23][6] ), .S0(
        n5574), .Y(\i_MIPS/Register/n378 ) );
  CLKMX2X2 U12508 ( .A(n5491), .B(\i_MIPS/Register/register[23][5] ), .S0(
        n5574), .Y(\i_MIPS/Register/n377 ) );
  CLKMX2X2 U12509 ( .A(n5487), .B(\i_MIPS/Register/register[23][4] ), .S0(
        n5574), .Y(\i_MIPS/Register/n376 ) );
  CLKMX2X2 U12510 ( .A(n4775), .B(\i_MIPS/Register/register[23][3] ), .S0(
        n5574), .Y(\i_MIPS/Register/n375 ) );
  CLKMX2X2 U12511 ( .A(n5479), .B(\i_MIPS/Register/register[23][2] ), .S0(
        n5574), .Y(\i_MIPS/Register/n374 ) );
  CLKMX2X2 U12512 ( .A(n5476), .B(\i_MIPS/Register/register[23][1] ), .S0(
        n5575), .Y(\i_MIPS/Register/n373 ) );
  CLKMX2X2 U12513 ( .A(n5485), .B(\i_MIPS/Register/register[23][0] ), .S0(
        n5575), .Y(\i_MIPS/Register/n372 ) );
  CLKMX2X2 U12514 ( .A(n5470), .B(\i_MIPS/Register/register[24][31] ), .S0(
        n5572), .Y(\i_MIPS/Register/n371 ) );
  CLKMX2X2 U12515 ( .A(n5411), .B(\i_MIPS/Register/register[24][28] ), .S0(
        n5573), .Y(\i_MIPS/Register/n368 ) );
  CLKMX2X2 U12516 ( .A(n5408), .B(\i_MIPS/Register/register[24][27] ), .S0(
        n5572), .Y(\i_MIPS/Register/n367 ) );
  CLKMX2X2 U12517 ( .A(n5405), .B(\i_MIPS/Register/register[24][26] ), .S0(
        n5572), .Y(\i_MIPS/Register/n366 ) );
  CLKMX2X2 U12518 ( .A(n5414), .B(\i_MIPS/Register/register[24][25] ), .S0(
        n5573), .Y(\i_MIPS/Register/n365 ) );
  CLKMX2X2 U12519 ( .A(n5483), .B(\i_MIPS/Register/register[24][23] ), .S0(
        n5573), .Y(\i_MIPS/Register/n363 ) );
  CLKMX2X2 U12520 ( .A(n5423), .B(\i_MIPS/Register/register[24][22] ), .S0(
        n5572), .Y(\i_MIPS/Register/n362 ) );
  CLKMX2X2 U12521 ( .A(n5432), .B(\i_MIPS/Register/register[24][19] ), .S0(
        n5572), .Y(\i_MIPS/Register/n359 ) );
  CLKMX2X2 U12522 ( .A(n5417), .B(\i_MIPS/Register/register[24][18] ), .S0(
        n5573), .Y(\i_MIPS/Register/n358 ) );
  CLKMX2X2 U12523 ( .A(n5458), .B(\i_MIPS/Register/register[24][17] ), .S0(
        n5573), .Y(\i_MIPS/Register/n357 ) );
  CLKMX2X2 U12524 ( .A(n5456), .B(\i_MIPS/Register/register[24][15] ), .S0(
        n5573), .Y(\i_MIPS/Register/n355 ) );
  CLKMX2X2 U12525 ( .A(n5454), .B(\i_MIPS/Register/register[24][14] ), .S0(
        n5573), .Y(\i_MIPS/Register/n354 ) );
  CLKMX2X2 U12526 ( .A(n5452), .B(\i_MIPS/Register/register[24][13] ), .S0(
        n5573), .Y(\i_MIPS/Register/n353 ) );
  CLKMX2X2 U12527 ( .A(n5449), .B(\i_MIPS/Register/register[24][12] ), .S0(
        n5573), .Y(\i_MIPS/Register/n352 ) );
  CLKMX2X2 U12528 ( .A(n5446), .B(\i_MIPS/Register/register[24][11] ), .S0(
        n5572), .Y(\i_MIPS/Register/n351 ) );
  CLKMX2X2 U12529 ( .A(n5420), .B(\i_MIPS/Register/register[24][10] ), .S0(
        n5572), .Y(\i_MIPS/Register/n350 ) );
  CLKMX2X2 U12530 ( .A(n5475), .B(\i_MIPS/Register/register[24][8] ), .S0(
        n5573), .Y(\i_MIPS/Register/n348 ) );
  CLKMX2X2 U12531 ( .A(n5472), .B(\i_MIPS/Register/register[24][7] ), .S0(
        n5573), .Y(\i_MIPS/Register/n347 ) );
  CLKMX2X2 U12532 ( .A(n5043), .B(\i_MIPS/Register/register[24][6] ), .S0(
        n5572), .Y(\i_MIPS/Register/n346 ) );
  CLKMX2X2 U12533 ( .A(n5491), .B(\i_MIPS/Register/register[24][5] ), .S0(
        n5572), .Y(\i_MIPS/Register/n345 ) );
  CLKMX2X2 U12534 ( .A(n5488), .B(\i_MIPS/Register/register[24][4] ), .S0(
        n5572), .Y(\i_MIPS/Register/n344 ) );
  CLKMX2X2 U12535 ( .A(n4776), .B(\i_MIPS/Register/register[24][3] ), .S0(
        n5572), .Y(\i_MIPS/Register/n343 ) );
  CLKMX2X2 U12536 ( .A(n5480), .B(\i_MIPS/Register/register[24][2] ), .S0(
        n5572), .Y(\i_MIPS/Register/n342 ) );
  CLKMX2X2 U12537 ( .A(n5477), .B(\i_MIPS/Register/register[24][1] ), .S0(
        n5573), .Y(\i_MIPS/Register/n341 ) );
  CLKMX2X2 U12538 ( .A(n5485), .B(\i_MIPS/Register/register[24][0] ), .S0(
        n5573), .Y(\i_MIPS/Register/n340 ) );
  CLKMX2X2 U12539 ( .A(n5470), .B(\i_MIPS/Register/register[25][31] ), .S0(
        n5570), .Y(\i_MIPS/Register/n339 ) );
  CLKMX2X2 U12540 ( .A(n5411), .B(\i_MIPS/Register/register[25][28] ), .S0(
        n5571), .Y(\i_MIPS/Register/n336 ) );
  CLKMX2X2 U12541 ( .A(n5408), .B(\i_MIPS/Register/register[25][27] ), .S0(
        n5570), .Y(\i_MIPS/Register/n335 ) );
  CLKMX2X2 U12542 ( .A(n5405), .B(\i_MIPS/Register/register[25][26] ), .S0(
        n5570), .Y(\i_MIPS/Register/n334 ) );
  CLKMX2X2 U12543 ( .A(n5414), .B(\i_MIPS/Register/register[25][25] ), .S0(
        n5571), .Y(\i_MIPS/Register/n333 ) );
  CLKMX2X2 U12544 ( .A(n5483), .B(\i_MIPS/Register/register[25][23] ), .S0(
        n5571), .Y(\i_MIPS/Register/n331 ) );
  CLKMX2X2 U12545 ( .A(n5423), .B(\i_MIPS/Register/register[25][22] ), .S0(
        n5570), .Y(\i_MIPS/Register/n330 ) );
  CLKMX2X2 U12546 ( .A(n5432), .B(\i_MIPS/Register/register[25][19] ), .S0(
        n5570), .Y(\i_MIPS/Register/n327 ) );
  CLKMX2X2 U12547 ( .A(n5417), .B(\i_MIPS/Register/register[25][18] ), .S0(
        n5571), .Y(\i_MIPS/Register/n326 ) );
  CLKMX2X2 U12548 ( .A(n5458), .B(\i_MIPS/Register/register[25][17] ), .S0(
        n5571), .Y(\i_MIPS/Register/n325 ) );
  CLKMX2X2 U12549 ( .A(n5456), .B(\i_MIPS/Register/register[25][15] ), .S0(
        n5571), .Y(\i_MIPS/Register/n323 ) );
  CLKMX2X2 U12550 ( .A(n5454), .B(\i_MIPS/Register/register[25][14] ), .S0(
        n5571), .Y(\i_MIPS/Register/n322 ) );
  CLKMX2X2 U12551 ( .A(n5452), .B(\i_MIPS/Register/register[25][13] ), .S0(
        n5571), .Y(\i_MIPS/Register/n321 ) );
  CLKMX2X2 U12552 ( .A(n5449), .B(\i_MIPS/Register/register[25][12] ), .S0(
        n5571), .Y(\i_MIPS/Register/n320 ) );
  CLKMX2X2 U12553 ( .A(n5446), .B(\i_MIPS/Register/register[25][11] ), .S0(
        n5570), .Y(\i_MIPS/Register/n319 ) );
  CLKMX2X2 U12554 ( .A(n5420), .B(\i_MIPS/Register/register[25][10] ), .S0(
        n5570), .Y(\i_MIPS/Register/n318 ) );
  CLKMX2X2 U12555 ( .A(n5475), .B(\i_MIPS/Register/register[25][8] ), .S0(
        n5571), .Y(\i_MIPS/Register/n316 ) );
  CLKMX2X2 U12556 ( .A(n5472), .B(\i_MIPS/Register/register[25][7] ), .S0(
        n5571), .Y(\i_MIPS/Register/n315 ) );
  CLKMX2X2 U12557 ( .A(n5042), .B(\i_MIPS/Register/register[25][6] ), .S0(
        n5570), .Y(\i_MIPS/Register/n314 ) );
  CLKMX2X2 U12558 ( .A(n5491), .B(\i_MIPS/Register/register[25][5] ), .S0(
        n5570), .Y(\i_MIPS/Register/n313 ) );
  CLKMX2X2 U12559 ( .A(n5488), .B(\i_MIPS/Register/register[25][4] ), .S0(
        n5570), .Y(\i_MIPS/Register/n312 ) );
  CLKMX2X2 U12560 ( .A(n4776), .B(\i_MIPS/Register/register[25][3] ), .S0(
        n5570), .Y(\i_MIPS/Register/n311 ) );
  CLKMX2X2 U12561 ( .A(n5480), .B(\i_MIPS/Register/register[25][2] ), .S0(
        n5570), .Y(\i_MIPS/Register/n310 ) );
  CLKMX2X2 U12562 ( .A(n5477), .B(\i_MIPS/Register/register[25][1] ), .S0(
        n5571), .Y(\i_MIPS/Register/n309 ) );
  CLKMX2X2 U12563 ( .A(n5485), .B(\i_MIPS/Register/register[25][0] ), .S0(
        n5571), .Y(\i_MIPS/Register/n308 ) );
  CLKMX2X2 U12564 ( .A(n5470), .B(\i_MIPS/Register/register[26][31] ), .S0(
        n5568), .Y(\i_MIPS/Register/n307 ) );
  CLKMX2X2 U12565 ( .A(n5411), .B(\i_MIPS/Register/register[26][28] ), .S0(
        n5569), .Y(\i_MIPS/Register/n304 ) );
  CLKMX2X2 U12566 ( .A(n5408), .B(\i_MIPS/Register/register[26][27] ), .S0(
        n5568), .Y(\i_MIPS/Register/n303 ) );
  CLKMX2X2 U12567 ( .A(n5405), .B(\i_MIPS/Register/register[26][26] ), .S0(
        n5568), .Y(\i_MIPS/Register/n302 ) );
  CLKMX2X2 U12568 ( .A(n5414), .B(\i_MIPS/Register/register[26][25] ), .S0(
        n5569), .Y(\i_MIPS/Register/n301 ) );
  CLKMX2X2 U12569 ( .A(n5483), .B(\i_MIPS/Register/register[26][23] ), .S0(
        n5569), .Y(\i_MIPS/Register/n299 ) );
  CLKMX2X2 U12570 ( .A(n5423), .B(\i_MIPS/Register/register[26][22] ), .S0(
        n5568), .Y(\i_MIPS/Register/n298 ) );
  CLKMX2X2 U12571 ( .A(n5432), .B(\i_MIPS/Register/register[26][19] ), .S0(
        n5568), .Y(\i_MIPS/Register/n295 ) );
  CLKMX2X2 U12572 ( .A(n5417), .B(\i_MIPS/Register/register[26][18] ), .S0(
        n5569), .Y(\i_MIPS/Register/n294 ) );
  CLKMX2X2 U12573 ( .A(n5458), .B(\i_MIPS/Register/register[26][17] ), .S0(
        n5569), .Y(\i_MIPS/Register/n293 ) );
  CLKMX2X2 U12574 ( .A(n5456), .B(\i_MIPS/Register/register[26][15] ), .S0(
        n5569), .Y(\i_MIPS/Register/n291 ) );
  CLKMX2X2 U12575 ( .A(n5454), .B(\i_MIPS/Register/register[26][14] ), .S0(
        n5569), .Y(\i_MIPS/Register/n290 ) );
  CLKMX2X2 U12576 ( .A(n5452), .B(\i_MIPS/Register/register[26][13] ), .S0(
        n5569), .Y(\i_MIPS/Register/n289 ) );
  CLKMX2X2 U12577 ( .A(n5449), .B(\i_MIPS/Register/register[26][12] ), .S0(
        n5569), .Y(\i_MIPS/Register/n288 ) );
  CLKMX2X2 U12578 ( .A(n5446), .B(\i_MIPS/Register/register[26][11] ), .S0(
        n5568), .Y(\i_MIPS/Register/n287 ) );
  CLKMX2X2 U12579 ( .A(n5420), .B(\i_MIPS/Register/register[26][10] ), .S0(
        n5568), .Y(\i_MIPS/Register/n286 ) );
  CLKMX2X2 U12580 ( .A(n5475), .B(\i_MIPS/Register/register[26][8] ), .S0(
        n5569), .Y(\i_MIPS/Register/n284 ) );
  CLKMX2X2 U12581 ( .A(n5472), .B(\i_MIPS/Register/register[26][7] ), .S0(
        n5569), .Y(\i_MIPS/Register/n283 ) );
  CLKMX2X2 U12582 ( .A(n5043), .B(\i_MIPS/Register/register[26][6] ), .S0(
        n5568), .Y(\i_MIPS/Register/n282 ) );
  CLKMX2X2 U12583 ( .A(n5491), .B(\i_MIPS/Register/register[26][5] ), .S0(
        n5568), .Y(\i_MIPS/Register/n281 ) );
  CLKMX2X2 U12584 ( .A(n5488), .B(\i_MIPS/Register/register[26][4] ), .S0(
        n5568), .Y(\i_MIPS/Register/n280 ) );
  CLKMX2X2 U12585 ( .A(n4776), .B(\i_MIPS/Register/register[26][3] ), .S0(
        n5568), .Y(\i_MIPS/Register/n279 ) );
  CLKMX2X2 U12586 ( .A(n5480), .B(\i_MIPS/Register/register[26][2] ), .S0(
        n5568), .Y(\i_MIPS/Register/n278 ) );
  CLKMX2X2 U12587 ( .A(n5477), .B(\i_MIPS/Register/register[26][1] ), .S0(
        n5569), .Y(\i_MIPS/Register/n277 ) );
  CLKMX2X2 U12588 ( .A(n5485), .B(\i_MIPS/Register/register[26][0] ), .S0(
        n5569), .Y(\i_MIPS/Register/n276 ) );
  CLKMX2X2 U12589 ( .A(n5470), .B(\i_MIPS/Register/register[27][31] ), .S0(
        n5566), .Y(\i_MIPS/Register/n275 ) );
  CLKMX2X2 U12590 ( .A(n5411), .B(\i_MIPS/Register/register[27][28] ), .S0(
        n5567), .Y(\i_MIPS/Register/n272 ) );
  CLKMX2X2 U12591 ( .A(n5408), .B(\i_MIPS/Register/register[27][27] ), .S0(
        n5566), .Y(\i_MIPS/Register/n271 ) );
  CLKMX2X2 U12592 ( .A(n5405), .B(\i_MIPS/Register/register[27][26] ), .S0(
        n5566), .Y(\i_MIPS/Register/n270 ) );
  CLKMX2X2 U12593 ( .A(n5414), .B(\i_MIPS/Register/register[27][25] ), .S0(
        n5567), .Y(\i_MIPS/Register/n269 ) );
  CLKMX2X2 U12594 ( .A(n5483), .B(\i_MIPS/Register/register[27][23] ), .S0(
        n5567), .Y(\i_MIPS/Register/n267 ) );
  CLKMX2X2 U12595 ( .A(n5423), .B(\i_MIPS/Register/register[27][22] ), .S0(
        n5566), .Y(\i_MIPS/Register/n266 ) );
  CLKMX2X2 U12596 ( .A(n5432), .B(\i_MIPS/Register/register[27][19] ), .S0(
        n5566), .Y(\i_MIPS/Register/n263 ) );
  CLKMX2X2 U12597 ( .A(n5416), .B(\i_MIPS/Register/register[27][18] ), .S0(
        n5567), .Y(\i_MIPS/Register/n262 ) );
  CLKMX2X2 U12598 ( .A(n5458), .B(\i_MIPS/Register/register[27][17] ), .S0(
        n5567), .Y(\i_MIPS/Register/n261 ) );
  CLKMX2X2 U12599 ( .A(n5456), .B(\i_MIPS/Register/register[27][15] ), .S0(
        n5567), .Y(\i_MIPS/Register/n259 ) );
  CLKMX2X2 U12600 ( .A(n5454), .B(\i_MIPS/Register/register[27][14] ), .S0(
        n5567), .Y(\i_MIPS/Register/n258 ) );
  CLKMX2X2 U12601 ( .A(n5452), .B(\i_MIPS/Register/register[27][13] ), .S0(
        n5567), .Y(\i_MIPS/Register/n257 ) );
  CLKMX2X2 U12602 ( .A(n5448), .B(\i_MIPS/Register/register[27][12] ), .S0(
        n5567), .Y(\i_MIPS/Register/n256 ) );
  CLKMX2X2 U12603 ( .A(n5446), .B(\i_MIPS/Register/register[27][11] ), .S0(
        n5566), .Y(\i_MIPS/Register/n255 ) );
  CLKMX2X2 U12604 ( .A(n5420), .B(\i_MIPS/Register/register[27][10] ), .S0(
        n5566), .Y(\i_MIPS/Register/n254 ) );
  CLKMX2X2 U12605 ( .A(n5475), .B(\i_MIPS/Register/register[27][8] ), .S0(
        n5567), .Y(\i_MIPS/Register/n252 ) );
  CLKMX2X2 U12606 ( .A(n5472), .B(\i_MIPS/Register/register[27][7] ), .S0(
        n5567), .Y(\i_MIPS/Register/n251 ) );
  CLKMX2X2 U12607 ( .A(n5043), .B(\i_MIPS/Register/register[27][6] ), .S0(
        n5566), .Y(\i_MIPS/Register/n250 ) );
  CLKMX2X2 U12608 ( .A(n5490), .B(\i_MIPS/Register/register[27][5] ), .S0(
        n5566), .Y(\i_MIPS/Register/n249 ) );
  CLKMX2X2 U12609 ( .A(n5488), .B(\i_MIPS/Register/register[27][4] ), .S0(
        n5566), .Y(\i_MIPS/Register/n248 ) );
  CLKMX2X2 U12610 ( .A(n4776), .B(\i_MIPS/Register/register[27][3] ), .S0(
        n5566), .Y(\i_MIPS/Register/n247 ) );
  CLKMX2X2 U12611 ( .A(n5480), .B(\i_MIPS/Register/register[27][2] ), .S0(
        n5566), .Y(\i_MIPS/Register/n246 ) );
  CLKMX2X2 U12612 ( .A(n5477), .B(\i_MIPS/Register/register[27][1] ), .S0(
        n5567), .Y(\i_MIPS/Register/n245 ) );
  CLKMX2X2 U12613 ( .A(n5484), .B(\i_MIPS/Register/register[27][0] ), .S0(
        n5567), .Y(\i_MIPS/Register/n244 ) );
  CLKMX2X2 U12614 ( .A(n5470), .B(\i_MIPS/Register/register[28][31] ), .S0(
        n5564), .Y(\i_MIPS/Register/n243 ) );
  CLKMX2X2 U12615 ( .A(n5411), .B(\i_MIPS/Register/register[28][28] ), .S0(
        n5565), .Y(\i_MIPS/Register/n240 ) );
  CLKMX2X2 U12616 ( .A(n5408), .B(\i_MIPS/Register/register[28][27] ), .S0(
        n5564), .Y(\i_MIPS/Register/n239 ) );
  CLKMX2X2 U12617 ( .A(n5405), .B(\i_MIPS/Register/register[28][26] ), .S0(
        n5564), .Y(\i_MIPS/Register/n238 ) );
  CLKMX2X2 U12618 ( .A(n5414), .B(\i_MIPS/Register/register[28][25] ), .S0(
        n5565), .Y(\i_MIPS/Register/n237 ) );
  CLKMX2X2 U12619 ( .A(n5483), .B(\i_MIPS/Register/register[28][23] ), .S0(
        n5565), .Y(\i_MIPS/Register/n235 ) );
  CLKMX2X2 U12620 ( .A(n5423), .B(\i_MIPS/Register/register[28][22] ), .S0(
        n5564), .Y(\i_MIPS/Register/n234 ) );
  CLKMX2X2 U12621 ( .A(n5432), .B(\i_MIPS/Register/register[28][19] ), .S0(
        n5564), .Y(\i_MIPS/Register/n231 ) );
  CLKMX2X2 U12622 ( .A(n5417), .B(\i_MIPS/Register/register[28][18] ), .S0(
        n5565), .Y(\i_MIPS/Register/n230 ) );
  CLKMX2X2 U12623 ( .A(n5458), .B(\i_MIPS/Register/register[28][17] ), .S0(
        n5565), .Y(\i_MIPS/Register/n229 ) );
  CLKMX2X2 U12624 ( .A(n5456), .B(\i_MIPS/Register/register[28][15] ), .S0(
        n5565), .Y(\i_MIPS/Register/n227 ) );
  CLKMX2X2 U12625 ( .A(n5454), .B(\i_MIPS/Register/register[28][14] ), .S0(
        n5565), .Y(\i_MIPS/Register/n226 ) );
  CLKMX2X2 U12626 ( .A(n5452), .B(\i_MIPS/Register/register[28][13] ), .S0(
        n5565), .Y(\i_MIPS/Register/n225 ) );
  CLKMX2X2 U12627 ( .A(n5449), .B(\i_MIPS/Register/register[28][12] ), .S0(
        n5565), .Y(\i_MIPS/Register/n224 ) );
  CLKMX2X2 U12628 ( .A(n5446), .B(\i_MIPS/Register/register[28][11] ), .S0(
        n5564), .Y(\i_MIPS/Register/n223 ) );
  CLKMX2X2 U12629 ( .A(n5420), .B(\i_MIPS/Register/register[28][10] ), .S0(
        n5564), .Y(\i_MIPS/Register/n222 ) );
  CLKMX2X2 U12630 ( .A(n5475), .B(\i_MIPS/Register/register[28][8] ), .S0(
        n5565), .Y(\i_MIPS/Register/n220 ) );
  CLKMX2X2 U12631 ( .A(n5472), .B(\i_MIPS/Register/register[28][7] ), .S0(
        n5565), .Y(\i_MIPS/Register/n219 ) );
  CLKMX2X2 U12632 ( .A(n5042), .B(\i_MIPS/Register/register[28][6] ), .S0(
        n5564), .Y(\i_MIPS/Register/n218 ) );
  CLKMX2X2 U12633 ( .A(n5491), .B(\i_MIPS/Register/register[28][5] ), .S0(
        n5564), .Y(\i_MIPS/Register/n217 ) );
  CLKMX2X2 U12634 ( .A(n5488), .B(\i_MIPS/Register/register[28][4] ), .S0(
        n5564), .Y(\i_MIPS/Register/n216 ) );
  CLKMX2X2 U12635 ( .A(n4776), .B(\i_MIPS/Register/register[28][3] ), .S0(
        n5564), .Y(\i_MIPS/Register/n215 ) );
  CLKMX2X2 U12636 ( .A(n5480), .B(\i_MIPS/Register/register[28][2] ), .S0(
        n5564), .Y(\i_MIPS/Register/n214 ) );
  CLKMX2X2 U12637 ( .A(n5477), .B(\i_MIPS/Register/register[28][1] ), .S0(
        n5565), .Y(\i_MIPS/Register/n213 ) );
  CLKMX2X2 U12638 ( .A(n5485), .B(\i_MIPS/Register/register[28][0] ), .S0(
        n5565), .Y(\i_MIPS/Register/n212 ) );
  CLKMX2X2 U12639 ( .A(n5469), .B(\i_MIPS/Register/register[29][31] ), .S0(
        n5562), .Y(\i_MIPS/Register/n211 ) );
  CLKMX2X2 U12640 ( .A(n5410), .B(\i_MIPS/Register/register[29][28] ), .S0(
        n5563), .Y(\i_MIPS/Register/n208 ) );
  CLKMX2X2 U12641 ( .A(n5407), .B(\i_MIPS/Register/register[29][27] ), .S0(
        n5562), .Y(\i_MIPS/Register/n207 ) );
  CLKMX2X2 U12642 ( .A(n5404), .B(\i_MIPS/Register/register[29][26] ), .S0(
        n5562), .Y(\i_MIPS/Register/n206 ) );
  CLKMX2X2 U12643 ( .A(n5413), .B(\i_MIPS/Register/register[29][25] ), .S0(
        n5563), .Y(\i_MIPS/Register/n205 ) );
  CLKMX2X2 U12644 ( .A(n5482), .B(\i_MIPS/Register/register[29][23] ), .S0(
        n5563), .Y(\i_MIPS/Register/n203 ) );
  CLKMX2X2 U12645 ( .A(n5422), .B(\i_MIPS/Register/register[29][22] ), .S0(
        n5562), .Y(\i_MIPS/Register/n202 ) );
  CLKMX2X2 U12646 ( .A(n5431), .B(\i_MIPS/Register/register[29][19] ), .S0(
        n5562), .Y(\i_MIPS/Register/n199 ) );
  CLKMX2X2 U12647 ( .A(n5417), .B(\i_MIPS/Register/register[29][18] ), .S0(
        n5563), .Y(\i_MIPS/Register/n198 ) );
  CLKMX2X2 U12648 ( .A(n5457), .B(\i_MIPS/Register/register[29][17] ), .S0(
        n5563), .Y(\i_MIPS/Register/n197 ) );
  CLKMX2X2 U12649 ( .A(n5455), .B(\i_MIPS/Register/register[29][15] ), .S0(
        n5563), .Y(\i_MIPS/Register/n195 ) );
  CLKMX2X2 U12650 ( .A(n5453), .B(\i_MIPS/Register/register[29][14] ), .S0(
        n5563), .Y(\i_MIPS/Register/n194 ) );
  CLKMX2X2 U12651 ( .A(n5451), .B(\i_MIPS/Register/register[29][13] ), .S0(
        n5563), .Y(\i_MIPS/Register/n193 ) );
  CLKMX2X2 U12652 ( .A(n5449), .B(\i_MIPS/Register/register[29][12] ), .S0(
        n5563), .Y(\i_MIPS/Register/n192 ) );
  CLKMX2X2 U12653 ( .A(n5445), .B(\i_MIPS/Register/register[29][11] ), .S0(
        n5562), .Y(\i_MIPS/Register/n191 ) );
  CLKMX2X2 U12654 ( .A(n5419), .B(\i_MIPS/Register/register[29][10] ), .S0(
        n5562), .Y(\i_MIPS/Register/n190 ) );
  CLKMX2X2 U12655 ( .A(n5474), .B(\i_MIPS/Register/register[29][8] ), .S0(
        n5563), .Y(\i_MIPS/Register/n188 ) );
  CLKMX2X2 U12656 ( .A(n5471), .B(\i_MIPS/Register/register[29][7] ), .S0(
        n5563), .Y(\i_MIPS/Register/n187 ) );
  CLKMX2X2 U12657 ( .A(n5043), .B(\i_MIPS/Register/register[29][6] ), .S0(
        n5562), .Y(\i_MIPS/Register/n186 ) );
  CLKMX2X2 U12658 ( .A(n5491), .B(\i_MIPS/Register/register[29][5] ), .S0(
        n5562), .Y(\i_MIPS/Register/n185 ) );
  CLKMX2X2 U12659 ( .A(n5487), .B(\i_MIPS/Register/register[29][4] ), .S0(
        n5562), .Y(\i_MIPS/Register/n184 ) );
  CLKMX2X2 U12660 ( .A(n4775), .B(\i_MIPS/Register/register[29][3] ), .S0(
        n5562), .Y(\i_MIPS/Register/n183 ) );
  CLKMX2X2 U12661 ( .A(n5479), .B(\i_MIPS/Register/register[29][2] ), .S0(
        n5562), .Y(\i_MIPS/Register/n182 ) );
  CLKMX2X2 U12662 ( .A(n5476), .B(\i_MIPS/Register/register[29][1] ), .S0(
        n5563), .Y(\i_MIPS/Register/n181 ) );
  CLKMX2X2 U12663 ( .A(n5485), .B(\i_MIPS/Register/register[29][0] ), .S0(
        n5563), .Y(\i_MIPS/Register/n180 ) );
  CLKMX2X2 U12664 ( .A(n5470), .B(\i_MIPS/Register/register[30][31] ), .S0(
        n5560), .Y(\i_MIPS/Register/n179 ) );
  CLKMX2X2 U12665 ( .A(n5411), .B(\i_MIPS/Register/register[30][28] ), .S0(
        n5561), .Y(\i_MIPS/Register/n176 ) );
  CLKMX2X2 U12666 ( .A(n5408), .B(\i_MIPS/Register/register[30][27] ), .S0(
        n5560), .Y(\i_MIPS/Register/n175 ) );
  CLKMX2X2 U12667 ( .A(n5405), .B(\i_MIPS/Register/register[30][26] ), .S0(
        n5560), .Y(\i_MIPS/Register/n174 ) );
  CLKMX2X2 U12668 ( .A(n5414), .B(\i_MIPS/Register/register[30][25] ), .S0(
        n5561), .Y(\i_MIPS/Register/n173 ) );
  CLKMX2X2 U12669 ( .A(n5483), .B(\i_MIPS/Register/register[30][23] ), .S0(
        n5561), .Y(\i_MIPS/Register/n171 ) );
  CLKMX2X2 U12670 ( .A(n5423), .B(\i_MIPS/Register/register[30][22] ), .S0(
        n5560), .Y(\i_MIPS/Register/n170 ) );
  CLKMX2X2 U12671 ( .A(n5432), .B(\i_MIPS/Register/register[30][19] ), .S0(
        n5560), .Y(\i_MIPS/Register/n167 ) );
  CLKMX2X2 U12672 ( .A(n5417), .B(\i_MIPS/Register/register[30][18] ), .S0(
        n5561), .Y(\i_MIPS/Register/n166 ) );
  CLKMX2X2 U12673 ( .A(n5458), .B(\i_MIPS/Register/register[30][17] ), .S0(
        n5561), .Y(\i_MIPS/Register/n165 ) );
  CLKMX2X2 U12674 ( .A(n5456), .B(\i_MIPS/Register/register[30][15] ), .S0(
        n5561), .Y(\i_MIPS/Register/n163 ) );
  CLKMX2X2 U12675 ( .A(n5454), .B(\i_MIPS/Register/register[30][14] ), .S0(
        n5561), .Y(\i_MIPS/Register/n162 ) );
  CLKMX2X2 U12676 ( .A(n5452), .B(\i_MIPS/Register/register[30][13] ), .S0(
        n5561), .Y(\i_MIPS/Register/n161 ) );
  CLKMX2X2 U12677 ( .A(n5449), .B(\i_MIPS/Register/register[30][12] ), .S0(
        n5561), .Y(\i_MIPS/Register/n160 ) );
  CLKMX2X2 U12678 ( .A(n5446), .B(\i_MIPS/Register/register[30][11] ), .S0(
        n5560), .Y(\i_MIPS/Register/n159 ) );
  CLKMX2X2 U12679 ( .A(n5420), .B(\i_MIPS/Register/register[30][10] ), .S0(
        n5560), .Y(\i_MIPS/Register/n158 ) );
  CLKMX2X2 U12680 ( .A(n5475), .B(\i_MIPS/Register/register[30][8] ), .S0(
        n5561), .Y(\i_MIPS/Register/n156 ) );
  CLKMX2X2 U12681 ( .A(n5472), .B(\i_MIPS/Register/register[30][7] ), .S0(
        n5561), .Y(\i_MIPS/Register/n155 ) );
  CLKMX2X2 U12682 ( .A(n5043), .B(\i_MIPS/Register/register[30][6] ), .S0(
        n5560), .Y(\i_MIPS/Register/n154 ) );
  CLKMX2X2 U12683 ( .A(n5491), .B(\i_MIPS/Register/register[30][5] ), .S0(
        n5560), .Y(\i_MIPS/Register/n153 ) );
  CLKMX2X2 U12684 ( .A(n5488), .B(\i_MIPS/Register/register[30][4] ), .S0(
        n5560), .Y(\i_MIPS/Register/n152 ) );
  CLKMX2X2 U12685 ( .A(n4776), .B(\i_MIPS/Register/register[30][3] ), .S0(
        n5560), .Y(\i_MIPS/Register/n151 ) );
  CLKMX2X2 U12686 ( .A(n5480), .B(\i_MIPS/Register/register[30][2] ), .S0(
        n5560), .Y(\i_MIPS/Register/n150 ) );
  CLKMX2X2 U12687 ( .A(n5477), .B(\i_MIPS/Register/register[30][1] ), .S0(
        n5561), .Y(\i_MIPS/Register/n149 ) );
  CLKMX2X2 U12688 ( .A(n5485), .B(\i_MIPS/Register/register[30][0] ), .S0(
        n5561), .Y(\i_MIPS/Register/n148 ) );
  MX2XL U12689 ( .A(n3604), .B(n14), .S0(n219), .Y(\i_MIPS/n399 ) );
  MXI2X1 U12690 ( .A(n4536), .B(\i_MIPS/n224 ), .S0(n207), .Y(\i_MIPS/n503 )
         );
  MX2XL U12691 ( .A(net107796), .B(\i_MIPS/Sign_Extend_ID[8] ), .S0(n222), .Y(
        \i_MIPS/n504 ) );
  MX2XL U12692 ( .A(\i_MIPS/ID_EX[67] ), .B(n4592), .S0(n205), .Y(
        \i_MIPS/n385 ) );
  MX2XL U12693 ( .A(n3597), .B(n225), .S0(n205), .Y(\i_MIPS/n395 ) );
  MX2XL U12694 ( .A(n3598), .B(n11176), .S0(n216), .Y(\i_MIPS/n377 ) );
  MXI2XL U12695 ( .A(n4537), .B(\i_MIPS/n226 ), .S0(n205), .Y(\i_MIPS/n501 )
         );
  MX2XL U12696 ( .A(\i_MIPS/ID_EX[78] ), .B(\i_MIPS/Sign_Extend_ID[5] ), .S0(
        n217), .Y(\i_MIPS/n507 ) );
  MX2XL U12697 ( .A(n3812), .B(\i_MIPS/Sign_Extend_ID[1] ), .S0(n213), .Y(
        \i_MIPS/n511 ) );
  MX2XL U12698 ( .A(\i_MIPS/ID_EX[79] ), .B(\i_MIPS/Sign_Extend_ID[6] ), .S0(
        n219), .Y(\i_MIPS/n506 ) );
  MX2XL U12699 ( .A(\i_MIPS/ID_EX[77] ), .B(\i_MIPS/Sign_Extend_ID[4] ), .S0(
        n220), .Y(\i_MIPS/n508 ) );
  MX2XL U12700 ( .A(n3696), .B(\i_MIPS/Sign_Extend_ID[3] ), .S0(n214), .Y(
        \i_MIPS/n509 ) );
  MX2XL U12701 ( .A(n3608), .B(n4488), .S0(n219), .Y(\i_MIPS/n530 ) );
  MXI2XL U12702 ( .A(n4539), .B(\i_MIPS/n227 ), .S0(n210), .Y(\i_MIPS/n500 )
         );
  MX2XL U12703 ( .A(n12939), .B(n10652), .S0(n205), .Y(\i_MIPS/n449 ) );
  BUFX20 U12704 ( .A(ICACHE_addr[3]), .Y(n4661) );
  AO22X1 U12705 ( .A0(\i_MIPS/control_out[7] ), .A1(net108200), .B0(
        \i_MIPS/ALUOp[1] ), .B1(n202), .Y(\i_MIPS/n471 ) );
  AO22XL U12706 ( .A0(net108200), .A1(n9614), .B0(\i_MIPS/ID_EX_5 ), .B1(n202), 
        .Y(\i_MIPS/n478 ) );
  AO22X1 U12707 ( .A0(n5545), .A1(n11124), .B0(net112406), .B1(
        \i_MIPS/IR_ID[19] ), .Y(\i_MIPS/N77 ) );
  AO22X1 U12708 ( .A0(n4072), .A1(n10628), .B0(net112406), .B1(n9737), .Y(
        \i_MIPS/N74 ) );
  CLKINVX1 U12709 ( .A(\i_MIPS/n312 ), .Y(n9737) );
  AO22X1 U12710 ( .A0(n4073), .A1(n10532), .B0(net112406), .B1(n9688), .Y(
        \i_MIPS/N76 ) );
  CLKINVX1 U12711 ( .A(\i_MIPS/n316 ), .Y(n9688) );
  AO22X1 U12712 ( .A0(\i_MIPS/control_out[0] ), .A1(net108200), .B0(n202), 
        .B1(\i_MIPS/ID_EX_0 ), .Y(\i_MIPS/n528 ) );
  NAND3BX1 U12713 ( .AN(\i_MIPS/control_out[7] ), .B(n5558), .C(
        \i_MIPS/Control_ID/n12 ), .Y(\i_MIPS/control_out[0] ) );
  INVX12 U12714 ( .A(n408), .Y(mem_addr_D[6]) );
  AO21XL U12715 ( .A0(\i_MIPS/ID_EX[94] ), .A1(n202), .B0(n4380), .Y(
        \i_MIPS/n491 ) );
  AO21XL U12716 ( .A0(\i_MIPS/ID_EX[95] ), .A1(n202), .B0(n4380), .Y(
        \i_MIPS/n490 ) );
  AO21XL U12717 ( .A0(\i_MIPS/ID_EX[96] ), .A1(n202), .B0(n4380), .Y(
        \i_MIPS/n489 ) );
  AO21XL U12718 ( .A0(\i_MIPS/ID_EX[97] ), .A1(n202), .B0(n4380), .Y(
        \i_MIPS/n488 ) );
  AO21XL U12719 ( .A0(\i_MIPS/ID_EX[89] ), .A1(n202), .B0(n4380), .Y(
        \i_MIPS/n496 ) );
  AO21XL U12720 ( .A0(\i_MIPS/ID_EX[93] ), .A1(n202), .B0(n4380), .Y(
        \i_MIPS/n492 ) );
  AO21XL U12721 ( .A0(\i_MIPS/ID_EX[98] ), .A1(n202), .B0(n4380), .Y(
        \i_MIPS/n487 ) );
  AO21XL U12722 ( .A0(\i_MIPS/ID_EX[99] ), .A1(n202), .B0(n4380), .Y(
        \i_MIPS/n486 ) );
  AO21XL U12723 ( .A0(\i_MIPS/ID_EX[100] ), .A1(n202), .B0(n4380), .Y(
        \i_MIPS/n485 ) );
  AO21XL U12724 ( .A0(\i_MIPS/ID_EX[101] ), .A1(n202), .B0(n4380), .Y(
        \i_MIPS/n484 ) );
  AO21XL U12725 ( .A0(\i_MIPS/ID_EX[103] ), .A1(n202), .B0(n4380), .Y(
        \i_MIPS/n482 ) );
  AO21XL U12726 ( .A0(\i_MIPS/ID_EX[104] ), .A1(n202), .B0(n4380), .Y(
        \i_MIPS/n481 ) );
  AO21XL U12727 ( .A0(n202), .A1(n3609), .B0(n4452), .Y(\i_MIPS/n527 ) );
  AO21XL U12728 ( .A0(n202), .A1(\i_MIPS/ID_EX_3 ), .B0(n4452), .Y(
        \i_MIPS/n525 ) );
  NAND4X1 U12729 ( .A(n6443), .B(n6442), .C(n6441), .D(n6440), .Y(n6456) );
  XOR2XL U12730 ( .A(n6604), .B(\i_MIPS/IR_ID[19] ), .Y(n6610) );
  AND3X2 U12731 ( .A(\i_MIPS/Register/n120 ), .B(n4542), .C(\i_MIPS/Reg_W[3] ), 
        .Y(\i_MIPS/Register/n131 ) );
  AND3X2 U12732 ( .A(\i_MIPS/Register/n120 ), .B(n4543), .C(\i_MIPS/Reg_W[4] ), 
        .Y(\i_MIPS/Register/n122 ) );
  AND3X2 U12733 ( .A(\i_MIPS/Register/n120 ), .B(\i_MIPS/Reg_W[3] ), .C(
        \i_MIPS/Reg_W[4] ), .Y(\i_MIPS/Register/n104 ) );
  NAND3BX1 U12734 ( .AN(n9890), .B(\i_MIPS/IR_ID[29] ), .C(n9889), .Y(
        \i_MIPS/Control_ID/n15 ) );
  NAND2X1 U12735 ( .A(\i_MIPS/IR_ID[28] ), .B(\i_MIPS/n324 ), .Y(n9888) );
  XOR2XL U12736 ( .A(\i_MIPS/n313 ), .B(\i_MIPS/IR_ID[21] ), .Y(n9554) );
  XOR2XL U12737 ( .A(\i_MIPS/n317 ), .B(\i_MIPS/IR_ID[23] ), .Y(n9555) );
  XOR2XL U12738 ( .A(\i_MIPS/n313 ), .B(\i_MIPS/IR_ID[16] ), .Y(n9552) );
  XOR2XL U12739 ( .A(\i_MIPS/n317 ), .B(\i_MIPS/IR_ID[18] ), .Y(n9553) );
  NOR2BX1 U12740 ( .AN(\i_MIPS/EX_MEM_0 ), .B(\i_MIPS/EX_MEM_74 ), .Y(
        \i_MIPS/Register/n120 ) );
  NAND3BX1 U12741 ( .AN(\i_MIPS/IR_ID[29] ), .B(\i_MIPS/n326 ), .C(
        \i_MIPS/n330 ), .Y(n9567) );
  NAND4X1 U12742 ( .A(n6239), .B(n6238), .C(\i_MIPS/n216 ), .D(n6237), .Y(
        n10375) );
  NOR2X1 U12743 ( .A(\i_MIPS/Sign_Extend_ID[0] ), .B(
        \i_MIPS/Sign_Extend_ID[5] ), .Y(n6238) );
  NOR2X1 U12744 ( .A(\i_MIPS/Sign_Extend_ID[4] ), .B(
        \i_MIPS/Sign_Extend_ID[2] ), .Y(n6237) );
  NAND2X1 U12745 ( .A(\i_MIPS/PHT_2/history_state[0] ), .B(\i_MIPS/PHT_2/n12 ), 
        .Y(n11046) );
  NAND2X1 U12746 ( .A(\i_MIPS/PHT_2/n12 ), .B(\i_MIPS/PHT_2/n13 ), .Y(n11047)
         );
  NOR2BX1 U12747 ( .AN(\i_MIPS/Sign_Extend_ID[3] ), .B(\i_MIPS/Control_ID/n10 ), .Y(n6239) );
  AND2X2 U12748 ( .A(\i_MIPS/IR_ID[27] ), .B(\i_MIPS/IR_ID[26] ), .Y(n4544) );
  CLKBUFX3 U12749 ( .A(\i_MIPS/IR_ID[25] ), .Y(net107816) );
  CLKBUFX3 U12750 ( .A(mem_ready_I), .Y(n4651) );
  NAND2X1 U12751 ( .A(\i_MIPS/PHT_2/current_state_0[1] ), .B(n11060), .Y(
        n11057) );
  NAND2X1 U12752 ( .A(\i_MIPS/PHT_2/current_state_1[1] ), .B(n11065), .Y(
        n11061) );
  AO21XL U12753 ( .A0(n4651), .A1(n5320), .B0(\I_cache/cache[7][154] ), .Y(
        n11548) );
  AO21XL U12754 ( .A0(n4651), .A1(n5362), .B0(\I_cache/cache[6][154] ), .Y(
        n11549) );
  AO21XL U12755 ( .A0(n4651), .A1(n5226), .B0(\I_cache/cache[5][154] ), .Y(
        n11550) );
  AO21XL U12756 ( .A0(n4651), .A1(n5273), .B0(\I_cache/cache[4][154] ), .Y(
        n11551) );
  AO21XL U12757 ( .A0(n4651), .A1(n5138), .B0(\I_cache/cache[3][154] ), .Y(
        n11552) );
  AO21XL U12758 ( .A0(n4651), .A1(n5184), .B0(\I_cache/cache[2][154] ), .Y(
        n11553) );
  AO21XL U12759 ( .A0(n4651), .A1(n5053), .B0(\I_cache/cache[1][154] ), .Y(
        n11554) );
  AO21XL U12760 ( .A0(n4651), .A1(n5098), .B0(\I_cache/cache[0][154] ), .Y(
        n11555) );
  AO22X1 U12761 ( .A0(ICACHE_addr[13]), .A1(n11512), .B0(n4657), .B1(n11328), 
        .Y(n12820) );
  AO22X1 U12762 ( .A0(ICACHE_addr[15]), .A1(n11512), .B0(n4656), .B1(n11330), 
        .Y(n12818) );
  AO22X1 U12763 ( .A0(ICACHE_addr[18]), .A1(n11512), .B0(mem_write_I), .B1(
        n11333), .Y(n12815) );
  AO22X1 U12764 ( .A0(ICACHE_addr[19]), .A1(n11512), .B0(mem_write_I), .B1(
        n11334), .Y(n12814) );
  AO22X1 U12765 ( .A0(ICACHE_addr[20]), .A1(n11512), .B0(mem_write_I), .B1(
        n11335), .Y(n12813) );
  AO22X1 U12766 ( .A0(ICACHE_addr[22]), .A1(n11512), .B0(mem_write_I), .B1(
        n11337), .Y(n12811) );
  AO22X1 U12767 ( .A0(ICACHE_addr[23]), .A1(n11512), .B0(mem_write_I), .B1(
        n11338), .Y(n12810) );
  AO22X1 U12768 ( .A0(ICACHE_addr[24]), .A1(n11512), .B0(mem_write_I), .B1(
        n11339), .Y(n12809) );
  AO22X1 U12769 ( .A0(ICACHE_addr[26]), .A1(n11512), .B0(mem_write_I), .B1(
        n11341), .Y(n12807) );
  AO22X1 U12770 ( .A0(ICACHE_addr[27]), .A1(n11512), .B0(mem_write_I), .B1(
        n11342), .Y(n12806) );
  AO22X1 U12771 ( .A0(ICACHE_addr[28]), .A1(n11512), .B0(mem_write_I), .B1(
        n11343), .Y(n12805) );
  AO22X1 U12772 ( .A0(ICACHE_addr[29]), .A1(n11512), .B0(mem_write_I), .B1(
        n11344), .Y(n12804) );
  MX2XL U12773 ( .A(n10680), .B(n3802), .S0(n211), .Y(\i_MIPS/n379 ) );
  NAND2XL U12774 ( .A(net112962), .B(n4673), .Y(net99002) );
  INVX12 U12775 ( .A(n4594), .Y(DCACHE_addr[10]) );
  INVX12 U12776 ( .A(n4596), .Y(DCACHE_addr[11]) );
  INVX12 U12777 ( .A(n4598), .Y(DCACHE_addr[15]) );
  OAI221XL U12778 ( .A0(net103249), .A1(net111624), .B0(net103250), .B1(
        net111636), .C0(net103251), .Y(n4601) );
  CLKINVX1 U12779 ( .A(n8239), .Y(n6569) );
  OAI221XL U12780 ( .A0(net105045), .A1(net111624), .B0(net105046), .B1(
        net111636), .C0(net105047), .Y(n4611) );
  OAI221XL U12781 ( .A0(n8724), .A1(net111622), .B0(n8723), .B1(net111634), 
        .C0(n8722), .Y(n4612) );
  OAI221XL U12782 ( .A0(net104251), .A1(net111624), .B0(net104252), .B1(
        net111636), .C0(net104253), .Y(n4613) );
  OAI221XL U12783 ( .A0(n8917), .A1(net111622), .B0(n3903), .B1(net111634), 
        .C0(n8916), .Y(n4619) );
  OAI221XL U12784 ( .A0(n8826), .A1(net111622), .B0(n8825), .B1(net111634), 
        .C0(n8824), .Y(n4621) );
  OAI221XL U12785 ( .A0(net103089), .A1(net111624), .B0(net103090), .B1(
        net111634), .C0(net103091), .Y(n4623) );
  NAND3BX4 U12786 ( .AN(\i_MIPS/PC/n22 ), .B(ICACHE_addr[17]), .C(n10283), .Y(
        n10328) );
  NAND3BX4 U12787 ( .AN(n11479), .B(n3854), .C(n11478), .Y(n11482) );
  OAI221XL U12788 ( .A0(net104105), .A1(net111624), .B0(net104106), .B1(
        net111636), .C0(net104107), .Y(n4627) );
  MX2XL U12789 ( .A(n3611), .B(n10208), .S0(n222), .Y(\i_MIPS/n393 ) );
  MX2XL U12790 ( .A(n12947), .B(n13), .S0(n204), .Y(\i_MIPS/n457 ) );
  INVX12 U12791 ( .A(n4629), .Y(DCACHE_addr[16]) );
  MX2XL U12792 ( .A(DCACHE_addr[12]), .B(net98029), .S0(n210), .Y(
        \i_MIPS/n455 ) );
  NAND2XL U12793 ( .A(n12943), .B(\i_MIPS/n336 ), .Y(n10287) );
  AO22X2 U12794 ( .A0(n5528), .A1(DCACHE_addr[23]), .B0(n5527), .B1(n11501), 
        .Y(n11033) );
  MX2XL U12795 ( .A(n12946), .B(n241), .S0(n223), .Y(\i_MIPS/n456 ) );
  INVX12 U12796 ( .A(n4631), .Y(DCACHE_addr[21]) );
  INVX12 U12797 ( .A(n4633), .Y(DCACHE_addr[17]) );
  MX2XL U12798 ( .A(n12943), .B(n3807), .S0(n214), .Y(\i_MIPS/n453 ) );
  MX2XL U12799 ( .A(n12940), .B(n3809), .S0(n208), .Y(\i_MIPS/n450 ) );
  NAND2XL U12800 ( .A(n12940), .B(n4673), .Y(n10152) );
  NAND2XL U12801 ( .A(n12936), .B(n4674), .Y(n10559) );
  XNOR2X4 U12802 ( .A(n11503), .B(DCACHE_addr[25]), .Y(n4638) );
  NAND2X1 U12803 ( .A(n7684), .B(n3688), .Y(n7414) );
  NAND2X1 U12804 ( .A(DCACHE_addr[1]), .B(\i_MIPS/n336 ), .Y(n9978) );
  OAI2BB2X4 U12805 ( .B0(n6601), .B1(n6602), .A0N(n6600), .A1N(n6599), .Y(
        n10787) );
  AOI2BB2X1 U12806 ( .B0(DCACHE_addr[29]), .B1(mem_read_D), .A0N(n4649), .A1N(
        n4650), .Y(n4648) );
  NAND2X4 U12807 ( .A(n6041), .B(n6040), .Y(n6042) );
  OA22X4 U12808 ( .A0(n5104), .A1(n1724), .B0(n5065), .B1(n3406), .Y(n6114) );
  OA22X4 U12809 ( .A0(n5195), .A1(n1725), .B0(n5152), .B1(n3407), .Y(n6113) );
  OA22X4 U12810 ( .A0(n5306), .A1(n3334), .B0(n5240), .B1(n1727), .Y(n6112) );
  OA22X4 U12811 ( .A0(n5394), .A1(n3408), .B0(n5331), .B1(n1775), .Y(n6111) );
  CLKINVX3 U12812 ( .A(n10223), .Y(n10065) );
  OR2X8 U12813 ( .A(n6312), .B(n6311), .Y(n11345) );
  NAND4X2 U12814 ( .A(n6320), .B(n6319), .C(n6318), .D(n6317), .Y(n11380) );
  OA22X4 U12815 ( .A0(n4837), .A1(n3372), .B0(n4883), .B1(n1743), .Y(n6325) );
  OAI221X2 U12816 ( .A0(n4764), .A1(n3346), .B0(n4798), .B1(n1731), .C0(n6325), 
        .Y(n6326) );
  OA22X4 U12817 ( .A0(n4989), .A1(n3373), .B0(n5035), .B1(n1744), .Y(n6327) );
  OAI221X2 U12818 ( .A0(n4770), .A1(n3347), .B0(n4797), .B1(n405), .C0(n6328), 
        .Y(n6329) );
  OAI221X2 U12819 ( .A0(n4902), .A1(n3344), .B0(n4945), .B1(n1730), .C0(n6330), 
        .Y(n6331) );
  OAI221X2 U12820 ( .A0(n4765), .A1(n3348), .B0(n4787), .B1(n1732), .C0(n6333), 
        .Y(n6334) );
  OA22X4 U12821 ( .A0(n4993), .A1(n3374), .B0(n5034), .B1(n1745), .Y(n6335) );
  OAI221X2 U12822 ( .A0(n4903), .A1(n3349), .B0(n4946), .B1(n1733), .C0(n6335), 
        .Y(n6336) );
  OA22X4 U12823 ( .A0(n4835), .A1(n3375), .B0(n4881), .B1(n1746), .Y(n6355) );
  OA22X4 U12824 ( .A0(n4988), .A1(n3377), .B0(n5036), .B1(n1748), .Y(n6353) );
  OA22X4 U12825 ( .A0(n4835), .A1(n3378), .B0(n4881), .B1(n1749), .Y(n6359) );
  OA22X4 U12826 ( .A0(n4926), .A1(n3379), .B0(n4953), .B1(n1750), .Y(n6358) );
  OA22X4 U12827 ( .A0(n4988), .A1(n3380), .B0(n5034), .B1(n1751), .Y(n6357) );
  OA22X4 U12828 ( .A0(n4835), .A1(n3381), .B0(n4881), .B1(n1752), .Y(n6362) );
  OA22X4 U12829 ( .A0(n4926), .A1(n3382), .B0(n4955), .B1(n1753), .Y(n6361) );
  OA22X4 U12830 ( .A0(n4988), .A1(n3383), .B0(n5037), .B1(n1754), .Y(n6360) );
  OA22X4 U12831 ( .A0(n4835), .A1(n3384), .B0(n4881), .B1(n1755), .Y(n6365) );
  OA22X4 U12832 ( .A0(n4926), .A1(n3385), .B0(n4955), .B1(n1756), .Y(n6364) );
  OA22X4 U12833 ( .A0(n4988), .A1(n3386), .B0(n5036), .B1(n1757), .Y(n6363) );
  OA22X4 U12834 ( .A0(n4763), .A1(n631), .B0(n4796), .B1(n3361), .Y(n6372) );
  OA22X4 U12835 ( .A0(n4835), .A1(n632), .B0(n4881), .B1(n3362), .Y(n6371) );
  OA22X4 U12836 ( .A0(n4925), .A1(n3387), .B0(n4950), .B1(n1758), .Y(n6370) );
  OA22X4 U12837 ( .A0(n4988), .A1(n3388), .B0(n5033), .B1(n1759), .Y(n6369) );
  XNOR2X4 U12838 ( .A(n12947), .B(n11488), .Y(n6388) );
  OA22X4 U12839 ( .A0(n4763), .A1(n633), .B0(n4796), .B1(n3363), .Y(n6376) );
  OA22X4 U12840 ( .A0(n4925), .A1(n3390), .B0(n4950), .B1(n1761), .Y(n6374) );
  XNOR2X4 U12841 ( .A(n11489), .B(n12946), .Y(n6387) );
  OA22X4 U12842 ( .A0(n4925), .A1(n3392), .B0(n4950), .B1(n1763), .Y(n6378) );
  OA22X4 U12843 ( .A0(n4763), .A1(n634), .B0(n4796), .B1(n3364), .Y(n6384) );
  OA22X4 U12844 ( .A0(n4925), .A1(n3393), .B0(n4955), .B1(n1764), .Y(n6382) );
  XNOR2X4 U12845 ( .A(n12942), .B(n11493), .Y(n6385) );
  OA22X4 U12846 ( .A0(n4986), .A1(n636), .B0(n5032), .B1(n3365), .Y(n6409) );
  OAI31X2 U12847 ( .A0(n6445), .A1(n9886), .A2(n9884), .B0(\i_MIPS/ID_EX_0 ), 
        .Y(n6446) );
  NAND4BBX4 U12848 ( .AN(n6456), .BN(n6455), .C(\i_MIPS/EX_MEM_0 ), .D(n6454), 
        .Y(net100478) );
  NAND2X2 U12849 ( .A(n6544), .B(\i_MIPS/ALUin1[10] ), .Y(n7308) );
  NAND2X2 U12850 ( .A(n3841), .B(\i_MIPS/n348 ), .Y(n8849) );
  NAND2X2 U12851 ( .A(n8849), .B(n8253), .Y(n6520) );
  NAND2X2 U12852 ( .A(n6571), .B(\i_MIPS/n350 ), .Y(n9487) );
  NAND2X2 U12853 ( .A(n6576), .B(\i_MIPS/n357 ), .Y(n7803) );
  NAND2X2 U12854 ( .A(\i_MIPS/ALUin1[22] ), .B(n6560), .Y(n9475) );
  NAND2X2 U12855 ( .A(\i_MIPS/ALUin1[24] ), .B(n6564), .Y(n8947) );
  OAI31X2 U12856 ( .A0(n9044), .A1(n11182), .A2(n8172), .B0(n6596), .Y(n6680)
         );
  AOI211X2 U12857 ( .A0(n6703), .A1(n6702), .B0(n6701), .C0(n6700), .Y(n6715)
         );
  XOR2X4 U12858 ( .A(n10880), .B(n10867), .Y(net105350) );
  CLKINVX3 U12859 ( .A(n6758), .Y(n6760) );
  NAND2X2 U12860 ( .A(net103354), .B(\i_MIPS/n340 ), .Y(n8350) );
  OAI221X2 U12861 ( .A0(net112366), .A1(\i_MIPS/n348 ), .B0(net112348), .B1(
        \i_MIPS/n349 ), .C0(n6837), .Y(n7473) );
  OA22X4 U12862 ( .A0(n4831), .A1(n2190), .B0(n4876), .B1(n616), .Y(n7007) );
  OA22X4 U12863 ( .A0(n4922), .A1(n3394), .B0(n4249), .B1(n1765), .Y(n7006) );
  OA22X4 U12864 ( .A0(n4983), .A1(n2191), .B0(n5029), .B1(n617), .Y(n7005) );
  OA22X4 U12865 ( .A0(n4758), .A1(n2192), .B0(n4794), .B1(n618), .Y(n7096) );
  OA22X4 U12866 ( .A0(n4830), .A1(n2193), .B0(n4875), .B1(n619), .Y(n7095) );
  OA22X4 U12867 ( .A0(n4982), .A1(n2194), .B0(n5028), .B1(n620), .Y(n7093) );
  OA22X4 U12868 ( .A0(n4921), .A1(n3396), .B0(n4949), .B1(n1767), .Y(n7269) );
  OA22X4 U12869 ( .A0(n4981), .A1(n2197), .B0(n5027), .B1(n623), .Y(n7268) );
  NAND4X2 U12870 ( .A(n7271), .B(n7270), .C(n7269), .D(n7268), .Y(n11425) );
  CLKINVX3 U12871 ( .A(net102427), .Y(net103891) );
  OA22X4 U12872 ( .A0(n4977), .A1(n2099), .B0(n5022), .B1(n514), .Y(n7841) );
  NAND4X2 U12873 ( .A(n7844), .B(n7843), .C(n7842), .D(n7841), .Y(n11431) );
  OA22X4 U12874 ( .A0(n4914), .A1(n3397), .B0(n4947), .B1(n1768), .Y(n8193) );
  OA22X4 U12875 ( .A0(n4975), .A1(n2072), .B0(n5020), .B1(n481), .Y(n8192) );
  OA22X4 U12876 ( .A0(n4913), .A1(n3398), .B0(n4249), .B1(n1769), .Y(n8389) );
  OA22X4 U12877 ( .A0(n4974), .A1(n2199), .B0(n5019), .B1(n625), .Y(n8388) );
  NAND4X2 U12878 ( .A(n8391), .B(n8390), .C(n8389), .D(n8388), .Y(n11449) );
  CLKINVX3 U12879 ( .A(n8864), .Y(n8548) );
  OA22X4 U12880 ( .A0(n4817), .A1(n2095), .B0(n4863), .B1(n508), .Y(n8887) );
  OA22X4 U12881 ( .A0(n4970), .A1(n2096), .B0(n5015), .B1(n509), .Y(n8885) );
  OA22X4 U12882 ( .A0(n4815), .A1(n2200), .B0(n4860), .B1(n626), .Y(n9294) );
  OA22X4 U12883 ( .A0(n4967), .A1(n2201), .B0(n185), .B1(n627), .Y(n9292) );
  OA22X4 U12884 ( .A0(n230), .A1(n3010), .B0(n5247), .B1(n1442), .Y(n9640) );
  OA22X4 U12885 ( .A0(n5111), .A1(n3011), .B0(n5072), .B1(n1443), .Y(n9647) );
  OA22X4 U12886 ( .A0(n5369), .A1(n3013), .B0(n5338), .B1(n1445), .Y(n9644) );
  OA22X4 U12887 ( .A0(n5112), .A1(n3323), .B0(n5054), .B1(n1722), .Y(n9657) );
  OA22X4 U12888 ( .A0(n9660), .A1(n5425), .B0(n9659), .B1(n5429), .Y(n9661) );
  NAND2X2 U12889 ( .A(n4462), .B(n10082), .Y(n10070) );
  AO21X4 U12890 ( .A0(n4303), .A1(n10072), .B0(n10070), .Y(n10990) );
  AO21X4 U12891 ( .A0(n4303), .A1(n10071), .B0(n10070), .Y(n10994) );
  CLKINVX3 U12892 ( .A(n10374), .Y(n10376) );
  NAND2X2 U12893 ( .A(\i_MIPS/IF_ID[97] ), .B(net108200), .Y(n11051) );
endmodule

