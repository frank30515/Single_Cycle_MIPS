
module CHIP ( clk, rst_n, mem_read_D, mem_write_D, mem_addr_D, mem_wdata_D, 
        mem_rdata_D, mem_ready_D, mem_read_I, mem_write_I, mem_addr_I, 
        mem_wdata_I, mem_rdata_I, mem_ready_I, DCACHE_addr, DCACHE_wdata, 
        DCACHE_wen );
  output [31:4] mem_addr_D;
  output [127:0] mem_wdata_D;
  input [127:0] mem_rdata_D;
  output [31:4] mem_addr_I;
  output [127:0] mem_wdata_I;
  input [127:0] mem_rdata_I;
  output [29:0] DCACHE_addr;
  output [31:0] DCACHE_wdata;
  input clk, rst_n, mem_ready_D, mem_ready_I;
  output mem_read_D, mem_write_D, mem_read_I, mem_write_I, DCACHE_wen;
  wire   n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831,
         n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839,
         n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847,
         n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855,
         n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863,
         n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871,
         n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879,
         n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
         n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895,
         n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903,
         n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911,
         n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919,
         n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927,
         n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935,
         n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943,
         n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951,
         n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959,
         n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967,
         n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975,
         n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983,
         n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991,
         n12992, n12993, n12994, n12995, n12996, n12997, DCACHE_ren,
         \i_MIPS/n563 , \i_MIPS/n562 , \i_MIPS/n561 , \i_MIPS/n560 ,
         \i_MIPS/n559 , \i_MIPS/n558 , \i_MIPS/n557 , \i_MIPS/n556 ,
         \i_MIPS/n555 , \i_MIPS/n554 , \i_MIPS/n553 , \i_MIPS/n552 ,
         \i_MIPS/n551 , \i_MIPS/n550 , \i_MIPS/n549 , \i_MIPS/n548 ,
         \i_MIPS/n547 , \i_MIPS/n546 , \i_MIPS/n545 , \i_MIPS/n544 ,
         \i_MIPS/n543 , \i_MIPS/n542 , \i_MIPS/n541 , \i_MIPS/n540 ,
         \i_MIPS/n539 , \i_MIPS/n538 , \i_MIPS/n537 , \i_MIPS/n536 ,
         \i_MIPS/n535 , \i_MIPS/n534 , \i_MIPS/n533 , \i_MIPS/n532 ,
         \i_MIPS/n531 , \i_MIPS/n530 , \i_MIPS/n529 , \i_MIPS/n528 ,
         \i_MIPS/n527 , \i_MIPS/n526 , \i_MIPS/n525 , \i_MIPS/n524 ,
         \i_MIPS/n523 , \i_MIPS/n522 , \i_MIPS/n521 , \i_MIPS/n520 ,
         \i_MIPS/n519 , \i_MIPS/n518 , \i_MIPS/n517 , \i_MIPS/n516 ,
         \i_MIPS/n515 , \i_MIPS/n514 , \i_MIPS/n513 , \i_MIPS/n512 ,
         \i_MIPS/n511 , \i_MIPS/n510 , \i_MIPS/n509 , \i_MIPS/n508 ,
         \i_MIPS/n507 , \i_MIPS/n506 , \i_MIPS/n505 , \i_MIPS/n504 ,
         \i_MIPS/n503 , \i_MIPS/n502 , \i_MIPS/n501 , \i_MIPS/n500 ,
         \i_MIPS/n499 , \i_MIPS/n498 , \i_MIPS/n497 , \i_MIPS/n496 ,
         \i_MIPS/n495 , \i_MIPS/n494 , \i_MIPS/n493 , \i_MIPS/n492 ,
         \i_MIPS/n491 , \i_MIPS/n490 , \i_MIPS/n489 , \i_MIPS/n488 ,
         \i_MIPS/n487 , \i_MIPS/n486 , \i_MIPS/n485 , \i_MIPS/n484 ,
         \i_MIPS/n483 , \i_MIPS/n482 , \i_MIPS/n481 , \i_MIPS/n480 ,
         \i_MIPS/n479 , \i_MIPS/n478 , \i_MIPS/n477 , \i_MIPS/n476 ,
         \i_MIPS/n475 , \i_MIPS/n474 , \i_MIPS/n473 , \i_MIPS/n472 ,
         \i_MIPS/n471 , \i_MIPS/n470 , \i_MIPS/n469 , \i_MIPS/n468 ,
         \i_MIPS/n467 , \i_MIPS/n466 , \i_MIPS/n465 , \i_MIPS/n464 ,
         \i_MIPS/n463 , \i_MIPS/n462 , \i_MIPS/n461 , \i_MIPS/n460 ,
         \i_MIPS/n459 , \i_MIPS/n458 , \i_MIPS/n457 , \i_MIPS/n456 ,
         \i_MIPS/n455 , \i_MIPS/n454 , \i_MIPS/n453 , \i_MIPS/n452 ,
         \i_MIPS/n451 , \i_MIPS/n450 , \i_MIPS/n449 , \i_MIPS/n448 ,
         \i_MIPS/n447 , \i_MIPS/n446 , \i_MIPS/n445 , \i_MIPS/n444 ,
         \i_MIPS/n443 , \i_MIPS/n442 , \i_MIPS/n441 , \i_MIPS/n440 ,
         \i_MIPS/n439 , \i_MIPS/n438 , \i_MIPS/n437 , \i_MIPS/n436 ,
         \i_MIPS/n435 , \i_MIPS/n434 , \i_MIPS/n433 , \i_MIPS/n432 ,
         \i_MIPS/n431 , \i_MIPS/n430 , \i_MIPS/n429 , \i_MIPS/n428 ,
         \i_MIPS/n427 , \i_MIPS/n426 , \i_MIPS/n425 , \i_MIPS/n424 ,
         \i_MIPS/n423 , \i_MIPS/n422 , \i_MIPS/n421 , \i_MIPS/n420 ,
         \i_MIPS/n419 , \i_MIPS/n418 , \i_MIPS/n417 , \i_MIPS/n416 ,
         \i_MIPS/n415 , \i_MIPS/n414 , \i_MIPS/n413 , \i_MIPS/n412 ,
         \i_MIPS/n411 , \i_MIPS/n410 , \i_MIPS/n409 , \i_MIPS/n408 ,
         \i_MIPS/n407 , \i_MIPS/n406 , \i_MIPS/n405 , \i_MIPS/n404 ,
         \i_MIPS/n403 , \i_MIPS/n402 , \i_MIPS/n401 , \i_MIPS/n400 ,
         \i_MIPS/n399 , \i_MIPS/n398 , \i_MIPS/n397 , \i_MIPS/n396 ,
         \i_MIPS/n395 , \i_MIPS/n394 , \i_MIPS/n393 , \i_MIPS/n392 ,
         \i_MIPS/n391 , \i_MIPS/n390 , \i_MIPS/n389 , \i_MIPS/n388 ,
         \i_MIPS/n387 , \i_MIPS/n386 , \i_MIPS/n385 , \i_MIPS/n384 ,
         \i_MIPS/n383 , \i_MIPS/n382 , \i_MIPS/n381 , \i_MIPS/n380 ,
         \i_MIPS/n379 , \i_MIPS/n378 , \i_MIPS/n377 , \i_MIPS/n376 ,
         \i_MIPS/n375 , \i_MIPS/n374 , \i_MIPS/n373 , \i_MIPS/n372 ,
         \i_MIPS/n371 , \i_MIPS/n370 , \i_MIPS/n369 , \i_MIPS/n368 ,
         \i_MIPS/n367 , \i_MIPS/n366 , \i_MIPS/n365 , \i_MIPS/n364 ,
         \i_MIPS/n363 , \i_MIPS/n362 , \i_MIPS/n361 , \i_MIPS/n360 ,
         \i_MIPS/n359 , \i_MIPS/n358 , \i_MIPS/n356 , \i_MIPS/n355 ,
         \i_MIPS/n354 , \i_MIPS/n353 , \i_MIPS/n352 , \i_MIPS/n351 ,
         \i_MIPS/n350 , \i_MIPS/n349 , \i_MIPS/n348 , \i_MIPS/n347 ,
         \i_MIPS/n346 , \i_MIPS/n345 , \i_MIPS/n344 , \i_MIPS/n343 ,
         \i_MIPS/n342 , \i_MIPS/n341 , \i_MIPS/n340 , \i_MIPS/n339 ,
         \i_MIPS/n338 , \i_MIPS/n337 , \i_MIPS/n336 , \i_MIPS/n335 ,
         \i_MIPS/n334 , \i_MIPS/n333 , \i_MIPS/n332 , \i_MIPS/n331 ,
         \i_MIPS/n330 , \i_MIPS/n329 , \i_MIPS/n328 , \i_MIPS/n327 ,
         \i_MIPS/n326 , \i_MIPS/n325 , \i_MIPS/n324 , \i_MIPS/n323 ,
         \i_MIPS/n322 , \i_MIPS/n321 , \i_MIPS/n320 , \i_MIPS/n319 ,
         \i_MIPS/n318 , \i_MIPS/n317 , \i_MIPS/n316 , \i_MIPS/n315 ,
         \i_MIPS/n314 , \i_MIPS/n313 , \i_MIPS/n312 , \i_MIPS/n311 ,
         \i_MIPS/n310 , \i_MIPS/n309 , \i_MIPS/n308 , \i_MIPS/n307 ,
         \i_MIPS/n306 , \i_MIPS/n305 , \i_MIPS/n304 , \i_MIPS/n303 ,
         \i_MIPS/n302 , \i_MIPS/n301 , \i_MIPS/n300 , \i_MIPS/n299 ,
         \i_MIPS/n298 , \i_MIPS/n296 , \i_MIPS/n295 , \i_MIPS/n294 ,
         \i_MIPS/n293 , \i_MIPS/n292 , \i_MIPS/n291 , \i_MIPS/n290 ,
         \i_MIPS/n289 , \i_MIPS/n288 , \i_MIPS/n287 , \i_MIPS/n286 ,
         \i_MIPS/n285 , \i_MIPS/n284 , \i_MIPS/n283 , \i_MIPS/n282 ,
         \i_MIPS/n281 , \i_MIPS/n280 , \i_MIPS/n279 , \i_MIPS/n278 ,
         \i_MIPS/n277 , \i_MIPS/n276 , \i_MIPS/n275 , \i_MIPS/n274 ,
         \i_MIPS/n273 , \i_MIPS/n272 , \i_MIPS/n271 , \i_MIPS/n270 ,
         \i_MIPS/n269 , \i_MIPS/n268 , \i_MIPS/n267 , \i_MIPS/n266 ,
         \i_MIPS/n265 , \i_MIPS/n264 , \i_MIPS/n263 , \i_MIPS/n262 ,
         \i_MIPS/n261 , \i_MIPS/n260 , \i_MIPS/n259 , \i_MIPS/n258 ,
         \i_MIPS/n257 , \i_MIPS/n256 , \i_MIPS/n255 , \i_MIPS/n254 ,
         \i_MIPS/n253 , \i_MIPS/n252 , \i_MIPS/n251 , \i_MIPS/n250 ,
         \i_MIPS/n249 , \i_MIPS/n248 , \i_MIPS/n247 , \i_MIPS/n246 ,
         \i_MIPS/n245 , \i_MIPS/n244 , \i_MIPS/n243 , \i_MIPS/n242 ,
         \i_MIPS/n241 , \i_MIPS/n240 , \i_MIPS/n239 , \i_MIPS/n238 ,
         \i_MIPS/n237 , \i_MIPS/n236 , \i_MIPS/n235 , \i_MIPS/n234 ,
         \i_MIPS/n233 , \i_MIPS/n232 , \i_MIPS/n231 , \i_MIPS/n230 ,
         \i_MIPS/n229 , \i_MIPS/n228 , \i_MIPS/n227 , \i_MIPS/n226 ,
         \i_MIPS/n225 , \i_MIPS/n224 , \i_MIPS/n223 , \i_MIPS/n222 ,
         \i_MIPS/n221 , \i_MIPS/n220 , \i_MIPS/n219 , \i_MIPS/n218 ,
         \i_MIPS/n217 , \i_MIPS/n216 , \i_MIPS/n215 , \i_MIPS/n214 ,
         \i_MIPS/n213 , \i_MIPS/n212 , \i_MIPS/n211 , \i_MIPS/n210 ,
         \i_MIPS/n209 , \i_MIPS/n208 , \i_MIPS/n207 , \i_MIPS/n206 ,
         \i_MIPS/n205 , \i_MIPS/n204 , \i_MIPS/n203 , \i_MIPS/n202 ,
         \i_MIPS/n201 , \i_MIPS/n200 , \i_MIPS/n199 , \i_MIPS/n198 ,
         \i_MIPS/n197 , \i_MIPS/n196 , \i_MIPS/n195 , \i_MIPS/n194 ,
         \i_MIPS/n193 , \i_MIPS/n192 , \i_MIPS/n191 , \i_MIPS/n190 ,
         \i_MIPS/n189 , \i_MIPS/n188 , \i_MIPS/n187 , \i_MIPS/n186 ,
         \i_MIPS/n185 , \i_MIPS/n184 , \i_MIPS/n183 , \i_MIPS/n182 ,
         \i_MIPS/n181 , \i_MIPS/n180 , \i_MIPS/n179 , \i_MIPS/n178 ,
         \i_MIPS/n177 , \i_MIPS/n176 , \i_MIPS/n175 , \i_MIPS/n174 ,
         \i_MIPS/n173 , \i_MIPS/n172 , \i_MIPS/n171 , \i_MIPS/n170 ,
         \i_MIPS/n169 , \i_MIPS/n168 , \i_MIPS/n167 , \i_MIPS/n166 ,
         \i_MIPS/n165 , \i_MIPS/n164 , \i_MIPS/n163 , \i_MIPS/n162 ,
         \i_MIPS/n161 , \i_MIPS/n160 , \i_MIPS/n159 , \i_MIPS/N120 ,
         \i_MIPS/N119 , \i_MIPS/N118 , \i_MIPS/N117 , \i_MIPS/N116 ,
         \i_MIPS/N115 , \i_MIPS/N114 , \i_MIPS/N113 , \i_MIPS/N112 ,
         \i_MIPS/N111 , \i_MIPS/N110 , \i_MIPS/N109 , \i_MIPS/N108 ,
         \i_MIPS/N107 , \i_MIPS/N106 , \i_MIPS/N105 , \i_MIPS/N104 ,
         \i_MIPS/N103 , \i_MIPS/N102 , \i_MIPS/N101 , \i_MIPS/N100 ,
         \i_MIPS/N99 , \i_MIPS/N98 , \i_MIPS/N97 , \i_MIPS/N96 , \i_MIPS/N95 ,
         \i_MIPS/N94 , \i_MIPS/N93 , \i_MIPS/N92 , \i_MIPS/N91 , \i_MIPS/N90 ,
         \i_MIPS/N89 , \i_MIPS/N88 , \i_MIPS/N87 , \i_MIPS/N86 , \i_MIPS/N85 ,
         \i_MIPS/N84 , \i_MIPS/N83 , \i_MIPS/N82 , \i_MIPS/N81 , \i_MIPS/N80 ,
         \i_MIPS/N79 , \i_MIPS/N78 , \i_MIPS/N77 , \i_MIPS/N76 , \i_MIPS/N75 ,
         \i_MIPS/N74 , \i_MIPS/N73 , \i_MIPS/N72 , \i_MIPS/N71 , \i_MIPS/N70 ,
         \i_MIPS/N69 , \i_MIPS/N68 , \i_MIPS/N67 , \i_MIPS/N66 , \i_MIPS/N65 ,
         \i_MIPS/N64 , \i_MIPS/N63 , \i_MIPS/N62 , \i_MIPS/N61 , \i_MIPS/N60 ,
         \i_MIPS/N59 , \i_MIPS/N58 , \i_MIPS/N57 , \i_MIPS/N56 , \i_MIPS/N55 ,
         \i_MIPS/N54 , \i_MIPS/N53 , \i_MIPS/N52 , \i_MIPS/N51 , \i_MIPS/N50 ,
         \i_MIPS/N49 , \i_MIPS/N48 , \i_MIPS/N47 , \i_MIPS/N46 , \i_MIPS/N45 ,
         \i_MIPS/N44 , \i_MIPS/N43 , \i_MIPS/N42 , \i_MIPS/N41 , \i_MIPS/N40 ,
         \i_MIPS/N39 , \i_MIPS/N38 , \i_MIPS/N37 , \i_MIPS/N36 , \i_MIPS/N35 ,
         \i_MIPS/N34 , \i_MIPS/N33 , \i_MIPS/N32 , \i_MIPS/N31 , \i_MIPS/N30 ,
         \i_MIPS/N29 , \i_MIPS/N28 , \i_MIPS/N27 , \i_MIPS/N26 , \i_MIPS/N25 ,
         \i_MIPS/N24 , \i_MIPS/N23 , \i_MIPS/ALUin1[30] , \i_MIPS/ALUin1[29] ,
         \i_MIPS/ALUin1[28] , \i_MIPS/ALUin1[27] , \i_MIPS/ALUin1[26] ,
         \i_MIPS/ALUin1[25] , \i_MIPS/ALUin1[24] , \i_MIPS/ALUin1[23] ,
         \i_MIPS/ALUin1[22] , \i_MIPS/ALUin1[21] , \i_MIPS/ALUin1[20] ,
         \i_MIPS/ALUin1[19] , \i_MIPS/ALUin1[18] , \i_MIPS/ALUin1[17] ,
         \i_MIPS/ALUin1[16] , \i_MIPS/ALUin1[15] , \i_MIPS/ALUin1[13] ,
         \i_MIPS/ALUin1[12] , \i_MIPS/ALUin1[11] , \i_MIPS/ALUin1[10] ,
         \i_MIPS/ALUin1[9] , \i_MIPS/ALUin1[8] , \i_MIPS/ALUin1[7] ,
         \i_MIPS/ALUin1[6] , \i_MIPS/ALUin1[5] , \i_MIPS/ALUin1[4] ,
         \i_MIPS/ALUin1[3] , \i_MIPS/ALUin1[2] , \i_MIPS/ALUin1[1] ,
         \i_MIPS/ALUin1[0] , \i_MIPS/ALUOp[1] , \i_MIPS/EX_MEM_0 ,
         \i_MIPS/EX_MEM_1 , \i_MIPS/EX_MEM[5] , \i_MIPS/EX_MEM[6] ,
         \i_MIPS/EX_MEM_74 , \i_MIPS/Sign_Extend_ID[31] ,
         \i_MIPS/Sign_Extend_ID[8] , \i_MIPS/Sign_Extend_ID[6] ,
         \i_MIPS/Sign_Extend_ID[5] , \i_MIPS/Sign_Extend_ID[4] ,
         \i_MIPS/Sign_Extend_ID[3] , \i_MIPS/Sign_Extend_ID[2] ,
         \i_MIPS/Sign_Extend_ID[1] , \i_MIPS/Sign_Extend_ID[0] ,
         \i_MIPS/ID_EX_0 , \i_MIPS/ID_EX_3 , \i_MIPS/ID_EX_5 ,
         \i_MIPS/ID_EX[41] , \i_MIPS/ID_EX[49] , \i_MIPS/ID_EX[50] ,
         \i_MIPS/ID_EX[55] , \i_MIPS/ID_EX[56] , \i_MIPS/ID_EX[68] ,
         \i_MIPS/ID_EX[69] , \i_MIPS/ID_EX[70] , \i_MIPS/ID_EX[72] ,
         \i_MIPS/ID_EX[73] , \i_MIPS/ID_EX[75] , \i_MIPS/ID_EX[78] ,
         \i_MIPS/ID_EX[80] , \i_MIPS/ID_EX[81] , \i_MIPS/ID_EX[82] ,
         \i_MIPS/ID_EX[83] , \i_MIPS/ID_EX[84] , \i_MIPS/ID_EX[85] ,
         \i_MIPS/ID_EX[86] , \i_MIPS/ID_EX[87] , \i_MIPS/ID_EX[88] ,
         \i_MIPS/ID_EX[89] , \i_MIPS/ID_EX[90] , \i_MIPS/ID_EX[91] ,
         \i_MIPS/ID_EX[92] , \i_MIPS/ID_EX[93] , \i_MIPS/ID_EX[94] ,
         \i_MIPS/ID_EX[95] , \i_MIPS/ID_EX[96] , \i_MIPS/ID_EX[97] ,
         \i_MIPS/ID_EX[98] , \i_MIPS/ID_EX[99] , \i_MIPS/ID_EX[100] ,
         \i_MIPS/ID_EX[101] , \i_MIPS/ID_EX[102] , \i_MIPS/ID_EX[103] ,
         \i_MIPS/ID_EX[104] , \i_MIPS/ID_EX[105] , \i_MIPS/ID_EX[106] ,
         \i_MIPS/ID_EX[107] , \i_MIPS/ID_EX[108] , \i_MIPS/ID_EX[111] ,
         \i_MIPS/ID_EX[112] , \i_MIPS/ID_EX[113] , \i_MIPS/ID_EX[114] ,
         \i_MIPS/ID_EX[115] , \i_MIPS/control_out[7] , \i_MIPS/control_out[0] ,
         \i_MIPS/Reg_W[0] , \i_MIPS/Reg_W[1] , \i_MIPS/Reg_W[2] ,
         \i_MIPS/Reg_W[3] , \i_MIPS/Reg_W[4] , \i_MIPS/IR_ID[16] ,
         \i_MIPS/IR_ID[17] , \i_MIPS/IR_ID[18] , \i_MIPS/IR_ID[19] ,
         \i_MIPS/IR_ID[20] , \i_MIPS/IR_ID[21] , \i_MIPS/IR_ID[22] ,
         \i_MIPS/IR_ID[23] , \i_MIPS/IR_ID[24] , \i_MIPS/IR_ID[25] ,
         \i_MIPS/IR_ID[26] , \i_MIPS/IR_ID[27] , \i_MIPS/IR_ID[28] ,
         \i_MIPS/IR_ID[29] , \i_MIPS/IR_ID[30] , \i_MIPS/IR_ID[31] ,
         \i_MIPS/PC_o[1] , \i_MIPS/IF_ID_1 , \i_MIPS/IF_ID_2 ,
         \i_MIPS/IF_ID_28 , \i_MIPS/IF_ID[64] , \i_MIPS/IF_ID[65] ,
         \i_MIPS/IF_ID[66] , \i_MIPS/IF_ID[67] , \i_MIPS/IF_ID[68] ,
         \i_MIPS/IF_ID[69] , \i_MIPS/IF_ID[70] , \i_MIPS/IF_ID[71] ,
         \i_MIPS/IF_ID[72] , \i_MIPS/IF_ID[73] , \i_MIPS/IF_ID[74] ,
         \i_MIPS/IF_ID[75] , \i_MIPS/IF_ID[76] , \i_MIPS/IF_ID[77] ,
         \i_MIPS/IF_ID[78] , \i_MIPS/IF_ID[79] , \i_MIPS/IF_ID[80] ,
         \i_MIPS/IF_ID[81] , \i_MIPS/IF_ID[82] , \i_MIPS/IF_ID[83] ,
         \i_MIPS/IF_ID[84] , \i_MIPS/IF_ID[85] , \i_MIPS/IF_ID[86] ,
         \i_MIPS/IF_ID[87] , \i_MIPS/IF_ID[88] , \i_MIPS/IF_ID[89] ,
         \i_MIPS/IF_ID[90] , \i_MIPS/IF_ID[91] , \i_MIPS/IF_ID[92] ,
         \i_MIPS/IF_ID[93] , \i_MIPS/IF_ID[94] , \i_MIPS/IF_ID[95] ,
         \i_MIPS/IF_ID[96] , \i_MIPS/IF_ID[97] , \i_MIPS/BranchAddr[0] ,
         \D_cache/n1796 , \D_cache/n1795 , \D_cache/n1794 , \D_cache/n1793 ,
         \D_cache/n1792 , \D_cache/n1791 , \D_cache/n1790 , \D_cache/n1789 ,
         \D_cache/n1788 , \D_cache/n1787 , \D_cache/n1786 , \D_cache/n1785 ,
         \D_cache/n1784 , \D_cache/n1783 , \D_cache/n1782 , \D_cache/n1781 ,
         \D_cache/n1780 , \D_cache/n1779 , \D_cache/n1778 , \D_cache/n1777 ,
         \D_cache/n1776 , \D_cache/n1775 , \D_cache/n1774 , \D_cache/n1773 ,
         \D_cache/n1772 , \D_cache/n1771 , \D_cache/n1770 , \D_cache/n1769 ,
         \D_cache/n1768 , \D_cache/n1767 , \D_cache/n1766 , \D_cache/n1765 ,
         \D_cache/n1764 , \D_cache/n1763 , \D_cache/n1762 , \D_cache/n1761 ,
         \D_cache/n1760 , \D_cache/n1759 , \D_cache/n1758 , \D_cache/n1757 ,
         \D_cache/n1756 , \D_cache/n1755 , \D_cache/n1754 , \D_cache/n1753 ,
         \D_cache/n1752 , \D_cache/n1751 , \D_cache/n1750 , \D_cache/n1749 ,
         \D_cache/n1748 , \D_cache/n1747 , \D_cache/n1746 , \D_cache/n1745 ,
         \D_cache/n1744 , \D_cache/n1743 , \D_cache/n1742 , \D_cache/n1741 ,
         \D_cache/n1740 , \D_cache/n1739 , \D_cache/n1738 , \D_cache/n1737 ,
         \D_cache/n1736 , \D_cache/n1735 , \D_cache/n1734 , \D_cache/n1733 ,
         \D_cache/n1732 , \D_cache/n1731 , \D_cache/n1730 , \D_cache/n1729 ,
         \D_cache/n1728 , \D_cache/n1727 , \D_cache/n1726 , \D_cache/n1725 ,
         \D_cache/n1724 , \D_cache/n1723 , \D_cache/n1722 , \D_cache/n1721 ,
         \D_cache/n1720 , \D_cache/n1719 , \D_cache/n1718 , \D_cache/n1717 ,
         \D_cache/n1716 , \D_cache/n1715 , \D_cache/n1714 , \D_cache/n1713 ,
         \D_cache/n1712 , \D_cache/n1711 , \D_cache/n1710 , \D_cache/n1709 ,
         \D_cache/n1708 , \D_cache/n1707 , \D_cache/n1706 , \D_cache/n1705 ,
         \D_cache/n1704 , \D_cache/n1703 , \D_cache/n1702 , \D_cache/n1701 ,
         \D_cache/n1700 , \D_cache/n1699 , \D_cache/n1698 , \D_cache/n1697 ,
         \D_cache/n1696 , \D_cache/n1695 , \D_cache/n1694 , \D_cache/n1693 ,
         \D_cache/n1692 , \D_cache/n1691 , \D_cache/n1690 , \D_cache/n1689 ,
         \D_cache/n1688 , \D_cache/n1687 , \D_cache/n1686 , \D_cache/n1685 ,
         \D_cache/n1684 , \D_cache/n1683 , \D_cache/n1682 , \D_cache/n1681 ,
         \D_cache/n1680 , \D_cache/n1679 , \D_cache/n1678 , \D_cache/n1677 ,
         \D_cache/n1676 , \D_cache/n1675 , \D_cache/n1674 , \D_cache/n1673 ,
         \D_cache/n1672 , \D_cache/n1671 , \D_cache/n1670 , \D_cache/n1669 ,
         \D_cache/n1668 , \D_cache/n1667 , \D_cache/n1666 , \D_cache/n1665 ,
         \D_cache/n1664 , \D_cache/n1663 , \D_cache/n1662 , \D_cache/n1661 ,
         \D_cache/n1660 , \D_cache/n1659 , \D_cache/n1658 , \D_cache/n1657 ,
         \D_cache/n1656 , \D_cache/n1655 , \D_cache/n1654 , \D_cache/n1653 ,
         \D_cache/n1652 , \D_cache/n1651 , \D_cache/n1650 , \D_cache/n1649 ,
         \D_cache/n1648 , \D_cache/n1647 , \D_cache/n1646 , \D_cache/n1645 ,
         \D_cache/n1644 , \D_cache/n1643 , \D_cache/n1642 , \D_cache/n1641 ,
         \D_cache/n1640 , \D_cache/n1639 , \D_cache/n1638 , \D_cache/n1637 ,
         \D_cache/n1636 , \D_cache/n1635 , \D_cache/n1634 , \D_cache/n1633 ,
         \D_cache/n1632 , \D_cache/n1631 , \D_cache/n1630 , \D_cache/n1629 ,
         \D_cache/n1628 , \D_cache/n1627 , \D_cache/n1626 , \D_cache/n1625 ,
         \D_cache/n1624 , \D_cache/n1623 , \D_cache/n1622 , \D_cache/n1621 ,
         \D_cache/n1620 , \D_cache/n1619 , \D_cache/n1618 , \D_cache/n1617 ,
         \D_cache/n1616 , \D_cache/n1615 , \D_cache/n1614 , \D_cache/n1613 ,
         \D_cache/n1612 , \D_cache/n1611 , \D_cache/n1610 , \D_cache/n1609 ,
         \D_cache/n1608 , \D_cache/n1607 , \D_cache/n1606 , \D_cache/n1605 ,
         \D_cache/n1604 , \D_cache/n1603 , \D_cache/n1602 , \D_cache/n1601 ,
         \D_cache/n1600 , \D_cache/n1599 , \D_cache/n1598 , \D_cache/n1597 ,
         \D_cache/n1596 , \D_cache/n1595 , \D_cache/n1594 , \D_cache/n1593 ,
         \D_cache/n1592 , \D_cache/n1591 , \D_cache/n1590 , \D_cache/n1589 ,
         \D_cache/n1588 , \D_cache/n1587 , \D_cache/n1586 , \D_cache/n1585 ,
         \D_cache/n1584 , \D_cache/n1583 , \D_cache/n1582 , \D_cache/n1581 ,
         \D_cache/n1580 , \D_cache/n1579 , \D_cache/n1578 , \D_cache/n1577 ,
         \D_cache/n1576 , \D_cache/n1575 , \D_cache/n1574 , \D_cache/n1573 ,
         \D_cache/n1572 , \D_cache/n1571 , \D_cache/n1570 , \D_cache/n1569 ,
         \D_cache/n1568 , \D_cache/n1567 , \D_cache/n1566 , \D_cache/n1565 ,
         \D_cache/n1564 , \D_cache/n1563 , \D_cache/n1562 , \D_cache/n1561 ,
         \D_cache/n1560 , \D_cache/n1559 , \D_cache/n1558 , \D_cache/n1557 ,
         \D_cache/n1556 , \D_cache/n1555 , \D_cache/n1554 , \D_cache/n1553 ,
         \D_cache/n1552 , \D_cache/n1551 , \D_cache/n1550 , \D_cache/n1549 ,
         \D_cache/n1548 , \D_cache/n1547 , \D_cache/n1546 , \D_cache/n1545 ,
         \D_cache/n1544 , \D_cache/n1543 , \D_cache/n1542 , \D_cache/n1541 ,
         \D_cache/n1540 , \D_cache/n1539 , \D_cache/n1538 , \D_cache/n1537 ,
         \D_cache/n1536 , \D_cache/n1535 , \D_cache/n1534 , \D_cache/n1533 ,
         \D_cache/n1532 , \D_cache/n1531 , \D_cache/n1530 , \D_cache/n1529 ,
         \D_cache/n1528 , \D_cache/n1527 , \D_cache/n1526 , \D_cache/n1525 ,
         \D_cache/n1524 , \D_cache/n1523 , \D_cache/n1522 , \D_cache/n1521 ,
         \D_cache/n1520 , \D_cache/n1519 , \D_cache/n1518 , \D_cache/n1517 ,
         \D_cache/n1516 , \D_cache/n1515 , \D_cache/n1514 , \D_cache/n1513 ,
         \D_cache/n1512 , \D_cache/n1511 , \D_cache/n1510 , \D_cache/n1509 ,
         \D_cache/n1508 , \D_cache/n1507 , \D_cache/n1506 , \D_cache/n1505 ,
         \D_cache/n1504 , \D_cache/n1503 , \D_cache/n1502 , \D_cache/n1501 ,
         \D_cache/n1500 , \D_cache/n1499 , \D_cache/n1498 , \D_cache/n1497 ,
         \D_cache/n1496 , \D_cache/n1495 , \D_cache/n1494 , \D_cache/n1493 ,
         \D_cache/n1492 , \D_cache/n1491 , \D_cache/n1490 , \D_cache/n1489 ,
         \D_cache/n1488 , \D_cache/n1487 , \D_cache/n1486 , \D_cache/n1485 ,
         \D_cache/n1484 , \D_cache/n1483 , \D_cache/n1482 , \D_cache/n1481 ,
         \D_cache/n1480 , \D_cache/n1479 , \D_cache/n1478 , \D_cache/n1477 ,
         \D_cache/n1476 , \D_cache/n1475 , \D_cache/n1474 , \D_cache/n1473 ,
         \D_cache/n1472 , \D_cache/n1471 , \D_cache/n1470 , \D_cache/n1469 ,
         \D_cache/n1468 , \D_cache/n1467 , \D_cache/n1466 , \D_cache/n1465 ,
         \D_cache/n1464 , \D_cache/n1463 , \D_cache/n1462 , \D_cache/n1461 ,
         \D_cache/n1460 , \D_cache/n1459 , \D_cache/n1458 , \D_cache/n1457 ,
         \D_cache/n1456 , \D_cache/n1455 , \D_cache/n1454 , \D_cache/n1453 ,
         \D_cache/n1452 , \D_cache/n1451 , \D_cache/n1450 , \D_cache/n1449 ,
         \D_cache/n1448 , \D_cache/n1447 , \D_cache/n1446 , \D_cache/n1445 ,
         \D_cache/n1444 , \D_cache/n1443 , \D_cache/n1442 , \D_cache/n1441 ,
         \D_cache/n1440 , \D_cache/n1439 , \D_cache/n1438 , \D_cache/n1437 ,
         \D_cache/n1436 , \D_cache/n1435 , \D_cache/n1434 , \D_cache/n1433 ,
         \D_cache/n1432 , \D_cache/n1431 , \D_cache/n1430 , \D_cache/n1429 ,
         \D_cache/n1428 , \D_cache/n1427 , \D_cache/n1426 , \D_cache/n1425 ,
         \D_cache/n1424 , \D_cache/n1423 , \D_cache/n1422 , \D_cache/n1421 ,
         \D_cache/n1420 , \D_cache/n1419 , \D_cache/n1418 , \D_cache/n1417 ,
         \D_cache/n1416 , \D_cache/n1415 , \D_cache/n1414 , \D_cache/n1413 ,
         \D_cache/n1412 , \D_cache/n1411 , \D_cache/n1410 , \D_cache/n1409 ,
         \D_cache/n1408 , \D_cache/n1407 , \D_cache/n1406 , \D_cache/n1405 ,
         \D_cache/n1404 , \D_cache/n1403 , \D_cache/n1402 , \D_cache/n1401 ,
         \D_cache/n1400 , \D_cache/n1399 , \D_cache/n1398 , \D_cache/n1397 ,
         \D_cache/n1396 , \D_cache/n1395 , \D_cache/n1394 , \D_cache/n1393 ,
         \D_cache/n1392 , \D_cache/n1391 , \D_cache/n1390 , \D_cache/n1389 ,
         \D_cache/n1388 , \D_cache/n1387 , \D_cache/n1386 , \D_cache/n1385 ,
         \D_cache/n1384 , \D_cache/n1383 , \D_cache/n1382 , \D_cache/n1381 ,
         \D_cache/n1380 , \D_cache/n1379 , \D_cache/n1378 , \D_cache/n1377 ,
         \D_cache/n1376 , \D_cache/n1375 , \D_cache/n1374 , \D_cache/n1373 ,
         \D_cache/n1372 , \D_cache/n1371 , \D_cache/n1370 , \D_cache/n1369 ,
         \D_cache/n1368 , \D_cache/n1367 , \D_cache/n1366 , \D_cache/n1365 ,
         \D_cache/n1364 , \D_cache/n1363 , \D_cache/n1362 , \D_cache/n1361 ,
         \D_cache/n1360 , \D_cache/n1359 , \D_cache/n1358 , \D_cache/n1357 ,
         \D_cache/n1356 , \D_cache/n1355 , \D_cache/n1354 , \D_cache/n1353 ,
         \D_cache/n1352 , \D_cache/n1351 , \D_cache/n1350 , \D_cache/n1349 ,
         \D_cache/n1348 , \D_cache/n1347 , \D_cache/n1346 , \D_cache/n1345 ,
         \D_cache/n1344 , \D_cache/n1343 , \D_cache/n1342 , \D_cache/n1341 ,
         \D_cache/n1340 , \D_cache/n1339 , \D_cache/n1338 , \D_cache/n1337 ,
         \D_cache/n1336 , \D_cache/n1335 , \D_cache/n1334 , \D_cache/n1333 ,
         \D_cache/n1332 , \D_cache/n1331 , \D_cache/n1330 , \D_cache/n1329 ,
         \D_cache/n1328 , \D_cache/n1327 , \D_cache/n1326 , \D_cache/n1325 ,
         \D_cache/n1324 , \D_cache/n1323 , \D_cache/n1322 , \D_cache/n1321 ,
         \D_cache/n1320 , \D_cache/n1319 , \D_cache/n1318 , \D_cache/n1317 ,
         \D_cache/n1316 , \D_cache/n1315 , \D_cache/n1314 , \D_cache/n1313 ,
         \D_cache/n1312 , \D_cache/n1311 , \D_cache/n1310 , \D_cache/n1309 ,
         \D_cache/n1308 , \D_cache/n1307 , \D_cache/n1306 , \D_cache/n1305 ,
         \D_cache/n1304 , \D_cache/n1303 , \D_cache/n1302 , \D_cache/n1301 ,
         \D_cache/n1300 , \D_cache/n1299 , \D_cache/n1298 , \D_cache/n1297 ,
         \D_cache/n1296 , \D_cache/n1295 , \D_cache/n1294 , \D_cache/n1293 ,
         \D_cache/n1292 , \D_cache/n1291 , \D_cache/n1290 , \D_cache/n1289 ,
         \D_cache/n1288 , \D_cache/n1287 , \D_cache/n1286 , \D_cache/n1285 ,
         \D_cache/n1284 , \D_cache/n1283 , \D_cache/n1282 , \D_cache/n1281 ,
         \D_cache/n1280 , \D_cache/n1279 , \D_cache/n1278 , \D_cache/n1277 ,
         \D_cache/n1276 , \D_cache/n1275 , \D_cache/n1274 , \D_cache/n1273 ,
         \D_cache/n1272 , \D_cache/n1271 , \D_cache/n1270 , \D_cache/n1269 ,
         \D_cache/n1268 , \D_cache/n1267 , \D_cache/n1266 , \D_cache/n1265 ,
         \D_cache/n1264 , \D_cache/n1263 , \D_cache/n1262 , \D_cache/n1261 ,
         \D_cache/n1260 , \D_cache/n1259 , \D_cache/n1258 , \D_cache/n1257 ,
         \D_cache/n1256 , \D_cache/n1255 , \D_cache/n1254 , \D_cache/n1253 ,
         \D_cache/n1252 , \D_cache/n1251 , \D_cache/n1250 , \D_cache/n1249 ,
         \D_cache/n1248 , \D_cache/n1247 , \D_cache/n1246 , \D_cache/n1245 ,
         \D_cache/n1244 , \D_cache/n1243 , \D_cache/n1242 , \D_cache/n1241 ,
         \D_cache/n1240 , \D_cache/n1239 , \D_cache/n1238 , \D_cache/n1237 ,
         \D_cache/n1236 , \D_cache/n1235 , \D_cache/n1234 , \D_cache/n1233 ,
         \D_cache/n1232 , \D_cache/n1231 , \D_cache/n1230 , \D_cache/n1229 ,
         \D_cache/n1228 , \D_cache/n1227 , \D_cache/n1226 , \D_cache/n1225 ,
         \D_cache/n1224 , \D_cache/n1223 , \D_cache/n1222 , \D_cache/n1221 ,
         \D_cache/n1220 , \D_cache/n1219 , \D_cache/n1218 , \D_cache/n1217 ,
         \D_cache/n1216 , \D_cache/n1215 , \D_cache/n1214 , \D_cache/n1213 ,
         \D_cache/n1212 , \D_cache/n1211 , \D_cache/n1210 , \D_cache/n1209 ,
         \D_cache/n1208 , \D_cache/n1207 , \D_cache/n1206 , \D_cache/n1205 ,
         \D_cache/n1204 , \D_cache/n1203 , \D_cache/n1202 , \D_cache/n1201 ,
         \D_cache/n1200 , \D_cache/n1199 , \D_cache/n1198 , \D_cache/n1197 ,
         \D_cache/n1196 , \D_cache/n1195 , \D_cache/n1194 , \D_cache/n1193 ,
         \D_cache/n1192 , \D_cache/n1191 , \D_cache/n1190 , \D_cache/n1189 ,
         \D_cache/n1188 , \D_cache/n1187 , \D_cache/n1186 , \D_cache/n1185 ,
         \D_cache/n1184 , \D_cache/n1183 , \D_cache/n1182 , \D_cache/n1181 ,
         \D_cache/n1180 , \D_cache/n1179 , \D_cache/n1178 , \D_cache/n1177 ,
         \D_cache/n1176 , \D_cache/n1175 , \D_cache/n1174 , \D_cache/n1173 ,
         \D_cache/n1172 , \D_cache/n1171 , \D_cache/n1170 , \D_cache/n1169 ,
         \D_cache/n1168 , \D_cache/n1167 , \D_cache/n1166 , \D_cache/n1165 ,
         \D_cache/n1164 , \D_cache/n1163 , \D_cache/n1162 , \D_cache/n1161 ,
         \D_cache/n1160 , \D_cache/n1159 , \D_cache/n1158 , \D_cache/n1157 ,
         \D_cache/n1156 , \D_cache/n1155 , \D_cache/n1154 , \D_cache/n1153 ,
         \D_cache/n1152 , \D_cache/n1151 , \D_cache/n1150 , \D_cache/n1149 ,
         \D_cache/n1148 , \D_cache/n1147 , \D_cache/n1146 , \D_cache/n1145 ,
         \D_cache/n1144 , \D_cache/n1143 , \D_cache/n1142 , \D_cache/n1141 ,
         \D_cache/n1140 , \D_cache/n1139 , \D_cache/n1138 , \D_cache/n1137 ,
         \D_cache/n1136 , \D_cache/n1135 , \D_cache/n1134 , \D_cache/n1133 ,
         \D_cache/n1132 , \D_cache/n1131 , \D_cache/n1130 , \D_cache/n1129 ,
         \D_cache/n1128 , \D_cache/n1127 , \D_cache/n1126 , \D_cache/n1125 ,
         \D_cache/n1124 , \D_cache/n1123 , \D_cache/n1122 , \D_cache/n1121 ,
         \D_cache/n1120 , \D_cache/n1119 , \D_cache/n1118 , \D_cache/n1117 ,
         \D_cache/n1116 , \D_cache/n1115 , \D_cache/n1114 , \D_cache/n1113 ,
         \D_cache/n1112 , \D_cache/n1111 , \D_cache/n1110 , \D_cache/n1109 ,
         \D_cache/n1108 , \D_cache/n1107 , \D_cache/n1106 , \D_cache/n1105 ,
         \D_cache/n1104 , \D_cache/n1103 , \D_cache/n1102 , \D_cache/n1101 ,
         \D_cache/n1100 , \D_cache/n1099 , \D_cache/n1098 , \D_cache/n1097 ,
         \D_cache/n1096 , \D_cache/n1095 , \D_cache/n1094 , \D_cache/n1093 ,
         \D_cache/n1092 , \D_cache/n1091 , \D_cache/n1090 , \D_cache/n1089 ,
         \D_cache/n1088 , \D_cache/n1087 , \D_cache/n1086 , \D_cache/n1085 ,
         \D_cache/n1084 , \D_cache/n1083 , \D_cache/n1082 , \D_cache/n1081 ,
         \D_cache/n1080 , \D_cache/n1079 , \D_cache/n1078 , \D_cache/n1077 ,
         \D_cache/n1076 , \D_cache/n1075 , \D_cache/n1074 , \D_cache/n1073 ,
         \D_cache/n1072 , \D_cache/n1071 , \D_cache/n1070 , \D_cache/n1069 ,
         \D_cache/n1068 , \D_cache/n1067 , \D_cache/n1066 , \D_cache/n1065 ,
         \D_cache/n1064 , \D_cache/n1063 , \D_cache/n1062 , \D_cache/n1061 ,
         \D_cache/n1060 , \D_cache/n1059 , \D_cache/n1058 , \D_cache/n1057 ,
         \D_cache/n1056 , \D_cache/n1055 , \D_cache/n1054 , \D_cache/n1053 ,
         \D_cache/n1052 , \D_cache/n1051 , \D_cache/n1050 , \D_cache/n1049 ,
         \D_cache/n1048 , \D_cache/n1047 , \D_cache/n1046 , \D_cache/n1045 ,
         \D_cache/n1044 , \D_cache/n1043 , \D_cache/n1042 , \D_cache/n1041 ,
         \D_cache/n1040 , \D_cache/n1039 , \D_cache/n1038 , \D_cache/n1037 ,
         \D_cache/n1036 , \D_cache/n1035 , \D_cache/n1034 , \D_cache/n1033 ,
         \D_cache/n1032 , \D_cache/n1031 , \D_cache/n1030 , \D_cache/n1029 ,
         \D_cache/n1028 , \D_cache/n1027 , \D_cache/n1026 , \D_cache/n1025 ,
         \D_cache/n1024 , \D_cache/n1023 , \D_cache/n1022 , \D_cache/n1021 ,
         \D_cache/n1020 , \D_cache/n1019 , \D_cache/n1018 , \D_cache/n1017 ,
         \D_cache/n1016 , \D_cache/n1015 , \D_cache/n1014 , \D_cache/n1013 ,
         \D_cache/n1012 , \D_cache/n1011 , \D_cache/n1010 , \D_cache/n1009 ,
         \D_cache/n1008 , \D_cache/n1007 , \D_cache/n1006 , \D_cache/n1005 ,
         \D_cache/n1004 , \D_cache/n1003 , \D_cache/n1002 , \D_cache/n1001 ,
         \D_cache/n1000 , \D_cache/n999 , \D_cache/n998 , \D_cache/n997 ,
         \D_cache/n996 , \D_cache/n995 , \D_cache/n994 , \D_cache/n993 ,
         \D_cache/n992 , \D_cache/n991 , \D_cache/n990 , \D_cache/n989 ,
         \D_cache/n988 , \D_cache/n987 , \D_cache/n986 , \D_cache/n985 ,
         \D_cache/n984 , \D_cache/n983 , \D_cache/n982 , \D_cache/n981 ,
         \D_cache/n980 , \D_cache/n979 , \D_cache/n978 , \D_cache/n977 ,
         \D_cache/n976 , \D_cache/n975 , \D_cache/n974 , \D_cache/n973 ,
         \D_cache/n972 , \D_cache/n971 , \D_cache/n970 , \D_cache/n969 ,
         \D_cache/n968 , \D_cache/n967 , \D_cache/n966 , \D_cache/n965 ,
         \D_cache/n964 , \D_cache/n963 , \D_cache/n962 , \D_cache/n961 ,
         \D_cache/n960 , \D_cache/n959 , \D_cache/n958 , \D_cache/n957 ,
         \D_cache/n956 , \D_cache/n955 , \D_cache/n954 , \D_cache/n953 ,
         \D_cache/n952 , \D_cache/n951 , \D_cache/n950 , \D_cache/n949 ,
         \D_cache/n948 , \D_cache/n947 , \D_cache/n946 , \D_cache/n945 ,
         \D_cache/n944 , \D_cache/n943 , \D_cache/n942 , \D_cache/n941 ,
         \D_cache/n940 , \D_cache/n939 , \D_cache/n938 , \D_cache/n937 ,
         \D_cache/n936 , \D_cache/n935 , \D_cache/n934 , \D_cache/n933 ,
         \D_cache/n932 , \D_cache/n931 , \D_cache/n930 , \D_cache/n929 ,
         \D_cache/n928 , \D_cache/n927 , \D_cache/n926 , \D_cache/n925 ,
         \D_cache/n924 , \D_cache/n923 , \D_cache/n922 , \D_cache/n921 ,
         \D_cache/n920 , \D_cache/n919 , \D_cache/n918 , \D_cache/n917 ,
         \D_cache/n916 , \D_cache/n915 , \D_cache/n914 , \D_cache/n913 ,
         \D_cache/n912 , \D_cache/n911 , \D_cache/n910 , \D_cache/n909 ,
         \D_cache/n908 , \D_cache/n907 , \D_cache/n906 , \D_cache/n905 ,
         \D_cache/n904 , \D_cache/n903 , \D_cache/n902 , \D_cache/n901 ,
         \D_cache/n900 , \D_cache/n899 , \D_cache/n898 , \D_cache/n897 ,
         \D_cache/n896 , \D_cache/n895 , \D_cache/n894 , \D_cache/n893 ,
         \D_cache/n892 , \D_cache/n891 , \D_cache/n890 , \D_cache/n889 ,
         \D_cache/n888 , \D_cache/n887 , \D_cache/n886 , \D_cache/n885 ,
         \D_cache/n884 , \D_cache/n883 , \D_cache/n882 , \D_cache/n881 ,
         \D_cache/n880 , \D_cache/n879 , \D_cache/n878 , \D_cache/n877 ,
         \D_cache/n876 , \D_cache/n875 , \D_cache/n874 , \D_cache/n873 ,
         \D_cache/n872 , \D_cache/n871 , \D_cache/n870 , \D_cache/n869 ,
         \D_cache/n868 , \D_cache/n867 , \D_cache/n866 , \D_cache/n865 ,
         \D_cache/n864 , \D_cache/n863 , \D_cache/n862 , \D_cache/n861 ,
         \D_cache/n860 , \D_cache/n859 , \D_cache/n858 , \D_cache/n857 ,
         \D_cache/n856 , \D_cache/n855 , \D_cache/n854 , \D_cache/n853 ,
         \D_cache/n852 , \D_cache/n851 , \D_cache/n850 , \D_cache/n849 ,
         \D_cache/n848 , \D_cache/n847 , \D_cache/n846 , \D_cache/n845 ,
         \D_cache/n844 , \D_cache/n843 , \D_cache/n842 , \D_cache/n841 ,
         \D_cache/n840 , \D_cache/n839 , \D_cache/n838 , \D_cache/n837 ,
         \D_cache/n836 , \D_cache/n835 , \D_cache/n834 , \D_cache/n833 ,
         \D_cache/n832 , \D_cache/n831 , \D_cache/n830 , \D_cache/n829 ,
         \D_cache/n828 , \D_cache/n827 , \D_cache/n826 , \D_cache/n825 ,
         \D_cache/n824 , \D_cache/n823 , \D_cache/n822 , \D_cache/n821 ,
         \D_cache/n820 , \D_cache/n819 , \D_cache/n818 , \D_cache/n817 ,
         \D_cache/n816 , \D_cache/n815 , \D_cache/n814 , \D_cache/n813 ,
         \D_cache/n812 , \D_cache/n811 , \D_cache/n810 , \D_cache/n809 ,
         \D_cache/n808 , \D_cache/n807 , \D_cache/n806 , \D_cache/n805 ,
         \D_cache/n804 , \D_cache/n803 , \D_cache/n802 , \D_cache/n801 ,
         \D_cache/n800 , \D_cache/n799 , \D_cache/n798 , \D_cache/n797 ,
         \D_cache/n796 , \D_cache/n795 , \D_cache/n794 , \D_cache/n793 ,
         \D_cache/n792 , \D_cache/n791 , \D_cache/n790 , \D_cache/n789 ,
         \D_cache/n788 , \D_cache/n787 , \D_cache/n786 , \D_cache/n785 ,
         \D_cache/n784 , \D_cache/n783 , \D_cache/n782 , \D_cache/n781 ,
         \D_cache/n780 , \D_cache/n779 , \D_cache/n778 , \D_cache/n777 ,
         \D_cache/n776 , \D_cache/n775 , \D_cache/n774 , \D_cache/n773 ,
         \D_cache/n772 , \D_cache/n771 , \D_cache/n770 , \D_cache/n769 ,
         \D_cache/n768 , \D_cache/n767 , \D_cache/n766 , \D_cache/n765 ,
         \D_cache/n764 , \D_cache/n763 , \D_cache/n762 , \D_cache/n761 ,
         \D_cache/n760 , \D_cache/n759 , \D_cache/n758 , \D_cache/n757 ,
         \D_cache/n756 , \D_cache/n755 , \D_cache/n754 , \D_cache/n753 ,
         \D_cache/n752 , \D_cache/n751 , \D_cache/n750 , \D_cache/n749 ,
         \D_cache/n748 , \D_cache/n747 , \D_cache/n746 , \D_cache/n745 ,
         \D_cache/n744 , \D_cache/n743 , \D_cache/n742 , \D_cache/n741 ,
         \D_cache/n740 , \D_cache/n739 , \D_cache/n738 , \D_cache/n737 ,
         \D_cache/n736 , \D_cache/n735 , \D_cache/n734 , \D_cache/n733 ,
         \D_cache/n732 , \D_cache/n731 , \D_cache/n730 , \D_cache/n729 ,
         \D_cache/n728 , \D_cache/n727 , \D_cache/n726 , \D_cache/n725 ,
         \D_cache/n724 , \D_cache/n723 , \D_cache/n722 , \D_cache/n721 ,
         \D_cache/n720 , \D_cache/n719 , \D_cache/n718 , \D_cache/n717 ,
         \D_cache/n716 , \D_cache/n715 , \D_cache/n714 , \D_cache/n713 ,
         \D_cache/n712 , \D_cache/n711 , \D_cache/n710 , \D_cache/n709 ,
         \D_cache/n708 , \D_cache/n707 , \D_cache/n706 , \D_cache/n705 ,
         \D_cache/n704 , \D_cache/n703 , \D_cache/n702 , \D_cache/n701 ,
         \D_cache/n700 , \D_cache/n699 , \D_cache/n698 , \D_cache/n697 ,
         \D_cache/n696 , \D_cache/n695 , \D_cache/n694 , \D_cache/n693 ,
         \D_cache/n692 , \D_cache/n691 , \D_cache/n690 , \D_cache/n689 ,
         \D_cache/n688 , \D_cache/n687 , \D_cache/n686 , \D_cache/n685 ,
         \D_cache/n684 , \D_cache/n683 , \D_cache/n682 , \D_cache/n681 ,
         \D_cache/n680 , \D_cache/n679 , \D_cache/n678 , \D_cache/n677 ,
         \D_cache/n676 , \D_cache/n675 , \D_cache/n674 , \D_cache/n673 ,
         \D_cache/n672 , \D_cache/n671 , \D_cache/n670 , \D_cache/n669 ,
         \D_cache/n668 , \D_cache/n667 , \D_cache/n666 , \D_cache/n665 ,
         \D_cache/n664 , \D_cache/n663 , \D_cache/n662 , \D_cache/n661 ,
         \D_cache/n660 , \D_cache/n659 , \D_cache/n658 , \D_cache/n657 ,
         \D_cache/n656 , \D_cache/n655 , \D_cache/n654 , \D_cache/n653 ,
         \D_cache/n652 , \D_cache/n651 , \D_cache/n650 , \D_cache/n649 ,
         \D_cache/n648 , \D_cache/n647 , \D_cache/n646 , \D_cache/n645 ,
         \D_cache/n644 , \D_cache/n643 , \D_cache/n642 , \D_cache/n641 ,
         \D_cache/n640 , \D_cache/n639 , \D_cache/n638 , \D_cache/n637 ,
         \D_cache/n636 , \D_cache/n635 , \D_cache/n634 , \D_cache/n633 ,
         \D_cache/n632 , \D_cache/n631 , \D_cache/n630 , \D_cache/n629 ,
         \D_cache/n628 , \D_cache/n627 , \D_cache/n626 , \D_cache/n625 ,
         \D_cache/n624 , \D_cache/n623 , \D_cache/n622 , \D_cache/n621 ,
         \D_cache/n620 , \D_cache/n619 , \D_cache/n618 , \D_cache/n617 ,
         \D_cache/n616 , \D_cache/n615 , \D_cache/n614 , \D_cache/n613 ,
         \D_cache/n612 , \D_cache/n611 , \D_cache/n610 , \D_cache/n609 ,
         \D_cache/n608 , \D_cache/n607 , \D_cache/n606 , \D_cache/n605 ,
         \D_cache/n604 , \D_cache/n603 , \D_cache/n602 , \D_cache/n601 ,
         \D_cache/n600 , \D_cache/n599 , \D_cache/n598 , \D_cache/n597 ,
         \D_cache/n596 , \D_cache/n595 , \D_cache/n594 , \D_cache/n593 ,
         \D_cache/n592 , \D_cache/n591 , \D_cache/n590 , \D_cache/n589 ,
         \D_cache/n588 , \D_cache/n587 , \D_cache/n586 , \D_cache/n585 ,
         \D_cache/n584 , \D_cache/n583 , \D_cache/n582 , \D_cache/n581 ,
         \D_cache/n580 , \D_cache/n579 , \D_cache/n578 , \D_cache/n577 ,
         \D_cache/n576 , \D_cache/n575 , \D_cache/n574 , \D_cache/n573 ,
         \D_cache/n572 , \D_cache/n571 , \D_cache/n570 , \D_cache/n569 ,
         \D_cache/n568 , \D_cache/n567 , \D_cache/n566 , \D_cache/n565 ,
         \D_cache/n564 , \D_cache/n563 , \D_cache/n562 , \D_cache/n561 ,
         \D_cache/n560 , \D_cache/n559 , \D_cache/n558 , \D_cache/n557 ,
         \D_cache/cache[7][0] , \D_cache/cache[7][1] , \D_cache/cache[7][2] ,
         \D_cache/cache[7][3] , \D_cache/cache[7][4] , \D_cache/cache[7][5] ,
         \D_cache/cache[7][6] , \D_cache/cache[7][7] , \D_cache/cache[7][8] ,
         \D_cache/cache[7][9] , \D_cache/cache[7][10] , \D_cache/cache[7][11] ,
         \D_cache/cache[7][12] , \D_cache/cache[7][13] ,
         \D_cache/cache[7][14] , \D_cache/cache[7][15] ,
         \D_cache/cache[7][16] , \D_cache/cache[7][17] ,
         \D_cache/cache[7][18] , \D_cache/cache[7][19] ,
         \D_cache/cache[7][20] , \D_cache/cache[7][21] ,
         \D_cache/cache[7][22] , \D_cache/cache[7][23] ,
         \D_cache/cache[7][24] , \D_cache/cache[7][25] ,
         \D_cache/cache[7][26] , \D_cache/cache[7][27] ,
         \D_cache/cache[7][28] , \D_cache/cache[7][29] ,
         \D_cache/cache[7][30] , \D_cache/cache[7][31] ,
         \D_cache/cache[7][32] , \D_cache/cache[7][33] ,
         \D_cache/cache[7][34] , \D_cache/cache[7][35] ,
         \D_cache/cache[7][36] , \D_cache/cache[7][37] ,
         \D_cache/cache[7][38] , \D_cache/cache[7][39] ,
         \D_cache/cache[7][40] , \D_cache/cache[7][41] ,
         \D_cache/cache[7][42] , \D_cache/cache[7][43] ,
         \D_cache/cache[7][44] , \D_cache/cache[7][45] ,
         \D_cache/cache[7][46] , \D_cache/cache[7][47] ,
         \D_cache/cache[7][48] , \D_cache/cache[7][49] ,
         \D_cache/cache[7][50] , \D_cache/cache[7][51] ,
         \D_cache/cache[7][52] , \D_cache/cache[7][53] ,
         \D_cache/cache[7][54] , \D_cache/cache[7][55] ,
         \D_cache/cache[7][56] , \D_cache/cache[7][57] ,
         \D_cache/cache[7][58] , \D_cache/cache[7][59] ,
         \D_cache/cache[7][60] , \D_cache/cache[7][61] ,
         \D_cache/cache[7][62] , \D_cache/cache[7][63] ,
         \D_cache/cache[7][64] , \D_cache/cache[7][65] ,
         \D_cache/cache[7][66] , \D_cache/cache[7][67] ,
         \D_cache/cache[7][68] , \D_cache/cache[7][69] ,
         \D_cache/cache[7][70] , \D_cache/cache[7][71] ,
         \D_cache/cache[7][72] , \D_cache/cache[7][73] ,
         \D_cache/cache[7][74] , \D_cache/cache[7][75] ,
         \D_cache/cache[7][76] , \D_cache/cache[7][77] ,
         \D_cache/cache[7][78] , \D_cache/cache[7][79] ,
         \D_cache/cache[7][80] , \D_cache/cache[7][81] ,
         \D_cache/cache[7][82] , \D_cache/cache[7][83] ,
         \D_cache/cache[7][84] , \D_cache/cache[7][85] ,
         \D_cache/cache[7][86] , \D_cache/cache[7][87] ,
         \D_cache/cache[7][88] , \D_cache/cache[7][89] ,
         \D_cache/cache[7][90] , \D_cache/cache[7][91] ,
         \D_cache/cache[7][92] , \D_cache/cache[7][93] ,
         \D_cache/cache[7][94] , \D_cache/cache[7][95] ,
         \D_cache/cache[7][96] , \D_cache/cache[7][97] ,
         \D_cache/cache[7][98] , \D_cache/cache[7][99] ,
         \D_cache/cache[7][100] , \D_cache/cache[7][101] ,
         \D_cache/cache[7][102] , \D_cache/cache[7][103] ,
         \D_cache/cache[7][104] , \D_cache/cache[7][105] ,
         \D_cache/cache[7][106] , \D_cache/cache[7][107] ,
         \D_cache/cache[7][108] , \D_cache/cache[7][109] ,
         \D_cache/cache[7][110] , \D_cache/cache[7][111] ,
         \D_cache/cache[7][112] , \D_cache/cache[7][113] ,
         \D_cache/cache[7][114] , \D_cache/cache[7][115] ,
         \D_cache/cache[7][116] , \D_cache/cache[7][117] ,
         \D_cache/cache[7][118] , \D_cache/cache[7][119] ,
         \D_cache/cache[7][120] , \D_cache/cache[7][121] ,
         \D_cache/cache[7][122] , \D_cache/cache[7][123] ,
         \D_cache/cache[7][124] , \D_cache/cache[7][125] ,
         \D_cache/cache[7][126] , \D_cache/cache[7][127] ,
         \D_cache/cache[7][128] , \D_cache/cache[7][129] ,
         \D_cache/cache[7][130] , \D_cache/cache[7][131] ,
         \D_cache/cache[7][132] , \D_cache/cache[7][133] ,
         \D_cache/cache[7][134] , \D_cache/cache[7][135] ,
         \D_cache/cache[7][136] , \D_cache/cache[7][137] ,
         \D_cache/cache[7][138] , \D_cache/cache[7][139] ,
         \D_cache/cache[7][140] , \D_cache/cache[7][141] ,
         \D_cache/cache[7][142] , \D_cache/cache[7][143] ,
         \D_cache/cache[7][144] , \D_cache/cache[7][145] ,
         \D_cache/cache[7][146] , \D_cache/cache[7][147] ,
         \D_cache/cache[7][148] , \D_cache/cache[7][149] ,
         \D_cache/cache[7][150] , \D_cache/cache[7][151] ,
         \D_cache/cache[7][152] , \D_cache/cache[7][153] ,
         \D_cache/cache[7][154] , \D_cache/cache[6][0] , \D_cache/cache[6][1] ,
         \D_cache/cache[6][2] , \D_cache/cache[6][3] , \D_cache/cache[6][4] ,
         \D_cache/cache[6][5] , \D_cache/cache[6][6] , \D_cache/cache[6][7] ,
         \D_cache/cache[6][8] , \D_cache/cache[6][9] , \D_cache/cache[6][10] ,
         \D_cache/cache[6][11] , \D_cache/cache[6][12] ,
         \D_cache/cache[6][13] , \D_cache/cache[6][14] ,
         \D_cache/cache[6][15] , \D_cache/cache[6][16] ,
         \D_cache/cache[6][17] , \D_cache/cache[6][18] ,
         \D_cache/cache[6][19] , \D_cache/cache[6][20] ,
         \D_cache/cache[6][21] , \D_cache/cache[6][22] ,
         \D_cache/cache[6][23] , \D_cache/cache[6][24] ,
         \D_cache/cache[6][25] , \D_cache/cache[6][26] ,
         \D_cache/cache[6][27] , \D_cache/cache[6][28] ,
         \D_cache/cache[6][29] , \D_cache/cache[6][30] ,
         \D_cache/cache[6][31] , \D_cache/cache[6][32] ,
         \D_cache/cache[6][33] , \D_cache/cache[6][34] ,
         \D_cache/cache[6][35] , \D_cache/cache[6][36] ,
         \D_cache/cache[6][37] , \D_cache/cache[6][38] ,
         \D_cache/cache[6][39] , \D_cache/cache[6][40] ,
         \D_cache/cache[6][41] , \D_cache/cache[6][42] ,
         \D_cache/cache[6][43] , \D_cache/cache[6][44] ,
         \D_cache/cache[6][45] , \D_cache/cache[6][46] ,
         \D_cache/cache[6][47] , \D_cache/cache[6][48] ,
         \D_cache/cache[6][49] , \D_cache/cache[6][50] ,
         \D_cache/cache[6][51] , \D_cache/cache[6][52] ,
         \D_cache/cache[6][53] , \D_cache/cache[6][54] ,
         \D_cache/cache[6][55] , \D_cache/cache[6][56] ,
         \D_cache/cache[6][57] , \D_cache/cache[6][58] ,
         \D_cache/cache[6][59] , \D_cache/cache[6][60] ,
         \D_cache/cache[6][61] , \D_cache/cache[6][62] ,
         \D_cache/cache[6][63] , \D_cache/cache[6][64] ,
         \D_cache/cache[6][65] , \D_cache/cache[6][66] ,
         \D_cache/cache[6][67] , \D_cache/cache[6][68] ,
         \D_cache/cache[6][69] , \D_cache/cache[6][70] ,
         \D_cache/cache[6][71] , \D_cache/cache[6][72] ,
         \D_cache/cache[6][73] , \D_cache/cache[6][74] ,
         \D_cache/cache[6][75] , \D_cache/cache[6][76] ,
         \D_cache/cache[6][77] , \D_cache/cache[6][78] ,
         \D_cache/cache[6][79] , \D_cache/cache[6][80] ,
         \D_cache/cache[6][81] , \D_cache/cache[6][82] ,
         \D_cache/cache[6][83] , \D_cache/cache[6][84] ,
         \D_cache/cache[6][85] , \D_cache/cache[6][86] ,
         \D_cache/cache[6][87] , \D_cache/cache[6][88] ,
         \D_cache/cache[6][89] , \D_cache/cache[6][90] ,
         \D_cache/cache[6][91] , \D_cache/cache[6][92] ,
         \D_cache/cache[6][93] , \D_cache/cache[6][94] ,
         \D_cache/cache[6][95] , \D_cache/cache[6][96] ,
         \D_cache/cache[6][97] , \D_cache/cache[6][98] ,
         \D_cache/cache[6][99] , \D_cache/cache[6][100] ,
         \D_cache/cache[6][101] , \D_cache/cache[6][102] ,
         \D_cache/cache[6][103] , \D_cache/cache[6][104] ,
         \D_cache/cache[6][105] , \D_cache/cache[6][106] ,
         \D_cache/cache[6][107] , \D_cache/cache[6][108] ,
         \D_cache/cache[6][109] , \D_cache/cache[6][110] ,
         \D_cache/cache[6][111] , \D_cache/cache[6][112] ,
         \D_cache/cache[6][113] , \D_cache/cache[6][114] ,
         \D_cache/cache[6][115] , \D_cache/cache[6][116] ,
         \D_cache/cache[6][117] , \D_cache/cache[6][118] ,
         \D_cache/cache[6][119] , \D_cache/cache[6][120] ,
         \D_cache/cache[6][121] , \D_cache/cache[6][122] ,
         \D_cache/cache[6][123] , \D_cache/cache[6][124] ,
         \D_cache/cache[6][125] , \D_cache/cache[6][126] ,
         \D_cache/cache[6][127] , \D_cache/cache[6][128] ,
         \D_cache/cache[6][129] , \D_cache/cache[6][130] ,
         \D_cache/cache[6][131] , \D_cache/cache[6][132] ,
         \D_cache/cache[6][133] , \D_cache/cache[6][134] ,
         \D_cache/cache[6][135] , \D_cache/cache[6][136] ,
         \D_cache/cache[6][137] , \D_cache/cache[6][138] ,
         \D_cache/cache[6][139] , \D_cache/cache[6][140] ,
         \D_cache/cache[6][141] , \D_cache/cache[6][142] ,
         \D_cache/cache[6][143] , \D_cache/cache[6][144] ,
         \D_cache/cache[6][145] , \D_cache/cache[6][146] ,
         \D_cache/cache[6][147] , \D_cache/cache[6][148] ,
         \D_cache/cache[6][149] , \D_cache/cache[6][150] ,
         \D_cache/cache[6][151] , \D_cache/cache[6][152] ,
         \D_cache/cache[6][153] , \D_cache/cache[6][154] ,
         \D_cache/cache[5][0] , \D_cache/cache[5][1] , \D_cache/cache[5][2] ,
         \D_cache/cache[5][3] , \D_cache/cache[5][4] , \D_cache/cache[5][5] ,
         \D_cache/cache[5][6] , \D_cache/cache[5][7] , \D_cache/cache[5][8] ,
         \D_cache/cache[5][9] , \D_cache/cache[5][10] , \D_cache/cache[5][11] ,
         \D_cache/cache[5][12] , \D_cache/cache[5][13] ,
         \D_cache/cache[5][14] , \D_cache/cache[5][15] ,
         \D_cache/cache[5][16] , \D_cache/cache[5][17] ,
         \D_cache/cache[5][18] , \D_cache/cache[5][19] ,
         \D_cache/cache[5][20] , \D_cache/cache[5][21] ,
         \D_cache/cache[5][22] , \D_cache/cache[5][23] ,
         \D_cache/cache[5][24] , \D_cache/cache[5][25] ,
         \D_cache/cache[5][26] , \D_cache/cache[5][27] ,
         \D_cache/cache[5][28] , \D_cache/cache[5][29] ,
         \D_cache/cache[5][30] , \D_cache/cache[5][31] ,
         \D_cache/cache[5][32] , \D_cache/cache[5][33] ,
         \D_cache/cache[5][34] , \D_cache/cache[5][35] ,
         \D_cache/cache[5][36] , \D_cache/cache[5][37] ,
         \D_cache/cache[5][38] , \D_cache/cache[5][39] ,
         \D_cache/cache[5][40] , \D_cache/cache[5][41] ,
         \D_cache/cache[5][42] , \D_cache/cache[5][43] ,
         \D_cache/cache[5][44] , \D_cache/cache[5][45] ,
         \D_cache/cache[5][46] , \D_cache/cache[5][47] ,
         \D_cache/cache[5][48] , \D_cache/cache[5][49] ,
         \D_cache/cache[5][50] , \D_cache/cache[5][51] ,
         \D_cache/cache[5][52] , \D_cache/cache[5][53] ,
         \D_cache/cache[5][54] , \D_cache/cache[5][55] ,
         \D_cache/cache[5][56] , \D_cache/cache[5][57] ,
         \D_cache/cache[5][58] , \D_cache/cache[5][59] ,
         \D_cache/cache[5][60] , \D_cache/cache[5][61] ,
         \D_cache/cache[5][62] , \D_cache/cache[5][63] ,
         \D_cache/cache[5][64] , \D_cache/cache[5][65] ,
         \D_cache/cache[5][66] , \D_cache/cache[5][67] ,
         \D_cache/cache[5][68] , \D_cache/cache[5][69] ,
         \D_cache/cache[5][70] , \D_cache/cache[5][71] ,
         \D_cache/cache[5][72] , \D_cache/cache[5][73] ,
         \D_cache/cache[5][74] , \D_cache/cache[5][75] ,
         \D_cache/cache[5][76] , \D_cache/cache[5][77] ,
         \D_cache/cache[5][78] , \D_cache/cache[5][79] ,
         \D_cache/cache[5][80] , \D_cache/cache[5][81] ,
         \D_cache/cache[5][82] , \D_cache/cache[5][83] ,
         \D_cache/cache[5][84] , \D_cache/cache[5][85] ,
         \D_cache/cache[5][86] , \D_cache/cache[5][87] ,
         \D_cache/cache[5][88] , \D_cache/cache[5][89] ,
         \D_cache/cache[5][90] , \D_cache/cache[5][91] ,
         \D_cache/cache[5][92] , \D_cache/cache[5][93] ,
         \D_cache/cache[5][94] , \D_cache/cache[5][95] ,
         \D_cache/cache[5][96] , \D_cache/cache[5][97] ,
         \D_cache/cache[5][98] , \D_cache/cache[5][99] ,
         \D_cache/cache[5][100] , \D_cache/cache[5][101] ,
         \D_cache/cache[5][102] , \D_cache/cache[5][103] ,
         \D_cache/cache[5][104] , \D_cache/cache[5][105] ,
         \D_cache/cache[5][106] , \D_cache/cache[5][107] ,
         \D_cache/cache[5][108] , \D_cache/cache[5][109] ,
         \D_cache/cache[5][110] , \D_cache/cache[5][111] ,
         \D_cache/cache[5][112] , \D_cache/cache[5][113] ,
         \D_cache/cache[5][114] , \D_cache/cache[5][115] ,
         \D_cache/cache[5][116] , \D_cache/cache[5][117] ,
         \D_cache/cache[5][118] , \D_cache/cache[5][119] ,
         \D_cache/cache[5][120] , \D_cache/cache[5][121] ,
         \D_cache/cache[5][122] , \D_cache/cache[5][123] ,
         \D_cache/cache[5][124] , \D_cache/cache[5][125] ,
         \D_cache/cache[5][126] , \D_cache/cache[5][127] ,
         \D_cache/cache[5][128] , \D_cache/cache[5][129] ,
         \D_cache/cache[5][130] , \D_cache/cache[5][131] ,
         \D_cache/cache[5][132] , \D_cache/cache[5][133] ,
         \D_cache/cache[5][134] , \D_cache/cache[5][135] ,
         \D_cache/cache[5][136] , \D_cache/cache[5][137] ,
         \D_cache/cache[5][138] , \D_cache/cache[5][139] ,
         \D_cache/cache[5][140] , \D_cache/cache[5][141] ,
         \D_cache/cache[5][142] , \D_cache/cache[5][143] ,
         \D_cache/cache[5][144] , \D_cache/cache[5][145] ,
         \D_cache/cache[5][146] , \D_cache/cache[5][147] ,
         \D_cache/cache[5][148] , \D_cache/cache[5][149] ,
         \D_cache/cache[5][150] , \D_cache/cache[5][151] ,
         \D_cache/cache[5][152] , \D_cache/cache[5][153] ,
         \D_cache/cache[5][154] , \D_cache/cache[4][0] , \D_cache/cache[4][1] ,
         \D_cache/cache[4][2] , \D_cache/cache[4][3] , \D_cache/cache[4][4] ,
         \D_cache/cache[4][5] , \D_cache/cache[4][6] , \D_cache/cache[4][7] ,
         \D_cache/cache[4][8] , \D_cache/cache[4][9] , \D_cache/cache[4][10] ,
         \D_cache/cache[4][11] , \D_cache/cache[4][12] ,
         \D_cache/cache[4][13] , \D_cache/cache[4][14] ,
         \D_cache/cache[4][15] , \D_cache/cache[4][16] ,
         \D_cache/cache[4][17] , \D_cache/cache[4][18] ,
         \D_cache/cache[4][19] , \D_cache/cache[4][20] ,
         \D_cache/cache[4][21] , \D_cache/cache[4][22] ,
         \D_cache/cache[4][23] , \D_cache/cache[4][24] ,
         \D_cache/cache[4][25] , \D_cache/cache[4][26] ,
         \D_cache/cache[4][27] , \D_cache/cache[4][28] ,
         \D_cache/cache[4][29] , \D_cache/cache[4][30] ,
         \D_cache/cache[4][31] , \D_cache/cache[4][32] ,
         \D_cache/cache[4][33] , \D_cache/cache[4][34] ,
         \D_cache/cache[4][35] , \D_cache/cache[4][36] ,
         \D_cache/cache[4][37] , \D_cache/cache[4][38] ,
         \D_cache/cache[4][39] , \D_cache/cache[4][40] ,
         \D_cache/cache[4][41] , \D_cache/cache[4][42] ,
         \D_cache/cache[4][43] , \D_cache/cache[4][44] ,
         \D_cache/cache[4][45] , \D_cache/cache[4][46] ,
         \D_cache/cache[4][47] , \D_cache/cache[4][48] ,
         \D_cache/cache[4][49] , \D_cache/cache[4][50] ,
         \D_cache/cache[4][51] , \D_cache/cache[4][52] ,
         \D_cache/cache[4][53] , \D_cache/cache[4][54] ,
         \D_cache/cache[4][55] , \D_cache/cache[4][56] ,
         \D_cache/cache[4][57] , \D_cache/cache[4][58] ,
         \D_cache/cache[4][59] , \D_cache/cache[4][60] ,
         \D_cache/cache[4][61] , \D_cache/cache[4][62] ,
         \D_cache/cache[4][63] , \D_cache/cache[4][64] ,
         \D_cache/cache[4][65] , \D_cache/cache[4][66] ,
         \D_cache/cache[4][67] , \D_cache/cache[4][68] ,
         \D_cache/cache[4][69] , \D_cache/cache[4][70] ,
         \D_cache/cache[4][71] , \D_cache/cache[4][72] ,
         \D_cache/cache[4][73] , \D_cache/cache[4][74] ,
         \D_cache/cache[4][75] , \D_cache/cache[4][76] ,
         \D_cache/cache[4][77] , \D_cache/cache[4][78] ,
         \D_cache/cache[4][79] , \D_cache/cache[4][80] ,
         \D_cache/cache[4][81] , \D_cache/cache[4][82] ,
         \D_cache/cache[4][83] , \D_cache/cache[4][84] ,
         \D_cache/cache[4][85] , \D_cache/cache[4][86] ,
         \D_cache/cache[4][87] , \D_cache/cache[4][88] ,
         \D_cache/cache[4][89] , \D_cache/cache[4][90] ,
         \D_cache/cache[4][91] , \D_cache/cache[4][92] ,
         \D_cache/cache[4][93] , \D_cache/cache[4][94] ,
         \D_cache/cache[4][95] , \D_cache/cache[4][96] ,
         \D_cache/cache[4][97] , \D_cache/cache[4][98] ,
         \D_cache/cache[4][99] , \D_cache/cache[4][100] ,
         \D_cache/cache[4][101] , \D_cache/cache[4][102] ,
         \D_cache/cache[4][103] , \D_cache/cache[4][104] ,
         \D_cache/cache[4][105] , \D_cache/cache[4][106] ,
         \D_cache/cache[4][107] , \D_cache/cache[4][108] ,
         \D_cache/cache[4][109] , \D_cache/cache[4][110] ,
         \D_cache/cache[4][111] , \D_cache/cache[4][112] ,
         \D_cache/cache[4][113] , \D_cache/cache[4][114] ,
         \D_cache/cache[4][115] , \D_cache/cache[4][116] ,
         \D_cache/cache[4][117] , \D_cache/cache[4][118] ,
         \D_cache/cache[4][119] , \D_cache/cache[4][120] ,
         \D_cache/cache[4][121] , \D_cache/cache[4][122] ,
         \D_cache/cache[4][123] , \D_cache/cache[4][124] ,
         \D_cache/cache[4][125] , \D_cache/cache[4][126] ,
         \D_cache/cache[4][127] , \D_cache/cache[4][128] ,
         \D_cache/cache[4][129] , \D_cache/cache[4][130] ,
         \D_cache/cache[4][131] , \D_cache/cache[4][132] ,
         \D_cache/cache[4][133] , \D_cache/cache[4][134] ,
         \D_cache/cache[4][135] , \D_cache/cache[4][136] ,
         \D_cache/cache[4][137] , \D_cache/cache[4][138] ,
         \D_cache/cache[4][139] , \D_cache/cache[4][140] ,
         \D_cache/cache[4][141] , \D_cache/cache[4][142] ,
         \D_cache/cache[4][143] , \D_cache/cache[4][144] ,
         \D_cache/cache[4][145] , \D_cache/cache[4][146] ,
         \D_cache/cache[4][147] , \D_cache/cache[4][148] ,
         \D_cache/cache[4][149] , \D_cache/cache[4][150] ,
         \D_cache/cache[4][151] , \D_cache/cache[4][152] ,
         \D_cache/cache[4][153] , \D_cache/cache[4][154] ,
         \D_cache/cache[3][0] , \D_cache/cache[3][1] , \D_cache/cache[3][2] ,
         \D_cache/cache[3][3] , \D_cache/cache[3][4] , \D_cache/cache[3][5] ,
         \D_cache/cache[3][6] , \D_cache/cache[3][7] , \D_cache/cache[3][8] ,
         \D_cache/cache[3][9] , \D_cache/cache[3][10] , \D_cache/cache[3][11] ,
         \D_cache/cache[3][12] , \D_cache/cache[3][13] ,
         \D_cache/cache[3][14] , \D_cache/cache[3][15] ,
         \D_cache/cache[3][16] , \D_cache/cache[3][17] ,
         \D_cache/cache[3][18] , \D_cache/cache[3][19] ,
         \D_cache/cache[3][20] , \D_cache/cache[3][21] ,
         \D_cache/cache[3][22] , \D_cache/cache[3][23] ,
         \D_cache/cache[3][24] , \D_cache/cache[3][25] ,
         \D_cache/cache[3][26] , \D_cache/cache[3][27] ,
         \D_cache/cache[3][28] , \D_cache/cache[3][29] ,
         \D_cache/cache[3][30] , \D_cache/cache[3][31] ,
         \D_cache/cache[3][32] , \D_cache/cache[3][33] ,
         \D_cache/cache[3][34] , \D_cache/cache[3][35] ,
         \D_cache/cache[3][36] , \D_cache/cache[3][37] ,
         \D_cache/cache[3][38] , \D_cache/cache[3][39] ,
         \D_cache/cache[3][40] , \D_cache/cache[3][41] ,
         \D_cache/cache[3][42] , \D_cache/cache[3][43] ,
         \D_cache/cache[3][44] , \D_cache/cache[3][45] ,
         \D_cache/cache[3][46] , \D_cache/cache[3][47] ,
         \D_cache/cache[3][48] , \D_cache/cache[3][49] ,
         \D_cache/cache[3][50] , \D_cache/cache[3][51] ,
         \D_cache/cache[3][52] , \D_cache/cache[3][53] ,
         \D_cache/cache[3][54] , \D_cache/cache[3][55] ,
         \D_cache/cache[3][56] , \D_cache/cache[3][57] ,
         \D_cache/cache[3][58] , \D_cache/cache[3][59] ,
         \D_cache/cache[3][60] , \D_cache/cache[3][61] ,
         \D_cache/cache[3][62] , \D_cache/cache[3][63] ,
         \D_cache/cache[3][64] , \D_cache/cache[3][65] ,
         \D_cache/cache[3][66] , \D_cache/cache[3][67] ,
         \D_cache/cache[3][68] , \D_cache/cache[3][69] ,
         \D_cache/cache[3][70] , \D_cache/cache[3][71] ,
         \D_cache/cache[3][72] , \D_cache/cache[3][73] ,
         \D_cache/cache[3][74] , \D_cache/cache[3][75] ,
         \D_cache/cache[3][76] , \D_cache/cache[3][77] ,
         \D_cache/cache[3][78] , \D_cache/cache[3][79] ,
         \D_cache/cache[3][80] , \D_cache/cache[3][81] ,
         \D_cache/cache[3][82] , \D_cache/cache[3][83] ,
         \D_cache/cache[3][84] , \D_cache/cache[3][85] ,
         \D_cache/cache[3][86] , \D_cache/cache[3][87] ,
         \D_cache/cache[3][88] , \D_cache/cache[3][89] ,
         \D_cache/cache[3][90] , \D_cache/cache[3][91] ,
         \D_cache/cache[3][92] , \D_cache/cache[3][93] ,
         \D_cache/cache[3][94] , \D_cache/cache[3][95] ,
         \D_cache/cache[3][96] , \D_cache/cache[3][97] ,
         \D_cache/cache[3][98] , \D_cache/cache[3][99] ,
         \D_cache/cache[3][100] , \D_cache/cache[3][101] ,
         \D_cache/cache[3][102] , \D_cache/cache[3][103] ,
         \D_cache/cache[3][104] , \D_cache/cache[3][105] ,
         \D_cache/cache[3][106] , \D_cache/cache[3][107] ,
         \D_cache/cache[3][108] , \D_cache/cache[3][109] ,
         \D_cache/cache[3][110] , \D_cache/cache[3][111] ,
         \D_cache/cache[3][112] , \D_cache/cache[3][113] ,
         \D_cache/cache[3][114] , \D_cache/cache[3][115] ,
         \D_cache/cache[3][116] , \D_cache/cache[3][117] ,
         \D_cache/cache[3][118] , \D_cache/cache[3][119] ,
         \D_cache/cache[3][120] , \D_cache/cache[3][121] ,
         \D_cache/cache[3][122] , \D_cache/cache[3][123] ,
         \D_cache/cache[3][124] , \D_cache/cache[3][125] ,
         \D_cache/cache[3][126] , \D_cache/cache[3][127] ,
         \D_cache/cache[3][128] , \D_cache/cache[3][129] ,
         \D_cache/cache[3][130] , \D_cache/cache[3][131] ,
         \D_cache/cache[3][132] , \D_cache/cache[3][133] ,
         \D_cache/cache[3][134] , \D_cache/cache[3][135] ,
         \D_cache/cache[3][136] , \D_cache/cache[3][137] ,
         \D_cache/cache[3][138] , \D_cache/cache[3][139] ,
         \D_cache/cache[3][140] , \D_cache/cache[3][141] ,
         \D_cache/cache[3][142] , \D_cache/cache[3][143] ,
         \D_cache/cache[3][144] , \D_cache/cache[3][145] ,
         \D_cache/cache[3][146] , \D_cache/cache[3][147] ,
         \D_cache/cache[3][148] , \D_cache/cache[3][149] ,
         \D_cache/cache[3][150] , \D_cache/cache[3][151] ,
         \D_cache/cache[3][152] , \D_cache/cache[3][153] ,
         \D_cache/cache[3][154] , \D_cache/cache[2][0] , \D_cache/cache[2][1] ,
         \D_cache/cache[2][2] , \D_cache/cache[2][3] , \D_cache/cache[2][4] ,
         \D_cache/cache[2][5] , \D_cache/cache[2][6] , \D_cache/cache[2][7] ,
         \D_cache/cache[2][8] , \D_cache/cache[2][9] , \D_cache/cache[2][10] ,
         \D_cache/cache[2][11] , \D_cache/cache[2][12] ,
         \D_cache/cache[2][13] , \D_cache/cache[2][14] ,
         \D_cache/cache[2][15] , \D_cache/cache[2][16] ,
         \D_cache/cache[2][17] , \D_cache/cache[2][18] ,
         \D_cache/cache[2][19] , \D_cache/cache[2][20] ,
         \D_cache/cache[2][21] , \D_cache/cache[2][22] ,
         \D_cache/cache[2][23] , \D_cache/cache[2][24] ,
         \D_cache/cache[2][25] , \D_cache/cache[2][26] ,
         \D_cache/cache[2][27] , \D_cache/cache[2][28] ,
         \D_cache/cache[2][29] , \D_cache/cache[2][30] ,
         \D_cache/cache[2][31] , \D_cache/cache[2][32] ,
         \D_cache/cache[2][33] , \D_cache/cache[2][34] ,
         \D_cache/cache[2][35] , \D_cache/cache[2][36] ,
         \D_cache/cache[2][37] , \D_cache/cache[2][38] ,
         \D_cache/cache[2][39] , \D_cache/cache[2][40] ,
         \D_cache/cache[2][41] , \D_cache/cache[2][42] ,
         \D_cache/cache[2][43] , \D_cache/cache[2][44] ,
         \D_cache/cache[2][45] , \D_cache/cache[2][46] ,
         \D_cache/cache[2][47] , \D_cache/cache[2][48] ,
         \D_cache/cache[2][49] , \D_cache/cache[2][50] ,
         \D_cache/cache[2][51] , \D_cache/cache[2][52] ,
         \D_cache/cache[2][53] , \D_cache/cache[2][54] ,
         \D_cache/cache[2][55] , \D_cache/cache[2][56] ,
         \D_cache/cache[2][57] , \D_cache/cache[2][58] ,
         \D_cache/cache[2][59] , \D_cache/cache[2][60] ,
         \D_cache/cache[2][61] , \D_cache/cache[2][62] ,
         \D_cache/cache[2][63] , \D_cache/cache[2][64] ,
         \D_cache/cache[2][65] , \D_cache/cache[2][66] ,
         \D_cache/cache[2][67] , \D_cache/cache[2][68] ,
         \D_cache/cache[2][69] , \D_cache/cache[2][70] ,
         \D_cache/cache[2][71] , \D_cache/cache[2][72] ,
         \D_cache/cache[2][73] , \D_cache/cache[2][74] ,
         \D_cache/cache[2][75] , \D_cache/cache[2][76] ,
         \D_cache/cache[2][77] , \D_cache/cache[2][78] ,
         \D_cache/cache[2][79] , \D_cache/cache[2][80] ,
         \D_cache/cache[2][81] , \D_cache/cache[2][82] ,
         \D_cache/cache[2][83] , \D_cache/cache[2][84] ,
         \D_cache/cache[2][85] , \D_cache/cache[2][86] ,
         \D_cache/cache[2][87] , \D_cache/cache[2][88] ,
         \D_cache/cache[2][89] , \D_cache/cache[2][90] ,
         \D_cache/cache[2][91] , \D_cache/cache[2][92] ,
         \D_cache/cache[2][93] , \D_cache/cache[2][94] ,
         \D_cache/cache[2][95] , \D_cache/cache[2][96] ,
         \D_cache/cache[2][97] , \D_cache/cache[2][98] ,
         \D_cache/cache[2][99] , \D_cache/cache[2][100] ,
         \D_cache/cache[2][101] , \D_cache/cache[2][102] ,
         \D_cache/cache[2][103] , \D_cache/cache[2][104] ,
         \D_cache/cache[2][105] , \D_cache/cache[2][106] ,
         \D_cache/cache[2][107] , \D_cache/cache[2][108] ,
         \D_cache/cache[2][109] , \D_cache/cache[2][110] ,
         \D_cache/cache[2][111] , \D_cache/cache[2][112] ,
         \D_cache/cache[2][113] , \D_cache/cache[2][114] ,
         \D_cache/cache[2][115] , \D_cache/cache[2][116] ,
         \D_cache/cache[2][117] , \D_cache/cache[2][118] ,
         \D_cache/cache[2][119] , \D_cache/cache[2][120] ,
         \D_cache/cache[2][121] , \D_cache/cache[2][122] ,
         \D_cache/cache[2][123] , \D_cache/cache[2][124] ,
         \D_cache/cache[2][125] , \D_cache/cache[2][126] ,
         \D_cache/cache[2][127] , \D_cache/cache[2][128] ,
         \D_cache/cache[2][129] , \D_cache/cache[2][130] ,
         \D_cache/cache[2][131] , \D_cache/cache[2][132] ,
         \D_cache/cache[2][133] , \D_cache/cache[2][134] ,
         \D_cache/cache[2][135] , \D_cache/cache[2][136] ,
         \D_cache/cache[2][137] , \D_cache/cache[2][138] ,
         \D_cache/cache[2][139] , \D_cache/cache[2][140] ,
         \D_cache/cache[2][141] , \D_cache/cache[2][142] ,
         \D_cache/cache[2][143] , \D_cache/cache[2][144] ,
         \D_cache/cache[2][145] , \D_cache/cache[2][146] ,
         \D_cache/cache[2][147] , \D_cache/cache[2][148] ,
         \D_cache/cache[2][149] , \D_cache/cache[2][150] ,
         \D_cache/cache[2][151] , \D_cache/cache[2][152] ,
         \D_cache/cache[2][153] , \D_cache/cache[2][154] ,
         \D_cache/cache[1][0] , \D_cache/cache[1][1] , \D_cache/cache[1][2] ,
         \D_cache/cache[1][3] , \D_cache/cache[1][4] , \D_cache/cache[1][5] ,
         \D_cache/cache[1][6] , \D_cache/cache[1][7] , \D_cache/cache[1][8] ,
         \D_cache/cache[1][9] , \D_cache/cache[1][10] , \D_cache/cache[1][11] ,
         \D_cache/cache[1][12] , \D_cache/cache[1][13] ,
         \D_cache/cache[1][14] , \D_cache/cache[1][15] ,
         \D_cache/cache[1][16] , \D_cache/cache[1][17] ,
         \D_cache/cache[1][18] , \D_cache/cache[1][19] ,
         \D_cache/cache[1][20] , \D_cache/cache[1][21] ,
         \D_cache/cache[1][22] , \D_cache/cache[1][23] ,
         \D_cache/cache[1][24] , \D_cache/cache[1][25] ,
         \D_cache/cache[1][26] , \D_cache/cache[1][27] ,
         \D_cache/cache[1][28] , \D_cache/cache[1][29] ,
         \D_cache/cache[1][30] , \D_cache/cache[1][31] ,
         \D_cache/cache[1][32] , \D_cache/cache[1][33] ,
         \D_cache/cache[1][34] , \D_cache/cache[1][35] ,
         \D_cache/cache[1][36] , \D_cache/cache[1][37] ,
         \D_cache/cache[1][38] , \D_cache/cache[1][39] ,
         \D_cache/cache[1][40] , \D_cache/cache[1][41] ,
         \D_cache/cache[1][42] , \D_cache/cache[1][43] ,
         \D_cache/cache[1][44] , \D_cache/cache[1][45] ,
         \D_cache/cache[1][46] , \D_cache/cache[1][47] ,
         \D_cache/cache[1][48] , \D_cache/cache[1][49] ,
         \D_cache/cache[1][50] , \D_cache/cache[1][51] ,
         \D_cache/cache[1][52] , \D_cache/cache[1][53] ,
         \D_cache/cache[1][54] , \D_cache/cache[1][55] ,
         \D_cache/cache[1][56] , \D_cache/cache[1][57] ,
         \D_cache/cache[1][58] , \D_cache/cache[1][59] ,
         \D_cache/cache[1][60] , \D_cache/cache[1][61] ,
         \D_cache/cache[1][62] , \D_cache/cache[1][63] ,
         \D_cache/cache[1][64] , \D_cache/cache[1][65] ,
         \D_cache/cache[1][66] , \D_cache/cache[1][67] ,
         \D_cache/cache[1][68] , \D_cache/cache[1][69] ,
         \D_cache/cache[1][70] , \D_cache/cache[1][71] ,
         \D_cache/cache[1][72] , \D_cache/cache[1][73] ,
         \D_cache/cache[1][74] , \D_cache/cache[1][75] ,
         \D_cache/cache[1][76] , \D_cache/cache[1][77] ,
         \D_cache/cache[1][78] , \D_cache/cache[1][79] ,
         \D_cache/cache[1][80] , \D_cache/cache[1][81] ,
         \D_cache/cache[1][82] , \D_cache/cache[1][83] ,
         \D_cache/cache[1][84] , \D_cache/cache[1][85] ,
         \D_cache/cache[1][86] , \D_cache/cache[1][87] ,
         \D_cache/cache[1][88] , \D_cache/cache[1][89] ,
         \D_cache/cache[1][90] , \D_cache/cache[1][91] ,
         \D_cache/cache[1][92] , \D_cache/cache[1][93] ,
         \D_cache/cache[1][94] , \D_cache/cache[1][95] ,
         \D_cache/cache[1][96] , \D_cache/cache[1][97] ,
         \D_cache/cache[1][98] , \D_cache/cache[1][99] ,
         \D_cache/cache[1][100] , \D_cache/cache[1][101] ,
         \D_cache/cache[1][102] , \D_cache/cache[1][103] ,
         \D_cache/cache[1][104] , \D_cache/cache[1][105] ,
         \D_cache/cache[1][106] , \D_cache/cache[1][107] ,
         \D_cache/cache[1][108] , \D_cache/cache[1][109] ,
         \D_cache/cache[1][110] , \D_cache/cache[1][111] ,
         \D_cache/cache[1][112] , \D_cache/cache[1][113] ,
         \D_cache/cache[1][114] , \D_cache/cache[1][115] ,
         \D_cache/cache[1][116] , \D_cache/cache[1][117] ,
         \D_cache/cache[1][118] , \D_cache/cache[1][119] ,
         \D_cache/cache[1][120] , \D_cache/cache[1][121] ,
         \D_cache/cache[1][122] , \D_cache/cache[1][123] ,
         \D_cache/cache[1][124] , \D_cache/cache[1][125] ,
         \D_cache/cache[1][126] , \D_cache/cache[1][127] ,
         \D_cache/cache[1][128] , \D_cache/cache[1][129] ,
         \D_cache/cache[1][130] , \D_cache/cache[1][131] ,
         \D_cache/cache[1][132] , \D_cache/cache[1][133] ,
         \D_cache/cache[1][134] , \D_cache/cache[1][135] ,
         \D_cache/cache[1][136] , \D_cache/cache[1][137] ,
         \D_cache/cache[1][138] , \D_cache/cache[1][139] ,
         \D_cache/cache[1][140] , \D_cache/cache[1][141] ,
         \D_cache/cache[1][142] , \D_cache/cache[1][143] ,
         \D_cache/cache[1][144] , \D_cache/cache[1][145] ,
         \D_cache/cache[1][146] , \D_cache/cache[1][147] ,
         \D_cache/cache[1][148] , \D_cache/cache[1][149] ,
         \D_cache/cache[1][150] , \D_cache/cache[1][151] ,
         \D_cache/cache[1][152] , \D_cache/cache[1][153] ,
         \D_cache/cache[1][154] , \D_cache/cache[0][0] , \D_cache/cache[0][1] ,
         \D_cache/cache[0][2] , \D_cache/cache[0][3] , \D_cache/cache[0][4] ,
         \D_cache/cache[0][5] , \D_cache/cache[0][6] , \D_cache/cache[0][7] ,
         \D_cache/cache[0][8] , \D_cache/cache[0][9] , \D_cache/cache[0][10] ,
         \D_cache/cache[0][11] , \D_cache/cache[0][12] ,
         \D_cache/cache[0][13] , \D_cache/cache[0][14] ,
         \D_cache/cache[0][15] , \D_cache/cache[0][16] ,
         \D_cache/cache[0][17] , \D_cache/cache[0][18] ,
         \D_cache/cache[0][19] , \D_cache/cache[0][20] ,
         \D_cache/cache[0][21] , \D_cache/cache[0][22] ,
         \D_cache/cache[0][23] , \D_cache/cache[0][24] ,
         \D_cache/cache[0][25] , \D_cache/cache[0][26] ,
         \D_cache/cache[0][27] , \D_cache/cache[0][28] ,
         \D_cache/cache[0][29] , \D_cache/cache[0][30] ,
         \D_cache/cache[0][31] , \D_cache/cache[0][32] ,
         \D_cache/cache[0][33] , \D_cache/cache[0][34] ,
         \D_cache/cache[0][35] , \D_cache/cache[0][36] ,
         \D_cache/cache[0][37] , \D_cache/cache[0][38] ,
         \D_cache/cache[0][39] , \D_cache/cache[0][40] ,
         \D_cache/cache[0][41] , \D_cache/cache[0][42] ,
         \D_cache/cache[0][43] , \D_cache/cache[0][44] ,
         \D_cache/cache[0][45] , \D_cache/cache[0][46] ,
         \D_cache/cache[0][47] , \D_cache/cache[0][48] ,
         \D_cache/cache[0][49] , \D_cache/cache[0][50] ,
         \D_cache/cache[0][51] , \D_cache/cache[0][52] ,
         \D_cache/cache[0][53] , \D_cache/cache[0][54] ,
         \D_cache/cache[0][55] , \D_cache/cache[0][56] ,
         \D_cache/cache[0][57] , \D_cache/cache[0][58] ,
         \D_cache/cache[0][59] , \D_cache/cache[0][60] ,
         \D_cache/cache[0][61] , \D_cache/cache[0][62] ,
         \D_cache/cache[0][63] , \D_cache/cache[0][64] ,
         \D_cache/cache[0][65] , \D_cache/cache[0][66] ,
         \D_cache/cache[0][67] , \D_cache/cache[0][68] ,
         \D_cache/cache[0][69] , \D_cache/cache[0][70] ,
         \D_cache/cache[0][71] , \D_cache/cache[0][72] ,
         \D_cache/cache[0][73] , \D_cache/cache[0][74] ,
         \D_cache/cache[0][75] , \D_cache/cache[0][76] ,
         \D_cache/cache[0][77] , \D_cache/cache[0][78] ,
         \D_cache/cache[0][79] , \D_cache/cache[0][80] ,
         \D_cache/cache[0][81] , \D_cache/cache[0][82] ,
         \D_cache/cache[0][83] , \D_cache/cache[0][84] ,
         \D_cache/cache[0][85] , \D_cache/cache[0][86] ,
         \D_cache/cache[0][87] , \D_cache/cache[0][88] ,
         \D_cache/cache[0][89] , \D_cache/cache[0][90] ,
         \D_cache/cache[0][91] , \D_cache/cache[0][92] ,
         \D_cache/cache[0][93] , \D_cache/cache[0][94] ,
         \D_cache/cache[0][95] , \D_cache/cache[0][96] ,
         \D_cache/cache[0][97] , \D_cache/cache[0][98] ,
         \D_cache/cache[0][99] , \D_cache/cache[0][100] ,
         \D_cache/cache[0][101] , \D_cache/cache[0][102] ,
         \D_cache/cache[0][103] , \D_cache/cache[0][104] ,
         \D_cache/cache[0][105] , \D_cache/cache[0][106] ,
         \D_cache/cache[0][107] , \D_cache/cache[0][108] ,
         \D_cache/cache[0][109] , \D_cache/cache[0][110] ,
         \D_cache/cache[0][111] , \D_cache/cache[0][112] ,
         \D_cache/cache[0][113] , \D_cache/cache[0][114] ,
         \D_cache/cache[0][115] , \D_cache/cache[0][116] ,
         \D_cache/cache[0][117] , \D_cache/cache[0][118] ,
         \D_cache/cache[0][119] , \D_cache/cache[0][120] ,
         \D_cache/cache[0][121] , \D_cache/cache[0][122] ,
         \D_cache/cache[0][123] , \D_cache/cache[0][124] ,
         \D_cache/cache[0][125] , \D_cache/cache[0][126] ,
         \D_cache/cache[0][127] , \D_cache/cache[0][128] ,
         \D_cache/cache[0][129] , \D_cache/cache[0][130] ,
         \D_cache/cache[0][131] , \D_cache/cache[0][132] ,
         \D_cache/cache[0][133] , \D_cache/cache[0][134] ,
         \D_cache/cache[0][135] , \D_cache/cache[0][136] ,
         \D_cache/cache[0][137] , \D_cache/cache[0][138] ,
         \D_cache/cache[0][139] , \D_cache/cache[0][140] ,
         \D_cache/cache[0][141] , \D_cache/cache[0][142] ,
         \D_cache/cache[0][143] , \D_cache/cache[0][144] ,
         \D_cache/cache[0][145] , \D_cache/cache[0][146] ,
         \D_cache/cache[0][147] , \D_cache/cache[0][148] ,
         \D_cache/cache[0][149] , \D_cache/cache[0][150] ,
         \D_cache/cache[0][151] , \D_cache/cache[0][152] ,
         \D_cache/cache[0][153] , \D_cache/cache[0][154] ,
         \i_MIPS/Pred_2bit/n8 , \i_MIPS/Pred_2bit/n7 , \i_MIPS/Pred_2bit/n1 ,
         \i_MIPS/Pred_2bit/current_state[0] ,
         \i_MIPS/Pred_2bit/current_state[1] , \i_MIPS/PC/n62 , \i_MIPS/PC/n61 ,
         \i_MIPS/PC/n60 , \i_MIPS/PC/n59 , \i_MIPS/PC/n58 , \i_MIPS/PC/n57 ,
         \i_MIPS/PC/n56 , \i_MIPS/PC/n55 , \i_MIPS/PC/n54 , \i_MIPS/PC/n53 ,
         \i_MIPS/PC/n52 , \i_MIPS/PC/n51 , \i_MIPS/PC/n50 , \i_MIPS/PC/n49 ,
         \i_MIPS/PC/n48 , \i_MIPS/PC/n47 , \i_MIPS/PC/n46 , \i_MIPS/PC/n45 ,
         \i_MIPS/PC/n44 , \i_MIPS/PC/n43 , \i_MIPS/PC/n42 , \i_MIPS/PC/n41 ,
         \i_MIPS/PC/n40 , \i_MIPS/PC/n39 , \i_MIPS/PC/n38 , \i_MIPS/PC/n37 ,
         \i_MIPS/PC/n36 , \i_MIPS/PC/n35 , \i_MIPS/PC/n34 , \i_MIPS/PC/n33 ,
         \i_MIPS/PC/n32 , \i_MIPS/PC/n31 , \i_MIPS/PC/n30 , \i_MIPS/PC/n29 ,
         \i_MIPS/PC/n28 , \i_MIPS/PC/n27 , \i_MIPS/PC/n26 , \i_MIPS/PC/n25 ,
         \i_MIPS/PC/n24 , \i_MIPS/PC/n23 , \i_MIPS/PC/n22 , \i_MIPS/PC/n21 ,
         \i_MIPS/PC/n20 , \i_MIPS/PC/n19 , \i_MIPS/PC/n18 , \i_MIPS/PC/n17 ,
         \i_MIPS/PC/n16 , \i_MIPS/PC/n15 , \i_MIPS/PC/n14 , \i_MIPS/PC/n13 ,
         \i_MIPS/PC/n9 , \i_MIPS/PC/n5 , \i_MIPS/PC/n4 , \i_MIPS/PC/n3 ,
         \i_MIPS/Register/n1139 , \i_MIPS/Register/n1138 ,
         \i_MIPS/Register/n1137 , \i_MIPS/Register/n1136 ,
         \i_MIPS/Register/n1135 , \i_MIPS/Register/n1134 ,
         \i_MIPS/Register/n1133 , \i_MIPS/Register/n1132 ,
         \i_MIPS/Register/n1131 , \i_MIPS/Register/n1130 ,
         \i_MIPS/Register/n1129 , \i_MIPS/Register/n1128 ,
         \i_MIPS/Register/n1127 , \i_MIPS/Register/n1126 ,
         \i_MIPS/Register/n1125 , \i_MIPS/Register/n1124 ,
         \i_MIPS/Register/n1123 , \i_MIPS/Register/n1122 ,
         \i_MIPS/Register/n1121 , \i_MIPS/Register/n1120 ,
         \i_MIPS/Register/n1119 , \i_MIPS/Register/n1118 ,
         \i_MIPS/Register/n1117 , \i_MIPS/Register/n1116 ,
         \i_MIPS/Register/n1115 , \i_MIPS/Register/n1114 ,
         \i_MIPS/Register/n1113 , \i_MIPS/Register/n1112 ,
         \i_MIPS/Register/n1111 , \i_MIPS/Register/n1110 ,
         \i_MIPS/Register/n1109 , \i_MIPS/Register/n1108 ,
         \i_MIPS/Register/n1107 , \i_MIPS/Register/n1106 ,
         \i_MIPS/Register/n1105 , \i_MIPS/Register/n1104 ,
         \i_MIPS/Register/n1103 , \i_MIPS/Register/n1102 ,
         \i_MIPS/Register/n1101 , \i_MIPS/Register/n1100 ,
         \i_MIPS/Register/n1099 , \i_MIPS/Register/n1098 ,
         \i_MIPS/Register/n1097 , \i_MIPS/Register/n1096 ,
         \i_MIPS/Register/n1095 , \i_MIPS/Register/n1094 ,
         \i_MIPS/Register/n1093 , \i_MIPS/Register/n1092 ,
         \i_MIPS/Register/n1091 , \i_MIPS/Register/n1090 ,
         \i_MIPS/Register/n1089 , \i_MIPS/Register/n1088 ,
         \i_MIPS/Register/n1087 , \i_MIPS/Register/n1086 ,
         \i_MIPS/Register/n1085 , \i_MIPS/Register/n1084 ,
         \i_MIPS/Register/n1083 , \i_MIPS/Register/n1082 ,
         \i_MIPS/Register/n1081 , \i_MIPS/Register/n1080 ,
         \i_MIPS/Register/n1079 , \i_MIPS/Register/n1078 ,
         \i_MIPS/Register/n1077 , \i_MIPS/Register/n1076 ,
         \i_MIPS/Register/n1075 , \i_MIPS/Register/n1074 ,
         \i_MIPS/Register/n1073 , \i_MIPS/Register/n1072 ,
         \i_MIPS/Register/n1071 , \i_MIPS/Register/n1070 ,
         \i_MIPS/Register/n1069 , \i_MIPS/Register/n1068 ,
         \i_MIPS/Register/n1067 , \i_MIPS/Register/n1066 ,
         \i_MIPS/Register/n1065 , \i_MIPS/Register/n1064 ,
         \i_MIPS/Register/n1063 , \i_MIPS/Register/n1062 ,
         \i_MIPS/Register/n1061 , \i_MIPS/Register/n1060 ,
         \i_MIPS/Register/n1059 , \i_MIPS/Register/n1058 ,
         \i_MIPS/Register/n1057 , \i_MIPS/Register/n1056 ,
         \i_MIPS/Register/n1055 , \i_MIPS/Register/n1054 ,
         \i_MIPS/Register/n1053 , \i_MIPS/Register/n1052 ,
         \i_MIPS/Register/n1051 , \i_MIPS/Register/n1050 ,
         \i_MIPS/Register/n1049 , \i_MIPS/Register/n1048 ,
         \i_MIPS/Register/n1047 , \i_MIPS/Register/n1046 ,
         \i_MIPS/Register/n1045 , \i_MIPS/Register/n1044 ,
         \i_MIPS/Register/n1043 , \i_MIPS/Register/n1042 ,
         \i_MIPS/Register/n1041 , \i_MIPS/Register/n1040 ,
         \i_MIPS/Register/n1039 , \i_MIPS/Register/n1038 ,
         \i_MIPS/Register/n1037 , \i_MIPS/Register/n1036 ,
         \i_MIPS/Register/n1035 , \i_MIPS/Register/n1034 ,
         \i_MIPS/Register/n1033 , \i_MIPS/Register/n1032 ,
         \i_MIPS/Register/n1031 , \i_MIPS/Register/n1030 ,
         \i_MIPS/Register/n1029 , \i_MIPS/Register/n1028 ,
         \i_MIPS/Register/n1027 , \i_MIPS/Register/n1026 ,
         \i_MIPS/Register/n1025 , \i_MIPS/Register/n1024 ,
         \i_MIPS/Register/n1023 , \i_MIPS/Register/n1022 ,
         \i_MIPS/Register/n1021 , \i_MIPS/Register/n1020 ,
         \i_MIPS/Register/n1019 , \i_MIPS/Register/n1018 ,
         \i_MIPS/Register/n1017 , \i_MIPS/Register/n1016 ,
         \i_MIPS/Register/n1015 , \i_MIPS/Register/n1014 ,
         \i_MIPS/Register/n1013 , \i_MIPS/Register/n1012 ,
         \i_MIPS/Register/n1011 , \i_MIPS/Register/n1010 ,
         \i_MIPS/Register/n1009 , \i_MIPS/Register/n1008 ,
         \i_MIPS/Register/n1007 , \i_MIPS/Register/n1006 ,
         \i_MIPS/Register/n1005 , \i_MIPS/Register/n1004 ,
         \i_MIPS/Register/n1003 , \i_MIPS/Register/n1002 ,
         \i_MIPS/Register/n1001 , \i_MIPS/Register/n1000 ,
         \i_MIPS/Register/n999 , \i_MIPS/Register/n998 ,
         \i_MIPS/Register/n997 , \i_MIPS/Register/n996 ,
         \i_MIPS/Register/n995 , \i_MIPS/Register/n994 ,
         \i_MIPS/Register/n993 , \i_MIPS/Register/n992 ,
         \i_MIPS/Register/n991 , \i_MIPS/Register/n990 ,
         \i_MIPS/Register/n989 , \i_MIPS/Register/n988 ,
         \i_MIPS/Register/n987 , \i_MIPS/Register/n986 ,
         \i_MIPS/Register/n985 , \i_MIPS/Register/n984 ,
         \i_MIPS/Register/n983 , \i_MIPS/Register/n982 ,
         \i_MIPS/Register/n981 , \i_MIPS/Register/n980 ,
         \i_MIPS/Register/n979 , \i_MIPS/Register/n978 ,
         \i_MIPS/Register/n977 , \i_MIPS/Register/n976 ,
         \i_MIPS/Register/n975 , \i_MIPS/Register/n974 ,
         \i_MIPS/Register/n973 , \i_MIPS/Register/n972 ,
         \i_MIPS/Register/n971 , \i_MIPS/Register/n970 ,
         \i_MIPS/Register/n969 , \i_MIPS/Register/n968 ,
         \i_MIPS/Register/n967 , \i_MIPS/Register/n966 ,
         \i_MIPS/Register/n965 , \i_MIPS/Register/n964 ,
         \i_MIPS/Register/n963 , \i_MIPS/Register/n962 ,
         \i_MIPS/Register/n961 , \i_MIPS/Register/n960 ,
         \i_MIPS/Register/n959 , \i_MIPS/Register/n958 ,
         \i_MIPS/Register/n957 , \i_MIPS/Register/n956 ,
         \i_MIPS/Register/n955 , \i_MIPS/Register/n954 ,
         \i_MIPS/Register/n953 , \i_MIPS/Register/n952 ,
         \i_MIPS/Register/n951 , \i_MIPS/Register/n950 ,
         \i_MIPS/Register/n949 , \i_MIPS/Register/n948 ,
         \i_MIPS/Register/n947 , \i_MIPS/Register/n946 ,
         \i_MIPS/Register/n945 , \i_MIPS/Register/n944 ,
         \i_MIPS/Register/n943 , \i_MIPS/Register/n942 ,
         \i_MIPS/Register/n941 , \i_MIPS/Register/n940 ,
         \i_MIPS/Register/n939 , \i_MIPS/Register/n938 ,
         \i_MIPS/Register/n937 , \i_MIPS/Register/n936 ,
         \i_MIPS/Register/n935 , \i_MIPS/Register/n934 ,
         \i_MIPS/Register/n933 , \i_MIPS/Register/n932 ,
         \i_MIPS/Register/n931 , \i_MIPS/Register/n930 ,
         \i_MIPS/Register/n929 , \i_MIPS/Register/n928 ,
         \i_MIPS/Register/n927 , \i_MIPS/Register/n926 ,
         \i_MIPS/Register/n925 , \i_MIPS/Register/n924 ,
         \i_MIPS/Register/n923 , \i_MIPS/Register/n922 ,
         \i_MIPS/Register/n921 , \i_MIPS/Register/n920 ,
         \i_MIPS/Register/n919 , \i_MIPS/Register/n918 ,
         \i_MIPS/Register/n917 , \i_MIPS/Register/n916 ,
         \i_MIPS/Register/n915 , \i_MIPS/Register/n914 ,
         \i_MIPS/Register/n913 , \i_MIPS/Register/n912 ,
         \i_MIPS/Register/n911 , \i_MIPS/Register/n910 ,
         \i_MIPS/Register/n909 , \i_MIPS/Register/n908 ,
         \i_MIPS/Register/n907 , \i_MIPS/Register/n906 ,
         \i_MIPS/Register/n905 , \i_MIPS/Register/n904 ,
         \i_MIPS/Register/n903 , \i_MIPS/Register/n902 ,
         \i_MIPS/Register/n901 , \i_MIPS/Register/n900 ,
         \i_MIPS/Register/n899 , \i_MIPS/Register/n898 ,
         \i_MIPS/Register/n897 , \i_MIPS/Register/n896 ,
         \i_MIPS/Register/n895 , \i_MIPS/Register/n894 ,
         \i_MIPS/Register/n893 , \i_MIPS/Register/n892 ,
         \i_MIPS/Register/n891 , \i_MIPS/Register/n890 ,
         \i_MIPS/Register/n889 , \i_MIPS/Register/n888 ,
         \i_MIPS/Register/n887 , \i_MIPS/Register/n886 ,
         \i_MIPS/Register/n885 , \i_MIPS/Register/n884 ,
         \i_MIPS/Register/n883 , \i_MIPS/Register/n882 ,
         \i_MIPS/Register/n881 , \i_MIPS/Register/n880 ,
         \i_MIPS/Register/n879 , \i_MIPS/Register/n878 ,
         \i_MIPS/Register/n877 , \i_MIPS/Register/n876 ,
         \i_MIPS/Register/n875 , \i_MIPS/Register/n874 ,
         \i_MIPS/Register/n873 , \i_MIPS/Register/n872 ,
         \i_MIPS/Register/n871 , \i_MIPS/Register/n870 ,
         \i_MIPS/Register/n869 , \i_MIPS/Register/n868 ,
         \i_MIPS/Register/n867 , \i_MIPS/Register/n866 ,
         \i_MIPS/Register/n865 , \i_MIPS/Register/n864 ,
         \i_MIPS/Register/n863 , \i_MIPS/Register/n862 ,
         \i_MIPS/Register/n861 , \i_MIPS/Register/n860 ,
         \i_MIPS/Register/n859 , \i_MIPS/Register/n858 ,
         \i_MIPS/Register/n857 , \i_MIPS/Register/n856 ,
         \i_MIPS/Register/n855 , \i_MIPS/Register/n854 ,
         \i_MIPS/Register/n853 , \i_MIPS/Register/n852 ,
         \i_MIPS/Register/n851 , \i_MIPS/Register/n850 ,
         \i_MIPS/Register/n849 , \i_MIPS/Register/n848 ,
         \i_MIPS/Register/n847 , \i_MIPS/Register/n846 ,
         \i_MIPS/Register/n845 , \i_MIPS/Register/n844 ,
         \i_MIPS/Register/n843 , \i_MIPS/Register/n842 ,
         \i_MIPS/Register/n841 , \i_MIPS/Register/n840 ,
         \i_MIPS/Register/n839 , \i_MIPS/Register/n838 ,
         \i_MIPS/Register/n837 , \i_MIPS/Register/n836 ,
         \i_MIPS/Register/n835 , \i_MIPS/Register/n834 ,
         \i_MIPS/Register/n833 , \i_MIPS/Register/n832 ,
         \i_MIPS/Register/n831 , \i_MIPS/Register/n830 ,
         \i_MIPS/Register/n829 , \i_MIPS/Register/n828 ,
         \i_MIPS/Register/n827 , \i_MIPS/Register/n826 ,
         \i_MIPS/Register/n825 , \i_MIPS/Register/n824 ,
         \i_MIPS/Register/n823 , \i_MIPS/Register/n822 ,
         \i_MIPS/Register/n821 , \i_MIPS/Register/n820 ,
         \i_MIPS/Register/n819 , \i_MIPS/Register/n818 ,
         \i_MIPS/Register/n817 , \i_MIPS/Register/n816 ,
         \i_MIPS/Register/n815 , \i_MIPS/Register/n814 ,
         \i_MIPS/Register/n813 , \i_MIPS/Register/n812 ,
         \i_MIPS/Register/n811 , \i_MIPS/Register/n810 ,
         \i_MIPS/Register/n809 , \i_MIPS/Register/n808 ,
         \i_MIPS/Register/n807 , \i_MIPS/Register/n806 ,
         \i_MIPS/Register/n805 , \i_MIPS/Register/n804 ,
         \i_MIPS/Register/n803 , \i_MIPS/Register/n802 ,
         \i_MIPS/Register/n801 , \i_MIPS/Register/n800 ,
         \i_MIPS/Register/n799 , \i_MIPS/Register/n798 ,
         \i_MIPS/Register/n797 , \i_MIPS/Register/n796 ,
         \i_MIPS/Register/n795 , \i_MIPS/Register/n794 ,
         \i_MIPS/Register/n793 , \i_MIPS/Register/n792 ,
         \i_MIPS/Register/n791 , \i_MIPS/Register/n790 ,
         \i_MIPS/Register/n789 , \i_MIPS/Register/n788 ,
         \i_MIPS/Register/n787 , \i_MIPS/Register/n786 ,
         \i_MIPS/Register/n785 , \i_MIPS/Register/n784 ,
         \i_MIPS/Register/n783 , \i_MIPS/Register/n782 ,
         \i_MIPS/Register/n781 , \i_MIPS/Register/n780 ,
         \i_MIPS/Register/n779 , \i_MIPS/Register/n778 ,
         \i_MIPS/Register/n777 , \i_MIPS/Register/n776 ,
         \i_MIPS/Register/n775 , \i_MIPS/Register/n774 ,
         \i_MIPS/Register/n773 , \i_MIPS/Register/n772 ,
         \i_MIPS/Register/n771 , \i_MIPS/Register/n770 ,
         \i_MIPS/Register/n769 , \i_MIPS/Register/n768 ,
         \i_MIPS/Register/n767 , \i_MIPS/Register/n766 ,
         \i_MIPS/Register/n765 , \i_MIPS/Register/n764 ,
         \i_MIPS/Register/n763 , \i_MIPS/Register/n762 ,
         \i_MIPS/Register/n761 , \i_MIPS/Register/n760 ,
         \i_MIPS/Register/n759 , \i_MIPS/Register/n758 ,
         \i_MIPS/Register/n757 , \i_MIPS/Register/n756 ,
         \i_MIPS/Register/n755 , \i_MIPS/Register/n754 ,
         \i_MIPS/Register/n753 , \i_MIPS/Register/n752 ,
         \i_MIPS/Register/n751 , \i_MIPS/Register/n750 ,
         \i_MIPS/Register/n749 , \i_MIPS/Register/n748 ,
         \i_MIPS/Register/n747 , \i_MIPS/Register/n746 ,
         \i_MIPS/Register/n745 , \i_MIPS/Register/n744 ,
         \i_MIPS/Register/n743 , \i_MIPS/Register/n742 ,
         \i_MIPS/Register/n741 , \i_MIPS/Register/n740 ,
         \i_MIPS/Register/n739 , \i_MIPS/Register/n738 ,
         \i_MIPS/Register/n737 , \i_MIPS/Register/n736 ,
         \i_MIPS/Register/n735 , \i_MIPS/Register/n734 ,
         \i_MIPS/Register/n733 , \i_MIPS/Register/n732 ,
         \i_MIPS/Register/n731 , \i_MIPS/Register/n730 ,
         \i_MIPS/Register/n729 , \i_MIPS/Register/n728 ,
         \i_MIPS/Register/n727 , \i_MIPS/Register/n726 ,
         \i_MIPS/Register/n725 , \i_MIPS/Register/n724 ,
         \i_MIPS/Register/n723 , \i_MIPS/Register/n722 ,
         \i_MIPS/Register/n721 , \i_MIPS/Register/n720 ,
         \i_MIPS/Register/n719 , \i_MIPS/Register/n718 ,
         \i_MIPS/Register/n717 , \i_MIPS/Register/n716 ,
         \i_MIPS/Register/n715 , \i_MIPS/Register/n714 ,
         \i_MIPS/Register/n713 , \i_MIPS/Register/n712 ,
         \i_MIPS/Register/n711 , \i_MIPS/Register/n710 ,
         \i_MIPS/Register/n709 , \i_MIPS/Register/n708 ,
         \i_MIPS/Register/n707 , \i_MIPS/Register/n706 ,
         \i_MIPS/Register/n705 , \i_MIPS/Register/n704 ,
         \i_MIPS/Register/n703 , \i_MIPS/Register/n702 ,
         \i_MIPS/Register/n701 , \i_MIPS/Register/n700 ,
         \i_MIPS/Register/n699 , \i_MIPS/Register/n698 ,
         \i_MIPS/Register/n697 , \i_MIPS/Register/n696 ,
         \i_MIPS/Register/n695 , \i_MIPS/Register/n694 ,
         \i_MIPS/Register/n693 , \i_MIPS/Register/n692 ,
         \i_MIPS/Register/n691 , \i_MIPS/Register/n690 ,
         \i_MIPS/Register/n689 , \i_MIPS/Register/n688 ,
         \i_MIPS/Register/n687 , \i_MIPS/Register/n686 ,
         \i_MIPS/Register/n685 , \i_MIPS/Register/n684 ,
         \i_MIPS/Register/n683 , \i_MIPS/Register/n682 ,
         \i_MIPS/Register/n681 , \i_MIPS/Register/n680 ,
         \i_MIPS/Register/n679 , \i_MIPS/Register/n678 ,
         \i_MIPS/Register/n677 , \i_MIPS/Register/n676 ,
         \i_MIPS/Register/n675 , \i_MIPS/Register/n674 ,
         \i_MIPS/Register/n673 , \i_MIPS/Register/n672 ,
         \i_MIPS/Register/n671 , \i_MIPS/Register/n670 ,
         \i_MIPS/Register/n669 , \i_MIPS/Register/n668 ,
         \i_MIPS/Register/n667 , \i_MIPS/Register/n666 ,
         \i_MIPS/Register/n665 , \i_MIPS/Register/n664 ,
         \i_MIPS/Register/n663 , \i_MIPS/Register/n662 ,
         \i_MIPS/Register/n661 , \i_MIPS/Register/n660 ,
         \i_MIPS/Register/n659 , \i_MIPS/Register/n658 ,
         \i_MIPS/Register/n657 , \i_MIPS/Register/n656 ,
         \i_MIPS/Register/n655 , \i_MIPS/Register/n654 ,
         \i_MIPS/Register/n653 , \i_MIPS/Register/n652 ,
         \i_MIPS/Register/n651 , \i_MIPS/Register/n650 ,
         \i_MIPS/Register/n649 , \i_MIPS/Register/n648 ,
         \i_MIPS/Register/n647 , \i_MIPS/Register/n646 ,
         \i_MIPS/Register/n645 , \i_MIPS/Register/n644 ,
         \i_MIPS/Register/n643 , \i_MIPS/Register/n642 ,
         \i_MIPS/Register/n641 , \i_MIPS/Register/n640 ,
         \i_MIPS/Register/n639 , \i_MIPS/Register/n638 ,
         \i_MIPS/Register/n637 , \i_MIPS/Register/n636 ,
         \i_MIPS/Register/n635 , \i_MIPS/Register/n634 ,
         \i_MIPS/Register/n633 , \i_MIPS/Register/n632 ,
         \i_MIPS/Register/n631 , \i_MIPS/Register/n630 ,
         \i_MIPS/Register/n629 , \i_MIPS/Register/n628 ,
         \i_MIPS/Register/n627 , \i_MIPS/Register/n626 ,
         \i_MIPS/Register/n625 , \i_MIPS/Register/n624 ,
         \i_MIPS/Register/n623 , \i_MIPS/Register/n622 ,
         \i_MIPS/Register/n621 , \i_MIPS/Register/n620 ,
         \i_MIPS/Register/n619 , \i_MIPS/Register/n618 ,
         \i_MIPS/Register/n617 , \i_MIPS/Register/n616 ,
         \i_MIPS/Register/n615 , \i_MIPS/Register/n614 ,
         \i_MIPS/Register/n613 , \i_MIPS/Register/n612 ,
         \i_MIPS/Register/n611 , \i_MIPS/Register/n610 ,
         \i_MIPS/Register/n609 , \i_MIPS/Register/n608 ,
         \i_MIPS/Register/n607 , \i_MIPS/Register/n606 ,
         \i_MIPS/Register/n605 , \i_MIPS/Register/n604 ,
         \i_MIPS/Register/n603 , \i_MIPS/Register/n602 ,
         \i_MIPS/Register/n601 , \i_MIPS/Register/n600 ,
         \i_MIPS/Register/n599 , \i_MIPS/Register/n598 ,
         \i_MIPS/Register/n597 , \i_MIPS/Register/n596 ,
         \i_MIPS/Register/n595 , \i_MIPS/Register/n594 ,
         \i_MIPS/Register/n593 , \i_MIPS/Register/n592 ,
         \i_MIPS/Register/n591 , \i_MIPS/Register/n590 ,
         \i_MIPS/Register/n589 , \i_MIPS/Register/n588 ,
         \i_MIPS/Register/n587 , \i_MIPS/Register/n586 ,
         \i_MIPS/Register/n585 , \i_MIPS/Register/n584 ,
         \i_MIPS/Register/n583 , \i_MIPS/Register/n582 ,
         \i_MIPS/Register/n581 , \i_MIPS/Register/n580 ,
         \i_MIPS/Register/n579 , \i_MIPS/Register/n578 ,
         \i_MIPS/Register/n577 , \i_MIPS/Register/n576 ,
         \i_MIPS/Register/n575 , \i_MIPS/Register/n574 ,
         \i_MIPS/Register/n573 , \i_MIPS/Register/n572 ,
         \i_MIPS/Register/n571 , \i_MIPS/Register/n570 ,
         \i_MIPS/Register/n569 , \i_MIPS/Register/n568 ,
         \i_MIPS/Register/n567 , \i_MIPS/Register/n566 ,
         \i_MIPS/Register/n565 , \i_MIPS/Register/n564 ,
         \i_MIPS/Register/n563 , \i_MIPS/Register/n562 ,
         \i_MIPS/Register/n561 , \i_MIPS/Register/n560 ,
         \i_MIPS/Register/n559 , \i_MIPS/Register/n558 ,
         \i_MIPS/Register/n557 , \i_MIPS/Register/n556 ,
         \i_MIPS/Register/n555 , \i_MIPS/Register/n554 ,
         \i_MIPS/Register/n553 , \i_MIPS/Register/n552 ,
         \i_MIPS/Register/n551 , \i_MIPS/Register/n550 ,
         \i_MIPS/Register/n549 , \i_MIPS/Register/n548 ,
         \i_MIPS/Register/n547 , \i_MIPS/Register/n546 ,
         \i_MIPS/Register/n545 , \i_MIPS/Register/n544 ,
         \i_MIPS/Register/n543 , \i_MIPS/Register/n542 ,
         \i_MIPS/Register/n541 , \i_MIPS/Register/n540 ,
         \i_MIPS/Register/n539 , \i_MIPS/Register/n538 ,
         \i_MIPS/Register/n537 , \i_MIPS/Register/n536 ,
         \i_MIPS/Register/n535 , \i_MIPS/Register/n534 ,
         \i_MIPS/Register/n533 , \i_MIPS/Register/n532 ,
         \i_MIPS/Register/n531 , \i_MIPS/Register/n530 ,
         \i_MIPS/Register/n529 , \i_MIPS/Register/n528 ,
         \i_MIPS/Register/n527 , \i_MIPS/Register/n526 ,
         \i_MIPS/Register/n525 , \i_MIPS/Register/n524 ,
         \i_MIPS/Register/n523 , \i_MIPS/Register/n522 ,
         \i_MIPS/Register/n521 , \i_MIPS/Register/n520 ,
         \i_MIPS/Register/n519 , \i_MIPS/Register/n518 ,
         \i_MIPS/Register/n517 , \i_MIPS/Register/n516 ,
         \i_MIPS/Register/n515 , \i_MIPS/Register/n514 ,
         \i_MIPS/Register/n513 , \i_MIPS/Register/n512 ,
         \i_MIPS/Register/n511 , \i_MIPS/Register/n510 ,
         \i_MIPS/Register/n509 , \i_MIPS/Register/n508 ,
         \i_MIPS/Register/n507 , \i_MIPS/Register/n506 ,
         \i_MIPS/Register/n505 , \i_MIPS/Register/n504 ,
         \i_MIPS/Register/n503 , \i_MIPS/Register/n502 ,
         \i_MIPS/Register/n501 , \i_MIPS/Register/n500 ,
         \i_MIPS/Register/n499 , \i_MIPS/Register/n498 ,
         \i_MIPS/Register/n497 , \i_MIPS/Register/n496 ,
         \i_MIPS/Register/n495 , \i_MIPS/Register/n494 ,
         \i_MIPS/Register/n493 , \i_MIPS/Register/n492 ,
         \i_MIPS/Register/n491 , \i_MIPS/Register/n490 ,
         \i_MIPS/Register/n489 , \i_MIPS/Register/n488 ,
         \i_MIPS/Register/n487 , \i_MIPS/Register/n486 ,
         \i_MIPS/Register/n485 , \i_MIPS/Register/n484 ,
         \i_MIPS/Register/n483 , \i_MIPS/Register/n482 ,
         \i_MIPS/Register/n481 , \i_MIPS/Register/n480 ,
         \i_MIPS/Register/n479 , \i_MIPS/Register/n478 ,
         \i_MIPS/Register/n477 , \i_MIPS/Register/n476 ,
         \i_MIPS/Register/n475 , \i_MIPS/Register/n474 ,
         \i_MIPS/Register/n473 , \i_MIPS/Register/n472 ,
         \i_MIPS/Register/n471 , \i_MIPS/Register/n470 ,
         \i_MIPS/Register/n469 , \i_MIPS/Register/n468 ,
         \i_MIPS/Register/n467 , \i_MIPS/Register/n466 ,
         \i_MIPS/Register/n465 , \i_MIPS/Register/n464 ,
         \i_MIPS/Register/n463 , \i_MIPS/Register/n462 ,
         \i_MIPS/Register/n461 , \i_MIPS/Register/n460 ,
         \i_MIPS/Register/n459 , \i_MIPS/Register/n458 ,
         \i_MIPS/Register/n457 , \i_MIPS/Register/n456 ,
         \i_MIPS/Register/n455 , \i_MIPS/Register/n454 ,
         \i_MIPS/Register/n453 , \i_MIPS/Register/n452 ,
         \i_MIPS/Register/n451 , \i_MIPS/Register/n450 ,
         \i_MIPS/Register/n449 , \i_MIPS/Register/n448 ,
         \i_MIPS/Register/n447 , \i_MIPS/Register/n446 ,
         \i_MIPS/Register/n445 , \i_MIPS/Register/n444 ,
         \i_MIPS/Register/n443 , \i_MIPS/Register/n442 ,
         \i_MIPS/Register/n441 , \i_MIPS/Register/n440 ,
         \i_MIPS/Register/n439 , \i_MIPS/Register/n438 ,
         \i_MIPS/Register/n437 , \i_MIPS/Register/n436 ,
         \i_MIPS/Register/n435 , \i_MIPS/Register/n434 ,
         \i_MIPS/Register/n433 , \i_MIPS/Register/n432 ,
         \i_MIPS/Register/n431 , \i_MIPS/Register/n430 ,
         \i_MIPS/Register/n429 , \i_MIPS/Register/n428 ,
         \i_MIPS/Register/n427 , \i_MIPS/Register/n426 ,
         \i_MIPS/Register/n425 , \i_MIPS/Register/n424 ,
         \i_MIPS/Register/n423 , \i_MIPS/Register/n422 ,
         \i_MIPS/Register/n421 , \i_MIPS/Register/n420 ,
         \i_MIPS/Register/n419 , \i_MIPS/Register/n418 ,
         \i_MIPS/Register/n417 , \i_MIPS/Register/n416 ,
         \i_MIPS/Register/n415 , \i_MIPS/Register/n414 ,
         \i_MIPS/Register/n413 , \i_MIPS/Register/n412 ,
         \i_MIPS/Register/n411 , \i_MIPS/Register/n410 ,
         \i_MIPS/Register/n409 , \i_MIPS/Register/n408 ,
         \i_MIPS/Register/n407 , \i_MIPS/Register/n406 ,
         \i_MIPS/Register/n405 , \i_MIPS/Register/n404 ,
         \i_MIPS/Register/n403 , \i_MIPS/Register/n402 ,
         \i_MIPS/Register/n401 , \i_MIPS/Register/n400 ,
         \i_MIPS/Register/n399 , \i_MIPS/Register/n398 ,
         \i_MIPS/Register/n397 , \i_MIPS/Register/n396 ,
         \i_MIPS/Register/n395 , \i_MIPS/Register/n394 ,
         \i_MIPS/Register/n393 , \i_MIPS/Register/n392 ,
         \i_MIPS/Register/n391 , \i_MIPS/Register/n390 ,
         \i_MIPS/Register/n389 , \i_MIPS/Register/n388 ,
         \i_MIPS/Register/n387 , \i_MIPS/Register/n386 ,
         \i_MIPS/Register/n385 , \i_MIPS/Register/n384 ,
         \i_MIPS/Register/n383 , \i_MIPS/Register/n382 ,
         \i_MIPS/Register/n381 , \i_MIPS/Register/n380 ,
         \i_MIPS/Register/n379 , \i_MIPS/Register/n378 ,
         \i_MIPS/Register/n377 , \i_MIPS/Register/n376 ,
         \i_MIPS/Register/n375 , \i_MIPS/Register/n374 ,
         \i_MIPS/Register/n373 , \i_MIPS/Register/n372 ,
         \i_MIPS/Register/n371 , \i_MIPS/Register/n370 ,
         \i_MIPS/Register/n369 , \i_MIPS/Register/n368 ,
         \i_MIPS/Register/n367 , \i_MIPS/Register/n366 ,
         \i_MIPS/Register/n365 , \i_MIPS/Register/n364 ,
         \i_MIPS/Register/n363 , \i_MIPS/Register/n362 ,
         \i_MIPS/Register/n361 , \i_MIPS/Register/n360 ,
         \i_MIPS/Register/n359 , \i_MIPS/Register/n358 ,
         \i_MIPS/Register/n357 , \i_MIPS/Register/n356 ,
         \i_MIPS/Register/n355 , \i_MIPS/Register/n354 ,
         \i_MIPS/Register/n353 , \i_MIPS/Register/n352 ,
         \i_MIPS/Register/n351 , \i_MIPS/Register/n350 ,
         \i_MIPS/Register/n349 , \i_MIPS/Register/n348 ,
         \i_MIPS/Register/n347 , \i_MIPS/Register/n346 ,
         \i_MIPS/Register/n345 , \i_MIPS/Register/n344 ,
         \i_MIPS/Register/n343 , \i_MIPS/Register/n342 ,
         \i_MIPS/Register/n341 , \i_MIPS/Register/n340 ,
         \i_MIPS/Register/n339 , \i_MIPS/Register/n338 ,
         \i_MIPS/Register/n337 , \i_MIPS/Register/n336 ,
         \i_MIPS/Register/n335 , \i_MIPS/Register/n334 ,
         \i_MIPS/Register/n333 , \i_MIPS/Register/n332 ,
         \i_MIPS/Register/n331 , \i_MIPS/Register/n330 ,
         \i_MIPS/Register/n329 , \i_MIPS/Register/n328 ,
         \i_MIPS/Register/n327 , \i_MIPS/Register/n326 ,
         \i_MIPS/Register/n325 , \i_MIPS/Register/n324 ,
         \i_MIPS/Register/n323 , \i_MIPS/Register/n322 ,
         \i_MIPS/Register/n321 , \i_MIPS/Register/n320 ,
         \i_MIPS/Register/n319 , \i_MIPS/Register/n318 ,
         \i_MIPS/Register/n317 , \i_MIPS/Register/n316 ,
         \i_MIPS/Register/n315 , \i_MIPS/Register/n314 ,
         \i_MIPS/Register/n313 , \i_MIPS/Register/n312 ,
         \i_MIPS/Register/n311 , \i_MIPS/Register/n310 ,
         \i_MIPS/Register/n309 , \i_MIPS/Register/n308 ,
         \i_MIPS/Register/n307 , \i_MIPS/Register/n306 ,
         \i_MIPS/Register/n305 , \i_MIPS/Register/n304 ,
         \i_MIPS/Register/n303 , \i_MIPS/Register/n302 ,
         \i_MIPS/Register/n301 , \i_MIPS/Register/n300 ,
         \i_MIPS/Register/n299 , \i_MIPS/Register/n298 ,
         \i_MIPS/Register/n297 , \i_MIPS/Register/n296 ,
         \i_MIPS/Register/n295 , \i_MIPS/Register/n294 ,
         \i_MIPS/Register/n293 , \i_MIPS/Register/n292 ,
         \i_MIPS/Register/n291 , \i_MIPS/Register/n290 ,
         \i_MIPS/Register/n289 , \i_MIPS/Register/n288 ,
         \i_MIPS/Register/n287 , \i_MIPS/Register/n286 ,
         \i_MIPS/Register/n285 , \i_MIPS/Register/n284 ,
         \i_MIPS/Register/n283 , \i_MIPS/Register/n282 ,
         \i_MIPS/Register/n281 , \i_MIPS/Register/n280 ,
         \i_MIPS/Register/n279 , \i_MIPS/Register/n278 ,
         \i_MIPS/Register/n277 , \i_MIPS/Register/n276 ,
         \i_MIPS/Register/n275 , \i_MIPS/Register/n274 ,
         \i_MIPS/Register/n273 , \i_MIPS/Register/n272 ,
         \i_MIPS/Register/n271 , \i_MIPS/Register/n270 ,
         \i_MIPS/Register/n269 , \i_MIPS/Register/n268 ,
         \i_MIPS/Register/n267 , \i_MIPS/Register/n266 ,
         \i_MIPS/Register/n265 , \i_MIPS/Register/n264 ,
         \i_MIPS/Register/n263 , \i_MIPS/Register/n262 ,
         \i_MIPS/Register/n261 , \i_MIPS/Register/n260 ,
         \i_MIPS/Register/n259 , \i_MIPS/Register/n258 ,
         \i_MIPS/Register/n257 , \i_MIPS/Register/n256 ,
         \i_MIPS/Register/n255 , \i_MIPS/Register/n254 ,
         \i_MIPS/Register/n253 , \i_MIPS/Register/n252 ,
         \i_MIPS/Register/n251 , \i_MIPS/Register/n250 ,
         \i_MIPS/Register/n249 , \i_MIPS/Register/n248 ,
         \i_MIPS/Register/n247 , \i_MIPS/Register/n246 ,
         \i_MIPS/Register/n245 , \i_MIPS/Register/n244 ,
         \i_MIPS/Register/n243 , \i_MIPS/Register/n242 ,
         \i_MIPS/Register/n241 , \i_MIPS/Register/n240 ,
         \i_MIPS/Register/n239 , \i_MIPS/Register/n238 ,
         \i_MIPS/Register/n237 , \i_MIPS/Register/n236 ,
         \i_MIPS/Register/n235 , \i_MIPS/Register/n234 ,
         \i_MIPS/Register/n233 , \i_MIPS/Register/n232 ,
         \i_MIPS/Register/n231 , \i_MIPS/Register/n230 ,
         \i_MIPS/Register/n229 , \i_MIPS/Register/n228 ,
         \i_MIPS/Register/n227 , \i_MIPS/Register/n226 ,
         \i_MIPS/Register/n225 , \i_MIPS/Register/n224 ,
         \i_MIPS/Register/n223 , \i_MIPS/Register/n222 ,
         \i_MIPS/Register/n221 , \i_MIPS/Register/n220 ,
         \i_MIPS/Register/n219 , \i_MIPS/Register/n218 ,
         \i_MIPS/Register/n217 , \i_MIPS/Register/n216 ,
         \i_MIPS/Register/n215 , \i_MIPS/Register/n214 ,
         \i_MIPS/Register/n213 , \i_MIPS/Register/n212 ,
         \i_MIPS/Register/n211 , \i_MIPS/Register/n210 ,
         \i_MIPS/Register/n209 , \i_MIPS/Register/n208 ,
         \i_MIPS/Register/n207 , \i_MIPS/Register/n206 ,
         \i_MIPS/Register/n205 , \i_MIPS/Register/n204 ,
         \i_MIPS/Register/n203 , \i_MIPS/Register/n202 ,
         \i_MIPS/Register/n201 , \i_MIPS/Register/n200 ,
         \i_MIPS/Register/n199 , \i_MIPS/Register/n198 ,
         \i_MIPS/Register/n197 , \i_MIPS/Register/n196 ,
         \i_MIPS/Register/n195 , \i_MIPS/Register/n194 ,
         \i_MIPS/Register/n193 , \i_MIPS/Register/n192 ,
         \i_MIPS/Register/n191 , \i_MIPS/Register/n190 ,
         \i_MIPS/Register/n189 , \i_MIPS/Register/n188 ,
         \i_MIPS/Register/n187 , \i_MIPS/Register/n186 ,
         \i_MIPS/Register/n185 , \i_MIPS/Register/n184 ,
         \i_MIPS/Register/n183 , \i_MIPS/Register/n182 ,
         \i_MIPS/Register/n181 , \i_MIPS/Register/n180 ,
         \i_MIPS/Register/n179 , \i_MIPS/Register/n178 ,
         \i_MIPS/Register/n177 , \i_MIPS/Register/n176 ,
         \i_MIPS/Register/n175 , \i_MIPS/Register/n174 ,
         \i_MIPS/Register/n173 , \i_MIPS/Register/n172 ,
         \i_MIPS/Register/n171 , \i_MIPS/Register/n170 ,
         \i_MIPS/Register/n169 , \i_MIPS/Register/n168 ,
         \i_MIPS/Register/n167 , \i_MIPS/Register/n166 ,
         \i_MIPS/Register/n165 , \i_MIPS/Register/n164 ,
         \i_MIPS/Register/n163 , \i_MIPS/Register/n162 ,
         \i_MIPS/Register/n161 , \i_MIPS/Register/n160 ,
         \i_MIPS/Register/n159 , \i_MIPS/Register/n158 ,
         \i_MIPS/Register/n157 , \i_MIPS/Register/n156 ,
         \i_MIPS/Register/n155 , \i_MIPS/Register/n154 ,
         \i_MIPS/Register/n153 , \i_MIPS/Register/n152 ,
         \i_MIPS/Register/n151 , \i_MIPS/Register/n150 ,
         \i_MIPS/Register/n149 , \i_MIPS/Register/n148 ,
         \i_MIPS/Register/n147 , \i_MIPS/Register/n146 ,
         \i_MIPS/Register/n145 , \i_MIPS/Register/n144 ,
         \i_MIPS/Register/n143 , \i_MIPS/Register/n142 ,
         \i_MIPS/Register/n141 , \i_MIPS/Register/n140 ,
         \i_MIPS/Register/n139 , \i_MIPS/Register/n138 ,
         \i_MIPS/Register/n137 , \i_MIPS/Register/n136 ,
         \i_MIPS/Register/n135 , \i_MIPS/Register/n134 ,
         \i_MIPS/Register/n133 , \i_MIPS/Register/n132 ,
         \i_MIPS/Register/n131 , \i_MIPS/Register/n130 ,
         \i_MIPS/Register/n129 , \i_MIPS/Register/n128 ,
         \i_MIPS/Register/n127 , \i_MIPS/Register/n126 ,
         \i_MIPS/Register/n125 , \i_MIPS/Register/n124 ,
         \i_MIPS/Register/n123 , \i_MIPS/Register/n122 ,
         \i_MIPS/Register/n121 , \i_MIPS/Register/n120 ,
         \i_MIPS/Register/n119 , \i_MIPS/Register/n118 ,
         \i_MIPS/Register/n117 , \i_MIPS/Register/n116 ,
         \i_MIPS/Register/n115 , \i_MIPS/Register/n114 ,
         \i_MIPS/Register/n113 , \i_MIPS/Register/n112 ,
         \i_MIPS/Register/n111 , \i_MIPS/Register/n110 ,
         \i_MIPS/Register/n109 , \i_MIPS/Register/n108 ,
         \i_MIPS/Register/n107 , \i_MIPS/Register/n106 ,
         \i_MIPS/Register/n105 , \i_MIPS/Register/n104 ,
         \i_MIPS/Register/register[31][0] , \i_MIPS/Register/register[31][2] ,
         \i_MIPS/Register/register[31][3] , \i_MIPS/Register/register[31][4] ,
         \i_MIPS/Register/register[31][5] , \i_MIPS/Register/register[31][6] ,
         \i_MIPS/Register/register[31][7] , \i_MIPS/Register/register[31][8] ,
         \i_MIPS/Register/register[31][9] , \i_MIPS/Register/register[31][10] ,
         \i_MIPS/Register/register[31][11] ,
         \i_MIPS/Register/register[31][12] ,
         \i_MIPS/Register/register[31][13] ,
         \i_MIPS/Register/register[31][14] ,
         \i_MIPS/Register/register[31][15] ,
         \i_MIPS/Register/register[31][16] ,
         \i_MIPS/Register/register[31][17] ,
         \i_MIPS/Register/register[31][18] ,
         \i_MIPS/Register/register[31][20] ,
         \i_MIPS/Register/register[31][21] ,
         \i_MIPS/Register/register[31][22] ,
         \i_MIPS/Register/register[31][23] ,
         \i_MIPS/Register/register[31][24] ,
         \i_MIPS/Register/register[31][25] ,
         \i_MIPS/Register/register[31][26] ,
         \i_MIPS/Register/register[31][27] ,
         \i_MIPS/Register/register[31][28] ,
         \i_MIPS/Register/register[31][29] ,
         \i_MIPS/Register/register[31][31] , \i_MIPS/Register/register[30][0] ,
         \i_MIPS/Register/register[30][1] , \i_MIPS/Register/register[30][2] ,
         \i_MIPS/Register/register[30][3] , \i_MIPS/Register/register[30][4] ,
         \i_MIPS/Register/register[30][5] , \i_MIPS/Register/register[30][6] ,
         \i_MIPS/Register/register[30][7] , \i_MIPS/Register/register[30][8] ,
         \i_MIPS/Register/register[30][9] , \i_MIPS/Register/register[30][10] ,
         \i_MIPS/Register/register[30][11] ,
         \i_MIPS/Register/register[30][12] ,
         \i_MIPS/Register/register[30][13] ,
         \i_MIPS/Register/register[30][14] ,
         \i_MIPS/Register/register[30][15] ,
         \i_MIPS/Register/register[30][16] ,
         \i_MIPS/Register/register[30][17] ,
         \i_MIPS/Register/register[30][18] ,
         \i_MIPS/Register/register[30][19] ,
         \i_MIPS/Register/register[30][20] ,
         \i_MIPS/Register/register[30][21] ,
         \i_MIPS/Register/register[30][22] ,
         \i_MIPS/Register/register[30][23] ,
         \i_MIPS/Register/register[30][24] ,
         \i_MIPS/Register/register[30][25] ,
         \i_MIPS/Register/register[30][26] ,
         \i_MIPS/Register/register[30][27] ,
         \i_MIPS/Register/register[30][28] ,
         \i_MIPS/Register/register[30][29] ,
         \i_MIPS/Register/register[30][30] ,
         \i_MIPS/Register/register[30][31] , \i_MIPS/Register/register[29][0] ,
         \i_MIPS/Register/register[29][1] , \i_MIPS/Register/register[29][2] ,
         \i_MIPS/Register/register[29][3] , \i_MIPS/Register/register[29][4] ,
         \i_MIPS/Register/register[29][5] , \i_MIPS/Register/register[29][6] ,
         \i_MIPS/Register/register[29][7] , \i_MIPS/Register/register[29][8] ,
         \i_MIPS/Register/register[29][9] , \i_MIPS/Register/register[29][10] ,
         \i_MIPS/Register/register[29][11] ,
         \i_MIPS/Register/register[29][12] ,
         \i_MIPS/Register/register[29][13] ,
         \i_MIPS/Register/register[29][14] ,
         \i_MIPS/Register/register[29][15] ,
         \i_MIPS/Register/register[29][16] ,
         \i_MIPS/Register/register[29][17] ,
         \i_MIPS/Register/register[29][18] ,
         \i_MIPS/Register/register[29][19] ,
         \i_MIPS/Register/register[29][20] ,
         \i_MIPS/Register/register[29][21] ,
         \i_MIPS/Register/register[29][22] ,
         \i_MIPS/Register/register[29][23] ,
         \i_MIPS/Register/register[29][24] ,
         \i_MIPS/Register/register[29][25] ,
         \i_MIPS/Register/register[29][26] ,
         \i_MIPS/Register/register[29][27] ,
         \i_MIPS/Register/register[29][28] ,
         \i_MIPS/Register/register[29][29] ,
         \i_MIPS/Register/register[29][30] ,
         \i_MIPS/Register/register[29][31] , \i_MIPS/Register/register[28][0] ,
         \i_MIPS/Register/register[28][1] , \i_MIPS/Register/register[28][2] ,
         \i_MIPS/Register/register[28][3] , \i_MIPS/Register/register[28][4] ,
         \i_MIPS/Register/register[28][5] , \i_MIPS/Register/register[28][6] ,
         \i_MIPS/Register/register[28][7] , \i_MIPS/Register/register[28][8] ,
         \i_MIPS/Register/register[28][9] , \i_MIPS/Register/register[28][10] ,
         \i_MIPS/Register/register[28][11] ,
         \i_MIPS/Register/register[28][12] ,
         \i_MIPS/Register/register[28][13] ,
         \i_MIPS/Register/register[28][14] ,
         \i_MIPS/Register/register[28][15] ,
         \i_MIPS/Register/register[28][16] ,
         \i_MIPS/Register/register[28][17] ,
         \i_MIPS/Register/register[28][18] ,
         \i_MIPS/Register/register[28][19] ,
         \i_MIPS/Register/register[28][20] ,
         \i_MIPS/Register/register[28][21] ,
         \i_MIPS/Register/register[28][22] ,
         \i_MIPS/Register/register[28][23] ,
         \i_MIPS/Register/register[28][24] ,
         \i_MIPS/Register/register[28][25] ,
         \i_MIPS/Register/register[28][26] ,
         \i_MIPS/Register/register[28][27] ,
         \i_MIPS/Register/register[28][28] ,
         \i_MIPS/Register/register[28][29] ,
         \i_MIPS/Register/register[28][30] ,
         \i_MIPS/Register/register[28][31] , \i_MIPS/Register/register[27][0] ,
         \i_MIPS/Register/register[27][1] , \i_MIPS/Register/register[27][2] ,
         \i_MIPS/Register/register[27][3] , \i_MIPS/Register/register[27][4] ,
         \i_MIPS/Register/register[27][5] , \i_MIPS/Register/register[27][6] ,
         \i_MIPS/Register/register[27][7] , \i_MIPS/Register/register[27][8] ,
         \i_MIPS/Register/register[27][9] , \i_MIPS/Register/register[27][10] ,
         \i_MIPS/Register/register[27][11] ,
         \i_MIPS/Register/register[27][12] ,
         \i_MIPS/Register/register[27][13] ,
         \i_MIPS/Register/register[27][14] ,
         \i_MIPS/Register/register[27][15] ,
         \i_MIPS/Register/register[27][16] ,
         \i_MIPS/Register/register[27][17] ,
         \i_MIPS/Register/register[27][18] ,
         \i_MIPS/Register/register[27][19] ,
         \i_MIPS/Register/register[27][20] ,
         \i_MIPS/Register/register[27][21] ,
         \i_MIPS/Register/register[27][22] ,
         \i_MIPS/Register/register[27][23] ,
         \i_MIPS/Register/register[27][24] ,
         \i_MIPS/Register/register[27][25] ,
         \i_MIPS/Register/register[27][26] ,
         \i_MIPS/Register/register[27][27] ,
         \i_MIPS/Register/register[27][28] ,
         \i_MIPS/Register/register[27][29] ,
         \i_MIPS/Register/register[27][30] ,
         \i_MIPS/Register/register[27][31] , \i_MIPS/Register/register[26][0] ,
         \i_MIPS/Register/register[26][1] , \i_MIPS/Register/register[26][2] ,
         \i_MIPS/Register/register[26][3] , \i_MIPS/Register/register[26][4] ,
         \i_MIPS/Register/register[26][5] , \i_MIPS/Register/register[26][6] ,
         \i_MIPS/Register/register[26][7] , \i_MIPS/Register/register[26][8] ,
         \i_MIPS/Register/register[26][9] , \i_MIPS/Register/register[26][10] ,
         \i_MIPS/Register/register[26][11] ,
         \i_MIPS/Register/register[26][12] ,
         \i_MIPS/Register/register[26][13] ,
         \i_MIPS/Register/register[26][14] ,
         \i_MIPS/Register/register[26][15] ,
         \i_MIPS/Register/register[26][16] ,
         \i_MIPS/Register/register[26][17] ,
         \i_MIPS/Register/register[26][18] ,
         \i_MIPS/Register/register[26][19] ,
         \i_MIPS/Register/register[26][20] ,
         \i_MIPS/Register/register[26][21] ,
         \i_MIPS/Register/register[26][22] ,
         \i_MIPS/Register/register[26][23] ,
         \i_MIPS/Register/register[26][24] ,
         \i_MIPS/Register/register[26][25] ,
         \i_MIPS/Register/register[26][26] ,
         \i_MIPS/Register/register[26][27] ,
         \i_MIPS/Register/register[26][28] ,
         \i_MIPS/Register/register[26][29] ,
         \i_MIPS/Register/register[26][30] ,
         \i_MIPS/Register/register[26][31] , \i_MIPS/Register/register[25][0] ,
         \i_MIPS/Register/register[25][1] , \i_MIPS/Register/register[25][2] ,
         \i_MIPS/Register/register[25][3] , \i_MIPS/Register/register[25][4] ,
         \i_MIPS/Register/register[25][5] , \i_MIPS/Register/register[25][6] ,
         \i_MIPS/Register/register[25][7] , \i_MIPS/Register/register[25][8] ,
         \i_MIPS/Register/register[25][9] , \i_MIPS/Register/register[25][10] ,
         \i_MIPS/Register/register[25][11] ,
         \i_MIPS/Register/register[25][12] ,
         \i_MIPS/Register/register[25][13] ,
         \i_MIPS/Register/register[25][14] ,
         \i_MIPS/Register/register[25][15] ,
         \i_MIPS/Register/register[25][16] ,
         \i_MIPS/Register/register[25][17] ,
         \i_MIPS/Register/register[25][18] ,
         \i_MIPS/Register/register[25][19] ,
         \i_MIPS/Register/register[25][20] ,
         \i_MIPS/Register/register[25][21] ,
         \i_MIPS/Register/register[25][22] ,
         \i_MIPS/Register/register[25][23] ,
         \i_MIPS/Register/register[25][24] ,
         \i_MIPS/Register/register[25][25] ,
         \i_MIPS/Register/register[25][26] ,
         \i_MIPS/Register/register[25][27] ,
         \i_MIPS/Register/register[25][28] ,
         \i_MIPS/Register/register[25][29] ,
         \i_MIPS/Register/register[25][30] ,
         \i_MIPS/Register/register[25][31] , \i_MIPS/Register/register[24][0] ,
         \i_MIPS/Register/register[24][1] , \i_MIPS/Register/register[24][2] ,
         \i_MIPS/Register/register[24][3] , \i_MIPS/Register/register[24][4] ,
         \i_MIPS/Register/register[24][5] , \i_MIPS/Register/register[24][6] ,
         \i_MIPS/Register/register[24][7] , \i_MIPS/Register/register[24][8] ,
         \i_MIPS/Register/register[24][9] , \i_MIPS/Register/register[24][10] ,
         \i_MIPS/Register/register[24][11] ,
         \i_MIPS/Register/register[24][12] ,
         \i_MIPS/Register/register[24][13] ,
         \i_MIPS/Register/register[24][14] ,
         \i_MIPS/Register/register[24][15] ,
         \i_MIPS/Register/register[24][16] ,
         \i_MIPS/Register/register[24][17] ,
         \i_MIPS/Register/register[24][18] ,
         \i_MIPS/Register/register[24][19] ,
         \i_MIPS/Register/register[24][20] ,
         \i_MIPS/Register/register[24][21] ,
         \i_MIPS/Register/register[24][22] ,
         \i_MIPS/Register/register[24][23] ,
         \i_MIPS/Register/register[24][24] ,
         \i_MIPS/Register/register[24][25] ,
         \i_MIPS/Register/register[24][26] ,
         \i_MIPS/Register/register[24][27] ,
         \i_MIPS/Register/register[24][28] ,
         \i_MIPS/Register/register[24][29] ,
         \i_MIPS/Register/register[24][30] ,
         \i_MIPS/Register/register[24][31] , \i_MIPS/Register/register[23][0] ,
         \i_MIPS/Register/register[23][1] , \i_MIPS/Register/register[23][2] ,
         \i_MIPS/Register/register[23][3] , \i_MIPS/Register/register[23][4] ,
         \i_MIPS/Register/register[23][5] , \i_MIPS/Register/register[23][6] ,
         \i_MIPS/Register/register[23][7] , \i_MIPS/Register/register[23][8] ,
         \i_MIPS/Register/register[23][9] , \i_MIPS/Register/register[23][10] ,
         \i_MIPS/Register/register[23][11] ,
         \i_MIPS/Register/register[23][12] ,
         \i_MIPS/Register/register[23][13] ,
         \i_MIPS/Register/register[23][14] ,
         \i_MIPS/Register/register[23][15] ,
         \i_MIPS/Register/register[23][16] ,
         \i_MIPS/Register/register[23][17] ,
         \i_MIPS/Register/register[23][18] ,
         \i_MIPS/Register/register[23][19] ,
         \i_MIPS/Register/register[23][20] ,
         \i_MIPS/Register/register[23][21] ,
         \i_MIPS/Register/register[23][22] ,
         \i_MIPS/Register/register[23][23] ,
         \i_MIPS/Register/register[23][24] ,
         \i_MIPS/Register/register[23][25] ,
         \i_MIPS/Register/register[23][26] ,
         \i_MIPS/Register/register[23][27] ,
         \i_MIPS/Register/register[23][28] ,
         \i_MIPS/Register/register[23][29] ,
         \i_MIPS/Register/register[23][30] ,
         \i_MIPS/Register/register[23][31] , \i_MIPS/Register/register[22][0] ,
         \i_MIPS/Register/register[22][1] , \i_MIPS/Register/register[22][2] ,
         \i_MIPS/Register/register[22][3] , \i_MIPS/Register/register[22][4] ,
         \i_MIPS/Register/register[22][5] , \i_MIPS/Register/register[22][6] ,
         \i_MIPS/Register/register[22][7] , \i_MIPS/Register/register[22][8] ,
         \i_MIPS/Register/register[22][9] , \i_MIPS/Register/register[22][10] ,
         \i_MIPS/Register/register[22][11] ,
         \i_MIPS/Register/register[22][12] ,
         \i_MIPS/Register/register[22][13] ,
         \i_MIPS/Register/register[22][14] ,
         \i_MIPS/Register/register[22][15] ,
         \i_MIPS/Register/register[22][16] ,
         \i_MIPS/Register/register[22][17] ,
         \i_MIPS/Register/register[22][18] ,
         \i_MIPS/Register/register[22][19] ,
         \i_MIPS/Register/register[22][20] ,
         \i_MIPS/Register/register[22][21] ,
         \i_MIPS/Register/register[22][22] ,
         \i_MIPS/Register/register[22][23] ,
         \i_MIPS/Register/register[22][24] ,
         \i_MIPS/Register/register[22][25] ,
         \i_MIPS/Register/register[22][26] ,
         \i_MIPS/Register/register[22][27] ,
         \i_MIPS/Register/register[22][28] ,
         \i_MIPS/Register/register[22][29] ,
         \i_MIPS/Register/register[22][30] ,
         \i_MIPS/Register/register[22][31] , \i_MIPS/Register/register[21][0] ,
         \i_MIPS/Register/register[21][1] , \i_MIPS/Register/register[21][2] ,
         \i_MIPS/Register/register[21][3] , \i_MIPS/Register/register[21][4] ,
         \i_MIPS/Register/register[21][5] , \i_MIPS/Register/register[21][6] ,
         \i_MIPS/Register/register[21][7] , \i_MIPS/Register/register[21][8] ,
         \i_MIPS/Register/register[21][9] , \i_MIPS/Register/register[21][10] ,
         \i_MIPS/Register/register[21][11] ,
         \i_MIPS/Register/register[21][12] ,
         \i_MIPS/Register/register[21][13] ,
         \i_MIPS/Register/register[21][14] ,
         \i_MIPS/Register/register[21][15] ,
         \i_MIPS/Register/register[21][16] ,
         \i_MIPS/Register/register[21][17] ,
         \i_MIPS/Register/register[21][18] ,
         \i_MIPS/Register/register[21][19] ,
         \i_MIPS/Register/register[21][20] ,
         \i_MIPS/Register/register[21][21] ,
         \i_MIPS/Register/register[21][22] ,
         \i_MIPS/Register/register[21][23] ,
         \i_MIPS/Register/register[21][24] ,
         \i_MIPS/Register/register[21][25] ,
         \i_MIPS/Register/register[21][26] ,
         \i_MIPS/Register/register[21][27] ,
         \i_MIPS/Register/register[21][28] ,
         \i_MIPS/Register/register[21][29] ,
         \i_MIPS/Register/register[21][30] ,
         \i_MIPS/Register/register[21][31] , \i_MIPS/Register/register[20][0] ,
         \i_MIPS/Register/register[20][1] , \i_MIPS/Register/register[20][2] ,
         \i_MIPS/Register/register[20][3] , \i_MIPS/Register/register[20][4] ,
         \i_MIPS/Register/register[20][5] , \i_MIPS/Register/register[20][6] ,
         \i_MIPS/Register/register[20][7] , \i_MIPS/Register/register[20][8] ,
         \i_MIPS/Register/register[20][9] , \i_MIPS/Register/register[20][10] ,
         \i_MIPS/Register/register[20][11] ,
         \i_MIPS/Register/register[20][12] ,
         \i_MIPS/Register/register[20][13] ,
         \i_MIPS/Register/register[20][14] ,
         \i_MIPS/Register/register[20][15] ,
         \i_MIPS/Register/register[20][16] ,
         \i_MIPS/Register/register[20][17] ,
         \i_MIPS/Register/register[20][18] ,
         \i_MIPS/Register/register[20][19] ,
         \i_MIPS/Register/register[20][20] ,
         \i_MIPS/Register/register[20][21] ,
         \i_MIPS/Register/register[20][22] ,
         \i_MIPS/Register/register[20][23] ,
         \i_MIPS/Register/register[20][24] ,
         \i_MIPS/Register/register[20][25] ,
         \i_MIPS/Register/register[20][26] ,
         \i_MIPS/Register/register[20][27] ,
         \i_MIPS/Register/register[20][28] ,
         \i_MIPS/Register/register[20][29] ,
         \i_MIPS/Register/register[20][30] ,
         \i_MIPS/Register/register[20][31] , \i_MIPS/Register/register[19][0] ,
         \i_MIPS/Register/register[19][1] , \i_MIPS/Register/register[19][2] ,
         \i_MIPS/Register/register[19][3] , \i_MIPS/Register/register[19][4] ,
         \i_MIPS/Register/register[19][5] , \i_MIPS/Register/register[19][6] ,
         \i_MIPS/Register/register[19][7] , \i_MIPS/Register/register[19][8] ,
         \i_MIPS/Register/register[19][9] , \i_MIPS/Register/register[19][10] ,
         \i_MIPS/Register/register[19][11] ,
         \i_MIPS/Register/register[19][12] ,
         \i_MIPS/Register/register[19][13] ,
         \i_MIPS/Register/register[19][14] ,
         \i_MIPS/Register/register[19][15] ,
         \i_MIPS/Register/register[19][16] ,
         \i_MIPS/Register/register[19][17] ,
         \i_MIPS/Register/register[19][18] ,
         \i_MIPS/Register/register[19][19] ,
         \i_MIPS/Register/register[19][20] ,
         \i_MIPS/Register/register[19][21] ,
         \i_MIPS/Register/register[19][22] ,
         \i_MIPS/Register/register[19][23] ,
         \i_MIPS/Register/register[19][24] ,
         \i_MIPS/Register/register[19][25] ,
         \i_MIPS/Register/register[19][26] ,
         \i_MIPS/Register/register[19][27] ,
         \i_MIPS/Register/register[19][28] ,
         \i_MIPS/Register/register[19][29] ,
         \i_MIPS/Register/register[19][30] ,
         \i_MIPS/Register/register[19][31] , \i_MIPS/Register/register[18][0] ,
         \i_MIPS/Register/register[18][1] , \i_MIPS/Register/register[18][2] ,
         \i_MIPS/Register/register[18][3] , \i_MIPS/Register/register[18][4] ,
         \i_MIPS/Register/register[18][5] , \i_MIPS/Register/register[18][6] ,
         \i_MIPS/Register/register[18][7] , \i_MIPS/Register/register[18][8] ,
         \i_MIPS/Register/register[18][9] , \i_MIPS/Register/register[18][10] ,
         \i_MIPS/Register/register[18][11] ,
         \i_MIPS/Register/register[18][12] ,
         \i_MIPS/Register/register[18][13] ,
         \i_MIPS/Register/register[18][14] ,
         \i_MIPS/Register/register[18][15] ,
         \i_MIPS/Register/register[18][16] ,
         \i_MIPS/Register/register[18][17] ,
         \i_MIPS/Register/register[18][18] ,
         \i_MIPS/Register/register[18][19] ,
         \i_MIPS/Register/register[18][20] ,
         \i_MIPS/Register/register[18][21] ,
         \i_MIPS/Register/register[18][22] ,
         \i_MIPS/Register/register[18][23] ,
         \i_MIPS/Register/register[18][24] ,
         \i_MIPS/Register/register[18][25] ,
         \i_MIPS/Register/register[18][26] ,
         \i_MIPS/Register/register[18][27] ,
         \i_MIPS/Register/register[18][28] ,
         \i_MIPS/Register/register[18][29] ,
         \i_MIPS/Register/register[18][30] ,
         \i_MIPS/Register/register[18][31] , \i_MIPS/Register/register[17][0] ,
         \i_MIPS/Register/register[17][1] , \i_MIPS/Register/register[17][2] ,
         \i_MIPS/Register/register[17][3] , \i_MIPS/Register/register[17][4] ,
         \i_MIPS/Register/register[17][5] , \i_MIPS/Register/register[17][6] ,
         \i_MIPS/Register/register[17][7] , \i_MIPS/Register/register[17][8] ,
         \i_MIPS/Register/register[17][9] , \i_MIPS/Register/register[17][10] ,
         \i_MIPS/Register/register[17][11] ,
         \i_MIPS/Register/register[17][12] ,
         \i_MIPS/Register/register[17][13] ,
         \i_MIPS/Register/register[17][14] ,
         \i_MIPS/Register/register[17][15] ,
         \i_MIPS/Register/register[17][16] ,
         \i_MIPS/Register/register[17][17] ,
         \i_MIPS/Register/register[17][18] ,
         \i_MIPS/Register/register[17][19] ,
         \i_MIPS/Register/register[17][20] ,
         \i_MIPS/Register/register[17][21] ,
         \i_MIPS/Register/register[17][22] ,
         \i_MIPS/Register/register[17][23] ,
         \i_MIPS/Register/register[17][24] ,
         \i_MIPS/Register/register[17][25] ,
         \i_MIPS/Register/register[17][26] ,
         \i_MIPS/Register/register[17][27] ,
         \i_MIPS/Register/register[17][28] ,
         \i_MIPS/Register/register[17][29] ,
         \i_MIPS/Register/register[17][30] ,
         \i_MIPS/Register/register[17][31] , \i_MIPS/Register/register[16][0] ,
         \i_MIPS/Register/register[16][1] , \i_MIPS/Register/register[16][2] ,
         \i_MIPS/Register/register[16][3] , \i_MIPS/Register/register[16][4] ,
         \i_MIPS/Register/register[16][5] , \i_MIPS/Register/register[16][6] ,
         \i_MIPS/Register/register[16][7] , \i_MIPS/Register/register[16][8] ,
         \i_MIPS/Register/register[16][9] , \i_MIPS/Register/register[16][10] ,
         \i_MIPS/Register/register[16][11] ,
         \i_MIPS/Register/register[16][12] ,
         \i_MIPS/Register/register[16][13] ,
         \i_MIPS/Register/register[16][14] ,
         \i_MIPS/Register/register[16][15] ,
         \i_MIPS/Register/register[16][16] ,
         \i_MIPS/Register/register[16][17] ,
         \i_MIPS/Register/register[16][18] ,
         \i_MIPS/Register/register[16][19] ,
         \i_MIPS/Register/register[16][20] ,
         \i_MIPS/Register/register[16][21] ,
         \i_MIPS/Register/register[16][22] ,
         \i_MIPS/Register/register[16][23] ,
         \i_MIPS/Register/register[16][24] ,
         \i_MIPS/Register/register[16][25] ,
         \i_MIPS/Register/register[16][26] ,
         \i_MIPS/Register/register[16][27] ,
         \i_MIPS/Register/register[16][28] ,
         \i_MIPS/Register/register[16][29] ,
         \i_MIPS/Register/register[16][30] ,
         \i_MIPS/Register/register[16][31] , \i_MIPS/Register/register[15][0] ,
         \i_MIPS/Register/register[15][1] , \i_MIPS/Register/register[15][2] ,
         \i_MIPS/Register/register[15][3] , \i_MIPS/Register/register[15][4] ,
         \i_MIPS/Register/register[15][5] , \i_MIPS/Register/register[15][6] ,
         \i_MIPS/Register/register[15][7] , \i_MIPS/Register/register[15][8] ,
         \i_MIPS/Register/register[15][9] , \i_MIPS/Register/register[15][10] ,
         \i_MIPS/Register/register[15][11] ,
         \i_MIPS/Register/register[15][12] ,
         \i_MIPS/Register/register[15][13] ,
         \i_MIPS/Register/register[15][14] ,
         \i_MIPS/Register/register[15][15] ,
         \i_MIPS/Register/register[15][16] ,
         \i_MIPS/Register/register[15][17] ,
         \i_MIPS/Register/register[15][18] ,
         \i_MIPS/Register/register[15][19] ,
         \i_MIPS/Register/register[15][20] ,
         \i_MIPS/Register/register[15][21] ,
         \i_MIPS/Register/register[15][22] ,
         \i_MIPS/Register/register[15][23] ,
         \i_MIPS/Register/register[15][24] ,
         \i_MIPS/Register/register[15][25] ,
         \i_MIPS/Register/register[15][26] ,
         \i_MIPS/Register/register[15][27] ,
         \i_MIPS/Register/register[15][28] ,
         \i_MIPS/Register/register[15][29] ,
         \i_MIPS/Register/register[15][30] ,
         \i_MIPS/Register/register[15][31] , \i_MIPS/Register/register[14][0] ,
         \i_MIPS/Register/register[14][1] , \i_MIPS/Register/register[14][2] ,
         \i_MIPS/Register/register[14][3] , \i_MIPS/Register/register[14][4] ,
         \i_MIPS/Register/register[14][5] , \i_MIPS/Register/register[14][6] ,
         \i_MIPS/Register/register[14][7] , \i_MIPS/Register/register[14][8] ,
         \i_MIPS/Register/register[14][9] , \i_MIPS/Register/register[14][10] ,
         \i_MIPS/Register/register[14][11] ,
         \i_MIPS/Register/register[14][12] ,
         \i_MIPS/Register/register[14][13] ,
         \i_MIPS/Register/register[14][14] ,
         \i_MIPS/Register/register[14][15] ,
         \i_MIPS/Register/register[14][16] ,
         \i_MIPS/Register/register[14][17] ,
         \i_MIPS/Register/register[14][18] ,
         \i_MIPS/Register/register[14][19] ,
         \i_MIPS/Register/register[14][20] ,
         \i_MIPS/Register/register[14][21] ,
         \i_MIPS/Register/register[14][22] ,
         \i_MIPS/Register/register[14][23] ,
         \i_MIPS/Register/register[14][24] ,
         \i_MIPS/Register/register[14][25] ,
         \i_MIPS/Register/register[14][26] ,
         \i_MIPS/Register/register[14][27] ,
         \i_MIPS/Register/register[14][28] ,
         \i_MIPS/Register/register[14][29] ,
         \i_MIPS/Register/register[14][30] ,
         \i_MIPS/Register/register[14][31] , \i_MIPS/Register/register[13][0] ,
         \i_MIPS/Register/register[13][1] , \i_MIPS/Register/register[13][2] ,
         \i_MIPS/Register/register[13][3] , \i_MIPS/Register/register[13][4] ,
         \i_MIPS/Register/register[13][5] , \i_MIPS/Register/register[13][6] ,
         \i_MIPS/Register/register[13][7] , \i_MIPS/Register/register[13][8] ,
         \i_MIPS/Register/register[13][9] , \i_MIPS/Register/register[13][10] ,
         \i_MIPS/Register/register[13][11] ,
         \i_MIPS/Register/register[13][12] ,
         \i_MIPS/Register/register[13][13] ,
         \i_MIPS/Register/register[13][14] ,
         \i_MIPS/Register/register[13][15] ,
         \i_MIPS/Register/register[13][16] ,
         \i_MIPS/Register/register[13][17] ,
         \i_MIPS/Register/register[13][18] ,
         \i_MIPS/Register/register[13][19] ,
         \i_MIPS/Register/register[13][20] ,
         \i_MIPS/Register/register[13][21] ,
         \i_MIPS/Register/register[13][22] ,
         \i_MIPS/Register/register[13][23] ,
         \i_MIPS/Register/register[13][24] ,
         \i_MIPS/Register/register[13][25] ,
         \i_MIPS/Register/register[13][26] ,
         \i_MIPS/Register/register[13][27] ,
         \i_MIPS/Register/register[13][28] ,
         \i_MIPS/Register/register[13][29] ,
         \i_MIPS/Register/register[13][30] ,
         \i_MIPS/Register/register[13][31] , \i_MIPS/Register/register[12][0] ,
         \i_MIPS/Register/register[12][1] , \i_MIPS/Register/register[12][2] ,
         \i_MIPS/Register/register[12][3] , \i_MIPS/Register/register[12][4] ,
         \i_MIPS/Register/register[12][5] , \i_MIPS/Register/register[12][6] ,
         \i_MIPS/Register/register[12][7] , \i_MIPS/Register/register[12][8] ,
         \i_MIPS/Register/register[12][9] , \i_MIPS/Register/register[12][10] ,
         \i_MIPS/Register/register[12][11] ,
         \i_MIPS/Register/register[12][12] ,
         \i_MIPS/Register/register[12][13] ,
         \i_MIPS/Register/register[12][14] ,
         \i_MIPS/Register/register[12][15] ,
         \i_MIPS/Register/register[12][16] ,
         \i_MIPS/Register/register[12][17] ,
         \i_MIPS/Register/register[12][18] ,
         \i_MIPS/Register/register[12][19] ,
         \i_MIPS/Register/register[12][20] ,
         \i_MIPS/Register/register[12][21] ,
         \i_MIPS/Register/register[12][22] ,
         \i_MIPS/Register/register[12][23] ,
         \i_MIPS/Register/register[12][24] ,
         \i_MIPS/Register/register[12][25] ,
         \i_MIPS/Register/register[12][26] ,
         \i_MIPS/Register/register[12][27] ,
         \i_MIPS/Register/register[12][28] ,
         \i_MIPS/Register/register[12][29] ,
         \i_MIPS/Register/register[12][30] ,
         \i_MIPS/Register/register[12][31] , \i_MIPS/Register/register[11][0] ,
         \i_MIPS/Register/register[11][1] , \i_MIPS/Register/register[11][2] ,
         \i_MIPS/Register/register[11][3] , \i_MIPS/Register/register[11][4] ,
         \i_MIPS/Register/register[11][5] , \i_MIPS/Register/register[11][6] ,
         \i_MIPS/Register/register[11][7] , \i_MIPS/Register/register[11][8] ,
         \i_MIPS/Register/register[11][9] , \i_MIPS/Register/register[11][10] ,
         \i_MIPS/Register/register[11][11] ,
         \i_MIPS/Register/register[11][12] ,
         \i_MIPS/Register/register[11][13] ,
         \i_MIPS/Register/register[11][14] ,
         \i_MIPS/Register/register[11][15] ,
         \i_MIPS/Register/register[11][16] ,
         \i_MIPS/Register/register[11][17] ,
         \i_MIPS/Register/register[11][18] ,
         \i_MIPS/Register/register[11][19] ,
         \i_MIPS/Register/register[11][20] ,
         \i_MIPS/Register/register[11][21] ,
         \i_MIPS/Register/register[11][22] ,
         \i_MIPS/Register/register[11][23] ,
         \i_MIPS/Register/register[11][24] ,
         \i_MIPS/Register/register[11][25] ,
         \i_MIPS/Register/register[11][26] ,
         \i_MIPS/Register/register[11][27] ,
         \i_MIPS/Register/register[11][28] ,
         \i_MIPS/Register/register[11][29] ,
         \i_MIPS/Register/register[11][30] ,
         \i_MIPS/Register/register[11][31] , \i_MIPS/Register/register[10][0] ,
         \i_MIPS/Register/register[10][1] , \i_MIPS/Register/register[10][2] ,
         \i_MIPS/Register/register[10][3] , \i_MIPS/Register/register[10][4] ,
         \i_MIPS/Register/register[10][5] , \i_MIPS/Register/register[10][6] ,
         \i_MIPS/Register/register[10][7] , \i_MIPS/Register/register[10][8] ,
         \i_MIPS/Register/register[10][9] , \i_MIPS/Register/register[10][10] ,
         \i_MIPS/Register/register[10][11] ,
         \i_MIPS/Register/register[10][12] ,
         \i_MIPS/Register/register[10][13] ,
         \i_MIPS/Register/register[10][14] ,
         \i_MIPS/Register/register[10][15] ,
         \i_MIPS/Register/register[10][16] ,
         \i_MIPS/Register/register[10][17] ,
         \i_MIPS/Register/register[10][18] ,
         \i_MIPS/Register/register[10][19] ,
         \i_MIPS/Register/register[10][20] ,
         \i_MIPS/Register/register[10][21] ,
         \i_MIPS/Register/register[10][22] ,
         \i_MIPS/Register/register[10][23] ,
         \i_MIPS/Register/register[10][24] ,
         \i_MIPS/Register/register[10][25] ,
         \i_MIPS/Register/register[10][26] ,
         \i_MIPS/Register/register[10][27] ,
         \i_MIPS/Register/register[10][28] ,
         \i_MIPS/Register/register[10][29] ,
         \i_MIPS/Register/register[10][30] ,
         \i_MIPS/Register/register[10][31] , \i_MIPS/Register/register[9][0] ,
         \i_MIPS/Register/register[9][1] , \i_MIPS/Register/register[9][2] ,
         \i_MIPS/Register/register[9][3] , \i_MIPS/Register/register[9][4] ,
         \i_MIPS/Register/register[9][5] , \i_MIPS/Register/register[9][6] ,
         \i_MIPS/Register/register[9][7] , \i_MIPS/Register/register[9][8] ,
         \i_MIPS/Register/register[9][9] , \i_MIPS/Register/register[9][10] ,
         \i_MIPS/Register/register[9][11] , \i_MIPS/Register/register[9][12] ,
         \i_MIPS/Register/register[9][13] , \i_MIPS/Register/register[9][14] ,
         \i_MIPS/Register/register[9][15] , \i_MIPS/Register/register[9][16] ,
         \i_MIPS/Register/register[9][17] , \i_MIPS/Register/register[9][18] ,
         \i_MIPS/Register/register[9][19] , \i_MIPS/Register/register[9][20] ,
         \i_MIPS/Register/register[9][21] , \i_MIPS/Register/register[9][22] ,
         \i_MIPS/Register/register[9][23] , \i_MIPS/Register/register[9][24] ,
         \i_MIPS/Register/register[9][25] , \i_MIPS/Register/register[9][26] ,
         \i_MIPS/Register/register[9][27] , \i_MIPS/Register/register[9][28] ,
         \i_MIPS/Register/register[9][29] , \i_MIPS/Register/register[9][30] ,
         \i_MIPS/Register/register[9][31] , \i_MIPS/Register/register[8][0] ,
         \i_MIPS/Register/register[8][1] , \i_MIPS/Register/register[8][2] ,
         \i_MIPS/Register/register[8][3] , \i_MIPS/Register/register[8][4] ,
         \i_MIPS/Register/register[8][5] , \i_MIPS/Register/register[8][6] ,
         \i_MIPS/Register/register[8][7] , \i_MIPS/Register/register[8][8] ,
         \i_MIPS/Register/register[8][9] , \i_MIPS/Register/register[8][10] ,
         \i_MIPS/Register/register[8][11] , \i_MIPS/Register/register[8][12] ,
         \i_MIPS/Register/register[8][13] , \i_MIPS/Register/register[8][14] ,
         \i_MIPS/Register/register[8][15] , \i_MIPS/Register/register[8][16] ,
         \i_MIPS/Register/register[8][17] , \i_MIPS/Register/register[8][18] ,
         \i_MIPS/Register/register[8][19] , \i_MIPS/Register/register[8][20] ,
         \i_MIPS/Register/register[8][21] , \i_MIPS/Register/register[8][22] ,
         \i_MIPS/Register/register[8][23] , \i_MIPS/Register/register[8][24] ,
         \i_MIPS/Register/register[8][25] , \i_MIPS/Register/register[8][26] ,
         \i_MIPS/Register/register[8][27] , \i_MIPS/Register/register[8][28] ,
         \i_MIPS/Register/register[8][29] , \i_MIPS/Register/register[8][30] ,
         \i_MIPS/Register/register[8][31] , \i_MIPS/Register/register[7][0] ,
         \i_MIPS/Register/register[7][1] , \i_MIPS/Register/register[7][2] ,
         \i_MIPS/Register/register[7][3] , \i_MIPS/Register/register[7][4] ,
         \i_MIPS/Register/register[7][5] , \i_MIPS/Register/register[7][6] ,
         \i_MIPS/Register/register[7][7] , \i_MIPS/Register/register[7][8] ,
         \i_MIPS/Register/register[7][9] , \i_MIPS/Register/register[7][10] ,
         \i_MIPS/Register/register[7][11] , \i_MIPS/Register/register[7][12] ,
         \i_MIPS/Register/register[7][13] , \i_MIPS/Register/register[7][14] ,
         \i_MIPS/Register/register[7][15] , \i_MIPS/Register/register[7][16] ,
         \i_MIPS/Register/register[7][17] , \i_MIPS/Register/register[7][18] ,
         \i_MIPS/Register/register[7][19] , \i_MIPS/Register/register[7][20] ,
         \i_MIPS/Register/register[7][21] , \i_MIPS/Register/register[7][22] ,
         \i_MIPS/Register/register[7][23] , \i_MIPS/Register/register[7][24] ,
         \i_MIPS/Register/register[7][25] , \i_MIPS/Register/register[7][26] ,
         \i_MIPS/Register/register[7][27] , \i_MIPS/Register/register[7][28] ,
         \i_MIPS/Register/register[7][29] , \i_MIPS/Register/register[7][30] ,
         \i_MIPS/Register/register[7][31] , \i_MIPS/Register/register[6][0] ,
         \i_MIPS/Register/register[6][1] , \i_MIPS/Register/register[6][2] ,
         \i_MIPS/Register/register[6][3] , \i_MIPS/Register/register[6][4] ,
         \i_MIPS/Register/register[6][5] , \i_MIPS/Register/register[6][6] ,
         \i_MIPS/Register/register[6][7] , \i_MIPS/Register/register[6][8] ,
         \i_MIPS/Register/register[6][9] , \i_MIPS/Register/register[6][10] ,
         \i_MIPS/Register/register[6][11] , \i_MIPS/Register/register[6][12] ,
         \i_MIPS/Register/register[6][13] , \i_MIPS/Register/register[6][14] ,
         \i_MIPS/Register/register[6][15] , \i_MIPS/Register/register[6][16] ,
         \i_MIPS/Register/register[6][17] , \i_MIPS/Register/register[6][18] ,
         \i_MIPS/Register/register[6][19] , \i_MIPS/Register/register[6][20] ,
         \i_MIPS/Register/register[6][21] , \i_MIPS/Register/register[6][22] ,
         \i_MIPS/Register/register[6][23] , \i_MIPS/Register/register[6][24] ,
         \i_MIPS/Register/register[6][25] , \i_MIPS/Register/register[6][26] ,
         \i_MIPS/Register/register[6][27] , \i_MIPS/Register/register[6][28] ,
         \i_MIPS/Register/register[6][29] , \i_MIPS/Register/register[6][30] ,
         \i_MIPS/Register/register[6][31] , \i_MIPS/Register/register[5][0] ,
         \i_MIPS/Register/register[5][1] , \i_MIPS/Register/register[5][2] ,
         \i_MIPS/Register/register[5][3] , \i_MIPS/Register/register[5][4] ,
         \i_MIPS/Register/register[5][5] , \i_MIPS/Register/register[5][6] ,
         \i_MIPS/Register/register[5][7] , \i_MIPS/Register/register[5][8] ,
         \i_MIPS/Register/register[5][9] , \i_MIPS/Register/register[5][10] ,
         \i_MIPS/Register/register[5][11] , \i_MIPS/Register/register[5][12] ,
         \i_MIPS/Register/register[5][13] , \i_MIPS/Register/register[5][14] ,
         \i_MIPS/Register/register[5][15] , \i_MIPS/Register/register[5][16] ,
         \i_MIPS/Register/register[5][17] , \i_MIPS/Register/register[5][18] ,
         \i_MIPS/Register/register[5][19] , \i_MIPS/Register/register[5][20] ,
         \i_MIPS/Register/register[5][21] , \i_MIPS/Register/register[5][22] ,
         \i_MIPS/Register/register[5][23] , \i_MIPS/Register/register[5][24] ,
         \i_MIPS/Register/register[5][25] , \i_MIPS/Register/register[5][26] ,
         \i_MIPS/Register/register[5][27] , \i_MIPS/Register/register[5][28] ,
         \i_MIPS/Register/register[5][29] , \i_MIPS/Register/register[5][30] ,
         \i_MIPS/Register/register[5][31] , \i_MIPS/Register/register[4][0] ,
         \i_MIPS/Register/register[4][1] , \i_MIPS/Register/register[4][2] ,
         \i_MIPS/Register/register[4][3] , \i_MIPS/Register/register[4][4] ,
         \i_MIPS/Register/register[4][5] , \i_MIPS/Register/register[4][6] ,
         \i_MIPS/Register/register[4][7] , \i_MIPS/Register/register[4][8] ,
         \i_MIPS/Register/register[4][9] , \i_MIPS/Register/register[4][10] ,
         \i_MIPS/Register/register[4][11] , \i_MIPS/Register/register[4][12] ,
         \i_MIPS/Register/register[4][13] , \i_MIPS/Register/register[4][14] ,
         \i_MIPS/Register/register[4][15] , \i_MIPS/Register/register[4][16] ,
         \i_MIPS/Register/register[4][17] , \i_MIPS/Register/register[4][18] ,
         \i_MIPS/Register/register[4][19] , \i_MIPS/Register/register[4][20] ,
         \i_MIPS/Register/register[4][21] , \i_MIPS/Register/register[4][22] ,
         \i_MIPS/Register/register[4][23] , \i_MIPS/Register/register[4][24] ,
         \i_MIPS/Register/register[4][25] , \i_MIPS/Register/register[4][26] ,
         \i_MIPS/Register/register[4][27] , \i_MIPS/Register/register[4][28] ,
         \i_MIPS/Register/register[4][29] , \i_MIPS/Register/register[4][30] ,
         \i_MIPS/Register/register[4][31] , \i_MIPS/Register/register[3][0] ,
         \i_MIPS/Register/register[3][1] , \i_MIPS/Register/register[3][2] ,
         \i_MIPS/Register/register[3][3] , \i_MIPS/Register/register[3][4] ,
         \i_MIPS/Register/register[3][5] , \i_MIPS/Register/register[3][6] ,
         \i_MIPS/Register/register[3][7] , \i_MIPS/Register/register[3][8] ,
         \i_MIPS/Register/register[3][9] , \i_MIPS/Register/register[3][10] ,
         \i_MIPS/Register/register[3][11] , \i_MIPS/Register/register[3][12] ,
         \i_MIPS/Register/register[3][13] , \i_MIPS/Register/register[3][14] ,
         \i_MIPS/Register/register[3][15] , \i_MIPS/Register/register[3][16] ,
         \i_MIPS/Register/register[3][17] , \i_MIPS/Register/register[3][18] ,
         \i_MIPS/Register/register[3][19] , \i_MIPS/Register/register[3][20] ,
         \i_MIPS/Register/register[3][21] , \i_MIPS/Register/register[3][22] ,
         \i_MIPS/Register/register[3][23] , \i_MIPS/Register/register[3][24] ,
         \i_MIPS/Register/register[3][25] , \i_MIPS/Register/register[3][26] ,
         \i_MIPS/Register/register[3][27] , \i_MIPS/Register/register[3][28] ,
         \i_MIPS/Register/register[3][29] , \i_MIPS/Register/register[3][30] ,
         \i_MIPS/Register/register[3][31] , \i_MIPS/Register/register[2][0] ,
         \i_MIPS/Register/register[2][1] , \i_MIPS/Register/register[2][2] ,
         \i_MIPS/Register/register[2][3] , \i_MIPS/Register/register[2][4] ,
         \i_MIPS/Register/register[2][5] , \i_MIPS/Register/register[2][6] ,
         \i_MIPS/Register/register[2][7] , \i_MIPS/Register/register[2][8] ,
         \i_MIPS/Register/register[2][9] , \i_MIPS/Register/register[2][10] ,
         \i_MIPS/Register/register[2][11] , \i_MIPS/Register/register[2][12] ,
         \i_MIPS/Register/register[2][13] , \i_MIPS/Register/register[2][14] ,
         \i_MIPS/Register/register[2][15] , \i_MIPS/Register/register[2][16] ,
         \i_MIPS/Register/register[2][17] , \i_MIPS/Register/register[2][18] ,
         \i_MIPS/Register/register[2][19] , \i_MIPS/Register/register[2][20] ,
         \i_MIPS/Register/register[2][21] , \i_MIPS/Register/register[2][22] ,
         \i_MIPS/Register/register[2][23] , \i_MIPS/Register/register[2][24] ,
         \i_MIPS/Register/register[2][25] , \i_MIPS/Register/register[2][26] ,
         \i_MIPS/Register/register[2][27] , \i_MIPS/Register/register[2][28] ,
         \i_MIPS/Register/register[2][29] , \i_MIPS/Register/register[2][30] ,
         \i_MIPS/Register/register[2][31] , \i_MIPS/Register/register[1][0] ,
         \i_MIPS/Register/register[1][1] , \i_MIPS/Register/register[1][2] ,
         \i_MIPS/Register/register[1][3] , \i_MIPS/Register/register[1][4] ,
         \i_MIPS/Register/register[1][5] , \i_MIPS/Register/register[1][6] ,
         \i_MIPS/Register/register[1][7] , \i_MIPS/Register/register[1][8] ,
         \i_MIPS/Register/register[1][9] , \i_MIPS/Register/register[1][10] ,
         \i_MIPS/Register/register[1][11] , \i_MIPS/Register/register[1][12] ,
         \i_MIPS/Register/register[1][13] , \i_MIPS/Register/register[1][14] ,
         \i_MIPS/Register/register[1][15] , \i_MIPS/Register/register[1][16] ,
         \i_MIPS/Register/register[1][17] , \i_MIPS/Register/register[1][18] ,
         \i_MIPS/Register/register[1][19] , \i_MIPS/Register/register[1][20] ,
         \i_MIPS/Register/register[1][21] , \i_MIPS/Register/register[1][22] ,
         \i_MIPS/Register/register[1][23] , \i_MIPS/Register/register[1][24] ,
         \i_MIPS/Register/register[1][25] , \i_MIPS/Register/register[1][26] ,
         \i_MIPS/Register/register[1][27] , \i_MIPS/Register/register[1][28] ,
         \i_MIPS/Register/register[1][29] , \i_MIPS/Register/register[1][30] ,
         \i_MIPS/Register/register[1][31] , \i_MIPS/Register/register[0][0] ,
         \i_MIPS/Register/register[0][1] , \i_MIPS/Register/register[0][2] ,
         \i_MIPS/Register/register[0][3] , \i_MIPS/Register/register[0][4] ,
         \i_MIPS/Register/register[0][5] , \i_MIPS/Register/register[0][6] ,
         \i_MIPS/Register/register[0][7] , \i_MIPS/Register/register[0][8] ,
         \i_MIPS/Register/register[0][9] , \i_MIPS/Register/register[0][10] ,
         \i_MIPS/Register/register[0][11] , \i_MIPS/Register/register[0][12] ,
         \i_MIPS/Register/register[0][13] , \i_MIPS/Register/register[0][14] ,
         \i_MIPS/Register/register[0][15] , \i_MIPS/Register/register[0][16] ,
         \i_MIPS/Register/register[0][17] , \i_MIPS/Register/register[0][18] ,
         \i_MIPS/Register/register[0][19] , \i_MIPS/Register/register[0][20] ,
         \i_MIPS/Register/register[0][21] , \i_MIPS/Register/register[0][22] ,
         \i_MIPS/Register/register[0][23] , \i_MIPS/Register/register[0][24] ,
         \i_MIPS/Register/register[0][25] , \i_MIPS/Register/register[0][26] ,
         \i_MIPS/Register/register[0][27] , \i_MIPS/Register/register[0][28] ,
         \i_MIPS/Register/register[0][29] , \i_MIPS/Register/register[0][30] ,
         \i_MIPS/Register/register[0][31] , \i_MIPS/Control_ID/n15 ,
         \i_MIPS/Control_ID/n12 , \i_MIPS/Control_ID/n10 ,
         \i_MIPS/Hazard_detection/n13 , \i_MIPS/Hazard_detection/n12 ,
         \i_MIPS/Hazard_detection/n11 , \i_MIPS/Hazard_detection/n10 ,
         \i_MIPS/Hazard_detection/n9 , \i_MIPS/Hazard_detection/n8 ,
         \i_MIPS/Hazard_detection/n7 , \i_MIPS/Hazard_detection/n4 ,
         \i_MIPS/forward_unit/n25 , \i_MIPS/forward_unit/n10 ,
         \i_MIPS/ALU_Control/n20 , \i_MIPS/ALU_Control/n15 ,
         \i_MIPS/ALU_Control/n11 , \i_MIPS/ALU_Control/n10 , \i_MIPS/ALU/N303 ,
         \I_cache/cache[7][0] , \I_cache/cache[7][1] , \I_cache/cache[7][2] ,
         \I_cache/cache[7][3] , \I_cache/cache[7][4] , \I_cache/cache[7][5] ,
         \I_cache/cache[7][6] , \I_cache/cache[7][7] , \I_cache/cache[7][8] ,
         \I_cache/cache[7][9] , \I_cache/cache[7][10] , \I_cache/cache[7][11] ,
         \I_cache/cache[7][12] , \I_cache/cache[7][13] ,
         \I_cache/cache[7][14] , \I_cache/cache[7][15] ,
         \I_cache/cache[7][16] , \I_cache/cache[7][17] ,
         \I_cache/cache[7][18] , \I_cache/cache[7][19] ,
         \I_cache/cache[7][20] , \I_cache/cache[7][21] ,
         \I_cache/cache[7][22] , \I_cache/cache[7][23] ,
         \I_cache/cache[7][24] , \I_cache/cache[7][25] ,
         \I_cache/cache[7][26] , \I_cache/cache[7][27] ,
         \I_cache/cache[7][28] , \I_cache/cache[7][29] ,
         \I_cache/cache[7][30] , \I_cache/cache[7][31] ,
         \I_cache/cache[7][32] , \I_cache/cache[7][33] ,
         \I_cache/cache[7][34] , \I_cache/cache[7][35] ,
         \I_cache/cache[7][36] , \I_cache/cache[7][37] ,
         \I_cache/cache[7][38] , \I_cache/cache[7][39] ,
         \I_cache/cache[7][40] , \I_cache/cache[7][41] ,
         \I_cache/cache[7][42] , \I_cache/cache[7][43] ,
         \I_cache/cache[7][44] , \I_cache/cache[7][45] ,
         \I_cache/cache[7][46] , \I_cache/cache[7][47] ,
         \I_cache/cache[7][48] , \I_cache/cache[7][49] ,
         \I_cache/cache[7][50] , \I_cache/cache[7][51] ,
         \I_cache/cache[7][52] , \I_cache/cache[7][53] ,
         \I_cache/cache[7][54] , \I_cache/cache[7][55] ,
         \I_cache/cache[7][56] , \I_cache/cache[7][57] ,
         \I_cache/cache[7][58] , \I_cache/cache[7][59] ,
         \I_cache/cache[7][60] , \I_cache/cache[7][61] ,
         \I_cache/cache[7][62] , \I_cache/cache[7][63] ,
         \I_cache/cache[7][64] , \I_cache/cache[7][65] ,
         \I_cache/cache[7][66] , \I_cache/cache[7][67] ,
         \I_cache/cache[7][68] , \I_cache/cache[7][69] ,
         \I_cache/cache[7][70] , \I_cache/cache[7][71] ,
         \I_cache/cache[7][72] , \I_cache/cache[7][73] ,
         \I_cache/cache[7][74] , \I_cache/cache[7][75] ,
         \I_cache/cache[7][76] , \I_cache/cache[7][77] ,
         \I_cache/cache[7][78] , \I_cache/cache[7][79] ,
         \I_cache/cache[7][80] , \I_cache/cache[7][81] ,
         \I_cache/cache[7][82] , \I_cache/cache[7][83] ,
         \I_cache/cache[7][84] , \I_cache/cache[7][85] ,
         \I_cache/cache[7][86] , \I_cache/cache[7][87] ,
         \I_cache/cache[7][88] , \I_cache/cache[7][89] ,
         \I_cache/cache[7][90] , \I_cache/cache[7][91] ,
         \I_cache/cache[7][92] , \I_cache/cache[7][93] ,
         \I_cache/cache[7][94] , \I_cache/cache[7][95] ,
         \I_cache/cache[7][96] , \I_cache/cache[7][97] ,
         \I_cache/cache[7][98] , \I_cache/cache[7][99] ,
         \I_cache/cache[7][100] , \I_cache/cache[7][101] ,
         \I_cache/cache[7][102] , \I_cache/cache[7][103] ,
         \I_cache/cache[7][104] , \I_cache/cache[7][105] ,
         \I_cache/cache[7][106] , \I_cache/cache[7][107] ,
         \I_cache/cache[7][108] , \I_cache/cache[7][109] ,
         \I_cache/cache[7][110] , \I_cache/cache[7][111] ,
         \I_cache/cache[7][112] , \I_cache/cache[7][113] ,
         \I_cache/cache[7][114] , \I_cache/cache[7][115] ,
         \I_cache/cache[7][116] , \I_cache/cache[7][117] ,
         \I_cache/cache[7][118] , \I_cache/cache[7][119] ,
         \I_cache/cache[7][120] , \I_cache/cache[7][121] ,
         \I_cache/cache[7][122] , \I_cache/cache[7][123] ,
         \I_cache/cache[7][124] , \I_cache/cache[7][125] ,
         \I_cache/cache[7][126] , \I_cache/cache[7][127] ,
         \I_cache/cache[7][128] , \I_cache/cache[7][129] ,
         \I_cache/cache[7][130] , \I_cache/cache[7][131] ,
         \I_cache/cache[7][132] , \I_cache/cache[7][133] ,
         \I_cache/cache[7][134] , \I_cache/cache[7][135] ,
         \I_cache/cache[7][136] , \I_cache/cache[7][137] ,
         \I_cache/cache[7][138] , \I_cache/cache[7][139] ,
         \I_cache/cache[7][140] , \I_cache/cache[7][141] ,
         \I_cache/cache[7][142] , \I_cache/cache[7][143] ,
         \I_cache/cache[7][144] , \I_cache/cache[7][145] ,
         \I_cache/cache[7][146] , \I_cache/cache[7][147] ,
         \I_cache/cache[7][148] , \I_cache/cache[7][149] ,
         \I_cache/cache[7][150] , \I_cache/cache[7][151] ,
         \I_cache/cache[7][152] , \I_cache/cache[7][153] ,
         \I_cache/cache[7][154] , \I_cache/cache[6][0] , \I_cache/cache[6][1] ,
         \I_cache/cache[6][2] , \I_cache/cache[6][3] , \I_cache/cache[6][4] ,
         \I_cache/cache[6][5] , \I_cache/cache[6][6] , \I_cache/cache[6][7] ,
         \I_cache/cache[6][8] , \I_cache/cache[6][9] , \I_cache/cache[6][10] ,
         \I_cache/cache[6][11] , \I_cache/cache[6][12] ,
         \I_cache/cache[6][13] , \I_cache/cache[6][14] ,
         \I_cache/cache[6][15] , \I_cache/cache[6][16] ,
         \I_cache/cache[6][17] , \I_cache/cache[6][18] ,
         \I_cache/cache[6][19] , \I_cache/cache[6][20] ,
         \I_cache/cache[6][21] , \I_cache/cache[6][22] ,
         \I_cache/cache[6][23] , \I_cache/cache[6][24] ,
         \I_cache/cache[6][25] , \I_cache/cache[6][26] ,
         \I_cache/cache[6][27] , \I_cache/cache[6][28] ,
         \I_cache/cache[6][29] , \I_cache/cache[6][30] ,
         \I_cache/cache[6][31] , \I_cache/cache[6][32] ,
         \I_cache/cache[6][33] , \I_cache/cache[6][34] ,
         \I_cache/cache[6][35] , \I_cache/cache[6][36] ,
         \I_cache/cache[6][37] , \I_cache/cache[6][38] ,
         \I_cache/cache[6][39] , \I_cache/cache[6][40] ,
         \I_cache/cache[6][41] , \I_cache/cache[6][42] ,
         \I_cache/cache[6][43] , \I_cache/cache[6][44] ,
         \I_cache/cache[6][45] , \I_cache/cache[6][46] ,
         \I_cache/cache[6][47] , \I_cache/cache[6][48] ,
         \I_cache/cache[6][49] , \I_cache/cache[6][50] ,
         \I_cache/cache[6][51] , \I_cache/cache[6][52] ,
         \I_cache/cache[6][53] , \I_cache/cache[6][54] ,
         \I_cache/cache[6][55] , \I_cache/cache[6][56] ,
         \I_cache/cache[6][57] , \I_cache/cache[6][58] ,
         \I_cache/cache[6][59] , \I_cache/cache[6][60] ,
         \I_cache/cache[6][61] , \I_cache/cache[6][62] ,
         \I_cache/cache[6][63] , \I_cache/cache[6][64] ,
         \I_cache/cache[6][65] , \I_cache/cache[6][66] ,
         \I_cache/cache[6][67] , \I_cache/cache[6][68] ,
         \I_cache/cache[6][69] , \I_cache/cache[6][70] ,
         \I_cache/cache[6][71] , \I_cache/cache[6][72] ,
         \I_cache/cache[6][73] , \I_cache/cache[6][74] ,
         \I_cache/cache[6][75] , \I_cache/cache[6][76] ,
         \I_cache/cache[6][77] , \I_cache/cache[6][78] ,
         \I_cache/cache[6][79] , \I_cache/cache[6][80] ,
         \I_cache/cache[6][81] , \I_cache/cache[6][82] ,
         \I_cache/cache[6][83] , \I_cache/cache[6][84] ,
         \I_cache/cache[6][85] , \I_cache/cache[6][86] ,
         \I_cache/cache[6][87] , \I_cache/cache[6][88] ,
         \I_cache/cache[6][89] , \I_cache/cache[6][90] ,
         \I_cache/cache[6][91] , \I_cache/cache[6][92] ,
         \I_cache/cache[6][93] , \I_cache/cache[6][94] ,
         \I_cache/cache[6][95] , \I_cache/cache[6][96] ,
         \I_cache/cache[6][97] , \I_cache/cache[6][98] ,
         \I_cache/cache[6][99] , \I_cache/cache[6][100] ,
         \I_cache/cache[6][101] , \I_cache/cache[6][102] ,
         \I_cache/cache[6][103] , \I_cache/cache[6][104] ,
         \I_cache/cache[6][105] , \I_cache/cache[6][106] ,
         \I_cache/cache[6][107] , \I_cache/cache[6][108] ,
         \I_cache/cache[6][109] , \I_cache/cache[6][110] ,
         \I_cache/cache[6][111] , \I_cache/cache[6][112] ,
         \I_cache/cache[6][113] , \I_cache/cache[6][114] ,
         \I_cache/cache[6][115] , \I_cache/cache[6][116] ,
         \I_cache/cache[6][117] , \I_cache/cache[6][118] ,
         \I_cache/cache[6][119] , \I_cache/cache[6][120] ,
         \I_cache/cache[6][121] , \I_cache/cache[6][122] ,
         \I_cache/cache[6][123] , \I_cache/cache[6][124] ,
         \I_cache/cache[6][125] , \I_cache/cache[6][126] ,
         \I_cache/cache[6][127] , \I_cache/cache[6][128] ,
         \I_cache/cache[6][129] , \I_cache/cache[6][130] ,
         \I_cache/cache[6][131] , \I_cache/cache[6][132] ,
         \I_cache/cache[6][133] , \I_cache/cache[6][134] ,
         \I_cache/cache[6][135] , \I_cache/cache[6][136] ,
         \I_cache/cache[6][137] , \I_cache/cache[6][138] ,
         \I_cache/cache[6][139] , \I_cache/cache[6][140] ,
         \I_cache/cache[6][141] , \I_cache/cache[6][142] ,
         \I_cache/cache[6][143] , \I_cache/cache[6][144] ,
         \I_cache/cache[6][145] , \I_cache/cache[6][146] ,
         \I_cache/cache[6][147] , \I_cache/cache[6][148] ,
         \I_cache/cache[6][149] , \I_cache/cache[6][150] ,
         \I_cache/cache[6][151] , \I_cache/cache[6][152] ,
         \I_cache/cache[6][153] , \I_cache/cache[6][154] ,
         \I_cache/cache[5][0] , \I_cache/cache[5][1] , \I_cache/cache[5][2] ,
         \I_cache/cache[5][3] , \I_cache/cache[5][4] , \I_cache/cache[5][5] ,
         \I_cache/cache[5][6] , \I_cache/cache[5][7] , \I_cache/cache[5][8] ,
         \I_cache/cache[5][9] , \I_cache/cache[5][10] , \I_cache/cache[5][11] ,
         \I_cache/cache[5][12] , \I_cache/cache[5][13] ,
         \I_cache/cache[5][14] , \I_cache/cache[5][15] ,
         \I_cache/cache[5][16] , \I_cache/cache[5][17] ,
         \I_cache/cache[5][18] , \I_cache/cache[5][19] ,
         \I_cache/cache[5][20] , \I_cache/cache[5][21] ,
         \I_cache/cache[5][22] , \I_cache/cache[5][23] ,
         \I_cache/cache[5][24] , \I_cache/cache[5][25] ,
         \I_cache/cache[5][26] , \I_cache/cache[5][27] ,
         \I_cache/cache[5][28] , \I_cache/cache[5][29] ,
         \I_cache/cache[5][30] , \I_cache/cache[5][31] ,
         \I_cache/cache[5][32] , \I_cache/cache[5][33] ,
         \I_cache/cache[5][34] , \I_cache/cache[5][35] ,
         \I_cache/cache[5][36] , \I_cache/cache[5][37] ,
         \I_cache/cache[5][38] , \I_cache/cache[5][39] ,
         \I_cache/cache[5][40] , \I_cache/cache[5][41] ,
         \I_cache/cache[5][42] , \I_cache/cache[5][43] ,
         \I_cache/cache[5][44] , \I_cache/cache[5][45] ,
         \I_cache/cache[5][46] , \I_cache/cache[5][47] ,
         \I_cache/cache[5][48] , \I_cache/cache[5][49] ,
         \I_cache/cache[5][50] , \I_cache/cache[5][51] ,
         \I_cache/cache[5][52] , \I_cache/cache[5][53] ,
         \I_cache/cache[5][54] , \I_cache/cache[5][55] ,
         \I_cache/cache[5][56] , \I_cache/cache[5][57] ,
         \I_cache/cache[5][58] , \I_cache/cache[5][59] ,
         \I_cache/cache[5][60] , \I_cache/cache[5][61] ,
         \I_cache/cache[5][62] , \I_cache/cache[5][63] ,
         \I_cache/cache[5][64] , \I_cache/cache[5][65] ,
         \I_cache/cache[5][66] , \I_cache/cache[5][67] ,
         \I_cache/cache[5][68] , \I_cache/cache[5][69] ,
         \I_cache/cache[5][70] , \I_cache/cache[5][71] ,
         \I_cache/cache[5][72] , \I_cache/cache[5][73] ,
         \I_cache/cache[5][74] , \I_cache/cache[5][75] ,
         \I_cache/cache[5][76] , \I_cache/cache[5][77] ,
         \I_cache/cache[5][78] , \I_cache/cache[5][79] ,
         \I_cache/cache[5][80] , \I_cache/cache[5][81] ,
         \I_cache/cache[5][82] , \I_cache/cache[5][83] ,
         \I_cache/cache[5][84] , \I_cache/cache[5][85] ,
         \I_cache/cache[5][86] , \I_cache/cache[5][87] ,
         \I_cache/cache[5][88] , \I_cache/cache[5][89] ,
         \I_cache/cache[5][90] , \I_cache/cache[5][91] ,
         \I_cache/cache[5][92] , \I_cache/cache[5][93] ,
         \I_cache/cache[5][94] , \I_cache/cache[5][95] ,
         \I_cache/cache[5][96] , \I_cache/cache[5][97] ,
         \I_cache/cache[5][98] , \I_cache/cache[5][99] ,
         \I_cache/cache[5][100] , \I_cache/cache[5][101] ,
         \I_cache/cache[5][102] , \I_cache/cache[5][103] ,
         \I_cache/cache[5][104] , \I_cache/cache[5][105] ,
         \I_cache/cache[5][106] , \I_cache/cache[5][107] ,
         \I_cache/cache[5][108] , \I_cache/cache[5][109] ,
         \I_cache/cache[5][110] , \I_cache/cache[5][111] ,
         \I_cache/cache[5][112] , \I_cache/cache[5][113] ,
         \I_cache/cache[5][114] , \I_cache/cache[5][115] ,
         \I_cache/cache[5][116] , \I_cache/cache[5][117] ,
         \I_cache/cache[5][118] , \I_cache/cache[5][119] ,
         \I_cache/cache[5][120] , \I_cache/cache[5][121] ,
         \I_cache/cache[5][122] , \I_cache/cache[5][123] ,
         \I_cache/cache[5][124] , \I_cache/cache[5][125] ,
         \I_cache/cache[5][126] , \I_cache/cache[5][127] ,
         \I_cache/cache[5][128] , \I_cache/cache[5][129] ,
         \I_cache/cache[5][130] , \I_cache/cache[5][131] ,
         \I_cache/cache[5][132] , \I_cache/cache[5][133] ,
         \I_cache/cache[5][134] , \I_cache/cache[5][135] ,
         \I_cache/cache[5][136] , \I_cache/cache[5][137] ,
         \I_cache/cache[5][138] , \I_cache/cache[5][139] ,
         \I_cache/cache[5][140] , \I_cache/cache[5][141] ,
         \I_cache/cache[5][142] , \I_cache/cache[5][143] ,
         \I_cache/cache[5][144] , \I_cache/cache[5][145] ,
         \I_cache/cache[5][146] , \I_cache/cache[5][147] ,
         \I_cache/cache[5][148] , \I_cache/cache[5][149] ,
         \I_cache/cache[5][150] , \I_cache/cache[5][151] ,
         \I_cache/cache[5][152] , \I_cache/cache[5][153] ,
         \I_cache/cache[5][154] , \I_cache/cache[4][0] , \I_cache/cache[4][1] ,
         \I_cache/cache[4][2] , \I_cache/cache[4][3] , \I_cache/cache[4][4] ,
         \I_cache/cache[4][5] , \I_cache/cache[4][6] , \I_cache/cache[4][7] ,
         \I_cache/cache[4][8] , \I_cache/cache[4][9] , \I_cache/cache[4][10] ,
         \I_cache/cache[4][11] , \I_cache/cache[4][12] ,
         \I_cache/cache[4][13] , \I_cache/cache[4][14] ,
         \I_cache/cache[4][15] , \I_cache/cache[4][16] ,
         \I_cache/cache[4][17] , \I_cache/cache[4][18] ,
         \I_cache/cache[4][19] , \I_cache/cache[4][20] ,
         \I_cache/cache[4][21] , \I_cache/cache[4][22] ,
         \I_cache/cache[4][23] , \I_cache/cache[4][24] ,
         \I_cache/cache[4][25] , \I_cache/cache[4][26] ,
         \I_cache/cache[4][27] , \I_cache/cache[4][28] ,
         \I_cache/cache[4][29] , \I_cache/cache[4][30] ,
         \I_cache/cache[4][31] , \I_cache/cache[4][32] ,
         \I_cache/cache[4][33] , \I_cache/cache[4][34] ,
         \I_cache/cache[4][35] , \I_cache/cache[4][36] ,
         \I_cache/cache[4][37] , \I_cache/cache[4][38] ,
         \I_cache/cache[4][39] , \I_cache/cache[4][40] ,
         \I_cache/cache[4][41] , \I_cache/cache[4][42] ,
         \I_cache/cache[4][43] , \I_cache/cache[4][44] ,
         \I_cache/cache[4][45] , \I_cache/cache[4][46] ,
         \I_cache/cache[4][47] , \I_cache/cache[4][48] ,
         \I_cache/cache[4][49] , \I_cache/cache[4][50] ,
         \I_cache/cache[4][51] , \I_cache/cache[4][52] ,
         \I_cache/cache[4][53] , \I_cache/cache[4][54] ,
         \I_cache/cache[4][55] , \I_cache/cache[4][56] ,
         \I_cache/cache[4][57] , \I_cache/cache[4][58] ,
         \I_cache/cache[4][59] , \I_cache/cache[4][60] ,
         \I_cache/cache[4][61] , \I_cache/cache[4][62] ,
         \I_cache/cache[4][63] , \I_cache/cache[4][64] ,
         \I_cache/cache[4][65] , \I_cache/cache[4][66] ,
         \I_cache/cache[4][67] , \I_cache/cache[4][68] ,
         \I_cache/cache[4][69] , \I_cache/cache[4][70] ,
         \I_cache/cache[4][71] , \I_cache/cache[4][72] ,
         \I_cache/cache[4][73] , \I_cache/cache[4][74] ,
         \I_cache/cache[4][75] , \I_cache/cache[4][76] ,
         \I_cache/cache[4][77] , \I_cache/cache[4][78] ,
         \I_cache/cache[4][79] , \I_cache/cache[4][80] ,
         \I_cache/cache[4][81] , \I_cache/cache[4][82] ,
         \I_cache/cache[4][83] , \I_cache/cache[4][84] ,
         \I_cache/cache[4][85] , \I_cache/cache[4][86] ,
         \I_cache/cache[4][87] , \I_cache/cache[4][88] ,
         \I_cache/cache[4][89] , \I_cache/cache[4][90] ,
         \I_cache/cache[4][91] , \I_cache/cache[4][92] ,
         \I_cache/cache[4][93] , \I_cache/cache[4][94] ,
         \I_cache/cache[4][95] , \I_cache/cache[4][96] ,
         \I_cache/cache[4][97] , \I_cache/cache[4][98] ,
         \I_cache/cache[4][99] , \I_cache/cache[4][100] ,
         \I_cache/cache[4][101] , \I_cache/cache[4][102] ,
         \I_cache/cache[4][103] , \I_cache/cache[4][104] ,
         \I_cache/cache[4][105] , \I_cache/cache[4][106] ,
         \I_cache/cache[4][107] , \I_cache/cache[4][108] ,
         \I_cache/cache[4][109] , \I_cache/cache[4][110] ,
         \I_cache/cache[4][111] , \I_cache/cache[4][112] ,
         \I_cache/cache[4][113] , \I_cache/cache[4][114] ,
         \I_cache/cache[4][115] , \I_cache/cache[4][116] ,
         \I_cache/cache[4][117] , \I_cache/cache[4][118] ,
         \I_cache/cache[4][119] , \I_cache/cache[4][120] ,
         \I_cache/cache[4][121] , \I_cache/cache[4][122] ,
         \I_cache/cache[4][123] , \I_cache/cache[4][124] ,
         \I_cache/cache[4][125] , \I_cache/cache[4][126] ,
         \I_cache/cache[4][127] , \I_cache/cache[4][128] ,
         \I_cache/cache[4][129] , \I_cache/cache[4][130] ,
         \I_cache/cache[4][131] , \I_cache/cache[4][132] ,
         \I_cache/cache[4][133] , \I_cache/cache[4][134] ,
         \I_cache/cache[4][135] , \I_cache/cache[4][136] ,
         \I_cache/cache[4][137] , \I_cache/cache[4][138] ,
         \I_cache/cache[4][139] , \I_cache/cache[4][140] ,
         \I_cache/cache[4][141] , \I_cache/cache[4][142] ,
         \I_cache/cache[4][143] , \I_cache/cache[4][144] ,
         \I_cache/cache[4][145] , \I_cache/cache[4][146] ,
         \I_cache/cache[4][147] , \I_cache/cache[4][148] ,
         \I_cache/cache[4][149] , \I_cache/cache[4][150] ,
         \I_cache/cache[4][151] , \I_cache/cache[4][152] ,
         \I_cache/cache[4][153] , \I_cache/cache[4][154] ,
         \I_cache/cache[3][0] , \I_cache/cache[3][1] , \I_cache/cache[3][2] ,
         \I_cache/cache[3][3] , \I_cache/cache[3][4] , \I_cache/cache[3][5] ,
         \I_cache/cache[3][6] , \I_cache/cache[3][7] , \I_cache/cache[3][8] ,
         \I_cache/cache[3][9] , \I_cache/cache[3][10] , \I_cache/cache[3][11] ,
         \I_cache/cache[3][12] , \I_cache/cache[3][13] ,
         \I_cache/cache[3][14] , \I_cache/cache[3][15] ,
         \I_cache/cache[3][16] , \I_cache/cache[3][17] ,
         \I_cache/cache[3][18] , \I_cache/cache[3][19] ,
         \I_cache/cache[3][20] , \I_cache/cache[3][21] ,
         \I_cache/cache[3][22] , \I_cache/cache[3][23] ,
         \I_cache/cache[3][24] , \I_cache/cache[3][25] ,
         \I_cache/cache[3][26] , \I_cache/cache[3][27] ,
         \I_cache/cache[3][28] , \I_cache/cache[3][29] ,
         \I_cache/cache[3][30] , \I_cache/cache[3][31] ,
         \I_cache/cache[3][32] , \I_cache/cache[3][33] ,
         \I_cache/cache[3][34] , \I_cache/cache[3][35] ,
         \I_cache/cache[3][36] , \I_cache/cache[3][37] ,
         \I_cache/cache[3][38] , \I_cache/cache[3][39] ,
         \I_cache/cache[3][40] , \I_cache/cache[3][41] ,
         \I_cache/cache[3][42] , \I_cache/cache[3][43] ,
         \I_cache/cache[3][44] , \I_cache/cache[3][45] ,
         \I_cache/cache[3][46] , \I_cache/cache[3][47] ,
         \I_cache/cache[3][48] , \I_cache/cache[3][49] ,
         \I_cache/cache[3][50] , \I_cache/cache[3][51] ,
         \I_cache/cache[3][52] , \I_cache/cache[3][53] ,
         \I_cache/cache[3][54] , \I_cache/cache[3][55] ,
         \I_cache/cache[3][56] , \I_cache/cache[3][57] ,
         \I_cache/cache[3][58] , \I_cache/cache[3][59] ,
         \I_cache/cache[3][60] , \I_cache/cache[3][61] ,
         \I_cache/cache[3][62] , \I_cache/cache[3][63] ,
         \I_cache/cache[3][64] , \I_cache/cache[3][65] ,
         \I_cache/cache[3][66] , \I_cache/cache[3][67] ,
         \I_cache/cache[3][68] , \I_cache/cache[3][69] ,
         \I_cache/cache[3][70] , \I_cache/cache[3][71] ,
         \I_cache/cache[3][72] , \I_cache/cache[3][73] ,
         \I_cache/cache[3][74] , \I_cache/cache[3][75] ,
         \I_cache/cache[3][76] , \I_cache/cache[3][77] ,
         \I_cache/cache[3][78] , \I_cache/cache[3][79] ,
         \I_cache/cache[3][80] , \I_cache/cache[3][81] ,
         \I_cache/cache[3][82] , \I_cache/cache[3][83] ,
         \I_cache/cache[3][84] , \I_cache/cache[3][85] ,
         \I_cache/cache[3][86] , \I_cache/cache[3][87] ,
         \I_cache/cache[3][88] , \I_cache/cache[3][89] ,
         \I_cache/cache[3][90] , \I_cache/cache[3][91] ,
         \I_cache/cache[3][92] , \I_cache/cache[3][93] ,
         \I_cache/cache[3][94] , \I_cache/cache[3][95] ,
         \I_cache/cache[3][96] , \I_cache/cache[3][97] ,
         \I_cache/cache[3][98] , \I_cache/cache[3][99] ,
         \I_cache/cache[3][100] , \I_cache/cache[3][101] ,
         \I_cache/cache[3][102] , \I_cache/cache[3][103] ,
         \I_cache/cache[3][104] , \I_cache/cache[3][105] ,
         \I_cache/cache[3][106] , \I_cache/cache[3][107] ,
         \I_cache/cache[3][108] , \I_cache/cache[3][109] ,
         \I_cache/cache[3][110] , \I_cache/cache[3][111] ,
         \I_cache/cache[3][112] , \I_cache/cache[3][113] ,
         \I_cache/cache[3][114] , \I_cache/cache[3][115] ,
         \I_cache/cache[3][116] , \I_cache/cache[3][117] ,
         \I_cache/cache[3][118] , \I_cache/cache[3][119] ,
         \I_cache/cache[3][120] , \I_cache/cache[3][121] ,
         \I_cache/cache[3][122] , \I_cache/cache[3][123] ,
         \I_cache/cache[3][124] , \I_cache/cache[3][125] ,
         \I_cache/cache[3][126] , \I_cache/cache[3][127] ,
         \I_cache/cache[3][128] , \I_cache/cache[3][129] ,
         \I_cache/cache[3][130] , \I_cache/cache[3][131] ,
         \I_cache/cache[3][132] , \I_cache/cache[3][133] ,
         \I_cache/cache[3][134] , \I_cache/cache[3][135] ,
         \I_cache/cache[3][136] , \I_cache/cache[3][137] ,
         \I_cache/cache[3][138] , \I_cache/cache[3][139] ,
         \I_cache/cache[3][140] , \I_cache/cache[3][141] ,
         \I_cache/cache[3][142] , \I_cache/cache[3][143] ,
         \I_cache/cache[3][144] , \I_cache/cache[3][145] ,
         \I_cache/cache[3][146] , \I_cache/cache[3][147] ,
         \I_cache/cache[3][148] , \I_cache/cache[3][149] ,
         \I_cache/cache[3][150] , \I_cache/cache[3][151] ,
         \I_cache/cache[3][152] , \I_cache/cache[3][153] ,
         \I_cache/cache[3][154] , \I_cache/cache[2][0] , \I_cache/cache[2][1] ,
         \I_cache/cache[2][2] , \I_cache/cache[2][3] , \I_cache/cache[2][4] ,
         \I_cache/cache[2][5] , \I_cache/cache[2][6] , \I_cache/cache[2][7] ,
         \I_cache/cache[2][8] , \I_cache/cache[2][9] , \I_cache/cache[2][10] ,
         \I_cache/cache[2][11] , \I_cache/cache[2][12] ,
         \I_cache/cache[2][13] , \I_cache/cache[2][14] ,
         \I_cache/cache[2][15] , \I_cache/cache[2][16] ,
         \I_cache/cache[2][17] , \I_cache/cache[2][18] ,
         \I_cache/cache[2][19] , \I_cache/cache[2][20] ,
         \I_cache/cache[2][21] , \I_cache/cache[2][22] ,
         \I_cache/cache[2][23] , \I_cache/cache[2][24] ,
         \I_cache/cache[2][25] , \I_cache/cache[2][26] ,
         \I_cache/cache[2][27] , \I_cache/cache[2][28] ,
         \I_cache/cache[2][29] , \I_cache/cache[2][30] ,
         \I_cache/cache[2][31] , \I_cache/cache[2][32] ,
         \I_cache/cache[2][33] , \I_cache/cache[2][34] ,
         \I_cache/cache[2][35] , \I_cache/cache[2][36] ,
         \I_cache/cache[2][37] , \I_cache/cache[2][38] ,
         \I_cache/cache[2][39] , \I_cache/cache[2][40] ,
         \I_cache/cache[2][41] , \I_cache/cache[2][42] ,
         \I_cache/cache[2][43] , \I_cache/cache[2][44] ,
         \I_cache/cache[2][45] , \I_cache/cache[2][46] ,
         \I_cache/cache[2][47] , \I_cache/cache[2][48] ,
         \I_cache/cache[2][49] , \I_cache/cache[2][50] ,
         \I_cache/cache[2][51] , \I_cache/cache[2][52] ,
         \I_cache/cache[2][53] , \I_cache/cache[2][54] ,
         \I_cache/cache[2][55] , \I_cache/cache[2][56] ,
         \I_cache/cache[2][57] , \I_cache/cache[2][58] ,
         \I_cache/cache[2][59] , \I_cache/cache[2][60] ,
         \I_cache/cache[2][61] , \I_cache/cache[2][62] ,
         \I_cache/cache[2][63] , \I_cache/cache[2][64] ,
         \I_cache/cache[2][65] , \I_cache/cache[2][66] ,
         \I_cache/cache[2][67] , \I_cache/cache[2][68] ,
         \I_cache/cache[2][69] , \I_cache/cache[2][70] ,
         \I_cache/cache[2][71] , \I_cache/cache[2][72] ,
         \I_cache/cache[2][73] , \I_cache/cache[2][74] ,
         \I_cache/cache[2][75] , \I_cache/cache[2][76] ,
         \I_cache/cache[2][77] , \I_cache/cache[2][78] ,
         \I_cache/cache[2][79] , \I_cache/cache[2][80] ,
         \I_cache/cache[2][81] , \I_cache/cache[2][82] ,
         \I_cache/cache[2][83] , \I_cache/cache[2][84] ,
         \I_cache/cache[2][85] , \I_cache/cache[2][86] ,
         \I_cache/cache[2][87] , \I_cache/cache[2][88] ,
         \I_cache/cache[2][89] , \I_cache/cache[2][90] ,
         \I_cache/cache[2][91] , \I_cache/cache[2][92] ,
         \I_cache/cache[2][93] , \I_cache/cache[2][94] ,
         \I_cache/cache[2][95] , \I_cache/cache[2][96] ,
         \I_cache/cache[2][97] , \I_cache/cache[2][98] ,
         \I_cache/cache[2][99] , \I_cache/cache[2][100] ,
         \I_cache/cache[2][101] , \I_cache/cache[2][102] ,
         \I_cache/cache[2][103] , \I_cache/cache[2][104] ,
         \I_cache/cache[2][105] , \I_cache/cache[2][106] ,
         \I_cache/cache[2][107] , \I_cache/cache[2][108] ,
         \I_cache/cache[2][109] , \I_cache/cache[2][110] ,
         \I_cache/cache[2][111] , \I_cache/cache[2][112] ,
         \I_cache/cache[2][113] , \I_cache/cache[2][114] ,
         \I_cache/cache[2][115] , \I_cache/cache[2][116] ,
         \I_cache/cache[2][117] , \I_cache/cache[2][118] ,
         \I_cache/cache[2][119] , \I_cache/cache[2][120] ,
         \I_cache/cache[2][121] , \I_cache/cache[2][122] ,
         \I_cache/cache[2][123] , \I_cache/cache[2][124] ,
         \I_cache/cache[2][125] , \I_cache/cache[2][126] ,
         \I_cache/cache[2][127] , \I_cache/cache[2][128] ,
         \I_cache/cache[2][129] , \I_cache/cache[2][130] ,
         \I_cache/cache[2][131] , \I_cache/cache[2][132] ,
         \I_cache/cache[2][133] , \I_cache/cache[2][134] ,
         \I_cache/cache[2][135] , \I_cache/cache[2][136] ,
         \I_cache/cache[2][137] , \I_cache/cache[2][138] ,
         \I_cache/cache[2][139] , \I_cache/cache[2][140] ,
         \I_cache/cache[2][141] , \I_cache/cache[2][142] ,
         \I_cache/cache[2][143] , \I_cache/cache[2][144] ,
         \I_cache/cache[2][145] , \I_cache/cache[2][146] ,
         \I_cache/cache[2][147] , \I_cache/cache[2][148] ,
         \I_cache/cache[2][149] , \I_cache/cache[2][150] ,
         \I_cache/cache[2][151] , \I_cache/cache[2][152] ,
         \I_cache/cache[2][153] , \I_cache/cache[2][154] ,
         \I_cache/cache[1][0] , \I_cache/cache[1][1] , \I_cache/cache[1][2] ,
         \I_cache/cache[1][3] , \I_cache/cache[1][4] , \I_cache/cache[1][5] ,
         \I_cache/cache[1][6] , \I_cache/cache[1][7] , \I_cache/cache[1][8] ,
         \I_cache/cache[1][9] , \I_cache/cache[1][10] , \I_cache/cache[1][11] ,
         \I_cache/cache[1][12] , \I_cache/cache[1][13] ,
         \I_cache/cache[1][14] , \I_cache/cache[1][15] ,
         \I_cache/cache[1][16] , \I_cache/cache[1][17] ,
         \I_cache/cache[1][18] , \I_cache/cache[1][19] ,
         \I_cache/cache[1][20] , \I_cache/cache[1][21] ,
         \I_cache/cache[1][22] , \I_cache/cache[1][23] ,
         \I_cache/cache[1][24] , \I_cache/cache[1][25] ,
         \I_cache/cache[1][26] , \I_cache/cache[1][27] ,
         \I_cache/cache[1][28] , \I_cache/cache[1][29] ,
         \I_cache/cache[1][30] , \I_cache/cache[1][31] ,
         \I_cache/cache[1][32] , \I_cache/cache[1][33] ,
         \I_cache/cache[1][34] , \I_cache/cache[1][35] ,
         \I_cache/cache[1][36] , \I_cache/cache[1][37] ,
         \I_cache/cache[1][38] , \I_cache/cache[1][39] ,
         \I_cache/cache[1][40] , \I_cache/cache[1][41] ,
         \I_cache/cache[1][42] , \I_cache/cache[1][43] ,
         \I_cache/cache[1][44] , \I_cache/cache[1][45] ,
         \I_cache/cache[1][46] , \I_cache/cache[1][47] ,
         \I_cache/cache[1][48] , \I_cache/cache[1][49] ,
         \I_cache/cache[1][50] , \I_cache/cache[1][51] ,
         \I_cache/cache[1][52] , \I_cache/cache[1][53] ,
         \I_cache/cache[1][54] , \I_cache/cache[1][55] ,
         \I_cache/cache[1][56] , \I_cache/cache[1][57] ,
         \I_cache/cache[1][58] , \I_cache/cache[1][59] ,
         \I_cache/cache[1][60] , \I_cache/cache[1][61] ,
         \I_cache/cache[1][62] , \I_cache/cache[1][63] ,
         \I_cache/cache[1][64] , \I_cache/cache[1][65] ,
         \I_cache/cache[1][66] , \I_cache/cache[1][67] ,
         \I_cache/cache[1][68] , \I_cache/cache[1][69] ,
         \I_cache/cache[1][70] , \I_cache/cache[1][71] ,
         \I_cache/cache[1][72] , \I_cache/cache[1][73] ,
         \I_cache/cache[1][74] , \I_cache/cache[1][75] ,
         \I_cache/cache[1][76] , \I_cache/cache[1][77] ,
         \I_cache/cache[1][78] , \I_cache/cache[1][79] ,
         \I_cache/cache[1][80] , \I_cache/cache[1][81] ,
         \I_cache/cache[1][82] , \I_cache/cache[1][83] ,
         \I_cache/cache[1][84] , \I_cache/cache[1][85] ,
         \I_cache/cache[1][86] , \I_cache/cache[1][87] ,
         \I_cache/cache[1][88] , \I_cache/cache[1][89] ,
         \I_cache/cache[1][90] , \I_cache/cache[1][91] ,
         \I_cache/cache[1][92] , \I_cache/cache[1][93] ,
         \I_cache/cache[1][94] , \I_cache/cache[1][95] ,
         \I_cache/cache[1][96] , \I_cache/cache[1][97] ,
         \I_cache/cache[1][98] , \I_cache/cache[1][99] ,
         \I_cache/cache[1][100] , \I_cache/cache[1][101] ,
         \I_cache/cache[1][102] , \I_cache/cache[1][103] ,
         \I_cache/cache[1][104] , \I_cache/cache[1][105] ,
         \I_cache/cache[1][106] , \I_cache/cache[1][107] ,
         \I_cache/cache[1][108] , \I_cache/cache[1][109] ,
         \I_cache/cache[1][110] , \I_cache/cache[1][111] ,
         \I_cache/cache[1][112] , \I_cache/cache[1][113] ,
         \I_cache/cache[1][114] , \I_cache/cache[1][115] ,
         \I_cache/cache[1][116] , \I_cache/cache[1][117] ,
         \I_cache/cache[1][118] , \I_cache/cache[1][119] ,
         \I_cache/cache[1][120] , \I_cache/cache[1][121] ,
         \I_cache/cache[1][122] , \I_cache/cache[1][123] ,
         \I_cache/cache[1][124] , \I_cache/cache[1][125] ,
         \I_cache/cache[1][126] , \I_cache/cache[1][127] ,
         \I_cache/cache[1][128] , \I_cache/cache[1][129] ,
         \I_cache/cache[1][130] , \I_cache/cache[1][131] ,
         \I_cache/cache[1][132] , \I_cache/cache[1][133] ,
         \I_cache/cache[1][134] , \I_cache/cache[1][135] ,
         \I_cache/cache[1][136] , \I_cache/cache[1][137] ,
         \I_cache/cache[1][138] , \I_cache/cache[1][139] ,
         \I_cache/cache[1][140] , \I_cache/cache[1][141] ,
         \I_cache/cache[1][142] , \I_cache/cache[1][143] ,
         \I_cache/cache[1][144] , \I_cache/cache[1][145] ,
         \I_cache/cache[1][146] , \I_cache/cache[1][147] ,
         \I_cache/cache[1][148] , \I_cache/cache[1][149] ,
         \I_cache/cache[1][150] , \I_cache/cache[1][151] ,
         \I_cache/cache[1][152] , \I_cache/cache[1][153] ,
         \I_cache/cache[1][154] , \I_cache/cache[0][0] , \I_cache/cache[0][1] ,
         \I_cache/cache[0][2] , \I_cache/cache[0][3] , \I_cache/cache[0][4] ,
         \I_cache/cache[0][5] , \I_cache/cache[0][6] , \I_cache/cache[0][7] ,
         \I_cache/cache[0][8] , \I_cache/cache[0][9] , \I_cache/cache[0][10] ,
         \I_cache/cache[0][11] , \I_cache/cache[0][12] ,
         \I_cache/cache[0][13] , \I_cache/cache[0][14] ,
         \I_cache/cache[0][15] , \I_cache/cache[0][16] ,
         \I_cache/cache[0][17] , \I_cache/cache[0][18] ,
         \I_cache/cache[0][19] , \I_cache/cache[0][20] ,
         \I_cache/cache[0][21] , \I_cache/cache[0][22] ,
         \I_cache/cache[0][23] , \I_cache/cache[0][24] ,
         \I_cache/cache[0][25] , \I_cache/cache[0][26] ,
         \I_cache/cache[0][27] , \I_cache/cache[0][28] ,
         \I_cache/cache[0][29] , \I_cache/cache[0][30] ,
         \I_cache/cache[0][31] , \I_cache/cache[0][32] ,
         \I_cache/cache[0][33] , \I_cache/cache[0][34] ,
         \I_cache/cache[0][35] , \I_cache/cache[0][36] ,
         \I_cache/cache[0][37] , \I_cache/cache[0][38] ,
         \I_cache/cache[0][39] , \I_cache/cache[0][40] ,
         \I_cache/cache[0][41] , \I_cache/cache[0][42] ,
         \I_cache/cache[0][43] , \I_cache/cache[0][44] ,
         \I_cache/cache[0][45] , \I_cache/cache[0][46] ,
         \I_cache/cache[0][47] , \I_cache/cache[0][48] ,
         \I_cache/cache[0][49] , \I_cache/cache[0][50] ,
         \I_cache/cache[0][51] , \I_cache/cache[0][52] ,
         \I_cache/cache[0][53] , \I_cache/cache[0][54] ,
         \I_cache/cache[0][55] , \I_cache/cache[0][56] ,
         \I_cache/cache[0][57] , \I_cache/cache[0][58] ,
         \I_cache/cache[0][59] , \I_cache/cache[0][60] ,
         \I_cache/cache[0][61] , \I_cache/cache[0][62] ,
         \I_cache/cache[0][63] , \I_cache/cache[0][64] ,
         \I_cache/cache[0][65] , \I_cache/cache[0][66] ,
         \I_cache/cache[0][67] , \I_cache/cache[0][68] ,
         \I_cache/cache[0][69] , \I_cache/cache[0][70] ,
         \I_cache/cache[0][71] , \I_cache/cache[0][72] ,
         \I_cache/cache[0][73] , \I_cache/cache[0][74] ,
         \I_cache/cache[0][75] , \I_cache/cache[0][76] ,
         \I_cache/cache[0][77] , \I_cache/cache[0][78] ,
         \I_cache/cache[0][79] , \I_cache/cache[0][80] ,
         \I_cache/cache[0][81] , \I_cache/cache[0][82] ,
         \I_cache/cache[0][83] , \I_cache/cache[0][84] ,
         \I_cache/cache[0][85] , \I_cache/cache[0][86] ,
         \I_cache/cache[0][87] , \I_cache/cache[0][88] ,
         \I_cache/cache[0][89] , \I_cache/cache[0][90] ,
         \I_cache/cache[0][91] , \I_cache/cache[0][92] ,
         \I_cache/cache[0][93] , \I_cache/cache[0][94] ,
         \I_cache/cache[0][95] , \I_cache/cache[0][96] ,
         \I_cache/cache[0][97] , \I_cache/cache[0][98] ,
         \I_cache/cache[0][99] , \I_cache/cache[0][100] ,
         \I_cache/cache[0][101] , \I_cache/cache[0][102] ,
         \I_cache/cache[0][103] , \I_cache/cache[0][104] ,
         \I_cache/cache[0][105] , \I_cache/cache[0][106] ,
         \I_cache/cache[0][107] , \I_cache/cache[0][108] ,
         \I_cache/cache[0][109] , \I_cache/cache[0][110] ,
         \I_cache/cache[0][111] , \I_cache/cache[0][112] ,
         \I_cache/cache[0][113] , \I_cache/cache[0][114] ,
         \I_cache/cache[0][115] , \I_cache/cache[0][116] ,
         \I_cache/cache[0][117] , \I_cache/cache[0][118] ,
         \I_cache/cache[0][119] , \I_cache/cache[0][120] ,
         \I_cache/cache[0][121] , \I_cache/cache[0][122] ,
         \I_cache/cache[0][123] , \I_cache/cache[0][124] ,
         \I_cache/cache[0][125] , \I_cache/cache[0][126] ,
         \I_cache/cache[0][127] , \I_cache/cache[0][128] ,
         \I_cache/cache[0][129] , \I_cache/cache[0][130] ,
         \I_cache/cache[0][131] , \I_cache/cache[0][132] ,
         \I_cache/cache[0][133] , \I_cache/cache[0][134] ,
         \I_cache/cache[0][135] , \I_cache/cache[0][136] ,
         \I_cache/cache[0][137] , \I_cache/cache[0][138] ,
         \I_cache/cache[0][139] , \I_cache/cache[0][140] ,
         \I_cache/cache[0][141] , \I_cache/cache[0][142] ,
         \I_cache/cache[0][143] , \I_cache/cache[0][144] ,
         \I_cache/cache[0][145] , \I_cache/cache[0][146] ,
         \I_cache/cache[0][147] , \I_cache/cache[0][148] ,
         \I_cache/cache[0][149] , \I_cache/cache[0][150] ,
         \I_cache/cache[0][151] , \I_cache/cache[0][152] ,
         \I_cache/cache[0][153] , \I_cache/cache[0][154] , net98089, net98121,
         net98153, net98375, net98391, net98396, net98429, net98430, net98432,
         net98436, net98447, net98449, net98472, net98501, net98564, net98880,
         net98881, net98897, net98898, net98899, net98900, net98901, net98915,
         net98929, net98932, net98946, net98950, net98951, net98952, net98964,
         net98965, net98966, net98967, net98968, net98970, net98971, net98973,
         net98974, net98988, net98992, net98993, net98994, net99009, net99014,
         net99015, net99016, net99019, net99037, net99038, net99039, net99042,
         net99056, net99060, net99061, net99062, net99064, net99078, net99080,
         net99087, net99089, net99090, net99104, net99108, net99109, net99110,
         net99146, net99254, net99267, net99270, net99284, net99288, net99289,
         net99290, net99293, net99307, net99311, net99312, net99313, net99316,
         net99330, net99334, net99335, net99336, net99354, net99359, net99360,
         net99363, net99364, net99378, net99382, net99383, net99384, net99386,
         net99387, net99401, net99405, net99406, net99407, net99410, net99424,
         net99428, net99429, net99430, net99432, net99447, net99450, net99461,
         net99464, net99475, net99476, net99477, net99502, net99503, net99504,
         net99531, net99536, net99537, net99538, net99541, net99555, net99576,
         net99581, net99582, net99583, net99603, net99604, net99605, net99607,
         net99609, net99624, net99634, net99637, net99638, net99639, net99654,
         net99664, net99671, net99693, net99711, net99712, net99734, net99737,
         net99753, net99759, net99760, net99765, net99814, net99815, net99845,
         net99849, net99855, net99932, net99933, net99935, net99936, net99962,
         net99969, net99970, net99971, net99974, net99977, net99978, net99991,
         net100015, net100023, net100025, net100026, net100029, net100032,
         net100035, net100038, net100039, net100042, net100044, net100048,
         net100049, net100079, net100081, net100082, net100084, net100087,
         net100093, net100095, net100096, net100099, net100103, net100104,
         net100748, net100749, net100750, net100751, net100866, net101969,
         net101970, net101971, net101973, net101981, net101983, net102036,
         net102087, net102088, net102094, net102095, net102120, net102121,
         net102183, net102300, net102344, net102345, net102346, net102371,
         net102372, net102413, net102500, net102565, net102651, net102744,
         net102745, net102746, net102899, net102900, net102901, net103059,
         net103060, net103061, net103218, net103220, net103390, net103391,
         net103392, net103393, net103394, net103479, net103630, net103707,
         net103708, net103709, net103795, net103869, net103871, net104023,
         net104024, net104025, net104183, net104184, net104185, net104271,
         net104351, net104352, net104353, net104440, net104524, net104525,
         net104526, net104563, net104564, net104704, net104705, net104706,
         net104829, net104831, net104868, net104869, net105003, net105004,
         net105008, net105009, net105010, net105011, net105020, net105021,
         net105022, net105023, net105044, net105045, net105046, net105047,
         net105120, net105150, net105151, net105152, net105284, net105285,
         net105286, net105373, net105425, net105426, net105427, net105577,
         net105578, net105579, net105666, net105735, net105736, net105737,
         net105824, net105929, net105930, net105931, net106078, net106108,
         net106109, net106110, net106270, net106271, net106272, net106418,
         net106419, net106420, net106535, net106564, net106565, net106566,
         net106801, net106881, net106977, net107011, net107041, net107042,
         net107043, net107168, net107236, net107237, net107238, net108204,
         net108963, net108959, net109183, net109181, net109179, net109185,
         net109795, net109791, net109805, net109801, net110191, net110189,
         net110205, net110227, net110225, net110221, net110219, net110217,
         net110215, net110213, net110239, net110233, net110231, net110229,
         net110243, net110241, net110259, net110257, net110255, net110253,
         net110251, net110249, net110247, net111405, net111409, net111845,
         net111837, net111835, net111983, net111979, net111977, net111969,
         net111967, net111965, net111963, net111961, net111959, net111957,
         net111955, net111953, net111951, net111949, net111947, net111945,
         net111943, net111941, net111939, net111937, net111935, net111933,
         net111931, net111929, net111927, net111925, net111923, net111921,
         net111919, net111917, net111915, net111905, net111889, net111885,
         net111883, net111881, net111879, net111877, net111873, net111871,
         net111867, net111865, net112107, net112105, net112101, net112097,
         net112095, net112093, net112091, net112089, net112087, net112085,
         net112083, net112081, net112079, net112077, net112075, net112073,
         net112071, net112069, net112067, net112065, net112063, net112061,
         net112059, net112057, net112055, net112053, net112051, net112049,
         net112047, net112045, net112043, net112041, net112037, net112033,
         net112019, net112011, net112009, net112005, net112003, net111999,
         net111995, net111993, net111991, net111989, net112187, net112169,
         net112165, net112163, net112161, net112159, net112155, net112153,
         net112151, net112147, net112145, net112143, net112139, net112137,
         net112131, net112129, net112127, net112125, net112123, net112121,
         net112119, net112117, net112115, net112113, net112271, net112269,
         net112265, net112263, net112259, net112257, net112245, net112241,
         net112239, net112237, net112235, net112233, net112231, net112229,
         net112221, net112217, net112215, net112213, net112211, net112201,
         net112199, net112197, net112195, net112385, net112383, net112381,
         net112379, net112377, net112369, net112367, net112363, net112361,
         net112359, net112357, net112355, net112353, net112351, net112349,
         net112347, net112345, net112343, net112341, net112339, net112337,
         net112335, net112333, net112331, net112329, net112325, net112319,
         net112303, net112301, net112295, net112293, net112291, net112289,
         net112285, net112283, net112281, net112279, net112277, net112519,
         net112517, net112515, net112511, net112509, net112507, net112505,
         net112503, net112499, net112497, net112493, net112491, net112489,
         net112487, net112485, net112483, net112481, net112477, net112473,
         net112471, net112469, net112467, net112465, net112463, net112461,
         net112459, net112457, net112455, net112453, net112449, net112443,
         net112431, net112429, net112427, net112425, net112423, net112419,
         net112417, net112415, net112411, net112409, net112405, net112403,
         net112401, net112601, net112599, net112593, net112589, net112587,
         net112585, net112583, net112577, net112575, net112573, net112571,
         net112569, net112565, net112563, net112561, net112555, net112547,
         net112545, net112543, net112541, net112539, net112537, net112535,
         net112533, net112531, net112529, net112527, net112525, net112609,
         net112607, net112701, net112697, net112695, net112693, net112691,
         net112687, net112681, net112679, net112673, net112671, net112667,
         net112665, net112663, net112659, net112657, net112655, net112651,
         net112649, net112647, net112645, net112643, net112641, net112639,
         net112637, net112635, net112633, net112631, net112629, net112627,
         net112713, net112709, net112707, net112723, net112721, net112725,
         net112731, net112729, net112727, net113041, net113039, net113047,
         net113083, net113081, net113079, net113077, net113075, net113089,
         net113087, net113169, net113167, net113439, net113437, net113447,
         net113445, net113457, net113455, net113463, net113461, net113533,
         net113532, net113537, net113541, net113540, net113551, net113592,
         net113608, net113607, net113606, net113605, net113667, net113725,
         net113916, net113919, net113983, net114031, net114085, net114092,
         net114113, net126164, net130301, net130420, net130474, net130509,
         net130576, net130594, net131142, net134088, net134093, net134103,
         net134107, net134109, net134117, net134118, net134133, net137471,
         net137470, net138398, net139669, net139682, net139681, net139803,
         net140281, net140280, net140278, net140424, net140423, net140445,
         net140444, net140551, net99850, net102400, net102398, net102397,
         net105006, net105005, net100020, net100019, net100013, net98185,
         net105035, net105034, net105033, net105032, net112705, net112703,
         net100105, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3518, n3520, n3521, n3522, n3523, n3524,
         n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533, n3534,
         n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543, n3544,
         n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553, n3554,
         n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563, n3564,
         n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3685,
         n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694, n3695,
         n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704, n3705,
         n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714, n3715,
         n3716, n3718, n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726,
         n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736,
         n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746,
         n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756,
         n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
         n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776,
         n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786,
         n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796,
         n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806,
         n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816,
         n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826,
         n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836,
         n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846,
         n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856,
         n3857, n3858, n3859, n3860, n3861, n3862, n3864, n3865, n3866, n3867,
         n3868, n3869, n3870, n3871, n3872, n3881, n3883, n3884, n3885, n3889,
         n3890, n3891, n3892, n3893, n3961, n3964, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4028, n4029,
         n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039,
         n4040, n4041, n4042, n4043, n4044, n4045, n4047, n4048, n4049, n4050,
         n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4060, n4061,
         n4062, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
         n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329,
         n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339,
         n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349,
         n4350, n4351, n4385, n4393, n4395, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4719,
         n4722, n4723, n4724, n4727, n4728, n4743, n4746, n4747, n4748, n4750,
         n4751, n4752, n4754, n4756, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4780, n4782, n4783, n4784, n4787,
         n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797,
         n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807,
         n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
         n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
         n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
         n4838, n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847,
         n4848, n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857,
         n4858, n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867,
         n4868, n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877,
         n4878, n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887,
         n4888, n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897,
         n4898, n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907,
         n4908, n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917,
         n4918, n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927,
         n4928, n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937,
         n4938, n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947,
         n4948, n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957,
         n4958, n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967,
         n4968, n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977,
         n4978, n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987,
         n4988, n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997,
         n4998, n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007,
         n5008, n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017,
         n5018, n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027,
         n5028, n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037,
         n5038, n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047,
         n5048, n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057,
         n5058, n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067,
         n5068, n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077,
         n5078, n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087,
         n5088, n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097,
         n5098, n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107,
         n5108, n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117,
         n5118, n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127,
         n5128, n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137,
         n5138, n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147,
         n5148, n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157,
         n5158, n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167,
         n5168, n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177,
         n5178, n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187,
         n5188, n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197,
         n5198, n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207,
         n5208, n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217,
         n5218, n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227,
         n5228, n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237,
         n5238, n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247,
         n5248, n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257,
         n5258, n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267,
         n5268, n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277,
         n5278, n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287,
         n5288, n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297,
         n5298, n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307,
         n5308, n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317,
         n5318, n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327,
         n5328, n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337,
         n5338, n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347,
         n5348, n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357,
         n5358, n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367,
         n5368, n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377,
         n5378, n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387,
         n5388, n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397,
         n5398, n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407,
         n5408, n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417,
         n5418, n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427,
         n5428, n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437,
         n5438, n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447,
         n5448, n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457,
         n5458, n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467,
         n5468, n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477,
         n5478, n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487,
         n5488, n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497,
         n5498, n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507,
         n5508, n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517,
         n5518, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530,
         n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
         n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
         n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
         n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
         n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
         n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
         n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
         n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
         n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
         n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
         n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
         n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
         n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
         n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
         n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
         n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
         n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
         n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
         n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
         n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
         n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
         n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
         n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
         n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
         n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
         n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
         n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
         n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
         n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850,
         n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
         n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
         n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
         n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950,
         n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960,
         n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970,
         n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980,
         n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990,
         n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000,
         n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010,
         n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020,
         n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030,
         n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040,
         n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050,
         n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060,
         n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070,
         n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080,
         n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090,
         n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100,
         n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110,
         n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120,
         n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130,
         n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140,
         n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150,
         n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160,
         n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170,
         n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180,
         n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190,
         n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200,
         n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210,
         n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220,
         n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230,
         n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240,
         n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250,
         n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260,
         n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270,
         n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280,
         n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290,
         n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300,
         n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310,
         n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320,
         n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330,
         n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340,
         n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350,
         n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360,
         n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370,
         n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380,
         n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390,
         n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400,
         n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410,
         n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420,
         n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430,
         n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440,
         n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450,
         n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460,
         n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470,
         n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480,
         n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490,
         n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500,
         n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510,
         n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520,
         n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530,
         n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540,
         n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550,
         n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560,
         n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570,
         n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580,
         n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590,
         n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600,
         n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610,
         n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620,
         n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630,
         n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640,
         n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650,
         n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660,
         n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670,
         n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680,
         n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690,
         n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700,
         n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710,
         n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720,
         n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730,
         n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740,
         n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750,
         n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760,
         n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770,
         n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780,
         n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790,
         n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800,
         n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810,
         n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820,
         n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830,
         n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840,
         n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850,
         n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860,
         n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870,
         n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880,
         n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890,
         n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900,
         n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910,
         n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920,
         n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930,
         n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940,
         n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950,
         n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960,
         n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970,
         n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980,
         n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990,
         n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000,
         n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010,
         n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020,
         n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030,
         n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040,
         n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050,
         n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060,
         n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070,
         n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080,
         n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090,
         n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100,
         n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110,
         n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120,
         n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130,
         n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140,
         n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150,
         n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160,
         n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170,
         n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180,
         n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190,
         n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200,
         n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210,
         n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220,
         n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230,
         n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240,
         n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250,
         n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260,
         n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270,
         n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280,
         n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290,
         n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300,
         n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310,
         n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320,
         n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330,
         n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340,
         n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350,
         n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360,
         n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370,
         n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380,
         n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390,
         n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400,
         n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410,
         n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420,
         n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430,
         n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440,
         n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450,
         n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460,
         n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470,
         n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480,
         n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490,
         n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500,
         n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510,
         n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520,
         n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530,
         n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540,
         n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550,
         n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560,
         n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570,
         n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580,
         n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590,
         n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600,
         n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610,
         n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620,
         n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630,
         n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640,
         n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650,
         n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660,
         n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670,
         n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680,
         n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690,
         n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700,
         n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710,
         n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720,
         n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730,
         n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740,
         n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750,
         n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760,
         n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770,
         n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780,
         n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790,
         n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800,
         n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810,
         n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820,
         n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830,
         n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840,
         n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850,
         n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860,
         n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870,
         n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880,
         n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890,
         n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900,
         n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910,
         n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920,
         n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930,
         n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940,
         n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950,
         n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960,
         n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970,
         n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980,
         n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990,
         n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000,
         n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010,
         n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020,
         n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030,
         n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040,
         n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050,
         n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060,
         n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070,
         n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080,
         n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090,
         n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100,
         n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110,
         n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120,
         n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130,
         n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140,
         n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150,
         n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160,
         n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170,
         n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180,
         n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190,
         n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200,
         n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210,
         n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220,
         n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230,
         n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240,
         n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250,
         n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260,
         n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270,
         n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280,
         n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290,
         n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300,
         n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310,
         n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320,
         n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330,
         n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340,
         n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350,
         n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360,
         n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370,
         n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380,
         n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390,
         n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400,
         n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410,
         n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420,
         n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430,
         n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440,
         n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450,
         n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460,
         n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470,
         n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480,
         n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490,
         n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500,
         n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510,
         n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520,
         n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530,
         n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540,
         n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550,
         n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560,
         n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570,
         n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580,
         n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588, n8589, n8590,
         n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598, n8599, n8600,
         n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608, n8609, n8610,
         n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618, n8619, n8620,
         n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628, n8629, n8630,
         n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638, n8639, n8640,
         n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648, n8649, n8650,
         n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658, n8659, n8660,
         n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668, n8669, n8670,
         n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678, n8679, n8680,
         n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688, n8689, n8690,
         n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698, n8699, n8700,
         n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708, n8709, n8710,
         n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718, n8719, n8720,
         n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728, n8729, n8730,
         n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738, n8739, n8740,
         n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748, n8749, n8750,
         n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758, n8759, n8760,
         n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768, n8769, n8770,
         n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778, n8779, n8780,
         n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788, n8789, n8790,
         n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798, n8799, n8800,
         n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808, n8809, n8810,
         n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818, n8819, n8820,
         n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828, n8829, n8830,
         n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838, n8839, n8840,
         n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848, n8849, n8850,
         n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858, n8859, n8860,
         n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868, n8869, n8870,
         n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878, n8879, n8880,
         n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888, n8889, n8890,
         n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898, n8899, n8900,
         n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908, n8909, n8910,
         n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918, n8919, n8920,
         n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928, n8929, n8930,
         n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938, n8939, n8940,
         n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948, n8949, n8950,
         n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958, n8959, n8960,
         n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968, n8969, n8970,
         n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978, n8979, n8980,
         n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988, n8989, n8990,
         n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998, n8999, n9000,
         n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008, n9009, n9010,
         n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018, n9019, n9020,
         n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028, n9029, n9030,
         n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038, n9039, n9040,
         n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048, n9049, n9050,
         n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058, n9059, n9060,
         n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068, n9069, n9070,
         n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078, n9079, n9080,
         n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088, n9089, n9090,
         n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098, n9099, n9100,
         n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108, n9109, n9110,
         n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118, n9119, n9120,
         n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128, n9129, n9130,
         n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138, n9139, n9140,
         n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148, n9149, n9150,
         n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158, n9159, n9160,
         n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168, n9169, n9170,
         n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178, n9179, n9180,
         n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188, n9189, n9190,
         n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198, n9199, n9200,
         n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208, n9209, n9210,
         n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218, n9219, n9220,
         n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228, n9229, n9230,
         n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238, n9239, n9240,
         n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248, n9249, n9250,
         n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258, n9259, n9260,
         n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268, n9269, n9270,
         n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278, n9279, n9280,
         n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288, n9289, n9290,
         n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298, n9299, n9300,
         n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308, n9309, n9310,
         n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318, n9319, n9320,
         n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328, n9329, n9330,
         n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338, n9339, n9340,
         n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348, n9349, n9350,
         n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358, n9359, n9360,
         n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368, n9369, n9370,
         n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378, n9379, n9380,
         n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388, n9389, n9390,
         n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398, n9399, n9400,
         n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408, n9409, n9410,
         n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418, n9419, n9420,
         n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428, n9429, n9430,
         n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438, n9439, n9440,
         n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448, n9449, n9450,
         n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458, n9459, n9460,
         n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468, n9469, n9470,
         n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478, n9479, n9480,
         n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488, n9489, n9490,
         n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498, n9499, n9500,
         n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508, n9509, n9510,
         n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518, n9519, n9520,
         n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528, n9529, n9530,
         n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538, n9539, n9540,
         n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548, n9549, n9550,
         n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558, n9559, n9560,
         n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568, n9569, n9570,
         n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578, n9579, n9580,
         n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588, n9589, n9590,
         n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598, n9599, n9600,
         n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608, n9609, n9610,
         n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618, n9619, n9620,
         n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628, n9629, n9630,
         n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638, n9639, n9640,
         n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648, n9649, n9650,
         n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658, n9659, n9660,
         n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668, n9669, n9670,
         n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678, n9679, n9680,
         n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688, n9689, n9690,
         n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698, n9699, n9700,
         n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708, n9709, n9710,
         n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718, n9719, n9720,
         n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728, n9729, n9730,
         n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738, n9739, n9740,
         n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748, n9749, n9750,
         n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758, n9759, n9760,
         n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768, n9769, n9770,
         n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778, n9779, n9780,
         n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788, n9789, n9790,
         n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798, n9799, n9800,
         n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808, n9809, n9810,
         n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818, n9819, n9820,
         n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828, n9829, n9830,
         n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838, n9839, n9840,
         n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848, n9849, n9850,
         n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858, n9859, n9860,
         n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868, n9869, n9870,
         n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878, n9879, n9880,
         n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888, n9889, n9890,
         n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898, n9899, n9900,
         n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908, n9909, n9910,
         n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918, n9919, n9920,
         n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928, n9929, n9930,
         n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938, n9939, n9940,
         n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948, n9949, n9950,
         n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958, n9959, n9960,
         n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968, n9969, n9970,
         n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978, n9979, n9980,
         n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988, n9989, n9990,
         n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998, n9999, n10000,
         n10001, n10002, n10003, n10004, n10005, n10006, n10007, n10008,
         n10009, n10010, n10011, n10012, n10013, n10014, n10015, n10016,
         n10017, n10018, n10019, n10020, n10021, n10022, n10023, n10024,
         n10025, n10026, n10027, n10028, n10029, n10030, n10031, n10032,
         n10033, n10034, n10035, n10036, n10037, n10038, n10039, n10040,
         n10041, n10042, n10043, n10044, n10045, n10046, n10047, n10048,
         n10049, n10050, n10051, n10052, n10053, n10054, n10055, n10056,
         n10057, n10058, n10059, n10060, n10061, n10062, n10063, n10064,
         n10065, n10066, n10067, n10068, n10069, n10070, n10071, n10072,
         n10073, n10074, n10075, n10076, n10077, n10078, n10079, n10080,
         n10081, n10082, n10083, n10084, n10085, n10086, n10087, n10088,
         n10089, n10090, n10091, n10092, n10093, n10094, n10095, n10096,
         n10097, n10098, n10099, n10100, n10101, n10102, n10103, n10104,
         n10105, n10106, n10107, n10108, n10109, n10110, n10111, n10112,
         n10113, n10114, n10115, n10116, n10117, n10118, n10119, n10120,
         n10121, n10122, n10123, n10124, n10125, n10126, n10127, n10128,
         n10129, n10130, n10131, n10132, n10133, n10134, n10135, n10136,
         n10137, n10138, n10139, n10140, n10141, n10142, n10143, n10144,
         n10145, n10146, n10147, n10148, n10149, n10150, n10151, n10152,
         n10153, n10154, n10155, n10156, n10157, n10158, n10159, n10160,
         n10161, n10162, n10163, n10164, n10165, n10166, n10167, n10168,
         n10169, n10170, n10171, n10172, n10173, n10174, n10175, n10176,
         n10177, n10178, n10179, n10180, n10181, n10182, n10183, n10184,
         n10185, n10186, n10187, n10188, n10189, n10190, n10191, n10192,
         n10193, n10194, n10195, n10196, n10197, n10198, n10199, n10200,
         n10201, n10202, n10203, n10204, n10205, n10206, n10207, n10208,
         n10209, n10210, n10211, n10212, n10213, n10214, n10215, n10216,
         n10217, n10218, n10219, n10220, n10221, n10222, n10223, n10224,
         n10225, n10226, n10227, n10228, n10229, n10230, n10231, n10232,
         n10233, n10234, n10235, n10236, n10237, n10238, n10239, n10240,
         n10241, n10242, n10243, n10244, n10245, n10246, n10247, n10248,
         n10249, n10250, n10251, n10252, n10253, n10254, n10255, n10256,
         n10257, n10258, n10259, n10260, n10261, n10262, n10263, n10264,
         n10265, n10266, n10267, n10268, n10269, n10270, n10271, n10272,
         n10273, n10274, n10275, n10276, n10277, n10278, n10279, n10280,
         n10281, n10282, n10283, n10284, n10285, n10286, n10287, n10288,
         n10289, n10290, n10291, n10292, n10293, n10294, n10295, n10296,
         n10297, n10298, n10299, n10300, n10301, n10302, n10303, n10304,
         n10305, n10306, n10307, n10308, n10309, n10310, n10311, n10312,
         n10313, n10314, n10315, n10316, n10317, n10318, n10319, n10320,
         n10321, n10322, n10323, n10324, n10325, n10326, n10327, n10328,
         n10329, n10330, n10331, n10332, n10333, n10334, n10335, n10336,
         n10337, n10338, n10339, n10340, n10341, n10342, n10343, n10344,
         n10345, n10346, n10347, n10348, n10349, n10350, n10351, n10352,
         n10353, n10354, n10355, n10356, n10357, n10358, n10359, n10360,
         n10361, n10362, n10363, n10364, n10365, n10366, n10367, n10368,
         n10369, n10370, n10371, n10372, n10373, n10374, n10375, n10376,
         n10377, n10378, n10379, n10380, n10381, n10382, n10383, n10384,
         n10385, n10386, n10387, n10388, n10389, n10390, n10391, n10392,
         n10393, n10394, n10395, n10396, n10397, n10398, n10399, n10400,
         n10401, n10402, n10403, n10404, n10405, n10406, n10407, n10408,
         n10409, n10410, n10411, n10412, n10413, n10414, n10415, n10416,
         n10417, n10418, n10419, n10420, n10421, n10422, n10423, n10424,
         n10425, n10426, n10427, n10428, n10429, n10430, n10431, n10432,
         n10433, n10434, n10435, n10436, n10437, n10438, n10439, n10440,
         n10441, n10442, n10443, n10444, n10445, n10446, n10447, n10448,
         n10449, n10450, n10451, n10452, n10453, n10454, n10455, n10456,
         n10457, n10458, n10459, n10460, n10461, n10462, n10463, n10464,
         n10465, n10466, n10467, n10468, n10469, n10470, n10471, n10472,
         n10473, n10474, n10475, n10476, n10477, n10478, n10479, n10480,
         n10481, n10482, n10483, n10484, n10485, n10486, n10487, n10488,
         n10489, n10490, n10491, n10492, n10493, n10494, n10495, n10496,
         n10497, n10498, n10499, n10500, n10501, n10502, n10503, n10504,
         n10505, n10506, n10507, n10508, n10509, n10510, n10511, n10512,
         n10513, n10514, n10515, n10516, n10517, n10518, n10519, n10520,
         n10521, n10522, n10523, n10524, n10525, n10526, n10527, n10528,
         n10529, n10530, n10531, n10532, n10533, n10534, n10535, n10536,
         n10537, n10538, n10539, n10540, n10541, n10542, n10543, n10544,
         n10545, n10546, n10547, n10548, n10549, n10550, n10551, n10552,
         n10553, n10554, n10555, n10556, n10557, n10558, n10559, n10560,
         n10561, n10562, n10563, n10564, n10565, n10566, n10567, n10568,
         n10569, n10570, n10571, n10572, n10573, n10574, n10575, n10576,
         n10577, n10578, n10579, n10580, n10581, n10582, n10583, n10584,
         n10585, n10586, n10587, n10588, n10589, n10590, n10591, n10592,
         n10593, n10594, n10595, n10596, n10597, n10598, n10599, n10600,
         n10601, n10602, n10603, n10604, n10605, n10606, n10607, n10608,
         n10609, n10610, n10611, n10612, n10613, n10614, n10615, n10616,
         n10617, n10618, n10619, n10620, n10621, n10622, n10623, n10624,
         n10625, n10626, n10627, n10628, n10629, n10630, n10631, n10632,
         n10633, n10634, n10635, n10636, n10637, n10638, n10639, n10640,
         n10641, n10642, n10643, n10644, n10645, n10646, n10647, n10648,
         n10649, n10650, n10651, n10652, n10653, n10654, n10655, n10656,
         n10657, n10658, n10659, n10660, n10661, n10662, n10663, n10664,
         n10665, n10666, n10667, n10668, n10669, n10670, n10671, n10672,
         n10673, n10674, n10675, n10676, n10677, n10678, n10679, n10680,
         n10681, n10682, n10683, n10684, n10685, n10686, n10687, n10688,
         n10689, n10690, n10691, n10692, n10693, n10694, n10695, n10696,
         n10697, n10698, n10699, n10700, n10701, n10702, n10703, n10704,
         n10705, n10706, n10707, n10708, n10709, n10710, n10711, n10712,
         n10713, n10714, n10715, n10716, n10717, n10718, n10719, n10720,
         n10721, n10722, n10723, n10724, n10725, n10726, n10727, n10728,
         n10729, n10730, n10731, n10732, n10733, n10734, n10735, n10736,
         n10737, n10738, n10739, n10740, n10741, n10742, n10743, n10744,
         n10745, n10746, n10747, n10748, n10749, n10750, n10751, n10752,
         n10753, n10754, n10755, n10756, n10757, n10758, n10759, n10760,
         n10761, n10762, n10763, n10764, n10765, n10766, n10767, n10768,
         n10769, n10770, n10771, n10772, n10773, n10774, n10775, n10776,
         n10777, n10778, n10779, n10780, n10781, n10782, n10783, n10784,
         n10785, n10786, n10787, n10788, n10789, n10790, n10791, n10792,
         n10793, n10794, n10795, n10796, n10797, n10798, n10799, n10800,
         n10801, n10802, n10803, n10804, n10805, n10806, n10807, n10808,
         n10809, n10810, n10811, n10812, n10813, n10814, n10815, n10816,
         n10817, n10818, n10819, n10820, n10821, n10822, n10823, n10824,
         n10825, n10826, n10827, n10828, n10829, n10830, n10831, n10832,
         n10833, n10834, n10835, n10836, n10837, n10838, n10839, n10840,
         n10841, n10842, n10843, n10844, n10845, n10846, n10847, n10848,
         n10849, n10850, n10851, n10852, n10853, n10854, n10855, n10856,
         n10857, n10858, n10859, n10860, n10861, n10862, n10863, n10864,
         n10865, n10866, n10867, n10868, n10869, n10870, n10871, n10872,
         n10873, n10874, n10875, n10876, n10877, n10878, n10879, n10880,
         n10881, n10882, n10883, n10884, n10885, n10886, n10887, n10888,
         n10889, n10890, n10891, n10892, n10893, n10894, n10895, n10896,
         n10897, n10898, n10899, n10900, n10901, n10902, n10903, n10904,
         n10905, n10906, n10907, n10908, n10909, n10910, n10911, n10912,
         n10913, n10914, n10915, n10916, n10917, n10918, n10919, n10920,
         n10921, n10922, n10923, n10924, n10925, n10926, n10927, n10928,
         n10929, n10930, n10931, n10932, n10933, n10934, n10935, n10936,
         n10937, n10938, n10939, n10940, n10941, n10942, n10943, n10944,
         n10945, n10946, n10947, n10948, n10949, n10950, n10951, n10952,
         n10953, n10954, n10955, n10956, n10957, n10958, n10959, n10960,
         n10961, n10962, n10963, n10964, n10965, n10966, n10967, n10968,
         n10969, n10970, n10971, n10972, n10973, n10974, n10975, n10976,
         n10977, n10978, n10979, n10980, n10981, n10982, n10983, n10984,
         n10985, n10986, n10987, n10988, n10989, n10990, n10991, n10992,
         n10993, n10994, n10995, n10996, n10997, n10998, n10999, n11000,
         n11001, n11002, n11003, n11004, n11005, n11006, n11007, n11008,
         n11009, n11010, n11011, n11012, n11013, n11014, n11015, n11016,
         n11017, n11018, n11019, n11020, n11021, n11022, n11023, n11024,
         n11025, n11026, n11027, n11028, n11029, n11030, n11031, n11032,
         n11033, n11034, n11035, n11036, n11037, n11038, n11039, n11040,
         n11041, n11042, n11043, n11044, n11045, n11046, n11047, n11048,
         n11049, n11050, n11051, n11052, n11053, n11054, n11055, n11056,
         n11057, n11058, n11059, n11060, n11061, n11062, n11063, n11064,
         n11065, n11066, n11067, n11068, n11069, n11070, n11071, n11072,
         n11073, n11074, n11075, n11076, n11077, n11078, n11079, n11080,
         n11081, n11082, n11083, n11084, n11085, n11086, n11087, n11088,
         n11089, n11090, n11091, n11092, n11093, n11094, n11095, n11096,
         n11097, n11098, n11099, n11100, n11101, n11102, n11103, n11104,
         n11105, n11106, n11107, n11108, n11109, n11110, n11111, n11112,
         n11113, n11114, n11115, n11116, n11117, n11118, n11119, n11120,
         n11121, n11122, n11123, n11124, n11125, n11126, n11127, n11128,
         n11129, n11130, n11131, n11132, n11133, n11134, n11135, n11136,
         n11137, n11138, n11139, n11140, n11141, n11142, n11143, n11144,
         n11145, n11146, n11147, n11148, n11149, n11150, n11151, n11152,
         n11153, n11154, n11155, n11156, n11157, n11158, n11159, n11160,
         n11161, n11162, n11163, n11164, n11165, n11166, n11167, n11168,
         n11169, n11170, n11171, n11172, n11173, n11174, n11175, n11176,
         n11177, n11178, n11179, n11180, n11181, n11182, n11183, n11184,
         n11185, n11186, n11187, n11188, n11189, n11190, n11191, n11192,
         n11193, n11194, n11195, n11196, n11197, n11198, n11199, n11200,
         n11201, n11202, n11203, n11204, n11205, n11206, n11207, n11208,
         n11209, n11210, n11211, n11212, n11213, n11214, n11215, n11216,
         n11217, n11218, n11219, n11220, n11221, n11222, n11223, n11224,
         n11225, n11226, n11227, n11228, n11229, n11230, n11231, n11232,
         n11233, n11234, n11235, n11236, n11237, n11238, n11239, n11240,
         n11241, n11242, n11243, n11244, n11245, n11246, n11247, n11248,
         n11249, n11250, n11251, n11252, n11253, n11254, n11255, n11256,
         n11257, n11258, n11259, n11260, n11261, n11262, n11263, n11264,
         n11265, n11266, n11267, n11268, n11269, n11270, n11271, n11272,
         n11273, n11274, n11275, n11276, n11277, n11278, n11279, n11280,
         n11281, n11282, n11283, n11284, n11285, n11286, n11287, n11288,
         n11289, n11290, n11291, n11292, n11293, n11294, n11295, n11296,
         n11297, n11298, n11299, n11300, n11301, n11302, n11303, n11304,
         n11305, n11306, n11307, n11308, n11309, n11310, n11311, n11312,
         n11313, n11314, n11315, n11316, n11317, n11318, n11319, n11320,
         n11321, n11322, n11323, n11324, n11325, n11326, n11327, n11328,
         n11329, n11330, n11331, n11332, n11333, n11334, n11335, n11336,
         n11337, n11338, n11339, n11340, n11341, n11342, n11343, n11344,
         n11345, n11346, n11347, n11348, n11349, n11350, n11351, n11352,
         n11353, n11354, n11355, n11356, n11357, n11358, n11359, n11360,
         n11361, n11362, n11363, n11364, n11365, n11366, n11367, n11368,
         n11369, n11370, n11371, n11372, n11373, n11374, n11375, n11376,
         n11377, n11378, n11379, n11380, n11381, n11382, n11383, n11384,
         n11385, n11386, n11387, n11388, n11389, n11390, n11391, n11392,
         n11393, n11394, n11395, n11396, n11397, n11398, n11399, n11400,
         n11401, n11402, n11403, n11404, n11405, n11406, n11407, n11408,
         n11409, n11410, n11411, n11412, n11413, n11414, n11415, n11416,
         n11417, n11418, n11419, n11420, n11421, n11422, n11423, n11424,
         n11425, n11426, n11427, n11428, n11429, n11430, n11431, n11432,
         n11433, n11434, n11435, n11436, n11437, n11438, n11439, n11440,
         n11441, n11442, n11443, n11444, n11445, n11446, n11447, n11448,
         n11449, n11450, n11451, n11452, n11453, n11454, n11455, n11456,
         n11457, n11458, n11459, n11460, n11461, n11462, n11463, n11464,
         n11465, n11466, n11467, n11468, n11469, n11470, n11471, n11472,
         n11473, n11474, n11475, n11476, n11477, n11478, n11479, n11480,
         n11481, n11482, n11483, n11484, n11485, n11486, n11487, n11488,
         n11489, n11490, n11491, n11492, n11493, n11494, n11495, n11496,
         n11497, n11498, n11499, n11500, n11501, n11502, n11503, n11504,
         n11505, n11506, n11507, n11508, n11509, n11510, n11511, n11512,
         n11513, n11514, n11515, n11516, n11517, n11518, n11519, n11520,
         n11521, n11522, n11523, n11524, n11525, n11526, n11527, n11528,
         n11529, n11530, n11531, n11532, n11533, n11534, n11535, n11536,
         n11537, n11538, n11539, n11540, n11541, n11542, n11543, n11544,
         n11545, n11546, n11547, n11548, n11549, n11550, n11551, n11552,
         n11553, n11554, n11555, n11556, n11557, n11558, n11559, n11560,
         n11561, n11562, n11563, n11564, n11565, n11566, n11567, n11568,
         n11569, n11570, n11571, n11572, n11573, n11574, n11575, n11576,
         n11577, n11578, n11579, n11580, n11581, n11582, n11583, n11584,
         n11585, n11586, n11587, n11588, n11589, n11590, n11591, n11592,
         n11593, n11594, n11595, n11596, n11597, n11598, n11599, n11600,
         n11601, n11602, n11603, n11604, n11605, n11606, n11607, n11608,
         n11609, n11610, n11611, n11612, n11613, n11614, n11615, n11616,
         n11617, n11618, n11619, n11620, n11621, n11622, n11623, n11624,
         n11625, n11626, n11627, n11628, n11629, n11630, n11631, n11632,
         n11633, n11634, n11635, n11636, n11637, n11638, n11639, n11640,
         n11641, n11642, n11643, n11644, n11645, n11646, n11647, n11648,
         n11649, n11650, n11651, n11652, n11653, n11654, n11655, n11656,
         n11657, n11658, n11659, n11660, n11661, n11662, n11663, n11664,
         n11665, n11666, n11667, n11668, n11669, n11670, n11671, n11672,
         n11673, n11674, n11675, n11676, n11677, n11678, n11679, n11680,
         n11681, n11682, n11683, n11684, n11685, n11686, n11687, n11688,
         n11689, n11690, n11691, n11692, n11693, n11694, n11695, n11696,
         n11697, n11698, n11699, n11700, n11701, n11702, n11703, n11704,
         n11705, n11706, n11707, n11708, n11709, n11710, n11711, n11712,
         n11713, n11714, n11715, n11716, n11717, n11718, n11719, n11720,
         n11721, n11722, n11723, n11724, n11725, n11726, n11727, n11728,
         n11729, n11730, n11731, n11732, n11733, n11734, n11735, n11736,
         n11737, n11738, n11739, n11740, n11741, n11742, n11743, n11744,
         n11745, n11746, n11747, n11748, n11749, n11750, n11751, n11752,
         n11753, n11754, n11755, n11756, n11757, n11758, n11759, n11760,
         n11761, n11762, n11763, n11764, n11765, n11766, n11767, n11768,
         n11769, n11770, n11771, n11772, n11773, n11774, n11775, n11776,
         n11777, n11778, n11779, n11780, n11781, n11782, n11783, n11784,
         n11785, n11786, n11787, n11788, n11789, n11790, n11791, n11792,
         n11793, n11794, n11795, n11796, n11797, n11798, n11799, n11800,
         n11801, n11802, n11803, n11804, n11805, n11806, n11807, n11808,
         n11809, n11810, n11811, n11812, n11813, n11814, n11815, n11816,
         n11817, n11818, n11819, n11820, n11821, n11822, n11823, n11824,
         n11825, n11826, n11827, n11828, n11829, n11830, n11831, n11832,
         n11833, n11834, n11835, n11836, n11837, n11838, n11839, n11840,
         n11841, n11842, n11843, n11844, n11845, n11846, n11847, n11848,
         n11849, n11850, n11851, n11852, n11853, n11854, n11855, n11856,
         n11857, n11858, n11859, n11860, n11861, n11862, n11863, n11864,
         n11865, n11866, n11867, n11868, n11869, n11870, n11871, n11872,
         n11873, n11874, n11875, n11876, n11877, n11878, n11879, n11880,
         n11881, n11882, n11883, n11884, n11885, n11886, n11887, n11888,
         n11889, n11890, n11891, n11892, n11893, n11894, n11895, n11896,
         n11897, n11898, n11899, n11900, n11901, n11902, n11903, n11904,
         n11905, n11906, n11907, n11908, n11909, n11910, n11911, n11912,
         n11913, n11914, n11915, n11916, n11917, n11918, n11919, n11920,
         n11921, n11922, n11923, n11924, n11925, n11926, n11927, n11928,
         n11929, n11930, n11931, n11932, n11933, n11934, n11935, n11936,
         n11937, n11938, n11939, n11940, n11941, n11942, n11943, n11944,
         n11945, n11946, n11947, n11948, n11949, n11950, n11951, n11952,
         n11953, n11954, n11955, n11956, n11957, n11958, n11959, n11960,
         n11961, n11962, n11963, n11964, n11965, n11966, n11967, n11968,
         n11969, n11970, n11971, n11972, n11973, n11974, n11975, n11976,
         n11977, n11978, n11979, n11980, n11981, n11982, n11983, n11984,
         n11985, n11986, n11987, n11988, n11989, n11990, n11991, n11992,
         n11993, n11994, n11995, n11996, n11997, n11998, n11999, n12000,
         n12001, n12002, n12003, n12004, n12005, n12006, n12007, n12008,
         n12009, n12010, n12011, n12012, n12013, n12014, n12015, n12016,
         n12017, n12018, n12019, n12020, n12021, n12022, n12023, n12024,
         n12025, n12026, n12027, n12028, n12029, n12030, n12031, n12032,
         n12033, n12034, n12035, n12036, n12037, n12038, n12039, n12040,
         n12041, n12042, n12043, n12044, n12045, n12046, n12047, n12048,
         n12049, n12050, n12051, n12052, n12053, n12054, n12055, n12056,
         n12057, n12058, n12059, n12060, n12061, n12062, n12063, n12064,
         n12065, n12066, n12067, n12068, n12069, n12070, n12071, n12072,
         n12073, n12074, n12075, n12076, n12077, n12078, n12079, n12080,
         n12081, n12082, n12083, n12084, n12085, n12086, n12087, n12088,
         n12089, n12090, n12091, n12092, n12093, n12094, n12095, n12096,
         n12097, n12098, n12099, n12100, n12101, n12102, n12103, n12104,
         n12105, n12106, n12107, n12108, n12109, n12110, n12111, n12112,
         n12113, n12114, n12115, n12116, n12117, n12118, n12119, n12120,
         n12121, n12122, n12123, n12124, n12125, n12126, n12127, n12128,
         n12129, n12130, n12131, n12132, n12133, n12134, n12135, n12136,
         n12137, n12138, n12139, n12140, n12141, n12142, n12143, n12144,
         n12145, n12146, n12147, n12148, n12149, n12150, n12151, n12152,
         n12153, n12154, n12155, n12156, n12157, n12158, n12159, n12160,
         n12161, n12162, n12163, n12164, n12165, n12166, n12167, n12168,
         n12169, n12170, n12171, n12172, n12173, n12174, n12175, n12176,
         n12177, n12178, n12179, n12180, n12181, n12182, n12183, n12184,
         n12185, n12186, n12187, n12188, n12189, n12190, n12191, n12192,
         n12193, n12194, n12195, n12196, n12197, n12198, n12199, n12200,
         n12201, n12202, n12203, n12204, n12205, n12206, n12207, n12208,
         n12209, n12210, n12211, n12212, n12213, n12214, n12215, n12216,
         n12217, n12218, n12219, n12220, n12221, n12222, n12223, n12224,
         n12225, n12226, n12227, n12228, n12229, n12230, n12231, n12232,
         n12233, n12234, n12235, n12236, n12237, n12238, n12239, n12240,
         n12241, n12242, n12243, n12244, n12245, n12246, n12247, n12248,
         n12249, n12250, n12251, n12252, n12253, n12254, n12255, n12256,
         n12257, n12258, n12259, n12260, n12261, n12262, n12263, n12264,
         n12265, n12266, n12267, n12268, n12269, n12270, n12271, n12272,
         n12273, n12274, n12275, n12276, n12277, n12278, n12279, n12280,
         n12281, n12282, n12283, n12284, n12285, n12286, n12287, n12288,
         n12289, n12290, n12291, n12292, n12293, n12294, n12295, n12296,
         n12297, n12298, n12299, n12300, n12301, n12302, n12303, n12304,
         n12305, n12306, n12307, n12308, n12309, n12310, n12311, n12312,
         n12313, n12314, n12315, n12316, n12317, n12318, n12319, n12320,
         n12321, n12322, n12323, n12324, n12325, n12326, n12327, n12328,
         n12329, n12330, n12331, n12332, n12333, n12334, n12335, n12336,
         n12337, n12338, n12339, n12340, n12341, n12342, n12343, n12344,
         n12345, n12346, n12347, n12348, n12349, n12350, n12351, n12352,
         n12353, n12354, n12355, n12356, n12357, n12358, n12359, n12360,
         n12361, n12362, n12363, n12364, n12365, n12366, n12367, n12368,
         n12369, n12370, n12371, n12372, n12373, n12374, n12375, n12376,
         n12377, n12378, n12379, n12380, n12381, n12382, n12383, n12384,
         n12385, n12386, n12387, n12388, n12389, n12390, n12391, n12392,
         n12393, n12394, n12395, n12396, n12397, n12398, n12399, n12400,
         n12401, n12402, n12403, n12404, n12405, n12406, n12407, n12408,
         n12409, n12410, n12411, n12412, n12413, n12414, n12415, n12416,
         n12417, n12418, n12419, n12420, n12421, n12422, n12423, n12424,
         n12425, n12426, n12427, n12428, n12429, n12430, n12431, n12432,
         n12433, n12434, n12435, n12436, n12437, n12438, n12439, n12440,
         n12441, n12442, n12443, n12444, n12445, n12446, n12447, n12448,
         n12449, n12450, n12451, n12452, n12453, n12454, n12455, n12456,
         n12457, n12458, n12459, n12460, n12461, n12462, n12463, n12464,
         n12465, n12466, n12467, n12468, n12469, n12470, n12471, n12472,
         n12473, n12474, n12475, n12476, n12477, n12478, n12479, n12480,
         n12481, n12482, n12483, n12484, n12485, n12486, n12487, n12488,
         n12489, n12490, n12491, n12492, n12493, n12494, n12495, n12496,
         n12497, n12498, n12499, n12500, n12501, n12502, n12503, n12504,
         n12505, n12506, n12507, n12508, n12509, n12510, n12511, n12512,
         n12513, n12514, n12515, n12516, n12517, n12518, n12519, n12520,
         n12521, n12522, n12523, n12524, n12525, n12526, n12527, n12528,
         n12529, n12530, n12531, n12532, n12533, n12534, n12535, n12536,
         n12537, n12538, n12539, n12540, n12541, n12542, n12543, n12544,
         n12545, n12546, n12547, n12548, n12549, n12550, n12551, n12552,
         n12553, n12554, n12555, n12556, n12557, n12558, n12559, n12560,
         n12561, n12562, n12563, n12564, n12565, n12566, n12567, n12568,
         n12569, n12570, n12571, n12572, n12573, n12574, n12575, n12576,
         n12577, n12578, n12579, n12580, n12581, n12582, n12583, n12584,
         n12585, n12586, n12587, n12588, n12589, n12590, n12591, n12592,
         n12593, n12594, n12595, n12596, n12597, n12598, n12599, n12600,
         n12601, n12602, n12603, n12604, n12605, n12606, n12607, n12608,
         n12609, n12610, n12611, n12612, n12613, n12614, n12615, n12616,
         n12617, n12618, n12619, n12620, n12621, n12622, n12623, n12624,
         n12625, n12626, n12627, n12628, n12629, n12630, n12631, n12632,
         n12633, n12634, n12635, n12636, n12637, n12638, n12639, n12640,
         n12641, n12642, n12643, n12644, n12645, n12646, n12647, n12648,
         n12649, n12650, n12651, n12652, n12653, n12654, n12655, n12656,
         n12657, n12658, n12659, n12660, n12661, n12662, n12663, n12664,
         n12665, n12666, n12667, n12668, n12669, n12670, n12671, n12672,
         n12673, n12674, n12675, n12676, n12677, n12678, n12679, n12680,
         n12681, n12682, n12683, n12684, n12685, n12686, n12687, n12688,
         n12689, n12690, n12691, n12692, n12693, n12694, n12695, n12696,
         n12697, n12698, n12699, n12700, n12701, n12702, n12703, n12704,
         n12705, n12706, n12707, n12708, n12709, n12710, n12711, n12712,
         n12713, n12714, n12715, n12716, n12717, n12718, n12719, n12720,
         n12721, n12722, n12723, n12724, n12725, n12726, n12727, n12728,
         n12729, n12730, n12731, n12732, n12733, n12734, n12735, n12736,
         n12737, n12738, n12739, n12740, n12741, n12742, n12743, n12744,
         n12745, n12746, n12747, n12748, n12749, n12750, n12751, n12752,
         n12753, n12754, n12755, n12756, n12757, n12758, n12759, n12760,
         n12761, n12762, n12763, n12764, n12765, n12766, n12767, n12768,
         n12769, n12770, n12771, n12772, n12773, n12774, n12775, n12776,
         n12777, n12778, n12779, n12780, n12781, n12782, n12783, n12784,
         n12785, n12786, n12787, n12788, n12789, n12790, n12791, n12792,
         n12793, n12794, n12795, n12796, n12797, n12798, n12799, n12800,
         n12801, n12802, n12803, n12804, n12805, n12806, n12807, n12808,
         n12809, n12810, n12811, n12812, n12813, n12814, n12815, n12816,
         n12817, n12818, n12819, n12820, n12821, n12822, n12823;
  wire   [29:0] ICACHE_addr;
  assign mem_write_D = net109179;
  assign DCACHE_addr[3] = net113537;
  assign DCACHE_wdata[6] = net139803;

  DFFRX4 \i_MIPS/ID_EX_reg[7]  ( .D(\i_MIPS/n471 ), .CK(clk), .RN(n5609), .Q(
        \i_MIPS/ALUOp[1] ), .QN(n3526) );
  DFFRX4 \i_MIPS/ID_EX_reg[5]  ( .D(\i_MIPS/n478 ), .CK(clk), .RN(n5610), .Q(
        \i_MIPS/ID_EX_5 ) );
  DFFRX4 \i_MIPS/ID_EX_reg[83]  ( .D(\i_MIPS/n502 ), .CK(clk), .RN(n5612), .Q(
        \i_MIPS/ID_EX[83] ), .QN(n4704) );
  DFFRX4 \i_MIPS/ID_EX_reg[82]  ( .D(\i_MIPS/n503 ), .CK(clk), .RN(n5612), .Q(
        \i_MIPS/ID_EX[82] ), .QN(n4707) );
  DFFRX4 \i_MIPS/ID_EX_reg[81]  ( .D(\i_MIPS/n504 ), .CK(clk), .RN(n5612), .Q(
        \i_MIPS/ID_EX[81] ), .QN(n3787) );
  DFFRX4 \i_MIPS/ID_EX_reg[80]  ( .D(\i_MIPS/n505 ), .CK(clk), .RN(n5612), .Q(
        \i_MIPS/ID_EX[80] ), .QN(n4706) );
  DFFRX4 \i_MIPS/ID_EX_reg[78]  ( .D(\i_MIPS/n507 ), .CK(clk), .RN(n5612), .Q(
        \i_MIPS/ID_EX[78] ), .QN(n4641) );
  DFFRX4 \i_MIPS/ID_EX_reg[75]  ( .D(\i_MIPS/n510 ), .CK(clk), .RN(n5612), .Q(
        \i_MIPS/ID_EX[75] ), .QN(n3755) );
  DFFRX4 \i_MIPS/ID_EX_reg[73]  ( .D(\i_MIPS/n512 ), .CK(clk), .RN(n5613), .Q(
        \i_MIPS/ID_EX[73] ), .QN(n3800) );
  DFFRX4 \i_MIPS/IF_ID_reg[48]  ( .D(\i_MIPS/N71 ), .CK(clk), .RN(n5614), .Q(
        \i_MIPS/IR_ID[16] ), .QN(\i_MIPS/n312 ) );
  DFFRX4 \i_MIPS/IF_ID_reg[51]  ( .D(\i_MIPS/N74 ), .CK(clk), .RN(n5614), .Q(
        \i_MIPS/IR_ID[19] ), .QN(\i_MIPS/n318 ) );
  DFFRX4 \i_MIPS/IF_ID_reg[54]  ( .D(\i_MIPS/N77 ), .CK(clk), .RN(n5615), .Q(
        \i_MIPS/IR_ID[22] ), .QN(\i_MIPS/n229 ) );
  DFFRX4 \i_MIPS/IF_ID_reg[55]  ( .D(\i_MIPS/N78 ), .CK(clk), .RN(n5615), .Q(
        \i_MIPS/IR_ID[23] ), .QN(\i_MIPS/n230 ) );
  DFFRX4 \i_MIPS/IF_ID_reg[57]  ( .D(\i_MIPS/N80 ), .CK(clk), .RN(n5615), .Q(
        \i_MIPS/IR_ID[25] ), .QN(\i_MIPS/n232 ) );
  DFFRX4 \i_MIPS/ID_EX_reg[24]  ( .D(\i_MIPS/n547 ), .CK(clk), .RN(n5618), .Q(
        \i_MIPS/ALUin1[15] ), .QN(\i_MIPS/n356 ) );
  DFFRX4 \i_MIPS/ID_EX_reg[18]  ( .D(\i_MIPS/n553 ), .CK(clk), .RN(n5619), .Q(
        \i_MIPS/ALUin1[9] ), .QN(\i_MIPS/n362 ) );
  DFFRX4 \i_MIPS/ID_EX_reg[15]  ( .D(\i_MIPS/n556 ), .CK(clk), .RN(n5619), .Q(
        \i_MIPS/ALUin1[6] ), .QN(\i_MIPS/n365 ) );
  DFFRX4 \i_MIPS/ID_EX_reg[14]  ( .D(\i_MIPS/n557 ), .CK(clk), .RN(n5619), .Q(
        \i_MIPS/ALUin1[5] ), .QN(\i_MIPS/n366 ) );
  DFFRX4 \i_MIPS/ID_EX_reg[13]  ( .D(\i_MIPS/n558 ), .CK(clk), .RN(n5619), .Q(
        \i_MIPS/ALUin1[4] ), .QN(\i_MIPS/n367 ) );
  NAND4BX4 \i_MIPS/ALU_Control/U16  ( .AN(\i_MIPS/ID_EX[106] ), .B(
        \i_MIPS/ID_EX[105] ), .C(\i_MIPS/ID_EX[107] ), .D(
        \i_MIPS/ALU_Control/n11 ), .Y(\i_MIPS/ALU_Control/n20 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[30]  ( .D(\i_MIPS/n444 ), .CK(clk), .RN(n5607), 
        .Q(n12945), .QN(n4754) );
  DFFRX1 \i_MIPS/EX_MEM_reg[22]  ( .D(\i_MIPS/n452 ), .CK(clk), .RN(n5608), 
        .Q(n12953), .QN(n4752) );
  DFFRX1 \i_MIPS/EX_MEM_reg[17]  ( .D(\i_MIPS/n457 ), .CK(clk), .RN(n5608), 
        .Q(n12958), .QN(n4748) );
  DFFRX1 \i_MIPS/EX_MEM_reg[23]  ( .D(\i_MIPS/n451 ), .CK(clk), .RN(n5607), 
        .Q(n12952), .QN(n1877) );
  DFFRX1 \i_MIPS/EX_MEM_reg[36]  ( .D(\i_MIPS/n438 ), .CK(clk), .RN(n5606), 
        .Q(n12939) );
  DFFRX1 \i_MIPS/IF_ID_reg[40]  ( .D(\i_MIPS/N63 ), .CK(clk), .RN(n5613), .Q(
        \i_MIPS/Sign_Extend_ID[8] ), .QN(\i_MIPS/n220 ) );
  DFFRX1 \i_MIPS/Pred_2bit/current_state_reg[0]  ( .D(\i_MIPS/Pred_2bit/n8 ), 
        .CK(clk), .RN(n5620), .Q(\i_MIPS/Pred_2bit/current_state[0] ), .QN(
        \i_MIPS/Pred_2bit/n1 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[5]  ( .D(\i_MIPS/N28 ), .CK(clk), .RN(n5600), .QN(
        \i_MIPS/n185 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[86]  ( .D(\i_MIPS/N109 ), .CK(clk), .RN(n5596), .Q(
        \i_MIPS/IF_ID[86] ), .QN(\i_MIPS/n168 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[82]  ( .D(\i_MIPS/N105 ), .CK(clk), .RN(n5597), .Q(
        \i_MIPS/IF_ID[82] ), .QN(\i_MIPS/n164 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[78]  ( .D(\i_MIPS/N101 ), .CK(clk), .RN(n5597), .Q(
        \i_MIPS/IF_ID[78] ), .QN(\i_MIPS/n160 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[93]  ( .D(\i_MIPS/N116 ), .CK(clk), .RN(n5596), .Q(
        \i_MIPS/IF_ID[93] ), .QN(\i_MIPS/n175 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[85]  ( .D(\i_MIPS/N108 ), .CK(clk), .RN(n5597), .Q(
        \i_MIPS/IF_ID[85] ), .QN(\i_MIPS/n167 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[4]  ( .D(\i_MIPS/n480 ), .CK(clk), .RN(n5610), .Q(
        n3507), .QN(\i_MIPS/n311 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[1]  ( .D(\i_MIPS/n527 ), .CK(clk), .RN(n5616), .Q(
        n3504), .QN(\i_MIPS/n337 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[116]  ( .D(\i_MIPS/n530 ), .CK(clk), .RN(n5617), 
        .Q(n3505), .QN(\i_MIPS/n339 ) );
  DFFSX1 \i_MIPS/Pred_2bit/current_state_reg[1]  ( .D(\i_MIPS/Pred_2bit/n7 ), 
        .CK(clk), .SN(n5914), .Q(\i_MIPS/Pred_2bit/current_state[1] ), .QN(
        n4699) );
  DFFRX1 \i_MIPS/ID_EX_reg[3]  ( .D(\i_MIPS/n525 ), .CK(clk), .RN(n5616), .Q(
        \i_MIPS/ID_EX_3 ), .QN(\i_MIPS/n335 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[74]  ( .D(\i_MIPS/n529 ), .CK(clk), .RN(n5617), 
        .Q(\i_MIPS/EX_MEM_74 ), .QN(\i_MIPS/n338 ) );
  DFFRX1 \i_MIPS/Register/register_reg[28][0]  ( .D(\i_MIPS/Register/n212 ), 
        .CK(clk), .RN(n5630), .Q(\i_MIPS/Register/register[28][0] ), .QN(n298)
         );
  DFFRX1 \i_MIPS/Register/register_reg[24][0]  ( .D(\i_MIPS/Register/n340 ), 
        .CK(clk), .RN(n5641), .Q(\i_MIPS/Register/register[24][0] ), .QN(n296)
         );
  DFFRX1 \i_MIPS/Register/register_reg[20][0]  ( .D(\i_MIPS/Register/n468 ), 
        .CK(clk), .RN(n5652), .Q(\i_MIPS/Register/register[20][0] ), .QN(n1871) );
  DFFRX1 \i_MIPS/Register/register_reg[16][0]  ( .D(\i_MIPS/Register/n596 ), 
        .CK(clk), .RN(n5662), .Q(\i_MIPS/Register/register[16][0] ), .QN(n1869) );
  DFFRX1 \i_MIPS/Register/register_reg[15][1]  ( .D(\i_MIPS/Register/n629 ), 
        .CK(clk), .RN(n5665), .Q(\i_MIPS/Register/register[15][1] ), .QN(n198)
         );
  DFFRX1 \i_MIPS/Register/register_reg[12][0]  ( .D(\i_MIPS/Register/n724 ), 
        .CK(clk), .RN(n5673), .Q(\i_MIPS/Register/register[12][0] ), .QN(n299)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][0]  ( .D(\i_MIPS/Register/n852 ), 
        .CK(clk), .RN(n5684), .Q(\i_MIPS/Register/register[8][0] ), .QN(n297)
         );
  DFFRX1 \i_MIPS/Register/register_reg[4][0]  ( .D(\i_MIPS/Register/n980 ), 
        .CK(clk), .RN(n5694), .Q(\i_MIPS/Register/register[4][0] ), .QN(n1872)
         );
  DFFRX1 \i_MIPS/Register/register_reg[0][0]  ( .D(\i_MIPS/Register/n1108 ), 
        .CK(clk), .RN(n5705), .Q(\i_MIPS/Register/register[0][0] ), .QN(n1870)
         );
  DFFRX1 \i_MIPS/Register/register_reg[31][8]  ( .D(n11572), .CK(clk), .RN(
        n5623), .Q(\i_MIPS/Register/register[31][8] ), .QN(n226) );
  DFFRX1 \i_MIPS/Register/register_reg[31][9]  ( .D(n11571), .CK(clk), .RN(
        n5623), .Q(\i_MIPS/Register/register[31][9] ), .QN(n225) );
  DFFRX1 \i_MIPS/Register/register_reg[31][12]  ( .D(n11568), .CK(clk), .RN(
        n5623), .Q(\i_MIPS/Register/register[31][12] ), .QN(n237) );
  DFFRX1 \i_MIPS/Register/register_reg[31][15]  ( .D(n11565), .CK(clk), .RN(
        n5624), .Q(\i_MIPS/Register/register[31][15] ), .QN(n239) );
  DFFRX1 \i_MIPS/Register/register_reg[31][17]  ( .D(n11563), .CK(clk), .RN(
        n5624), .Q(\i_MIPS/Register/register[31][17] ), .QN(n189) );
  DFFRX1 \i_MIPS/Register/register_reg[31][31]  ( .D(n11549), .CK(clk), .RN(
        n5625), .Q(\i_MIPS/Register/register[31][31] ), .QN(n190) );
  DFFRX1 \i_MIPS/EX_MEM_reg[6]  ( .D(\i_MIPS/n468 ), .CK(clk), .RN(n5609), .Q(
        \i_MIPS/EX_MEM[6] ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[5]  ( .D(\i_MIPS/n469 ), .CK(clk), .RN(n5609), .Q(
        \i_MIPS/EX_MEM[5] ), .QN(n4710) );
  DFFRX1 \I_cache/cache_reg[0][16]  ( .D(n12695), .CK(clk), .RN(n5822), .Q(
        \I_cache/cache[0][16] ), .QN(n1701) );
  DFFRX1 \I_cache/cache_reg[1][16]  ( .D(n12694), .CK(clk), .RN(n5822), .Q(
        \I_cache/cache[1][16] ), .QN(n3385) );
  DFFRX1 \I_cache/cache_reg[2][16]  ( .D(n12693), .CK(clk), .RN(n5822), .Q(
        \I_cache/cache[2][16] ), .QN(n1702) );
  DFFRX1 \I_cache/cache_reg[5][16]  ( .D(n12690), .CK(clk), .RN(n5822), .Q(
        \I_cache/cache[5][16] ), .QN(n3415) );
  DFFRX1 \I_cache/cache_reg[6][16]  ( .D(n12689), .CK(clk), .RN(n5822), .Q(
        \I_cache/cache[6][16] ), .QN(n1703) );
  DFFRX1 \I_cache/cache_reg[7][16]  ( .D(n12688), .CK(clk), .RN(n5822), .Q(
        \I_cache/cache[7][16] ), .QN(n3387) );
  DFFRX1 \I_cache/cache_reg[0][17]  ( .D(n12687), .CK(clk), .RN(n5822), .Q(
        \I_cache/cache[0][17] ), .QN(n1782) );
  DFFRX1 \I_cache/cache_reg[1][17]  ( .D(n12686), .CK(clk), .RN(n5822), .Q(
        \I_cache/cache[1][17] ), .QN(n3466) );
  DFFRX1 \I_cache/cache_reg[2][17]  ( .D(n12685), .CK(clk), .RN(n5822), .Q(
        \I_cache/cache[2][17] ), .QN(n1783) );
  DFFRX1 \I_cache/cache_reg[3][17]  ( .D(n12684), .CK(clk), .RN(n5823), .Q(
        \I_cache/cache[3][17] ), .QN(n3467) );
  DFFRX1 \I_cache/cache_reg[4][17]  ( .D(n12683), .CK(clk), .RN(n5823), .Q(
        \I_cache/cache[4][17] ), .QN(n1796) );
  DFFRX1 \I_cache/cache_reg[5][17]  ( .D(n12682), .CK(clk), .RN(n5823), .Q(
        \I_cache/cache[5][17] ), .QN(n3480) );
  DFFRX1 \I_cache/cache_reg[6][17]  ( .D(n12681), .CK(clk), .RN(n5823), .Q(
        \I_cache/cache[6][17] ), .QN(n1784) );
  DFFRX1 \I_cache/cache_reg[7][17]  ( .D(n12680), .CK(clk), .RN(n5823), .Q(
        \I_cache/cache[7][17] ), .QN(n3468) );
  DFFRX1 \I_cache/cache_reg[0][18]  ( .D(n12679), .CK(clk), .RN(n5823), .Q(
        \I_cache/cache[0][18] ), .QN(n1689) );
  DFFRX1 \I_cache/cache_reg[1][18]  ( .D(n12678), .CK(clk), .RN(n5823), .Q(
        \I_cache/cache[1][18] ), .QN(n3373) );
  DFFRX1 \I_cache/cache_reg[2][18]  ( .D(n12677), .CK(clk), .RN(n5823), .Q(
        \I_cache/cache[2][18] ), .QN(n1690) );
  DFFRX1 \I_cache/cache_reg[3][18]  ( .D(n12676), .CK(clk), .RN(n5823), .Q(
        \I_cache/cache[3][18] ), .QN(n3374) );
  DFFRX1 \I_cache/cache_reg[4][18]  ( .D(n12675), .CK(clk), .RN(n5823), .Q(
        \I_cache/cache[4][18] ), .QN(n1727) );
  DFFRX1 \I_cache/cache_reg[5][18]  ( .D(n12674), .CK(clk), .RN(n5823), .Q(
        \I_cache/cache[5][18] ), .QN(n3411) );
  DFFRX1 \I_cache/cache_reg[6][18]  ( .D(n12673), .CK(clk), .RN(n5823), .Q(
        \I_cache/cache[6][18] ), .QN(n1691) );
  DFFRX1 \I_cache/cache_reg[7][18]  ( .D(n12672), .CK(clk), .RN(n5824), .Q(
        \I_cache/cache[7][18] ), .QN(n3375) );
  DFFRX1 \I_cache/cache_reg[0][19]  ( .D(n12671), .CK(clk), .RN(n5824), .Q(
        \I_cache/cache[0][19] ), .QN(n1776) );
  DFFRX1 \I_cache/cache_reg[1][19]  ( .D(n12670), .CK(clk), .RN(n5824), .Q(
        \I_cache/cache[1][19] ), .QN(n3460) );
  DFFRX1 \I_cache/cache_reg[2][19]  ( .D(n12669), .CK(clk), .RN(n5824), .Q(
        \I_cache/cache[2][19] ), .QN(n1777) );
  DFFRX1 \I_cache/cache_reg[3][19]  ( .D(n12668), .CK(clk), .RN(n5824), .Q(
        \I_cache/cache[3][19] ), .QN(n3461) );
  DFFRX1 \I_cache/cache_reg[4][19]  ( .D(n12667), .CK(clk), .RN(n5824), .Q(
        \I_cache/cache[4][19] ), .QN(n1791) );
  DFFRX1 \I_cache/cache_reg[5][19]  ( .D(n12666), .CK(clk), .RN(n5824), .Q(
        \I_cache/cache[5][19] ), .QN(n3475) );
  DFFRX1 \I_cache/cache_reg[6][19]  ( .D(n12665), .CK(clk), .RN(n5824), .Q(
        \I_cache/cache[6][19] ), .QN(n1778) );
  DFFRX1 \I_cache/cache_reg[7][19]  ( .D(n12664), .CK(clk), .RN(n5824), .Q(
        \I_cache/cache[7][19] ), .QN(n3462) );
  DFFRX1 \I_cache/cache_reg[0][20]  ( .D(n12663), .CK(clk), .RN(n5824), .Q(
        \I_cache/cache[0][20] ), .QN(n1674) );
  DFFRX1 \I_cache/cache_reg[1][20]  ( .D(n12662), .CK(clk), .RN(n5824), .Q(
        \I_cache/cache[1][20] ), .QN(n3358) );
  DFFRX1 \I_cache/cache_reg[2][20]  ( .D(n12661), .CK(clk), .RN(n5824), .Q(
        \I_cache/cache[2][20] ), .QN(n1675) );
  DFFRX1 \I_cache/cache_reg[3][20]  ( .D(n12660), .CK(clk), .RN(n5825), .Q(
        \I_cache/cache[3][20] ), .QN(n3359) );
  DFFRX1 \I_cache/cache_reg[4][20]  ( .D(n12659), .CK(clk), .RN(n5825), .Q(
        \I_cache/cache[4][20] ), .QN(n1722) );
  DFFRX1 \I_cache/cache_reg[5][20]  ( .D(n12658), .CK(clk), .RN(n5825), .Q(
        \I_cache/cache[5][20] ), .QN(n3406) );
  DFFRX1 \I_cache/cache_reg[6][20]  ( .D(n12657), .CK(clk), .RN(n5825), .Q(
        \I_cache/cache[6][20] ), .QN(n1676) );
  DFFRX1 \I_cache/cache_reg[7][20]  ( .D(n12656), .CK(clk), .RN(n5825), .Q(
        \I_cache/cache[7][20] ), .QN(n3360) );
  DFFRX1 \I_cache/cache_reg[0][21]  ( .D(n12655), .CK(clk), .RN(n5825), .Q(
        \I_cache/cache[0][21] ), .QN(n1662) );
  DFFRX1 \I_cache/cache_reg[1][21]  ( .D(n12654), .CK(clk), .RN(n5825), .Q(
        \I_cache/cache[1][21] ), .QN(n3346) );
  DFFRX1 \I_cache/cache_reg[2][21]  ( .D(n12653), .CK(clk), .RN(n5825), .Q(
        \I_cache/cache[2][21] ), .QN(n1663) );
  DFFRX1 \I_cache/cache_reg[3][21]  ( .D(n12652), .CK(clk), .RN(n5825), .Q(
        \I_cache/cache[3][21] ), .QN(n3347) );
  DFFRX1 \I_cache/cache_reg[4][21]  ( .D(n12651), .CK(clk), .RN(n5825), .Q(
        \I_cache/cache[4][21] ), .QN(n1718) );
  DFFRX1 \I_cache/cache_reg[5][21]  ( .D(n12650), .CK(clk), .RN(n5825), .Q(
        \I_cache/cache[5][21] ), .QN(n3402) );
  DFFRX1 \I_cache/cache_reg[6][21]  ( .D(n12649), .CK(clk), .RN(n5825), .Q(
        \I_cache/cache[6][21] ), .QN(n1664) );
  DFFRX1 \I_cache/cache_reg[7][21]  ( .D(n12648), .CK(clk), .RN(n5826), .Q(
        \I_cache/cache[7][21] ), .QN(n3348) );
  DFFRX1 \I_cache/cache_reg[0][22]  ( .D(n12647), .CK(clk), .RN(n5826), .Q(
        \I_cache/cache[0][22] ), .QN(n1773) );
  DFFRX1 \I_cache/cache_reg[1][22]  ( .D(n12646), .CK(clk), .RN(n5826), .Q(
        \I_cache/cache[1][22] ), .QN(n3457) );
  DFFRX1 \I_cache/cache_reg[2][22]  ( .D(n12645), .CK(clk), .RN(n5826), .Q(
        \I_cache/cache[2][22] ), .QN(n1774) );
  DFFRX1 \I_cache/cache_reg[3][22]  ( .D(n12644), .CK(clk), .RN(n5826), .Q(
        \I_cache/cache[3][22] ), .QN(n3458) );
  DFFRX1 \I_cache/cache_reg[4][22]  ( .D(n12643), .CK(clk), .RN(n5826), .Q(
        \I_cache/cache[4][22] ), .QN(n1789) );
  DFFRX1 \I_cache/cache_reg[5][22]  ( .D(n12642), .CK(clk), .RN(n5826), .Q(
        \I_cache/cache[5][22] ), .QN(n3473) );
  DFFRX1 \I_cache/cache_reg[6][22]  ( .D(n12641), .CK(clk), .RN(n5826), .Q(
        \I_cache/cache[6][22] ), .QN(n1775) );
  DFFRX1 \I_cache/cache_reg[7][22]  ( .D(n12640), .CK(clk), .RN(n5826), .Q(
        \I_cache/cache[7][22] ), .QN(n3459) );
  DFFRX1 \I_cache/cache_reg[0][23]  ( .D(n12639), .CK(clk), .RN(n5826), .Q(
        \I_cache/cache[0][23] ), .QN(n1650) );
  DFFRX1 \I_cache/cache_reg[1][23]  ( .D(n12638), .CK(clk), .RN(n5826), .Q(
        \I_cache/cache[1][23] ), .QN(n3334) );
  DFFRX1 \I_cache/cache_reg[2][23]  ( .D(n12637), .CK(clk), .RN(n5826), .Q(
        \I_cache/cache[2][23] ), .QN(n1651) );
  DFFRX1 \I_cache/cache_reg[3][23]  ( .D(n12636), .CK(clk), .RN(n5827), .Q(
        \I_cache/cache[3][23] ), .QN(n3335) );
  DFFRX1 \I_cache/cache_reg[4][23]  ( .D(n12635), .CK(clk), .RN(n5827), .Q(
        \I_cache/cache[4][23] ), .QN(n1714) );
  DFFRX1 \I_cache/cache_reg[5][23]  ( .D(n12634), .CK(clk), .RN(n5827), .Q(
        \I_cache/cache[5][23] ), .QN(n3398) );
  DFFRX1 \I_cache/cache_reg[6][23]  ( .D(n12633), .CK(clk), .RN(n5827), .Q(
        \I_cache/cache[6][23] ), .QN(n1652) );
  DFFRX1 \I_cache/cache_reg[7][23]  ( .D(n12632), .CK(clk), .RN(n5827), .Q(
        \I_cache/cache[7][23] ), .QN(n3336) );
  DFFRX1 \I_cache/cache_reg[0][24]  ( .D(n12631), .CK(clk), .RN(n5827), .Q(
        \I_cache/cache[0][24] ), .QN(n1638) );
  DFFRX1 \I_cache/cache_reg[1][24]  ( .D(n12630), .CK(clk), .RN(n5827), .Q(
        \I_cache/cache[1][24] ), .QN(n3322) );
  DFFRX1 \I_cache/cache_reg[2][24]  ( .D(n12629), .CK(clk), .RN(n5827), .Q(
        \I_cache/cache[2][24] ), .QN(n1639) );
  DFFRX1 \I_cache/cache_reg[3][24]  ( .D(n12628), .CK(clk), .RN(n5827), .Q(
        \I_cache/cache[3][24] ), .QN(n3323) );
  DFFRX1 \I_cache/cache_reg[4][24]  ( .D(n12627), .CK(clk), .RN(n5827), .Q(
        \I_cache/cache[4][24] ), .QN(n1710) );
  DFFRX1 \I_cache/cache_reg[5][24]  ( .D(n12626), .CK(clk), .RN(n5827), .Q(
        \I_cache/cache[5][24] ), .QN(n3394) );
  DFFRX1 \I_cache/cache_reg[6][24]  ( .D(n12625), .CK(clk), .RN(n5827), .Q(
        \I_cache/cache[6][24] ), .QN(n1640) );
  DFFRX1 \I_cache/cache_reg[7][24]  ( .D(n12624), .CK(clk), .RN(n5828), .Q(
        \I_cache/cache[7][24] ), .QN(n3324) );
  DFFRX1 \I_cache/cache_reg[0][25]  ( .D(n12623), .CK(clk), .RN(n5828), .Q(
        \I_cache/cache[0][25] ), .QN(n1764) );
  DFFRX1 \I_cache/cache_reg[1][25]  ( .D(n12622), .CK(clk), .RN(n5828), .Q(
        \I_cache/cache[1][25] ), .QN(n3448) );
  DFFRX1 \I_cache/cache_reg[2][25]  ( .D(n12621), .CK(clk), .RN(n5828), .Q(
        \I_cache/cache[2][25] ), .QN(n1765) );
  DFFRX1 \I_cache/cache_reg[3][25]  ( .D(n12620), .CK(clk), .RN(n5828), .Q(
        \I_cache/cache[3][25] ), .QN(n3449) );
  DFFRX1 \I_cache/cache_reg[4][25]  ( .D(n12619), .CK(clk), .RN(n5828), .Q(
        \I_cache/cache[4][25] ), .QN(n1785) );
  DFFRX1 \I_cache/cache_reg[6][25]  ( .D(n12617), .CK(clk), .RN(n5828), .Q(
        \I_cache/cache[6][25] ), .QN(n1766) );
  DFFRX1 \I_cache/cache_reg[0][26]  ( .D(n12615), .CK(clk), .RN(n5828), .Q(
        \I_cache/cache[0][26] ), .QN(n2509) );
  DFFRX1 \I_cache/cache_reg[1][26]  ( .D(n12614), .CK(clk), .RN(n5828), .Q(
        \I_cache/cache[1][26] ), .QN(n758) );
  DFFRX1 \I_cache/cache_reg[2][26]  ( .D(n12613), .CK(clk), .RN(n5828), .Q(
        \I_cache/cache[2][26] ), .QN(n2510) );
  DFFRX1 \I_cache/cache_reg[3][26]  ( .D(n12612), .CK(clk), .RN(n5829), .Q(
        \I_cache/cache[3][26] ), .QN(n759) );
  DFFRX1 \I_cache/cache_reg[4][26]  ( .D(n12611), .CK(clk), .RN(n5829), .Q(
        \I_cache/cache[4][26] ), .QN(n1211) );
  DFFRX1 \I_cache/cache_reg[5][26]  ( .D(n12610), .CK(clk), .RN(n5829), .Q(
        \I_cache/cache[5][26] ), .QN(n2783) );
  DFFRX1 \I_cache/cache_reg[6][26]  ( .D(n12609), .CK(clk), .RN(n5829), .Q(
        \I_cache/cache[6][26] ), .QN(n2511) );
  DFFRX1 \I_cache/cache_reg[7][26]  ( .D(n12608), .CK(clk), .RN(n5829), .Q(
        \I_cache/cache[7][26] ), .QN(n760) );
  DFFRX1 \I_cache/cache_reg[0][27]  ( .D(n12607), .CK(clk), .RN(n5829), .Q(
        \I_cache/cache[0][27] ), .QN(n1168) );
  DFFRX1 \I_cache/cache_reg[1][27]  ( .D(n12606), .CK(clk), .RN(n5829), .Q(
        \I_cache/cache[1][27] ), .QN(n2740) );
  DFFRX1 \I_cache/cache_reg[2][27]  ( .D(n12605), .CK(clk), .RN(n5829), .Q(
        \I_cache/cache[2][27] ), .QN(n1169) );
  DFFRX1 \I_cache/cache_reg[3][27]  ( .D(n12604), .CK(clk), .RN(n5829), .Q(
        \I_cache/cache[3][27] ), .QN(n2741) );
  DFFRX1 \I_cache/cache_reg[4][27]  ( .D(n12603), .CK(clk), .RN(n5829), .Q(
        \I_cache/cache[4][27] ), .QN(n1216) );
  DFFRX1 \I_cache/cache_reg[5][27]  ( .D(n12602), .CK(clk), .RN(n5829), .Q(
        \I_cache/cache[5][27] ), .QN(n2788) );
  DFFRX1 \I_cache/cache_reg[6][27]  ( .D(n12601), .CK(clk), .RN(n5829), .Q(
        \I_cache/cache[6][27] ), .QN(n1170) );
  DFFRX1 \I_cache/cache_reg[7][27]  ( .D(n12600), .CK(clk), .RN(n5830), .Q(
        \I_cache/cache[7][27] ), .QN(n2742) );
  DFFRX1 \I_cache/cache_reg[0][28]  ( .D(n12599), .CK(clk), .RN(n5830), .Q(
        \I_cache/cache[0][28] ), .QN(n1074) );
  DFFRX1 \I_cache/cache_reg[1][28]  ( .D(n12598), .CK(clk), .RN(n5830), .Q(
        \I_cache/cache[1][28] ), .QN(n2646) );
  DFFRX1 \I_cache/cache_reg[2][28]  ( .D(n12597), .CK(clk), .RN(n5830), .Q(
        \I_cache/cache[2][28] ), .QN(n981) );
  DFFRX1 \I_cache/cache_reg[3][28]  ( .D(n12596), .CK(clk), .RN(n5830), .Q(
        \I_cache/cache[3][28] ), .QN(n2529) );
  DFFRX1 \I_cache/cache_reg[4][28]  ( .D(n12595), .CK(clk), .RN(n5830), .Q(
        \I_cache/cache[4][28] ), .QN(n1210) );
  DFFRX1 \I_cache/cache_reg[5][28]  ( .D(n12594), .CK(clk), .RN(n5830), .Q(
        \I_cache/cache[5][28] ), .QN(n2782) );
  DFFRX1 \I_cache/cache_reg[6][28]  ( .D(n12593), .CK(clk), .RN(n5830), .Q(
        \I_cache/cache[6][28] ), .QN(n982) );
  DFFRX1 \I_cache/cache_reg[7][28]  ( .D(n12592), .CK(clk), .RN(n5830), .Q(
        \I_cache/cache[7][28] ), .QN(n2530) );
  DFFRX1 \I_cache/cache_reg[0][29]  ( .D(n12591), .CK(clk), .RN(n5830), .Q(
        \I_cache/cache[0][29] ), .QN(n1073) );
  DFFRX1 \I_cache/cache_reg[1][29]  ( .D(n12590), .CK(clk), .RN(n5830), .Q(
        \I_cache/cache[1][29] ), .QN(n2645) );
  DFFRX1 \I_cache/cache_reg[2][29]  ( .D(n12589), .CK(clk), .RN(n5830), .Q(
        \I_cache/cache[2][29] ), .QN(n980) );
  DFFRX1 \I_cache/cache_reg[3][29]  ( .D(n12588), .CK(clk), .RN(n5831), .Q(
        \I_cache/cache[3][29] ), .QN(n2528) );
  DFFRX1 \I_cache/cache_reg[4][29]  ( .D(n12587), .CK(clk), .RN(n5831), .Q(
        \I_cache/cache[4][29] ), .QN(n1063) );
  DFFRX1 \I_cache/cache_reg[5][29]  ( .D(n12586), .CK(clk), .RN(n5831), .Q(
        \I_cache/cache[5][29] ), .QN(n2635) );
  DFFRX1 \I_cache/cache_reg[6][29]  ( .D(n12585), .CK(clk), .RN(n5831), .Q(
        \I_cache/cache[6][29] ), .QN(n1057) );
  DFFRX1 \I_cache/cache_reg[7][29]  ( .D(n12584), .CK(clk), .RN(n5831), .Q(
        \I_cache/cache[7][29] ), .QN(n2629) );
  DFFRX1 \I_cache/cache_reg[0][30]  ( .D(n12583), .CK(clk), .RN(n5831), .Q(
        \I_cache/cache[0][30] ), .QN(n1017) );
  DFFRX1 \I_cache/cache_reg[1][30]  ( .D(n12582), .CK(clk), .RN(n5831), .Q(
        \I_cache/cache[1][30] ), .QN(n2589) );
  DFFRX1 \I_cache/cache_reg[2][30]  ( .D(n12581), .CK(clk), .RN(n5831), .Q(
        \I_cache/cache[2][30] ), .QN(n1018) );
  DFFRX1 \I_cache/cache_reg[3][30]  ( .D(n12580), .CK(clk), .RN(n5831), .Q(
        \I_cache/cache[3][30] ), .QN(n2590) );
  DFFRX1 \I_cache/cache_reg[4][30]  ( .D(n12579), .CK(clk), .RN(n5831), .Q(
        \I_cache/cache[4][30] ), .QN(n1049) );
  DFFRX1 \I_cache/cache_reg[5][30]  ( .D(n12578), .CK(clk), .RN(n5831), .Q(
        \I_cache/cache[5][30] ), .QN(n2621) );
  DFFRX1 \I_cache/cache_reg[6][30]  ( .D(n12577), .CK(clk), .RN(n5831), .Q(
        \I_cache/cache[6][30] ), .QN(n1019) );
  DFFRX1 \I_cache/cache_reg[7][30]  ( .D(n12576), .CK(clk), .RN(n5832), .Q(
        \I_cache/cache[7][30] ), .QN(n2591) );
  DFFRX1 \I_cache/cache_reg[0][31]  ( .D(n12575), .CK(clk), .RN(n5832), .Q(
        \I_cache/cache[0][31] ), .QN(n1009) );
  DFFRX1 \I_cache/cache_reg[1][31]  ( .D(n12574), .CK(clk), .RN(n5832), .Q(
        \I_cache/cache[1][31] ), .QN(n2581) );
  DFFRX1 \I_cache/cache_reg[2][31]  ( .D(n12573), .CK(clk), .RN(n5832), .Q(
        \I_cache/cache[2][31] ), .QN(n1010) );
  DFFRX1 \I_cache/cache_reg[3][31]  ( .D(n12572), .CK(clk), .RN(n5832), .Q(
        \I_cache/cache[3][31] ), .QN(n2582) );
  DFFRX1 \I_cache/cache_reg[4][31]  ( .D(n12571), .CK(clk), .RN(n5832), .Q(
        \I_cache/cache[4][31] ), .QN(n1047) );
  DFFRX1 \I_cache/cache_reg[6][31]  ( .D(n12569), .CK(clk), .RN(n5832), .Q(
        \I_cache/cache[6][31] ), .QN(n1011) );
  DFFRX1 \I_cache/cache_reg[0][48]  ( .D(n12439), .CK(clk), .RN(n5843), .Q(
        \I_cache/cache[0][48] ), .QN(n1707) );
  DFFRX1 \I_cache/cache_reg[1][48]  ( .D(n12438), .CK(clk), .RN(n5843), .Q(
        \I_cache/cache[1][48] ), .QN(n3391) );
  DFFRX1 \I_cache/cache_reg[2][48]  ( .D(n12437), .CK(clk), .RN(n5843), .Q(
        \I_cache/cache[2][48] ), .QN(n1708) );
  DFFRX1 \I_cache/cache_reg[4][48]  ( .D(n12435), .CK(clk), .RN(n5843), .Q(
        \I_cache/cache[4][48] ), .QN(n1733) );
  DFFRX1 \I_cache/cache_reg[5][48]  ( .D(n12434), .CK(clk), .RN(n5843), .Q(
        \I_cache/cache[5][48] ), .QN(n3417) );
  DFFRX1 \I_cache/cache_reg[6][48]  ( .D(n12433), .CK(clk), .RN(n5843), .Q(
        \I_cache/cache[6][48] ), .QN(n1709) );
  DFFRX1 \I_cache/cache_reg[0][49]  ( .D(n12431), .CK(clk), .RN(n5844), .Q(
        \I_cache/cache[0][49] ), .QN(n1755) );
  DFFRX1 \I_cache/cache_reg[1][49]  ( .D(n12430), .CK(clk), .RN(n5844), .Q(
        \I_cache/cache[1][49] ), .QN(n3439) );
  DFFRX1 \I_cache/cache_reg[2][49]  ( .D(n12429), .CK(clk), .RN(n5844), .Q(
        \I_cache/cache[2][49] ), .QN(n1756) );
  DFFRX1 \I_cache/cache_reg[3][49]  ( .D(n12428), .CK(clk), .RN(n5844), .Q(
        \I_cache/cache[3][49] ), .QN(n3440) );
  DFFRX1 \I_cache/cache_reg[4][49]  ( .D(n12427), .CK(clk), .RN(n5844), .Q(
        \I_cache/cache[4][49] ), .QN(n1799) );
  DFFRX1 \I_cache/cache_reg[5][49]  ( .D(n12426), .CK(clk), .RN(n5844), .Q(
        \I_cache/cache[5][49] ), .QN(n3483) );
  DFFRX1 \I_cache/cache_reg[6][49]  ( .D(n12425), .CK(clk), .RN(n5844), .Q(
        \I_cache/cache[6][49] ), .QN(n1757) );
  DFFRX1 \I_cache/cache_reg[7][49]  ( .D(n12424), .CK(clk), .RN(n5844), .Q(
        \I_cache/cache[7][49] ), .QN(n3441) );
  DFFRX1 \I_cache/cache_reg[0][50]  ( .D(n12423), .CK(clk), .RN(n5844), .Q(
        \I_cache/cache[0][50] ), .QN(n1698) );
  DFFRX1 \I_cache/cache_reg[1][50]  ( .D(n12422), .CK(clk), .RN(n5844), .Q(
        \I_cache/cache[1][50] ), .QN(n3382) );
  DFFRX1 \I_cache/cache_reg[2][50]  ( .D(n12421), .CK(clk), .RN(n5844), .Q(
        \I_cache/cache[2][50] ), .QN(n1699) );
  DFFRX1 \I_cache/cache_reg[4][50]  ( .D(n12419), .CK(clk), .RN(n5845), .Q(
        \I_cache/cache[4][50] ), .QN(n1730) );
  DFFRX1 \I_cache/cache_reg[5][50]  ( .D(n12418), .CK(clk), .RN(n5845), .Q(
        \I_cache/cache[5][50] ), .QN(n3414) );
  DFFRX1 \I_cache/cache_reg[6][50]  ( .D(n12417), .CK(clk), .RN(n5845), .Q(
        \I_cache/cache[6][50] ), .QN(n1700) );
  DFFRX1 \I_cache/cache_reg[0][51]  ( .D(n12415), .CK(clk), .RN(n5845), .Q(
        \I_cache/cache[0][51] ), .QN(n1746) );
  DFFRX1 \I_cache/cache_reg[1][51]  ( .D(n12414), .CK(clk), .RN(n5845), .Q(
        \I_cache/cache[1][51] ), .QN(n3430) );
  DFFRX1 \I_cache/cache_reg[2][51]  ( .D(n12413), .CK(clk), .RN(n5845), .Q(
        \I_cache/cache[2][51] ), .QN(n1747) );
  DFFRX1 \I_cache/cache_reg[3][51]  ( .D(n12412), .CK(clk), .RN(n5845), .Q(
        \I_cache/cache[3][51] ), .QN(n3431) );
  DFFRX1 \I_cache/cache_reg[4][51]  ( .D(n12411), .CK(clk), .RN(n5845), .Q(
        \I_cache/cache[4][51] ), .QN(n1793) );
  DFFRX1 \I_cache/cache_reg[5][51]  ( .D(n12410), .CK(clk), .RN(n5845), .Q(
        \I_cache/cache[5][51] ), .QN(n3477) );
  DFFRX1 \I_cache/cache_reg[6][51]  ( .D(n12409), .CK(clk), .RN(n5845), .Q(
        \I_cache/cache[6][51] ), .QN(n1748) );
  DFFRX1 \I_cache/cache_reg[7][51]  ( .D(n12408), .CK(clk), .RN(n5846), .Q(
        \I_cache/cache[7][51] ), .QN(n3432) );
  DFFRX1 \I_cache/cache_reg[0][52]  ( .D(n12407), .CK(clk), .RN(n5846), .Q(
        \I_cache/cache[0][52] ), .QN(n1683) );
  DFFRX1 \I_cache/cache_reg[1][52]  ( .D(n12406), .CK(clk), .RN(n5846), .Q(
        \I_cache/cache[1][52] ), .QN(n3367) );
  DFFRX1 \I_cache/cache_reg[2][52]  ( .D(n12405), .CK(clk), .RN(n5846), .Q(
        \I_cache/cache[2][52] ), .QN(n1684) );
  DFFRX1 \I_cache/cache_reg[3][52]  ( .D(n12404), .CK(clk), .RN(n5846), .Q(
        \I_cache/cache[3][52] ), .QN(n3368) );
  DFFRX1 \I_cache/cache_reg[4][52]  ( .D(n12403), .CK(clk), .RN(n5846), .Q(
        \I_cache/cache[4][52] ), .QN(n1725) );
  DFFRX1 \I_cache/cache_reg[5][52]  ( .D(n12402), .CK(clk), .RN(n5846), .Q(
        \I_cache/cache[5][52] ), .QN(n3409) );
  DFFRX1 \I_cache/cache_reg[6][52]  ( .D(n12401), .CK(clk), .RN(n5846), .Q(
        \I_cache/cache[6][52] ), .QN(n1685) );
  DFFRX1 \I_cache/cache_reg[7][52]  ( .D(n12400), .CK(clk), .RN(n5846), .Q(
        \I_cache/cache[7][52] ), .QN(n3369) );
  DFFRX1 \I_cache/cache_reg[0][53]  ( .D(n12399), .CK(clk), .RN(n5846), .Q(
        \I_cache/cache[0][53] ), .QN(n1671) );
  DFFRX1 \I_cache/cache_reg[1][53]  ( .D(n12398), .CK(clk), .RN(n5846), .Q(
        \I_cache/cache[1][53] ), .QN(n3355) );
  DFFRX1 \I_cache/cache_reg[2][53]  ( .D(n12397), .CK(clk), .RN(n5846), .Q(
        \I_cache/cache[2][53] ), .QN(n1672) );
  DFFRX1 \I_cache/cache_reg[3][53]  ( .D(n12396), .CK(clk), .RN(n5847), .Q(
        \I_cache/cache[3][53] ), .QN(n3356) );
  DFFRX1 \I_cache/cache_reg[4][53]  ( .D(n12395), .CK(clk), .RN(n5847), .Q(
        \I_cache/cache[4][53] ), .QN(n1721) );
  DFFRX1 \I_cache/cache_reg[5][53]  ( .D(n12394), .CK(clk), .RN(n5847), .Q(
        \I_cache/cache[5][53] ), .QN(n3405) );
  DFFRX1 \I_cache/cache_reg[6][53]  ( .D(n12393), .CK(clk), .RN(n5847), .Q(
        \I_cache/cache[6][53] ), .QN(n1673) );
  DFFRX1 \I_cache/cache_reg[7][53]  ( .D(n12392), .CK(clk), .RN(n5847), .Q(
        \I_cache/cache[7][53] ), .QN(n3357) );
  DFFRX1 \I_cache/cache_reg[0][54]  ( .D(n12391), .CK(clk), .RN(n5847), .Q(
        \I_cache/cache[0][54] ), .QN(n1743) );
  DFFRX1 \I_cache/cache_reg[1][54]  ( .D(n12390), .CK(clk), .RN(n5847), .Q(
        \I_cache/cache[1][54] ), .QN(n3427) );
  DFFRX1 \I_cache/cache_reg[2][54]  ( .D(n12389), .CK(clk), .RN(n5847), .Q(
        \I_cache/cache[2][54] ), .QN(n1744) );
  DFFRX1 \I_cache/cache_reg[3][54]  ( .D(n12388), .CK(clk), .RN(n5847), .Q(
        \I_cache/cache[3][54] ), .QN(n3428) );
  DFFRX1 \I_cache/cache_reg[4][54]  ( .D(n12387), .CK(clk), .RN(n5847), .Q(
        \I_cache/cache[4][54] ), .QN(n1790) );
  DFFRX1 \I_cache/cache_reg[5][54]  ( .D(n12386), .CK(clk), .RN(n5847), .Q(
        \I_cache/cache[5][54] ), .QN(n3474) );
  DFFRX1 \I_cache/cache_reg[6][54]  ( .D(n12385), .CK(clk), .RN(n5847), .Q(
        \I_cache/cache[6][54] ), .QN(n1745) );
  DFFRX1 \I_cache/cache_reg[7][54]  ( .D(n12384), .CK(clk), .RN(n5848), .Q(
        \I_cache/cache[7][54] ), .QN(n3429) );
  DFFRX1 \I_cache/cache_reg[0][55]  ( .D(n12383), .CK(clk), .RN(n5848), .Q(
        \I_cache/cache[0][55] ), .QN(n1653) );
  DFFRX1 \I_cache/cache_reg[1][55]  ( .D(n12382), .CK(clk), .RN(n5848), .Q(
        \I_cache/cache[1][55] ), .QN(n3337) );
  DFFRX1 \I_cache/cache_reg[2][55]  ( .D(n12381), .CK(clk), .RN(n5848), .Q(
        \I_cache/cache[2][55] ), .QN(n1654) );
  DFFRX1 \I_cache/cache_reg[3][55]  ( .D(n12380), .CK(clk), .RN(n5848), .Q(
        \I_cache/cache[3][55] ), .QN(n3338) );
  DFFRX1 \I_cache/cache_reg[4][55]  ( .D(n12379), .CK(clk), .RN(n5848), .Q(
        \I_cache/cache[4][55] ), .QN(n1715) );
  DFFRX1 \I_cache/cache_reg[5][55]  ( .D(n12378), .CK(clk), .RN(n5848), .Q(
        \I_cache/cache[5][55] ), .QN(n3399) );
  DFFRX1 \I_cache/cache_reg[6][55]  ( .D(n12377), .CK(clk), .RN(n5848), .Q(
        \I_cache/cache[6][55] ), .QN(n1655) );
  DFFRX1 \I_cache/cache_reg[7][55]  ( .D(n12376), .CK(clk), .RN(n5848), .Q(
        \I_cache/cache[7][55] ), .QN(n3339) );
  DFFRX1 \I_cache/cache_reg[0][56]  ( .D(n12375), .CK(clk), .RN(n5848), .Q(
        \I_cache/cache[0][56] ), .QN(n1647) );
  DFFRX1 \I_cache/cache_reg[1][56]  ( .D(n12374), .CK(clk), .RN(n5848), .Q(
        \I_cache/cache[1][56] ), .QN(n3331) );
  DFFRX1 \I_cache/cache_reg[2][56]  ( .D(n12373), .CK(clk), .RN(n5848), .Q(
        \I_cache/cache[2][56] ), .QN(n1648) );
  DFFRX1 \I_cache/cache_reg[3][56]  ( .D(n12372), .CK(clk), .RN(n5849), .Q(
        \I_cache/cache[3][56] ), .QN(n3332) );
  DFFRX1 \I_cache/cache_reg[4][56]  ( .D(n12371), .CK(clk), .RN(n5849), .Q(
        \I_cache/cache[4][56] ), .QN(n1713) );
  DFFRX1 \I_cache/cache_reg[5][56]  ( .D(n12370), .CK(clk), .RN(n5849), .Q(
        \I_cache/cache[5][56] ), .QN(n3397) );
  DFFRX1 \I_cache/cache_reg[6][56]  ( .D(n12369), .CK(clk), .RN(n5849), .Q(
        \I_cache/cache[6][56] ), .QN(n1649) );
  DFFRX1 \I_cache/cache_reg[7][56]  ( .D(n12368), .CK(clk), .RN(n5849), .Q(
        \I_cache/cache[7][56] ), .QN(n3333) );
  DFFRX1 \I_cache/cache_reg[0][57]  ( .D(n12367), .CK(clk), .RN(n5849), .Q(
        \I_cache/cache[0][57] ), .QN(n1737) );
  DFFRX1 \I_cache/cache_reg[1][57]  ( .D(n12366), .CK(clk), .RN(n5849), .Q(
        \I_cache/cache[1][57] ), .QN(n3421) );
  DFFRX1 \I_cache/cache_reg[2][57]  ( .D(n12365), .CK(clk), .RN(n5849), .Q(
        \I_cache/cache[2][57] ), .QN(n1738) );
  DFFRX1 \I_cache/cache_reg[3][57]  ( .D(n12364), .CK(clk), .RN(n5849), .Q(
        \I_cache/cache[3][57] ), .QN(n3422) );
  DFFRX1 \I_cache/cache_reg[4][57]  ( .D(n12363), .CK(clk), .RN(n5849), .Q(
        \I_cache/cache[4][57] ), .QN(n1788) );
  DFFRX1 \I_cache/cache_reg[5][57]  ( .D(n12362), .CK(clk), .RN(n5849), .Q(
        \I_cache/cache[5][57] ), .QN(n3472) );
  DFFRX1 \I_cache/cache_reg[6][57]  ( .D(n12361), .CK(clk), .RN(n5849), .Q(
        \I_cache/cache[6][57] ), .QN(n1739) );
  DFFRX1 \I_cache/cache_reg[7][57]  ( .D(n12360), .CK(clk), .RN(n5850), .Q(
        \I_cache/cache[7][57] ), .QN(n3423) );
  DFFRX1 \I_cache/cache_reg[0][58]  ( .D(n12359), .CK(clk), .RN(n5850), .Q(
        \I_cache/cache[0][58] ), .QN(n1015) );
  DFFRX1 \I_cache/cache_reg[1][58]  ( .D(n12358), .CK(clk), .RN(n5850), .Q(
        \I_cache/cache[1][58] ), .QN(n2587) );
  DFFRX1 \I_cache/cache_reg[2][58]  ( .D(n12357), .CK(clk), .RN(n5850), .Q(
        \I_cache/cache[2][58] ), .QN(n1016) );
  DFFRX1 \I_cache/cache_reg[3][58]  ( .D(n12356), .CK(clk), .RN(n5850), .Q(
        \I_cache/cache[3][58] ), .QN(n2588) );
  DFFRX1 \I_cache/cache_reg[4][58]  ( .D(n12355), .CK(clk), .RN(n5850), .Q(
        \I_cache/cache[4][58] ), .QN(n1215) );
  DFFRX1 \I_cache/cache_reg[5][58]  ( .D(n12354), .CK(clk), .RN(n5850), .Q(
        \I_cache/cache[5][58] ), .QN(n2787) );
  DFFRX1 \I_cache/cache_reg[6][58]  ( .D(n12353), .CK(clk), .RN(n5850), .Q(
        \I_cache/cache[6][58] ), .QN(n2515) );
  DFFRX1 \I_cache/cache_reg[7][58]  ( .D(n12352), .CK(clk), .RN(n5850), .Q(
        \I_cache/cache[7][58] ), .QN(n764) );
  DFFRX1 \I_cache/cache_reg[0][59]  ( .D(n12351), .CK(clk), .RN(n5850), .Q(
        \I_cache/cache[0][59] ), .QN(n1162) );
  DFFRX1 \I_cache/cache_reg[1][59]  ( .D(n12350), .CK(clk), .RN(n5850), .Q(
        \I_cache/cache[1][59] ), .QN(n2734) );
  DFFRX1 \I_cache/cache_reg[2][59]  ( .D(n12349), .CK(clk), .RN(n5850), .Q(
        \I_cache/cache[2][59] ), .QN(n1163) );
  DFFRX1 \I_cache/cache_reg[3][59]  ( .D(n12348), .CK(clk), .RN(n5851), .Q(
        \I_cache/cache[3][59] ), .QN(n2735) );
  DFFRX1 \I_cache/cache_reg[4][59]  ( .D(n12347), .CK(clk), .RN(n5851), .Q(
        \I_cache/cache[4][59] ), .QN(n1219) );
  DFFRX1 \I_cache/cache_reg[5][59]  ( .D(n12346), .CK(clk), .RN(n5851), .Q(
        \I_cache/cache[5][59] ), .QN(n2791) );
  DFFRX1 \I_cache/cache_reg[6][59]  ( .D(n12345), .CK(clk), .RN(n5851), .Q(
        \I_cache/cache[6][59] ), .QN(n1164) );
  DFFRX1 \I_cache/cache_reg[7][59]  ( .D(n12344), .CK(clk), .RN(n5851), .Q(
        \I_cache/cache[7][59] ), .QN(n2736) );
  DFFRX1 \I_cache/cache_reg[0][60]  ( .D(n12343), .CK(clk), .RN(n5851), .Q(
        \I_cache/cache[0][60] ), .QN(n2561) );
  DFFRX1 \I_cache/cache_reg[1][60]  ( .D(n12342), .CK(clk), .RN(n5851), .Q(
        \I_cache/cache[1][60] ), .QN(n790) );
  DFFRX1 \I_cache/cache_reg[2][60]  ( .D(n12341), .CK(clk), .RN(n5851), .Q(
        \I_cache/cache[2][60] ), .QN(n2562) );
  DFFRX1 \I_cache/cache_reg[3][60]  ( .D(n12340), .CK(clk), .RN(n5851), .Q(
        \I_cache/cache[3][60] ), .QN(n791) );
  DFFRX1 \I_cache/cache_reg[4][60]  ( .D(n12339), .CK(clk), .RN(n5851), .Q(
        \I_cache/cache[4][60] ), .QN(n1214) );
  DFFRX1 \I_cache/cache_reg[5][60]  ( .D(n12338), .CK(clk), .RN(n5851), .Q(
        \I_cache/cache[5][60] ), .QN(n2786) );
  DFFRX1 \I_cache/cache_reg[6][60]  ( .D(n12337), .CK(clk), .RN(n5851), .Q(
        \I_cache/cache[6][60] ), .QN(n2563) );
  DFFRX1 \I_cache/cache_reg[7][60]  ( .D(n12336), .CK(clk), .RN(n5852), .Q(
        \I_cache/cache[7][60] ), .QN(n792) );
  DFFRX1 \I_cache/cache_reg[0][61]  ( .D(n12335), .CK(clk), .RN(n5852), .Q(
        \I_cache/cache[0][61] ), .QN(n1156) );
  DFFRX1 \I_cache/cache_reg[1][61]  ( .D(n12334), .CK(clk), .RN(n5852), .Q(
        \I_cache/cache[1][61] ), .QN(n2728) );
  DFFRX1 \I_cache/cache_reg[2][61]  ( .D(n12333), .CK(clk), .RN(n5852), .Q(
        \I_cache/cache[2][61] ), .QN(n1157) );
  DFFRX1 \I_cache/cache_reg[3][61]  ( .D(n12332), .CK(clk), .RN(n5852), .Q(
        \I_cache/cache[3][61] ), .QN(n2729) );
  DFFRX1 \I_cache/cache_reg[4][61]  ( .D(n12331), .CK(clk), .RN(n5852), .Q(
        \I_cache/cache[4][61] ), .QN(n1207) );
  DFFRX1 \I_cache/cache_reg[5][61]  ( .D(n12330), .CK(clk), .RN(n5852), .Q(
        \I_cache/cache[5][61] ), .QN(n2779) );
  DFFRX1 \I_cache/cache_reg[6][61]  ( .D(n12329), .CK(clk), .RN(n5852), .Q(
        \I_cache/cache[6][61] ), .QN(n1158) );
  DFFRX1 \I_cache/cache_reg[7][61]  ( .D(n12328), .CK(clk), .RN(n5852), .Q(
        \I_cache/cache[7][61] ), .QN(n2730) );
  DFFRX1 \I_cache/cache_reg[0][62]  ( .D(n12327), .CK(clk), .RN(n5852), .Q(
        \I_cache/cache[0][62] ), .QN(n1180) );
  DFFRX1 \I_cache/cache_reg[1][62]  ( .D(n12326), .CK(clk), .RN(n5852), .Q(
        \I_cache/cache[1][62] ), .QN(n2752) );
  DFFRX1 \I_cache/cache_reg[2][62]  ( .D(n12325), .CK(clk), .RN(n5852), .Q(
        \I_cache/cache[2][62] ), .QN(n1181) );
  DFFRX1 \I_cache/cache_reg[3][62]  ( .D(n12324), .CK(clk), .RN(n5853), .Q(
        \I_cache/cache[3][62] ), .QN(n2753) );
  DFFRX1 \I_cache/cache_reg[4][62]  ( .D(n12323), .CK(clk), .RN(n5853), .Q(
        \I_cache/cache[4][62] ), .QN(n1212) );
  DFFRX1 \I_cache/cache_reg[5][62]  ( .D(n12322), .CK(clk), .RN(n5853), .Q(
        \I_cache/cache[5][62] ), .QN(n2784) );
  DFFRX1 \I_cache/cache_reg[6][62]  ( .D(n12321), .CK(clk), .RN(n5853), .Q(
        \I_cache/cache[6][62] ), .QN(n1182) );
  DFFRX1 \I_cache/cache_reg[7][62]  ( .D(n12320), .CK(clk), .RN(n5853), .Q(
        \I_cache/cache[7][62] ), .QN(n2754) );
  DFFRX1 \I_cache/cache_reg[0][63]  ( .D(n12319), .CK(clk), .RN(n5853), .Q(
        \I_cache/cache[0][63] ), .QN(n1183) );
  DFFRX1 \I_cache/cache_reg[1][63]  ( .D(n12318), .CK(clk), .RN(n5853), .Q(
        \I_cache/cache[1][63] ), .QN(n2755) );
  DFFRX1 \I_cache/cache_reg[2][63]  ( .D(n12317), .CK(clk), .RN(n5853), .Q(
        \I_cache/cache[2][63] ), .QN(n1184) );
  DFFRX1 \I_cache/cache_reg[3][63]  ( .D(n12316), .CK(clk), .RN(n5853), .Q(
        \I_cache/cache[3][63] ), .QN(n2756) );
  DFFRX1 \I_cache/cache_reg[4][63]  ( .D(n12315), .CK(clk), .RN(n5853), .Q(
        \I_cache/cache[4][63] ), .QN(n1209) );
  DFFRX1 \I_cache/cache_reg[5][63]  ( .D(n12314), .CK(clk), .RN(n5853), .Q(
        \I_cache/cache[5][63] ), .QN(n2781) );
  DFFRX1 \I_cache/cache_reg[6][63]  ( .D(n12313), .CK(clk), .RN(n5853), .Q(
        \I_cache/cache[6][63] ), .QN(n1185) );
  DFFRX1 \I_cache/cache_reg[7][63]  ( .D(n12312), .CK(clk), .RN(n5854), .Q(
        \I_cache/cache[7][63] ), .QN(n2757) );
  DFFRX1 \I_cache/cache_reg[0][64]  ( .D(n12311), .CK(clk), .RN(n5854), .Q(
        \I_cache/cache[0][64] ), .QN(n1761) );
  DFFRX1 \I_cache/cache_reg[1][64]  ( .D(n12310), .CK(clk), .RN(n5854), .Q(
        \I_cache/cache[1][64] ), .QN(n3445) );
  DFFRX1 \I_cache/cache_reg[2][64]  ( .D(n12309), .CK(clk), .RN(n5854), .Q(
        \I_cache/cache[2][64] ), .QN(n1762) );
  DFFRX1 \I_cache/cache_reg[3][64]  ( .D(n12308), .CK(clk), .RN(n5854), .Q(
        \I_cache/cache[3][64] ), .QN(n3446) );
  DFFRX1 \I_cache/cache_reg[6][64]  ( .D(n12305), .CK(clk), .RN(n5854), .Q(
        \I_cache/cache[6][64] ), .QN(n1763) );
  DFFRX1 \I_cache/cache_reg[7][64]  ( .D(n12304), .CK(clk), .RN(n5854), .Q(
        \I_cache/cache[7][64] ), .QN(n3447) );
  DFFRX1 \I_cache/cache_reg[0][80]  ( .D(n12183), .CK(clk), .RN(n5864), .Q(
        \I_cache/cache[0][80] ), .QN(n1758) );
  DFFRX1 \I_cache/cache_reg[1][80]  ( .D(n12182), .CK(clk), .RN(n5864), .Q(
        \I_cache/cache[1][80] ), .QN(n3442) );
  DFFRX1 \I_cache/cache_reg[2][80]  ( .D(n12181), .CK(clk), .RN(n5864), .Q(
        \I_cache/cache[2][80] ), .QN(n1759) );
  DFFRX1 \I_cache/cache_reg[4][80]  ( .D(n12179), .CK(clk), .RN(n5865), .Q(
        \I_cache/cache[4][80] ), .QN(n1794) );
  DFFRX1 \I_cache/cache_reg[5][80]  ( .D(n12178), .CK(clk), .RN(n5865), .Q(
        \I_cache/cache[5][80] ), .QN(n3478) );
  DFFRX1 \I_cache/cache_reg[6][80]  ( .D(n12177), .CK(clk), .RN(n5865), .Q(
        \I_cache/cache[6][80] ), .QN(n1760) );
  DFFRX1 \I_cache/cache_reg[0][81]  ( .D(n12175), .CK(clk), .RN(n5865), .Q(
        \I_cache/cache[0][81] ), .QN(n1752) );
  DFFRX1 \I_cache/cache_reg[1][81]  ( .D(n12174), .CK(clk), .RN(n5865), .Q(
        \I_cache/cache[1][81] ), .QN(n3436) );
  DFFRX1 \I_cache/cache_reg[2][81]  ( .D(n12173), .CK(clk), .RN(n5865), .Q(
        \I_cache/cache[2][81] ), .QN(n1753) );
  DFFRX1 \I_cache/cache_reg[3][81]  ( .D(n12172), .CK(clk), .RN(n5865), .Q(
        \I_cache/cache[3][81] ), .QN(n3437) );
  DFFRX1 \I_cache/cache_reg[4][81]  ( .D(n12171), .CK(clk), .RN(n5865), .Q(
        \I_cache/cache[4][81] ), .QN(n1798) );
  DFFRX1 \I_cache/cache_reg[5][81]  ( .D(n12170), .CK(clk), .RN(n5865), .Q(
        \I_cache/cache[5][81] ), .QN(n3482) );
  DFFRX1 \I_cache/cache_reg[6][81]  ( .D(n12169), .CK(clk), .RN(n5865), .Q(
        \I_cache/cache[6][81] ), .QN(n1754) );
  DFFRX1 \I_cache/cache_reg[7][81]  ( .D(n12168), .CK(clk), .RN(n5866), .Q(
        \I_cache/cache[7][81] ), .QN(n3438) );
  DFFRX1 \I_cache/cache_reg[0][82]  ( .D(n12167), .CK(clk), .RN(n5866), .Q(
        \I_cache/cache[0][82] ), .QN(n1695) );
  DFFRX1 \I_cache/cache_reg[2][82]  ( .D(n12165), .CK(clk), .RN(n5866), .Q(
        \I_cache/cache[2][82] ), .QN(n1696) );
  DFFRX1 \I_cache/cache_reg[3][82]  ( .D(n12164), .CK(clk), .RN(n5866), .Q(
        \I_cache/cache[3][82] ), .QN(n3380) );
  DFFRX1 \I_cache/cache_reg[4][82]  ( .D(n12163), .CK(clk), .RN(n5866), .Q(
        \I_cache/cache[4][82] ), .QN(n1729) );
  DFFRX1 \I_cache/cache_reg[5][82]  ( .D(n12162), .CK(clk), .RN(n5866), .Q(
        \I_cache/cache[5][82] ), .QN(n3413) );
  DFFRX1 \I_cache/cache_reg[6][82]  ( .D(n12161), .CK(clk), .RN(n5866), .Q(
        \I_cache/cache[6][82] ), .QN(n1697) );
  DFFRX1 \I_cache/cache_reg[0][83]  ( .D(n12159), .CK(clk), .RN(n5866), .Q(
        \I_cache/cache[0][83] ), .QN(n1686) );
  DFFRX1 \I_cache/cache_reg[1][83]  ( .D(n12158), .CK(clk), .RN(n5866), .Q(
        \I_cache/cache[1][83] ), .QN(n3370) );
  DFFRX1 \I_cache/cache_reg[2][83]  ( .D(n12157), .CK(clk), .RN(n5866), .Q(
        \I_cache/cache[2][83] ), .QN(n1687) );
  DFFRX1 \I_cache/cache_reg[3][83]  ( .D(n12156), .CK(clk), .RN(n5867), .Q(
        \I_cache/cache[3][83] ), .QN(n3371) );
  DFFRX1 \I_cache/cache_reg[4][83]  ( .D(n12155), .CK(clk), .RN(n5867), .Q(
        \I_cache/cache[4][83] ), .QN(n1726) );
  DFFRX1 \I_cache/cache_reg[5][83]  ( .D(n12154), .CK(clk), .RN(n5867), .Q(
        \I_cache/cache[5][83] ), .QN(n3410) );
  DFFRX1 \I_cache/cache_reg[6][83]  ( .D(n12153), .CK(clk), .RN(n5867), .Q(
        \I_cache/cache[6][83] ), .QN(n1688) );
  DFFRX1 \I_cache/cache_reg[7][83]  ( .D(n12152), .CK(clk), .RN(n5867), .Q(
        \I_cache/cache[7][83] ), .QN(n3372) );
  DFFRX1 \I_cache/cache_reg[0][84]  ( .D(n12151), .CK(clk), .RN(n5867), .Q(
        \I_cache/cache[0][84] ), .QN(n1680) );
  DFFRX1 \I_cache/cache_reg[1][84]  ( .D(n12150), .CK(clk), .RN(n5867), .Q(
        \I_cache/cache[1][84] ), .QN(n3364) );
  DFFRX1 \I_cache/cache_reg[2][84]  ( .D(n12149), .CK(clk), .RN(n5867), .Q(
        \I_cache/cache[2][84] ), .QN(n1681) );
  DFFRX1 \I_cache/cache_reg[3][84]  ( .D(n12148), .CK(clk), .RN(n5867), .Q(
        \I_cache/cache[3][84] ), .QN(n3365) );
  DFFRX1 \I_cache/cache_reg[4][84]  ( .D(n12147), .CK(clk), .RN(n5867), .Q(
        \I_cache/cache[4][84] ), .QN(n1724) );
  DFFRX1 \I_cache/cache_reg[5][84]  ( .D(n12146), .CK(clk), .RN(n5867), .Q(
        \I_cache/cache[5][84] ), .QN(n3408) );
  DFFRX1 \I_cache/cache_reg[6][84]  ( .D(n12145), .CK(clk), .RN(n5867), .Q(
        \I_cache/cache[6][84] ), .QN(n1682) );
  DFFRX1 \I_cache/cache_reg[7][84]  ( .D(n12144), .CK(clk), .RN(n5868), .Q(
        \I_cache/cache[7][84] ), .QN(n3366) );
  DFFRX1 \I_cache/cache_reg[0][85]  ( .D(n12143), .CK(clk), .RN(n5868), .Q(
        \I_cache/cache[0][85] ), .QN(n1668) );
  DFFRX1 \I_cache/cache_reg[1][85]  ( .D(n12142), .CK(clk), .RN(n5868), .Q(
        \I_cache/cache[1][85] ), .QN(n3352) );
  DFFRX1 \I_cache/cache_reg[2][85]  ( .D(n12141), .CK(clk), .RN(n5868), .Q(
        \I_cache/cache[2][85] ), .QN(n1669) );
  DFFRX1 \I_cache/cache_reg[3][85]  ( .D(n12140), .CK(clk), .RN(n5868), .Q(
        \I_cache/cache[3][85] ), .QN(n3353) );
  DFFRX1 \I_cache/cache_reg[4][85]  ( .D(n12139), .CK(clk), .RN(n5868), .Q(
        \I_cache/cache[4][85] ), .QN(n1720) );
  DFFRX1 \I_cache/cache_reg[5][85]  ( .D(n12138), .CK(clk), .RN(n5868), .Q(
        \I_cache/cache[5][85] ), .QN(n3404) );
  DFFRX1 \I_cache/cache_reg[6][85]  ( .D(n12137), .CK(clk), .RN(n5868), .Q(
        \I_cache/cache[6][85] ), .QN(n1670) );
  DFFRX1 \I_cache/cache_reg[7][85]  ( .D(n12136), .CK(clk), .RN(n5868), .Q(
        \I_cache/cache[7][85] ), .QN(n3354) );
  DFFRX1 \I_cache/cache_reg[0][86]  ( .D(n12135), .CK(clk), .RN(n5868), .Q(
        \I_cache/cache[0][86] ), .QN(n1659) );
  DFFRX1 \I_cache/cache_reg[1][86]  ( .D(n12134), .CK(clk), .RN(n5868), .Q(
        \I_cache/cache[1][86] ), .QN(n3343) );
  DFFRX1 \I_cache/cache_reg[2][86]  ( .D(n12133), .CK(clk), .RN(n5868), .Q(
        \I_cache/cache[2][86] ), .QN(n1660) );
  DFFRX1 \I_cache/cache_reg[3][86]  ( .D(n12132), .CK(clk), .RN(n5869), .Q(
        \I_cache/cache[3][86] ), .QN(n3344) );
  DFFRX1 \I_cache/cache_reg[4][86]  ( .D(n12131), .CK(clk), .RN(n5869), .Q(
        \I_cache/cache[4][86] ), .QN(n1717) );
  DFFRX1 \I_cache/cache_reg[5][86]  ( .D(n12130), .CK(clk), .RN(n5869), .Q(
        \I_cache/cache[5][86] ), .QN(n3401) );
  DFFRX1 \I_cache/cache_reg[6][86]  ( .D(n12129), .CK(clk), .RN(n5869), .Q(
        \I_cache/cache[6][86] ), .QN(n1661) );
  DFFRX1 \I_cache/cache_reg[7][86]  ( .D(n12128), .CK(clk), .RN(n5869), .Q(
        \I_cache/cache[7][86] ), .QN(n3345) );
  DFFRX1 \I_cache/cache_reg[0][87]  ( .D(n12127), .CK(clk), .RN(n5869), .Q(
        \I_cache/cache[0][87] ), .QN(n1740) );
  DFFRX1 \I_cache/cache_reg[1][87]  ( .D(n12126), .CK(clk), .RN(n5869), .Q(
        \I_cache/cache[1][87] ), .QN(n3424) );
  DFFRX1 \I_cache/cache_reg[2][87]  ( .D(n12125), .CK(clk), .RN(n5869), .Q(
        \I_cache/cache[2][87] ), .QN(n1741) );
  DFFRX1 \I_cache/cache_reg[3][87]  ( .D(n12124), .CK(clk), .RN(n5869), .Q(
        \I_cache/cache[3][87] ), .QN(n3425) );
  DFFRX1 \I_cache/cache_reg[4][87]  ( .D(n12123), .CK(clk), .RN(n5869), .Q(
        \I_cache/cache[4][87] ), .QN(n1801) );
  DFFRX1 \I_cache/cache_reg[5][87]  ( .D(n12122), .CK(clk), .RN(n5869), .Q(
        \I_cache/cache[5][87] ), .QN(n3485) );
  DFFRX1 \I_cache/cache_reg[6][87]  ( .D(n12121), .CK(clk), .RN(n5869), .Q(
        \I_cache/cache[6][87] ), .QN(n1742) );
  DFFRX1 \I_cache/cache_reg[7][87]  ( .D(n12120), .CK(clk), .RN(n5870), .Q(
        \I_cache/cache[7][87] ), .QN(n3426) );
  DFFRX1 \I_cache/cache_reg[0][88]  ( .D(n12119), .CK(clk), .RN(n5870), .Q(
        \I_cache/cache[0][88] ), .QN(n1644) );
  DFFRX1 \I_cache/cache_reg[1][88]  ( .D(n12118), .CK(clk), .RN(n5870), .Q(
        \I_cache/cache[1][88] ), .QN(n3328) );
  DFFRX1 \I_cache/cache_reg[2][88]  ( .D(n12117), .CK(clk), .RN(n5870), .Q(
        \I_cache/cache[2][88] ), .QN(n1645) );
  DFFRX1 \I_cache/cache_reg[3][88]  ( .D(n12116), .CK(clk), .RN(n5870), .Q(
        \I_cache/cache[3][88] ), .QN(n3329) );
  DFFRX1 \I_cache/cache_reg[4][88]  ( .D(n12115), .CK(clk), .RN(n5870), .Q(
        \I_cache/cache[4][88] ), .QN(n1712) );
  DFFRX1 \I_cache/cache_reg[5][88]  ( .D(n12114), .CK(clk), .RN(n5870), .Q(
        \I_cache/cache[5][88] ), .QN(n3396) );
  DFFRX1 \I_cache/cache_reg[6][88]  ( .D(n12113), .CK(clk), .RN(n5870), .Q(
        \I_cache/cache[6][88] ), .QN(n1646) );
  DFFRX1 \I_cache/cache_reg[7][88]  ( .D(n12112), .CK(clk), .RN(n5870), .Q(
        \I_cache/cache[7][88] ), .QN(n3330) );
  DFFRX1 \I_cache/cache_reg[0][89]  ( .D(n12111), .CK(clk), .RN(n5870), .Q(
        \I_cache/cache[0][89] ), .QN(n1734) );
  DFFRX1 \I_cache/cache_reg[1][89]  ( .D(n12110), .CK(clk), .RN(n5870), .Q(
        \I_cache/cache[1][89] ), .QN(n3418) );
  DFFRX1 \I_cache/cache_reg[2][89]  ( .D(n12109), .CK(clk), .RN(n5870), .Q(
        \I_cache/cache[2][89] ), .QN(n1735) );
  DFFRX1 \I_cache/cache_reg[3][89]  ( .D(n12108), .CK(clk), .RN(n5871), .Q(
        \I_cache/cache[3][89] ), .QN(n3419) );
  DFFRX1 \I_cache/cache_reg[4][89]  ( .D(n12107), .CK(clk), .RN(n5871), .Q(
        \I_cache/cache[4][89] ), .QN(n1787) );
  DFFRX1 \I_cache/cache_reg[5][89]  ( .D(n12106), .CK(clk), .RN(n5871), .Q(
        \I_cache/cache[5][89] ), .QN(n3471) );
  DFFRX1 \I_cache/cache_reg[6][89]  ( .D(n12105), .CK(clk), .RN(n5871), .Q(
        \I_cache/cache[6][89] ), .QN(n1736) );
  DFFRX1 \I_cache/cache_reg[7][89]  ( .D(n12104), .CK(clk), .RN(n5871), .Q(
        \I_cache/cache[7][89] ), .QN(n3420) );
  DFFRX1 \I_cache/cache_reg[0][90]  ( .D(n12103), .CK(clk), .RN(n5871), .Q(
        \I_cache/cache[0][90] ), .QN(n1014) );
  DFFRX1 \I_cache/cache_reg[1][90]  ( .D(n12102), .CK(clk), .RN(n5871), .Q(
        \I_cache/cache[1][90] ), .QN(n2586) );
  DFFRX1 \I_cache/cache_reg[2][90]  ( .D(n12101), .CK(clk), .RN(n5871), .Q(
        \I_cache/cache[2][90] ), .QN(n2513) );
  DFFRX1 \I_cache/cache_reg[3][90]  ( .D(n12100), .CK(clk), .RN(n5871), .Q(
        \I_cache/cache[3][90] ), .QN(n762) );
  DFFRX1 \I_cache/cache_reg[6][90]  ( .D(n12097), .CK(clk), .RN(n5871), .Q(
        \I_cache/cache[6][90] ), .QN(n2514) );
  DFFRX1 \I_cache/cache_reg[7][90]  ( .D(n12096), .CK(clk), .RN(n5872), .Q(
        \I_cache/cache[7][90] ), .QN(n763) );
  DFFRX1 \I_cache/cache_reg[0][91]  ( .D(n12095), .CK(clk), .RN(n5872), .Q(
        \I_cache/cache[0][91] ), .QN(n1159) );
  DFFRX1 \I_cache/cache_reg[1][91]  ( .D(n12094), .CK(clk), .RN(n5872), .Q(
        \I_cache/cache[1][91] ), .QN(n2731) );
  DFFRX1 \I_cache/cache_reg[2][91]  ( .D(n12093), .CK(clk), .RN(n5872), .Q(
        \I_cache/cache[2][91] ), .QN(n1160) );
  DFFRX1 \I_cache/cache_reg[3][91]  ( .D(n12092), .CK(clk), .RN(n5872), .Q(
        \I_cache/cache[3][91] ), .QN(n2732) );
  DFFRX1 \I_cache/cache_reg[4][91]  ( .D(n12091), .CK(clk), .RN(n5872), .Q(
        \I_cache/cache[4][91] ), .QN(n1217) );
  DFFRX1 \I_cache/cache_reg[5][91]  ( .D(n12090), .CK(clk), .RN(n5872), .Q(
        \I_cache/cache[5][91] ), .QN(n2789) );
  DFFRX1 \I_cache/cache_reg[6][91]  ( .D(n12089), .CK(clk), .RN(n5872), .Q(
        \I_cache/cache[6][91] ), .QN(n1161) );
  DFFRX1 \I_cache/cache_reg[7][91]  ( .D(n12088), .CK(clk), .RN(n5872), .Q(
        \I_cache/cache[7][91] ), .QN(n2733) );
  DFFRX1 \I_cache/cache_reg[0][92]  ( .D(n12087), .CK(clk), .RN(n5872), .Q(
        \I_cache/cache[0][92] ), .QN(n2558) );
  DFFRX1 \I_cache/cache_reg[1][92]  ( .D(n12086), .CK(clk), .RN(n5872), .Q(
        \I_cache/cache[1][92] ), .QN(n787) );
  DFFRX1 \I_cache/cache_reg[2][92]  ( .D(n12085), .CK(clk), .RN(n5872), .Q(
        \I_cache/cache[2][92] ), .QN(n2559) );
  DFFRX1 \I_cache/cache_reg[3][92]  ( .D(n12084), .CK(clk), .RN(n5873), .Q(
        \I_cache/cache[3][92] ), .QN(n788) );
  DFFRX1 \I_cache/cache_reg[4][92]  ( .D(n12083), .CK(clk), .RN(n5873), .Q(
        \I_cache/cache[4][92] ), .QN(n1213) );
  DFFRX1 \I_cache/cache_reg[5][92]  ( .D(n12082), .CK(clk), .RN(n5873), .Q(
        \I_cache/cache[5][92] ), .QN(n2785) );
  DFFRX1 \I_cache/cache_reg[6][92]  ( .D(n12081), .CK(clk), .RN(n5873), .Q(
        \I_cache/cache[6][92] ), .QN(n2560) );
  DFFRX1 \I_cache/cache_reg[7][92]  ( .D(n12080), .CK(clk), .RN(n5873), .Q(
        \I_cache/cache[7][92] ), .QN(n789) );
  DFFRX1 \I_cache/cache_reg[0][93]  ( .D(n12079), .CK(clk), .RN(n5873), .Q(
        \I_cache/cache[0][93] ), .QN(n1006) );
  DFFRX1 \I_cache/cache_reg[1][93]  ( .D(n12078), .CK(clk), .RN(n5873), .Q(
        \I_cache/cache[1][93] ), .QN(n2578) );
  DFFRX1 \I_cache/cache_reg[2][93]  ( .D(n12077), .CK(clk), .RN(n5873), .Q(
        \I_cache/cache[2][93] ), .QN(n1007) );
  DFFRX1 \I_cache/cache_reg[3][93]  ( .D(n12076), .CK(clk), .RN(n5873), .Q(
        \I_cache/cache[3][93] ), .QN(n2579) );
  DFFRX1 \I_cache/cache_reg[4][93]  ( .D(n12075), .CK(clk), .RN(n5873), .Q(
        \I_cache/cache[4][93] ), .QN(n1046) );
  DFFRX1 \I_cache/cache_reg[5][93]  ( .D(n12074), .CK(clk), .RN(n5873), .Q(
        \I_cache/cache[5][93] ), .QN(n2618) );
  DFFRX1 \I_cache/cache_reg[6][93]  ( .D(n12073), .CK(clk), .RN(n5873), .Q(
        \I_cache/cache[6][93] ), .QN(n1008) );
  DFFRX1 \I_cache/cache_reg[7][93]  ( .D(n12072), .CK(clk), .RN(n5874), .Q(
        \I_cache/cache[7][93] ), .QN(n2580) );
  DFFRX1 \I_cache/cache_reg[0][94]  ( .D(n12071), .CK(clk), .RN(n5874), .Q(
        \I_cache/cache[0][94] ), .QN(n1171) );
  DFFRX1 \I_cache/cache_reg[1][94]  ( .D(n12070), .CK(clk), .RN(n5874), .Q(
        \I_cache/cache[1][94] ), .QN(n2743) );
  DFFRX1 \I_cache/cache_reg[2][94]  ( .D(n12069), .CK(clk), .RN(n5874), .Q(
        \I_cache/cache[2][94] ), .QN(n1172) );
  DFFRX1 \I_cache/cache_reg[3][94]  ( .D(n12068), .CK(clk), .RN(n5874), .Q(
        \I_cache/cache[3][94] ), .QN(n2744) );
  DFFRX1 \I_cache/cache_reg[4][94]  ( .D(n12067), .CK(clk), .RN(n5874), .Q(
        \I_cache/cache[4][94] ), .QN(n1208) );
  DFFRX1 \I_cache/cache_reg[5][94]  ( .D(n12066), .CK(clk), .RN(n5874), .Q(
        \I_cache/cache[5][94] ), .QN(n2780) );
  DFFRX1 \I_cache/cache_reg[6][94]  ( .D(n12065), .CK(clk), .RN(n5874), .Q(
        \I_cache/cache[6][94] ), .QN(n1173) );
  DFFRX1 \I_cache/cache_reg[7][94]  ( .D(n12064), .CK(clk), .RN(n5874), .Q(
        \I_cache/cache[7][94] ), .QN(n2745) );
  DFFRX1 \I_cache/cache_reg[0][95]  ( .D(n12063), .CK(clk), .RN(n5874), .Q(
        \I_cache/cache[0][95] ), .QN(n1174) );
  DFFRX1 \I_cache/cache_reg[1][95]  ( .D(n12062), .CK(clk), .RN(n5874), .Q(
        \I_cache/cache[1][95] ), .QN(n2746) );
  DFFRX1 \I_cache/cache_reg[2][95]  ( .D(n12061), .CK(clk), .RN(n5874), .Q(
        \I_cache/cache[2][95] ), .QN(n1175) );
  DFFRX1 \I_cache/cache_reg[3][95]  ( .D(n12060), .CK(clk), .RN(n5875), .Q(
        \I_cache/cache[3][95] ), .QN(n2747) );
  DFFRX1 \I_cache/cache_reg[4][95]  ( .D(n12059), .CK(clk), .RN(n5875), .Q(
        \I_cache/cache[4][95] ), .QN(n1206) );
  DFFRX1 \I_cache/cache_reg[5][95]  ( .D(n12058), .CK(clk), .RN(n5875), .Q(
        \I_cache/cache[5][95] ), .QN(n2778) );
  DFFRX1 \I_cache/cache_reg[6][95]  ( .D(n12057), .CK(clk), .RN(n5875), .Q(
        \I_cache/cache[6][95] ), .QN(n1176) );
  DFFRX1 \I_cache/cache_reg[7][95]  ( .D(n12056), .CK(clk), .RN(n5875), .Q(
        \I_cache/cache[7][95] ), .QN(n2748) );
  DFFRX1 \I_cache/cache_reg[0][112]  ( .D(n11927), .CK(clk), .RN(n5886), .Q(
        \I_cache/cache[0][112] ), .QN(n1704) );
  DFFRX1 \I_cache/cache_reg[2][112]  ( .D(n11925), .CK(clk), .RN(n5886), .Q(
        \I_cache/cache[2][112] ), .QN(n1705) );
  DFFRX1 \I_cache/cache_reg[3][112]  ( .D(n11924), .CK(clk), .RN(n5886), .Q(
        \I_cache/cache[3][112] ), .QN(n3389) );
  DFFRX1 \I_cache/cache_reg[4][112]  ( .D(n11923), .CK(clk), .RN(n5886), .Q(
        \I_cache/cache[4][112] ), .QN(n1732) );
  DFFRX1 \I_cache/cache_reg[5][112]  ( .D(n11922), .CK(clk), .RN(n5886), .Q(
        \I_cache/cache[5][112] ), .QN(n3416) );
  DFFRX1 \I_cache/cache_reg[6][112]  ( .D(n11921), .CK(clk), .RN(n5886), .Q(
        \I_cache/cache[6][112] ), .QN(n1706) );
  DFFRX1 \I_cache/cache_reg[0][113]  ( .D(n11919), .CK(clk), .RN(n5886), .Q(
        \I_cache/cache[0][113] ), .QN(n1749) );
  DFFRX1 \I_cache/cache_reg[1][113]  ( .D(n11918), .CK(clk), .RN(n5886), .Q(
        \I_cache/cache[1][113] ), .QN(n3433) );
  DFFRX1 \I_cache/cache_reg[2][113]  ( .D(n11917), .CK(clk), .RN(n5886), .Q(
        \I_cache/cache[2][113] ), .QN(n1750) );
  DFFRX1 \I_cache/cache_reg[3][113]  ( .D(n11916), .CK(clk), .RN(n5887), .Q(
        \I_cache/cache[3][113] ), .QN(n3434) );
  DFFRX1 \I_cache/cache_reg[4][113]  ( .D(n11915), .CK(clk), .RN(n5887), .Q(
        \I_cache/cache[4][113] ), .QN(n1797) );
  DFFRX1 \I_cache/cache_reg[5][113]  ( .D(n11914), .CK(clk), .RN(n5887), .Q(
        \I_cache/cache[5][113] ), .QN(n3481) );
  DFFRX1 \I_cache/cache_reg[6][113]  ( .D(n11913), .CK(clk), .RN(n5887), .Q(
        \I_cache/cache[6][113] ), .QN(n1751) );
  DFFRX1 \I_cache/cache_reg[7][113]  ( .D(n11912), .CK(clk), .RN(n5887), .Q(
        \I_cache/cache[7][113] ), .QN(n3435) );
  DFFRX1 \I_cache/cache_reg[0][114]  ( .D(n11911), .CK(clk), .RN(n5887), .Q(
        \I_cache/cache[0][114] ), .QN(n1692) );
  DFFRX1 \I_cache/cache_reg[1][114]  ( .D(n11910), .CK(clk), .RN(n5887), .Q(
        \I_cache/cache[1][114] ), .QN(n3376) );
  DFFRX1 \I_cache/cache_reg[2][114]  ( .D(n11909), .CK(clk), .RN(n5887), .Q(
        \I_cache/cache[2][114] ), .QN(n1693) );
  DFFRX1 \I_cache/cache_reg[5][114]  ( .D(n11906), .CK(clk), .RN(n5887), .Q(
        \I_cache/cache[5][114] ), .QN(n3412) );
  DFFRX1 \I_cache/cache_reg[6][114]  ( .D(n11905), .CK(clk), .RN(n5887), .Q(
        \I_cache/cache[6][114] ), .QN(n1694) );
  DFFRX1 \I_cache/cache_reg[7][114]  ( .D(n11904), .CK(clk), .RN(n5888), .Q(
        \I_cache/cache[7][114] ), .QN(n3378) );
  DFFRX1 \I_cache/cache_reg[0][115]  ( .D(n11903), .CK(clk), .RN(n5888), .Q(
        \I_cache/cache[0][115] ), .QN(n1779) );
  DFFRX1 \I_cache/cache_reg[1][115]  ( .D(n11902), .CK(clk), .RN(n5888), .Q(
        \I_cache/cache[1][115] ), .QN(n3463) );
  DFFRX1 \I_cache/cache_reg[2][115]  ( .D(n11901), .CK(clk), .RN(n5888), .Q(
        \I_cache/cache[2][115] ), .QN(n1780) );
  DFFRX1 \I_cache/cache_reg[3][115]  ( .D(n11900), .CK(clk), .RN(n5888), .Q(
        \I_cache/cache[3][115] ), .QN(n3464) );
  DFFRX1 \I_cache/cache_reg[4][115]  ( .D(n11899), .CK(clk), .RN(n5888), .Q(
        \I_cache/cache[4][115] ), .QN(n1792) );
  DFFRX1 \I_cache/cache_reg[5][115]  ( .D(n11898), .CK(clk), .RN(n5888), .Q(
        \I_cache/cache[5][115] ), .QN(n3476) );
  DFFRX1 \I_cache/cache_reg[6][115]  ( .D(n11897), .CK(clk), .RN(n5888), .Q(
        \I_cache/cache[6][115] ), .QN(n1781) );
  DFFRX1 \I_cache/cache_reg[7][115]  ( .D(n11896), .CK(clk), .RN(n5888), .Q(
        \I_cache/cache[7][115] ), .QN(n3465) );
  DFFRX1 \I_cache/cache_reg[0][116]  ( .D(n11895), .CK(clk), .RN(n5888), .Q(
        \I_cache/cache[0][116] ), .QN(n1677) );
  DFFRX1 \I_cache/cache_reg[1][116]  ( .D(n11894), .CK(clk), .RN(n5888), .Q(
        \I_cache/cache[1][116] ), .QN(n3361) );
  DFFRX1 \I_cache/cache_reg[2][116]  ( .D(n11893), .CK(clk), .RN(n5888), .Q(
        \I_cache/cache[2][116] ), .QN(n1678) );
  DFFRX1 \I_cache/cache_reg[3][116]  ( .D(n11892), .CK(clk), .RN(n5889), .Q(
        \I_cache/cache[3][116] ), .QN(n3362) );
  DFFRX1 \I_cache/cache_reg[4][116]  ( .D(n11891), .CK(clk), .RN(n5889), .Q(
        \I_cache/cache[4][116] ), .QN(n1723) );
  DFFRX1 \I_cache/cache_reg[5][116]  ( .D(n11890), .CK(clk), .RN(n5889), .Q(
        \I_cache/cache[5][116] ), .QN(n3407) );
  DFFRX1 \I_cache/cache_reg[6][116]  ( .D(n11889), .CK(clk), .RN(n5889), .Q(
        \I_cache/cache[6][116] ), .QN(n1679) );
  DFFRX1 \I_cache/cache_reg[7][116]  ( .D(n11888), .CK(clk), .RN(n5889), .Q(
        \I_cache/cache[7][116] ), .QN(n3363) );
  DFFRX1 \I_cache/cache_reg[0][117]  ( .D(n11887), .CK(clk), .RN(n5889), .Q(
        \I_cache/cache[0][117] ), .QN(n1665) );
  DFFRX1 \I_cache/cache_reg[1][117]  ( .D(n11886), .CK(clk), .RN(n5889), .Q(
        \I_cache/cache[1][117] ), .QN(n3349) );
  DFFRX1 \I_cache/cache_reg[2][117]  ( .D(n11885), .CK(clk), .RN(n5889), .Q(
        \I_cache/cache[2][117] ), .QN(n1666) );
  DFFRX1 \I_cache/cache_reg[3][117]  ( .D(n11884), .CK(clk), .RN(n5889), .Q(
        \I_cache/cache[3][117] ), .QN(n3350) );
  DFFRX1 \I_cache/cache_reg[4][117]  ( .D(n11883), .CK(clk), .RN(n5889), .Q(
        \I_cache/cache[4][117] ), .QN(n1719) );
  DFFRX1 \I_cache/cache_reg[5][117]  ( .D(n11882), .CK(clk), .RN(n5889), .Q(
        \I_cache/cache[5][117] ), .QN(n3403) );
  DFFRX1 \I_cache/cache_reg[6][117]  ( .D(n11881), .CK(clk), .RN(n5889), .Q(
        \I_cache/cache[6][117] ), .QN(n1667) );
  DFFRX1 \I_cache/cache_reg[7][117]  ( .D(n11880), .CK(clk), .RN(n5890), .Q(
        \I_cache/cache[7][117] ), .QN(n3351) );
  DFFRX1 \I_cache/cache_reg[0][118]  ( .D(n11879), .CK(clk), .RN(n5890), .Q(
        \I_cache/cache[0][118] ), .QN(n1656) );
  DFFRX1 \I_cache/cache_reg[1][118]  ( .D(n11878), .CK(clk), .RN(n5890), .Q(
        \I_cache/cache[1][118] ), .QN(n3340) );
  DFFRX1 \I_cache/cache_reg[2][118]  ( .D(n11877), .CK(clk), .RN(n5890), .Q(
        \I_cache/cache[2][118] ), .QN(n1657) );
  DFFRX1 \I_cache/cache_reg[3][118]  ( .D(n11876), .CK(clk), .RN(n5890), .Q(
        \I_cache/cache[3][118] ), .QN(n3341) );
  DFFRX1 \I_cache/cache_reg[4][118]  ( .D(n11875), .CK(clk), .RN(n5890), .Q(
        \I_cache/cache[4][118] ), .QN(n1716) );
  DFFRX1 \I_cache/cache_reg[5][118]  ( .D(n11874), .CK(clk), .RN(n5890), .Q(
        \I_cache/cache[5][118] ), .QN(n3400) );
  DFFRX1 \I_cache/cache_reg[6][118]  ( .D(n11873), .CK(clk), .RN(n5890), .Q(
        \I_cache/cache[6][118] ), .QN(n1658) );
  DFFRX1 \I_cache/cache_reg[7][118]  ( .D(n11872), .CK(clk), .RN(n5890), .Q(
        \I_cache/cache[7][118] ), .QN(n3342) );
  DFFRX1 \I_cache/cache_reg[0][119]  ( .D(n11871), .CK(clk), .RN(n5890), .Q(
        \I_cache/cache[0][119] ), .QN(n1770) );
  DFFRX1 \I_cache/cache_reg[1][119]  ( .D(n11870), .CK(clk), .RN(n5890), .Q(
        \I_cache/cache[1][119] ), .QN(n3454) );
  DFFRX1 \I_cache/cache_reg[2][119]  ( .D(n11869), .CK(clk), .RN(n5890), .Q(
        \I_cache/cache[2][119] ), .QN(n1771) );
  DFFRX1 \I_cache/cache_reg[3][119]  ( .D(n11868), .CK(clk), .RN(n5891), .Q(
        \I_cache/cache[3][119] ), .QN(n3455) );
  DFFRX1 \I_cache/cache_reg[4][119]  ( .D(n11867), .CK(clk), .RN(n5891), .Q(
        \I_cache/cache[4][119] ), .QN(n1800) );
  DFFRX1 \I_cache/cache_reg[5][119]  ( .D(n11866), .CK(clk), .RN(n5891), .Q(
        \I_cache/cache[5][119] ), .QN(n3484) );
  DFFRX1 \I_cache/cache_reg[6][119]  ( .D(n11865), .CK(clk), .RN(n5891), .Q(
        \I_cache/cache[6][119] ), .QN(n1772) );
  DFFRX1 \I_cache/cache_reg[7][119]  ( .D(n11864), .CK(clk), .RN(n5891), .Q(
        \I_cache/cache[7][119] ), .QN(n3456) );
  DFFRX1 \I_cache/cache_reg[0][120]  ( .D(n11863), .CK(clk), .RN(n5891), .Q(
        \I_cache/cache[0][120] ), .QN(n1641) );
  DFFRX1 \I_cache/cache_reg[1][120]  ( .D(n11862), .CK(clk), .RN(n5891), .Q(
        \I_cache/cache[1][120] ), .QN(n3325) );
  DFFRX1 \I_cache/cache_reg[2][120]  ( .D(n11861), .CK(clk), .RN(n5891), .Q(
        \I_cache/cache[2][120] ), .QN(n1642) );
  DFFRX1 \I_cache/cache_reg[3][120]  ( .D(n11860), .CK(clk), .RN(n5891), .Q(
        \I_cache/cache[3][120] ), .QN(n3326) );
  DFFRX1 \I_cache/cache_reg[4][120]  ( .D(n11859), .CK(clk), .RN(n5891), .Q(
        \I_cache/cache[4][120] ), .QN(n1711) );
  DFFRX1 \I_cache/cache_reg[5][120]  ( .D(n11858), .CK(clk), .RN(n5891), .Q(
        \I_cache/cache[5][120] ), .QN(n3395) );
  DFFRX1 \I_cache/cache_reg[6][120]  ( .D(n11857), .CK(clk), .RN(n5891), .Q(
        \I_cache/cache[6][120] ), .QN(n1643) );
  DFFRX1 \I_cache/cache_reg[7][120]  ( .D(n11856), .CK(clk), .RN(n5892), .Q(
        \I_cache/cache[7][120] ), .QN(n3327) );
  DFFRX1 \I_cache/cache_reg[0][121]  ( .D(n11855), .CK(clk), .RN(n5892), .Q(
        \I_cache/cache[0][121] ), .QN(n1767) );
  DFFRX1 \I_cache/cache_reg[1][121]  ( .D(n11854), .CK(clk), .RN(n5892), .Q(
        \I_cache/cache[1][121] ), .QN(n3451) );
  DFFRX1 \I_cache/cache_reg[2][121]  ( .D(n11853), .CK(clk), .RN(n5892), .Q(
        \I_cache/cache[2][121] ), .QN(n1768) );
  DFFRX1 \I_cache/cache_reg[3][121]  ( .D(n11852), .CK(clk), .RN(n5892), .Q(
        \I_cache/cache[3][121] ), .QN(n3452) );
  DFFRX1 \I_cache/cache_reg[4][121]  ( .D(n11851), .CK(clk), .RN(n5892), .Q(
        \I_cache/cache[4][121] ), .QN(n1786) );
  DFFRX1 \I_cache/cache_reg[6][121]  ( .D(n11849), .CK(clk), .RN(n5892), .Q(
        \I_cache/cache[6][121] ), .QN(n1769) );
  DFFRX1 \I_cache/cache_reg[0][122]  ( .D(n11847), .CK(clk), .RN(n5892), .Q(
        \I_cache/cache[0][122] ), .QN(n1012) );
  DFFRX1 \I_cache/cache_reg[1][122]  ( .D(n11846), .CK(clk), .RN(n5892), .Q(
        \I_cache/cache[1][122] ), .QN(n2584) );
  DFFRX1 \I_cache/cache_reg[2][122]  ( .D(n11845), .CK(clk), .RN(n5892), .Q(
        \I_cache/cache[2][122] ), .QN(n1013) );
  DFFRX1 \I_cache/cache_reg[3][122]  ( .D(n11844), .CK(clk), .RN(n5893), .Q(
        \I_cache/cache[3][122] ), .QN(n2585) );
  DFFRX1 \I_cache/cache_reg[4][122]  ( .D(n11843), .CK(clk), .RN(n5893), .Q(
        \I_cache/cache[4][122] ), .QN(n2527) );
  DFFRX1 \I_cache/cache_reg[5][122]  ( .D(n11842), .CK(clk), .RN(n5893), .Q(
        \I_cache/cache[5][122] ), .QN(n775) );
  DFFRX1 \I_cache/cache_reg[6][122]  ( .D(n11841), .CK(clk), .RN(n5893), .Q(
        \I_cache/cache[6][122] ), .QN(n2512) );
  DFFRX1 \I_cache/cache_reg[7][122]  ( .D(n11840), .CK(clk), .RN(n5893), .Q(
        \I_cache/cache[7][122] ), .QN(n761) );
  DFFRX1 \I_cache/cache_reg[0][123]  ( .D(n11839), .CK(clk), .RN(n5893), .Q(
        \I_cache/cache[0][123] ), .QN(n1165) );
  DFFRX1 \I_cache/cache_reg[1][123]  ( .D(n11838), .CK(clk), .RN(n5893), .Q(
        \I_cache/cache[1][123] ), .QN(n2737) );
  DFFRX1 \I_cache/cache_reg[2][123]  ( .D(n11837), .CK(clk), .RN(n5893), .Q(
        \I_cache/cache[2][123] ), .QN(n1166) );
  DFFRX1 \I_cache/cache_reg[3][123]  ( .D(n11836), .CK(clk), .RN(n5893), .Q(
        \I_cache/cache[3][123] ), .QN(n2738) );
  DFFRX1 \I_cache/cache_reg[4][123]  ( .D(n11835), .CK(clk), .RN(n5893), .Q(
        \I_cache/cache[4][123] ), .QN(n1218) );
  DFFRX1 \I_cache/cache_reg[5][123]  ( .D(n11834), .CK(clk), .RN(n5893), .Q(
        \I_cache/cache[5][123] ), .QN(n2790) );
  DFFRX1 \I_cache/cache_reg[6][123]  ( .D(n11833), .CK(clk), .RN(n5893), .Q(
        \I_cache/cache[6][123] ), .QN(n1167) );
  DFFRX1 \I_cache/cache_reg[7][123]  ( .D(n11832), .CK(clk), .RN(n5894), .Q(
        \I_cache/cache[7][123] ), .QN(n2739) );
  DFFRX1 \I_cache/cache_reg[0][124]  ( .D(n11831), .CK(clk), .RN(n5894), .Q(
        \I_cache/cache[0][124] ), .QN(n1186) );
  DFFRX1 \I_cache/cache_reg[1][124]  ( .D(n11830), .CK(clk), .RN(n5894), .Q(
        \I_cache/cache[1][124] ), .QN(n2758) );
  DFFRX1 \I_cache/cache_reg[2][124]  ( .D(n11829), .CK(clk), .RN(n5894), .Q(
        \I_cache/cache[2][124] ), .QN(n1187) );
  DFFRX1 \I_cache/cache_reg[3][124]  ( .D(n11828), .CK(clk), .RN(n5894), .Q(
        \I_cache/cache[3][124] ), .QN(n2759) );
  DFFRX1 \I_cache/cache_reg[4][124]  ( .D(n11827), .CK(clk), .RN(n5894), .Q(
        \I_cache/cache[4][124] ), .QN(n2508) );
  DFFRX1 \I_cache/cache_reg[5][124]  ( .D(n11826), .CK(clk), .RN(n5894), .Q(
        \I_cache/cache[5][124] ), .QN(n748) );
  DFFRX1 \I_cache/cache_reg[6][124]  ( .D(n11825), .CK(clk), .RN(n5894), .Q(
        \I_cache/cache[6][124] ), .QN(n2564) );
  DFFRX1 \I_cache/cache_reg[7][124]  ( .D(n11824), .CK(clk), .RN(n5894), .Q(
        \I_cache/cache[7][124] ), .QN(n793) );
  DFFRX1 \I_cache/cache_reg[0][125]  ( .D(n11823), .CK(clk), .RN(n5894), .Q(
        \I_cache/cache[0][125] ), .QN(n1003) );
  DFFRX1 \I_cache/cache_reg[1][125]  ( .D(n11822), .CK(clk), .RN(n5894), .Q(
        \I_cache/cache[1][125] ), .QN(n2575) );
  DFFRX1 \I_cache/cache_reg[2][125]  ( .D(n11821), .CK(clk), .RN(n5894), .Q(
        \I_cache/cache[2][125] ), .QN(n1004) );
  DFFRX1 \I_cache/cache_reg[3][125]  ( .D(n11820), .CK(clk), .RN(n5895), .Q(
        \I_cache/cache[3][125] ), .QN(n2576) );
  DFFRX1 \I_cache/cache_reg[4][125]  ( .D(n11819), .CK(clk), .RN(n5895), .Q(
        \I_cache/cache[4][125] ), .QN(n1045) );
  DFFRX1 \I_cache/cache_reg[5][125]  ( .D(n11818), .CK(clk), .RN(n5895), .Q(
        \I_cache/cache[5][125] ), .QN(n2617) );
  DFFRX1 \I_cache/cache_reg[6][125]  ( .D(n11817), .CK(clk), .RN(n5895), .Q(
        \I_cache/cache[6][125] ), .QN(n1005) );
  DFFRX1 \I_cache/cache_reg[7][125]  ( .D(n11816), .CK(clk), .RN(n5895), .Q(
        \I_cache/cache[7][125] ), .QN(n2577) );
  DFFRX1 \I_cache/cache_reg[0][126]  ( .D(n11815), .CK(clk), .RN(n5895), .Q(
        \I_cache/cache[0][126] ), .QN(n1177) );
  DFFRX1 \I_cache/cache_reg[1][126]  ( .D(n11814), .CK(clk), .RN(n5895), .Q(
        \I_cache/cache[1][126] ), .QN(n2749) );
  DFFRX1 \I_cache/cache_reg[2][126]  ( .D(n11813), .CK(clk), .RN(n5895), .Q(
        \I_cache/cache[2][126] ), .QN(n987) );
  DFFRX1 \I_cache/cache_reg[3][126]  ( .D(n11812), .CK(clk), .RN(n5895), .Q(
        \I_cache/cache[3][126] ), .QN(n2539) );
  DFFRX1 \I_cache/cache_reg[4][126]  ( .D(n11811), .CK(clk), .RN(n5895), .Q(
        \I_cache/cache[4][126] ), .QN(n1062) );
  DFFRX1 \I_cache/cache_reg[5][126]  ( .D(n11810), .CK(clk), .RN(n5895), .Q(
        \I_cache/cache[5][126] ), .QN(n2634) );
  DFFRX1 \I_cache/cache_reg[6][126]  ( .D(n11809), .CK(clk), .RN(n5895), .Q(
        \I_cache/cache[6][126] ), .QN(n1178) );
  DFFRX1 \I_cache/cache_reg[7][126]  ( .D(n11808), .CK(clk), .RN(n5896), .Q(
        \I_cache/cache[7][126] ), .QN(n2750) );
  DFFRX1 \I_cache/cache_reg[0][127]  ( .D(n11807), .CK(clk), .RN(n5896), .Q(
        \I_cache/cache[0][127] ), .QN(n1179) );
  DFFRX1 \I_cache/cache_reg[1][127]  ( .D(n11806), .CK(clk), .RN(n5896), .Q(
        \I_cache/cache[1][127] ), .QN(n2751) );
  DFFRX1 \I_cache/cache_reg[2][127]  ( .D(n11805), .CK(clk), .RN(n5896), .Q(
        \I_cache/cache[2][127] ), .QN(n989) );
  DFFRX1 \I_cache/cache_reg[3][127]  ( .D(n11804), .CK(clk), .RN(n5896), .Q(
        \I_cache/cache[3][127] ), .QN(n2541) );
  DFFRX1 \I_cache/cache_reg[4][127]  ( .D(n11803), .CK(clk), .RN(n5896), .Q(
        \I_cache/cache[4][127] ), .QN(n998) );
  DFFRX1 \I_cache/cache_reg[5][127]  ( .D(n11802), .CK(clk), .RN(n5896), .Q(
        \I_cache/cache[5][127] ), .QN(n2550) );
  DFFRX1 \I_cache/cache_reg[6][127]  ( .D(n11801), .CK(clk), .RN(n5896), .Q(
        \I_cache/cache[6][127] ), .QN(n988) );
  DFFRX1 \I_cache/cache_reg[7][127]  ( .D(n11800), .CK(clk), .RN(n5896), .Q(
        \I_cache/cache[7][127] ), .QN(n2540) );
  DFFRX1 \i_MIPS/Register/register_reg[30][0]  ( .D(\i_MIPS/Register/n148 ), 
        .CK(clk), .RN(n5625), .Q(\i_MIPS/Register/register[30][0] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][1]  ( .D(\i_MIPS/Register/n149 ), 
        .CK(clk), .RN(n5625), .Q(\i_MIPS/Register/register[30][1] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][4]  ( .D(\i_MIPS/Register/n152 ), 
        .CK(clk), .RN(n5625), .Q(\i_MIPS/Register/register[30][4] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][5]  ( .D(\i_MIPS/Register/n153 ), 
        .CK(clk), .RN(n5625), .Q(\i_MIPS/Register/register[30][5] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][8]  ( .D(\i_MIPS/Register/n156 ), 
        .CK(clk), .RN(n5626), .Q(\i_MIPS/Register/register[30][8] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][10]  ( .D(\i_MIPS/Register/n158 ), 
        .CK(clk), .RN(n5626), .Q(\i_MIPS/Register/register[30][10] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][11]  ( .D(\i_MIPS/Register/n159 ), 
        .CK(clk), .RN(n5626), .Q(\i_MIPS/Register/register[30][11] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][12]  ( .D(\i_MIPS/Register/n160 ), 
        .CK(clk), .RN(n5626), .Q(\i_MIPS/Register/register[30][12] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][15]  ( .D(\i_MIPS/Register/n163 ), 
        .CK(clk), .RN(n5626), .Q(\i_MIPS/Register/register[30][15] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][17]  ( .D(\i_MIPS/Register/n165 ), 
        .CK(clk), .RN(n5626), .Q(\i_MIPS/Register/register[30][17] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][18]  ( .D(\i_MIPS/Register/n166 ), 
        .CK(clk), .RN(n5626), .Q(\i_MIPS/Register/register[30][18] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][19]  ( .D(\i_MIPS/Register/n167 ), 
        .CK(clk), .RN(n5627), .Q(\i_MIPS/Register/register[30][19] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][26]  ( .D(\i_MIPS/Register/n174 ), 
        .CK(clk), .RN(n5627), .Q(\i_MIPS/Register/register[30][26] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][29]  ( .D(\i_MIPS/Register/n177 ), 
        .CK(clk), .RN(n5627), .Q(\i_MIPS/Register/register[30][29] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][30]  ( .D(\i_MIPS/Register/n178 ), 
        .CK(clk), .RN(n5627), .Q(\i_MIPS/Register/register[30][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][31]  ( .D(\i_MIPS/Register/n179 ), 
        .CK(clk), .RN(n5628), .Q(\i_MIPS/Register/register[30][31] ) );
  DFFRX1 \i_MIPS/Register/register_reg[29][0]  ( .D(\i_MIPS/Register/n180 ), 
        .CK(clk), .RN(n5628), .Q(\i_MIPS/Register/register[29][0] ) );
  DFFRX1 \i_MIPS/Register/register_reg[28][1]  ( .D(\i_MIPS/Register/n213 ), 
        .CK(clk), .RN(n5630), .Q(\i_MIPS/Register/register[28][1] ) );
  DFFRX1 \i_MIPS/Register/register_reg[28][19]  ( .D(\i_MIPS/Register/n231 ), 
        .CK(clk), .RN(n5632), .Q(\i_MIPS/Register/register[28][19] ) );
  DFFRX1 \i_MIPS/Register/register_reg[28][30]  ( .D(\i_MIPS/Register/n242 ), 
        .CK(clk), .RN(n5633), .Q(\i_MIPS/Register/register[28][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[27][0]  ( .D(\i_MIPS/Register/n244 ), 
        .CK(clk), .RN(n5633), .Q(\i_MIPS/Register/register[27][0] ) );
  DFFRX1 \i_MIPS/Register/register_reg[25][0]  ( .D(\i_MIPS/Register/n308 ), 
        .CK(clk), .RN(n5638), .Q(\i_MIPS/Register/register[25][0] ) );
  DFFRX1 \i_MIPS/Register/register_reg[24][1]  ( .D(\i_MIPS/Register/n341 ), 
        .CK(clk), .RN(n5641), .Q(\i_MIPS/Register/register[24][1] ) );
  DFFRX1 \i_MIPS/Register/register_reg[24][19]  ( .D(\i_MIPS/Register/n359 ), 
        .CK(clk), .RN(n5643), .Q(\i_MIPS/Register/register[24][19] ) );
  DFFRX1 \i_MIPS/Register/register_reg[24][30]  ( .D(\i_MIPS/Register/n370 ), 
        .CK(clk), .RN(n5643), .Q(\i_MIPS/Register/register[24][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[15][0]  ( .D(\i_MIPS/Register/n628 ), 
        .CK(clk), .RN(n5665), .Q(\i_MIPS/Register/register[15][0] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][0]  ( .D(\i_MIPS/Register/n660 ), 
        .CK(clk), .RN(n5668), .Q(\i_MIPS/Register/register[14][0] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][1]  ( .D(\i_MIPS/Register/n661 ), 
        .CK(clk), .RN(n5668), .Q(\i_MIPS/Register/register[14][1] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][4]  ( .D(\i_MIPS/Register/n664 ), 
        .CK(clk), .RN(n5668), .Q(\i_MIPS/Register/register[14][4] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][5]  ( .D(\i_MIPS/Register/n665 ), 
        .CK(clk), .RN(n5668), .Q(\i_MIPS/Register/register[14][5] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][8]  ( .D(\i_MIPS/Register/n668 ), 
        .CK(clk), .RN(n5668), .Q(\i_MIPS/Register/register[14][8] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][9]  ( .D(\i_MIPS/Register/n669 ), 
        .CK(clk), .RN(n5668), .Q(\i_MIPS/Register/register[14][9] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][10]  ( .D(\i_MIPS/Register/n670 ), 
        .CK(clk), .RN(n5668), .Q(\i_MIPS/Register/register[14][10] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][11]  ( .D(\i_MIPS/Register/n671 ), 
        .CK(clk), .RN(n5669), .Q(\i_MIPS/Register/register[14][11] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][12]  ( .D(\i_MIPS/Register/n672 ), 
        .CK(clk), .RN(n5669), .Q(\i_MIPS/Register/register[14][12] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][15]  ( .D(\i_MIPS/Register/n675 ), 
        .CK(clk), .RN(n5669), .Q(\i_MIPS/Register/register[14][15] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][17]  ( .D(\i_MIPS/Register/n677 ), 
        .CK(clk), .RN(n5669), .Q(\i_MIPS/Register/register[14][17] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][18]  ( .D(\i_MIPS/Register/n678 ), 
        .CK(clk), .RN(n5669), .Q(\i_MIPS/Register/register[14][18] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][19]  ( .D(\i_MIPS/Register/n679 ), 
        .CK(clk), .RN(n5669), .Q(\i_MIPS/Register/register[14][19] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][26]  ( .D(\i_MIPS/Register/n686 ), 
        .CK(clk), .RN(n5670), .Q(\i_MIPS/Register/register[14][26] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][29]  ( .D(\i_MIPS/Register/n689 ), 
        .CK(clk), .RN(n5670), .Q(\i_MIPS/Register/register[14][29] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][30]  ( .D(\i_MIPS/Register/n690 ), 
        .CK(clk), .RN(n5670), .Q(\i_MIPS/Register/register[14][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][31]  ( .D(\i_MIPS/Register/n691 ), 
        .CK(clk), .RN(n5670), .Q(\i_MIPS/Register/register[14][31] ) );
  DFFRX1 \i_MIPS/Register/register_reg[13][0]  ( .D(\i_MIPS/Register/n692 ), 
        .CK(clk), .RN(n5670), .Q(\i_MIPS/Register/register[13][0] ) );
  DFFRX1 \i_MIPS/Register/register_reg[12][1]  ( .D(\i_MIPS/Register/n725 ), 
        .CK(clk), .RN(n5673), .Q(\i_MIPS/Register/register[12][1] ) );
  DFFRX1 \i_MIPS/Register/register_reg[12][19]  ( .D(\i_MIPS/Register/n743 ), 
        .CK(clk), .RN(n5675), .Q(\i_MIPS/Register/register[12][19] ) );
  DFFRX1 \i_MIPS/Register/register_reg[12][30]  ( .D(\i_MIPS/Register/n754 ), 
        .CK(clk), .RN(n5675), .Q(\i_MIPS/Register/register[12][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[11][0]  ( .D(\i_MIPS/Register/n756 ), 
        .CK(clk), .RN(n5676), .Q(\i_MIPS/Register/register[11][0] ) );
  DFFRX1 \i_MIPS/Register/register_reg[9][0]  ( .D(\i_MIPS/Register/n820 ), 
        .CK(clk), .RN(n5681), .Q(\i_MIPS/Register/register[9][0] ) );
  DFFRX1 \i_MIPS/Register/register_reg[8][1]  ( .D(\i_MIPS/Register/n853 ), 
        .CK(clk), .RN(n5684), .Q(\i_MIPS/Register/register[8][1] ) );
  DFFRX1 \i_MIPS/Register/register_reg[8][19]  ( .D(\i_MIPS/Register/n871 ), 
        .CK(clk), .RN(n5685), .Q(\i_MIPS/Register/register[8][19] ) );
  DFFRX1 \i_MIPS/Register/register_reg[8][30]  ( .D(\i_MIPS/Register/n882 ), 
        .CK(clk), .RN(n5686), .Q(\i_MIPS/Register/register[8][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[23][0]  ( .D(\i_MIPS/Register/n372 ), 
        .CK(clk), .RN(n5644), .Q(\i_MIPS/Register/register[23][0] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][0]  ( .D(\i_MIPS/Register/n404 ), 
        .CK(clk), .RN(n5646), .Q(\i_MIPS/Register/register[22][0] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][1]  ( .D(\i_MIPS/Register/n405 ), 
        .CK(clk), .RN(n5646), .Q(\i_MIPS/Register/register[22][1] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][2]  ( .D(\i_MIPS/Register/n406 ), 
        .CK(clk), .RN(n5646), .Q(\i_MIPS/Register/register[22][2] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][4]  ( .D(\i_MIPS/Register/n408 ), 
        .CK(clk), .RN(n5647), .Q(\i_MIPS/Register/register[22][4] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][5]  ( .D(\i_MIPS/Register/n409 ), 
        .CK(clk), .RN(n5647), .Q(\i_MIPS/Register/register[22][5] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][6]  ( .D(\i_MIPS/Register/n410 ), 
        .CK(clk), .RN(n5647), .Q(\i_MIPS/Register/register[22][6] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][7]  ( .D(\i_MIPS/Register/n411 ), 
        .CK(clk), .RN(n5647), .Q(\i_MIPS/Register/register[22][7] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][8]  ( .D(\i_MIPS/Register/n412 ), 
        .CK(clk), .RN(n5647), .Q(\i_MIPS/Register/register[22][8] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][9]  ( .D(\i_MIPS/Register/n413 ), 
        .CK(clk), .RN(n5647), .Q(\i_MIPS/Register/register[22][9] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][10]  ( .D(\i_MIPS/Register/n414 ), 
        .CK(clk), .RN(n5647), .Q(\i_MIPS/Register/register[22][10] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][11]  ( .D(\i_MIPS/Register/n415 ), 
        .CK(clk), .RN(n5647), .Q(\i_MIPS/Register/register[22][11] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][12]  ( .D(\i_MIPS/Register/n416 ), 
        .CK(clk), .RN(n5647), .Q(\i_MIPS/Register/register[22][12] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][13]  ( .D(\i_MIPS/Register/n417 ), 
        .CK(clk), .RN(n5647), .Q(\i_MIPS/Register/register[22][13] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][14]  ( .D(\i_MIPS/Register/n418 ), 
        .CK(clk), .RN(n5647), .Q(\i_MIPS/Register/register[22][14] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][15]  ( .D(\i_MIPS/Register/n419 ), 
        .CK(clk), .RN(n5648), .Q(\i_MIPS/Register/register[22][15] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][17]  ( .D(\i_MIPS/Register/n421 ), 
        .CK(clk), .RN(n5648), .Q(\i_MIPS/Register/register[22][17] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][18]  ( .D(\i_MIPS/Register/n422 ), 
        .CK(clk), .RN(n5648), .Q(\i_MIPS/Register/register[22][18] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][19]  ( .D(\i_MIPS/Register/n423 ), 
        .CK(clk), .RN(n5648), .Q(\i_MIPS/Register/register[22][19] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][21]  ( .D(\i_MIPS/Register/n425 ), 
        .CK(clk), .RN(n5648), .Q(\i_MIPS/Register/register[22][21] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][25]  ( .D(\i_MIPS/Register/n429 ), 
        .CK(clk), .RN(n5648), .Q(\i_MIPS/Register/register[22][25] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][26]  ( .D(\i_MIPS/Register/n430 ), 
        .CK(clk), .RN(n5648), .Q(\i_MIPS/Register/register[22][26] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][27]  ( .D(\i_MIPS/Register/n431 ), 
        .CK(clk), .RN(n5649), .Q(\i_MIPS/Register/register[22][27] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][28]  ( .D(\i_MIPS/Register/n432 ), 
        .CK(clk), .RN(n5649), .Q(\i_MIPS/Register/register[22][28] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][29]  ( .D(\i_MIPS/Register/n433 ), 
        .CK(clk), .RN(n5649), .Q(\i_MIPS/Register/register[22][29] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][30]  ( .D(\i_MIPS/Register/n434 ), 
        .CK(clk), .RN(n5649), .Q(\i_MIPS/Register/register[22][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][31]  ( .D(\i_MIPS/Register/n435 ), 
        .CK(clk), .RN(n5649), .Q(\i_MIPS/Register/register[22][31] ) );
  DFFRX1 \i_MIPS/Register/register_reg[21][0]  ( .D(\i_MIPS/Register/n436 ), 
        .CK(clk), .RN(n5649), .Q(\i_MIPS/Register/register[21][0] ) );
  DFFRX1 \i_MIPS/Register/register_reg[20][1]  ( .D(\i_MIPS/Register/n469 ), 
        .CK(clk), .RN(n5652), .Q(\i_MIPS/Register/register[20][1] ) );
  DFFRX1 \i_MIPS/Register/register_reg[20][19]  ( .D(\i_MIPS/Register/n487 ), 
        .CK(clk), .RN(n5653), .Q(\i_MIPS/Register/register[20][19] ) );
  DFFRX1 \i_MIPS/Register/register_reg[20][30]  ( .D(\i_MIPS/Register/n498 ), 
        .CK(clk), .RN(n5654), .Q(\i_MIPS/Register/register[20][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[19][0]  ( .D(\i_MIPS/Register/n500 ), 
        .CK(clk), .RN(n5654), .Q(\i_MIPS/Register/register[19][0] ) );
  DFFRX1 \i_MIPS/Register/register_reg[17][0]  ( .D(\i_MIPS/Register/n564 ), 
        .CK(clk), .RN(n5660), .Q(\i_MIPS/Register/register[17][0] ) );
  DFFRX1 \i_MIPS/Register/register_reg[16][1]  ( .D(\i_MIPS/Register/n597 ), 
        .CK(clk), .RN(n5662), .Q(\i_MIPS/Register/register[16][1] ) );
  DFFRX1 \i_MIPS/Register/register_reg[16][19]  ( .D(\i_MIPS/Register/n615 ), 
        .CK(clk), .RN(n5664), .Q(\i_MIPS/Register/register[16][19] ) );
  DFFRX1 \i_MIPS/Register/register_reg[16][30]  ( .D(\i_MIPS/Register/n626 ), 
        .CK(clk), .RN(n5665), .Q(\i_MIPS/Register/register[16][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[7][0]  ( .D(\i_MIPS/Register/n884 ), 
        .CK(clk), .RN(n5686), .Q(\i_MIPS/Register/register[7][0] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][0]  ( .D(\i_MIPS/Register/n916 ), 
        .CK(clk), .RN(n5689), .Q(\i_MIPS/Register/register[6][0] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][1]  ( .D(\i_MIPS/Register/n917 ), 
        .CK(clk), .RN(n5689), .Q(\i_MIPS/Register/register[6][1] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][2]  ( .D(\i_MIPS/Register/n918 ), 
        .CK(clk), .RN(n5689), .Q(\i_MIPS/Register/register[6][2] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][4]  ( .D(\i_MIPS/Register/n920 ), 
        .CK(clk), .RN(n5689), .Q(\i_MIPS/Register/register[6][4] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][5]  ( .D(\i_MIPS/Register/n921 ), 
        .CK(clk), .RN(n5689), .Q(\i_MIPS/Register/register[6][5] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][6]  ( .D(\i_MIPS/Register/n922 ), 
        .CK(clk), .RN(n5689), .Q(\i_MIPS/Register/register[6][6] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][7]  ( .D(\i_MIPS/Register/n923 ), 
        .CK(clk), .RN(n5690), .Q(\i_MIPS/Register/register[6][7] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][8]  ( .D(\i_MIPS/Register/n924 ), 
        .CK(clk), .RN(n5690), .Q(\i_MIPS/Register/register[6][8] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][9]  ( .D(\i_MIPS/Register/n925 ), 
        .CK(clk), .RN(n5690), .Q(\i_MIPS/Register/register[6][9] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][10]  ( .D(\i_MIPS/Register/n926 ), 
        .CK(clk), .RN(n5690), .Q(\i_MIPS/Register/register[6][10] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][11]  ( .D(\i_MIPS/Register/n927 ), 
        .CK(clk), .RN(n5690), .Q(\i_MIPS/Register/register[6][11] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][12]  ( .D(\i_MIPS/Register/n928 ), 
        .CK(clk), .RN(n5690), .Q(\i_MIPS/Register/register[6][12] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][13]  ( .D(\i_MIPS/Register/n929 ), 
        .CK(clk), .RN(n5690), .Q(\i_MIPS/Register/register[6][13] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][14]  ( .D(\i_MIPS/Register/n930 ), 
        .CK(clk), .RN(n5690), .Q(\i_MIPS/Register/register[6][14] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][15]  ( .D(\i_MIPS/Register/n931 ), 
        .CK(clk), .RN(n5690), .Q(\i_MIPS/Register/register[6][15] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][17]  ( .D(\i_MIPS/Register/n933 ), 
        .CK(clk), .RN(n5690), .Q(\i_MIPS/Register/register[6][17] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][18]  ( .D(\i_MIPS/Register/n934 ), 
        .CK(clk), .RN(n5690), .Q(\i_MIPS/Register/register[6][18] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][19]  ( .D(\i_MIPS/Register/n935 ), 
        .CK(clk), .RN(n5691), .Q(\i_MIPS/Register/register[6][19] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][21]  ( .D(\i_MIPS/Register/n937 ), 
        .CK(clk), .RN(n5691), .Q(\i_MIPS/Register/register[6][21] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][25]  ( .D(\i_MIPS/Register/n941 ), 
        .CK(clk), .RN(n5691), .Q(\i_MIPS/Register/register[6][25] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][26]  ( .D(\i_MIPS/Register/n942 ), 
        .CK(clk), .RN(n5691), .Q(\i_MIPS/Register/register[6][26] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][27]  ( .D(\i_MIPS/Register/n943 ), 
        .CK(clk), .RN(n5691), .Q(\i_MIPS/Register/register[6][27] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][28]  ( .D(\i_MIPS/Register/n944 ), 
        .CK(clk), .RN(n5691), .Q(\i_MIPS/Register/register[6][28] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][29]  ( .D(\i_MIPS/Register/n945 ), 
        .CK(clk), .RN(n5691), .Q(\i_MIPS/Register/register[6][29] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][30]  ( .D(\i_MIPS/Register/n946 ), 
        .CK(clk), .RN(n5691), .Q(\i_MIPS/Register/register[6][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][31]  ( .D(\i_MIPS/Register/n947 ), 
        .CK(clk), .RN(n5692), .Q(\i_MIPS/Register/register[6][31] ) );
  DFFRX1 \i_MIPS/Register/register_reg[5][0]  ( .D(\i_MIPS/Register/n948 ), 
        .CK(clk), .RN(n5692), .Q(\i_MIPS/Register/register[5][0] ) );
  DFFRX1 \i_MIPS/Register/register_reg[4][1]  ( .D(\i_MIPS/Register/n981 ), 
        .CK(clk), .RN(n5694), .Q(\i_MIPS/Register/register[4][1] ) );
  DFFRX1 \i_MIPS/Register/register_reg[4][19]  ( .D(\i_MIPS/Register/n999 ), 
        .CK(clk), .RN(n5696), .Q(\i_MIPS/Register/register[4][19] ) );
  DFFRX1 \i_MIPS/Register/register_reg[4][30]  ( .D(\i_MIPS/Register/n1010 ), 
        .CK(clk), .RN(n5697), .Q(\i_MIPS/Register/register[4][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[3][0]  ( .D(\i_MIPS/Register/n1012 ), 
        .CK(clk), .RN(n5697), .Q(\i_MIPS/Register/register[3][0] ) );
  DFFRX1 \i_MIPS/Register/register_reg[1][0]  ( .D(\i_MIPS/Register/n1076 ), 
        .CK(clk), .RN(n5702), .Q(\i_MIPS/Register/register[1][0] ) );
  DFFRX1 \i_MIPS/Register/register_reg[0][1]  ( .D(\i_MIPS/Register/n1109 ), 
        .CK(clk), .RN(n5705), .Q(\i_MIPS/Register/register[0][1] ) );
  DFFRX1 \i_MIPS/Register/register_reg[0][19]  ( .D(\i_MIPS/Register/n1127 ), 
        .CK(clk), .RN(n5707), .Q(\i_MIPS/Register/register[0][19] ) );
  DFFRX1 \i_MIPS/Register/register_reg[0][30]  ( .D(\i_MIPS/Register/n1138 ), 
        .CK(clk), .RN(n5707), .Q(\i_MIPS/Register/register[0][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[28][2]  ( .D(\i_MIPS/Register/n214 ), 
        .CK(clk), .RN(n5630), .Q(\i_MIPS/Register/register[28][2] ), .QN(n604)
         );
  DFFRX1 \i_MIPS/Register/register_reg[28][3]  ( .D(\i_MIPS/Register/n215 ), 
        .CK(clk), .RN(n5631), .Q(\i_MIPS/Register/register[28][3] ), .QN(n601)
         );
  DFFRX1 \i_MIPS/Register/register_reg[28][4]  ( .D(\i_MIPS/Register/n216 ), 
        .CK(clk), .RN(n5631), .Q(\i_MIPS/Register/register[28][4] ), .QN(n605)
         );
  DFFRX1 \i_MIPS/Register/register_reg[28][5]  ( .D(\i_MIPS/Register/n217 ), 
        .CK(clk), .RN(n5631), .Q(\i_MIPS/Register/register[28][5] ), .QN(n670)
         );
  DFFRX1 \i_MIPS/Register/register_reg[28][6]  ( .D(\i_MIPS/Register/n218 ), 
        .CK(clk), .RN(n5631), .Q(\i_MIPS/Register/register[28][6] ), .QN(n674)
         );
  DFFRX1 \i_MIPS/Register/register_reg[28][7]  ( .D(\i_MIPS/Register/n219 ), 
        .CK(clk), .RN(n5631), .Q(\i_MIPS/Register/register[28][7] ), .QN(n671)
         );
  DFFRX1 \i_MIPS/Register/register_reg[28][8]  ( .D(\i_MIPS/Register/n220 ), 
        .CK(clk), .RN(n5631), .Q(\i_MIPS/Register/register[28][8] ), .QN(n676)
         );
  DFFRX1 \i_MIPS/Register/register_reg[28][9]  ( .D(\i_MIPS/Register/n221 ), 
        .CK(clk), .RN(n5631), .Q(\i_MIPS/Register/register[28][9] ), .QN(n675)
         );
  DFFRX1 \i_MIPS/Register/register_reg[28][10]  ( .D(\i_MIPS/Register/n222 ), 
        .CK(clk), .RN(n5631), .Q(\i_MIPS/Register/register[28][10] ), .QN(n678) );
  DFFRX1 \i_MIPS/Register/register_reg[28][11]  ( .D(\i_MIPS/Register/n223 ), 
        .CK(clk), .RN(n5631), .Q(\i_MIPS/Register/register[28][11] ), .QN(n607) );
  DFFRX1 \i_MIPS/Register/register_reg[28][12]  ( .D(\i_MIPS/Register/n224 ), 
        .CK(clk), .RN(n5631), .Q(\i_MIPS/Register/register[28][12] ), .QN(n677) );
  DFFRX1 \i_MIPS/Register/register_reg[28][13]  ( .D(\i_MIPS/Register/n225 ), 
        .CK(clk), .RN(n5631), .Q(\i_MIPS/Register/register[28][13] ), .QN(n598) );
  DFFRX1 \i_MIPS/Register/register_reg[28][14]  ( .D(\i_MIPS/Register/n226 ), 
        .CK(clk), .RN(n5631), .Q(\i_MIPS/Register/register[28][14] ), .QN(n673) );
  DFFRX1 \i_MIPS/Register/register_reg[28][15]  ( .D(\i_MIPS/Register/n227 ), 
        .CK(clk), .RN(n5632), .Q(\i_MIPS/Register/register[28][15] ), .QN(n672) );
  DFFRX1 \i_MIPS/Register/register_reg[28][16]  ( .D(\i_MIPS/Register/n228 ), 
        .CK(clk), .RN(n5632), .Q(\i_MIPS/Register/register[28][16] ), .QN(n330) );
  DFFRX1 \i_MIPS/Register/register_reg[28][17]  ( .D(\i_MIPS/Register/n229 ), 
        .CK(clk), .RN(n5632), .Q(\i_MIPS/Register/register[28][17] ), .QN(n679) );
  DFFRX1 \i_MIPS/Register/register_reg[28][18]  ( .D(\i_MIPS/Register/n230 ), 
        .CK(clk), .RN(n5632), .Q(\i_MIPS/Register/register[28][18] ), .QN(n680) );
  DFFRX1 \i_MIPS/Register/register_reg[28][20]  ( .D(\i_MIPS/Register/n232 ), 
        .CK(clk), .RN(n5632), .Q(\i_MIPS/Register/register[28][20] ), .QN(n602) );
  DFFRX1 \i_MIPS/Register/register_reg[28][21]  ( .D(\i_MIPS/Register/n233 ), 
        .CK(clk), .RN(n5632), .Q(\i_MIPS/Register/register[28][21] ), .QN(n603) );
  DFFRX1 \i_MIPS/Register/register_reg[28][22]  ( .D(\i_MIPS/Register/n234 ), 
        .CK(clk), .RN(n5632), .Q(\i_MIPS/Register/register[28][22] ), .QN(n600) );
  DFFRX1 \i_MIPS/Register/register_reg[28][23]  ( .D(\i_MIPS/Register/n235 ), 
        .CK(clk), .RN(n5632), .Q(\i_MIPS/Register/register[28][23] ), .QN(n327) );
  DFFRX1 \i_MIPS/Register/register_reg[28][25]  ( .D(\i_MIPS/Register/n237 ), 
        .CK(clk), .RN(n5632), .Q(\i_MIPS/Register/register[28][25] ), .QN(n346) );
  DFFRX1 \i_MIPS/Register/register_reg[28][26]  ( .D(\i_MIPS/Register/n238 ), 
        .CK(clk), .RN(n5632), .Q(\i_MIPS/Register/register[28][26] ), .QN(n331) );
  DFFRX1 \i_MIPS/Register/register_reg[28][27]  ( .D(\i_MIPS/Register/n239 ), 
        .CK(clk), .RN(n5633), .Q(\i_MIPS/Register/register[28][27] ), .QN(n608) );
  DFFRX1 \i_MIPS/Register/register_reg[28][28]  ( .D(\i_MIPS/Register/n240 ), 
        .CK(clk), .RN(n5633), .Q(\i_MIPS/Register/register[28][28] ), .QN(n606) );
  DFFRX1 \i_MIPS/Register/register_reg[28][29]  ( .D(\i_MIPS/Register/n241 ), 
        .CK(clk), .RN(n5633), .Q(\i_MIPS/Register/register[28][29] ), .QN(n635) );
  DFFRX1 \i_MIPS/Register/register_reg[28][31]  ( .D(\i_MIPS/Register/n243 ), 
        .CK(clk), .RN(n5633), .Q(\i_MIPS/Register/register[28][31] ), .QN(n431) );
  DFFRX1 \i_MIPS/Register/register_reg[27][8]  ( .D(\i_MIPS/Register/n252 ), 
        .CK(clk), .RN(n5634), .Q(\i_MIPS/Register/register[27][8] ), .QN(n499)
         );
  DFFRX1 \i_MIPS/Register/register_reg[27][15]  ( .D(\i_MIPS/Register/n259 ), 
        .CK(clk), .RN(n5634), .Q(\i_MIPS/Register/register[27][15] ), .QN(n537) );
  DFFRX1 \i_MIPS/Register/register_reg[27][17]  ( .D(\i_MIPS/Register/n261 ), 
        .CK(clk), .RN(n5634), .Q(\i_MIPS/Register/register[27][17] ), .QN(n494) );
  DFFRX1 \i_MIPS/Register/register_reg[27][31]  ( .D(\i_MIPS/Register/n275 ), 
        .CK(clk), .RN(n5636), .Q(\i_MIPS/Register/register[27][31] ), .QN(n543) );
  DFFRX1 \i_MIPS/Register/register_reg[24][2]  ( .D(\i_MIPS/Register/n342 ), 
        .CK(clk), .RN(n5641), .Q(\i_MIPS/Register/register[24][2] ), .QN(n626)
         );
  DFFRX1 \i_MIPS/Register/register_reg[24][4]  ( .D(\i_MIPS/Register/n344 ), 
        .CK(clk), .RN(n5641), .Q(\i_MIPS/Register/register[24][4] ), .QN(n268)
         );
  DFFRX1 \i_MIPS/Register/register_reg[24][5]  ( .D(\i_MIPS/Register/n345 ), 
        .CK(clk), .RN(n5641), .Q(\i_MIPS/Register/register[24][5] ), .QN(n275)
         );
  DFFRX1 \i_MIPS/Register/register_reg[24][6]  ( .D(\i_MIPS/Register/n346 ), 
        .CK(clk), .RN(n5641), .Q(\i_MIPS/Register/register[24][6] ), .QN(n686)
         );
  DFFRX1 \i_MIPS/Register/register_reg[24][7]  ( .D(\i_MIPS/Register/n347 ), 
        .CK(clk), .RN(n5642), .Q(\i_MIPS/Register/register[24][7] ), .QN(n685)
         );
  DFFRX1 \i_MIPS/Register/register_reg[24][8]  ( .D(\i_MIPS/Register/n348 ), 
        .CK(clk), .RN(n5642), .Q(\i_MIPS/Register/register[24][8] ), .QN(n479)
         );
  DFFRX1 \i_MIPS/Register/register_reg[24][9]  ( .D(\i_MIPS/Register/n349 ), 
        .CK(clk), .RN(n5642), .Q(\i_MIPS/Register/register[24][9] ), .QN(n687)
         );
  DFFRX1 \i_MIPS/Register/register_reg[24][10]  ( .D(\i_MIPS/Register/n350 ), 
        .CK(clk), .RN(n5642), .Q(\i_MIPS/Register/register[24][10] ), .QN(n276) );
  DFFRX1 \i_MIPS/Register/register_reg[24][11]  ( .D(\i_MIPS/Register/n351 ), 
        .CK(clk), .RN(n5642), .Q(\i_MIPS/Register/register[24][11] ), .QN(n270) );
  DFFRX1 \i_MIPS/Register/register_reg[24][12]  ( .D(\i_MIPS/Register/n352 ), 
        .CK(clk), .RN(n5642), .Q(\i_MIPS/Register/register[24][12] ), .QN(n513) );
  DFFRX1 \i_MIPS/Register/register_reg[24][13]  ( .D(\i_MIPS/Register/n353 ), 
        .CK(clk), .RN(n5642), .Q(\i_MIPS/Register/register[24][13] ), .QN(n628) );
  DFFRX1 \i_MIPS/Register/register_reg[24][14]  ( .D(\i_MIPS/Register/n354 ), 
        .CK(clk), .RN(n5642), .Q(\i_MIPS/Register/register[24][14] ), .QN(n274) );
  DFFRX1 \i_MIPS/Register/register_reg[24][15]  ( .D(\i_MIPS/Register/n355 ), 
        .CK(clk), .RN(n5642), .Q(\i_MIPS/Register/register[24][15] ), .QN(n277) );
  DFFRX1 \i_MIPS/Register/register_reg[24][16]  ( .D(\i_MIPS/Register/n356 ), 
        .CK(clk), .RN(n5642), .Q(\i_MIPS/Register/register[24][16] ), .QN(n614) );
  DFFRX1 \i_MIPS/Register/register_reg[24][17]  ( .D(\i_MIPS/Register/n357 ), 
        .CK(clk), .RN(n5642), .Q(\i_MIPS/Register/register[24][17] ), .QN(n688) );
  DFFRX1 \i_MIPS/Register/register_reg[24][18]  ( .D(\i_MIPS/Register/n358 ), 
        .CK(clk), .RN(n5642), .Q(\i_MIPS/Register/register[24][18] ), .QN(n690) );
  DFFRX1 \i_MIPS/Register/register_reg[24][20]  ( .D(\i_MIPS/Register/n360 ), 
        .CK(clk), .RN(n5643), .Q(\i_MIPS/Register/register[24][20] ), .QN(n622) );
  DFFRX1 \i_MIPS/Register/register_reg[24][21]  ( .D(\i_MIPS/Register/n361 ), 
        .CK(clk), .RN(n5643), .Q(\i_MIPS/Register/register[24][21] ), .QN(n623) );
  DFFRX1 \i_MIPS/Register/register_reg[24][22]  ( .D(\i_MIPS/Register/n362 ), 
        .CK(clk), .RN(n5643), .Q(\i_MIPS/Register/register[24][22] ), .QN(n618) );
  DFFRX1 \i_MIPS/Register/register_reg[24][23]  ( .D(\i_MIPS/Register/n363 ), 
        .CK(clk), .RN(n5643), .Q(\i_MIPS/Register/register[24][23] ), .QN(n616) );
  DFFRX1 \i_MIPS/Register/register_reg[24][25]  ( .D(\i_MIPS/Register/n365 ), 
        .CK(clk), .RN(n5643), .Q(\i_MIPS/Register/register[24][25] ), .QN(n477) );
  DFFRX1 \i_MIPS/Register/register_reg[24][26]  ( .D(\i_MIPS/Register/n366 ), 
        .CK(clk), .RN(n5643), .Q(\i_MIPS/Register/register[24][26] ), .QN(n629) );
  DFFRX1 \i_MIPS/Register/register_reg[24][27]  ( .D(\i_MIPS/Register/n367 ), 
        .CK(clk), .RN(n5643), .Q(\i_MIPS/Register/register[24][27] ), .QN(n633) );
  DFFRX1 \i_MIPS/Register/register_reg[24][28]  ( .D(\i_MIPS/Register/n368 ), 
        .CK(clk), .RN(n5643), .Q(\i_MIPS/Register/register[24][28] ), .QN(n631) );
  DFFRX1 \i_MIPS/Register/register_reg[24][29]  ( .D(\i_MIPS/Register/n369 ), 
        .CK(clk), .RN(n5643), .Q(\i_MIPS/Register/register[24][29] ), .QN(n609) );
  DFFRX1 \i_MIPS/Register/register_reg[24][31]  ( .D(\i_MIPS/Register/n371 ), 
        .CK(clk), .RN(n5644), .Q(\i_MIPS/Register/register[24][31] ), .QN(n474) );
  DFFRX1 \i_MIPS/Register/register_reg[15][8]  ( .D(\i_MIPS/Register/n636 ), 
        .CK(clk), .RN(n5666), .Q(\i_MIPS/Register/register[15][8] ), .QN(n310)
         );
  DFFRX1 \i_MIPS/Register/register_reg[15][9]  ( .D(\i_MIPS/Register/n637 ), 
        .CK(clk), .RN(n5666), .Q(\i_MIPS/Register/register[15][9] ), .QN(n309)
         );
  DFFRX1 \i_MIPS/Register/register_reg[15][12]  ( .D(\i_MIPS/Register/n640 ), 
        .CK(clk), .RN(n5666), .Q(\i_MIPS/Register/register[15][12] ), .QN(n662) );
  DFFRX1 \i_MIPS/Register/register_reg[15][15]  ( .D(\i_MIPS/Register/n643 ), 
        .CK(clk), .RN(n5666), .Q(\i_MIPS/Register/register[15][15] ), .QN(n665) );
  DFFRX1 \i_MIPS/Register/register_reg[15][17]  ( .D(\i_MIPS/Register/n645 ), 
        .CK(clk), .RN(n5666), .Q(\i_MIPS/Register/register[15][17] ), .QN(n215) );
  DFFRX1 \i_MIPS/Register/register_reg[15][18]  ( .D(\i_MIPS/Register/n646 ), 
        .CK(clk), .RN(n5666), .Q(\i_MIPS/Register/register[15][18] ), .QN(n214) );
  DFFRX1 \i_MIPS/Register/register_reg[15][31]  ( .D(\i_MIPS/Register/n659 ), 
        .CK(clk), .RN(n5668), .Q(\i_MIPS/Register/register[15][31] ), .QN(n658) );
  DFFRX1 \i_MIPS/Register/register_reg[12][2]  ( .D(\i_MIPS/Register/n726 ), 
        .CK(clk), .RN(n5673), .Q(\i_MIPS/Register/register[12][2] ), .QN(n643)
         );
  DFFRX1 \i_MIPS/Register/register_reg[12][3]  ( .D(\i_MIPS/Register/n727 ), 
        .CK(clk), .RN(n5673), .Q(\i_MIPS/Register/register[12][3] ), .QN(n641)
         );
  DFFRX1 \i_MIPS/Register/register_reg[12][4]  ( .D(\i_MIPS/Register/n728 ), 
        .CK(clk), .RN(n5673), .Q(\i_MIPS/Register/register[12][4] ), .QN(n644)
         );
  DFFRX1 \i_MIPS/Register/register_reg[12][5]  ( .D(\i_MIPS/Register/n729 ), 
        .CK(clk), .RN(n5673), .Q(\i_MIPS/Register/register[12][5] ), .QN(n693)
         );
  DFFRX1 \i_MIPS/Register/register_reg[12][6]  ( .D(\i_MIPS/Register/n730 ), 
        .CK(clk), .RN(n5673), .Q(\i_MIPS/Register/register[12][6] ), .QN(n695)
         );
  DFFRX1 \i_MIPS/Register/register_reg[12][7]  ( .D(\i_MIPS/Register/n731 ), 
        .CK(clk), .RN(n5674), .Q(\i_MIPS/Register/register[12][7] ), .QN(n694)
         );
  DFFRX1 \i_MIPS/Register/register_reg[12][8]  ( .D(\i_MIPS/Register/n732 ), 
        .CK(clk), .RN(n5674), .Q(\i_MIPS/Register/register[12][8] ), .QN(n473)
         );
  DFFRX1 \i_MIPS/Register/register_reg[12][9]  ( .D(\i_MIPS/Register/n733 ), 
        .CK(clk), .RN(n5674), .Q(\i_MIPS/Register/register[12][9] ), .QN(n696)
         );
  DFFRX1 \i_MIPS/Register/register_reg[12][10]  ( .D(\i_MIPS/Register/n734 ), 
        .CK(clk), .RN(n5674), .Q(\i_MIPS/Register/register[12][10] ), .QN(n698) );
  DFFRX1 \i_MIPS/Register/register_reg[12][11]  ( .D(\i_MIPS/Register/n735 ), 
        .CK(clk), .RN(n5674), .Q(\i_MIPS/Register/register[12][11] ), .QN(n699) );
  DFFRX1 \i_MIPS/Register/register_reg[12][12]  ( .D(\i_MIPS/Register/n736 ), 
        .CK(clk), .RN(n5674), .Q(\i_MIPS/Register/register[12][12] ), .QN(n697) );
  DFFRX1 \i_MIPS/Register/register_reg[12][13]  ( .D(\i_MIPS/Register/n737 ), 
        .CK(clk), .RN(n5674), .Q(\i_MIPS/Register/register[12][13] ), .QN(n638) );
  DFFRX1 \i_MIPS/Register/register_reg[12][14]  ( .D(\i_MIPS/Register/n738 ), 
        .CK(clk), .RN(n5674), .Q(\i_MIPS/Register/register[12][14] ), .QN(n436) );
  DFFRX1 \i_MIPS/Register/register_reg[12][15]  ( .D(\i_MIPS/Register/n739 ), 
        .CK(clk), .RN(n5674), .Q(\i_MIPS/Register/register[12][15] ), .QN(n637) );
  DFFRX1 \i_MIPS/Register/register_reg[12][16]  ( .D(\i_MIPS/Register/n740 ), 
        .CK(clk), .RN(n5674), .Q(\i_MIPS/Register/register[12][16] ), .QN(n329) );
  DFFRX1 \i_MIPS/Register/register_reg[12][17]  ( .D(\i_MIPS/Register/n741 ), 
        .CK(clk), .RN(n5674), .Q(\i_MIPS/Register/register[12][17] ), .QN(n700) );
  DFFRX1 \i_MIPS/Register/register_reg[12][18]  ( .D(\i_MIPS/Register/n742 ), 
        .CK(clk), .RN(n5674), .Q(\i_MIPS/Register/register[12][18] ), .QN(n701) );
  DFFRX1 \i_MIPS/Register/register_reg[12][20]  ( .D(\i_MIPS/Register/n744 ), 
        .CK(clk), .RN(n5675), .Q(\i_MIPS/Register/register[12][20] ), .QN(n332) );
  DFFRX1 \i_MIPS/Register/register_reg[12][21]  ( .D(\i_MIPS/Register/n745 ), 
        .CK(clk), .RN(n5675), .Q(\i_MIPS/Register/register[12][21] ), .QN(n642) );
  DFFRX1 \i_MIPS/Register/register_reg[12][22]  ( .D(\i_MIPS/Register/n746 ), 
        .CK(clk), .RN(n5675), .Q(\i_MIPS/Register/register[12][22] ), .QN(n640) );
  DFFRX1 \i_MIPS/Register/register_reg[12][23]  ( .D(\i_MIPS/Register/n747 ), 
        .CK(clk), .RN(n5675), .Q(\i_MIPS/Register/register[12][23] ), .QN(n328) );
  DFFRX1 \i_MIPS/Register/register_reg[12][25]  ( .D(\i_MIPS/Register/n749 ), 
        .CK(clk), .RN(n5675), .Q(\i_MIPS/Register/register[12][25] ), .QN(n429) );
  DFFRX1 \i_MIPS/Register/register_reg[12][26]  ( .D(\i_MIPS/Register/n750 ), 
        .CK(clk), .RN(n5675), .Q(\i_MIPS/Register/register[12][26] ), .QN(n489) );
  DFFRX1 \i_MIPS/Register/register_reg[12][27]  ( .D(\i_MIPS/Register/n751 ), 
        .CK(clk), .RN(n5675), .Q(\i_MIPS/Register/register[12][27] ), .QN(n646) );
  DFFRX1 \i_MIPS/Register/register_reg[12][28]  ( .D(\i_MIPS/Register/n752 ), 
        .CK(clk), .RN(n5675), .Q(\i_MIPS/Register/register[12][28] ), .QN(n645) );
  DFFRX1 \i_MIPS/Register/register_reg[12][29]  ( .D(\i_MIPS/Register/n753 ), 
        .CK(clk), .RN(n5675), .Q(\i_MIPS/Register/register[12][29] ), .QN(n636) );
  DFFRX1 \i_MIPS/Register/register_reg[12][31]  ( .D(\i_MIPS/Register/n755 ), 
        .CK(clk), .RN(n5676), .Q(\i_MIPS/Register/register[12][31] ), .QN(n430) );
  DFFRX1 \i_MIPS/Register/register_reg[11][8]  ( .D(\i_MIPS/Register/n764 ), 
        .CK(clk), .RN(n5676), .Q(\i_MIPS/Register/register[11][8] ), .QN(n500)
         );
  DFFRX1 \i_MIPS/Register/register_reg[11][15]  ( .D(\i_MIPS/Register/n771 ), 
        .CK(clk), .RN(n5677), .Q(\i_MIPS/Register/register[11][15] ), .QN(n538) );
  DFFRX1 \i_MIPS/Register/register_reg[11][17]  ( .D(\i_MIPS/Register/n773 ), 
        .CK(clk), .RN(n5677), .Q(\i_MIPS/Register/register[11][17] ), .QN(n495) );
  DFFRX1 \i_MIPS/Register/register_reg[11][31]  ( .D(\i_MIPS/Register/n787 ), 
        .CK(clk), .RN(n5678), .Q(\i_MIPS/Register/register[11][31] ), .QN(n544) );
  DFFRX1 \i_MIPS/Register/register_reg[8][2]  ( .D(\i_MIPS/Register/n854 ), 
        .CK(clk), .RN(n5684), .Q(\i_MIPS/Register/register[8][2] ), .QN(n627)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][4]  ( .D(\i_MIPS/Register/n856 ), 
        .CK(clk), .RN(n5684), .Q(\i_MIPS/Register/register[8][4] ), .QN(n269)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][5]  ( .D(\i_MIPS/Register/n857 ), 
        .CK(clk), .RN(n5684), .Q(\i_MIPS/Register/register[8][5] ), .QN(n272)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][6]  ( .D(\i_MIPS/Register/n858 ), 
        .CK(clk), .RN(n5684), .Q(\i_MIPS/Register/register[8][6] ), .QN(n682)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][7]  ( .D(\i_MIPS/Register/n859 ), 
        .CK(clk), .RN(n5684), .Q(\i_MIPS/Register/register[8][7] ), .QN(n681)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][8]  ( .D(\i_MIPS/Register/n860 ), 
        .CK(clk), .RN(n5684), .Q(\i_MIPS/Register/register[8][8] ), .QN(n476)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][9]  ( .D(\i_MIPS/Register/n861 ), 
        .CK(clk), .RN(n5684), .Q(\i_MIPS/Register/register[8][9] ), .QN(n683)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][10]  ( .D(\i_MIPS/Register/n862 ), 
        .CK(clk), .RN(n5684), .Q(\i_MIPS/Register/register[8][10] ), .QN(n278)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][11]  ( .D(\i_MIPS/Register/n863 ), 
        .CK(clk), .RN(n5685), .Q(\i_MIPS/Register/register[8][11] ), .QN(n271)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][12]  ( .D(\i_MIPS/Register/n864 ), 
        .CK(clk), .RN(n5685), .Q(\i_MIPS/Register/register[8][12] ), .QN(n684)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][13]  ( .D(\i_MIPS/Register/n865 ), 
        .CK(clk), .RN(n5685), .Q(\i_MIPS/Register/register[8][13] ), .QN(n611)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][14]  ( .D(\i_MIPS/Register/n866 ), 
        .CK(clk), .RN(n5685), .Q(\i_MIPS/Register/register[8][14] ), .QN(n273)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][15]  ( .D(\i_MIPS/Register/n867 ), 
        .CK(clk), .RN(n5685), .Q(\i_MIPS/Register/register[8][15] ), .QN(n267)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][16]  ( .D(\i_MIPS/Register/n868 ), 
        .CK(clk), .RN(n5685), .Q(\i_MIPS/Register/register[8][16] ), .QN(n615)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][17]  ( .D(\i_MIPS/Register/n869 ), 
        .CK(clk), .RN(n5685), .Q(\i_MIPS/Register/register[8][17] ), .QN(n689)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][18]  ( .D(\i_MIPS/Register/n870 ), 
        .CK(clk), .RN(n5685), .Q(\i_MIPS/Register/register[8][18] ), .QN(n691)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][20]  ( .D(\i_MIPS/Register/n872 ), 
        .CK(clk), .RN(n5685), .Q(\i_MIPS/Register/register[8][20] ), .QN(n624)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][21]  ( .D(\i_MIPS/Register/n873 ), 
        .CK(clk), .RN(n5685), .Q(\i_MIPS/Register/register[8][21] ), .QN(n625)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][22]  ( .D(\i_MIPS/Register/n874 ), 
        .CK(clk), .RN(n5685), .Q(\i_MIPS/Register/register[8][22] ), .QN(n619)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][23]  ( .D(\i_MIPS/Register/n875 ), 
        .CK(clk), .RN(n5686), .Q(\i_MIPS/Register/register[8][23] ), .QN(n617)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][25]  ( .D(\i_MIPS/Register/n877 ), 
        .CK(clk), .RN(n5686), .Q(\i_MIPS/Register/register[8][25] ), .QN(n478)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][26]  ( .D(\i_MIPS/Register/n878 ), 
        .CK(clk), .RN(n5686), .Q(\i_MIPS/Register/register[8][26] ), .QN(n630)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][27]  ( .D(\i_MIPS/Register/n879 ), 
        .CK(clk), .RN(n5686), .Q(\i_MIPS/Register/register[8][27] ), .QN(n634)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][28]  ( .D(\i_MIPS/Register/n880 ), 
        .CK(clk), .RN(n5686), .Q(\i_MIPS/Register/register[8][28] ), .QN(n632)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][29]  ( .D(\i_MIPS/Register/n881 ), 
        .CK(clk), .RN(n5686), .Q(\i_MIPS/Register/register[8][29] ), .QN(n610)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][31]  ( .D(\i_MIPS/Register/n883 ), 
        .CK(clk), .RN(n5686), .Q(\i_MIPS/Register/register[8][31] ), .QN(n475)
         );
  DFFRX1 \i_MIPS/Register/register_reg[23][8]  ( .D(\i_MIPS/Register/n380 ), 
        .CK(clk), .RN(n5644), .Q(\i_MIPS/Register/register[23][8] ), .QN(n2070) );
  DFFRX1 \i_MIPS/Register/register_reg[23][9]  ( .D(\i_MIPS/Register/n381 ), 
        .CK(clk), .RN(n5644), .Q(\i_MIPS/Register/register[23][9] ), .QN(n2066) );
  DFFRX1 \i_MIPS/Register/register_reg[23][12]  ( .D(\i_MIPS/Register/n384 ), 
        .CK(clk), .RN(n5645), .Q(\i_MIPS/Register/register[23][12] ), .QN(
        n2186) );
  DFFRX1 \i_MIPS/Register/register_reg[23][15]  ( .D(\i_MIPS/Register/n387 ), 
        .CK(clk), .RN(n5645), .Q(\i_MIPS/Register/register[23][15] ), .QN(
        n2191) );
  DFFRX1 \i_MIPS/Register/register_reg[23][17]  ( .D(\i_MIPS/Register/n389 ), 
        .CK(clk), .RN(n5645), .Q(\i_MIPS/Register/register[23][17] ), .QN(n734) );
  DFFRX1 \i_MIPS/Register/register_reg[23][31]  ( .D(\i_MIPS/Register/n403 ), 
        .CK(clk), .RN(n5646), .Q(\i_MIPS/Register/register[23][31] ), .QN(
        n2180) );
  DFFRX1 \i_MIPS/Register/register_reg[20][2]  ( .D(\i_MIPS/Register/n470 ), 
        .CK(clk), .RN(n5652), .Q(\i_MIPS/Register/register[20][2] ), .QN(n2124) );
  DFFRX1 \i_MIPS/Register/register_reg[20][4]  ( .D(\i_MIPS/Register/n472 ), 
        .CK(clk), .RN(n5652), .Q(\i_MIPS/Register/register[20][4] ), .QN(n2125) );
  DFFRX1 \i_MIPS/Register/register_reg[20][5]  ( .D(\i_MIPS/Register/n473 ), 
        .CK(clk), .RN(n5652), .Q(\i_MIPS/Register/register[20][5] ), .QN(n2199) );
  DFFRX1 \i_MIPS/Register/register_reg[20][6]  ( .D(\i_MIPS/Register/n474 ), 
        .CK(clk), .RN(n5652), .Q(\i_MIPS/Register/register[20][6] ), .QN(n2203) );
  DFFRX1 \i_MIPS/Register/register_reg[20][7]  ( .D(\i_MIPS/Register/n475 ), 
        .CK(clk), .RN(n5652), .Q(\i_MIPS/Register/register[20][7] ), .QN(n2200) );
  DFFRX1 \i_MIPS/Register/register_reg[20][8]  ( .D(\i_MIPS/Register/n476 ), 
        .CK(clk), .RN(n5652), .Q(\i_MIPS/Register/register[20][8] ), .QN(n2205) );
  DFFRX1 \i_MIPS/Register/register_reg[20][9]  ( .D(\i_MIPS/Register/n477 ), 
        .CK(clk), .RN(n5652), .Q(\i_MIPS/Register/register[20][9] ), .QN(n2204) );
  DFFRX1 \i_MIPS/Register/register_reg[20][10]  ( .D(\i_MIPS/Register/n478 ), 
        .CK(clk), .RN(n5652), .Q(\i_MIPS/Register/register[20][10] ), .QN(
        n2207) );
  DFFRX1 \i_MIPS/Register/register_reg[20][11]  ( .D(\i_MIPS/Register/n479 ), 
        .CK(clk), .RN(n5653), .Q(\i_MIPS/Register/register[20][11] ), .QN(
        n2127) );
  DFFRX1 \i_MIPS/Register/register_reg[20][12]  ( .D(\i_MIPS/Register/n480 ), 
        .CK(clk), .RN(n5653), .Q(\i_MIPS/Register/register[20][12] ), .QN(
        n2206) );
  DFFRX1 \i_MIPS/Register/register_reg[20][13]  ( .D(\i_MIPS/Register/n481 ), 
        .CK(clk), .RN(n5653), .Q(\i_MIPS/Register/register[20][13] ), .QN(
        n2118) );
  DFFRX1 \i_MIPS/Register/register_reg[20][14]  ( .D(\i_MIPS/Register/n482 ), 
        .CK(clk), .RN(n5653), .Q(\i_MIPS/Register/register[20][14] ), .QN(
        n2202) );
  DFFRX1 \i_MIPS/Register/register_reg[20][15]  ( .D(\i_MIPS/Register/n483 ), 
        .CK(clk), .RN(n5653), .Q(\i_MIPS/Register/register[20][15] ), .QN(
        n2201) );
  DFFRX1 \i_MIPS/Register/register_reg[20][17]  ( .D(\i_MIPS/Register/n485 ), 
        .CK(clk), .RN(n5653), .Q(\i_MIPS/Register/register[20][17] ), .QN(
        n2208) );
  DFFRX1 \i_MIPS/Register/register_reg[20][18]  ( .D(\i_MIPS/Register/n486 ), 
        .CK(clk), .RN(n5653), .Q(\i_MIPS/Register/register[20][18] ), .QN(
        n2209) );
  DFFRX1 \i_MIPS/Register/register_reg[20][20]  ( .D(\i_MIPS/Register/n488 ), 
        .CK(clk), .RN(n5653), .Q(\i_MIPS/Register/register[20][20] ), .QN(
        n2122) );
  DFFRX1 \i_MIPS/Register/register_reg[20][21]  ( .D(\i_MIPS/Register/n489 ), 
        .CK(clk), .RN(n5653), .Q(\i_MIPS/Register/register[20][21] ), .QN(
        n2123) );
  DFFRX1 \i_MIPS/Register/register_reg[20][25]  ( .D(\i_MIPS/Register/n493 ), 
        .CK(clk), .RN(n5654), .Q(\i_MIPS/Register/register[20][25] ), .QN(
        n1928) );
  DFFRX1 \i_MIPS/Register/register_reg[20][26]  ( .D(\i_MIPS/Register/n494 ), 
        .CK(clk), .RN(n5654), .Q(\i_MIPS/Register/register[20][26] ), .QN(
        n1908) );
  DFFRX1 \i_MIPS/Register/register_reg[20][27]  ( .D(\i_MIPS/Register/n495 ), 
        .CK(clk), .RN(n5654), .Q(\i_MIPS/Register/register[20][27] ), .QN(
        n2128) );
  DFFRX1 \i_MIPS/Register/register_reg[20][28]  ( .D(\i_MIPS/Register/n496 ), 
        .CK(clk), .RN(n5654), .Q(\i_MIPS/Register/register[20][28] ), .QN(
        n2126) );
  DFFRX1 \i_MIPS/Register/register_reg[20][29]  ( .D(\i_MIPS/Register/n497 ), 
        .CK(clk), .RN(n5654), .Q(\i_MIPS/Register/register[20][29] ), .QN(
        n2156) );
  DFFRX1 \i_MIPS/Register/register_reg[20][31]  ( .D(\i_MIPS/Register/n499 ), 
        .CK(clk), .RN(n5654), .Q(\i_MIPS/Register/register[20][31] ), .QN(
        n1994) );
  DFFRX1 \i_MIPS/Register/register_reg[16][4]  ( .D(\i_MIPS/Register/n600 ), 
        .CK(clk), .RN(n5663), .Q(\i_MIPS/Register/register[16][4] ), .QN(n720)
         );
  DFFRX1 \i_MIPS/Register/register_reg[16][5]  ( .D(\i_MIPS/Register/n601 ), 
        .CK(clk), .RN(n5663), .Q(\i_MIPS/Register/register[16][5] ), .QN(n730)
         );
  DFFRX1 \i_MIPS/Register/register_reg[16][6]  ( .D(\i_MIPS/Register/n602 ), 
        .CK(clk), .RN(n5663), .Q(\i_MIPS/Register/register[16][6] ), .QN(n2215) );
  DFFRX1 \i_MIPS/Register/register_reg[16][7]  ( .D(\i_MIPS/Register/n603 ), 
        .CK(clk), .RN(n5663), .Q(\i_MIPS/Register/register[16][7] ), .QN(n2214) );
  DFFRX1 \i_MIPS/Register/register_reg[16][8]  ( .D(\i_MIPS/Register/n604 ), 
        .CK(clk), .RN(n5663), .Q(\i_MIPS/Register/register[16][8] ), .QN(n2032) );
  DFFRX1 \i_MIPS/Register/register_reg[16][9]  ( .D(\i_MIPS/Register/n605 ), 
        .CK(clk), .RN(n5663), .Q(\i_MIPS/Register/register[16][9] ), .QN(n2216) );
  DFFRX1 \i_MIPS/Register/register_reg[16][10]  ( .D(\i_MIPS/Register/n606 ), 
        .CK(clk), .RN(n5663), .Q(\i_MIPS/Register/register[16][10] ), .QN(n731) );
  DFFRX1 \i_MIPS/Register/register_reg[16][11]  ( .D(\i_MIPS/Register/n607 ), 
        .CK(clk), .RN(n5663), .Q(\i_MIPS/Register/register[16][11] ), .QN(n722) );
  DFFRX1 \i_MIPS/Register/register_reg[16][12]  ( .D(\i_MIPS/Register/n608 ), 
        .CK(clk), .RN(n5663), .Q(\i_MIPS/Register/register[16][12] ), .QN(
        n2266) );
  DFFRX1 \i_MIPS/Register/register_reg[16][13]  ( .D(\i_MIPS/Register/n609 ), 
        .CK(clk), .RN(n5663), .Q(\i_MIPS/Register/register[16][13] ), .QN(
        n2148) );
  DFFRX1 \i_MIPS/Register/register_reg[16][14]  ( .D(\i_MIPS/Register/n610 ), 
        .CK(clk), .RN(n5663), .Q(\i_MIPS/Register/register[16][14] ), .QN(n729) );
  DFFRX1 \i_MIPS/Register/register_reg[16][15]  ( .D(\i_MIPS/Register/n611 ), 
        .CK(clk), .RN(n5664), .Q(\i_MIPS/Register/register[16][15] ), .QN(n732) );
  DFFRX1 \i_MIPS/Register/register_reg[16][17]  ( .D(\i_MIPS/Register/n613 ), 
        .CK(clk), .RN(n5664), .Q(\i_MIPS/Register/register[16][17] ), .QN(
        n2217) );
  DFFRX1 \i_MIPS/Register/register_reg[16][18]  ( .D(\i_MIPS/Register/n614 ), 
        .CK(clk), .RN(n5664), .Q(\i_MIPS/Register/register[16][18] ), .QN(
        n2219) );
  DFFRX1 \i_MIPS/Register/register_reg[16][25]  ( .D(\i_MIPS/Register/n621 ), 
        .CK(clk), .RN(n5664), .Q(\i_MIPS/Register/register[16][25] ), .QN(
        n2030) );
  DFFRX1 \i_MIPS/Register/register_reg[16][26]  ( .D(\i_MIPS/Register/n622 ), 
        .CK(clk), .RN(n5664), .Q(\i_MIPS/Register/register[16][26] ), .QN(
        n2149) );
  DFFRX1 \i_MIPS/Register/register_reg[16][27]  ( .D(\i_MIPS/Register/n623 ), 
        .CK(clk), .RN(n5665), .Q(\i_MIPS/Register/register[16][27] ), .QN(
        n2153) );
  DFFRX1 \i_MIPS/Register/register_reg[16][28]  ( .D(\i_MIPS/Register/n624 ), 
        .CK(clk), .RN(n5665), .Q(\i_MIPS/Register/register[16][28] ), .QN(
        n2151) );
  DFFRX1 \i_MIPS/Register/register_reg[16][29]  ( .D(\i_MIPS/Register/n625 ), 
        .CK(clk), .RN(n5665), .Q(\i_MIPS/Register/register[16][29] ), .QN(
        n2129) );
  DFFRX1 \i_MIPS/Register/register_reg[16][31]  ( .D(\i_MIPS/Register/n627 ), 
        .CK(clk), .RN(n5665), .Q(\i_MIPS/Register/register[16][31] ), .QN(
        n2027) );
  DFFRX1 \i_MIPS/Register/register_reg[7][8]  ( .D(\i_MIPS/Register/n892 ), 
        .CK(clk), .RN(n5687), .Q(\i_MIPS/Register/register[7][8] ), .QN(n2072)
         );
  DFFRX1 \i_MIPS/Register/register_reg[7][9]  ( .D(\i_MIPS/Register/n893 ), 
        .CK(clk), .RN(n5687), .Q(\i_MIPS/Register/register[7][9] ), .QN(n2068)
         );
  DFFRX1 \i_MIPS/Register/register_reg[7][12]  ( .D(\i_MIPS/Register/n896 ), 
        .CK(clk), .RN(n5687), .Q(\i_MIPS/Register/register[7][12] ), .QN(n2187) );
  DFFRX1 \i_MIPS/Register/register_reg[7][15]  ( .D(\i_MIPS/Register/n899 ), 
        .CK(clk), .RN(n5688), .Q(\i_MIPS/Register/register[7][15] ), .QN(n2192) );
  DFFRX1 \i_MIPS/Register/register_reg[7][17]  ( .D(\i_MIPS/Register/n901 ), 
        .CK(clk), .RN(n5688), .Q(\i_MIPS/Register/register[7][17] ), .QN(n716)
         );
  DFFRX1 \i_MIPS/Register/register_reg[7][31]  ( .D(\i_MIPS/Register/n915 ), 
        .CK(clk), .RN(n5689), .Q(\i_MIPS/Register/register[7][31] ), .QN(n2182) );
  DFFRX1 \i_MIPS/Register/register_reg[4][2]  ( .D(\i_MIPS/Register/n982 ), 
        .CK(clk), .RN(n5694), .Q(\i_MIPS/Register/register[4][2] ), .QN(n2164)
         );
  DFFRX1 \i_MIPS/Register/register_reg[4][4]  ( .D(\i_MIPS/Register/n984 ), 
        .CK(clk), .RN(n5695), .Q(\i_MIPS/Register/register[4][4] ), .QN(n2165)
         );
  DFFRX1 \i_MIPS/Register/register_reg[4][5]  ( .D(\i_MIPS/Register/n985 ), 
        .CK(clk), .RN(n5695), .Q(\i_MIPS/Register/register[4][5] ), .QN(n2222)
         );
  DFFRX1 \i_MIPS/Register/register_reg[4][6]  ( .D(\i_MIPS/Register/n986 ), 
        .CK(clk), .RN(n5695), .Q(\i_MIPS/Register/register[4][6] ), .QN(n2224)
         );
  DFFRX1 \i_MIPS/Register/register_reg[4][7]  ( .D(\i_MIPS/Register/n987 ), 
        .CK(clk), .RN(n5695), .Q(\i_MIPS/Register/register[4][7] ), .QN(n2223)
         );
  DFFRX1 \i_MIPS/Register/register_reg[4][8]  ( .D(\i_MIPS/Register/n988 ), 
        .CK(clk), .RN(n5695), .Q(\i_MIPS/Register/register[4][8] ), .QN(n2039)
         );
  DFFRX1 \i_MIPS/Register/register_reg[4][9]  ( .D(\i_MIPS/Register/n989 ), 
        .CK(clk), .RN(n5695), .Q(\i_MIPS/Register/register[4][9] ), .QN(n2225)
         );
  DFFRX1 \i_MIPS/Register/register_reg[4][10]  ( .D(\i_MIPS/Register/n990 ), 
        .CK(clk), .RN(n5695), .Q(\i_MIPS/Register/register[4][10] ), .QN(n2227) );
  DFFRX1 \i_MIPS/Register/register_reg[4][11]  ( .D(\i_MIPS/Register/n991 ), 
        .CK(clk), .RN(n5695), .Q(\i_MIPS/Register/register[4][11] ), .QN(n2228) );
  DFFRX1 \i_MIPS/Register/register_reg[4][12]  ( .D(\i_MIPS/Register/n992 ), 
        .CK(clk), .RN(n5695), .Q(\i_MIPS/Register/register[4][12] ), .QN(n2226) );
  DFFRX1 \i_MIPS/Register/register_reg[4][13]  ( .D(\i_MIPS/Register/n993 ), 
        .CK(clk), .RN(n5695), .Q(\i_MIPS/Register/register[4][13] ), .QN(n2159) );
  DFFRX1 \i_MIPS/Register/register_reg[4][14]  ( .D(\i_MIPS/Register/n994 ), 
        .CK(clk), .RN(n5695), .Q(\i_MIPS/Register/register[4][14] ), .QN(n1999) );
  DFFRX1 \i_MIPS/Register/register_reg[4][15]  ( .D(\i_MIPS/Register/n995 ), 
        .CK(clk), .RN(n5696), .Q(\i_MIPS/Register/register[4][15] ), .QN(n2158) );
  DFFRX1 \i_MIPS/Register/register_reg[4][17]  ( .D(\i_MIPS/Register/n997 ), 
        .CK(clk), .RN(n5696), .Q(\i_MIPS/Register/register[4][17] ), .QN(n2229) );
  DFFRX1 \i_MIPS/Register/register_reg[4][18]  ( .D(\i_MIPS/Register/n998 ), 
        .CK(clk), .RN(n5696), .Q(\i_MIPS/Register/register[4][18] ), .QN(n2230) );
  DFFRX1 \i_MIPS/Register/register_reg[4][20]  ( .D(\i_MIPS/Register/n1000 ), 
        .CK(clk), .RN(n5696), .Q(\i_MIPS/Register/register[4][20] ), .QN(n1909) );
  DFFRX1 \i_MIPS/Register/register_reg[4][21]  ( .D(\i_MIPS/Register/n1001 ), 
        .CK(clk), .RN(n5696), .Q(\i_MIPS/Register/register[4][21] ), .QN(n2163) );
  DFFRX1 \i_MIPS/Register/register_reg[4][25]  ( .D(\i_MIPS/Register/n1005 ), 
        .CK(clk), .RN(n5696), .Q(\i_MIPS/Register/register[4][25] ), .QN(n1992) );
  DFFRX1 \i_MIPS/Register/register_reg[4][26]  ( .D(\i_MIPS/Register/n1006 ), 
        .CK(clk), .RN(n5696), .Q(\i_MIPS/Register/register[4][26] ), .QN(n2233) );
  DFFRX1 \i_MIPS/Register/register_reg[4][27]  ( .D(\i_MIPS/Register/n1007 ), 
        .CK(clk), .RN(n5697), .Q(\i_MIPS/Register/register[4][27] ), .QN(n2167) );
  DFFRX1 \i_MIPS/Register/register_reg[4][28]  ( .D(\i_MIPS/Register/n1008 ), 
        .CK(clk), .RN(n5697), .Q(\i_MIPS/Register/register[4][28] ), .QN(n2166) );
  DFFRX1 \i_MIPS/Register/register_reg[4][29]  ( .D(\i_MIPS/Register/n1009 ), 
        .CK(clk), .RN(n5697), .Q(\i_MIPS/Register/register[4][29] ), .QN(n2157) );
  DFFRX1 \i_MIPS/Register/register_reg[4][31]  ( .D(\i_MIPS/Register/n1011 ), 
        .CK(clk), .RN(n5697), .Q(\i_MIPS/Register/register[4][31] ), .QN(n1993) );
  DFFRX1 \i_MIPS/Register/register_reg[0][4]  ( .D(\i_MIPS/Register/n1112 ), 
        .CK(clk), .RN(n5705), .Q(\i_MIPS/Register/register[0][4] ), .QN(n721)
         );
  DFFRX1 \i_MIPS/Register/register_reg[0][5]  ( .D(\i_MIPS/Register/n1113 ), 
        .CK(clk), .RN(n5705), .Q(\i_MIPS/Register/register[0][5] ), .QN(n727)
         );
  DFFRX1 \i_MIPS/Register/register_reg[0][6]  ( .D(\i_MIPS/Register/n1114 ), 
        .CK(clk), .RN(n5705), .Q(\i_MIPS/Register/register[0][6] ), .QN(n2211)
         );
  DFFRX1 \i_MIPS/Register/register_reg[0][7]  ( .D(\i_MIPS/Register/n1115 ), 
        .CK(clk), .RN(n5706), .Q(\i_MIPS/Register/register[0][7] ), .QN(n2210)
         );
  DFFRX1 \i_MIPS/Register/register_reg[0][8]  ( .D(\i_MIPS/Register/n1116 ), 
        .CK(clk), .RN(n5706), .Q(\i_MIPS/Register/register[0][8] ), .QN(n2029)
         );
  DFFRX1 \i_MIPS/Register/register_reg[0][9]  ( .D(\i_MIPS/Register/n1117 ), 
        .CK(clk), .RN(n5706), .Q(\i_MIPS/Register/register[0][9] ), .QN(n2212)
         );
  DFFRX1 \i_MIPS/Register/register_reg[0][10]  ( .D(\i_MIPS/Register/n1118 ), 
        .CK(clk), .RN(n5706), .Q(\i_MIPS/Register/register[0][10] ), .QN(n733)
         );
  DFFRX1 \i_MIPS/Register/register_reg[0][11]  ( .D(\i_MIPS/Register/n1119 ), 
        .CK(clk), .RN(n5706), .Q(\i_MIPS/Register/register[0][11] ), .QN(n723)
         );
  DFFRX1 \i_MIPS/Register/register_reg[0][12]  ( .D(\i_MIPS/Register/n1120 ), 
        .CK(clk), .RN(n5706), .Q(\i_MIPS/Register/register[0][12] ), .QN(n2213) );
  DFFRX1 \i_MIPS/Register/register_reg[0][13]  ( .D(\i_MIPS/Register/n1121 ), 
        .CK(clk), .RN(n5706), .Q(\i_MIPS/Register/register[0][13] ), .QN(n2131) );
  DFFRX1 \i_MIPS/Register/register_reg[0][14]  ( .D(\i_MIPS/Register/n1122 ), 
        .CK(clk), .RN(n5706), .Q(\i_MIPS/Register/register[0][14] ), .QN(n728)
         );
  DFFRX1 \i_MIPS/Register/register_reg[0][15]  ( .D(\i_MIPS/Register/n1123 ), 
        .CK(clk), .RN(n5706), .Q(\i_MIPS/Register/register[0][15] ), .QN(n719)
         );
  DFFRX1 \i_MIPS/Register/register_reg[0][17]  ( .D(\i_MIPS/Register/n1125 ), 
        .CK(clk), .RN(n5706), .Q(\i_MIPS/Register/register[0][17] ), .QN(n2218) );
  DFFRX1 \i_MIPS/Register/register_reg[0][18]  ( .D(\i_MIPS/Register/n1126 ), 
        .CK(clk), .RN(n5706), .Q(\i_MIPS/Register/register[0][18] ), .QN(n2220) );
  DFFRX1 \i_MIPS/Register/register_reg[0][25]  ( .D(\i_MIPS/Register/n1133 ), 
        .CK(clk), .RN(n5707), .Q(\i_MIPS/Register/register[0][25] ), .QN(n2031) );
  DFFRX1 \i_MIPS/Register/register_reg[0][26]  ( .D(\i_MIPS/Register/n1134 ), 
        .CK(clk), .RN(n5707), .Q(\i_MIPS/Register/register[0][26] ), .QN(n2150) );
  DFFRX1 \i_MIPS/Register/register_reg[0][27]  ( .D(\i_MIPS/Register/n1135 ), 
        .CK(clk), .RN(n5707), .Q(\i_MIPS/Register/register[0][27] ), .QN(n2154) );
  DFFRX1 \i_MIPS/Register/register_reg[0][28]  ( .D(\i_MIPS/Register/n1136 ), 
        .CK(clk), .RN(n5707), .Q(\i_MIPS/Register/register[0][28] ), .QN(n2152) );
  DFFRX1 \i_MIPS/Register/register_reg[0][29]  ( .D(\i_MIPS/Register/n1137 ), 
        .CK(clk), .RN(n5707), .Q(\i_MIPS/Register/register[0][29] ), .QN(n2130) );
  DFFRX1 \i_MIPS/Register/register_reg[0][31]  ( .D(\i_MIPS/Register/n1139 ), 
        .CK(clk), .RN(n5708), .Q(\i_MIPS/Register/register[0][31] ), .QN(n2028) );
  DFFRX1 \i_MIPS/Register/register_reg[31][0]  ( .D(n11580), .CK(clk), .RN(
        n5622), .Q(\i_MIPS/Register/register[31][0] ), .QN(n1802) );
  DFFRX1 \i_MIPS/Register/register_reg[18][0]  ( .D(\i_MIPS/Register/n532 ), 
        .CK(clk), .RN(n5657), .Q(\i_MIPS/Register/register[18][0] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][1]  ( .D(\i_MIPS/Register/n533 ), 
        .CK(clk), .RN(n5657), .Q(\i_MIPS/Register/register[18][1] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][2]  ( .D(\i_MIPS/Register/n534 ), 
        .CK(clk), .RN(n5657), .Q(\i_MIPS/Register/register[18][2] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][3]  ( .D(\i_MIPS/Register/n535 ), 
        .CK(clk), .RN(n5657), .Q(\i_MIPS/Register/register[18][3] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][4]  ( .D(\i_MIPS/Register/n536 ), 
        .CK(clk), .RN(n5657), .Q(\i_MIPS/Register/register[18][4] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][5]  ( .D(\i_MIPS/Register/n537 ), 
        .CK(clk), .RN(n5657), .Q(\i_MIPS/Register/register[18][5] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][6]  ( .D(\i_MIPS/Register/n538 ), 
        .CK(clk), .RN(n5657), .Q(\i_MIPS/Register/register[18][6] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][7]  ( .D(\i_MIPS/Register/n539 ), 
        .CK(clk), .RN(n5658), .Q(\i_MIPS/Register/register[18][7] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][8]  ( .D(\i_MIPS/Register/n540 ), 
        .CK(clk), .RN(n5658), .Q(\i_MIPS/Register/register[18][8] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][9]  ( .D(\i_MIPS/Register/n541 ), 
        .CK(clk), .RN(n5658), .Q(\i_MIPS/Register/register[18][9] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][10]  ( .D(\i_MIPS/Register/n542 ), 
        .CK(clk), .RN(n5658), .Q(\i_MIPS/Register/register[18][10] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][11]  ( .D(\i_MIPS/Register/n543 ), 
        .CK(clk), .RN(n5658), .Q(\i_MIPS/Register/register[18][11] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][12]  ( .D(\i_MIPS/Register/n544 ), 
        .CK(clk), .RN(n5658), .Q(\i_MIPS/Register/register[18][12] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][13]  ( .D(\i_MIPS/Register/n545 ), 
        .CK(clk), .RN(n5658), .Q(\i_MIPS/Register/register[18][13] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][14]  ( .D(\i_MIPS/Register/n546 ), 
        .CK(clk), .RN(n5658), .Q(\i_MIPS/Register/register[18][14] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][15]  ( .D(\i_MIPS/Register/n547 ), 
        .CK(clk), .RN(n5658), .Q(\i_MIPS/Register/register[18][15] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][16]  ( .D(\i_MIPS/Register/n548 ), 
        .CK(clk), .RN(n5658), .Q(\i_MIPS/Register/register[18][16] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][17]  ( .D(\i_MIPS/Register/n549 ), 
        .CK(clk), .RN(n5658), .Q(\i_MIPS/Register/register[18][17] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][18]  ( .D(\i_MIPS/Register/n550 ), 
        .CK(clk), .RN(n5658), .Q(\i_MIPS/Register/register[18][18] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][19]  ( .D(\i_MIPS/Register/n551 ), 
        .CK(clk), .RN(n5659), .Q(\i_MIPS/Register/register[18][19] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][20]  ( .D(\i_MIPS/Register/n552 ), 
        .CK(clk), .RN(n5659), .Q(\i_MIPS/Register/register[18][20] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][21]  ( .D(\i_MIPS/Register/n553 ), 
        .CK(clk), .RN(n5659), .Q(\i_MIPS/Register/register[18][21] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][22]  ( .D(\i_MIPS/Register/n554 ), 
        .CK(clk), .RN(n5659), .Q(\i_MIPS/Register/register[18][22] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][23]  ( .D(\i_MIPS/Register/n555 ), 
        .CK(clk), .RN(n5659), .Q(\i_MIPS/Register/register[18][23] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][24]  ( .D(\i_MIPS/Register/n556 ), 
        .CK(clk), .RN(n5659), .Q(\i_MIPS/Register/register[18][24] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][25]  ( .D(\i_MIPS/Register/n557 ), 
        .CK(clk), .RN(n5659), .Q(\i_MIPS/Register/register[18][25] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][26]  ( .D(\i_MIPS/Register/n558 ), 
        .CK(clk), .RN(n5659), .Q(\i_MIPS/Register/register[18][26] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][27]  ( .D(\i_MIPS/Register/n559 ), 
        .CK(clk), .RN(n5659), .Q(\i_MIPS/Register/register[18][27] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][28]  ( .D(\i_MIPS/Register/n560 ), 
        .CK(clk), .RN(n5659), .Q(\i_MIPS/Register/register[18][28] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][29]  ( .D(\i_MIPS/Register/n561 ), 
        .CK(clk), .RN(n5659), .Q(\i_MIPS/Register/register[18][29] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][30]  ( .D(\i_MIPS/Register/n562 ), 
        .CK(clk), .RN(n5659), .Q(\i_MIPS/Register/register[18][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][31]  ( .D(\i_MIPS/Register/n563 ), 
        .CK(clk), .RN(n5660), .Q(\i_MIPS/Register/register[18][31] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][0]  ( .D(\i_MIPS/Register/n1044 ), 
        .CK(clk), .RN(n5700), .Q(\i_MIPS/Register/register[2][0] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][1]  ( .D(\i_MIPS/Register/n1045 ), 
        .CK(clk), .RN(n5700), .Q(\i_MIPS/Register/register[2][1] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][2]  ( .D(\i_MIPS/Register/n1046 ), 
        .CK(clk), .RN(n5700), .Q(\i_MIPS/Register/register[2][2] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][3]  ( .D(\i_MIPS/Register/n1047 ), 
        .CK(clk), .RN(n5700), .Q(\i_MIPS/Register/register[2][3] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][4]  ( .D(\i_MIPS/Register/n1048 ), 
        .CK(clk), .RN(n5700), .Q(\i_MIPS/Register/register[2][4] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][5]  ( .D(\i_MIPS/Register/n1049 ), 
        .CK(clk), .RN(n5700), .Q(\i_MIPS/Register/register[2][5] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][6]  ( .D(\i_MIPS/Register/n1050 ), 
        .CK(clk), .RN(n5700), .Q(\i_MIPS/Register/register[2][6] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][7]  ( .D(\i_MIPS/Register/n1051 ), 
        .CK(clk), .RN(n5700), .Q(\i_MIPS/Register/register[2][7] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][8]  ( .D(\i_MIPS/Register/n1052 ), 
        .CK(clk), .RN(n5700), .Q(\i_MIPS/Register/register[2][8] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][9]  ( .D(\i_MIPS/Register/n1053 ), 
        .CK(clk), .RN(n5700), .Q(\i_MIPS/Register/register[2][9] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][10]  ( .D(\i_MIPS/Register/n1054 ), 
        .CK(clk), .RN(n5700), .Q(\i_MIPS/Register/register[2][10] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][11]  ( .D(\i_MIPS/Register/n1055 ), 
        .CK(clk), .RN(n5701), .Q(\i_MIPS/Register/register[2][11] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][12]  ( .D(\i_MIPS/Register/n1056 ), 
        .CK(clk), .RN(n5701), .Q(\i_MIPS/Register/register[2][12] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][13]  ( .D(\i_MIPS/Register/n1057 ), 
        .CK(clk), .RN(n5701), .Q(\i_MIPS/Register/register[2][13] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][14]  ( .D(\i_MIPS/Register/n1058 ), 
        .CK(clk), .RN(n5701), .Q(\i_MIPS/Register/register[2][14] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][15]  ( .D(\i_MIPS/Register/n1059 ), 
        .CK(clk), .RN(n5701), .Q(\i_MIPS/Register/register[2][15] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][16]  ( .D(\i_MIPS/Register/n1060 ), 
        .CK(clk), .RN(n5701), .Q(\i_MIPS/Register/register[2][16] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][17]  ( .D(\i_MIPS/Register/n1061 ), 
        .CK(clk), .RN(n5701), .Q(\i_MIPS/Register/register[2][17] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][18]  ( .D(\i_MIPS/Register/n1062 ), 
        .CK(clk), .RN(n5701), .Q(\i_MIPS/Register/register[2][18] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][19]  ( .D(\i_MIPS/Register/n1063 ), 
        .CK(clk), .RN(n5701), .Q(\i_MIPS/Register/register[2][19] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][20]  ( .D(\i_MIPS/Register/n1064 ), 
        .CK(clk), .RN(n5701), .Q(\i_MIPS/Register/register[2][20] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][21]  ( .D(\i_MIPS/Register/n1065 ), 
        .CK(clk), .RN(n5701), .Q(\i_MIPS/Register/register[2][21] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][22]  ( .D(\i_MIPS/Register/n1066 ), 
        .CK(clk), .RN(n5701), .Q(\i_MIPS/Register/register[2][22] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][23]  ( .D(\i_MIPS/Register/n1067 ), 
        .CK(clk), .RN(n5702), .Q(\i_MIPS/Register/register[2][23] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][24]  ( .D(\i_MIPS/Register/n1068 ), 
        .CK(clk), .RN(n5702), .Q(\i_MIPS/Register/register[2][24] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][25]  ( .D(\i_MIPS/Register/n1069 ), 
        .CK(clk), .RN(n5702), .Q(\i_MIPS/Register/register[2][25] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][26]  ( .D(\i_MIPS/Register/n1070 ), 
        .CK(clk), .RN(n5702), .Q(\i_MIPS/Register/register[2][26] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][27]  ( .D(\i_MIPS/Register/n1071 ), 
        .CK(clk), .RN(n5702), .Q(\i_MIPS/Register/register[2][27] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][28]  ( .D(\i_MIPS/Register/n1072 ), 
        .CK(clk), .RN(n5702), .Q(\i_MIPS/Register/register[2][28] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][29]  ( .D(\i_MIPS/Register/n1073 ), 
        .CK(clk), .RN(n5702), .Q(\i_MIPS/Register/register[2][29] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][30]  ( .D(\i_MIPS/Register/n1074 ), 
        .CK(clk), .RN(n5702), .Q(\i_MIPS/Register/register[2][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][31]  ( .D(\i_MIPS/Register/n1075 ), 
        .CK(clk), .RN(n5702), .Q(\i_MIPS/Register/register[2][31] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][0]  ( .D(\i_MIPS/Register/n276 ), 
        .CK(clk), .RN(n5636), .Q(\i_MIPS/Register/register[26][0] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][1]  ( .D(\i_MIPS/Register/n277 ), 
        .CK(clk), .RN(n5636), .Q(\i_MIPS/Register/register[26][1] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][2]  ( .D(\i_MIPS/Register/n278 ), 
        .CK(clk), .RN(n5636), .Q(\i_MIPS/Register/register[26][2] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][4]  ( .D(\i_MIPS/Register/n280 ), 
        .CK(clk), .RN(n5636), .Q(\i_MIPS/Register/register[26][4] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][5]  ( .D(\i_MIPS/Register/n281 ), 
        .CK(clk), .RN(n5636), .Q(\i_MIPS/Register/register[26][5] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][6]  ( .D(\i_MIPS/Register/n282 ), 
        .CK(clk), .RN(n5636), .Q(\i_MIPS/Register/register[26][6] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][7]  ( .D(\i_MIPS/Register/n283 ), 
        .CK(clk), .RN(n5636), .Q(\i_MIPS/Register/register[26][7] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][8]  ( .D(\i_MIPS/Register/n284 ), 
        .CK(clk), .RN(n5636), .Q(\i_MIPS/Register/register[26][8] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][9]  ( .D(\i_MIPS/Register/n285 ), 
        .CK(clk), .RN(n5636), .Q(\i_MIPS/Register/register[26][9] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][10]  ( .D(\i_MIPS/Register/n286 ), 
        .CK(clk), .RN(n5636), .Q(\i_MIPS/Register/register[26][10] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][11]  ( .D(\i_MIPS/Register/n287 ), 
        .CK(clk), .RN(n5637), .Q(\i_MIPS/Register/register[26][11] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][12]  ( .D(\i_MIPS/Register/n288 ), 
        .CK(clk), .RN(n5637), .Q(\i_MIPS/Register/register[26][12] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][13]  ( .D(\i_MIPS/Register/n289 ), 
        .CK(clk), .RN(n5637), .Q(\i_MIPS/Register/register[26][13] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][14]  ( .D(\i_MIPS/Register/n290 ), 
        .CK(clk), .RN(n5637), .Q(\i_MIPS/Register/register[26][14] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][15]  ( .D(\i_MIPS/Register/n291 ), 
        .CK(clk), .RN(n5637), .Q(\i_MIPS/Register/register[26][15] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][17]  ( .D(\i_MIPS/Register/n293 ), 
        .CK(clk), .RN(n5637), .Q(\i_MIPS/Register/register[26][17] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][18]  ( .D(\i_MIPS/Register/n294 ), 
        .CK(clk), .RN(n5637), .Q(\i_MIPS/Register/register[26][18] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][19]  ( .D(\i_MIPS/Register/n295 ), 
        .CK(clk), .RN(n5637), .Q(\i_MIPS/Register/register[26][19] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][20]  ( .D(\i_MIPS/Register/n296 ), 
        .CK(clk), .RN(n5637), .Q(\i_MIPS/Register/register[26][20] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][21]  ( .D(\i_MIPS/Register/n297 ), 
        .CK(clk), .RN(n5637), .Q(\i_MIPS/Register/register[26][21] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][22]  ( .D(\i_MIPS/Register/n298 ), 
        .CK(clk), .RN(n5637), .Q(\i_MIPS/Register/register[26][22] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][23]  ( .D(\i_MIPS/Register/n299 ), 
        .CK(clk), .RN(n5638), .Q(\i_MIPS/Register/register[26][23] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][24]  ( .D(\i_MIPS/Register/n300 ), 
        .CK(clk), .RN(n5638), .Q(\i_MIPS/Register/register[26][24] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][25]  ( .D(\i_MIPS/Register/n301 ), 
        .CK(clk), .RN(n5638), .Q(\i_MIPS/Register/register[26][25] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][26]  ( .D(\i_MIPS/Register/n302 ), 
        .CK(clk), .RN(n5638), .Q(\i_MIPS/Register/register[26][26] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][27]  ( .D(\i_MIPS/Register/n303 ), 
        .CK(clk), .RN(n5638), .Q(\i_MIPS/Register/register[26][27] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][28]  ( .D(\i_MIPS/Register/n304 ), 
        .CK(clk), .RN(n5638), .Q(\i_MIPS/Register/register[26][28] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][29]  ( .D(\i_MIPS/Register/n305 ), 
        .CK(clk), .RN(n5638), .Q(\i_MIPS/Register/register[26][29] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][30]  ( .D(\i_MIPS/Register/n306 ), 
        .CK(clk), .RN(n5638), .Q(\i_MIPS/Register/register[26][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][31]  ( .D(\i_MIPS/Register/n307 ), 
        .CK(clk), .RN(n5638), .Q(\i_MIPS/Register/register[26][31] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][0]  ( .D(\i_MIPS/Register/n788 ), 
        .CK(clk), .RN(n5678), .Q(\i_MIPS/Register/register[10][0] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][1]  ( .D(\i_MIPS/Register/n789 ), 
        .CK(clk), .RN(n5678), .Q(\i_MIPS/Register/register[10][1] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][2]  ( .D(\i_MIPS/Register/n790 ), 
        .CK(clk), .RN(n5678), .Q(\i_MIPS/Register/register[10][2] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][4]  ( .D(\i_MIPS/Register/n792 ), 
        .CK(clk), .RN(n5679), .Q(\i_MIPS/Register/register[10][4] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][5]  ( .D(\i_MIPS/Register/n793 ), 
        .CK(clk), .RN(n5679), .Q(\i_MIPS/Register/register[10][5] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][6]  ( .D(\i_MIPS/Register/n794 ), 
        .CK(clk), .RN(n5679), .Q(\i_MIPS/Register/register[10][6] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][7]  ( .D(\i_MIPS/Register/n795 ), 
        .CK(clk), .RN(n5679), .Q(\i_MIPS/Register/register[10][7] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][8]  ( .D(\i_MIPS/Register/n796 ), 
        .CK(clk), .RN(n5679), .Q(\i_MIPS/Register/register[10][8] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][9]  ( .D(\i_MIPS/Register/n797 ), 
        .CK(clk), .RN(n5679), .Q(\i_MIPS/Register/register[10][9] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][10]  ( .D(\i_MIPS/Register/n798 ), 
        .CK(clk), .RN(n5679), .Q(\i_MIPS/Register/register[10][10] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][11]  ( .D(\i_MIPS/Register/n799 ), 
        .CK(clk), .RN(n5679), .Q(\i_MIPS/Register/register[10][11] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][12]  ( .D(\i_MIPS/Register/n800 ), 
        .CK(clk), .RN(n5679), .Q(\i_MIPS/Register/register[10][12] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][13]  ( .D(\i_MIPS/Register/n801 ), 
        .CK(clk), .RN(n5679), .Q(\i_MIPS/Register/register[10][13] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][14]  ( .D(\i_MIPS/Register/n802 ), 
        .CK(clk), .RN(n5679), .Q(\i_MIPS/Register/register[10][14] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][15]  ( .D(\i_MIPS/Register/n803 ), 
        .CK(clk), .RN(n5680), .Q(\i_MIPS/Register/register[10][15] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][16]  ( .D(\i_MIPS/Register/n804 ), 
        .CK(clk), .RN(n5680), .Q(\i_MIPS/Register/register[10][16] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][17]  ( .D(\i_MIPS/Register/n805 ), 
        .CK(clk), .RN(n5680), .Q(\i_MIPS/Register/register[10][17] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][18]  ( .D(\i_MIPS/Register/n806 ), 
        .CK(clk), .RN(n5680), .Q(\i_MIPS/Register/register[10][18] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][19]  ( .D(\i_MIPS/Register/n807 ), 
        .CK(clk), .RN(n5680), .Q(\i_MIPS/Register/register[10][19] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][20]  ( .D(\i_MIPS/Register/n808 ), 
        .CK(clk), .RN(n5680), .Q(\i_MIPS/Register/register[10][20] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][21]  ( .D(\i_MIPS/Register/n809 ), 
        .CK(clk), .RN(n5680), .Q(\i_MIPS/Register/register[10][21] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][22]  ( .D(\i_MIPS/Register/n810 ), 
        .CK(clk), .RN(n5680), .Q(\i_MIPS/Register/register[10][22] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][23]  ( .D(\i_MIPS/Register/n811 ), 
        .CK(clk), .RN(n5680), .Q(\i_MIPS/Register/register[10][23] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][24]  ( .D(\i_MIPS/Register/n812 ), 
        .CK(clk), .RN(n5680), .Q(\i_MIPS/Register/register[10][24] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][25]  ( .D(\i_MIPS/Register/n813 ), 
        .CK(clk), .RN(n5680), .Q(\i_MIPS/Register/register[10][25] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][26]  ( .D(\i_MIPS/Register/n814 ), 
        .CK(clk), .RN(n5680), .Q(\i_MIPS/Register/register[10][26] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][27]  ( .D(\i_MIPS/Register/n815 ), 
        .CK(clk), .RN(n5681), .Q(\i_MIPS/Register/register[10][27] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][28]  ( .D(\i_MIPS/Register/n816 ), 
        .CK(clk), .RN(n5681), .Q(\i_MIPS/Register/register[10][28] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][29]  ( .D(\i_MIPS/Register/n817 ), 
        .CK(clk), .RN(n5681), .Q(\i_MIPS/Register/register[10][29] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][30]  ( .D(\i_MIPS/Register/n818 ), 
        .CK(clk), .RN(n5681), .Q(\i_MIPS/Register/register[10][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][31]  ( .D(\i_MIPS/Register/n819 ), 
        .CK(clk), .RN(n5681), .Q(\i_MIPS/Register/register[10][31] ) );
  DFFRX1 \i_MIPS/Register/register_reg[31][1]  ( .D(n11579), .CK(clk), .RN(
        n5622), .QN(n183) );
  DFFRX1 \i_MIPS/Register/register_reg[31][19]  ( .D(n11561), .CK(clk), .RN(
        n5624), .QN(n184) );
  DFFRX1 \i_MIPS/Register/register_reg[31][30]  ( .D(n11550), .CK(clk), .RN(
        n5625), .QN(n228) );
  DFFRX1 \i_MIPS/ID_EX_reg[0]  ( .D(\i_MIPS/n528 ), .CK(clk), .RN(n5616), .Q(
        \i_MIPS/ID_EX_0 ), .QN(\i_MIPS/n372 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[72]  ( .D(\i_MIPS/n375 ), .CK(clk), .RN(n5601), .Q(
        \i_MIPS/ID_EX[72] ), .QN(\i_MIPS/n247 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[69]  ( .D(\i_MIPS/n381 ), .CK(clk), .RN(n5602), .Q(
        \i_MIPS/ID_EX[69] ), .QN(\i_MIPS/n253 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[68]  ( .D(\i_MIPS/n383 ), .CK(clk), .RN(n5602), .Q(
        \i_MIPS/ID_EX[68] ), .QN(\i_MIPS/n255 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[67]  ( .D(\i_MIPS/n385 ), .CK(clk), .RN(n5602), .Q(
        n3503), .QN(\i_MIPS/n257 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[70]  ( .D(\i_MIPS/n379 ), .CK(clk), .RN(n5601), .Q(
        \i_MIPS/ID_EX[70] ), .QN(\i_MIPS/n251 ) );
  DFFRX1 \D_cache/cache_reg[0][154]  ( .D(\D_cache/n564 ), .CK(clk), .RN(n5810), .Q(\D_cache/cache[0][154] ), .QN(n2352) );
  DFFRX1 \D_cache/cache_reg[1][154]  ( .D(\D_cache/n563 ), .CK(clk), .RN(n5810), .Q(\D_cache/cache[1][154] ), .QN(n850) );
  DFFRX1 \D_cache/cache_reg[2][154]  ( .D(\D_cache/n562 ), .CK(clk), .RN(n5810), .Q(\D_cache/cache[2][154] ), .QN(n2353) );
  DFFRX1 \D_cache/cache_reg[3][154]  ( .D(\D_cache/n561 ), .CK(clk), .RN(n5811), .Q(\D_cache/cache[3][154] ), .QN(n851) );
  DFFRX1 \D_cache/cache_reg[4][154]  ( .D(\D_cache/n560 ), .CK(clk), .RN(n5811), .Q(\D_cache/cache[4][154] ), .QN(n2354) );
  DFFRX1 \D_cache/cache_reg[5][154]  ( .D(\D_cache/n559 ), .CK(clk), .RN(n5811), .Q(\D_cache/cache[5][154] ), .QN(n852) );
  DFFRX1 \D_cache/cache_reg[6][154]  ( .D(\D_cache/n558 ), .CK(clk), .RN(n5811), .Q(\D_cache/cache[6][154] ), .QN(n2355) );
  DFFRX1 \D_cache/cache_reg[7][154]  ( .D(\D_cache/n557 ), .CK(clk), .RN(n5811), .Q(\D_cache/cache[7][154] ), .QN(n853) );
  DFFRX1 \i_MIPS/Register/register_reg[29][1]  ( .D(\i_MIPS/Register/n181 ), 
        .CK(clk), .RN(n5628), .Q(\i_MIPS/Register/register[29][1] ), .QN(n251)
         );
  DFFRX1 \i_MIPS/Register/register_reg[29][19]  ( .D(\i_MIPS/Register/n199 ), 
        .CK(clk), .RN(n5629), .Q(\i_MIPS/Register/register[29][19] ), .QN(n289) );
  DFFRX1 \i_MIPS/Register/register_reg[29][30]  ( .D(\i_MIPS/Register/n210 ), 
        .CK(clk), .RN(n5630), .Q(\i_MIPS/Register/register[29][30] ), .QN(n197) );
  DFFRX1 \i_MIPS/Register/register_reg[27][1]  ( .D(\i_MIPS/Register/n245 ), 
        .CK(clk), .RN(n5633), .Q(\i_MIPS/Register/register[27][1] ), .QN(n248)
         );
  DFFRX1 \i_MIPS/Register/register_reg[27][19]  ( .D(\i_MIPS/Register/n263 ), 
        .CK(clk), .RN(n5635), .Q(\i_MIPS/Register/register[27][19] ), .QN(n295) );
  DFFRX1 \i_MIPS/Register/register_reg[27][30]  ( .D(\i_MIPS/Register/n274 ), 
        .CK(clk), .RN(n5635), .Q(\i_MIPS/Register/register[27][30] ), .QN(n185) );
  DFFRX1 \i_MIPS/Register/register_reg[25][1]  ( .D(\i_MIPS/Register/n309 ), 
        .CK(clk), .RN(n5638), .Q(\i_MIPS/Register/register[25][1] ), .QN(n246)
         );
  DFFRX1 \i_MIPS/Register/register_reg[25][19]  ( .D(\i_MIPS/Register/n327 ), 
        .CK(clk), .RN(n5640), .Q(\i_MIPS/Register/register[25][19] ), .QN(n234) );
  DFFRX1 \i_MIPS/Register/register_reg[25][30]  ( .D(\i_MIPS/Register/n338 ), 
        .CK(clk), .RN(n5641), .Q(\i_MIPS/Register/register[25][30] ), .QN(n200) );
  DFFRX1 \i_MIPS/Register/register_reg[23][1]  ( .D(\i_MIPS/Register/n373 ), 
        .CK(clk), .RN(n5644), .Q(\i_MIPS/Register/register[23][1] ), .QN(n202)
         );
  DFFRX1 \i_MIPS/Register/register_reg[23][19]  ( .D(\i_MIPS/Register/n391 ), 
        .CK(clk), .RN(n5645), .Q(\i_MIPS/Register/register[23][19] ), .QN(n203) );
  DFFRX1 \i_MIPS/Register/register_reg[23][30]  ( .D(\i_MIPS/Register/n402 ), 
        .CK(clk), .RN(n5646), .Q(\i_MIPS/Register/register[23][30] ), .QN(n302) );
  DFFRX1 \i_MIPS/Register/register_reg[21][1]  ( .D(\i_MIPS/Register/n437 ), 
        .CK(clk), .RN(n5649), .Q(\i_MIPS/Register/register[21][1] ), .QN(n304)
         );
  DFFRX1 \i_MIPS/Register/register_reg[21][19]  ( .D(\i_MIPS/Register/n455 ), 
        .CK(clk), .RN(n5651), .Q(\i_MIPS/Register/register[21][19] ), .QN(
        n1859) );
  DFFRX1 \i_MIPS/Register/register_reg[21][30]  ( .D(\i_MIPS/Register/n466 ), 
        .CK(clk), .RN(n5651), .Q(\i_MIPS/Register/register[21][30] ), .QN(n303) );
  DFFRX1 \i_MIPS/Register/register_reg[19][1]  ( .D(\i_MIPS/Register/n501 ), 
        .CK(clk), .RN(n5654), .Q(\i_MIPS/Register/register[19][1] ), .QN(n307)
         );
  DFFRX1 \i_MIPS/Register/register_reg[19][19]  ( .D(\i_MIPS/Register/n519 ), 
        .CK(clk), .RN(n5656), .Q(\i_MIPS/Register/register[19][19] ), .QN(
        n1867) );
  DFFRX1 \i_MIPS/Register/register_reg[19][30]  ( .D(\i_MIPS/Register/n530 ), 
        .CK(clk), .RN(n5657), .Q(\i_MIPS/Register/register[19][30] ), .QN(n201) );
  DFFRX1 \i_MIPS/Register/register_reg[17][1]  ( .D(\i_MIPS/Register/n565 ), 
        .CK(clk), .RN(n5660), .Q(\i_MIPS/Register/register[17][1] ), .QN(n1874) );
  DFFRX1 \i_MIPS/Register/register_reg[17][19]  ( .D(\i_MIPS/Register/n583 ), 
        .CK(clk), .RN(n5661), .Q(\i_MIPS/Register/register[17][19] ), .QN(
        n1832) );
  DFFRX1 \i_MIPS/Register/register_reg[17][30]  ( .D(\i_MIPS/Register/n594 ), 
        .CK(clk), .RN(n5662), .Q(\i_MIPS/Register/register[17][30] ), .QN(n252) );
  DFFRX1 \i_MIPS/Register/register_reg[15][19]  ( .D(\i_MIPS/Register/n647 ), 
        .CK(clk), .RN(n5667), .Q(\i_MIPS/Register/register[15][19] ), .QN(n199) );
  DFFRX1 \i_MIPS/Register/register_reg[15][30]  ( .D(\i_MIPS/Register/n658 ), 
        .CK(clk), .RN(n5667), .Q(\i_MIPS/Register/register[15][30] ), .QN(n300) );
  DFFRX1 \i_MIPS/Register/register_reg[13][1]  ( .D(\i_MIPS/Register/n693 ), 
        .CK(clk), .RN(n5670), .Q(\i_MIPS/Register/register[13][1] ), .QN(n294)
         );
  DFFRX1 \i_MIPS/Register/register_reg[13][19]  ( .D(\i_MIPS/Register/n711 ), 
        .CK(clk), .RN(n5672), .Q(\i_MIPS/Register/register[13][19] ), .QN(n236) );
  DFFRX1 \i_MIPS/Register/register_reg[13][30]  ( .D(\i_MIPS/Register/n722 ), 
        .CK(clk), .RN(n5673), .Q(\i_MIPS/Register/register[13][30] ), .QN(n250) );
  DFFRX1 \i_MIPS/Register/register_reg[11][1]  ( .D(\i_MIPS/Register/n757 ), 
        .CK(clk), .RN(n5676), .Q(\i_MIPS/Register/register[11][1] ), .QN(n293)
         );
  DFFRX1 \i_MIPS/Register/register_reg[11][19]  ( .D(\i_MIPS/Register/n775 ), 
        .CK(clk), .RN(n5677), .Q(\i_MIPS/Register/register[11][19] ), .QN(n290) );
  DFFRX1 \i_MIPS/Register/register_reg[11][30]  ( .D(\i_MIPS/Register/n786 ), 
        .CK(clk), .RN(n5678), .Q(\i_MIPS/Register/register[11][30] ), .QN(n301) );
  DFFRX1 \i_MIPS/Register/register_reg[9][1]  ( .D(\i_MIPS/Register/n821 ), 
        .CK(clk), .RN(n5681), .Q(\i_MIPS/Register/register[9][1] ), .QN(n247)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][19]  ( .D(\i_MIPS/Register/n839 ), 
        .CK(clk), .RN(n5683), .Q(\i_MIPS/Register/register[9][19] ), .QN(n235)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][30]  ( .D(\i_MIPS/Register/n850 ), 
        .CK(clk), .RN(n5683), .Q(\i_MIPS/Register/register[9][30] ), .QN(n249)
         );
  DFFRX1 \i_MIPS/Register/register_reg[7][1]  ( .D(\i_MIPS/Register/n885 ), 
        .CK(clk), .RN(n5686), .Q(\i_MIPS/Register/register[7][1] ), .QN(n305)
         );
  DFFRX1 \i_MIPS/Register/register_reg[7][19]  ( .D(\i_MIPS/Register/n903 ), 
        .CK(clk), .RN(n5688), .Q(\i_MIPS/Register/register[7][19] ), .QN(n306)
         );
  DFFRX1 \i_MIPS/Register/register_reg[7][30]  ( .D(\i_MIPS/Register/n914 ), 
        .CK(clk), .RN(n5689), .Q(\i_MIPS/Register/register[7][30] ), .QN(n1863) );
  DFFRX1 \i_MIPS/Register/register_reg[5][1]  ( .D(\i_MIPS/Register/n949 ), 
        .CK(clk), .RN(n5692), .Q(\i_MIPS/Register/register[5][1] ), .QN(n1866)
         );
  DFFRX1 \i_MIPS/Register/register_reg[5][19]  ( .D(\i_MIPS/Register/n967 ), 
        .CK(clk), .RN(n5693), .Q(\i_MIPS/Register/register[5][19] ), .QN(n1861) );
  DFFRX1 \i_MIPS/Register/register_reg[5][30]  ( .D(\i_MIPS/Register/n978 ), 
        .CK(clk), .RN(n5694), .Q(\i_MIPS/Register/register[5][30] ), .QN(n1865) );
  DFFRX1 \i_MIPS/Register/register_reg[3][1]  ( .D(\i_MIPS/Register/n1013 ), 
        .CK(clk), .RN(n5697), .Q(\i_MIPS/Register/register[3][1] ), .QN(n1873)
         );
  DFFRX1 \i_MIPS/Register/register_reg[3][19]  ( .D(\i_MIPS/Register/n1031 ), 
        .CK(clk), .RN(n5699), .Q(\i_MIPS/Register/register[3][19] ), .QN(n1860) );
  DFFRX1 \i_MIPS/Register/register_reg[3][30]  ( .D(\i_MIPS/Register/n1042 ), 
        .CK(clk), .RN(n5699), .Q(\i_MIPS/Register/register[3][30] ), .QN(n1864) );
  DFFRX1 \i_MIPS/Register/register_reg[1][1]  ( .D(\i_MIPS/Register/n1077 ), 
        .CK(clk), .RN(n5702), .Q(\i_MIPS/Register/register[1][1] ), .QN(n1875)
         );
  DFFRX1 \i_MIPS/Register/register_reg[1][19]  ( .D(\i_MIPS/Register/n1095 ), 
        .CK(clk), .RN(n5704), .Q(\i_MIPS/Register/register[1][19] ), .QN(n1833) );
  DFFRX1 \i_MIPS/Register/register_reg[1][30]  ( .D(\i_MIPS/Register/n1106 ), 
        .CK(clk), .RN(n5705), .Q(\i_MIPS/Register/register[1][30] ), .QN(n1868) );
  DFFRX1 \i_MIPS/Register/register_reg[31][2]  ( .D(n11578), .CK(clk), .RN(
        n5622), .Q(\i_MIPS/Register/register[31][2] ), .QN(n196) );
  DFFRX1 \i_MIPS/Register/register_reg[31][3]  ( .D(n11577), .CK(clk), .RN(
        n5623), .Q(\i_MIPS/Register/register[31][3] ), .QN(n243) );
  DFFRX1 \i_MIPS/Register/register_reg[31][4]  ( .D(n11576), .CK(clk), .RN(
        n5623), .Q(\i_MIPS/Register/register[31][4] ), .QN(n230) );
  DFFRX1 \i_MIPS/Register/register_reg[31][5]  ( .D(n11575), .CK(clk), .RN(
        n5623), .Q(\i_MIPS/Register/register[31][5] ), .QN(n195) );
  DFFRX1 \i_MIPS/Register/register_reg[31][6]  ( .D(n11574), .CK(clk), .RN(
        n5623), .Q(\i_MIPS/Register/register[31][6] ), .QN(n191) );
  DFFRX1 \i_MIPS/Register/register_reg[31][7]  ( .D(n11573), .CK(clk), .RN(
        n5623), .Q(\i_MIPS/Register/register[31][7] ), .QN(n238) );
  DFFRX1 \i_MIPS/Register/register_reg[31][10]  ( .D(n11570), .CK(clk), .RN(
        n5623), .Q(\i_MIPS/Register/register[31][10] ), .QN(n187) );
  DFFRX1 \i_MIPS/Register/register_reg[31][11]  ( .D(n11569), .CK(clk), .RN(
        n5623), .Q(\i_MIPS/Register/register[31][11] ), .QN(n233) );
  DFFRX1 \i_MIPS/Register/register_reg[31][13]  ( .D(n11567), .CK(clk), .RN(
        n5623), .Q(\i_MIPS/Register/register[31][13] ), .QN(n227) );
  DFFRX1 \i_MIPS/Register/register_reg[31][14]  ( .D(n11566), .CK(clk), .RN(
        n5623), .Q(\i_MIPS/Register/register[31][14] ), .QN(n232) );
  DFFRX1 \i_MIPS/Register/register_reg[31][16]  ( .D(n11564), .CK(clk), .RN(
        n5624), .Q(\i_MIPS/Register/register[31][16] ), .QN(n194) );
  DFFRX1 \i_MIPS/Register/register_reg[31][18]  ( .D(n11562), .CK(clk), .RN(
        n5624), .Q(\i_MIPS/Register/register[31][18] ), .QN(n192) );
  DFFRX1 \i_MIPS/Register/register_reg[31][20]  ( .D(n11560), .CK(clk), .RN(
        n5624), .Q(\i_MIPS/Register/register[31][20] ), .QN(n244) );
  DFFRX1 \i_MIPS/Register/register_reg[31][21]  ( .D(n11559), .CK(clk), .RN(
        n5624), .Q(\i_MIPS/Register/register[31][21] ), .QN(n291) );
  DFFRX1 \i_MIPS/Register/register_reg[31][22]  ( .D(n11558), .CK(clk), .RN(
        n5624), .Q(\i_MIPS/Register/register[31][22] ), .QN(n193) );
  DFFRX1 \i_MIPS/Register/register_reg[31][23]  ( .D(n11557), .CK(clk), .RN(
        n5624), .Q(\i_MIPS/Register/register[31][23] ), .QN(n241) );
  DFFRX1 \i_MIPS/Register/register_reg[31][24]  ( .D(n11556), .CK(clk), .RN(
        n5624), .Q(\i_MIPS/Register/register[31][24] ), .QN(n242) );
  DFFRX1 \i_MIPS/Register/register_reg[31][25]  ( .D(n11555), .CK(clk), .RN(
        n5624), .Q(\i_MIPS/Register/register[31][25] ), .QN(n240) );
  DFFRX1 \i_MIPS/Register/register_reg[31][26]  ( .D(n11554), .CK(clk), .RN(
        n5624), .Q(\i_MIPS/Register/register[31][26] ), .QN(n292) );
  DFFRX1 \i_MIPS/Register/register_reg[31][27]  ( .D(n11553), .CK(clk), .RN(
        n5625), .Q(\i_MIPS/Register/register[31][27] ), .QN(n188) );
  DFFRX1 \i_MIPS/Register/register_reg[31][28]  ( .D(n11552), .CK(clk), .RN(
        n5625), .Q(\i_MIPS/Register/register[31][28] ), .QN(n245) );
  DFFRX1 \i_MIPS/Register/register_reg[31][29]  ( .D(n11551), .CK(clk), .RN(
        n5625), .Q(\i_MIPS/Register/register[31][29] ), .QN(n231) );
  DFFRX1 \D_cache/cache_reg[0][0]  ( .D(\D_cache/n1795 ), .CK(clk), .RN(n5708), 
        .Q(\D_cache/cache[0][0] ), .QN(n1390) );
  DFFRX1 \D_cache/cache_reg[1][0]  ( .D(\D_cache/n1794 ), .CK(clk), .RN(n5708), 
        .Q(\D_cache/cache[1][0] ), .QN(n3003) );
  DFFRX1 \D_cache/cache_reg[2][0]  ( .D(\D_cache/n1793 ), .CK(clk), .RN(n5708), 
        .Q(\D_cache/cache[2][0] ), .QN(n1391) );
  DFFRX1 \D_cache/cache_reg[3][0]  ( .D(\D_cache/n1792 ), .CK(clk), .RN(n5708), 
        .Q(\D_cache/cache[3][0] ), .QN(n3004) );
  DFFRX1 \D_cache/cache_reg[4][0]  ( .D(\D_cache/n1791 ), .CK(clk), .RN(n5708), 
        .Q(\D_cache/cache[4][0] ), .QN(n2368) );
  DFFRX1 \D_cache/cache_reg[5][0]  ( .D(\D_cache/n1790 ), .CK(clk), .RN(n5708), 
        .Q(\D_cache/cache[5][0] ), .QN(n865) );
  DFFRX1 \D_cache/cache_reg[6][0]  ( .D(\D_cache/n1789 ), .CK(clk), .RN(n5708), 
        .Q(\D_cache/cache[6][0] ), .QN(n2858) );
  DFFRX1 \D_cache/cache_reg[7][0]  ( .D(\D_cache/n1796 ), .CK(clk), .RN(n5708), 
        .Q(\D_cache/cache[7][0] ), .QN(n849) );
  DFFRX1 \D_cache/cache_reg[0][1]  ( .D(\D_cache/n1788 ), .CK(clk), .RN(n5708), 
        .Q(\D_cache/cache[0][1] ), .QN(n1570) );
  DFFRX1 \D_cache/cache_reg[1][1]  ( .D(\D_cache/n1787 ), .CK(clk), .RN(n5708), 
        .Q(\D_cache/cache[1][1] ), .QN(n3183) );
  DFFRX1 \D_cache/cache_reg[2][1]  ( .D(\D_cache/n1786 ), .CK(clk), .RN(n5708), 
        .Q(\D_cache/cache[2][1] ), .QN(n931) );
  DFFRX1 \D_cache/cache_reg[3][1]  ( .D(\D_cache/n1785 ), .CK(clk), .RN(n5709), 
        .Q(\D_cache/cache[3][1] ), .QN(n2455) );
  DFFRX1 \D_cache/cache_reg[4][1]  ( .D(\D_cache/n1784 ), .CK(clk), .RN(n5709), 
        .Q(\D_cache/cache[4][1] ), .QN(n1571) );
  DFFRX1 \D_cache/cache_reg[5][1]  ( .D(\D_cache/n1783 ), .CK(clk), .RN(n5709), 
        .Q(\D_cache/cache[5][1] ), .QN(n3184) );
  DFFRX1 \D_cache/cache_reg[6][1]  ( .D(\D_cache/n1782 ), .CK(clk), .RN(n5709), 
        .Q(\D_cache/cache[6][1] ), .QN(n1549) );
  DFFRX1 \D_cache/cache_reg[7][1]  ( .D(\D_cache/n1781 ), .CK(clk), .RN(n5709), 
        .Q(\D_cache/cache[7][1] ), .QN(n3162) );
  DFFRX1 \D_cache/cache_reg[0][2]  ( .D(\D_cache/n1780 ), .CK(clk), .RN(n5709), 
        .Q(\D_cache/cache[0][2] ), .QN(n1424) );
  DFFRX1 \D_cache/cache_reg[1][2]  ( .D(\D_cache/n1779 ), .CK(clk), .RN(n5709), 
        .Q(\D_cache/cache[1][2] ), .QN(n3037) );
  DFFRX1 \D_cache/cache_reg[2][2]  ( .D(\D_cache/n1778 ), .CK(clk), .RN(n5709), 
        .Q(\D_cache/cache[2][2] ), .QN(n1425) );
  DFFRX1 \D_cache/cache_reg[3][2]  ( .D(\D_cache/n1777 ), .CK(clk), .RN(n5709), 
        .Q(\D_cache/cache[3][2] ), .QN(n3038) );
  DFFRX1 \D_cache/cache_reg[4][2]  ( .D(\D_cache/n1776 ), .CK(clk), .RN(n5709), 
        .Q(\D_cache/cache[4][2] ), .QN(n1426) );
  DFFRX1 \D_cache/cache_reg[5][2]  ( .D(\D_cache/n1775 ), .CK(clk), .RN(n5709), 
        .Q(\D_cache/cache[5][2] ), .QN(n3039) );
  DFFRX1 \D_cache/cache_reg[6][2]  ( .D(\D_cache/n1774 ), .CK(clk), .RN(n5709), 
        .Q(\D_cache/cache[6][2] ), .QN(n1441) );
  DFFRX1 \D_cache/cache_reg[7][2]  ( .D(\D_cache/n1773 ), .CK(clk), .RN(n5710), 
        .Q(\D_cache/cache[7][2] ), .QN(n3054) );
  DFFRX1 \D_cache/cache_reg[0][3]  ( .D(\D_cache/n1772 ), .CK(clk), .RN(n5710), 
        .Q(\D_cache/cache[0][3] ), .QN(n1385) );
  DFFRX1 \D_cache/cache_reg[1][3]  ( .D(\D_cache/n1771 ), .CK(clk), .RN(n5710), 
        .Q(\D_cache/cache[1][3] ), .QN(n2998) );
  DFFRX1 \D_cache/cache_reg[2][3]  ( .D(\D_cache/n1770 ), .CK(clk), .RN(n5710), 
        .Q(\D_cache/cache[2][3] ), .QN(n1384) );
  DFFRX1 \D_cache/cache_reg[3][3]  ( .D(\D_cache/n1769 ), .CK(clk), .RN(n5710), 
        .Q(\D_cache/cache[3][3] ), .QN(n2997) );
  DFFRX1 \D_cache/cache_reg[4][3]  ( .D(\D_cache/n1768 ), .CK(clk), .RN(n5710), 
        .Q(\D_cache/cache[4][3] ), .QN(n2852) );
  DFFRX1 \D_cache/cache_reg[5][3]  ( .D(\D_cache/n1767 ), .CK(clk), .RN(n5710), 
        .Q(\D_cache/cache[5][3] ), .QN(n846) );
  DFFRX1 \D_cache/cache_reg[6][3]  ( .D(\D_cache/n1766 ), .CK(clk), .RN(n5710), 
        .Q(\D_cache/cache[6][3] ), .QN(n2357) );
  DFFRX1 \D_cache/cache_reg[7][3]  ( .D(\D_cache/n1765 ), .CK(clk), .RN(n5710), 
        .Q(\D_cache/cache[7][3] ), .QN(n854) );
  DFFRX1 \D_cache/cache_reg[0][4]  ( .D(\D_cache/n1764 ), .CK(clk), .RN(n5710), 
        .Q(\D_cache/cache[0][4] ), .QN(n1373) );
  DFFRX1 \D_cache/cache_reg[1][4]  ( .D(\D_cache/n1763 ), .CK(clk), .RN(n5710), 
        .Q(\D_cache/cache[1][4] ), .QN(n2986) );
  DFFRX1 \D_cache/cache_reg[2][4]  ( .D(\D_cache/n1762 ), .CK(clk), .RN(n5710), 
        .Q(\D_cache/cache[2][4] ), .QN(n1372) );
  DFFRX1 \D_cache/cache_reg[3][4]  ( .D(\D_cache/n1761 ), .CK(clk), .RN(n5711), 
        .Q(\D_cache/cache[3][4] ), .QN(n2985) );
  DFFRX1 \D_cache/cache_reg[4][4]  ( .D(\D_cache/n1760 ), .CK(clk), .RN(n5711), 
        .Q(\D_cache/cache[4][4] ), .QN(n2385) );
  DFFRX1 \D_cache/cache_reg[5][4]  ( .D(\D_cache/n1759 ), .CK(clk), .RN(n5711), 
        .Q(\D_cache/cache[5][4] ), .QN(n880) );
  DFFRX1 \D_cache/cache_reg[6][4]  ( .D(\D_cache/n1758 ), .CK(clk), .RN(n5711), 
        .Q(\D_cache/cache[6][4] ), .QN(n950) );
  DFFRX1 \D_cache/cache_reg[7][4]  ( .D(\D_cache/n1757 ), .CK(clk), .RN(n5711), 
        .Q(\D_cache/cache[7][4] ), .QN(n2475) );
  DFFRX1 \D_cache/cache_reg[1][5]  ( .D(\D_cache/n1755 ), .CK(clk), .RN(n5711), 
        .Q(\D_cache/cache[1][5] ), .QN(n2978) );
  DFFRX1 \D_cache/cache_reg[2][5]  ( .D(\D_cache/n1754 ), .CK(clk), .RN(n5711), 
        .Q(\D_cache/cache[2][5] ), .QN(n1364) );
  DFFRX1 \D_cache/cache_reg[3][5]  ( .D(\D_cache/n1753 ), .CK(clk), .RN(n5711), 
        .Q(\D_cache/cache[3][5] ), .QN(n2977) );
  DFFRX1 \D_cache/cache_reg[4][5]  ( .D(\D_cache/n1752 ), .CK(clk), .RN(n5711), 
        .Q(\D_cache/cache[4][5] ), .QN(n2380) );
  DFFRX1 \D_cache/cache_reg[5][5]  ( .D(\D_cache/n1751 ), .CK(clk), .RN(n5711), 
        .Q(\D_cache/cache[5][5] ), .QN(n876) );
  DFFRX1 \D_cache/cache_reg[6][5]  ( .D(\D_cache/n1750 ), .CK(clk), .RN(n5711), 
        .Q(\D_cache/cache[6][5] ), .QN(n1483) );
  DFFRX1 \D_cache/cache_reg[7][5]  ( .D(\D_cache/n1749 ), .CK(clk), .RN(n5712), 
        .Q(\D_cache/cache[7][5] ), .QN(n3096) );
  DFFRX1 \D_cache/cache_reg[0][6]  ( .D(\D_cache/n1748 ), .CK(clk), .RN(n5712), 
        .Q(\D_cache/cache[0][6] ), .QN(n1581) );
  DFFRX1 \D_cache/cache_reg[1][6]  ( .D(\D_cache/n1747 ), .CK(clk), .RN(n5712), 
        .Q(\D_cache/cache[1][6] ), .QN(n3194) );
  DFFRX1 \D_cache/cache_reg[2][6]  ( .D(\D_cache/n1746 ), .CK(clk), .RN(n5712), 
        .Q(\D_cache/cache[2][6] ), .QN(n1400) );
  DFFRX1 \D_cache/cache_reg[3][6]  ( .D(\D_cache/n1745 ), .CK(clk), .RN(n5712), 
        .Q(\D_cache/cache[3][6] ), .QN(n3013) );
  DFFRX1 \D_cache/cache_reg[4][6]  ( .D(\D_cache/n1744 ), .CK(clk), .RN(n5712), 
        .Q(\D_cache/cache[4][6] ), .QN(n1576) );
  DFFRX1 \D_cache/cache_reg[5][6]  ( .D(\D_cache/n1743 ), .CK(clk), .RN(n5712), 
        .Q(\D_cache/cache[5][6] ), .QN(n3189) );
  DFFRX1 \D_cache/cache_reg[6][6]  ( .D(\D_cache/n1742 ), .CK(clk), .RN(n5712), 
        .Q(\D_cache/cache[6][6] ), .QN(n1401) );
  DFFRX1 \D_cache/cache_reg[7][6]  ( .D(\D_cache/n1741 ), .CK(clk), .RN(n5712), 
        .Q(\D_cache/cache[7][6] ), .QN(n3014) );
  DFFRX1 \D_cache/cache_reg[0][7]  ( .D(\D_cache/n1740 ), .CK(clk), .RN(n5712), 
        .Q(\D_cache/cache[0][7] ), .QN(n1535) );
  DFFRX1 \D_cache/cache_reg[1][7]  ( .D(\D_cache/n1739 ), .CK(clk), .RN(n5712), 
        .Q(\D_cache/cache[1][7] ), .QN(n3148) );
  DFFRX1 \D_cache/cache_reg[2][7]  ( .D(\D_cache/n1738 ), .CK(clk), .RN(n5712), 
        .Q(\D_cache/cache[2][7] ), .QN(n1394) );
  DFFRX1 \D_cache/cache_reg[3][7]  ( .D(\D_cache/n1737 ), .CK(clk), .RN(n5713), 
        .Q(\D_cache/cache[3][7] ), .QN(n3007) );
  DFFRX1 \D_cache/cache_reg[4][7]  ( .D(\D_cache/n1736 ), .CK(clk), .RN(n5713), 
        .Q(\D_cache/cache[4][7] ), .QN(n2384) );
  DFFRX1 \D_cache/cache_reg[5][7]  ( .D(\D_cache/n1735 ), .CK(clk), .RN(n5713), 
        .Q(\D_cache/cache[5][7] ), .QN(n879) );
  DFFRX1 \D_cache/cache_reg[6][7]  ( .D(\D_cache/n1734 ), .CK(clk), .RN(n5713), 
        .Q(\D_cache/cache[6][7] ), .QN(n1395) );
  DFFRX1 \D_cache/cache_reg[7][7]  ( .D(\D_cache/n1733 ), .CK(clk), .RN(n5713), 
        .Q(\D_cache/cache[7][7] ), .QN(n3008) );
  DFFRX1 \D_cache/cache_reg[0][8]  ( .D(\D_cache/n1732 ), .CK(clk), .RN(n5713), 
        .Q(\D_cache/cache[0][8] ), .QN(n1533) );
  DFFRX1 \D_cache/cache_reg[1][8]  ( .D(\D_cache/n1731 ), .CK(clk), .RN(n5713), 
        .Q(\D_cache/cache[1][8] ), .QN(n3146) );
  DFFRX1 \D_cache/cache_reg[2][8]  ( .D(\D_cache/n1730 ), .CK(clk), .RN(n5713), 
        .Q(\D_cache/cache[2][8] ), .QN(n975) );
  DFFRX1 \D_cache/cache_reg[3][8]  ( .D(\D_cache/n1729 ), .CK(clk), .RN(n5713), 
        .Q(\D_cache/cache[3][8] ), .QN(n2502) );
  DFFRX1 \D_cache/cache_reg[4][8]  ( .D(\D_cache/n1728 ), .CK(clk), .RN(n5713), 
        .Q(\D_cache/cache[4][8] ), .QN(n976) );
  DFFRX1 \D_cache/cache_reg[5][8]  ( .D(\D_cache/n1727 ), .CK(clk), .RN(n5713), 
        .Q(\D_cache/cache[5][8] ), .QN(n2503) );
  DFFRX1 \D_cache/cache_reg[6][8]  ( .D(\D_cache/n1726 ), .CK(clk), .RN(n5713), 
        .Q(\D_cache/cache[6][8] ), .QN(n1439) );
  DFFRX1 \D_cache/cache_reg[7][8]  ( .D(\D_cache/n1725 ), .CK(clk), .RN(n5714), 
        .Q(\D_cache/cache[7][8] ), .QN(n3052) );
  DFFRX1 \D_cache/cache_reg[0][9]  ( .D(\D_cache/n1724 ), .CK(clk), .RN(n5714), 
        .Q(\D_cache/cache[0][9] ), .QN(n1532) );
  DFFRX1 \D_cache/cache_reg[1][9]  ( .D(\D_cache/n1723 ), .CK(clk), .RN(n5714), 
        .Q(\D_cache/cache[1][9] ), .QN(n3145) );
  DFFRX1 \D_cache/cache_reg[2][9]  ( .D(\D_cache/n1722 ), .CK(clk), .RN(n5714), 
        .Q(\D_cache/cache[2][9] ), .QN(n967) );
  DFFRX1 \D_cache/cache_reg[3][9]  ( .D(\D_cache/n1721 ), .CK(clk), .RN(n5714), 
        .Q(\D_cache/cache[3][9] ), .QN(n2492) );
  DFFRX1 \D_cache/cache_reg[4][9]  ( .D(\D_cache/n1720 ), .CK(clk), .RN(n5714), 
        .Q(\D_cache/cache[4][9] ), .QN(n922) );
  DFFRX1 \D_cache/cache_reg[5][9]  ( .D(\D_cache/n1719 ), .CK(clk), .RN(n5714), 
        .Q(\D_cache/cache[5][9] ), .QN(n2493) );
  DFFRX1 \D_cache/cache_reg[6][9]  ( .D(\D_cache/n1718 ), .CK(clk), .RN(n5714), 
        .Q(\D_cache/cache[6][9] ), .QN(n1433) );
  DFFRX1 \D_cache/cache_reg[7][9]  ( .D(\D_cache/n1717 ), .CK(clk), .RN(n5714), 
        .Q(\D_cache/cache[7][9] ), .QN(n3046) );
  DFFRX1 \D_cache/cache_reg[0][10]  ( .D(\D_cache/n1716 ), .CK(clk), .RN(n5714), .Q(\D_cache/cache[0][10] ), .QN(n2375) );
  DFFRX1 \D_cache/cache_reg[1][10]  ( .D(\D_cache/n1715 ), .CK(clk), .RN(n5714), .Q(\D_cache/cache[1][10] ), .QN(n871) );
  DFFRX1 \D_cache/cache_reg[2][10]  ( .D(\D_cache/n1714 ), .CK(clk), .RN(n5714), .Q(\D_cache/cache[2][10] ), .QN(n939) );
  DFFRX1 \D_cache/cache_reg[3][10]  ( .D(\D_cache/n1713 ), .CK(clk), .RN(n5715), .Q(\D_cache/cache[3][10] ), .QN(n2464) );
  DFFRX1 \D_cache/cache_reg[4][10]  ( .D(\D_cache/n1712 ), .CK(clk), .RN(n5715), .Q(\D_cache/cache[4][10] ), .QN(n2392) );
  DFFRX1 \D_cache/cache_reg[5][10]  ( .D(\D_cache/n1711 ), .CK(clk), .RN(n5715), .Q(\D_cache/cache[5][10] ), .QN(n887) );
  DFFRX1 \D_cache/cache_reg[6][10]  ( .D(\D_cache/n1710 ), .CK(clk), .RN(n5715), .Q(\D_cache/cache[6][10] ), .QN(n1487) );
  DFFRX1 \D_cache/cache_reg[7][10]  ( .D(\D_cache/n1709 ), .CK(clk), .RN(n5715), .Q(\D_cache/cache[7][10] ), .QN(n3100) );
  DFFRX1 \D_cache/cache_reg[0][11]  ( .D(\D_cache/n1708 ), .CK(clk), .RN(n5715), .Q(\D_cache/cache[0][11] ), .QN(n2374) );
  DFFRX1 \D_cache/cache_reg[1][11]  ( .D(\D_cache/n1707 ), .CK(clk), .RN(n5715), .Q(\D_cache/cache[1][11] ), .QN(n870) );
  DFFRX1 \D_cache/cache_reg[2][11]  ( .D(\D_cache/n1706 ), .CK(clk), .RN(n5715), .Q(\D_cache/cache[2][11] ), .QN(n1497) );
  DFFRX1 \D_cache/cache_reg[3][11]  ( .D(\D_cache/n1705 ), .CK(clk), .RN(n5715), .Q(\D_cache/cache[3][11] ), .QN(n3110) );
  DFFRX1 \D_cache/cache_reg[4][11]  ( .D(\D_cache/n1704 ), .CK(clk), .RN(n5715), .Q(\D_cache/cache[4][11] ), .QN(n2391) );
  DFFRX1 \D_cache/cache_reg[5][11]  ( .D(\D_cache/n1703 ), .CK(clk), .RN(n5715), .Q(\D_cache/cache[5][11] ), .QN(n886) );
  DFFRX1 \D_cache/cache_reg[6][11]  ( .D(\D_cache/n1702 ), .CK(clk), .RN(n5715), .Q(\D_cache/cache[6][11] ), .QN(n1490) );
  DFFRX1 \D_cache/cache_reg[7][11]  ( .D(\D_cache/n1701 ), .CK(clk), .RN(n5716), .Q(\D_cache/cache[7][11] ), .QN(n3103) );
  DFFRX1 \D_cache/cache_reg[0][12]  ( .D(\D_cache/n1700 ), .CK(clk), .RN(n5716), .Q(\D_cache/cache[0][12] ), .QN(n1538) );
  DFFRX1 \D_cache/cache_reg[1][12]  ( .D(\D_cache/n1699 ), .CK(clk), .RN(n5716), .Q(\D_cache/cache[1][12] ), .QN(n3151) );
  DFFRX1 \D_cache/cache_reg[2][12]  ( .D(\D_cache/n1698 ), .CK(clk), .RN(n5716), .Q(\D_cache/cache[2][12] ), .QN(n1499) );
  DFFRX1 \D_cache/cache_reg[3][12]  ( .D(\D_cache/n1697 ), .CK(clk), .RN(n5716), .Q(\D_cache/cache[3][12] ), .QN(n3112) );
  DFFRX1 \D_cache/cache_reg[4][12]  ( .D(\D_cache/n1696 ), .CK(clk), .RN(n5716), .Q(\D_cache/cache[4][12] ), .QN(n2364) );
  DFFRX1 \D_cache/cache_reg[5][12]  ( .D(\D_cache/n1695 ), .CK(clk), .RN(n5716), .Q(\D_cache/cache[5][12] ), .QN(n861) );
  DFFRX1 \D_cache/cache_reg[6][12]  ( .D(\D_cache/n1694 ), .CK(clk), .RN(n5716), .Q(\D_cache/cache[6][12] ), .QN(n1500) );
  DFFRX1 \D_cache/cache_reg[7][12]  ( .D(\D_cache/n1693 ), .CK(clk), .RN(n5716), .Q(\D_cache/cache[7][12] ), .QN(n3113) );
  DFFRX1 \D_cache/cache_reg[0][13]  ( .D(\D_cache/n1692 ), .CK(clk), .RN(n5716), .Q(\D_cache/cache[0][13] ), .QN(n1241) );
  DFFRX1 \D_cache/cache_reg[1][13]  ( .D(\D_cache/n1691 ), .CK(clk), .RN(n5716), .Q(\D_cache/cache[1][13] ), .QN(n2846) );
  DFFRX1 \D_cache/cache_reg[2][13]  ( .D(\D_cache/n1690 ), .CK(clk), .RN(n5716), .Q(\D_cache/cache[2][13] ), .QN(n1402) );
  DFFRX1 \D_cache/cache_reg[3][13]  ( .D(\D_cache/n1689 ), .CK(clk), .RN(n5717), .Q(\D_cache/cache[3][13] ), .QN(n3015) );
  DFFRX1 \D_cache/cache_reg[4][13]  ( .D(\D_cache/n1688 ), .CK(clk), .RN(n5717), .Q(\D_cache/cache[4][13] ), .QN(n2362) );
  DFFRX1 \D_cache/cache_reg[5][13]  ( .D(\D_cache/n1687 ), .CK(clk), .RN(n5717), .Q(\D_cache/cache[5][13] ), .QN(n859) );
  DFFRX1 \D_cache/cache_reg[6][13]  ( .D(\D_cache/n1686 ), .CK(clk), .RN(n5717), .Q(\D_cache/cache[6][13] ), .QN(n1403) );
  DFFRX1 \D_cache/cache_reg[7][13]  ( .D(\D_cache/n1685 ), .CK(clk), .RN(n5717), .Q(\D_cache/cache[7][13] ), .QN(n3016) );
  DFFRX1 \D_cache/cache_reg[0][14]  ( .D(\D_cache/n1684 ), .CK(clk), .RN(n5717), .Q(\D_cache/cache[0][14] ), .QN(n804) );
  DFFRX1 \D_cache/cache_reg[1][14]  ( .D(\D_cache/n1683 ), .CK(clk), .RN(n5717), .Q(\D_cache/cache[1][14] ), .QN(n2351) );
  DFFRX1 \D_cache/cache_reg[2][14]  ( .D(\D_cache/n1682 ), .CK(clk), .RN(n5717), .Q(\D_cache/cache[2][14] ), .QN(n974) );
  DFFRX1 \D_cache/cache_reg[3][14]  ( .D(\D_cache/n1681 ), .CK(clk), .RN(n5717), .Q(\D_cache/cache[3][14] ), .QN(n2501) );
  DFFRX1 \D_cache/cache_reg[4][14]  ( .D(\D_cache/n1680 ), .CK(clk), .RN(n5717), .Q(\D_cache/cache[4][14] ), .QN(n2398) );
  DFFRX1 \D_cache/cache_reg[5][14]  ( .D(\D_cache/n1679 ), .CK(clk), .RN(n5717), .Q(\D_cache/cache[5][14] ), .QN(n893) );
  DFFRX1 \D_cache/cache_reg[6][14]  ( .D(\D_cache/n1678 ), .CK(clk), .RN(n5717), .Q(\D_cache/cache[6][14] ), .QN(n1438) );
  DFFRX1 \D_cache/cache_reg[7][14]  ( .D(\D_cache/n1677 ), .CK(clk), .RN(n5718), .Q(\D_cache/cache[7][14] ), .QN(n3051) );
  DFFRX1 \D_cache/cache_reg[0][15]  ( .D(\D_cache/n1676 ), .CK(clk), .RN(n5718), .Q(\D_cache/cache[0][15] ), .QN(n2370) );
  DFFRX1 \D_cache/cache_reg[1][15]  ( .D(\D_cache/n1675 ), .CK(clk), .RN(n5718), .Q(\D_cache/cache[1][15] ), .QN(n866) );
  DFFRX1 \D_cache/cache_reg[2][15]  ( .D(\D_cache/n1674 ), .CK(clk), .RN(n5718), .Q(\D_cache/cache[2][15] ), .QN(n1436) );
  DFFRX1 \D_cache/cache_reg[3][15]  ( .D(\D_cache/n1673 ), .CK(clk), .RN(n5718), .Q(\D_cache/cache[3][15] ), .QN(n3049) );
  DFFRX1 \D_cache/cache_reg[4][15]  ( .D(\D_cache/n1672 ), .CK(clk), .RN(n5718), .Q(\D_cache/cache[4][15] ), .QN(n2389) );
  DFFRX1 \D_cache/cache_reg[5][15]  ( .D(\D_cache/n1671 ), .CK(clk), .RN(n5718), .Q(\D_cache/cache[5][15] ), .QN(n884) );
  DFFRX1 \D_cache/cache_reg[6][15]  ( .D(\D_cache/n1670 ), .CK(clk), .RN(n5718), .Q(\D_cache/cache[6][15] ), .QN(n1437) );
  DFFRX1 \D_cache/cache_reg[7][15]  ( .D(\D_cache/n1669 ), .CK(clk), .RN(n5718), .Q(\D_cache/cache[7][15] ), .QN(n3050) );
  DFFRX1 \D_cache/cache_reg[0][16]  ( .D(\D_cache/n1668 ), .CK(clk), .RN(n5718), .Q(\D_cache/cache[0][16] ), .QN(n973) );
  DFFRX1 \D_cache/cache_reg[1][16]  ( .D(\D_cache/n1667 ), .CK(clk), .RN(n5718), .Q(\D_cache/cache[1][16] ), .QN(n2500) );
  DFFRX1 \D_cache/cache_reg[2][16]  ( .D(\D_cache/n1666 ), .CK(clk), .RN(n5718), .Q(\D_cache/cache[2][16] ), .QN(n1435) );
  DFFRX1 \D_cache/cache_reg[3][16]  ( .D(\D_cache/n1665 ), .CK(clk), .RN(n5719), .Q(\D_cache/cache[3][16] ), .QN(n3048) );
  DFFRX1 \D_cache/cache_reg[4][16]  ( .D(\D_cache/n1664 ), .CK(clk), .RN(n5719), .Q(\D_cache/cache[4][16] ), .QN(n972) );
  DFFRX1 \D_cache/cache_reg[5][16]  ( .D(\D_cache/n1663 ), .CK(clk), .RN(n5719), .Q(\D_cache/cache[5][16] ), .QN(n2499) );
  DFFRX1 \D_cache/cache_reg[6][16]  ( .D(\D_cache/n1662 ), .CK(clk), .RN(n5719), .Q(\D_cache/cache[6][16] ), .QN(n1508) );
  DFFRX1 \D_cache/cache_reg[7][16]  ( .D(\D_cache/n1661 ), .CK(clk), .RN(n5719), .Q(\D_cache/cache[7][16] ), .QN(n3121) );
  DFFRX1 \D_cache/cache_reg[0][17]  ( .D(\D_cache/n1660 ), .CK(clk), .RN(n5719), .Q(\D_cache/cache[0][17] ), .QN(n1579) );
  DFFRX1 \D_cache/cache_reg[1][17]  ( .D(\D_cache/n1659 ), .CK(clk), .RN(n5719), .Q(\D_cache/cache[1][17] ), .QN(n3192) );
  DFFRX1 \D_cache/cache_reg[2][17]  ( .D(\D_cache/n1658 ), .CK(clk), .RN(n5719), .Q(\D_cache/cache[2][17] ), .QN(n2833) );
  DFFRX1 \D_cache/cache_reg[3][17]  ( .D(\D_cache/n1657 ), .CK(clk), .RN(n5719), .Q(\D_cache/cache[3][17] ), .QN(n841) );
  DFFRX1 \D_cache/cache_reg[4][17]  ( .D(\D_cache/n1656 ), .CK(clk), .RN(n5719), .Q(\D_cache/cache[4][17] ), .QN(n1578) );
  DFFRX1 \D_cache/cache_reg[5][17]  ( .D(\D_cache/n1655 ), .CK(clk), .RN(n5719), .Q(\D_cache/cache[5][17] ), .QN(n3191) );
  DFFRX1 \D_cache/cache_reg[6][17]  ( .D(\D_cache/n1654 ), .CK(clk), .RN(n5719), .Q(\D_cache/cache[6][17] ), .QN(n2834) );
  DFFRX1 \D_cache/cache_reg[7][17]  ( .D(\D_cache/n1653 ), .CK(clk), .RN(n5720), .Q(\D_cache/cache[7][17] ), .QN(n842) );
  DFFRX1 \D_cache/cache_reg[0][18]  ( .D(\D_cache/n1652 ), .CK(clk), .RN(n5720), .Q(\D_cache/cache[0][18] ), .QN(n927) );
  DFFRX1 \D_cache/cache_reg[1][18]  ( .D(\D_cache/n1651 ), .CK(clk), .RN(n5720), .Q(\D_cache/cache[1][18] ), .QN(n2451) );
  DFFRX1 \D_cache/cache_reg[2][18]  ( .D(\D_cache/n1650 ), .CK(clk), .RN(n5720), .Q(\D_cache/cache[2][18] ), .QN(n929) );
  DFFRX1 \D_cache/cache_reg[3][18]  ( .D(\D_cache/n1649 ), .CK(clk), .RN(n5720), .Q(\D_cache/cache[3][18] ), .QN(n2453) );
  DFFRX1 \D_cache/cache_reg[4][18]  ( .D(\D_cache/n1648 ), .CK(clk), .RN(n5720), .Q(\D_cache/cache[4][18] ), .QN(n1498) );
  DFFRX1 \D_cache/cache_reg[5][18]  ( .D(\D_cache/n1647 ), .CK(clk), .RN(n5720), .Q(\D_cache/cache[5][18] ), .QN(n3111) );
  DFFRX1 \D_cache/cache_reg[6][18]  ( .D(\D_cache/n1646 ), .CK(clk), .RN(n5720), .Q(\D_cache/cache[6][18] ), .QN(n2316) );
  DFFRX1 \D_cache/cache_reg[0][19]  ( .D(\D_cache/n1644 ), .CK(clk), .RN(n5720), .Q(\D_cache/cache[0][19] ), .QN(n957) );
  DFFRX1 \D_cache/cache_reg[1][19]  ( .D(\D_cache/n1643 ), .CK(clk), .RN(n5720), .Q(\D_cache/cache[1][19] ), .QN(n2482) );
  DFFRX1 \D_cache/cache_reg[2][19]  ( .D(\D_cache/n1642 ), .CK(clk), .RN(n5720), .Q(\D_cache/cache[2][19] ), .QN(n956) );
  DFFRX1 \D_cache/cache_reg[3][19]  ( .D(\D_cache/n1641 ), .CK(clk), .RN(n5721), .Q(\D_cache/cache[3][19] ), .QN(n2481) );
  DFFRX1 \D_cache/cache_reg[4][19]  ( .D(\D_cache/n1640 ), .CK(clk), .RN(n5721), .Q(\D_cache/cache[4][19] ), .QN(n1572) );
  DFFRX1 \D_cache/cache_reg[5][19]  ( .D(\D_cache/n1639 ), .CK(clk), .RN(n5721), .Q(\D_cache/cache[5][19] ), .QN(n3185) );
  DFFRX1 \D_cache/cache_reg[6][19]  ( .D(\D_cache/n1638 ), .CK(clk), .RN(n5721), .Q(\D_cache/cache[6][19] ), .QN(n937) );
  DFFRX1 \D_cache/cache_reg[7][19]  ( .D(\D_cache/n1637 ), .CK(clk), .RN(n5721), .Q(\D_cache/cache[7][19] ), .QN(n2462) );
  DFFRX1 \D_cache/cache_reg[0][20]  ( .D(\D_cache/n1636 ), .CK(clk), .RN(n5721), .Q(\D_cache/cache[0][20] ), .QN(n966) );
  DFFRX1 \D_cache/cache_reg[1][20]  ( .D(\D_cache/n1635 ), .CK(clk), .RN(n5721), .Q(\D_cache/cache[1][20] ), .QN(n2491) );
  DFFRX1 \D_cache/cache_reg[2][20]  ( .D(\D_cache/n1634 ), .CK(clk), .RN(n5721), .Q(\D_cache/cache[2][20] ), .QN(n965) );
  DFFRX1 \D_cache/cache_reg[3][20]  ( .D(\D_cache/n1633 ), .CK(clk), .RN(n5721), .Q(\D_cache/cache[3][20] ), .QN(n2490) );
  DFFRX1 \D_cache/cache_reg[4][20]  ( .D(\D_cache/n1632 ), .CK(clk), .RN(n5721), .Q(\D_cache/cache[4][20] ), .QN(n1432) );
  DFFRX1 \D_cache/cache_reg[5][20]  ( .D(\D_cache/n1631 ), .CK(clk), .RN(n5721), .Q(\D_cache/cache[5][20] ), .QN(n3045) );
  DFFRX1 \D_cache/cache_reg[6][20]  ( .D(\D_cache/n1630 ), .CK(clk), .RN(n5721), .Q(\D_cache/cache[6][20] ), .QN(n1509) );
  DFFRX1 \D_cache/cache_reg[7][20]  ( .D(\D_cache/n1629 ), .CK(clk), .RN(n5722), .Q(\D_cache/cache[7][20] ), .QN(n3122) );
  DFFRX1 \D_cache/cache_reg[0][21]  ( .D(\D_cache/n1628 ), .CK(clk), .RN(n5722), .Q(\D_cache/cache[0][21] ), .QN(n1246) );
  DFFRX1 \D_cache/cache_reg[1][21]  ( .D(\D_cache/n1627 ), .CK(clk), .RN(n5722), .Q(\D_cache/cache[1][21] ), .QN(n2853) );
  DFFRX1 \D_cache/cache_reg[2][21]  ( .D(\D_cache/n1626 ), .CK(clk), .RN(n5722), .Q(\D_cache/cache[2][21] ), .QN(n2824) );
  DFFRX1 \D_cache/cache_reg[3][21]  ( .D(\D_cache/n1625 ), .CK(clk), .RN(n5722), .Q(\D_cache/cache[3][21] ), .QN(n832) );
  DFFRX1 \D_cache/cache_reg[4][21]  ( .D(\D_cache/n1624 ), .CK(clk), .RN(n5722), .Q(\D_cache/cache[4][21] ), .QN(n2825) );
  DFFRX1 \D_cache/cache_reg[5][21]  ( .D(\D_cache/n1623 ), .CK(clk), .RN(n5722), .Q(\D_cache/cache[5][21] ), .QN(n833) );
  DFFRX1 \D_cache/cache_reg[6][21]  ( .D(\D_cache/n1622 ), .CK(clk), .RN(n5722), .Q(\D_cache/cache[6][21] ), .QN(n2826) );
  DFFRX1 \D_cache/cache_reg[7][21]  ( .D(\D_cache/n1621 ), .CK(clk), .RN(n5722), .Q(\D_cache/cache[7][21] ), .QN(n834) );
  DFFRX1 \D_cache/cache_reg[0][22]  ( .D(\D_cache/n1620 ), .CK(clk), .RN(n5722), .Q(\D_cache/cache[0][22] ), .QN(n928) );
  DFFRX1 \D_cache/cache_reg[1][22]  ( .D(\D_cache/n1619 ), .CK(clk), .RN(n5722), .Q(\D_cache/cache[1][22] ), .QN(n2452) );
  DFFRX1 \D_cache/cache_reg[2][22]  ( .D(\D_cache/n1618 ), .CK(clk), .RN(n5722), .Q(\D_cache/cache[2][22] ), .QN(n1423) );
  DFFRX1 \D_cache/cache_reg[3][22]  ( .D(\D_cache/n1617 ), .CK(clk), .RN(n5723), .Q(\D_cache/cache[3][22] ), .QN(n3036) );
  DFFRX1 \D_cache/cache_reg[4][22]  ( .D(\D_cache/n1616 ), .CK(clk), .RN(n5723), .Q(\D_cache/cache[4][22] ), .QN(n2410) );
  DFFRX1 \D_cache/cache_reg[5][22]  ( .D(\D_cache/n1615 ), .CK(clk), .RN(n5723), .Q(\D_cache/cache[5][22] ), .QN(n382) );
  DFFRX1 \D_cache/cache_reg[6][22]  ( .D(\D_cache/n1614 ), .CK(clk), .RN(n5723), .Q(\D_cache/cache[6][22] ), .QN(n1448) );
  DFFRX1 \D_cache/cache_reg[7][22]  ( .D(\D_cache/n1613 ), .CK(clk), .RN(n5723), .Q(\D_cache/cache[7][22] ), .QN(n3061) );
  DFFRX1 \D_cache/cache_reg[0][23]  ( .D(\D_cache/n1612 ), .CK(clk), .RN(n5723), .Q(\D_cache/cache[0][23] ), .QN(n1464) );
  DFFRX1 \D_cache/cache_reg[1][23]  ( .D(\D_cache/n1611 ), .CK(clk), .RN(n5723), .Q(\D_cache/cache[1][23] ), .QN(n3077) );
  DFFRX1 \D_cache/cache_reg[2][23]  ( .D(\D_cache/n1610 ), .CK(clk), .RN(n5723), .Q(\D_cache/cache[2][23] ), .QN(n1427) );
  DFFRX1 \D_cache/cache_reg[3][23]  ( .D(\D_cache/n1609 ), .CK(clk), .RN(n5723), .Q(\D_cache/cache[3][23] ), .QN(n3040) );
  DFFRX1 \D_cache/cache_reg[4][23]  ( .D(\D_cache/n1608 ), .CK(clk), .RN(n5723), .Q(\D_cache/cache[4][23] ), .QN(n943) );
  DFFRX1 \D_cache/cache_reg[5][23]  ( .D(\D_cache/n1607 ), .CK(clk), .RN(n5723), .Q(\D_cache/cache[5][23] ), .QN(n2468) );
  DFFRX1 \D_cache/cache_reg[6][23]  ( .D(\D_cache/n1606 ), .CK(clk), .RN(n5723), .Q(\D_cache/cache[6][23] ), .QN(n1510) );
  DFFRX1 \D_cache/cache_reg[7][23]  ( .D(\D_cache/n1605 ), .CK(clk), .RN(n5724), .Q(\D_cache/cache[7][23] ), .QN(n3123) );
  DFFRX1 \D_cache/cache_reg[0][24]  ( .D(\D_cache/n1604 ), .CK(clk), .RN(n5724), .Q(\D_cache/cache[0][24] ), .QN(n969) );
  DFFRX1 \D_cache/cache_reg[1][24]  ( .D(\D_cache/n1603 ), .CK(clk), .RN(n5724), .Q(\D_cache/cache[1][24] ), .QN(n2495) );
  DFFRX1 \D_cache/cache_reg[2][24]  ( .D(\D_cache/n1602 ), .CK(clk), .RN(n5724), .Q(\D_cache/cache[2][24] ), .QN(n968) );
  DFFRX1 \D_cache/cache_reg[3][24]  ( .D(\D_cache/n1601 ), .CK(clk), .RN(n5724), .Q(\D_cache/cache[3][24] ), .QN(n2494) );
  DFFRX1 \D_cache/cache_reg[4][24]  ( .D(\D_cache/n1600 ), .CK(clk), .RN(n5724), .Q(\D_cache/cache[4][24] ), .QN(n2835) );
  DFFRX1 \D_cache/cache_reg[5][24]  ( .D(\D_cache/n1599 ), .CK(clk), .RN(n5724), .Q(\D_cache/cache[5][24] ), .QN(n843) );
  DFFRX1 \D_cache/cache_reg[6][24]  ( .D(\D_cache/n1598 ), .CK(clk), .RN(n5724), .Q(\D_cache/cache[6][24] ), .QN(n1493) );
  DFFRX1 \D_cache/cache_reg[7][24]  ( .D(\D_cache/n1597 ), .CK(clk), .RN(n5724), .Q(\D_cache/cache[7][24] ), .QN(n3106) );
  DFFRX1 \D_cache/cache_reg[0][25]  ( .D(\D_cache/n1596 ), .CK(clk), .RN(n5724), .Q(\D_cache/cache[0][25] ), .QN(n941) );
  DFFRX1 \D_cache/cache_reg[1][25]  ( .D(\D_cache/n1595 ), .CK(clk), .RN(n5724), .Q(\D_cache/cache[1][25] ), .QN(n2466) );
  DFFRX1 \D_cache/cache_reg[2][25]  ( .D(\D_cache/n1594 ), .CK(clk), .RN(n5724), .Q(\D_cache/cache[2][25] ), .QN(n1249) );
  DFFRX1 \D_cache/cache_reg[3][25]  ( .D(\D_cache/n1593 ), .CK(clk), .RN(n5725), .Q(\D_cache/cache[3][25] ), .QN(n2860) );
  DFFRX1 \D_cache/cache_reg[4][25]  ( .D(\D_cache/n1592 ), .CK(clk), .RN(n5725), .Q(\D_cache/cache[4][25] ), .QN(n940) );
  DFFRX1 \D_cache/cache_reg[5][25]  ( .D(\D_cache/n1591 ), .CK(clk), .RN(n5725), .Q(\D_cache/cache[5][25] ), .QN(n2465) );
  DFFRX1 \D_cache/cache_reg[6][25]  ( .D(\D_cache/n1590 ), .CK(clk), .RN(n5725), .Q(\D_cache/cache[6][25] ), .QN(n1250) );
  DFFRX1 \D_cache/cache_reg[7][25]  ( .D(\D_cache/n1589 ), .CK(clk), .RN(n5725), .Q(\D_cache/cache[7][25] ), .QN(n2861) );
  DFFRX1 \D_cache/cache_reg[0][26]  ( .D(\D_cache/n1588 ), .CK(clk), .RN(n5725), .Q(\D_cache/cache[0][26] ), .QN(n2409) );
  DFFRX1 \D_cache/cache_reg[1][26]  ( .D(\D_cache/n1587 ), .CK(clk), .RN(n5725), .Q(\D_cache/cache[1][26] ), .QN(n903) );
  DFFRX1 \D_cache/cache_reg[2][26]  ( .D(\D_cache/n1586 ), .CK(clk), .RN(n5725), .Q(\D_cache/cache[2][26] ), .QN(n920) );
  DFFRX1 \D_cache/cache_reg[3][26]  ( .D(\D_cache/n1585 ), .CK(clk), .RN(n5725), .Q(\D_cache/cache[3][26] ), .QN(n2498) );
  DFFRX1 \D_cache/cache_reg[4][26]  ( .D(\D_cache/n1584 ), .CK(clk), .RN(n5725), .Q(\D_cache/cache[4][26] ), .QN(n2836) );
  DFFRX1 \D_cache/cache_reg[5][26]  ( .D(\D_cache/n1583 ), .CK(clk), .RN(n5725), .Q(\D_cache/cache[5][26] ), .QN(n844) );
  DFFRX1 \D_cache/cache_reg[6][26]  ( .D(\D_cache/n1582 ), .CK(clk), .RN(n5725), .Q(\D_cache/cache[6][26] ), .QN(n1239) );
  DFFRX1 \D_cache/cache_reg[7][26]  ( .D(\D_cache/n1581 ), .CK(clk), .RN(n5726), .Q(\D_cache/cache[7][26] ), .QN(n2844) );
  DFFRX1 \D_cache/cache_reg[0][27]  ( .D(\D_cache/n1580 ), .CK(clk), .RN(n5726), .Q(\D_cache/cache[0][27] ), .QN(n971) );
  DFFRX1 \D_cache/cache_reg[1][27]  ( .D(\D_cache/n1579 ), .CK(clk), .RN(n5726), .Q(\D_cache/cache[1][27] ), .QN(n2497) );
  DFFRX1 \D_cache/cache_reg[2][27]  ( .D(\D_cache/n1578 ), .CK(clk), .RN(n5726), .Q(\D_cache/cache[2][27] ), .QN(n970) );
  DFFRX1 \D_cache/cache_reg[3][27]  ( .D(\D_cache/n1577 ), .CK(clk), .RN(n5726), .Q(\D_cache/cache[3][27] ), .QN(n2496) );
  DFFRX1 \D_cache/cache_reg[4][27]  ( .D(\D_cache/n1576 ), .CK(clk), .RN(n5726), .Q(\D_cache/cache[4][27] ), .QN(n1434) );
  DFFRX1 \D_cache/cache_reg[5][27]  ( .D(\D_cache/n1575 ), .CK(clk), .RN(n5726), .Q(\D_cache/cache[5][27] ), .QN(n3047) );
  DFFRX1 \D_cache/cache_reg[6][27]  ( .D(\D_cache/n1574 ), .CK(clk), .RN(n5726), .Q(\D_cache/cache[6][27] ), .QN(n2399) );
  DFFRX1 \D_cache/cache_reg[7][27]  ( .D(\D_cache/n1573 ), .CK(clk), .RN(n5726), .Q(\D_cache/cache[7][27] ), .QN(n894) );
  DFFRX1 \D_cache/cache_reg[0][28]  ( .D(\D_cache/n1572 ), .CK(clk), .RN(n5726), .Q(\D_cache/cache[0][28] ), .QN(n935) );
  DFFRX1 \D_cache/cache_reg[1][28]  ( .D(\D_cache/n1571 ), .CK(clk), .RN(n5726), .Q(\D_cache/cache[1][28] ), .QN(n2460) );
  DFFRX1 \D_cache/cache_reg[2][28]  ( .D(\D_cache/n1570 ), .CK(clk), .RN(n5726), .Q(\D_cache/cache[2][28] ), .QN(n2810) );
  DFFRX1 \D_cache/cache_reg[3][28]  ( .D(\D_cache/n1569 ), .CK(clk), .RN(n5727), .Q(\D_cache/cache[3][28] ), .QN(n818) );
  DFFRX1 \D_cache/cache_reg[4][28]  ( .D(\D_cache/n1568 ), .CK(clk), .RN(n5727), .Q(\D_cache/cache[4][28] ), .QN(n2811) );
  DFFRX1 \D_cache/cache_reg[5][28]  ( .D(\D_cache/n1567 ), .CK(clk), .RN(n5727), .Q(\D_cache/cache[5][28] ), .QN(n819) );
  DFFRX1 \D_cache/cache_reg[6][28]  ( .D(\D_cache/n1566 ), .CK(clk), .RN(n5727), .Q(\D_cache/cache[6][28] ), .QN(n2446) );
  DFFRX1 \D_cache/cache_reg[7][28]  ( .D(\D_cache/n1565 ), .CK(clk), .RN(n5727), .Q(\D_cache/cache[7][28] ), .QN(n471) );
  DFFRX1 \D_cache/cache_reg[0][29]  ( .D(\D_cache/n1564 ), .CK(clk), .RN(n5727), .Q(\D_cache/cache[0][29] ), .QN(n1503) );
  DFFRX1 \D_cache/cache_reg[1][29]  ( .D(\D_cache/n1563 ), .CK(clk), .RN(n5727), .Q(\D_cache/cache[1][29] ), .QN(n3116) );
  DFFRX1 \D_cache/cache_reg[2][29]  ( .D(\D_cache/n1562 ), .CK(clk), .RN(n5727), .Q(\D_cache/cache[2][29] ), .QN(n1501) );
  DFFRX1 \D_cache/cache_reg[3][29]  ( .D(\D_cache/n1561 ), .CK(clk), .RN(n5727), .Q(\D_cache/cache[3][29] ), .QN(n3114) );
  DFFRX1 \D_cache/cache_reg[4][29]  ( .D(\D_cache/n1560 ), .CK(clk), .RN(n5727), .Q(\D_cache/cache[4][29] ), .QN(n1502) );
  DFFRX1 \D_cache/cache_reg[5][29]  ( .D(\D_cache/n1559 ), .CK(clk), .RN(n5727), .Q(\D_cache/cache[5][29] ), .QN(n3115) );
  DFFRX1 \D_cache/cache_reg[6][29]  ( .D(\D_cache/n1558 ), .CK(clk), .RN(n5727), .Q(\D_cache/cache[6][29] ), .QN(n1491) );
  DFFRX1 \D_cache/cache_reg[7][29]  ( .D(\D_cache/n1557 ), .CK(clk), .RN(n5728), .Q(\D_cache/cache[7][29] ), .QN(n3104) );
  DFFRX1 \D_cache/cache_reg[0][30]  ( .D(\D_cache/n1556 ), .CK(clk), .RN(n5728), .Q(\D_cache/cache[0][30] ), .QN(n816) );
  DFFRX1 \D_cache/cache_reg[1][30]  ( .D(\D_cache/n1555 ), .CK(clk), .RN(n5728), .Q(\D_cache/cache[1][30] ), .QN(n2348) );
  DFFRX1 \D_cache/cache_reg[2][30]  ( .D(\D_cache/n1554 ), .CK(clk), .RN(n5728), .Q(\D_cache/cache[2][30] ), .QN(n812) );
  DFFRX1 \D_cache/cache_reg[3][30]  ( .D(\D_cache/n1553 ), .CK(clk), .RN(n5728), .Q(\D_cache/cache[3][30] ), .QN(n2345) );
  DFFRX1 \D_cache/cache_reg[4][30]  ( .D(\D_cache/n1552 ), .CK(clk), .RN(n5728), .Q(\D_cache/cache[4][30] ), .QN(n813) );
  DFFRX1 \D_cache/cache_reg[5][30]  ( .D(\D_cache/n1551 ), .CK(clk), .RN(n5728), .Q(\D_cache/cache[5][30] ), .QN(n2346) );
  DFFRX1 \D_cache/cache_reg[6][30]  ( .D(\D_cache/n1550 ), .CK(clk), .RN(n5728), .Q(\D_cache/cache[6][30] ), .QN(n811) );
  DFFRX1 \D_cache/cache_reg[7][30]  ( .D(\D_cache/n1549 ), .CK(clk), .RN(n5728), .Q(\D_cache/cache[7][30] ), .QN(n2344) );
  DFFRX1 \D_cache/cache_reg[0][31]  ( .D(\D_cache/n1548 ), .CK(clk), .RN(n5728), .Q(\D_cache/cache[0][31] ), .QN(n1420) );
  DFFRX1 \D_cache/cache_reg[1][31]  ( .D(\D_cache/n1547 ), .CK(clk), .RN(n5728), .Q(\D_cache/cache[1][31] ), .QN(n3033) );
  DFFRX1 \D_cache/cache_reg[2][31]  ( .D(\D_cache/n1546 ), .CK(clk), .RN(n5728), .Q(\D_cache/cache[2][31] ), .QN(n1421) );
  DFFRX1 \D_cache/cache_reg[3][31]  ( .D(\D_cache/n1545 ), .CK(clk), .RN(n5729), .Q(\D_cache/cache[3][31] ), .QN(n3034) );
  DFFRX1 \D_cache/cache_reg[4][31]  ( .D(\D_cache/n1544 ), .CK(clk), .RN(n5729), .Q(\D_cache/cache[4][31] ), .QN(n1422) );
  DFFRX1 \D_cache/cache_reg[5][31]  ( .D(\D_cache/n1543 ), .CK(clk), .RN(n5729), .Q(\D_cache/cache[5][31] ), .QN(n3035) );
  DFFRX1 \D_cache/cache_reg[6][31]  ( .D(\D_cache/n1542 ), .CK(clk), .RN(n5729), .Q(\D_cache/cache[6][31] ), .QN(n1235) );
  DFFRX1 \D_cache/cache_reg[7][31]  ( .D(\D_cache/n1541 ), .CK(clk), .RN(n5729), .Q(\D_cache/cache[7][31] ), .QN(n2840) );
  DFFRX1 \D_cache/cache_reg[0][32]  ( .D(\D_cache/n1540 ), .CK(clk), .RN(n5729), .Q(\D_cache/cache[0][32] ), .QN(n1328) );
  DFFRX1 \D_cache/cache_reg[1][32]  ( .D(\D_cache/n1539 ), .CK(clk), .RN(n5729), .Q(\D_cache/cache[1][32] ), .QN(n2940) );
  DFFRX1 \D_cache/cache_reg[2][32]  ( .D(\D_cache/n1538 ), .CK(clk), .RN(n5729), .Q(\D_cache/cache[2][32] ), .QN(n1329) );
  DFFRX1 \D_cache/cache_reg[3][32]  ( .D(\D_cache/n1537 ), .CK(clk), .RN(n5729), .Q(\D_cache/cache[3][32] ), .QN(n2941) );
  DFFRX1 \D_cache/cache_reg[4][32]  ( .D(\D_cache/n1536 ), .CK(clk), .RN(n5729), .Q(\D_cache/cache[4][32] ), .QN(n1330) );
  DFFRX1 \D_cache/cache_reg[5][32]  ( .D(\D_cache/n1535 ), .CK(clk), .RN(n5729), .Q(\D_cache/cache[5][32] ), .QN(n2942) );
  DFFRX1 \D_cache/cache_reg[6][32]  ( .D(\D_cache/n1534 ), .CK(clk), .RN(n5729), .Q(\D_cache/cache[6][32] ), .QN(n1551) );
  DFFRX1 \D_cache/cache_reg[7][32]  ( .D(\D_cache/n1533 ), .CK(clk), .RN(n5730), .Q(\D_cache/cache[7][32] ), .QN(n3164) );
  DFFRX1 \D_cache/cache_reg[0][33]  ( .D(\D_cache/n1532 ), .CK(clk), .RN(n5730), .Q(\D_cache/cache[0][33] ), .QN(n1563) );
  DFFRX1 \D_cache/cache_reg[1][33]  ( .D(\D_cache/n1531 ), .CK(clk), .RN(n5730), .Q(\D_cache/cache[1][33] ), .QN(n3176) );
  DFFRX1 \D_cache/cache_reg[2][33]  ( .D(\D_cache/n1530 ), .CK(clk), .RN(n5730), .Q(\D_cache/cache[2][33] ), .QN(n1304) );
  DFFRX1 \D_cache/cache_reg[3][33]  ( .D(\D_cache/n1529 ), .CK(clk), .RN(n5730), .Q(\D_cache/cache[3][33] ), .QN(n2916) );
  DFFRX1 \D_cache/cache_reg[4][33]  ( .D(\D_cache/n1528 ), .CK(clk), .RN(n5730), .Q(\D_cache/cache[4][33] ), .QN(n1564) );
  DFFRX1 \D_cache/cache_reg[5][33]  ( .D(\D_cache/n1527 ), .CK(clk), .RN(n5730), .Q(\D_cache/cache[5][33] ), .QN(n3177) );
  DFFRX1 \D_cache/cache_reg[6][33]  ( .D(\D_cache/n1526 ), .CK(clk), .RN(n5730), .Q(\D_cache/cache[6][33] ), .QN(n1550) );
  DFFRX1 \D_cache/cache_reg[7][33]  ( .D(\D_cache/n1525 ), .CK(clk), .RN(n5730), .Q(\D_cache/cache[7][33] ), .QN(n3163) );
  DFFRX1 \D_cache/cache_reg[0][34]  ( .D(\D_cache/n1524 ), .CK(clk), .RN(n5730), .Q(\D_cache/cache[0][34] ), .QN(n1471) );
  DFFRX1 \D_cache/cache_reg[1][34]  ( .D(\D_cache/n1523 ), .CK(clk), .RN(n5730), .Q(\D_cache/cache[1][34] ), .QN(n3084) );
  DFFRX1 \D_cache/cache_reg[2][34]  ( .D(\D_cache/n1522 ), .CK(clk), .RN(n5730), .Q(\D_cache/cache[2][34] ), .QN(n1417) );
  DFFRX1 \D_cache/cache_reg[3][34]  ( .D(\D_cache/n1521 ), .CK(clk), .RN(n5731), .Q(\D_cache/cache[3][34] ), .QN(n3030) );
  DFFRX1 \D_cache/cache_reg[4][34]  ( .D(\D_cache/n1520 ), .CK(clk), .RN(n5731), .Q(\D_cache/cache[4][34] ), .QN(n1472) );
  DFFRX1 \D_cache/cache_reg[5][34]  ( .D(\D_cache/n1519 ), .CK(clk), .RN(n5731), .Q(\D_cache/cache[5][34] ), .QN(n3085) );
  DFFRX1 \D_cache/cache_reg[6][34]  ( .D(\D_cache/n1518 ), .CK(clk), .RN(n5731), .Q(\D_cache/cache[6][34] ), .QN(n1237) );
  DFFRX1 \D_cache/cache_reg[7][34]  ( .D(\D_cache/n1517 ), .CK(clk), .RN(n5731), .Q(\D_cache/cache[7][34] ), .QN(n2842) );
  DFFRX1 \D_cache/cache_reg[0][35]  ( .D(\D_cache/n1516 ), .CK(clk), .RN(n5731), .Q(\D_cache/cache[0][35] ), .QN(n1275) );
  DFFRX1 \D_cache/cache_reg[1][35]  ( .D(\D_cache/n1515 ), .CK(clk), .RN(n5731), .Q(\D_cache/cache[1][35] ), .QN(n2887) );
  DFFRX1 \D_cache/cache_reg[2][35]  ( .D(\D_cache/n1514 ), .CK(clk), .RN(n5731), .Q(\D_cache/cache[2][35] ), .QN(n1274) );
  DFFRX1 \D_cache/cache_reg[3][35]  ( .D(\D_cache/n1513 ), .CK(clk), .RN(n5731), .Q(\D_cache/cache[3][35] ), .QN(n2886) );
  DFFRX1 \D_cache/cache_reg[4][35]  ( .D(\D_cache/n1512 ), .CK(clk), .RN(n5731), .Q(\D_cache/cache[4][35] ), .QN(n1276) );
  DFFRX1 \D_cache/cache_reg[5][35]  ( .D(\D_cache/n1511 ), .CK(clk), .RN(n5731), .Q(\D_cache/cache[5][35] ), .QN(n2888) );
  DFFRX1 \D_cache/cache_reg[6][35]  ( .D(\D_cache/n1510 ), .CK(clk), .RN(n5731), .Q(\D_cache/cache[6][35] ), .QN(n1517) );
  DFFRX1 \D_cache/cache_reg[7][35]  ( .D(\D_cache/n1509 ), .CK(clk), .RN(n5732), .Q(\D_cache/cache[7][35] ), .QN(n3130) );
  DFFRX1 \D_cache/cache_reg[0][36]  ( .D(\D_cache/n1508 ), .CK(clk), .RN(n5732), .Q(\D_cache/cache[0][36] ), .QN(n1289) );
  DFFRX1 \D_cache/cache_reg[1][36]  ( .D(\D_cache/n1507 ), .CK(clk), .RN(n5732), .Q(\D_cache/cache[1][36] ), .QN(n2901) );
  DFFRX1 \D_cache/cache_reg[2][36]  ( .D(\D_cache/n1506 ), .CK(clk), .RN(n5732), .Q(\D_cache/cache[2][36] ), .QN(n1290) );
  DFFRX1 \D_cache/cache_reg[3][36]  ( .D(\D_cache/n1505 ), .CK(clk), .RN(n5732), .Q(\D_cache/cache[3][36] ), .QN(n2902) );
  DFFRX1 \D_cache/cache_reg[4][36]  ( .D(\D_cache/n1504 ), .CK(clk), .RN(n5732), .Q(\D_cache/cache[4][36] ), .QN(n2388) );
  DFFRX1 \D_cache/cache_reg[5][36]  ( .D(\D_cache/n1503 ), .CK(clk), .RN(n5732), .Q(\D_cache/cache[5][36] ), .QN(n883) );
  DFFRX1 \D_cache/cache_reg[6][36]  ( .D(\D_cache/n1502 ), .CK(clk), .RN(n5732), .Q(\D_cache/cache[6][36] ), .QN(n1476) );
  DFFRX1 \D_cache/cache_reg[7][36]  ( .D(\D_cache/n1501 ), .CK(clk), .RN(n5732), .Q(\D_cache/cache[7][36] ), .QN(n3089) );
  DFFRX1 \D_cache/cache_reg[0][37]  ( .D(\D_cache/n1500 ), .CK(clk), .RN(n5732), .Q(\D_cache/cache[0][37] ), .QN(n1277) );
  DFFRX1 \D_cache/cache_reg[1][37]  ( .D(\D_cache/n1499 ), .CK(clk), .RN(n5732), .Q(\D_cache/cache[1][37] ), .QN(n2889) );
  DFFRX1 \D_cache/cache_reg[2][37]  ( .D(\D_cache/n1498 ), .CK(clk), .RN(n5732), .Q(\D_cache/cache[2][37] ), .QN(n1278) );
  DFFRX1 \D_cache/cache_reg[3][37]  ( .D(\D_cache/n1497 ), .CK(clk), .RN(n5733), .Q(\D_cache/cache[3][37] ), .QN(n2890) );
  DFFRX1 \D_cache/cache_reg[4][37]  ( .D(\D_cache/n1496 ), .CK(clk), .RN(n5733), .Q(\D_cache/cache[4][37] ), .QN(n2387) );
  DFFRX1 \D_cache/cache_reg[5][37]  ( .D(\D_cache/n1495 ), .CK(clk), .RN(n5733), .Q(\D_cache/cache[5][37] ), .QN(n882) );
  DFFRX1 \D_cache/cache_reg[6][37]  ( .D(\D_cache/n1494 ), .CK(clk), .RN(n5733), .Q(\D_cache/cache[6][37] ), .QN(n1546) );
  DFFRX1 \D_cache/cache_reg[7][37]  ( .D(\D_cache/n1493 ), .CK(clk), .RN(n5733), .Q(\D_cache/cache[7][37] ), .QN(n3159) );
  DFFRX1 \D_cache/cache_reg[0][38]  ( .D(\D_cache/n1492 ), .CK(clk), .RN(n5733), .Q(\D_cache/cache[0][38] ), .QN(n1582) );
  DFFRX1 \D_cache/cache_reg[1][38]  ( .D(\D_cache/n1491 ), .CK(clk), .RN(n5733), .Q(\D_cache/cache[1][38] ), .QN(n3195) );
  DFFRX1 \D_cache/cache_reg[2][38]  ( .D(\D_cache/n1490 ), .CK(clk), .RN(n5733), .Q(\D_cache/cache[2][38] ), .QN(n1342) );
  DFFRX1 \D_cache/cache_reg[3][38]  ( .D(\D_cache/n1489 ), .CK(clk), .RN(n5733), .Q(\D_cache/cache[3][38] ), .QN(n2954) );
  DFFRX1 \D_cache/cache_reg[4][38]  ( .D(\D_cache/n1488 ), .CK(clk), .RN(n5733), .Q(\D_cache/cache[4][38] ), .QN(n1569) );
  DFFRX1 \D_cache/cache_reg[5][38]  ( .D(\D_cache/n1487 ), .CK(clk), .RN(n5733), .Q(\D_cache/cache[5][38] ), .QN(n3182) );
  DFFRX1 \D_cache/cache_reg[6][38]  ( .D(\D_cache/n1486 ), .CK(clk), .RN(n5733), .Q(\D_cache/cache[6][38] ), .QN(n1343) );
  DFFRX1 \D_cache/cache_reg[7][38]  ( .D(\D_cache/n1485 ), .CK(clk), .RN(n5734), .Q(\D_cache/cache[7][38] ), .QN(n2955) );
  DFFRX1 \D_cache/cache_reg[0][39]  ( .D(\D_cache/n1484 ), .CK(clk), .RN(n5734), .Q(\D_cache/cache[0][39] ), .QN(n1240) );
  DFFRX1 \D_cache/cache_reg[1][39]  ( .D(\D_cache/n1483 ), .CK(clk), .RN(n5734), .Q(\D_cache/cache[1][39] ), .QN(n2845) );
  DFFRX1 \D_cache/cache_reg[2][39]  ( .D(\D_cache/n1482 ), .CK(clk), .RN(n5734), .Q(\D_cache/cache[2][39] ), .QN(n1337) );
  DFFRX1 \D_cache/cache_reg[3][39]  ( .D(\D_cache/n1481 ), .CK(clk), .RN(n5734), .Q(\D_cache/cache[3][39] ), .QN(n2949) );
  DFFRX1 \D_cache/cache_reg[4][39]  ( .D(\D_cache/n1480 ), .CK(clk), .RN(n5734), .Q(\D_cache/cache[4][39] ), .QN(n1338) );
  DFFRX1 \D_cache/cache_reg[5][39]  ( .D(\D_cache/n1479 ), .CK(clk), .RN(n5734), .Q(\D_cache/cache[5][39] ), .QN(n2950) );
  DFFRX1 \D_cache/cache_reg[6][39]  ( .D(\D_cache/n1478 ), .CK(clk), .RN(n5734), .Q(\D_cache/cache[6][39] ), .QN(n1339) );
  DFFRX1 \D_cache/cache_reg[7][39]  ( .D(\D_cache/n1477 ), .CK(clk), .RN(n5734), .Q(\D_cache/cache[7][39] ), .QN(n2951) );
  DFFRX1 \D_cache/cache_reg[0][40]  ( .D(\D_cache/n1476 ), .CK(clk), .RN(n5734), .Q(\D_cache/cache[0][40] ), .QN(n1358) );
  DFFRX1 \D_cache/cache_reg[1][40]  ( .D(\D_cache/n1475 ), .CK(clk), .RN(n5734), .Q(\D_cache/cache[1][40] ), .QN(n2971) );
  DFFRX1 \D_cache/cache_reg[2][40]  ( .D(\D_cache/n1474 ), .CK(clk), .RN(n5734), .Q(\D_cache/cache[2][40] ), .QN(n1357) );
  DFFRX1 \D_cache/cache_reg[3][40]  ( .D(\D_cache/n1473 ), .CK(clk), .RN(n5735), .Q(\D_cache/cache[3][40] ), .QN(n2970) );
  DFFRX1 \D_cache/cache_reg[4][40]  ( .D(\D_cache/n1472 ), .CK(clk), .RN(n5735), .Q(\D_cache/cache[4][40] ), .QN(n936) );
  DFFRX1 \D_cache/cache_reg[5][40]  ( .D(\D_cache/n1471 ), .CK(clk), .RN(n5735), .Q(\D_cache/cache[5][40] ), .QN(n2461) );
  DFFRX1 \D_cache/cache_reg[6][40]  ( .D(\D_cache/n1470 ), .CK(clk), .RN(n5735), .Q(\D_cache/cache[6][40] ), .QN(n1455) );
  DFFRX1 \D_cache/cache_reg[7][40]  ( .D(\D_cache/n1469 ), .CK(clk), .RN(n5735), .Q(\D_cache/cache[7][40] ), .QN(n3068) );
  DFFRX1 \D_cache/cache_reg[0][41]  ( .D(\D_cache/n1468 ), .CK(clk), .RN(n5735), .Q(\D_cache/cache[0][41] ), .QN(n1350) );
  DFFRX1 \D_cache/cache_reg[1][41]  ( .D(\D_cache/n1467 ), .CK(clk), .RN(n5735), .Q(\D_cache/cache[1][41] ), .QN(n2963) );
  DFFRX1 \D_cache/cache_reg[2][41]  ( .D(\D_cache/n1466 ), .CK(clk), .RN(n5735), .Q(\D_cache/cache[2][41] ), .QN(n1349) );
  DFFRX1 \D_cache/cache_reg[3][41]  ( .D(\D_cache/n1465 ), .CK(clk), .RN(n5735), .Q(\D_cache/cache[3][41] ), .QN(n2961) );
  DFFRX1 \D_cache/cache_reg[4][41]  ( .D(\D_cache/n1464 ), .CK(clk), .RN(n5735), .Q(\D_cache/cache[4][41] ), .QN(n1229) );
  DFFRX1 \D_cache/cache_reg[5][41]  ( .D(\D_cache/n1463 ), .CK(clk), .RN(n5735), .Q(\D_cache/cache[5][41] ), .QN(n2962) );
  DFFRX1 \D_cache/cache_reg[6][41]  ( .D(\D_cache/n1462 ), .CK(clk), .RN(n5735), .Q(\D_cache/cache[6][41] ), .QN(n1453) );
  DFFRX1 \D_cache/cache_reg[7][41]  ( .D(\D_cache/n1461 ), .CK(clk), .RN(n5736), .Q(\D_cache/cache[7][41] ), .QN(n3066) );
  DFFRX1 \D_cache/cache_reg[0][42]  ( .D(\D_cache/n1460 ), .CK(clk), .RN(n5736), .Q(\D_cache/cache[0][42] ), .QN(n2377) );
  DFFRX1 \D_cache/cache_reg[1][42]  ( .D(\D_cache/n1459 ), .CK(clk), .RN(n5736), .Q(\D_cache/cache[1][42] ), .QN(n873) );
  DFFRX1 \D_cache/cache_reg[2][42]  ( .D(\D_cache/n1458 ), .CK(clk), .RN(n5736), .Q(\D_cache/cache[2][42] ), .QN(n1283) );
  DFFRX1 \D_cache/cache_reg[3][42]  ( .D(\D_cache/n1457 ), .CK(clk), .RN(n5736), .Q(\D_cache/cache[3][42] ), .QN(n2895) );
  DFFRX1 \D_cache/cache_reg[4][42]  ( .D(\D_cache/n1456 ), .CK(clk), .RN(n5736), .Q(\D_cache/cache[4][42] ), .QN(n2397) );
  DFFRX1 \D_cache/cache_reg[5][42]  ( .D(\D_cache/n1455 ), .CK(clk), .RN(n5736), .Q(\D_cache/cache[5][42] ), .QN(n892) );
  DFFRX1 \D_cache/cache_reg[6][42]  ( .D(\D_cache/n1454 ), .CK(clk), .RN(n5736), .Q(\D_cache/cache[6][42] ), .QN(n1543) );
  DFFRX1 \D_cache/cache_reg[7][42]  ( .D(\D_cache/n1453 ), .CK(clk), .RN(n5736), .Q(\D_cache/cache[7][42] ), .QN(n3156) );
  DFFRX1 \D_cache/cache_reg[0][43]  ( .D(\D_cache/n1452 ), .CK(clk), .RN(n5736), .Q(\D_cache/cache[0][43] ), .QN(n1286) );
  DFFRX1 \D_cache/cache_reg[1][43]  ( .D(\D_cache/n1451 ), .CK(clk), .RN(n5736), .Q(\D_cache/cache[1][43] ), .QN(n2898) );
  DFFRX1 \D_cache/cache_reg[2][43]  ( .D(\D_cache/n1450 ), .CK(clk), .RN(n5736), .Q(\D_cache/cache[2][43] ), .QN(n1287) );
  DFFRX1 \D_cache/cache_reg[3][43]  ( .D(\D_cache/n1449 ), .CK(clk), .RN(n5737), .Q(\D_cache/cache[3][43] ), .QN(n2899) );
  DFFRX1 \D_cache/cache_reg[4][43]  ( .D(\D_cache/n1448 ), .CK(clk), .RN(n5737), .Q(\D_cache/cache[4][43] ), .QN(n1288) );
  DFFRX1 \D_cache/cache_reg[5][43]  ( .D(\D_cache/n1447 ), .CK(clk), .RN(n5737), .Q(\D_cache/cache[5][43] ), .QN(n2900) );
  DFFRX1 \D_cache/cache_reg[6][43]  ( .D(\D_cache/n1446 ), .CK(clk), .RN(n5737), .Q(\D_cache/cache[6][43] ), .QN(n1247) );
  DFFRX1 \D_cache/cache_reg[7][43]  ( .D(\D_cache/n1445 ), .CK(clk), .RN(n5737), .Q(\D_cache/cache[7][43] ), .QN(n2855) );
  DFFRX1 \D_cache/cache_reg[0][44]  ( .D(\D_cache/n1444 ), .CK(clk), .RN(n5737), .Q(\D_cache/cache[0][44] ), .QN(n1352) );
  DFFRX1 \D_cache/cache_reg[1][44]  ( .D(\D_cache/n1443 ), .CK(clk), .RN(n5737), .Q(\D_cache/cache[1][44] ), .QN(n2965) );
  DFFRX1 \D_cache/cache_reg[2][44]  ( .D(\D_cache/n1442 ), .CK(clk), .RN(n5737), .Q(\D_cache/cache[2][44] ), .QN(n1351) );
  DFFRX1 \D_cache/cache_reg[3][44]  ( .D(\D_cache/n1441 ), .CK(clk), .RN(n5737), .Q(\D_cache/cache[3][44] ), .QN(n2964) );
  DFFRX1 \D_cache/cache_reg[4][44]  ( .D(\D_cache/n1440 ), .CK(clk), .RN(n5737), .Q(\D_cache/cache[4][44] ), .QN(n2363) );
  DFFRX1 \D_cache/cache_reg[5][44]  ( .D(\D_cache/n1439 ), .CK(clk), .RN(n5737), .Q(\D_cache/cache[5][44] ), .QN(n860) );
  DFFRX1 \D_cache/cache_reg[6][44]  ( .D(\D_cache/n1438 ), .CK(clk), .RN(n5737), .Q(\D_cache/cache[6][44] ), .QN(n1539) );
  DFFRX1 \D_cache/cache_reg[7][44]  ( .D(\D_cache/n1437 ), .CK(clk), .RN(n5738), .Q(\D_cache/cache[7][44] ), .QN(n3152) );
  DFFRX1 \D_cache/cache_reg[0][45]  ( .D(\D_cache/n1436 ), .CK(clk), .RN(n5738), .Q(\D_cache/cache[0][45] ), .QN(n1345) );
  DFFRX1 \D_cache/cache_reg[1][45]  ( .D(\D_cache/n1435 ), .CK(clk), .RN(n5738), .Q(\D_cache/cache[1][45] ), .QN(n2957) );
  DFFRX1 \D_cache/cache_reg[2][45]  ( .D(\D_cache/n1434 ), .CK(clk), .RN(n5738), .Q(\D_cache/cache[2][45] ), .QN(n1344) );
  DFFRX1 \D_cache/cache_reg[3][45]  ( .D(\D_cache/n1433 ), .CK(clk), .RN(n5738), .Q(\D_cache/cache[3][45] ), .QN(n2956) );
  DFFRX1 \D_cache/cache_reg[4][45]  ( .D(\D_cache/n1432 ), .CK(clk), .RN(n5738), .Q(\D_cache/cache[4][45] ), .QN(n2367) );
  DFFRX1 \D_cache/cache_reg[5][45]  ( .D(\D_cache/n1431 ), .CK(clk), .RN(n5738), .Q(\D_cache/cache[5][45] ), .QN(n864) );
  DFFRX1 \D_cache/cache_reg[6][45]  ( .D(\D_cache/n1430 ), .CK(clk), .RN(n5738), .Q(\D_cache/cache[6][45] ), .QN(n1486) );
  DFFRX1 \D_cache/cache_reg[7][45]  ( .D(\D_cache/n1429 ), .CK(clk), .RN(n5738), .Q(\D_cache/cache[7][45] ), .QN(n3099) );
  DFFRX1 \D_cache/cache_reg[0][46]  ( .D(\D_cache/n1428 ), .CK(clk), .RN(n5738), .Q(\D_cache/cache[0][46] ), .QN(n2378) );
  DFFRX1 \D_cache/cache_reg[1][46]  ( .D(\D_cache/n1427 ), .CK(clk), .RN(n5738), .Q(\D_cache/cache[1][46] ), .QN(n874) );
  DFFRX1 \D_cache/cache_reg[2][46]  ( .D(\D_cache/n1426 ), .CK(clk), .RN(n5738), .Q(\D_cache/cache[2][46] ), .QN(n1457) );
  DFFRX1 \D_cache/cache_reg[3][46]  ( .D(\D_cache/n1425 ), .CK(clk), .RN(n5739), .Q(\D_cache/cache[3][46] ), .QN(n3070) );
  DFFRX1 \D_cache/cache_reg[4][46]  ( .D(\D_cache/n1424 ), .CK(clk), .RN(n5739), .Q(\D_cache/cache[4][46] ), .QN(n2394) );
  DFFRX1 \D_cache/cache_reg[5][46]  ( .D(\D_cache/n1423 ), .CK(clk), .RN(n5739), .Q(\D_cache/cache[5][46] ), .QN(n889) );
  DFFRX1 \D_cache/cache_reg[6][46]  ( .D(\D_cache/n1422 ), .CK(clk), .RN(n5739), .Q(\D_cache/cache[6][46] ), .QN(n1452) );
  DFFRX1 \D_cache/cache_reg[7][46]  ( .D(\D_cache/n1421 ), .CK(clk), .RN(n5739), .Q(\D_cache/cache[7][46] ), .QN(n3065) );
  DFFRX1 \D_cache/cache_reg[0][47]  ( .D(\D_cache/n1420 ), .CK(clk), .RN(n5739), .Q(\D_cache/cache[0][47] ), .QN(n2372) );
  DFFRX1 \D_cache/cache_reg[1][47]  ( .D(\D_cache/n1419 ), .CK(clk), .RN(n5739), .Q(\D_cache/cache[1][47] ), .QN(n868) );
  DFFRX1 \D_cache/cache_reg[2][47]  ( .D(\D_cache/n1418 ), .CK(clk), .RN(n5739), .Q(\D_cache/cache[2][47] ), .QN(n1233) );
  DFFRX1 \D_cache/cache_reg[3][47]  ( .D(\D_cache/n1417 ), .CK(clk), .RN(n5739), .Q(\D_cache/cache[3][47] ), .QN(n2838) );
  DFFRX1 \D_cache/cache_reg[4][47]  ( .D(\D_cache/n1416 ), .CK(clk), .RN(n5739), .Q(\D_cache/cache[4][47] ), .QN(n2390) );
  DFFRX1 \D_cache/cache_reg[5][47]  ( .D(\D_cache/n1415 ), .CK(clk), .RN(n5739), .Q(\D_cache/cache[5][47] ), .QN(n885) );
  DFFRX1 \D_cache/cache_reg[6][47]  ( .D(\D_cache/n1414 ), .CK(clk), .RN(n5739), .Q(\D_cache/cache[6][47] ), .QN(n1440) );
  DFFRX1 \D_cache/cache_reg[7][47]  ( .D(\D_cache/n1413 ), .CK(clk), .RN(n5740), .Q(\D_cache/cache[7][47] ), .QN(n3053) );
  DFFRX1 \D_cache/cache_reg[0][48]  ( .D(\D_cache/n1412 ), .CK(clk), .RN(n5740), .Q(\D_cache/cache[0][48] ), .QN(n1292) );
  DFFRX1 \D_cache/cache_reg[1][48]  ( .D(\D_cache/n1411 ), .CK(clk), .RN(n5740), .Q(\D_cache/cache[1][48] ), .QN(n2904) );
  DFFRX1 \D_cache/cache_reg[2][48]  ( .D(\D_cache/n1410 ), .CK(clk), .RN(n5740), .Q(\D_cache/cache[2][48] ), .QN(n1291) );
  DFFRX1 \D_cache/cache_reg[3][48]  ( .D(\D_cache/n1409 ), .CK(clk), .RN(n5740), .Q(\D_cache/cache[3][48] ), .QN(n2903) );
  DFFRX1 \D_cache/cache_reg[4][48]  ( .D(\D_cache/n1408 ), .CK(clk), .RN(n5740), .Q(\D_cache/cache[4][48] ), .QN(n1293) );
  DFFRX1 \D_cache/cache_reg[5][48]  ( .D(\D_cache/n1407 ), .CK(clk), .RN(n5740), .Q(\D_cache/cache[5][48] ), .QN(n2905) );
  DFFRX1 \D_cache/cache_reg[6][48]  ( .D(\D_cache/n1406 ), .CK(clk), .RN(n5740), .Q(\D_cache/cache[6][48] ), .QN(n1480) );
  DFFRX1 \D_cache/cache_reg[7][48]  ( .D(\D_cache/n1405 ), .CK(clk), .RN(n5740), .Q(\D_cache/cache[7][48] ), .QN(n3093) );
  DFFRX1 \D_cache/cache_reg[0][49]  ( .D(\D_cache/n1404 ), .CK(clk), .RN(n5740), .Q(\D_cache/cache[0][49] ), .QN(n1562) );
  DFFRX1 \D_cache/cache_reg[1][49]  ( .D(\D_cache/n1403 ), .CK(clk), .RN(n5740), .Q(\D_cache/cache[1][49] ), .QN(n3175) );
  DFFRX1 \D_cache/cache_reg[2][49]  ( .D(\D_cache/n1402 ), .CK(clk), .RN(n5740), .Q(\D_cache/cache[2][49] ), .QN(n2358) );
  DFFRX1 \D_cache/cache_reg[3][49]  ( .D(\D_cache/n1401 ), .CK(clk), .RN(n5741), .Q(\D_cache/cache[3][49] ), .QN(n855) );
  DFFRX1 \D_cache/cache_reg[4][49]  ( .D(\D_cache/n1400 ), .CK(clk), .RN(n5741), .Q(\D_cache/cache[4][49] ), .QN(n1561) );
  DFFRX1 \D_cache/cache_reg[5][49]  ( .D(\D_cache/n1399 ), .CK(clk), .RN(n5741), .Q(\D_cache/cache[5][49] ), .QN(n3174) );
  DFFRX1 \D_cache/cache_reg[6][49]  ( .D(\D_cache/n1398 ), .CK(clk), .RN(n5741), .Q(\D_cache/cache[6][49] ), .QN(n1512) );
  DFFRX1 \D_cache/cache_reg[7][49]  ( .D(\D_cache/n1397 ), .CK(clk), .RN(n5741), .Q(\D_cache/cache[7][49] ), .QN(n3125) );
  DFFRX1 \D_cache/cache_reg[0][50]  ( .D(\D_cache/n1396 ), .CK(clk), .RN(n5741), .Q(\D_cache/cache[0][50] ), .QN(n1324) );
  DFFRX1 \D_cache/cache_reg[1][50]  ( .D(\D_cache/n1395 ), .CK(clk), .RN(n5741), .Q(\D_cache/cache[1][50] ), .QN(n2936) );
  DFFRX1 \D_cache/cache_reg[2][50]  ( .D(\D_cache/n1394 ), .CK(clk), .RN(n5741), .Q(\D_cache/cache[2][50] ), .QN(n1325) );
  DFFRX1 \D_cache/cache_reg[3][50]  ( .D(\D_cache/n1393 ), .CK(clk), .RN(n5741), .Q(\D_cache/cache[3][50] ), .QN(n2937) );
  DFFRX1 \D_cache/cache_reg[4][50]  ( .D(\D_cache/n1392 ), .CK(clk), .RN(n5741), .Q(\D_cache/cache[4][50] ), .QN(n2814) );
  DFFRX1 \D_cache/cache_reg[5][50]  ( .D(\D_cache/n1391 ), .CK(clk), .RN(n5741), .Q(\D_cache/cache[5][50] ), .QN(n822) );
  DFFRX1 \D_cache/cache_reg[6][50]  ( .D(\D_cache/n1390 ), .CK(clk), .RN(n5741), .Q(\D_cache/cache[6][50] ), .QN(n1451) );
  DFFRX1 \D_cache/cache_reg[7][50]  ( .D(\D_cache/n1389 ), .CK(clk), .RN(n5742), .Q(\D_cache/cache[7][50] ), .QN(n3064) );
  DFFRX1 \D_cache/cache_reg[0][51]  ( .D(\D_cache/n1388 ), .CK(clk), .RN(n5742), .Q(\D_cache/cache[0][51] ), .QN(n953) );
  DFFRX1 \D_cache/cache_reg[1][51]  ( .D(\D_cache/n1387 ), .CK(clk), .RN(n5742), .Q(\D_cache/cache[1][51] ), .QN(n2478) );
  DFFRX1 \D_cache/cache_reg[2][51]  ( .D(\D_cache/n1386 ), .CK(clk), .RN(n5742), .Q(\D_cache/cache[2][51] ), .QN(n952) );
  DFFRX1 \D_cache/cache_reg[3][51]  ( .D(\D_cache/n1385 ), .CK(clk), .RN(n5742), .Q(\D_cache/cache[3][51] ), .QN(n2477) );
  DFFRX1 \D_cache/cache_reg[4][51]  ( .D(\D_cache/n1384 ), .CK(clk), .RN(n5742), .Q(\D_cache/cache[4][51] ), .QN(n1567) );
  DFFRX1 \D_cache/cache_reg[5][51]  ( .D(\D_cache/n1383 ), .CK(clk), .RN(n5742), .Q(\D_cache/cache[5][51] ), .QN(n3180) );
  DFFRX1 \D_cache/cache_reg[6][51]  ( .D(\D_cache/n1382 ), .CK(clk), .RN(n5742), .Q(\D_cache/cache[6][51] ), .QN(n1526) );
  DFFRX1 \D_cache/cache_reg[7][51]  ( .D(\D_cache/n1381 ), .CK(clk), .RN(n5742), .Q(\D_cache/cache[7][51] ), .QN(n3139) );
  DFFRX1 \D_cache/cache_reg[0][52]  ( .D(\D_cache/n1380 ), .CK(clk), .RN(n5742), .Q(\D_cache/cache[0][52] ), .QN(n1307) );
  DFFRX1 \D_cache/cache_reg[1][52]  ( .D(\D_cache/n1379 ), .CK(clk), .RN(n5742), .Q(\D_cache/cache[1][52] ), .QN(n2919) );
  DFFRX1 \D_cache/cache_reg[2][52]  ( .D(\D_cache/n1378 ), .CK(clk), .RN(n5742), .Q(\D_cache/cache[2][52] ), .QN(n1306) );
  DFFRX1 \D_cache/cache_reg[3][52]  ( .D(\D_cache/n1377 ), .CK(clk), .RN(n5743), .Q(\D_cache/cache[3][52] ), .QN(n2918) );
  DFFRX1 \D_cache/cache_reg[4][52]  ( .D(\D_cache/n1376 ), .CK(clk), .RN(n5743), .Q(\D_cache/cache[4][52] ), .QN(n1308) );
  DFFRX1 \D_cache/cache_reg[5][52]  ( .D(\D_cache/n1375 ), .CK(clk), .RN(n5743), .Q(\D_cache/cache[5][52] ), .QN(n2920) );
  DFFRX1 \D_cache/cache_reg[6][52]  ( .D(\D_cache/n1374 ), .CK(clk), .RN(n5743), .Q(\D_cache/cache[6][52] ), .QN(n1525) );
  DFFRX1 \D_cache/cache_reg[7][52]  ( .D(\D_cache/n1373 ), .CK(clk), .RN(n5743), .Q(\D_cache/cache[7][52] ), .QN(n3138) );
  DFFRX1 \D_cache/cache_reg[0][53]  ( .D(\D_cache/n1372 ), .CK(clk), .RN(n5743), .Q(\D_cache/cache[0][53] ), .QN(n1314) );
  DFFRX1 \D_cache/cache_reg[1][53]  ( .D(\D_cache/n1371 ), .CK(clk), .RN(n5743), .Q(\D_cache/cache[1][53] ), .QN(n2926) );
  DFFRX1 \D_cache/cache_reg[2][53]  ( .D(\D_cache/n1370 ), .CK(clk), .RN(n5743), .Q(\D_cache/cache[2][53] ), .QN(n1466) );
  DFFRX1 \D_cache/cache_reg[3][53]  ( .D(\D_cache/n1369 ), .CK(clk), .RN(n5743), .Q(\D_cache/cache[3][53] ), .QN(n3079) );
  DFFRX1 \D_cache/cache_reg[4][53]  ( .D(\D_cache/n1368 ), .CK(clk), .RN(n5743), .Q(\D_cache/cache[4][53] ), .QN(n2851) );
  DFFRX1 \D_cache/cache_reg[5][53]  ( .D(\D_cache/n1367 ), .CK(clk), .RN(n5743), .Q(\D_cache/cache[5][53] ), .QN(n845) );
  DFFRX1 \D_cache/cache_reg[6][53]  ( .D(\D_cache/n1366 ), .CK(clk), .RN(n5743), .Q(\D_cache/cache[6][53] ), .QN(n2859) );
  DFFRX1 \D_cache/cache_reg[7][53]  ( .D(\D_cache/n1365 ), .CK(clk), .RN(n5744), .Q(\D_cache/cache[7][53] ), .QN(n1230) );
  DFFRX1 \D_cache/cache_reg[0][54]  ( .D(\D_cache/n1364 ), .CK(clk), .RN(n5744), .Q(\D_cache/cache[0][54] ), .QN(n1318) );
  DFFRX1 \D_cache/cache_reg[1][54]  ( .D(\D_cache/n1363 ), .CK(clk), .RN(n5744), .Q(\D_cache/cache[1][54] ), .QN(n2930) );
  DFFRX1 \D_cache/cache_reg[2][54]  ( .D(\D_cache/n1362 ), .CK(clk), .RN(n5744), .Q(\D_cache/cache[2][54] ), .QN(n1316) );
  DFFRX1 \D_cache/cache_reg[3][54]  ( .D(\D_cache/n1361 ), .CK(clk), .RN(n5744), .Q(\D_cache/cache[3][54] ), .QN(n2928) );
  DFFRX1 \D_cache/cache_reg[4][54]  ( .D(\D_cache/n1360 ), .CK(clk), .RN(n5744), .Q(\D_cache/cache[4][54] ), .QN(n1317) );
  DFFRX1 \D_cache/cache_reg[5][54]  ( .D(\D_cache/n1359 ), .CK(clk), .RN(n5744), .Q(\D_cache/cache[5][54] ), .QN(n2929) );
  DFFRX1 \D_cache/cache_reg[6][54]  ( .D(\D_cache/n1358 ), .CK(clk), .RN(n5744), .Q(\D_cache/cache[6][54] ), .QN(n1529) );
  DFFRX1 \D_cache/cache_reg[7][54]  ( .D(\D_cache/n1357 ), .CK(clk), .RN(n5744), .Q(\D_cache/cache[7][54] ), .QN(n3142) );
  DFFRX1 \D_cache/cache_reg[0][55]  ( .D(\D_cache/n1356 ), .CK(clk), .RN(n5744), .Q(\D_cache/cache[0][55] ), .QN(n1462) );
  DFFRX1 \D_cache/cache_reg[1][55]  ( .D(\D_cache/n1355 ), .CK(clk), .RN(n5744), .Q(\D_cache/cache[1][55] ), .QN(n3075) );
  DFFRX1 \D_cache/cache_reg[2][55]  ( .D(\D_cache/n1354 ), .CK(clk), .RN(n5744), .Q(\D_cache/cache[2][55] ), .QN(n1418) );
  DFFRX1 \D_cache/cache_reg[3][55]  ( .D(\D_cache/n1353 ), .CK(clk), .RN(n5745), .Q(\D_cache/cache[3][55] ), .QN(n3031) );
  DFFRX1 \D_cache/cache_reg[4][55]  ( .D(\D_cache/n1352 ), .CK(clk), .RN(n5745), .Q(\D_cache/cache[4][55] ), .QN(n1419) );
  DFFRX1 \D_cache/cache_reg[5][55]  ( .D(\D_cache/n1351 ), .CK(clk), .RN(n5745), .Q(\D_cache/cache[5][55] ), .QN(n3032) );
  DFFRX1 \D_cache/cache_reg[6][55]  ( .D(\D_cache/n1350 ), .CK(clk), .RN(n5745), .Q(\D_cache/cache[6][55] ), .QN(n1511) );
  DFFRX1 \D_cache/cache_reg[7][55]  ( .D(\D_cache/n1349 ), .CK(clk), .RN(n5745), .Q(\D_cache/cache[7][55] ), .QN(n3124) );
  DFFRX1 \D_cache/cache_reg[0][56]  ( .D(\D_cache/n1348 ), .CK(clk), .RN(n5745), .Q(\D_cache/cache[0][56] ), .QN(n1270) );
  DFFRX1 \D_cache/cache_reg[1][56]  ( .D(\D_cache/n1347 ), .CK(clk), .RN(n5745), .Q(\D_cache/cache[1][56] ), .QN(n2881) );
  DFFRX1 \D_cache/cache_reg[2][56]  ( .D(\D_cache/n1346 ), .CK(clk), .RN(n5745), .Q(\D_cache/cache[2][56] ), .QN(n1269) );
  DFFRX1 \D_cache/cache_reg[3][56]  ( .D(\D_cache/n1345 ), .CK(clk), .RN(n5745), .Q(\D_cache/cache[3][56] ), .QN(n2880) );
  DFFRX1 \D_cache/cache_reg[4][56]  ( .D(\D_cache/n1344 ), .CK(clk), .RN(n5745), .Q(\D_cache/cache[4][56] ), .QN(n1271) );
  DFFRX1 \D_cache/cache_reg[5][56]  ( .D(\D_cache/n1343 ), .CK(clk), .RN(n5745), .Q(\D_cache/cache[5][56] ), .QN(n2882) );
  DFFRX1 \D_cache/cache_reg[6][56]  ( .D(\D_cache/n1342 ), .CK(clk), .RN(n5745), .Q(\D_cache/cache[6][56] ), .QN(n1515) );
  DFFRX1 \D_cache/cache_reg[7][56]  ( .D(\D_cache/n1341 ), .CK(clk), .RN(n5746), .Q(\D_cache/cache[7][56] ), .QN(n3128) );
  DFFRX1 \D_cache/cache_reg[0][57]  ( .D(\D_cache/n1340 ), .CK(clk), .RN(n5746), .Q(\D_cache/cache[0][57] ), .QN(n1333) );
  DFFRX1 \D_cache/cache_reg[1][57]  ( .D(\D_cache/n1339 ), .CK(clk), .RN(n5746), .Q(\D_cache/cache[1][57] ), .QN(n2945) );
  DFFRX1 \D_cache/cache_reg[2][57]  ( .D(\D_cache/n1338 ), .CK(clk), .RN(n5746), .Q(\D_cache/cache[2][57] ), .QN(n1331) );
  DFFRX1 \D_cache/cache_reg[3][57]  ( .D(\D_cache/n1337 ), .CK(clk), .RN(n5746), .Q(\D_cache/cache[3][57] ), .QN(n2943) );
  DFFRX1 \D_cache/cache_reg[4][57]  ( .D(\D_cache/n1336 ), .CK(clk), .RN(n5746), .Q(\D_cache/cache[4][57] ), .QN(n1332) );
  DFFRX1 \D_cache/cache_reg[5][57]  ( .D(\D_cache/n1335 ), .CK(clk), .RN(n5746), .Q(\D_cache/cache[5][57] ), .QN(n2944) );
  DFFRX1 \D_cache/cache_reg[6][57]  ( .D(\D_cache/n1334 ), .CK(clk), .RN(n5746), .Q(\D_cache/cache[6][57] ), .QN(n1481) );
  DFFRX1 \D_cache/cache_reg[7][57]  ( .D(\D_cache/n1333 ), .CK(clk), .RN(n5746), .Q(\D_cache/cache[7][57] ), .QN(n3094) );
  DFFRX1 \D_cache/cache_reg[0][58]  ( .D(\D_cache/n1332 ), .CK(clk), .RN(n5746), .Q(\D_cache/cache[0][58] ), .QN(n2406) );
  DFFRX1 \D_cache/cache_reg[1][58]  ( .D(\D_cache/n1331 ), .CK(clk), .RN(n5746), .Q(\D_cache/cache[1][58] ), .QN(n900) );
  DFFRX1 \D_cache/cache_reg[2][58]  ( .D(\D_cache/n1330 ), .CK(clk), .RN(n5746), .Q(\D_cache/cache[2][58] ), .QN(n1296) );
  DFFRX1 \D_cache/cache_reg[3][58]  ( .D(\D_cache/n1329 ), .CK(clk), .RN(n5747), .Q(\D_cache/cache[3][58] ), .QN(n2908) );
  DFFRX1 \D_cache/cache_reg[4][58]  ( .D(\D_cache/n1328 ), .CK(clk), .RN(n5747), .Q(\D_cache/cache[4][58] ), .QN(n1297) );
  DFFRX1 \D_cache/cache_reg[5][58]  ( .D(\D_cache/n1327 ), .CK(clk), .RN(n5747), .Q(\D_cache/cache[5][58] ), .QN(n2909) );
  DFFRX1 \D_cache/cache_reg[6][58]  ( .D(\D_cache/n1326 ), .CK(clk), .RN(n5747), .Q(\D_cache/cache[6][58] ), .QN(n1521) );
  DFFRX1 \D_cache/cache_reg[7][58]  ( .D(\D_cache/n1325 ), .CK(clk), .RN(n5747), .Q(\D_cache/cache[7][58] ), .QN(n3134) );
  DFFRX1 \D_cache/cache_reg[0][59]  ( .D(\D_cache/n1324 ), .CK(clk), .RN(n5747), .Q(\D_cache/cache[0][59] ), .QN(n1298) );
  DFFRX1 \D_cache/cache_reg[1][59]  ( .D(\D_cache/n1323 ), .CK(clk), .RN(n5747), .Q(\D_cache/cache[1][59] ), .QN(n2910) );
  DFFRX1 \D_cache/cache_reg[2][59]  ( .D(\D_cache/n1322 ), .CK(clk), .RN(n5747), .Q(\D_cache/cache[2][59] ), .QN(n2405) );
  DFFRX1 \D_cache/cache_reg[3][59]  ( .D(\D_cache/n1321 ), .CK(clk), .RN(n5747), .Q(\D_cache/cache[3][59] ), .QN(n899) );
  DFFRX1 \D_cache/cache_reg[4][59]  ( .D(\D_cache/n1320 ), .CK(clk), .RN(n5747), .Q(\D_cache/cache[4][59] ), .QN(n2414) );
  DFFRX1 \D_cache/cache_reg[5][59]  ( .D(\D_cache/n1319 ), .CK(clk), .RN(n5747), .Q(\D_cache/cache[5][59] ), .QN(n905) );
  DFFRX1 \D_cache/cache_reg[6][59]  ( .D(\D_cache/n1318 ), .CK(clk), .RN(n5747), .Q(\D_cache/cache[6][59] ), .QN(n2403) );
  DFFRX1 \D_cache/cache_reg[7][59]  ( .D(\D_cache/n1317 ), .CK(clk), .RN(n5748), .Q(\D_cache/cache[7][59] ), .QN(n897) );
  DFFRX1 \D_cache/cache_reg[0][60]  ( .D(\D_cache/n1316 ), .CK(clk), .RN(n5748), .Q(\D_cache/cache[0][60] ), .QN(n1254) );
  DFFRX1 \D_cache/cache_reg[1][60]  ( .D(\D_cache/n1315 ), .CK(clk), .RN(n5748), .Q(\D_cache/cache[1][60] ), .QN(n2865) );
  DFFRX1 \D_cache/cache_reg[2][60]  ( .D(\D_cache/n1314 ), .CK(clk), .RN(n5748), .Q(\D_cache/cache[2][60] ), .QN(n1255) );
  DFFRX1 \D_cache/cache_reg[3][60]  ( .D(\D_cache/n1313 ), .CK(clk), .RN(n5748), .Q(\D_cache/cache[3][60] ), .QN(n2866) );
  DFFRX1 \D_cache/cache_reg[4][60]  ( .D(\D_cache/n1312 ), .CK(clk), .RN(n5748), .Q(\D_cache/cache[4][60] ), .QN(n1256) );
  DFFRX1 \D_cache/cache_reg[5][60]  ( .D(\D_cache/n1311 ), .CK(clk), .RN(n5748), .Q(\D_cache/cache[5][60] ), .QN(n2867) );
  DFFRX1 \D_cache/cache_reg[6][60]  ( .D(\D_cache/n1310 ), .CK(clk), .RN(n5748), .Q(\D_cache/cache[6][60] ), .QN(n1477) );
  DFFRX1 \D_cache/cache_reg[7][60]  ( .D(\D_cache/n1309 ), .CK(clk), .RN(n5748), .Q(\D_cache/cache[7][60] ), .QN(n3090) );
  DFFRX1 \D_cache/cache_reg[0][61]  ( .D(\D_cache/n1308 ), .CK(clk), .RN(n5748), .Q(\D_cache/cache[0][61] ), .QN(n1310) );
  DFFRX1 \D_cache/cache_reg[1][61]  ( .D(\D_cache/n1307 ), .CK(clk), .RN(n5748), .Q(\D_cache/cache[1][61] ), .QN(n2922) );
  DFFRX1 \D_cache/cache_reg[2][61]  ( .D(\D_cache/n1306 ), .CK(clk), .RN(n5748), .Q(\D_cache/cache[2][61] ), .QN(n1309) );
  DFFRX1 \D_cache/cache_reg[3][61]  ( .D(\D_cache/n1305 ), .CK(clk), .RN(n5749), .Q(\D_cache/cache[3][61] ), .QN(n2921) );
  DFFRX1 \D_cache/cache_reg[4][61]  ( .D(\D_cache/n1304 ), .CK(clk), .RN(n5749), .Q(\D_cache/cache[4][61] ), .QN(n1458) );
  DFFRX1 \D_cache/cache_reg[5][61]  ( .D(\D_cache/n1303 ), .CK(clk), .RN(n5749), .Q(\D_cache/cache[5][61] ), .QN(n3071) );
  DFFRX1 \D_cache/cache_reg[6][61]  ( .D(\D_cache/n1302 ), .CK(clk), .RN(n5749), .Q(\D_cache/cache[6][61] ), .QN(n1552) );
  DFFRX1 \D_cache/cache_reg[7][61]  ( .D(\D_cache/n1301 ), .CK(clk), .RN(n5749), .Q(\D_cache/cache[7][61] ), .QN(n3165) );
  DFFRX1 \D_cache/cache_reg[0][62]  ( .D(\D_cache/n1300 ), .CK(clk), .RN(n5749), .Q(\D_cache/cache[0][62] ), .QN(n459) );
  DFFRX1 \D_cache/cache_reg[1][62]  ( .D(\D_cache/n1299 ), .CK(clk), .RN(n5749), .Q(\D_cache/cache[1][62] ), .QN(n2013) );
  DFFRX1 \D_cache/cache_reg[2][62]  ( .D(\D_cache/n1298 ), .CK(clk), .RN(n5749), .Q(\D_cache/cache[2][62] ), .QN(n461) );
  DFFRX1 \D_cache/cache_reg[3][62]  ( .D(\D_cache/n1297 ), .CK(clk), .RN(n5749), .Q(\D_cache/cache[3][62] ), .QN(n2015) );
  DFFRX1 \D_cache/cache_reg[4][62]  ( .D(\D_cache/n1296 ), .CK(clk), .RN(n5749), .Q(\D_cache/cache[4][62] ), .QN(n462) );
  DFFRX1 \D_cache/cache_reg[5][62]  ( .D(\D_cache/n1295 ), .CK(clk), .RN(n5749), .Q(\D_cache/cache[5][62] ), .QN(n2016) );
  DFFRX1 \D_cache/cache_reg[6][62]  ( .D(\D_cache/n1294 ), .CK(clk), .RN(n5749), .Q(\D_cache/cache[6][62] ), .QN(n460) );
  DFFRX1 \D_cache/cache_reg[7][62]  ( .D(\D_cache/n1293 ), .CK(clk), .RN(n5750), .Q(\D_cache/cache[7][62] ), .QN(n2014) );
  DFFRX1 \D_cache/cache_reg[0][63]  ( .D(\D_cache/n1292 ), .CK(clk), .RN(n5750), .Q(\D_cache/cache[0][63] ), .QN(n1261) );
  DFFRX1 \D_cache/cache_reg[1][63]  ( .D(\D_cache/n1291 ), .CK(clk), .RN(n5750), .Q(\D_cache/cache[1][63] ), .QN(n2872) );
  DFFRX1 \D_cache/cache_reg[2][63]  ( .D(\D_cache/n1290 ), .CK(clk), .RN(n5750), .Q(\D_cache/cache[2][63] ), .QN(n1262) );
  DFFRX1 \D_cache/cache_reg[3][63]  ( .D(\D_cache/n1289 ), .CK(clk), .RN(n5750), .Q(\D_cache/cache[3][63] ), .QN(n2873) );
  DFFRX1 \D_cache/cache_reg[4][63]  ( .D(\D_cache/n1288 ), .CK(clk), .RN(n5750), .Q(\D_cache/cache[4][63] ), .QN(n1263) );
  DFFRX1 \D_cache/cache_reg[5][63]  ( .D(\D_cache/n1287 ), .CK(clk), .RN(n5750), .Q(\D_cache/cache[5][63] ), .QN(n2874) );
  DFFRX1 \D_cache/cache_reg[6][63]  ( .D(\D_cache/n1286 ), .CK(clk), .RN(n5750), .Q(\D_cache/cache[6][63] ), .QN(n1557) );
  DFFRX1 \D_cache/cache_reg[7][63]  ( .D(\D_cache/n1285 ), .CK(clk), .RN(n5750), .Q(\D_cache/cache[7][63] ), .QN(n3170) );
  DFFRX1 \D_cache/cache_reg[0][64]  ( .D(\D_cache/n1284 ), .CK(clk), .RN(n5750), .Q(\D_cache/cache[0][64] ), .QN(n1326) );
  DFFRX1 \D_cache/cache_reg[1][64]  ( .D(\D_cache/n1283 ), .CK(clk), .RN(n5750), .Q(\D_cache/cache[1][64] ), .QN(n2938) );
  DFFRX1 \D_cache/cache_reg[2][64]  ( .D(\D_cache/n1282 ), .CK(clk), .RN(n5750), .Q(\D_cache/cache[2][64] ), .QN(n1327) );
  DFFRX1 \D_cache/cache_reg[3][64]  ( .D(\D_cache/n1281 ), .CK(clk), .RN(n5751), .Q(\D_cache/cache[3][64] ), .QN(n2939) );
  DFFRX1 \D_cache/cache_reg[4][64]  ( .D(\D_cache/n1280 ), .CK(clk), .RN(n5751), .Q(\D_cache/cache[4][64] ), .QN(n2365) );
  DFFRX1 \D_cache/cache_reg[5][64]  ( .D(\D_cache/n1279 ), .CK(clk), .RN(n5751), .Q(\D_cache/cache[5][64] ), .QN(n862) );
  DFFRX1 \D_cache/cache_reg[6][64]  ( .D(\D_cache/n1278 ), .CK(clk), .RN(n5751), .Q(\D_cache/cache[6][64] ), .QN(n1484) );
  DFFRX1 \D_cache/cache_reg[7][64]  ( .D(\D_cache/n1277 ), .CK(clk), .RN(n5751), .Q(\D_cache/cache[7][64] ), .QN(n3097) );
  DFFRX1 \D_cache/cache_reg[0][65]  ( .D(\D_cache/n1276 ), .CK(clk), .RN(n5751), .Q(\D_cache/cache[0][65] ), .QN(n1565) );
  DFFRX1 \D_cache/cache_reg[1][65]  ( .D(\D_cache/n1275 ), .CK(clk), .RN(n5751), .Q(\D_cache/cache[1][65] ), .QN(n3178) );
  DFFRX1 \D_cache/cache_reg[2][65]  ( .D(\D_cache/n1274 ), .CK(clk), .RN(n5751), .Q(\D_cache/cache[2][65] ), .QN(n1305) );
  DFFRX1 \D_cache/cache_reg[3][65]  ( .D(\D_cache/n1273 ), .CK(clk), .RN(n5751), .Q(\D_cache/cache[3][65] ), .QN(n2917) );
  DFFRX1 \D_cache/cache_reg[4][65]  ( .D(\D_cache/n1272 ), .CK(clk), .RN(n5751), .Q(\D_cache/cache[4][65] ), .QN(n1566) );
  DFFRX1 \D_cache/cache_reg[5][65]  ( .D(\D_cache/n1271 ), .CK(clk), .RN(n5751), .Q(\D_cache/cache[5][65] ), .QN(n3179) );
  DFFRX1 \D_cache/cache_reg[6][65]  ( .D(\D_cache/n1270 ), .CK(clk), .RN(n5751), .Q(\D_cache/cache[6][65] ), .QN(n1449) );
  DFFRX1 \D_cache/cache_reg[7][65]  ( .D(\D_cache/n1269 ), .CK(clk), .RN(n5752), .Q(\D_cache/cache[7][65] ), .QN(n3062) );
  DFFRX1 \D_cache/cache_reg[0][66]  ( .D(\D_cache/n1268 ), .CK(clk), .RN(n5752), .Q(\D_cache/cache[0][66] ), .QN(n1469) );
  DFFRX1 \D_cache/cache_reg[1][66]  ( .D(\D_cache/n1267 ), .CK(clk), .RN(n5752), .Q(\D_cache/cache[1][66] ), .QN(n3082) );
  DFFRX1 \D_cache/cache_reg[2][66]  ( .D(\D_cache/n1266 ), .CK(clk), .RN(n5752), .Q(\D_cache/cache[2][66] ), .QN(n1251) );
  DFFRX1 \D_cache/cache_reg[3][66]  ( .D(\D_cache/n1265 ), .CK(clk), .RN(n5752), .Q(\D_cache/cache[3][66] ), .QN(n2862) );
  DFFRX1 \D_cache/cache_reg[4][66]  ( .D(\D_cache/n1264 ), .CK(clk), .RN(n5752), .Q(\D_cache/cache[4][66] ), .QN(n1470) );
  DFFRX1 \D_cache/cache_reg[5][66]  ( .D(\D_cache/n1263 ), .CK(clk), .RN(n5752), .Q(\D_cache/cache[5][66] ), .QN(n3083) );
  DFFRX1 \D_cache/cache_reg[6][66]  ( .D(\D_cache/n1262 ), .CK(clk), .RN(n5752), .Q(\D_cache/cache[6][66] ), .QN(n1514) );
  DFFRX1 \D_cache/cache_reg[7][66]  ( .D(\D_cache/n1261 ), .CK(clk), .RN(n5752), .Q(\D_cache/cache[7][66] ), .QN(n3127) );
  DFFRX1 \D_cache/cache_reg[0][67]  ( .D(\D_cache/n1260 ), .CK(clk), .RN(n5752), .Q(\D_cache/cache[0][67] ), .QN(n1267) );
  DFFRX1 \D_cache/cache_reg[1][67]  ( .D(\D_cache/n1259 ), .CK(clk), .RN(n5752), .Q(\D_cache/cache[1][67] ), .QN(n2878) );
  DFFRX1 \D_cache/cache_reg[2][67]  ( .D(\D_cache/n1258 ), .CK(clk), .RN(n5752), .Q(\D_cache/cache[2][67] ), .QN(n1268) );
  DFFRX1 \D_cache/cache_reg[3][67]  ( .D(\D_cache/n1257 ), .CK(clk), .RN(n5753), .Q(\D_cache/cache[3][67] ), .QN(n2879) );
  DFFRX1 \D_cache/cache_reg[4][67]  ( .D(\D_cache/n1256 ), .CK(clk), .RN(n5753), .Q(\D_cache/cache[4][67] ), .QN(n942) );
  DFFRX1 \D_cache/cache_reg[5][67]  ( .D(\D_cache/n1255 ), .CK(clk), .RN(n5753), .Q(\D_cache/cache[5][67] ), .QN(n2467) );
  DFFRX1 \D_cache/cache_reg[6][67]  ( .D(\D_cache/n1254 ), .CK(clk), .RN(n5753), .Q(\D_cache/cache[6][67] ), .QN(n1518) );
  DFFRX1 \D_cache/cache_reg[7][67]  ( .D(\D_cache/n1253 ), .CK(clk), .RN(n5753), .Q(\D_cache/cache[7][67] ), .QN(n3131) );
  DFFRX1 \D_cache/cache_reg[0][68]  ( .D(\D_cache/n1252 ), .CK(clk), .RN(n5753), .Q(\D_cache/cache[0][68] ), .QN(n1294) );
  DFFRX1 \D_cache/cache_reg[1][68]  ( .D(\D_cache/n1251 ), .CK(clk), .RN(n5753), .Q(\D_cache/cache[1][68] ), .QN(n2906) );
  DFFRX1 \D_cache/cache_reg[2][68]  ( .D(\D_cache/n1250 ), .CK(clk), .RN(n5753), .Q(\D_cache/cache[2][68] ), .QN(n1295) );
  DFFRX1 \D_cache/cache_reg[3][68]  ( .D(\D_cache/n1249 ), .CK(clk), .RN(n5753), .Q(\D_cache/cache[3][68] ), .QN(n2907) );
  DFFRX1 \D_cache/cache_reg[4][68]  ( .D(\D_cache/n1248 ), .CK(clk), .RN(n5753), .Q(\D_cache/cache[4][68] ), .QN(n2382) );
  DFFRX1 \D_cache/cache_reg[5][68]  ( .D(\D_cache/n1247 ), .CK(clk), .RN(n5753), .Q(\D_cache/cache[5][68] ), .QN(n877) );
  DFFRX1 \D_cache/cache_reg[6][68]  ( .D(\D_cache/n1246 ), .CK(clk), .RN(n5753), .Q(\D_cache/cache[6][68] ), .QN(n1541) );
  DFFRX1 \D_cache/cache_reg[7][68]  ( .D(\D_cache/n1245 ), .CK(clk), .RN(n5754), .Q(\D_cache/cache[7][68] ), .QN(n3154) );
  DFFRX1 \D_cache/cache_reg[0][69]  ( .D(\D_cache/n1244 ), .CK(clk), .RN(n5754), .Q(\D_cache/cache[0][69] ), .QN(n1272) );
  DFFRX1 \D_cache/cache_reg[1][69]  ( .D(\D_cache/n1243 ), .CK(clk), .RN(n5754), .Q(\D_cache/cache[1][69] ), .QN(n2883) );
  DFFRX1 \D_cache/cache_reg[2][69]  ( .D(\D_cache/n1242 ), .CK(clk), .RN(n5754), .Q(\D_cache/cache[2][69] ), .QN(n1273) );
  DFFRX1 \D_cache/cache_reg[3][69]  ( .D(\D_cache/n1241 ), .CK(clk), .RN(n5754), .Q(\D_cache/cache[3][69] ), .QN(n2884) );
  DFFRX1 \D_cache/cache_reg[4][69]  ( .D(\D_cache/n1240 ), .CK(clk), .RN(n5754), .Q(\D_cache/cache[4][69] ), .QN(n1228) );
  DFFRX1 \D_cache/cache_reg[5][69]  ( .D(\D_cache/n1239 ), .CK(clk), .RN(n5754), .Q(\D_cache/cache[5][69] ), .QN(n2885) );
  DFFRX1 \D_cache/cache_reg[6][69]  ( .D(\D_cache/n1238 ), .CK(clk), .RN(n5754), .Q(\D_cache/cache[6][69] ), .QN(n1547) );
  DFFRX1 \D_cache/cache_reg[7][69]  ( .D(\D_cache/n1237 ), .CK(clk), .RN(n5754), .Q(\D_cache/cache[7][69] ), .QN(n3160) );
  DFFRX1 \D_cache/cache_reg[0][70]  ( .D(\D_cache/n1236 ), .CK(clk), .RN(n5754), .Q(\D_cache/cache[0][70] ), .QN(n1348) );
  DFFRX1 \D_cache/cache_reg[1][70]  ( .D(\D_cache/n1235 ), .CK(clk), .RN(n5754), .Q(\D_cache/cache[1][70] ), .QN(n2960) );
  DFFRX1 \D_cache/cache_reg[2][70]  ( .D(\D_cache/n1234 ), .CK(clk), .RN(n5754), .Q(\D_cache/cache[2][70] ), .QN(n1346) );
  DFFRX1 \D_cache/cache_reg[3][70]  ( .D(\D_cache/n1233 ), .CK(clk), .RN(n5755), .Q(\D_cache/cache[3][70] ), .QN(n2958) );
  DFFRX1 \D_cache/cache_reg[4][70]  ( .D(\D_cache/n1232 ), .CK(clk), .RN(n5755), .Q(\D_cache/cache[4][70] ), .QN(n1347) );
  DFFRX1 \D_cache/cache_reg[5][70]  ( .D(\D_cache/n1231 ), .CK(clk), .RN(n5755), .Q(\D_cache/cache[5][70] ), .QN(n2959) );
  DFFRX1 \D_cache/cache_reg[6][70]  ( .D(\D_cache/n1230 ), .CK(clk), .RN(n5755), .Q(\D_cache/cache[6][70] ), .QN(n1555) );
  DFFRX1 \D_cache/cache_reg[7][70]  ( .D(\D_cache/n1229 ), .CK(clk), .RN(n5755), .Q(\D_cache/cache[7][70] ), .QN(n3168) );
  DFFRX1 \D_cache/cache_reg[0][71]  ( .D(\D_cache/n1228 ), .CK(clk), .RN(n5755), .Q(\D_cache/cache[0][71] ), .QN(n1341) );
  DFFRX1 \D_cache/cache_reg[1][71]  ( .D(\D_cache/n1227 ), .CK(clk), .RN(n5755), .Q(\D_cache/cache[1][71] ), .QN(n2953) );
  DFFRX1 \D_cache/cache_reg[2][71]  ( .D(\D_cache/n1226 ), .CK(clk), .RN(n5755), .Q(\D_cache/cache[2][71] ), .QN(n1340) );
  DFFRX1 \D_cache/cache_reg[3][71]  ( .D(\D_cache/n1225 ), .CK(clk), .RN(n5755), .Q(\D_cache/cache[3][71] ), .QN(n2952) );
  DFFRX1 \D_cache/cache_reg[4][71]  ( .D(\D_cache/n1224 ), .CK(clk), .RN(n5755), .Q(\D_cache/cache[4][71] ), .QN(n2386) );
  DFFRX1 \D_cache/cache_reg[5][71]  ( .D(\D_cache/n1223 ), .CK(clk), .RN(n5755), .Q(\D_cache/cache[5][71] ), .QN(n881) );
  DFFRX1 \D_cache/cache_reg[6][71]  ( .D(\D_cache/n1222 ), .CK(clk), .RN(n5755), .Q(\D_cache/cache[6][71] ), .QN(n1554) );
  DFFRX1 \D_cache/cache_reg[7][71]  ( .D(\D_cache/n1221 ), .CK(clk), .RN(n5756), .Q(\D_cache/cache[7][71] ), .QN(n3167) );
  DFFRX1 \D_cache/cache_reg[0][72]  ( .D(\D_cache/n1220 ), .CK(clk), .RN(n5756), .Q(\D_cache/cache[0][72] ), .QN(n1506) );
  DFFRX1 \D_cache/cache_reg[1][72]  ( .D(\D_cache/n1219 ), .CK(clk), .RN(n5756), .Q(\D_cache/cache[1][72] ), .QN(n3119) );
  DFFRX1 \D_cache/cache_reg[2][72]  ( .D(\D_cache/n1218 ), .CK(clk), .RN(n5756), .Q(\D_cache/cache[2][72] ), .QN(n1504) );
  DFFRX1 \D_cache/cache_reg[3][72]  ( .D(\D_cache/n1217 ), .CK(clk), .RN(n5756), .Q(\D_cache/cache[3][72] ), .QN(n3117) );
  DFFRX1 \D_cache/cache_reg[4][72]  ( .D(\D_cache/n1216 ), .CK(clk), .RN(n5756), .Q(\D_cache/cache[4][72] ), .QN(n1505) );
  DFFRX1 \D_cache/cache_reg[5][72]  ( .D(\D_cache/n1215 ), .CK(clk), .RN(n5756), .Q(\D_cache/cache[5][72] ), .QN(n3118) );
  DFFRX1 \D_cache/cache_reg[6][72]  ( .D(\D_cache/n1214 ), .CK(clk), .RN(n5756), .Q(\D_cache/cache[6][72] ), .QN(n1548) );
  DFFRX1 \D_cache/cache_reg[7][72]  ( .D(\D_cache/n1213 ), .CK(clk), .RN(n5756), .Q(\D_cache/cache[7][72] ), .QN(n3161) );
  DFFRX1 \D_cache/cache_reg[0][73]  ( .D(\D_cache/n1212 ), .CK(clk), .RN(n5756), .Q(\D_cache/cache[0][73] ), .QN(n1354) );
  DFFRX1 \D_cache/cache_reg[1][73]  ( .D(\D_cache/n1211 ), .CK(clk), .RN(n5756), .Q(\D_cache/cache[1][73] ), .QN(n2967) );
  DFFRX1 \D_cache/cache_reg[2][73]  ( .D(\D_cache/n1210 ), .CK(clk), .RN(n5756), .Q(\D_cache/cache[2][73] ), .QN(n1353) );
  DFFRX1 \D_cache/cache_reg[3][73]  ( .D(\D_cache/n1209 ), .CK(clk), .RN(n5757), .Q(\D_cache/cache[3][73] ), .QN(n2966) );
  DFFRX1 \D_cache/cache_reg[4][73]  ( .D(\D_cache/n1208 ), .CK(clk), .RN(n5757), .Q(\D_cache/cache[4][73] ), .QN(n921) );
  DFFRX1 \D_cache/cache_reg[5][73]  ( .D(\D_cache/n1207 ), .CK(clk), .RN(n5757), .Q(\D_cache/cache[5][73] ), .QN(n2458) );
  DFFRX1 \D_cache/cache_reg[6][73]  ( .D(\D_cache/n1206 ), .CK(clk), .RN(n5757), .Q(\D_cache/cache[6][73] ), .QN(n1454) );
  DFFRX1 \D_cache/cache_reg[7][73]  ( .D(\D_cache/n1205 ), .CK(clk), .RN(n5757), .Q(\D_cache/cache[7][73] ), .QN(n3067) );
  DFFRX1 \D_cache/cache_reg[0][74]  ( .D(\D_cache/n1204 ), .CK(clk), .RN(n5757), .Q(\D_cache/cache[0][74] ), .QN(n1279) );
  DFFRX1 \D_cache/cache_reg[1][74]  ( .D(\D_cache/n1203 ), .CK(clk), .RN(n5757), .Q(\D_cache/cache[1][74] ), .QN(n2891) );
  DFFRX1 \D_cache/cache_reg[2][74]  ( .D(\D_cache/n1202 ), .CK(clk), .RN(n5757), .Q(\D_cache/cache[2][74] ), .QN(n1280) );
  DFFRX1 \D_cache/cache_reg[3][74]  ( .D(\D_cache/n1201 ), .CK(clk), .RN(n5757), .Q(\D_cache/cache[3][74] ), .QN(n2892) );
  DFFRX1 \D_cache/cache_reg[4][74]  ( .D(\D_cache/n1200 ), .CK(clk), .RN(n5757), .Q(\D_cache/cache[4][74] ), .QN(n1281) );
  DFFRX1 \D_cache/cache_reg[5][74]  ( .D(\D_cache/n1199 ), .CK(clk), .RN(n5757), .Q(\D_cache/cache[5][74] ), .QN(n2893) );
  DFFRX1 \D_cache/cache_reg[6][74]  ( .D(\D_cache/n1198 ), .CK(clk), .RN(n5757), .Q(\D_cache/cache[6][74] ), .QN(n1544) );
  DFFRX1 \D_cache/cache_reg[7][74]  ( .D(\D_cache/n1197 ), .CK(clk), .RN(n5758), .Q(\D_cache/cache[7][74] ), .QN(n3157) );
  DFFRX1 \D_cache/cache_reg[0][75]  ( .D(\D_cache/n1196 ), .CK(clk), .RN(n5758), .Q(\D_cache/cache[0][75] ), .QN(n2376) );
  DFFRX1 \D_cache/cache_reg[1][75]  ( .D(\D_cache/n1195 ), .CK(clk), .RN(n5758), .Q(\D_cache/cache[1][75] ), .QN(n872) );
  DFFRX1 \D_cache/cache_reg[2][75]  ( .D(\D_cache/n1194 ), .CK(clk), .RN(n5758), .Q(\D_cache/cache[2][75] ), .QN(n1282) );
  DFFRX1 \D_cache/cache_reg[3][75]  ( .D(\D_cache/n1193 ), .CK(clk), .RN(n5758), .Q(\D_cache/cache[3][75] ), .QN(n2894) );
  DFFRX1 \D_cache/cache_reg[4][75]  ( .D(\D_cache/n1192 ), .CK(clk), .RN(n5758), .Q(\D_cache/cache[4][75] ), .QN(n2396) );
  DFFRX1 \D_cache/cache_reg[5][75]  ( .D(\D_cache/n1191 ), .CK(clk), .RN(n5758), .Q(\D_cache/cache[5][75] ), .QN(n891) );
  DFFRX1 \D_cache/cache_reg[6][75]  ( .D(\D_cache/n1190 ), .CK(clk), .RN(n5758), .Q(\D_cache/cache[6][75] ), .QN(n1475) );
  DFFRX1 \D_cache/cache_reg[7][75]  ( .D(\D_cache/n1189 ), .CK(clk), .RN(n5758), .Q(\D_cache/cache[7][75] ), .QN(n3088) );
  DFFRX1 \D_cache/cache_reg[0][76]  ( .D(\D_cache/n1188 ), .CK(clk), .RN(n5758), .Q(\D_cache/cache[0][76] ), .QN(n1356) );
  DFFRX1 \D_cache/cache_reg[1][76]  ( .D(\D_cache/n1187 ), .CK(clk), .RN(n5758), .Q(\D_cache/cache[1][76] ), .QN(n2969) );
  DFFRX1 \D_cache/cache_reg[2][76]  ( .D(\D_cache/n1186 ), .CK(clk), .RN(n5758), .Q(\D_cache/cache[2][76] ), .QN(n1355) );
  DFFRX1 \D_cache/cache_reg[3][76]  ( .D(\D_cache/n1185 ), .CK(clk), .RN(n5759), .Q(\D_cache/cache[3][76] ), .QN(n2968) );
  DFFRX1 \D_cache/cache_reg[4][76]  ( .D(\D_cache/n1184 ), .CK(clk), .RN(n5759), .Q(\D_cache/cache[4][76] ), .QN(n2366) );
  DFFRX1 \D_cache/cache_reg[5][76]  ( .D(\D_cache/n1183 ), .CK(clk), .RN(n5759), .Q(\D_cache/cache[5][76] ), .QN(n863) );
  DFFRX1 \D_cache/cache_reg[6][76]  ( .D(\D_cache/n1182 ), .CK(clk), .RN(n5759), .Q(\D_cache/cache[6][76] ), .QN(n1540) );
  DFFRX1 \D_cache/cache_reg[7][76]  ( .D(\D_cache/n1181 ), .CK(clk), .RN(n5759), .Q(\D_cache/cache[7][76] ), .QN(n3153) );
  DFFRX1 \D_cache/cache_reg[0][77]  ( .D(\D_cache/n1180 ), .CK(clk), .RN(n5759), .Q(\D_cache/cache[0][77] ), .QN(n1537) );
  DFFRX1 \D_cache/cache_reg[1][77]  ( .D(\D_cache/n1179 ), .CK(clk), .RN(n5759), .Q(\D_cache/cache[1][77] ), .QN(n3150) );
  DFFRX1 \D_cache/cache_reg[2][77]  ( .D(\D_cache/n1178 ), .CK(clk), .RN(n5759), .Q(\D_cache/cache[2][77] ), .QN(n961) );
  DFFRX1 \D_cache/cache_reg[3][77]  ( .D(\D_cache/n1177 ), .CK(clk), .RN(n5759), .Q(\D_cache/cache[3][77] ), .QN(n2486) );
  DFFRX1 \D_cache/cache_reg[4][77]  ( .D(\D_cache/n1176 ), .CK(clk), .RN(n5759), .Q(\D_cache/cache[4][77] ), .QN(n962) );
  DFFRX1 \D_cache/cache_reg[5][77]  ( .D(\D_cache/n1175 ), .CK(clk), .RN(n5759), .Q(\D_cache/cache[5][77] ), .QN(n2487) );
  DFFRX1 \D_cache/cache_reg[6][77]  ( .D(\D_cache/n1174 ), .CK(clk), .RN(n5759), .Q(\D_cache/cache[6][77] ), .QN(n1428) );
  DFFRX1 \D_cache/cache_reg[7][77]  ( .D(\D_cache/n1173 ), .CK(clk), .RN(n5760), .Q(\D_cache/cache[7][77] ), .QN(n3041) );
  DFFRX1 \D_cache/cache_reg[0][78]  ( .D(\D_cache/n1172 ), .CK(clk), .RN(n5760), .Q(\D_cache/cache[0][78] ), .QN(n1531) );
  DFFRX1 \D_cache/cache_reg[1][78]  ( .D(\D_cache/n1171 ), .CK(clk), .RN(n5760), .Q(\D_cache/cache[1][78] ), .QN(n3144) );
  DFFRX1 \D_cache/cache_reg[2][78]  ( .D(\D_cache/n1170 ), .CK(clk), .RN(n5760), .Q(\D_cache/cache[2][78] ), .QN(n963) );
  DFFRX1 \D_cache/cache_reg[3][78]  ( .D(\D_cache/n1169 ), .CK(clk), .RN(n5760), .Q(\D_cache/cache[3][78] ), .QN(n2488) );
  DFFRX1 \D_cache/cache_reg[4][78]  ( .D(\D_cache/n1168 ), .CK(clk), .RN(n5760), .Q(\D_cache/cache[4][78] ), .QN(n964) );
  DFFRX1 \D_cache/cache_reg[5][78]  ( .D(\D_cache/n1167 ), .CK(clk), .RN(n5760), .Q(\D_cache/cache[5][78] ), .QN(n2489) );
  DFFRX1 \D_cache/cache_reg[6][78]  ( .D(\D_cache/n1166 ), .CK(clk), .RN(n5760), .Q(\D_cache/cache[6][78] ), .QN(n1431) );
  DFFRX1 \D_cache/cache_reg[7][78]  ( .D(\D_cache/n1165 ), .CK(clk), .RN(n5760), .Q(\D_cache/cache[7][78] ), .QN(n3044) );
  DFFRX1 \D_cache/cache_reg[0][79]  ( .D(\D_cache/n1164 ), .CK(clk), .RN(n5760), .Q(\D_cache/cache[0][79] ), .QN(n2373) );
  DFFRX1 \D_cache/cache_reg[1][79]  ( .D(\D_cache/n1163 ), .CK(clk), .RN(n5760), .Q(\D_cache/cache[1][79] ), .QN(n869) );
  DFFRX1 \D_cache/cache_reg[2][79]  ( .D(\D_cache/n1162 ), .CK(clk), .RN(n5760), .Q(\D_cache/cache[2][79] ), .QN(n1429) );
  DFFRX1 \D_cache/cache_reg[3][79]  ( .D(\D_cache/n1161 ), .CK(clk), .RN(n5761), .Q(\D_cache/cache[3][79] ), .QN(n3042) );
  DFFRX1 \D_cache/cache_reg[4][79]  ( .D(\D_cache/n1160 ), .CK(clk), .RN(n5761), .Q(\D_cache/cache[4][79] ), .QN(n2393) );
  DFFRX1 \D_cache/cache_reg[5][79]  ( .D(\D_cache/n1159 ), .CK(clk), .RN(n5761), .Q(\D_cache/cache[5][79] ), .QN(n888) );
  DFFRX1 \D_cache/cache_reg[6][79]  ( .D(\D_cache/n1158 ), .CK(clk), .RN(n5761), .Q(\D_cache/cache[6][79] ), .QN(n1430) );
  DFFRX1 \D_cache/cache_reg[7][79]  ( .D(\D_cache/n1157 ), .CK(clk), .RN(n5761), .Q(\D_cache/cache[7][79] ), .QN(n3043) );
  DFFRX1 \D_cache/cache_reg[0][80]  ( .D(\D_cache/n1156 ), .CK(clk), .RN(n5761), .Q(\D_cache/cache[0][80] ), .QN(n1284) );
  DFFRX1 \D_cache/cache_reg[1][80]  ( .D(\D_cache/n1155 ), .CK(clk), .RN(n5761), .Q(\D_cache/cache[1][80] ), .QN(n2896) );
  DFFRX1 \D_cache/cache_reg[2][80]  ( .D(\D_cache/n1154 ), .CK(clk), .RN(n5761), .Q(\D_cache/cache[2][80] ), .QN(n1285) );
  DFFRX1 \D_cache/cache_reg[3][80]  ( .D(\D_cache/n1153 ), .CK(clk), .RN(n5761), .Q(\D_cache/cache[3][80] ), .QN(n2897) );
  DFFRX1 \D_cache/cache_reg[4][80]  ( .D(\D_cache/n1152 ), .CK(clk), .RN(n5761), .Q(\D_cache/cache[4][80] ), .QN(n2412) );
  DFFRX1 \D_cache/cache_reg[5][80]  ( .D(\D_cache/n1151 ), .CK(clk), .RN(n5761), .Q(\D_cache/cache[5][80] ), .QN(n904) );
  DFFRX1 \D_cache/cache_reg[6][80]  ( .D(\D_cache/n1150 ), .CK(clk), .RN(n5761), .Q(\D_cache/cache[6][80] ), .QN(n1520) );
  DFFRX1 \D_cache/cache_reg[7][80]  ( .D(\D_cache/n1149 ), .CK(clk), .RN(n5762), .Q(\D_cache/cache[7][80] ), .QN(n3133) );
  DFFRX1 \D_cache/cache_reg[0][81]  ( .D(\D_cache/n1148 ), .CK(clk), .RN(n5762), .Q(\D_cache/cache[0][81] ), .QN(n1560) );
  DFFRX1 \D_cache/cache_reg[1][81]  ( .D(\D_cache/n1147 ), .CK(clk), .RN(n5762), .Q(\D_cache/cache[1][81] ), .QN(n3173) );
  DFFRX1 \D_cache/cache_reg[2][81]  ( .D(\D_cache/n1146 ), .CK(clk), .RN(n5762), .Q(\D_cache/cache[2][81] ), .QN(n951) );
  DFFRX1 \D_cache/cache_reg[3][81]  ( .D(\D_cache/n1145 ), .CK(clk), .RN(n5762), .Q(\D_cache/cache[3][81] ), .QN(n2476) );
  DFFRX1 \D_cache/cache_reg[4][81]  ( .D(\D_cache/n1144 ), .CK(clk), .RN(n5762), .Q(\D_cache/cache[4][81] ), .QN(n1559) );
  DFFRX1 \D_cache/cache_reg[5][81]  ( .D(\D_cache/n1143 ), .CK(clk), .RN(n5762), .Q(\D_cache/cache[5][81] ), .QN(n3172) );
  DFFRX1 \D_cache/cache_reg[6][81]  ( .D(\D_cache/n1142 ), .CK(clk), .RN(n5762), .Q(\D_cache/cache[6][81] ), .QN(n1236) );
  DFFRX1 \D_cache/cache_reg[7][81]  ( .D(\D_cache/n1141 ), .CK(clk), .RN(n5762), .Q(\D_cache/cache[7][81] ), .QN(n2841) );
  DFFRX1 \D_cache/cache_reg[0][82]  ( .D(\D_cache/n1140 ), .CK(clk), .RN(n5762), .Q(\D_cache/cache[0][82] ), .QN(n954) );
  DFFRX1 \D_cache/cache_reg[1][82]  ( .D(\D_cache/n1139 ), .CK(clk), .RN(n5762), .Q(\D_cache/cache[1][82] ), .QN(n2479) );
  DFFRX1 \D_cache/cache_reg[2][82]  ( .D(\D_cache/n1138 ), .CK(clk), .RN(n5762), .Q(\D_cache/cache[2][82] ), .QN(n955) );
  DFFRX1 \D_cache/cache_reg[3][82]  ( .D(\D_cache/n1137 ), .CK(clk), .RN(n5763), .Q(\D_cache/cache[3][82] ), .QN(n2480) );
  DFFRX1 \D_cache/cache_reg[4][82]  ( .D(\D_cache/n1136 ), .CK(clk), .RN(n5763), .Q(\D_cache/cache[4][82] ), .QN(n1568) );
  DFFRX1 \D_cache/cache_reg[5][82]  ( .D(\D_cache/n1135 ), .CK(clk), .RN(n5763), .Q(\D_cache/cache[5][82] ), .QN(n3181) );
  DFFRX1 \D_cache/cache_reg[6][82]  ( .D(\D_cache/n1134 ), .CK(clk), .RN(n5763), .Q(\D_cache/cache[6][82] ), .QN(n2400) );
  DFFRX1 \D_cache/cache_reg[7][82]  ( .D(\D_cache/n1133 ), .CK(clk), .RN(n5763), .Q(\D_cache/cache[7][82] ), .QN(n895) );
  DFFRX1 \D_cache/cache_reg[0][83]  ( .D(\D_cache/n1132 ), .CK(clk), .RN(n5763), .Q(\D_cache/cache[0][83] ), .QN(n1460) );
  DFFRX1 \D_cache/cache_reg[1][83]  ( .D(\D_cache/n1131 ), .CK(clk), .RN(n5763), .Q(\D_cache/cache[1][83] ), .QN(n3073) );
  DFFRX1 \D_cache/cache_reg[2][83]  ( .D(\D_cache/n1130 ), .CK(clk), .RN(n5763), .Q(\D_cache/cache[2][83] ), .QN(n1303) );
  DFFRX1 \D_cache/cache_reg[3][83]  ( .D(\D_cache/n1129 ), .CK(clk), .RN(n5763), .Q(\D_cache/cache[3][83] ), .QN(n2915) );
  DFFRX1 \D_cache/cache_reg[4][83]  ( .D(\D_cache/n1128 ), .CK(clk), .RN(n5763), .Q(\D_cache/cache[4][83] ), .QN(n944) );
  DFFRX1 \D_cache/cache_reg[5][83]  ( .D(\D_cache/n1127 ), .CK(clk), .RN(n5763), .Q(\D_cache/cache[5][83] ), .QN(n2469) );
  DFFRX1 \D_cache/cache_reg[6][83]  ( .D(\D_cache/n1126 ), .CK(clk), .RN(n5763), .Q(\D_cache/cache[6][83] ), .QN(n1527) );
  DFFRX1 \D_cache/cache_reg[7][83]  ( .D(\D_cache/n1125 ), .CK(clk), .RN(n5764), .Q(\D_cache/cache[7][83] ), .QN(n3140) );
  DFFRX1 \D_cache/cache_reg[0][84]  ( .D(\D_cache/n1124 ), .CK(clk), .RN(n5764), .Q(\D_cache/cache[0][84] ), .QN(n1465) );
  DFFRX1 \D_cache/cache_reg[1][84]  ( .D(\D_cache/n1123 ), .CK(clk), .RN(n5764), .Q(\D_cache/cache[1][84] ), .QN(n3078) );
  DFFRX1 \D_cache/cache_reg[2][84]  ( .D(\D_cache/n1122 ), .CK(clk), .RN(n5764), .Q(\D_cache/cache[2][84] ), .QN(n2359) );
  DFFRX1 \D_cache/cache_reg[3][84]  ( .D(\D_cache/n1121 ), .CK(clk), .RN(n5764), .Q(\D_cache/cache[3][84] ), .QN(n856) );
  DFFRX1 \D_cache/cache_reg[4][84]  ( .D(\D_cache/n1120 ), .CK(clk), .RN(n5764), .Q(\D_cache/cache[4][84] ), .QN(n1315) );
  DFFRX1 \D_cache/cache_reg[5][84]  ( .D(\D_cache/n1119 ), .CK(clk), .RN(n5764), .Q(\D_cache/cache[5][84] ), .QN(n2927) );
  DFFRX1 \D_cache/cache_reg[6][84]  ( .D(\D_cache/n1118 ), .CK(clk), .RN(n5764), .Q(\D_cache/cache[6][84] ), .QN(n930) );
  DFFRX1 \D_cache/cache_reg[7][84]  ( .D(\D_cache/n1117 ), .CK(clk), .RN(n5764), .Q(\D_cache/cache[7][84] ), .QN(n2454) );
  DFFRX1 \D_cache/cache_reg[0][85]  ( .D(\D_cache/n1116 ), .CK(clk), .RN(n5764), .Q(\D_cache/cache[0][85] ), .QN(n1320) );
  DFFRX1 \D_cache/cache_reg[1][85]  ( .D(\D_cache/n1115 ), .CK(clk), .RN(n5764), .Q(\D_cache/cache[1][85] ), .QN(n2932) );
  DFFRX1 \D_cache/cache_reg[2][85]  ( .D(\D_cache/n1114 ), .CK(clk), .RN(n5764), .Q(\D_cache/cache[2][85] ), .QN(n1319) );
  DFFRX1 \D_cache/cache_reg[3][85]  ( .D(\D_cache/n1113 ), .CK(clk), .RN(n5765), .Q(\D_cache/cache[3][85] ), .QN(n2931) );
  DFFRX1 \D_cache/cache_reg[4][85]  ( .D(\D_cache/n1112 ), .CK(clk), .RN(n5765), .Q(\D_cache/cache[4][85] ), .QN(n2411) );
  DFFRX1 \D_cache/cache_reg[5][85]  ( .D(\D_cache/n1111 ), .CK(clk), .RN(n5765), .Q(\D_cache/cache[5][85] ), .QN(n383) );
  DFFRX1 \D_cache/cache_reg[6][85]  ( .D(\D_cache/n1110 ), .CK(clk), .RN(n5765), .Q(\D_cache/cache[6][85] ), .QN(n1524) );
  DFFRX1 \D_cache/cache_reg[7][85]  ( .D(\D_cache/n1109 ), .CK(clk), .RN(n5765), .Q(\D_cache/cache[7][85] ), .QN(n3137) );
  DFFRX1 \D_cache/cache_reg[0][86]  ( .D(\D_cache/n1108 ), .CK(clk), .RN(n5765), .Q(\D_cache/cache[0][86] ), .QN(n1323) );
  DFFRX1 \D_cache/cache_reg[1][86]  ( .D(\D_cache/n1107 ), .CK(clk), .RN(n5765), .Q(\D_cache/cache[1][86] ), .QN(n2935) );
  DFFRX1 \D_cache/cache_reg[2][86]  ( .D(\D_cache/n1106 ), .CK(clk), .RN(n5765), .Q(\D_cache/cache[2][86] ), .QN(n1321) );
  DFFRX1 \D_cache/cache_reg[3][86]  ( .D(\D_cache/n1105 ), .CK(clk), .RN(n5765), .Q(\D_cache/cache[3][86] ), .QN(n2933) );
  DFFRX1 \D_cache/cache_reg[4][86]  ( .D(\D_cache/n1104 ), .CK(clk), .RN(n5765), .Q(\D_cache/cache[4][86] ), .QN(n1322) );
  DFFRX1 \D_cache/cache_reg[5][86]  ( .D(\D_cache/n1103 ), .CK(clk), .RN(n5765), .Q(\D_cache/cache[5][86] ), .QN(n2934) );
  DFFRX1 \D_cache/cache_reg[6][86]  ( .D(\D_cache/n1102 ), .CK(clk), .RN(n5765), .Q(\D_cache/cache[6][86] ), .QN(n1530) );
  DFFRX1 \D_cache/cache_reg[7][86]  ( .D(\D_cache/n1101 ), .CK(clk), .RN(n5766), .Q(\D_cache/cache[7][86] ), .QN(n3143) );
  DFFRX1 \D_cache/cache_reg[0][87]  ( .D(\D_cache/n1100 ), .CK(clk), .RN(n5766), .Q(\D_cache/cache[0][87] ), .QN(n2408) );
  DFFRX1 \D_cache/cache_reg[1][87]  ( .D(\D_cache/n1099 ), .CK(clk), .RN(n5766), .Q(\D_cache/cache[1][87] ), .QN(n902) );
  DFFRX1 \D_cache/cache_reg[2][87]  ( .D(\D_cache/n1098 ), .CK(clk), .RN(n5766), .Q(\D_cache/cache[2][87] ), .QN(n1259) );
  DFFRX1 \D_cache/cache_reg[3][87]  ( .D(\D_cache/n1097 ), .CK(clk), .RN(n5766), .Q(\D_cache/cache[3][87] ), .QN(n2870) );
  DFFRX1 \D_cache/cache_reg[4][87]  ( .D(\D_cache/n1096 ), .CK(clk), .RN(n5766), .Q(\D_cache/cache[4][87] ), .QN(n1260) );
  DFFRX1 \D_cache/cache_reg[5][87]  ( .D(\D_cache/n1095 ), .CK(clk), .RN(n5766), .Q(\D_cache/cache[5][87] ), .QN(n2871) );
  DFFRX1 \D_cache/cache_reg[6][87]  ( .D(\D_cache/n1094 ), .CK(clk), .RN(n5766), .Q(\D_cache/cache[6][87] ), .QN(n1519) );
  DFFRX1 \D_cache/cache_reg[7][87]  ( .D(\D_cache/n1093 ), .CK(clk), .RN(n5766), .Q(\D_cache/cache[7][87] ), .QN(n3132) );
  DFFRX1 \D_cache/cache_reg[0][88]  ( .D(\D_cache/n1092 ), .CK(clk), .RN(n5766), .Q(\D_cache/cache[0][88] ), .QN(n1257) );
  DFFRX1 \D_cache/cache_reg[1][88]  ( .D(\D_cache/n1091 ), .CK(clk), .RN(n5766), .Q(\D_cache/cache[1][88] ), .QN(n2868) );
  DFFRX1 \D_cache/cache_reg[2][88]  ( .D(\D_cache/n1090 ), .CK(clk), .RN(n5766), .Q(\D_cache/cache[2][88] ), .QN(n1258) );
  DFFRX1 \D_cache/cache_reg[3][88]  ( .D(\D_cache/n1089 ), .CK(clk), .RN(n5767), .Q(\D_cache/cache[3][88] ), .QN(n2869) );
  DFFRX1 \D_cache/cache_reg[4][88]  ( .D(\D_cache/n1088 ), .CK(clk), .RN(n5767), .Q(\D_cache/cache[4][88] ), .QN(n2813) );
  DFFRX1 \D_cache/cache_reg[5][88]  ( .D(\D_cache/n1087 ), .CK(clk), .RN(n5767), .Q(\D_cache/cache[5][88] ), .QN(n821) );
  DFFRX1 \D_cache/cache_reg[6][88]  ( .D(\D_cache/n1086 ), .CK(clk), .RN(n5767), .Q(\D_cache/cache[6][88] ), .QN(n1516) );
  DFFRX1 \D_cache/cache_reg[7][88]  ( .D(\D_cache/n1085 ), .CK(clk), .RN(n5767), .Q(\D_cache/cache[7][88] ), .QN(n3129) );
  DFFRX1 \D_cache/cache_reg[0][89]  ( .D(\D_cache/n1084 ), .CK(clk), .RN(n5767), .Q(\D_cache/cache[0][89] ), .QN(n1336) );
  DFFRX1 \D_cache/cache_reg[1][89]  ( .D(\D_cache/n1083 ), .CK(clk), .RN(n5767), .Q(\D_cache/cache[1][89] ), .QN(n2948) );
  DFFRX1 \D_cache/cache_reg[2][89]  ( .D(\D_cache/n1082 ), .CK(clk), .RN(n5767), .Q(\D_cache/cache[2][89] ), .QN(n1334) );
  DFFRX1 \D_cache/cache_reg[3][89]  ( .D(\D_cache/n1081 ), .CK(clk), .RN(n5767), .Q(\D_cache/cache[3][89] ), .QN(n2946) );
  DFFRX1 \D_cache/cache_reg[4][89]  ( .D(\D_cache/n1080 ), .CK(clk), .RN(n5767), .Q(\D_cache/cache[4][89] ), .QN(n1335) );
  DFFRX1 \D_cache/cache_reg[5][89]  ( .D(\D_cache/n1079 ), .CK(clk), .RN(n5767), .Q(\D_cache/cache[5][89] ), .QN(n2947) );
  DFFRX1 \D_cache/cache_reg[6][89]  ( .D(\D_cache/n1078 ), .CK(clk), .RN(n5767), .Q(\D_cache/cache[6][89] ), .QN(n1528) );
  DFFRX1 \D_cache/cache_reg[7][89]  ( .D(\D_cache/n1077 ), .CK(clk), .RN(n5768), .Q(\D_cache/cache[7][89] ), .QN(n3141) );
  DFFRX1 \D_cache/cache_reg[0][90]  ( .D(\D_cache/n1076 ), .CK(clk), .RN(n5768), .Q(\D_cache/cache[0][90] ), .QN(n1463) );
  DFFRX1 \D_cache/cache_reg[1][90]  ( .D(\D_cache/n1075 ), .CK(clk), .RN(n5768), .Q(\D_cache/cache[1][90] ), .QN(n3076) );
  DFFRX1 \D_cache/cache_reg[2][90]  ( .D(\D_cache/n1074 ), .CK(clk), .RN(n5768), .Q(\D_cache/cache[2][90] ), .QN(n1299) );
  DFFRX1 \D_cache/cache_reg[3][90]  ( .D(\D_cache/n1073 ), .CK(clk), .RN(n5768), .Q(\D_cache/cache[3][90] ), .QN(n2911) );
  DFFRX1 \D_cache/cache_reg[4][90]  ( .D(\D_cache/n1072 ), .CK(clk), .RN(n5768), .Q(\D_cache/cache[4][90] ), .QN(n1300) );
  DFFRX1 \D_cache/cache_reg[5][90]  ( .D(\D_cache/n1071 ), .CK(clk), .RN(n5768), .Q(\D_cache/cache[5][90] ), .QN(n2912) );
  DFFRX1 \D_cache/cache_reg[6][90]  ( .D(\D_cache/n1070 ), .CK(clk), .RN(n5768), .Q(\D_cache/cache[6][90] ), .QN(n1522) );
  DFFRX1 \D_cache/cache_reg[7][90]  ( .D(\D_cache/n1069 ), .CK(clk), .RN(n5768), .Q(\D_cache/cache[7][90] ), .QN(n3135) );
  DFFRX1 \D_cache/cache_reg[0][91]  ( .D(\D_cache/n1068 ), .CK(clk), .RN(n5768), .Q(\D_cache/cache[0][91] ), .QN(n1302) );
  DFFRX1 \D_cache/cache_reg[1][91]  ( .D(\D_cache/n1067 ), .CK(clk), .RN(n5768), .Q(\D_cache/cache[1][91] ), .QN(n2914) );
  DFFRX1 \D_cache/cache_reg[2][91]  ( .D(\D_cache/n1066 ), .CK(clk), .RN(n5768), .Q(\D_cache/cache[2][91] ), .QN(n1301) );
  DFFRX1 \D_cache/cache_reg[3][91]  ( .D(\D_cache/n1065 ), .CK(clk), .RN(n5769), .Q(\D_cache/cache[3][91] ), .QN(n2913) );
  DFFRX1 \D_cache/cache_reg[4][91]  ( .D(\D_cache/n1064 ), .CK(clk), .RN(n5769), .Q(\D_cache/cache[4][91] ), .QN(n1468) );
  DFFRX1 \D_cache/cache_reg[5][91]  ( .D(\D_cache/n1063 ), .CK(clk), .RN(n5769), .Q(\D_cache/cache[5][91] ), .QN(n3081) );
  DFFRX1 \D_cache/cache_reg[6][91]  ( .D(\D_cache/n1062 ), .CK(clk), .RN(n5769), .Q(\D_cache/cache[6][91] ), .QN(n1447) );
  DFFRX1 \D_cache/cache_reg[7][91]  ( .D(\D_cache/n1061 ), .CK(clk), .RN(n5769), .Q(\D_cache/cache[7][91] ), .QN(n3060) );
  DFFRX1 \D_cache/cache_reg[0][92]  ( .D(\D_cache/n1060 ), .CK(clk), .RN(n5769), .Q(\D_cache/cache[0][92] ), .QN(n1252) );
  DFFRX1 \D_cache/cache_reg[1][92]  ( .D(\D_cache/n1059 ), .CK(clk), .RN(n5769), .Q(\D_cache/cache[1][92] ), .QN(n2863) );
  DFFRX1 \D_cache/cache_reg[2][92]  ( .D(\D_cache/n1058 ), .CK(clk), .RN(n5769), .Q(\D_cache/cache[2][92] ), .QN(n1253) );
  DFFRX1 \D_cache/cache_reg[3][92]  ( .D(\D_cache/n1057 ), .CK(clk), .RN(n5769), .Q(\D_cache/cache[3][92] ), .QN(n2864) );
  DFFRX1 \D_cache/cache_reg[4][92]  ( .D(\D_cache/n1056 ), .CK(clk), .RN(n5769), .Q(\D_cache/cache[4][92] ), .QN(n2812) );
  DFFRX1 \D_cache/cache_reg[5][92]  ( .D(\D_cache/n1055 ), .CK(clk), .RN(n5769), .Q(\D_cache/cache[5][92] ), .QN(n820) );
  DFFRX1 \D_cache/cache_reg[6][92]  ( .D(\D_cache/n1054 ), .CK(clk), .RN(n5769), .Q(\D_cache/cache[6][92] ), .QN(n1482) );
  DFFRX1 \D_cache/cache_reg[7][92]  ( .D(\D_cache/n1053 ), .CK(clk), .RN(n5770), .Q(\D_cache/cache[7][92] ), .QN(n3095) );
  DFFRX1 \D_cache/cache_reg[0][93]  ( .D(\D_cache/n1052 ), .CK(clk), .RN(n5770), .Q(\D_cache/cache[0][93] ), .QN(n1312) );
  DFFRX1 \D_cache/cache_reg[1][93]  ( .D(\D_cache/n1051 ), .CK(clk), .RN(n5770), .Q(\D_cache/cache[1][93] ), .QN(n2924) );
  DFFRX1 \D_cache/cache_reg[2][93]  ( .D(\D_cache/n1050 ), .CK(clk), .RN(n5770), .Q(\D_cache/cache[2][93] ), .QN(n1311) );
  DFFRX1 \D_cache/cache_reg[3][93]  ( .D(\D_cache/n1049 ), .CK(clk), .RN(n5770), .Q(\D_cache/cache[3][93] ), .QN(n2923) );
  DFFRX1 \D_cache/cache_reg[4][93]  ( .D(\D_cache/n1048 ), .CK(clk), .RN(n5770), .Q(\D_cache/cache[4][93] ), .QN(n1313) );
  DFFRX1 \D_cache/cache_reg[5][93]  ( .D(\D_cache/n1047 ), .CK(clk), .RN(n5770), .Q(\D_cache/cache[5][93] ), .QN(n2925) );
  DFFRX1 \D_cache/cache_reg[6][93]  ( .D(\D_cache/n1046 ), .CK(clk), .RN(n5770), .Q(\D_cache/cache[6][93] ), .QN(n1553) );
  DFFRX1 \D_cache/cache_reg[7][93]  ( .D(\D_cache/n1045 ), .CK(clk), .RN(n5770), .Q(\D_cache/cache[7][93] ), .QN(n3166) );
  DFFRX1 \D_cache/cache_reg[0][94]  ( .D(\D_cache/n1044 ), .CK(clk), .RN(n5770), .Q(\D_cache/cache[0][94] ), .QN(n1958) );
  DFFRX1 \D_cache/cache_reg[1][94]  ( .D(\D_cache/n1043 ), .CK(clk), .RN(n5770), .Q(\D_cache/cache[1][94] ), .QN(n386) );
  DFFRX1 \D_cache/cache_reg[2][94]  ( .D(\D_cache/n1042 ), .CK(clk), .RN(n5770), .Q(\D_cache/cache[2][94] ), .QN(n454) );
  DFFRX1 \D_cache/cache_reg[3][94]  ( .D(\D_cache/n1041 ), .CK(clk), .RN(n5771), .Q(\D_cache/cache[3][94] ), .QN(n2010) );
  DFFRX1 \D_cache/cache_reg[4][94]  ( .D(\D_cache/n1040 ), .CK(clk), .RN(n5771), .Q(\D_cache/cache[4][94] ), .QN(n807) );
  DFFRX1 \D_cache/cache_reg[5][94]  ( .D(\D_cache/n1039 ), .CK(clk), .RN(n5771), .Q(\D_cache/cache[5][94] ), .QN(n2340) );
  DFFRX1 \D_cache/cache_reg[6][94]  ( .D(\D_cache/n1038 ), .CK(clk), .RN(n5771), .Q(\D_cache/cache[6][94] ), .QN(n1948) );
  DFFRX1 \D_cache/cache_reg[7][94]  ( .D(\D_cache/n1037 ), .CK(clk), .RN(n5771), .Q(\D_cache/cache[7][94] ), .QN(n370) );
  DFFRX1 \D_cache/cache_reg[0][95]  ( .D(\D_cache/n1036 ), .CK(clk), .RN(n5771), .Q(\D_cache/cache[0][95] ), .QN(n1264) );
  DFFRX1 \D_cache/cache_reg[1][95]  ( .D(\D_cache/n1035 ), .CK(clk), .RN(n5771), .Q(\D_cache/cache[1][95] ), .QN(n2875) );
  DFFRX1 \D_cache/cache_reg[2][95]  ( .D(\D_cache/n1034 ), .CK(clk), .RN(n5771), .Q(\D_cache/cache[2][95] ), .QN(n1265) );
  DFFRX1 \D_cache/cache_reg[3][95]  ( .D(\D_cache/n1033 ), .CK(clk), .RN(n5771), .Q(\D_cache/cache[3][95] ), .QN(n2876) );
  DFFRX1 \D_cache/cache_reg[4][95]  ( .D(\D_cache/n1032 ), .CK(clk), .RN(n5771), .Q(\D_cache/cache[4][95] ), .QN(n1266) );
  DFFRX1 \D_cache/cache_reg[5][95]  ( .D(\D_cache/n1031 ), .CK(clk), .RN(n5771), .Q(\D_cache/cache[5][95] ), .QN(n2877) );
  DFFRX1 \D_cache/cache_reg[6][95]  ( .D(\D_cache/n1030 ), .CK(clk), .RN(n5771), .Q(\D_cache/cache[6][95] ), .QN(n1558) );
  DFFRX1 \D_cache/cache_reg[7][95]  ( .D(\D_cache/n1029 ), .CK(clk), .RN(n5772), .Q(\D_cache/cache[7][95] ), .QN(n3171) );
  DFFRX1 \D_cache/cache_reg[0][96]  ( .D(\D_cache/n1028 ), .CK(clk), .RN(n5772), .Q(\D_cache/cache[0][96] ), .QN(n1392) );
  DFFRX1 \D_cache/cache_reg[1][96]  ( .D(\D_cache/n1027 ), .CK(clk), .RN(n5772), .Q(\D_cache/cache[1][96] ), .QN(n3005) );
  DFFRX1 \D_cache/cache_reg[2][96]  ( .D(\D_cache/n1026 ), .CK(clk), .RN(n5772), .Q(\D_cache/cache[2][96] ), .QN(n1393) );
  DFFRX1 \D_cache/cache_reg[3][96]  ( .D(\D_cache/n1025 ), .CK(clk), .RN(n5772), .Q(\D_cache/cache[3][96] ), .QN(n3006) );
  DFFRX1 \D_cache/cache_reg[4][96]  ( .D(\D_cache/n1024 ), .CK(clk), .RN(n5772), .Q(\D_cache/cache[4][96] ), .QN(n2369) );
  DFFRX1 \D_cache/cache_reg[5][96]  ( .D(\D_cache/n1023 ), .CK(clk), .RN(n5772), .Q(\D_cache/cache[5][96] ), .QN(n373) );
  DFFRX1 \D_cache/cache_reg[6][96]  ( .D(\D_cache/n1022 ), .CK(clk), .RN(n5772), .Q(\D_cache/cache[6][96] ), .QN(n1248) );
  DFFRX1 \D_cache/cache_reg[7][96]  ( .D(\D_cache/n1021 ), .CK(clk), .RN(n5772), .Q(\D_cache/cache[7][96] ), .QN(n2856) );
  DFFRX1 \D_cache/cache_reg[0][97]  ( .D(\D_cache/n1020 ), .CK(clk), .RN(n5772), .Q(\D_cache/cache[0][97] ), .QN(n925) );
  DFFRX1 \D_cache/cache_reg[1][97]  ( .D(\D_cache/n1019 ), .CK(clk), .RN(n5772), .Q(\D_cache/cache[1][97] ), .QN(n2448) );
  DFFRX1 \D_cache/cache_reg[2][97]  ( .D(\D_cache/n1018 ), .CK(clk), .RN(n5772), .Q(\D_cache/cache[2][97] ), .QN(n1381) );
  DFFRX1 \D_cache/cache_reg[3][97]  ( .D(\D_cache/n1017 ), .CK(clk), .RN(n5773), .Q(\D_cache/cache[3][97] ), .QN(n2994) );
  DFFRX1 \D_cache/cache_reg[4][97]  ( .D(\D_cache/n1016 ), .CK(clk), .RN(n5773), .Q(\D_cache/cache[4][97] ), .QN(n1574) );
  DFFRX1 \D_cache/cache_reg[5][97]  ( .D(\D_cache/n1015 ), .CK(clk), .RN(n5773), .Q(\D_cache/cache[5][97] ), .QN(n3187) );
  DFFRX1 \D_cache/cache_reg[6][97]  ( .D(\D_cache/n1014 ), .CK(clk), .RN(n5773), .Q(\D_cache/cache[6][97] ), .QN(n926) );
  DFFRX1 \D_cache/cache_reg[7][97]  ( .D(\D_cache/n1013 ), .CK(clk), .RN(n5773), .Q(\D_cache/cache[7][97] ), .QN(n2449) );
  DFFRX1 \D_cache/cache_reg[0][98]  ( .D(\D_cache/n1012 ), .CK(clk), .RN(n5773), .Q(\D_cache/cache[0][98] ), .QN(n1359) );
  DFFRX1 \D_cache/cache_reg[1][98]  ( .D(\D_cache/n1011 ), .CK(clk), .RN(n5773), .Q(\D_cache/cache[1][98] ), .QN(n2972) );
  DFFRX1 \D_cache/cache_reg[2][98]  ( .D(\D_cache/n1010 ), .CK(clk), .RN(n5773), .Q(\D_cache/cache[2][98] ), .QN(n1360) );
  DFFRX1 \D_cache/cache_reg[3][98]  ( .D(\D_cache/n1009 ), .CK(clk), .RN(n5773), .Q(\D_cache/cache[3][98] ), .QN(n2973) );
  DFFRX1 \D_cache/cache_reg[4][98]  ( .D(\D_cache/n1008 ), .CK(clk), .RN(n5773), .Q(\D_cache/cache[4][98] ), .QN(n2815) );
  DFFRX1 \D_cache/cache_reg[5][98]  ( .D(\D_cache/n1007 ), .CK(clk), .RN(n5773), .Q(\D_cache/cache[5][98] ), .QN(n823) );
  DFFRX1 \D_cache/cache_reg[6][98]  ( .D(\D_cache/n1006 ), .CK(clk), .RN(n5773), .Q(\D_cache/cache[6][98] ), .QN(n1442) );
  DFFRX1 \D_cache/cache_reg[7][98]  ( .D(\D_cache/n1005 ), .CK(clk), .RN(n5774), .Q(\D_cache/cache[7][98] ), .QN(n3055) );
  DFFRX1 \D_cache/cache_reg[0][99]  ( .D(\D_cache/n1004 ), .CK(clk), .RN(n5774), .Q(\D_cache/cache[0][99] ), .QN(n2823) );
  DFFRX1 \D_cache/cache_reg[1][99]  ( .D(\D_cache/n1003 ), .CK(clk), .RN(n5774), .Q(\D_cache/cache[1][99] ), .QN(n831) );
  DFFRX1 \D_cache/cache_reg[2][99]  ( .D(\D_cache/n1002 ), .CK(clk), .RN(n5774), .Q(\D_cache/cache[2][99] ), .QN(n2441) );
  DFFRX1 \D_cache/cache_reg[3][99]  ( .D(\D_cache/n1001 ), .CK(clk), .RN(n5774), .Q(\D_cache/cache[3][99] ), .QN(n466) );
  DFFRX1 \D_cache/cache_reg[4][99]  ( .D(\D_cache/n1000 ), .CK(clk), .RN(n5774), .Q(\D_cache/cache[4][99] ), .QN(n2442) );
  DFFRX1 \D_cache/cache_reg[5][99]  ( .D(\D_cache/n999 ), .CK(clk), .RN(n5774), 
        .Q(\D_cache/cache[5][99] ), .QN(n467) );
  DFFRX1 \D_cache/cache_reg[6][99]  ( .D(\D_cache/n998 ), .CK(clk), .RN(n5774), 
        .Q(\D_cache/cache[6][99] ), .QN(n2807) );
  DFFRX1 \D_cache/cache_reg[7][99]  ( .D(\D_cache/n997 ), .CK(clk), .RN(n5774), 
        .Q(\D_cache/cache[7][99] ), .QN(n805) );
  DFFRX1 \D_cache/cache_reg[0][100]  ( .D(\D_cache/n996 ), .CK(clk), .RN(n5774), .Q(\D_cache/cache[0][100] ), .QN(n1378) );
  DFFRX1 \D_cache/cache_reg[1][100]  ( .D(\D_cache/n995 ), .CK(clk), .RN(n5774), .Q(\D_cache/cache[1][100] ), .QN(n2991) );
  DFFRX1 \D_cache/cache_reg[2][100]  ( .D(\D_cache/n994 ), .CK(clk), .RN(n5774), .Q(\D_cache/cache[2][100] ), .QN(n1379) );
  DFFRX1 \D_cache/cache_reg[3][100]  ( .D(\D_cache/n993 ), .CK(clk), .RN(n5775), .Q(\D_cache/cache[3][100] ), .QN(n2992) );
  DFFRX1 \D_cache/cache_reg[4][100]  ( .D(\D_cache/n992 ), .CK(clk), .RN(n5775), .Q(\D_cache/cache[4][100] ), .QN(n2381) );
  DFFRX1 \D_cache/cache_reg[5][100]  ( .D(\D_cache/n991 ), .CK(clk), .RN(n5775), .Q(\D_cache/cache[5][100] ), .QN(n374) );
  DFFRX1 \D_cache/cache_reg[6][100]  ( .D(\D_cache/n990 ), .CK(clk), .RN(n5775), .Q(\D_cache/cache[6][100] ), .QN(n1494) );
  DFFRX1 \D_cache/cache_reg[7][100]  ( .D(\D_cache/n989 ), .CK(clk), .RN(n5775), .Q(\D_cache/cache[7][100] ), .QN(n3107) );
  DFFRX1 \D_cache/cache_reg[0][101]  ( .D(\D_cache/n988 ), .CK(clk), .RN(n5775), .Q(\D_cache/cache[0][101] ), .QN(n1368) );
  DFFRX1 \D_cache/cache_reg[1][101]  ( .D(\D_cache/n987 ), .CK(clk), .RN(n5775), .Q(\D_cache/cache[1][101] ), .QN(n2981) );
  DFFRX1 \D_cache/cache_reg[2][101]  ( .D(\D_cache/n986 ), .CK(clk), .RN(n5775), .Q(\D_cache/cache[2][101] ), .QN(n932) );
  DFFRX1 \D_cache/cache_reg[3][101]  ( .D(\D_cache/n985 ), .CK(clk), .RN(n5775), .Q(\D_cache/cache[3][101] ), .QN(n2456) );
  DFFRX1 \D_cache/cache_reg[4][101]  ( .D(\D_cache/n984 ), .CK(clk), .RN(n5775), .Q(\D_cache/cache[4][101] ), .QN(n2379) );
  DFFRX1 \D_cache/cache_reg[5][101]  ( .D(\D_cache/n983 ), .CK(clk), .RN(n5775), .Q(\D_cache/cache[5][101] ), .QN(n875) );
  DFFRX1 \D_cache/cache_reg[6][101]  ( .D(\D_cache/n982 ), .CK(clk), .RN(n5775), .Q(\D_cache/cache[6][101] ), .QN(n1545) );
  DFFRX1 \D_cache/cache_reg[7][101]  ( .D(\D_cache/n981 ), .CK(clk), .RN(n5776), .Q(\D_cache/cache[7][101] ), .QN(n3158) );
  DFFRX1 \D_cache/cache_reg[0][102]  ( .D(\D_cache/n980 ), .CK(clk), .RN(n5776), .Q(\D_cache/cache[0][102] ), .QN(n1459) );
  DFFRX1 \D_cache/cache_reg[1][102]  ( .D(\D_cache/n979 ), .CK(clk), .RN(n5776), .Q(\D_cache/cache[1][102] ), .QN(n3072) );
  DFFRX1 \D_cache/cache_reg[2][102]  ( .D(\D_cache/n978 ), .CK(clk), .RN(n5776), .Q(\D_cache/cache[2][102] ), .QN(n1242) );
  DFFRX1 \D_cache/cache_reg[3][102]  ( .D(\D_cache/n977 ), .CK(clk), .RN(n5776), .Q(\D_cache/cache[3][102] ), .QN(n2847) );
  DFFRX1 \D_cache/cache_reg[4][102]  ( .D(\D_cache/n976 ), .CK(clk), .RN(n5776), .Q(\D_cache/cache[4][102] ), .QN(n1243) );
  DFFRX1 \D_cache/cache_reg[5][102]  ( .D(\D_cache/n975 ), .CK(clk), .RN(n5776), .Q(\D_cache/cache[5][102] ), .QN(n2848) );
  DFFRX1 \D_cache/cache_reg[6][102]  ( .D(\D_cache/n974 ), .CK(clk), .RN(n5776), .Q(\D_cache/cache[6][102] ), .QN(n1244) );
  DFFRX1 \D_cache/cache_reg[7][102]  ( .D(\D_cache/n973 ), .CK(clk), .RN(n5776), .Q(\D_cache/cache[7][102] ), .QN(n2849) );
  DFFRX1 \D_cache/cache_reg[0][103]  ( .D(\D_cache/n972 ), .CK(clk), .RN(n5776), .Q(\D_cache/cache[0][103] ), .QN(n1536) );
  DFFRX1 \D_cache/cache_reg[1][103]  ( .D(\D_cache/n971 ), .CK(clk), .RN(n5776), .Q(\D_cache/cache[1][103] ), .QN(n3149) );
  DFFRX1 \D_cache/cache_reg[2][103]  ( .D(\D_cache/n970 ), .CK(clk), .RN(n5776), .Q(\D_cache/cache[2][103] ), .QN(n1398) );
  DFFRX1 \D_cache/cache_reg[3][103]  ( .D(\D_cache/n969 ), .CK(clk), .RN(n5777), .Q(\D_cache/cache[3][103] ), .QN(n3011) );
  DFFRX1 \D_cache/cache_reg[4][103]  ( .D(\D_cache/n968 ), .CK(clk), .RN(n5777), .Q(\D_cache/cache[4][103] ), .QN(n2383) );
  DFFRX1 \D_cache/cache_reg[5][103]  ( .D(\D_cache/n967 ), .CK(clk), .RN(n5777), .Q(\D_cache/cache[5][103] ), .QN(n878) );
  DFFRX1 \D_cache/cache_reg[6][103]  ( .D(\D_cache/n966 ), .CK(clk), .RN(n5777), .Q(\D_cache/cache[6][103] ), .QN(n1399) );
  DFFRX1 \D_cache/cache_reg[7][103]  ( .D(\D_cache/n965 ), .CK(clk), .RN(n5777), .Q(\D_cache/cache[7][103] ), .QN(n3012) );
  DFFRX1 \D_cache/cache_reg[0][104]  ( .D(\D_cache/n964 ), .CK(clk), .RN(n5777), .Q(\D_cache/cache[0][104] ), .QN(n1534) );
  DFFRX1 \D_cache/cache_reg[1][104]  ( .D(\D_cache/n963 ), .CK(clk), .RN(n5777), .Q(\D_cache/cache[1][104] ), .QN(n3147) );
  DFFRX1 \D_cache/cache_reg[2][104]  ( .D(\D_cache/n962 ), .CK(clk), .RN(n5777), .Q(\D_cache/cache[2][104] ), .QN(n1412) );
  DFFRX1 \D_cache/cache_reg[3][104]  ( .D(\D_cache/n961 ), .CK(clk), .RN(n5777), .Q(\D_cache/cache[3][104] ), .QN(n3025) );
  DFFRX1 \D_cache/cache_reg[4][104]  ( .D(\D_cache/n960 ), .CK(clk), .RN(n5777), .Q(\D_cache/cache[4][104] ), .QN(n1413) );
  DFFRX1 \D_cache/cache_reg[5][104]  ( .D(\D_cache/n959 ), .CK(clk), .RN(n5777), .Q(\D_cache/cache[5][104] ), .QN(n3026) );
  DFFRX1 \D_cache/cache_reg[6][104]  ( .D(\D_cache/n958 ), .CK(clk), .RN(n5777), .Q(\D_cache/cache[6][104] ), .QN(n1414) );
  DFFRX1 \D_cache/cache_reg[7][104]  ( .D(\D_cache/n957 ), .CK(clk), .RN(n5778), .Q(\D_cache/cache[7][104] ), .QN(n3027) );
  DFFRX1 \D_cache/cache_reg[0][105]  ( .D(\D_cache/n956 ), .CK(clk), .RN(n5778), .Q(\D_cache/cache[0][105] ), .QN(n1245) );
  DFFRX1 \D_cache/cache_reg[1][105]  ( .D(\D_cache/n955 ), .CK(clk), .RN(n5778), .Q(\D_cache/cache[1][105] ), .QN(n2850) );
  DFFRX1 \D_cache/cache_reg[2][105]  ( .D(\D_cache/n954 ), .CK(clk), .RN(n5778), .Q(\D_cache/cache[2][105] ), .QN(n1409) );
  DFFRX1 \D_cache/cache_reg[3][105]  ( .D(\D_cache/n953 ), .CK(clk), .RN(n5778), .Q(\D_cache/cache[3][105] ), .QN(n3022) );
  DFFRX1 \D_cache/cache_reg[4][105]  ( .D(\D_cache/n952 ), .CK(clk), .RN(n5778), .Q(\D_cache/cache[4][105] ), .QN(n938) );
  DFFRX1 \D_cache/cache_reg[5][105]  ( .D(\D_cache/n951 ), .CK(clk), .RN(n5778), .Q(\D_cache/cache[5][105] ), .QN(n2463) );
  DFFRX1 \D_cache/cache_reg[6][105]  ( .D(\D_cache/n950 ), .CK(clk), .RN(n5778), .Q(\D_cache/cache[6][105] ), .QN(n1410) );
  DFFRX1 \D_cache/cache_reg[7][105]  ( .D(\D_cache/n949 ), .CK(clk), .RN(n5778), .Q(\D_cache/cache[7][105] ), .QN(n3023) );
  DFFRX1 \D_cache/cache_reg[0][106]  ( .D(\D_cache/n948 ), .CK(clk), .RN(n5778), .Q(\D_cache/cache[0][106] ), .QN(n1369) );
  DFFRX1 \D_cache/cache_reg[1][106]  ( .D(\D_cache/n947 ), .CK(clk), .RN(n5778), .Q(\D_cache/cache[1][106] ), .QN(n2982) );
  DFFRX1 \D_cache/cache_reg[2][106]  ( .D(\D_cache/n946 ), .CK(clk), .RN(n5778), .Q(\D_cache/cache[2][106] ), .QN(n1370) );
  DFFRX1 \D_cache/cache_reg[3][106]  ( .D(\D_cache/n945 ), .CK(clk), .RN(n5779), .Q(\D_cache/cache[3][106] ), .QN(n2983) );
  DFFRX1 \D_cache/cache_reg[4][106]  ( .D(\D_cache/n944 ), .CK(clk), .RN(n5779), .Q(\D_cache/cache[4][106] ), .QN(n1371) );
  DFFRX1 \D_cache/cache_reg[5][106]  ( .D(\D_cache/n943 ), .CK(clk), .RN(n5779), .Q(\D_cache/cache[5][106] ), .QN(n2984) );
  DFFRX1 \D_cache/cache_reg[6][106]  ( .D(\D_cache/n942 ), .CK(clk), .RN(n5779), .Q(\D_cache/cache[6][106] ), .QN(n1542) );
  DFFRX1 \D_cache/cache_reg[7][106]  ( .D(\D_cache/n941 ), .CK(clk), .RN(n5779), .Q(\D_cache/cache[7][106] ), .QN(n3155) );
  DFFRX1 \D_cache/cache_reg[0][107]  ( .D(\D_cache/n940 ), .CK(clk), .RN(n5779), .Q(\D_cache/cache[0][107] ), .QN(n934) );
  DFFRX1 \D_cache/cache_reg[1][107]  ( .D(\D_cache/n939 ), .CK(clk), .RN(n5779), .Q(\D_cache/cache[1][107] ), .QN(n2459) );
  DFFRX1 \D_cache/cache_reg[2][107]  ( .D(\D_cache/n938 ), .CK(clk), .RN(n5779), .Q(\D_cache/cache[2][107] ), .QN(n1374) );
  DFFRX1 \D_cache/cache_reg[3][107]  ( .D(\D_cache/n937 ), .CK(clk), .RN(n5779), .Q(\D_cache/cache[3][107] ), .QN(n2987) );
  DFFRX1 \D_cache/cache_reg[4][107]  ( .D(\D_cache/n936 ), .CK(clk), .RN(n5779), .Q(\D_cache/cache[4][107] ), .QN(n2419) );
  DFFRX1 \D_cache/cache_reg[5][107]  ( .D(\D_cache/n935 ), .CK(clk), .RN(n5779), .Q(\D_cache/cache[5][107] ), .QN(n465) );
  DFFRX1 \D_cache/cache_reg[6][107]  ( .D(\D_cache/n934 ), .CK(clk), .RN(n5779), .Q(\D_cache/cache[6][107] ), .QN(n2445) );
  DFFRX1 \D_cache/cache_reg[7][107]  ( .D(\D_cache/n933 ), .CK(clk), .RN(n5780), .Q(\D_cache/cache[7][107] ), .QN(n470) );
  DFFRX1 \D_cache/cache_reg[0][108]  ( .D(\D_cache/n932 ), .CK(clk), .RN(n5780), .Q(\D_cache/cache[0][108] ), .QN(n923) );
  DFFRX1 \D_cache/cache_reg[1][108]  ( .D(\D_cache/n931 ), .CK(clk), .RN(n5780), .Q(\D_cache/cache[1][108] ), .QN(n2450) );
  DFFRX1 \D_cache/cache_reg[2][108]  ( .D(\D_cache/n930 ), .CK(clk), .RN(n5780), .Q(\D_cache/cache[2][108] ), .QN(n1411) );
  DFFRX1 \D_cache/cache_reg[3][108]  ( .D(\D_cache/n929 ), .CK(clk), .RN(n5780), .Q(\D_cache/cache[3][108] ), .QN(n3024) );
  DFFRX1 \D_cache/cache_reg[4][108]  ( .D(\D_cache/n928 ), .CK(clk), .RN(n5780), .Q(\D_cache/cache[4][108] ), .QN(n2360) );
  DFFRX1 \D_cache/cache_reg[5][108]  ( .D(\D_cache/n927 ), .CK(clk), .RN(n5780), .Q(\D_cache/cache[5][108] ), .QN(n857) );
  DFFRX1 \D_cache/cache_reg[6][108]  ( .D(\D_cache/n926 ), .CK(clk), .RN(n5780), .Q(\D_cache/cache[6][108] ), .QN(n1234) );
  DFFRX1 \D_cache/cache_reg[7][108]  ( .D(\D_cache/n925 ), .CK(clk), .RN(n5780), .Q(\D_cache/cache[7][108] ), .QN(n2839) );
  DFFRX1 \D_cache/cache_reg[0][109]  ( .D(\D_cache/n924 ), .CK(clk), .RN(n5780), .Q(\D_cache/cache[0][109] ), .QN(n1408) );
  DFFRX1 \D_cache/cache_reg[1][109]  ( .D(\D_cache/n923 ), .CK(clk), .RN(n5780), .Q(\D_cache/cache[1][109] ), .QN(n3021) );
  DFFRX1 \D_cache/cache_reg[2][109]  ( .D(\D_cache/n922 ), .CK(clk), .RN(n5780), .Q(\D_cache/cache[2][109] ), .QN(n1407) );
  DFFRX1 \D_cache/cache_reg[3][109]  ( .D(\D_cache/n921 ), .CK(clk), .RN(n5781), .Q(\D_cache/cache[3][109] ), .QN(n3020) );
  DFFRX1 \D_cache/cache_reg[4][109]  ( .D(\D_cache/n920 ), .CK(clk), .RN(n5781), .Q(\D_cache/cache[4][109] ), .QN(n2361) );
  DFFRX1 \D_cache/cache_reg[5][109]  ( .D(\D_cache/n919 ), .CK(clk), .RN(n5781), .Q(\D_cache/cache[5][109] ), .QN(n858) );
  DFFRX1 \D_cache/cache_reg[6][109]  ( .D(\D_cache/n918 ), .CK(clk), .RN(n5781), .Q(\D_cache/cache[6][109] ), .QN(n1485) );
  DFFRX1 \D_cache/cache_reg[7][109]  ( .D(\D_cache/n917 ), .CK(clk), .RN(n5781), .Q(\D_cache/cache[7][109] ), .QN(n3098) );
  DFFRX1 \D_cache/cache_reg[0][110]  ( .D(\D_cache/n916 ), .CK(clk), .RN(n5781), .Q(\D_cache/cache[0][110] ), .QN(n1479) );
  DFFRX1 \D_cache/cache_reg[1][110]  ( .D(\D_cache/n915 ), .CK(clk), .RN(n5781), .Q(\D_cache/cache[1][110] ), .QN(n3092) );
  DFFRX1 \D_cache/cache_reg[2][110]  ( .D(\D_cache/n914 ), .CK(clk), .RN(n5781), .Q(\D_cache/cache[2][110] ), .QN(n1404) );
  DFFRX1 \D_cache/cache_reg[3][110]  ( .D(\D_cache/n913 ), .CK(clk), .RN(n5781), .Q(\D_cache/cache[3][110] ), .QN(n3017) );
  DFFRX1 \D_cache/cache_reg[4][110]  ( .D(\D_cache/n912 ), .CK(clk), .RN(n5781), .Q(\D_cache/cache[4][110] ), .QN(n1405) );
  DFFRX1 \D_cache/cache_reg[5][110]  ( .D(\D_cache/n911 ), .CK(clk), .RN(n5781), .Q(\D_cache/cache[5][110] ), .QN(n3018) );
  DFFRX1 \D_cache/cache_reg[6][110]  ( .D(\D_cache/n910 ), .CK(clk), .RN(n5781), .Q(\D_cache/cache[6][110] ), .QN(n1406) );
  DFFRX1 \D_cache/cache_reg[7][110]  ( .D(\D_cache/n909 ), .CK(clk), .RN(n5782), .Q(\D_cache/cache[7][110] ), .QN(n3019) );
  DFFRX1 \D_cache/cache_reg[0][111]  ( .D(\D_cache/n908 ), .CK(clk), .RN(n5782), .Q(\D_cache/cache[0][111] ), .QN(n2371) );
  DFFRX1 \D_cache/cache_reg[1][111]  ( .D(\D_cache/n907 ), .CK(clk), .RN(n5782), .Q(\D_cache/cache[1][111] ), .QN(n867) );
  DFFRX1 \D_cache/cache_reg[2][111]  ( .D(\D_cache/n906 ), .CK(clk), .RN(n5782), .Q(\D_cache/cache[2][111] ), .QN(n1415) );
  DFFRX1 \D_cache/cache_reg[3][111]  ( .D(\D_cache/n905 ), .CK(clk), .RN(n5782), .Q(\D_cache/cache[3][111] ), .QN(n3028) );
  DFFRX1 \D_cache/cache_reg[4][111]  ( .D(\D_cache/n904 ), .CK(clk), .RN(n5782), .Q(\D_cache/cache[4][111] ), .QN(n2395) );
  DFFRX1 \D_cache/cache_reg[5][111]  ( .D(\D_cache/n903 ), .CK(clk), .RN(n5782), .Q(\D_cache/cache[5][111] ), .QN(n890) );
  DFFRX1 \D_cache/cache_reg[6][111]  ( .D(\D_cache/n902 ), .CK(clk), .RN(n5782), .Q(\D_cache/cache[6][111] ), .QN(n1416) );
  DFFRX1 \D_cache/cache_reg[7][111]  ( .D(\D_cache/n901 ), .CK(clk), .RN(n5782), .Q(\D_cache/cache[7][111] ), .QN(n3029) );
  DFFRX1 \D_cache/cache_reg[0][112]  ( .D(\D_cache/n900 ), .CK(clk), .RN(n5782), .Q(\D_cache/cache[0][112] ), .QN(n1376) );
  DFFRX1 \D_cache/cache_reg[1][112]  ( .D(\D_cache/n899 ), .CK(clk), .RN(n5782), .Q(\D_cache/cache[1][112] ), .QN(n2989) );
  DFFRX1 \D_cache/cache_reg[2][112]  ( .D(\D_cache/n898 ), .CK(clk), .RN(n5782), .Q(\D_cache/cache[2][112] ), .QN(n1375) );
  DFFRX1 \D_cache/cache_reg[3][112]  ( .D(\D_cache/n897 ), .CK(clk), .RN(n5783), .Q(\D_cache/cache[3][112] ), .QN(n2988) );
  DFFRX1 \D_cache/cache_reg[4][112]  ( .D(\D_cache/n896 ), .CK(clk), .RN(n5783), .Q(\D_cache/cache[4][112] ), .QN(n1377) );
  DFFRX1 \D_cache/cache_reg[5][112]  ( .D(\D_cache/n895 ), .CK(clk), .RN(n5783), .Q(\D_cache/cache[5][112] ), .QN(n2990) );
  DFFRX1 \D_cache/cache_reg[6][112]  ( .D(\D_cache/n894 ), .CK(clk), .RN(n5783), .Q(\D_cache/cache[6][112] ), .QN(n1444) );
  DFFRX1 \D_cache/cache_reg[7][112]  ( .D(\D_cache/n893 ), .CK(clk), .RN(n5783), .Q(\D_cache/cache[7][112] ), .QN(n3057) );
  DFFRX1 \D_cache/cache_reg[0][113]  ( .D(\D_cache/n892 ), .CK(clk), .RN(n5783), .Q(\D_cache/cache[0][113] ), .QN(n2809) );
  DFFRX1 \D_cache/cache_reg[1][113]  ( .D(\D_cache/n891 ), .CK(clk), .RN(n5783), .Q(\D_cache/cache[1][113] ), .QN(n814) );
  DFFRX1 \D_cache/cache_reg[2][113]  ( .D(\D_cache/n890 ), .CK(clk), .RN(n5783), .Q(\D_cache/cache[2][113] ), .QN(n2831) );
  DFFRX1 \D_cache/cache_reg[3][113]  ( .D(\D_cache/n889 ), .CK(clk), .RN(n5783), .Q(\D_cache/cache[3][113] ), .QN(n839) );
  DFFRX1 \D_cache/cache_reg[4][113]  ( .D(\D_cache/n888 ), .CK(clk), .RN(n5783), .Q(\D_cache/cache[4][113] ), .QN(n1577) );
  DFFRX1 \D_cache/cache_reg[5][113]  ( .D(\D_cache/n887 ), .CK(clk), .RN(n5783), .Q(\D_cache/cache[5][113] ), .QN(n3190) );
  DFFRX1 \D_cache/cache_reg[6][113]  ( .D(\D_cache/n886 ), .CK(clk), .RN(n5783), .Q(\D_cache/cache[6][113] ), .QN(n2832) );
  DFFRX1 \D_cache/cache_reg[7][113]  ( .D(\D_cache/n885 ), .CK(clk), .RN(n5784), .Q(\D_cache/cache[7][113] ), .QN(n840) );
  DFFRX1 \D_cache/cache_reg[0][114]  ( .D(\D_cache/n884 ), .CK(clk), .RN(n5784), .Q(\D_cache/cache[0][114] ), .QN(n960) );
  DFFRX1 \D_cache/cache_reg[1][114]  ( .D(\D_cache/n883 ), .CK(clk), .RN(n5784), .Q(\D_cache/cache[1][114] ), .QN(n2485) );
  DFFRX1 \D_cache/cache_reg[2][114]  ( .D(\D_cache/n882 ), .CK(clk), .RN(n5784), .Q(\D_cache/cache[2][114] ), .QN(n2447) );
  DFFRX1 \D_cache/cache_reg[3][114]  ( .D(\D_cache/n881 ), .CK(clk), .RN(n5784), .Q(\D_cache/cache[3][114] ), .QN(n472) );
  DFFRX1 \D_cache/cache_reg[4][114]  ( .D(\D_cache/n880 ), .CK(clk), .RN(n5784), .Q(\D_cache/cache[4][114] ), .QN(n1575) );
  DFFRX1 \D_cache/cache_reg[5][114]  ( .D(\D_cache/n879 ), .CK(clk), .RN(n5784), .Q(\D_cache/cache[5][114] ), .QN(n3188) );
  DFFRX1 \D_cache/cache_reg[6][114]  ( .D(\D_cache/n878 ), .CK(clk), .RN(n5784), .Q(\D_cache/cache[6][114] ), .QN(n1450) );
  DFFRX1 \D_cache/cache_reg[7][114]  ( .D(\D_cache/n877 ), .CK(clk), .RN(n5784), .Q(\D_cache/cache[7][114] ), .QN(n3063) );
  DFFRX1 \D_cache/cache_reg[0][115]  ( .D(\D_cache/n876 ), .CK(clk), .RN(n5784), .Q(\D_cache/cache[0][115] ), .QN(n959) );
  DFFRX1 \D_cache/cache_reg[1][115]  ( .D(\D_cache/n875 ), .CK(clk), .RN(n5784), .Q(\D_cache/cache[1][115] ), .QN(n2484) );
  DFFRX1 \D_cache/cache_reg[2][115]  ( .D(\D_cache/n874 ), .CK(clk), .RN(n5784), .Q(\D_cache/cache[2][115] ), .QN(n958) );
  DFFRX1 \D_cache/cache_reg[3][115]  ( .D(\D_cache/n873 ), .CK(clk), .RN(n5785), .Q(\D_cache/cache[3][115] ), .QN(n2483) );
  DFFRX1 \D_cache/cache_reg[4][115]  ( .D(\D_cache/n872 ), .CK(clk), .RN(n5785), .Q(\D_cache/cache[4][115] ), .QN(n1573) );
  DFFRX1 \D_cache/cache_reg[5][115]  ( .D(\D_cache/n871 ), .CK(clk), .RN(n5785), .Q(\D_cache/cache[5][115] ), .QN(n3186) );
  DFFRX1 \D_cache/cache_reg[6][115]  ( .D(\D_cache/n870 ), .CK(clk), .RN(n5785), .Q(\D_cache/cache[6][115] ), .QN(n1446) );
  DFFRX1 \D_cache/cache_reg[7][115]  ( .D(\D_cache/n869 ), .CK(clk), .RN(n5785), .Q(\D_cache/cache[7][115] ), .QN(n3059) );
  DFFRX1 \D_cache/cache_reg[0][116]  ( .D(\D_cache/n868 ), .CK(clk), .RN(n5785), .Q(\D_cache/cache[0][116] ), .QN(n1383) );
  DFFRX1 \D_cache/cache_reg[1][116]  ( .D(\D_cache/n867 ), .CK(clk), .RN(n5785), .Q(\D_cache/cache[1][116] ), .QN(n2996) );
  DFFRX1 \D_cache/cache_reg[2][116]  ( .D(\D_cache/n866 ), .CK(clk), .RN(n5785), .Q(\D_cache/cache[2][116] ), .QN(n1382) );
  DFFRX1 \D_cache/cache_reg[3][116]  ( .D(\D_cache/n865 ), .CK(clk), .RN(n5785), .Q(\D_cache/cache[3][116] ), .QN(n2995) );
  DFFRX1 \D_cache/cache_reg[4][116]  ( .D(\D_cache/n864 ), .CK(clk), .RN(n5785), .Q(\D_cache/cache[4][116] ), .QN(n1467) );
  DFFRX1 \D_cache/cache_reg[5][116]  ( .D(\D_cache/n863 ), .CK(clk), .RN(n5785), .Q(\D_cache/cache[5][116] ), .QN(n3080) );
  DFFRX1 \D_cache/cache_reg[6][116]  ( .D(\D_cache/n862 ), .CK(clk), .RN(n5785), .Q(\D_cache/cache[6][116] ), .QN(n1523) );
  DFFRX1 \D_cache/cache_reg[7][116]  ( .D(\D_cache/n861 ), .CK(clk), .RN(n5786), .Q(\D_cache/cache[7][116] ), .QN(n3136) );
  DFFRX1 \D_cache/cache_reg[0][117]  ( .D(\D_cache/n860 ), .CK(clk), .RN(n5786), .Q(\D_cache/cache[0][117] ), .QN(n1507) );
  DFFRX1 \D_cache/cache_reg[1][117]  ( .D(\D_cache/n859 ), .CK(clk), .RN(n5786), .Q(\D_cache/cache[1][117] ), .QN(n3120) );
  DFFRX1 \D_cache/cache_reg[2][117]  ( .D(\D_cache/n858 ), .CK(clk), .RN(n5786), .Q(\D_cache/cache[2][117] ), .QN(n2828) );
  DFFRX1 \D_cache/cache_reg[3][117]  ( .D(\D_cache/n857 ), .CK(clk), .RN(n5786), .Q(\D_cache/cache[3][117] ), .QN(n836) );
  DFFRX1 \D_cache/cache_reg[4][117]  ( .D(\D_cache/n856 ), .CK(clk), .RN(n5786), .Q(\D_cache/cache[4][117] ), .QN(n2413) );
  DFFRX1 \D_cache/cache_reg[5][117]  ( .D(\D_cache/n855 ), .CK(clk), .RN(n5786), .Q(\D_cache/cache[5][117] ), .QN(n384) );
  DFFRX1 \D_cache/cache_reg[6][117]  ( .D(\D_cache/n854 ), .CK(clk), .RN(n5786), .Q(\D_cache/cache[6][117] ), .QN(n2829) );
  DFFRX1 \D_cache/cache_reg[7][117]  ( .D(\D_cache/n853 ), .CK(clk), .RN(n5786), .Q(\D_cache/cache[7][117] ), .QN(n837) );
  DFFRX1 \D_cache/cache_reg[0][118]  ( .D(\D_cache/n852 ), .CK(clk), .RN(n5786), .Q(\D_cache/cache[0][118] ), .QN(n1389) );
  DFFRX1 \D_cache/cache_reg[1][118]  ( .D(\D_cache/n851 ), .CK(clk), .RN(n5786), .Q(\D_cache/cache[1][118] ), .QN(n3002) );
  DFFRX1 \D_cache/cache_reg[2][118]  ( .D(\D_cache/n850 ), .CK(clk), .RN(n5786), .Q(\D_cache/cache[2][118] ), .QN(n1388) );
  DFFRX1 \D_cache/cache_reg[3][118]  ( .D(\D_cache/n849 ), .CK(clk), .RN(n5787), .Q(\D_cache/cache[3][118] ), .QN(n3001) );
  DFFRX1 \D_cache/cache_reg[4][118]  ( .D(\D_cache/n848 ), .CK(clk), .RN(n5787), .Q(\D_cache/cache[4][118] ), .QN(n2830) );
  DFFRX1 \D_cache/cache_reg[5][118]  ( .D(\D_cache/n847 ), .CK(clk), .RN(n5787), .Q(\D_cache/cache[5][118] ), .QN(n838) );
  DFFRX1 \D_cache/cache_reg[6][118]  ( .D(\D_cache/n846 ), .CK(clk), .RN(n5787), .Q(\D_cache/cache[6][118] ), .QN(n1456) );
  DFFRX1 \D_cache/cache_reg[7][118]  ( .D(\D_cache/n845 ), .CK(clk), .RN(n5787), .Q(\D_cache/cache[7][118] ), .QN(n3069) );
  DFFRX1 \D_cache/cache_reg[0][119]  ( .D(\D_cache/n844 ), .CK(clk), .RN(n5787), .Q(\D_cache/cache[0][119] ), .QN(n1367) );
  DFFRX1 \D_cache/cache_reg[1][119]  ( .D(\D_cache/n843 ), .CK(clk), .RN(n5787), .Q(\D_cache/cache[1][119] ), .QN(n2980) );
  DFFRX1 \D_cache/cache_reg[2][119]  ( .D(\D_cache/n842 ), .CK(clk), .RN(n5787), .Q(\D_cache/cache[2][119] ), .QN(n1366) );
  DFFRX1 \D_cache/cache_reg[3][119]  ( .D(\D_cache/n841 ), .CK(clk), .RN(n5787), .Q(\D_cache/cache[3][119] ), .QN(n2979) );
  DFFRX1 \D_cache/cache_reg[4][119]  ( .D(\D_cache/n840 ), .CK(clk), .RN(n5787), .Q(\D_cache/cache[4][119] ), .QN(n2822) );
  DFFRX1 \D_cache/cache_reg[5][119]  ( .D(\D_cache/n839 ), .CK(clk), .RN(n5787), .Q(\D_cache/cache[5][119] ), .QN(n830) );
  DFFRX1 \D_cache/cache_reg[6][119]  ( .D(\D_cache/n838 ), .CK(clk), .RN(n5787), .Q(\D_cache/cache[6][119] ), .QN(n1443) );
  DFFRX1 \D_cache/cache_reg[7][119]  ( .D(\D_cache/n837 ), .CK(clk), .RN(n5788), .Q(\D_cache/cache[7][119] ), .QN(n3056) );
  DFFRX1 \D_cache/cache_reg[0][120]  ( .D(\D_cache/n836 ), .CK(clk), .RN(n5788), .Q(\D_cache/cache[0][120] ), .QN(n2820) );
  DFFRX1 \D_cache/cache_reg[1][120]  ( .D(\D_cache/n835 ), .CK(clk), .RN(n5788), .Q(\D_cache/cache[1][120] ), .QN(n828) );
  DFFRX1 \D_cache/cache_reg[2][120]  ( .D(\D_cache/n834 ), .CK(clk), .RN(n5788), .Q(\D_cache/cache[2][120] ), .QN(n2819) );
  DFFRX1 \D_cache/cache_reg[3][120]  ( .D(\D_cache/n833 ), .CK(clk), .RN(n5788), .Q(\D_cache/cache[3][120] ), .QN(n827) );
  DFFRX1 \D_cache/cache_reg[4][120]  ( .D(\D_cache/n832 ), .CK(clk), .RN(n5788), .Q(\D_cache/cache[4][120] ), .QN(n2821) );
  DFFRX1 \D_cache/cache_reg[5][120]  ( .D(\D_cache/n831 ), .CK(clk), .RN(n5788), .Q(\D_cache/cache[5][120] ), .QN(n829) );
  DFFRX1 \D_cache/cache_reg[6][120]  ( .D(\D_cache/n830 ), .CK(clk), .RN(n5788), .Q(\D_cache/cache[6][120] ), .QN(n1513) );
  DFFRX1 \D_cache/cache_reg[7][120]  ( .D(\D_cache/n829 ), .CK(clk), .RN(n5788), .Q(\D_cache/cache[7][120] ), .QN(n3126) );
  DFFRX1 \D_cache/cache_reg[0][121]  ( .D(\D_cache/n828 ), .CK(clk), .RN(n5788), .Q(\D_cache/cache[0][121] ), .QN(n1461) );
  DFFRX1 \D_cache/cache_reg[1][121]  ( .D(\D_cache/n827 ), .CK(clk), .RN(n5788), .Q(\D_cache/cache[1][121] ), .QN(n3074) );
  DFFRX1 \D_cache/cache_reg[2][121]  ( .D(\D_cache/n826 ), .CK(clk), .RN(n5788), .Q(\D_cache/cache[2][121] ), .QN(n1396) );
  DFFRX1 \D_cache/cache_reg[3][121]  ( .D(\D_cache/n825 ), .CK(clk), .RN(n5789), .Q(\D_cache/cache[3][121] ), .QN(n3009) );
  DFFRX1 \D_cache/cache_reg[4][121]  ( .D(\D_cache/n824 ), .CK(clk), .RN(n5789), .Q(\D_cache/cache[4][121] ), .QN(n1397) );
  DFFRX1 \D_cache/cache_reg[5][121]  ( .D(\D_cache/n823 ), .CK(clk), .RN(n5789), .Q(\D_cache/cache[5][121] ), .QN(n3010) );
  DFFRX1 \D_cache/cache_reg[6][121]  ( .D(\D_cache/n822 ), .CK(clk), .RN(n5789), .Q(\D_cache/cache[6][121] ), .QN(n1478) );
  DFFRX1 \D_cache/cache_reg[7][121]  ( .D(\D_cache/n821 ), .CK(clk), .RN(n5789), .Q(\D_cache/cache[7][121] ), .QN(n3091) );
  DFFRX1 \D_cache/cache_reg[0][122]  ( .D(\D_cache/n820 ), .CK(clk), .RN(n5789), .Q(\D_cache/cache[0][122] ), .QN(n2407) );
  DFFRX1 \D_cache/cache_reg[1][122]  ( .D(\D_cache/n819 ), .CK(clk), .RN(n5789), .Q(\D_cache/cache[1][122] ), .QN(n901) );
  DFFRX1 \D_cache/cache_reg[2][122]  ( .D(\D_cache/n818 ), .CK(clk), .RN(n5789), .Q(\D_cache/cache[2][122] ), .QN(n933) );
  DFFRX1 \D_cache/cache_reg[3][122]  ( .D(\D_cache/n817 ), .CK(clk), .RN(n5789), .Q(\D_cache/cache[3][122] ), .QN(n2457) );
  DFFRX1 \D_cache/cache_reg[4][122]  ( .D(\D_cache/n816 ), .CK(clk), .RN(n5789), .Q(\D_cache/cache[4][122] ), .QN(n2443) );
  DFFRX1 \D_cache/cache_reg[5][122]  ( .D(\D_cache/n815 ), .CK(clk), .RN(n5789), .Q(\D_cache/cache[5][122] ), .QN(n468) );
  DFFRX1 \D_cache/cache_reg[6][122]  ( .D(\D_cache/n814 ), .CK(clk), .RN(n5789), .Q(\D_cache/cache[6][122] ), .QN(n2440) );
  DFFRX1 \D_cache/cache_reg[7][122]  ( .D(\D_cache/n813 ), .CK(clk), .RN(n5790), .Q(\D_cache/cache[7][122] ), .QN(n464) );
  DFFRX1 \D_cache/cache_reg[0][123]  ( .D(\D_cache/n812 ), .CK(clk), .RN(n5790), .Q(\D_cache/cache[0][123] ), .QN(n945) );
  DFFRX1 \D_cache/cache_reg[1][123]  ( .D(\D_cache/n811 ), .CK(clk), .RN(n5790), .Q(\D_cache/cache[1][123] ), .QN(n2470) );
  DFFRX1 \D_cache/cache_reg[2][123]  ( .D(\D_cache/n810 ), .CK(clk), .RN(n5790), .Q(\D_cache/cache[2][123] ), .QN(n1380) );
  DFFRX1 \D_cache/cache_reg[3][123]  ( .D(\D_cache/n809 ), .CK(clk), .RN(n5790), .Q(\D_cache/cache[3][123] ), .QN(n2993) );
  DFFRX1 \D_cache/cache_reg[4][123]  ( .D(\D_cache/n808 ), .CK(clk), .RN(n5790), .Q(\D_cache/cache[4][123] ), .QN(n946) );
  DFFRX1 \D_cache/cache_reg[5][123]  ( .D(\D_cache/n807 ), .CK(clk), .RN(n5790), .Q(\D_cache/cache[5][123] ), .QN(n2471) );
  DFFRX1 \D_cache/cache_reg[6][123]  ( .D(\D_cache/n806 ), .CK(clk), .RN(n5790), .Q(\D_cache/cache[6][123] ), .QN(n1445) );
  DFFRX1 \D_cache/cache_reg[7][123]  ( .D(\D_cache/n805 ), .CK(clk), .RN(n5790), .Q(\D_cache/cache[7][123] ), .QN(n3058) );
  DFFRX1 \D_cache/cache_reg[0][124]  ( .D(\D_cache/n804 ), .CK(clk), .RN(n5790), .Q(\D_cache/cache[0][124] ), .QN(n2817) );
  DFFRX1 \D_cache/cache_reg[1][124]  ( .D(\D_cache/n803 ), .CK(clk), .RN(n5790), .Q(\D_cache/cache[1][124] ), .QN(n825) );
  DFFRX1 \D_cache/cache_reg[2][124]  ( .D(\D_cache/n802 ), .CK(clk), .RN(n5790), .Q(\D_cache/cache[2][124] ), .QN(n2816) );
  DFFRX1 \D_cache/cache_reg[3][124]  ( .D(\D_cache/n801 ), .CK(clk), .RN(n5791), .Q(\D_cache/cache[3][124] ), .QN(n824) );
  DFFRX1 \D_cache/cache_reg[4][124]  ( .D(\D_cache/n800 ), .CK(clk), .RN(n5791), .Q(\D_cache/cache[4][124] ), .QN(n2818) );
  DFFRX1 \D_cache/cache_reg[5][124]  ( .D(\D_cache/n799 ), .CK(clk), .RN(n5791), .Q(\D_cache/cache[5][124] ), .QN(n826) );
  DFFRX1 \D_cache/cache_reg[6][124]  ( .D(\D_cache/n798 ), .CK(clk), .RN(n5791), .Q(\D_cache/cache[6][124] ), .QN(n1492) );
  DFFRX1 \D_cache/cache_reg[7][124]  ( .D(\D_cache/n797 ), .CK(clk), .RN(n5791), .Q(\D_cache/cache[7][124] ), .QN(n3105) );
  DFFRX1 \D_cache/cache_reg[0][125]  ( .D(\D_cache/n796 ), .CK(clk), .RN(n5791), .Q(\D_cache/cache[0][125] ), .QN(n1387) );
  DFFRX1 \D_cache/cache_reg[1][125]  ( .D(\D_cache/n795 ), .CK(clk), .RN(n5791), .Q(\D_cache/cache[1][125] ), .QN(n3000) );
  DFFRX1 \D_cache/cache_reg[2][125]  ( .D(\D_cache/n794 ), .CK(clk), .RN(n5791), .Q(\D_cache/cache[2][125] ), .QN(n1386) );
  DFFRX1 \D_cache/cache_reg[3][125]  ( .D(\D_cache/n793 ), .CK(clk), .RN(n5791), .Q(\D_cache/cache[3][125] ), .QN(n2999) );
  DFFRX1 \D_cache/cache_reg[4][125]  ( .D(\D_cache/n792 ), .CK(clk), .RN(n5791), .Q(\D_cache/cache[4][125] ), .QN(n2827) );
  DFFRX1 \D_cache/cache_reg[5][125]  ( .D(\D_cache/n791 ), .CK(clk), .RN(n5791), .Q(\D_cache/cache[5][125] ), .QN(n835) );
  DFFRX1 \D_cache/cache_reg[6][125]  ( .D(\D_cache/n790 ), .CK(clk), .RN(n5791), .Q(\D_cache/cache[6][125] ), .QN(n2808) );
  DFFRX1 \D_cache/cache_reg[7][125]  ( .D(\D_cache/n789 ), .CK(clk), .RN(n5792), .Q(\D_cache/cache[7][125] ), .QN(n806) );
  DFFRX1 \D_cache/cache_reg[0][126]  ( .D(\D_cache/n788 ), .CK(clk), .RN(n5792), .Q(\D_cache/cache[0][126] ), .QN(n815) );
  DFFRX1 \D_cache/cache_reg[1][126]  ( .D(\D_cache/n787 ), .CK(clk), .RN(n5792), .Q(\D_cache/cache[1][126] ), .QN(n2347) );
  DFFRX1 \D_cache/cache_reg[2][126]  ( .D(\D_cache/n786 ), .CK(clk), .RN(n5792), .Q(\D_cache/cache[2][126] ), .QN(n809) );
  DFFRX1 \D_cache/cache_reg[3][126]  ( .D(\D_cache/n785 ), .CK(clk), .RN(n5792), .Q(\D_cache/cache[3][126] ), .QN(n2342) );
  DFFRX1 \D_cache/cache_reg[4][126]  ( .D(\D_cache/n784 ), .CK(clk), .RN(n5792), .Q(\D_cache/cache[4][126] ), .QN(n810) );
  DFFRX1 \D_cache/cache_reg[5][126]  ( .D(\D_cache/n783 ), .CK(clk), .RN(n5792), .Q(\D_cache/cache[5][126] ), .QN(n2343) );
  DFFRX1 \D_cache/cache_reg[6][126]  ( .D(\D_cache/n782 ), .CK(clk), .RN(n5792), .Q(\D_cache/cache[6][126] ), .QN(n808) );
  DFFRX1 \D_cache/cache_reg[7][126]  ( .D(\D_cache/n781 ), .CK(clk), .RN(n5792), .Q(\D_cache/cache[7][126] ), .QN(n2341) );
  DFFRX1 \D_cache/cache_reg[0][127]  ( .D(\D_cache/n780 ), .CK(clk), .RN(n5792), .Q(\D_cache/cache[0][127] ), .QN(n1361) );
  DFFRX1 \D_cache/cache_reg[1][127]  ( .D(\D_cache/n779 ), .CK(clk), .RN(n5792), .Q(\D_cache/cache[1][127] ), .QN(n2974) );
  DFFRX1 \D_cache/cache_reg[2][127]  ( .D(\D_cache/n778 ), .CK(clk), .RN(n5792), .Q(\D_cache/cache[2][127] ), .QN(n1362) );
  DFFRX1 \D_cache/cache_reg[3][127]  ( .D(\D_cache/n777 ), .CK(clk), .RN(n5793), .Q(\D_cache/cache[3][127] ), .QN(n2975) );
  DFFRX1 \D_cache/cache_reg[4][127]  ( .D(\D_cache/n776 ), .CK(clk), .RN(n5793), .Q(\D_cache/cache[4][127] ), .QN(n1363) );
  DFFRX1 \D_cache/cache_reg[5][127]  ( .D(\D_cache/n775 ), .CK(clk), .RN(n5793), .Q(\D_cache/cache[5][127] ), .QN(n2976) );
  DFFRX1 \D_cache/cache_reg[6][127]  ( .D(\D_cache/n774 ), .CK(clk), .RN(n5793), .Q(\D_cache/cache[6][127] ), .QN(n1556) );
  DFFRX1 \D_cache/cache_reg[7][127]  ( .D(\D_cache/n773 ), .CK(clk), .RN(n5793), .Q(\D_cache/cache[7][127] ), .QN(n3169) );
  DFFRX1 \D_cache/cache_reg[0][128]  ( .D(\D_cache/n772 ), .CK(clk), .RN(n5793), .Q(\D_cache/cache[0][128] ), .QN(n1226) );
  DFFRX1 \D_cache/cache_reg[1][128]  ( .D(\D_cache/n771 ), .CK(clk), .RN(n5793), .Q(\D_cache/cache[1][128] ), .QN(n2805) );
  DFFRX1 \D_cache/cache_reg[2][128]  ( .D(\D_cache/n770 ), .CK(clk), .RN(n5793), .Q(\D_cache/cache[2][128] ), .QN(n1960) );
  DFFRX1 \D_cache/cache_reg[3][128]  ( .D(\D_cache/n769 ), .CK(clk), .RN(n5793), .Q(\D_cache/cache[3][128] ), .QN(n388) );
  DFFRX1 \D_cache/cache_reg[6][128]  ( .D(\D_cache/n766 ), .CK(clk), .RN(n5793), .Q(\D_cache/cache[6][128] ), .QN(n1862) );
  DFFRX1 \D_cache/cache_reg[0][129]  ( .D(\D_cache/n764 ), .CK(clk), .RN(n5794), .Q(\D_cache/cache[0][129] ), .QN(n1882) );
  DFFRX1 \D_cache/cache_reg[1][129]  ( .D(\D_cache/n763 ), .CK(clk), .RN(n5794), .Q(\D_cache/cache[1][129] ), .QN(n316) );
  DFFRX1 \D_cache/cache_reg[4][129]  ( .D(\D_cache/n760 ), .CK(clk), .RN(n5794), .Q(\D_cache/cache[4][129] ), .QN(n2025) );
  DFFRX1 \D_cache/cache_reg[5][129]  ( .D(\D_cache/n759 ), .CK(clk), .RN(n5794), .Q(\D_cache/cache[5][129] ), .QN(n2023) );
  DFFRX1 \D_cache/cache_reg[0][130]  ( .D(\D_cache/n756 ), .CK(clk), .RN(n5794), .Q(\D_cache/cache[0][130] ), .QN(n1879) );
  DFFRX1 \D_cache/cache_reg[1][130]  ( .D(\D_cache/n755 ), .CK(clk), .RN(n5794), .Q(\D_cache/cache[1][130] ), .QN(n1892) );
  DFFRX1 \D_cache/cache_reg[4][130]  ( .D(\D_cache/n752 ), .CK(clk), .RN(n5795), .Q(\D_cache/cache[4][130] ), .QN(n322) );
  DFFRX1 \D_cache/cache_reg[0][131]  ( .D(\D_cache/n748 ), .CK(clk), .RN(n5795), .Q(\D_cache/cache[0][131] ), .QN(n2020) );
  DFFRX1 \D_cache/cache_reg[1][131]  ( .D(\D_cache/n747 ), .CK(clk), .RN(n5795), .Q(\D_cache/cache[1][131] ), .QN(n1989) );
  DFFRX1 \D_cache/cache_reg[4][131]  ( .D(\D_cache/n744 ), .CK(clk), .RN(n5795), .Q(\D_cache/cache[4][131] ), .QN(n2019) );
  DFFRX1 \D_cache/cache_reg[0][132]  ( .D(\D_cache/n740 ), .CK(clk), .RN(n5796), .Q(\D_cache/cache[0][132] ), .QN(n2046) );
  DFFRX1 \D_cache/cache_reg[1][132]  ( .D(\D_cache/n739 ), .CK(clk), .RN(n5796), .Q(\D_cache/cache[1][132] ), .QN(n706) );
  DFFRX1 \D_cache/cache_reg[2][132]  ( .D(\D_cache/n738 ), .CK(clk), .RN(n5796), .Q(\D_cache/cache[2][132] ), .QN(n1937) );
  DFFRX1 \D_cache/cache_reg[3][132]  ( .D(\D_cache/n737 ), .CK(clk), .RN(n5796), .Q(\D_cache/cache[3][132] ), .QN(n357) );
  DFFRX1 \D_cache/cache_reg[4][132]  ( .D(\D_cache/n736 ), .CK(clk), .RN(n5796), .Q(\D_cache/cache[4][132] ), .QN(n1616) );
  DFFRX1 \D_cache/cache_reg[5][132]  ( .D(\D_cache/n735 ), .CK(clk), .RN(n5796), .Q(\D_cache/cache[5][132] ), .QN(n281) );
  DFFRX1 \D_cache/cache_reg[6][132]  ( .D(\D_cache/n734 ), .CK(clk), .RN(n5796), .Q(\D_cache/cache[6][132] ), .QN(n1974) );
  DFFRX1 \D_cache/cache_reg[0][133]  ( .D(\D_cache/n732 ), .CK(clk), .RN(n5796), .Q(\D_cache/cache[0][133] ), .QN(n3196) );
  DFFRX1 \D_cache/cache_reg[1][133]  ( .D(\D_cache/n731 ), .CK(clk), .RN(n5796), .Q(\D_cache/cache[1][133] ), .QN(n1880) );
  DFFRX1 \D_cache/cache_reg[2][133]  ( .D(\D_cache/n730 ), .CK(clk), .RN(n5796), .Q(\D_cache/cache[2][133] ) );
  DFFRX1 \D_cache/cache_reg[4][133]  ( .D(\D_cache/n728 ), .CK(clk), .RN(n5797), .Q(\D_cache/cache[4][133] ), .QN(n2048) );
  DFFRX1 \D_cache/cache_reg[5][133]  ( .D(\D_cache/n727 ), .CK(clk), .RN(n5797), .Q(\D_cache/cache[5][133] ), .QN(n320) );
  DFFRX1 \D_cache/cache_reg[0][134]  ( .D(\D_cache/n724 ), .CK(clk), .RN(n5797), .Q(\D_cache/cache[0][134] ), .QN(n2798) );
  DFFRX1 \D_cache/cache_reg[1][134]  ( .D(\D_cache/n723 ), .CK(clk), .RN(n5797), .Q(\D_cache/cache[1][134] ), .QN(n2415) );
  DFFRX1 \D_cache/cache_reg[2][134]  ( .D(\D_cache/n722 ), .CK(clk), .RN(n5797), .Q(\D_cache/cache[2][134] ), .QN(n451) );
  DFFRX1 \D_cache/cache_reg[4][134]  ( .D(\D_cache/n720 ), .CK(clk), .RN(n5797), .Q(\D_cache/cache[4][134] ), .QN(n2795) );
  DFFRX1 \D_cache/cache_reg[5][134]  ( .D(\D_cache/n719 ), .CK(clk), .RN(n5797), .Q(\D_cache/cache[5][134] ), .QN(n2797) );
  DFFRX1 \D_cache/cache_reg[0][135]  ( .D(\D_cache/n716 ), .CK(clk), .RN(n5798), .Q(\D_cache/cache[0][135] ), .QN(n2041) );
  DFFRX1 \D_cache/cache_reg[1][135]  ( .D(\D_cache/n715 ), .CK(clk), .RN(n5798), .Q(\D_cache/cache[1][135] ), .QN(n279) );
  DFFRX1 \D_cache/cache_reg[2][135]  ( .D(\D_cache/n714 ), .CK(clk), .RN(n5798), .Q(\D_cache/cache[2][135] ), .QN(n1938) );
  DFFRX1 \D_cache/cache_reg[3][135]  ( .D(\D_cache/n713 ), .CK(clk), .RN(n5798), .Q(\D_cache/cache[3][135] ), .QN(n358) );
  DFFRX1 \D_cache/cache_reg[4][135]  ( .D(\D_cache/n712 ), .CK(clk), .RN(n5798), .Q(\D_cache/cache[4][135] ), .QN(n2045) );
  DFFRX1 \D_cache/cache_reg[5][135]  ( .D(\D_cache/n711 ), .CK(clk), .RN(n5798), .Q(\D_cache/cache[5][135] ), .QN(n705) );
  DFFRX1 \D_cache/cache_reg[6][135]  ( .D(\D_cache/n710 ), .CK(clk), .RN(n5798), .Q(\D_cache/cache[6][135] ), .QN(n424) );
  DFFRX1 \D_cache/cache_reg[0][136]  ( .D(\D_cache/n708 ), .CK(clk), .RN(n5798), .Q(\D_cache/cache[0][136] ), .QN(n2043) );
  DFFRX1 \D_cache/cache_reg[1][136]  ( .D(\D_cache/n707 ), .CK(clk), .RN(n5798), .Q(\D_cache/cache[1][136] ), .QN(n703) );
  DFFRX1 \D_cache/cache_reg[4][136]  ( .D(\D_cache/n704 ), .CK(clk), .RN(n5799), .Q(\D_cache/cache[4][136] ), .QN(n2044) );
  DFFRX1 \D_cache/cache_reg[5][136]  ( .D(\D_cache/n703 ), .CK(clk), .RN(n5799), .Q(\D_cache/cache[5][136] ), .QN(n704) );
  DFFRX1 \D_cache/cache_reg[6][136]  ( .D(\D_cache/n702 ), .CK(clk), .RN(n5799), .Q(\D_cache/cache[6][136] ), .QN(n421) );
  DFFRX1 \D_cache/cache_reg[7][136]  ( .D(\D_cache/n701 ), .CK(clk), .RN(n5799), .Q(\D_cache/cache[7][136] ), .QN(n3261) );
  DFFRX1 \D_cache/cache_reg[0][137]  ( .D(\D_cache/n700 ), .CK(clk), .RN(n5799), .Q(\D_cache/cache[0][137] ), .QN(n712) );
  DFFRX1 \D_cache/cache_reg[1][137]  ( .D(\D_cache/n699 ), .CK(clk), .RN(n5799), .Q(\D_cache/cache[1][137] ), .QN(n3249) );
  DFFRX1 \D_cache/cache_reg[2][137]  ( .D(\D_cache/n698 ), .CK(clk), .RN(n5799), .Q(\D_cache/cache[2][137] ), .QN(n1943) );
  DFFRX1 \D_cache/cache_reg[3][137]  ( .D(\D_cache/n697 ), .CK(clk), .RN(n5799), .Q(\D_cache/cache[3][137] ), .QN(n365) );
  DFFRX1 \D_cache/cache_reg[4][137]  ( .D(\D_cache/n696 ), .CK(clk), .RN(n5799), .Q(\D_cache/cache[4][137] ), .QN(n713) );
  DFFRX1 \D_cache/cache_reg[5][137]  ( .D(\D_cache/n695 ), .CK(clk), .RN(n5799), .Q(\D_cache/cache[5][137] ), .QN(n3250) );
  DFFRX1 \D_cache/cache_reg[6][137]  ( .D(\D_cache/n694 ), .CK(clk), .RN(n5799), .Q(\D_cache/cache[6][137] ), .QN(n423) );
  DFFRX1 \D_cache/cache_reg[0][138]  ( .D(\D_cache/n692 ), .CK(clk), .RN(n5800), .Q(\D_cache/cache[0][138] ), .QN(n2796) );
  DFFRX1 \D_cache/cache_reg[1][138]  ( .D(\D_cache/n691 ), .CK(clk), .RN(n5800), .Q(\D_cache/cache[1][138] ) );
  DFFRX1 \D_cache/cache_reg[4][138]  ( .D(\D_cache/n688 ), .CK(clk), .RN(n5800), .Q(\D_cache/cache[4][138] ), .QN(n2801) );
  DFFRX1 \D_cache/cache_reg[5][138]  ( .D(\D_cache/n687 ), .CK(clk), .RN(n5800), .Q(\D_cache/cache[5][138] ), .QN(n735) );
  DFFRX1 \D_cache/cache_reg[0][139]  ( .D(\D_cache/n684 ), .CK(clk), .RN(n5800), .Q(\D_cache/cache[0][139] ), .QN(n1887) );
  DFFRX1 \D_cache/cache_reg[4][139]  ( .D(\D_cache/n680 ), .CK(clk), .RN(n5801), .Q(\D_cache/cache[4][139] ), .QN(n1990) );
  DFFRX1 \D_cache/cache_reg[0][141]  ( .D(\D_cache/n668 ), .CK(clk), .RN(n5802), .Q(\D_cache/cache[0][141] ), .QN(n2350) );
  DFFRX1 \D_cache/cache_reg[1][141]  ( .D(\D_cache/n667 ), .CK(clk), .RN(n5802), .Q(\D_cache/cache[1][141] ) );
  DFFRX1 \D_cache/cache_reg[2][141]  ( .D(\D_cache/n666 ), .CK(clk), .RN(n5802), .Q(\D_cache/cache[2][141] ), .QN(n449) );
  DFFRX1 \D_cache/cache_reg[3][141]  ( .D(\D_cache/n665 ), .CK(clk), .RN(n5802), .Q(\D_cache/cache[3][141] ), .QN(n3291) );
  DFFRX1 \D_cache/cache_reg[4][141]  ( .D(\D_cache/n664 ), .CK(clk), .RN(n5802), .Q(\D_cache/cache[4][141] ), .QN(n1225) );
  DFFRX1 \D_cache/cache_reg[5][141]  ( .D(\D_cache/n663 ), .CK(clk), .RN(n5802), .Q(\D_cache/cache[5][141] ), .QN(n2804) );
  DFFRX1 \D_cache/cache_reg[6][141]  ( .D(\D_cache/n662 ), .CK(clk), .RN(n5802), .Q(\D_cache/cache[6][141] ), .QN(n1956) );
  DFFRX1 \D_cache/cache_reg[7][141]  ( .D(\D_cache/n661 ), .CK(clk), .RN(n5802), .Q(\D_cache/cache[7][141] ), .QN(n381) );
  DFFRX1 \D_cache/cache_reg[0][142]  ( .D(\D_cache/n660 ), .CK(clk), .RN(n5802), .Q(\D_cache/cache[0][142] ), .QN(n2018) );
  DFFRX1 \D_cache/cache_reg[4][142]  ( .D(\D_cache/n656 ), .CK(clk), .RN(n5803), .Q(\D_cache/cache[4][142] ), .QN(n2024) );
  DFFRX1 \D_cache/cache_reg[5][142]  ( .D(\D_cache/n655 ), .CK(clk), .RN(n5803), .Q(\D_cache/cache[5][142] ), .QN(n1988) );
  DFFRX1 \D_cache/cache_reg[0][143]  ( .D(\D_cache/n652 ), .CK(clk), .RN(n5803), .Q(\D_cache/cache[0][143] ), .QN(n2047) );
  DFFRX1 \D_cache/cache_reg[1][143]  ( .D(\D_cache/n651 ), .CK(clk), .RN(n5803), .Q(\D_cache/cache[1][143] ), .QN(n707) );
  DFFRX1 \D_cache/cache_reg[2][143]  ( .D(\D_cache/n650 ), .CK(clk), .RN(n5803), .Q(\D_cache/cache[2][143] ), .QN(n450) );
  DFFRX1 \D_cache/cache_reg[3][143]  ( .D(\D_cache/n649 ), .CK(clk), .RN(n5803), .Q(\D_cache/cache[3][143] ), .QN(n2006) );
  DFFRX1 \D_cache/cache_reg[4][143]  ( .D(\D_cache/n648 ), .CK(clk), .RN(n5803), .Q(\D_cache/cache[4][143] ), .QN(n1227) );
  DFFRX1 \D_cache/cache_reg[5][143]  ( .D(\D_cache/n647 ), .CK(clk), .RN(n5803), .Q(\D_cache/cache[5][143] ), .QN(n2806) );
  DFFRX1 \D_cache/cache_reg[6][143]  ( .D(\D_cache/n646 ), .CK(clk), .RN(n5803), .Q(\D_cache/cache[6][143] ), .QN(n1946) );
  DFFRX1 \D_cache/cache_reg[7][143]  ( .D(\D_cache/n645 ), .CK(clk), .RN(n5803), .Q(\D_cache/cache[7][143] ), .QN(n368) );
  DFFRX1 \D_cache/cache_reg[0][145]  ( .D(\D_cache/n636 ), .CK(clk), .RN(n5804), .Q(\D_cache/cache[0][145] ), .QN(n2040) );
  DFFRX1 \D_cache/cache_reg[1][145]  ( .D(\D_cache/n635 ), .CK(clk), .RN(n5804), .Q(\D_cache/cache[1][145] ), .QN(n702) );
  DFFRX1 \D_cache/cache_reg[2][145]  ( .D(\D_cache/n634 ), .CK(clk), .RN(n5804), .Q(\D_cache/cache[2][145] ), .QN(n1629) );
  DFFRX1 \D_cache/cache_reg[3][145]  ( .D(\D_cache/n633 ), .CK(clk), .RN(n5804), .Q(\D_cache/cache[3][145] ), .QN(n3292) );
  DFFRX1 \D_cache/cache_reg[4][145]  ( .D(\D_cache/n632 ), .CK(clk), .RN(n5805), .Q(\D_cache/cache[4][145] ) );
  DFFRX1 \D_cache/cache_reg[5][145]  ( .D(\D_cache/n631 ), .CK(clk), .RN(n5805), .Q(\D_cache/cache[5][145] ) );
  DFFRX1 \D_cache/cache_reg[6][145]  ( .D(\D_cache/n630 ), .CK(clk), .RN(n5805), .Q(\D_cache/cache[6][145] ), .QN(n3288) );
  DFFRX1 \D_cache/cache_reg[7][145]  ( .D(\D_cache/n629 ), .CK(clk), .RN(n5805), .Q(\D_cache/cache[7][145] ), .QN(n439) );
  DFFRX1 \D_cache/cache_reg[0][146]  ( .D(\D_cache/n628 ), .CK(clk), .RN(n5805), .Q(\D_cache/cache[0][146] ), .QN(n2799) );
  DFFRX1 \D_cache/cache_reg[1][146]  ( .D(\D_cache/n627 ), .CK(clk), .RN(n5805), .Q(\D_cache/cache[1][146] ), .QN(n1893) );
  DFFRX1 \D_cache/cache_reg[2][146]  ( .D(\D_cache/n626 ), .CK(clk), .RN(n5805), .Q(\D_cache/cache[2][146] ), .QN(n313) );
  DFFRX1 \D_cache/cache_reg[4][146]  ( .D(\D_cache/n624 ), .CK(clk), .RN(n5805), .Q(\D_cache/cache[4][146] ), .QN(n2042) );
  DFFRX1 \D_cache/cache_reg[5][146]  ( .D(\D_cache/n623 ), .CK(clk), .RN(n5805), .Q(\D_cache/cache[5][146] ), .QN(n315) );
  DFFRX1 \D_cache/cache_reg[0][147]  ( .D(\D_cache/n620 ), .CK(clk), .RN(n5806), .Q(\D_cache/cache[0][147] ), .QN(n2049) );
  DFFRX1 \D_cache/cache_reg[1][147]  ( .D(\D_cache/n619 ), .CK(clk), .RN(n5806), .Q(\D_cache/cache[1][147] ), .QN(n708) );
  DFFRX1 \D_cache/cache_reg[2][147]  ( .D(\D_cache/n618 ), .CK(clk), .RN(n5806), .Q(\D_cache/cache[2][147] ), .QN(n1964) );
  DFFRX1 \D_cache/cache_reg[3][147]  ( .D(\D_cache/n617 ), .CK(clk), .RN(n5806), .Q(\D_cache/cache[3][147] ), .QN(n392) );
  DFFRX1 \D_cache/cache_reg[4][147]  ( .D(\D_cache/n616 ), .CK(clk), .RN(n5806), .Q(\D_cache/cache[4][147] ), .QN(n2051) );
  DFFRX1 \D_cache/cache_reg[5][147]  ( .D(\D_cache/n615 ), .CK(clk), .RN(n5806), .Q(\D_cache/cache[5][147] ), .QN(n710) );
  DFFRX1 \D_cache/cache_reg[6][147]  ( .D(\D_cache/n614 ), .CK(clk), .RN(n5806), .Q(\D_cache/cache[6][147] ), .QN(n1965) );
  DFFRX1 \D_cache/cache_reg[7][147]  ( .D(\D_cache/n613 ), .CK(clk), .RN(n5806), .Q(\D_cache/cache[7][147] ), .QN(n393) );
  DFFRX1 \D_cache/cache_reg[0][148]  ( .D(\D_cache/n612 ), .CK(clk), .RN(n5806), .Q(\D_cache/cache[0][148] ), .QN(n254) );
  DFFRX1 \D_cache/cache_reg[1][148]  ( .D(\D_cache/n611 ), .CK(clk), .RN(n5806), .Q(\D_cache/cache[1][148] ), .QN(n204) );
  DFFRX1 \D_cache/cache_reg[2][148]  ( .D(\D_cache/n610 ), .CK(clk), .RN(n5806), .Q(\D_cache/cache[2][148] ) );
  DFFRX1 \D_cache/cache_reg[3][148]  ( .D(\D_cache/n609 ), .CK(clk), .RN(n5806), .Q(\D_cache/cache[3][148] ), .QN(n1895) );
  DFFRX1 \D_cache/cache_reg[4][148]  ( .D(\D_cache/n608 ), .CK(clk), .RN(n5807), .Q(\D_cache/cache[4][148] ), .QN(n2022) );
  DFFRX1 \D_cache/cache_reg[6][148]  ( .D(\D_cache/n606 ), .CK(clk), .RN(n5807), .Q(\D_cache/cache[6][148] ), .QN(n1967) );
  DFFRX1 \D_cache/cache_reg[7][148]  ( .D(\D_cache/n605 ), .CK(clk), .RN(n5807), .Q(\D_cache/cache[7][148] ), .QN(n395) );
  DFFRX1 \D_cache/cache_reg[0][149]  ( .D(\D_cache/n604 ), .CK(clk), .RN(n5807), .Q(\D_cache/cache[0][149] ), .QN(n2050) );
  DFFRX1 \D_cache/cache_reg[1][149]  ( .D(\D_cache/n603 ), .CK(clk), .RN(n5807), .Q(\D_cache/cache[1][149] ), .QN(n709) );
  DFFRX1 \D_cache/cache_reg[2][149]  ( .D(\D_cache/n602 ), .CK(clk), .RN(n5807), .Q(\D_cache/cache[2][149] ), .QN(n977) );
  DFFRX1 \D_cache/cache_reg[3][149]  ( .D(\D_cache/n601 ), .CK(clk), .RN(n5807), .Q(\D_cache/cache[3][149] ), .QN(n2504) );
  DFFRX1 \D_cache/cache_reg[4][149]  ( .D(\D_cache/n600 ), .CK(clk), .RN(n5807), .Q(\D_cache/cache[4][149] ), .QN(n3258) );
  DFFRX1 \D_cache/cache_reg[5][149]  ( .D(\D_cache/n599 ), .CK(clk), .RN(n5807), .Q(\D_cache/cache[5][149] ), .QN(n1615) );
  DFFRX1 \D_cache/cache_reg[6][149]  ( .D(\D_cache/n598 ), .CK(clk), .RN(n5807), .Q(\D_cache/cache[6][149] ), .QN(n978) );
  DFFRX1 \D_cache/cache_reg[7][149]  ( .D(\D_cache/n597 ), .CK(clk), .RN(n5807), .Q(\D_cache/cache[7][149] ), .QN(n2505) );
  DFFRX1 \D_cache/cache_reg[0][150]  ( .D(\D_cache/n596 ), .CK(clk), .RN(n5808), .Q(\D_cache/cache[0][150] ), .QN(n1631) );
  DFFRX1 \D_cache/cache_reg[1][150]  ( .D(\D_cache/n595 ), .CK(clk), .RN(n5808), .Q(\D_cache/cache[1][150] ), .QN(n3296) );
  DFFRX1 \D_cache/cache_reg[2][150]  ( .D(\D_cache/n594 ), .CK(clk), .RN(n5808), .Q(\D_cache/cache[2][150] ), .QN(n2402) );
  DFFRX1 \D_cache/cache_reg[3][150]  ( .D(\D_cache/n593 ), .CK(clk), .RN(n5808), .Q(\D_cache/cache[3][150] ), .QN(n896) );
  DFFRX1 \D_cache/cache_reg[4][150]  ( .D(\D_cache/n592 ), .CK(clk), .RN(n5808), .Q(\D_cache/cache[4][150] ), .QN(n1628) );
  DFFRX1 \D_cache/cache_reg[5][150]  ( .D(\D_cache/n591 ), .CK(clk), .RN(n5808), .Q(\D_cache/cache[5][150] ), .QN(n3287) );
  DFFRX1 \D_cache/cache_reg[6][150]  ( .D(\D_cache/n590 ), .CK(clk), .RN(n5808), .Q(\D_cache/cache[6][150] ), .QN(n2404) );
  DFFRX1 \D_cache/cache_reg[7][150]  ( .D(\D_cache/n589 ), .CK(clk), .RN(n5808), .Q(\D_cache/cache[7][150] ), .QN(n898) );
  DFFRX1 \D_cache/cache_reg[0][151]  ( .D(\D_cache/n588 ), .CK(clk), .RN(n5808), .Q(\D_cache/cache[0][151] ), .QN(n280) );
  DFFRX1 \D_cache/cache_reg[1][151]  ( .D(\D_cache/n587 ), .CK(clk), .RN(n5808), .Q(\D_cache/cache[1][151] ), .QN(n1231) );
  DFFRX1 \D_cache/cache_reg[2][151]  ( .D(\D_cache/n586 ), .CK(clk), .RN(n5808), .Q(\D_cache/cache[2][151] ), .QN(n1959) );
  DFFRX1 \D_cache/cache_reg[3][151]  ( .D(\D_cache/n585 ), .CK(clk), .RN(n5808), .Q(\D_cache/cache[3][151] ), .QN(n387) );
  DFFRX1 \D_cache/cache_reg[4][151]  ( .D(\D_cache/n584 ), .CK(clk), .RN(n5809), .Q(\D_cache/cache[4][151] ), .QN(n711) );
  DFFRX1 \D_cache/cache_reg[5][151]  ( .D(\D_cache/n583 ), .CK(clk), .RN(n5809), .Q(\D_cache/cache[5][151] ), .QN(n221) );
  DFFRX1 \D_cache/cache_reg[6][151]  ( .D(\D_cache/n582 ), .CK(clk), .RN(n5809), .Q(\D_cache/cache[6][151] ), .QN(n422) );
  DFFRX1 \D_cache/cache_reg[7][151]  ( .D(\D_cache/n581 ), .CK(clk), .RN(n5809), .Q(\D_cache/cache[7][151] ), .QN(n3262) );
  DFFRX1 \D_cache/cache_reg[0][152]  ( .D(\D_cache/n580 ), .CK(clk), .RN(n5809), .Q(\D_cache/cache[0][152] ), .QN(n2416) );
  DFFRX1 \D_cache/cache_reg[1][152]  ( .D(\D_cache/n579 ), .CK(clk), .RN(n5809), .Q(\D_cache/cache[1][152] ), .QN(n1614) );
  DFFRX1 \D_cache/cache_reg[4][152]  ( .D(\D_cache/n576 ), .CK(clk), .RN(n5809), .Q(\D_cache/cache[4][152] ), .QN(n1617) );
  DFFRX1 \D_cache/cache_reg[5][152]  ( .D(\D_cache/n575 ), .CK(clk), .RN(n5809), .Q(\D_cache/cache[5][152] ), .QN(n224) );
  DFFRX1 \D_cache/cache_reg[0][153]  ( .D(\D_cache/n572 ), .CK(clk), .RN(n5810), .Q(\D_cache/cache[0][153] ), .QN(n3239) );
  DFFRX1 \D_cache/cache_reg[1][153]  ( .D(\D_cache/n571 ), .CK(clk), .RN(n5810), .Q(\D_cache/cache[1][153] ), .QN(n1610) );
  DFFRX1 \D_cache/cache_reg[2][153]  ( .D(\D_cache/n570 ), .CK(clk), .RN(n5810), .Q(\D_cache/cache[2][153] ), .QN(n2339) );
  DFFRX1 \D_cache/cache_reg[3][153]  ( .D(\D_cache/n569 ), .CK(clk), .RN(n5810), .Q(\D_cache/cache[3][153] ), .QN(n803) );
  DFFRX1 \D_cache/cache_reg[4][153]  ( .D(\D_cache/n568 ), .CK(clk), .RN(n5810), .Q(\D_cache/cache[4][153] ), .QN(n2337) );
  DFFRX1 \D_cache/cache_reg[5][153]  ( .D(\D_cache/n567 ), .CK(clk), .RN(n5810), .Q(\D_cache/cache[5][153] ), .QN(n801) );
  DFFRX1 \D_cache/cache_reg[6][153]  ( .D(\D_cache/n566 ), .CK(clk), .RN(n5810), .Q(\D_cache/cache[6][153] ), .QN(n1155) );
  DFFRX1 \D_cache/cache_reg[7][153]  ( .D(\D_cache/n565 ), .CK(clk), .RN(n5810), .Q(\D_cache/cache[7][153] ), .QN(n2727) );
  DFFRX1 \I_cache/cache_reg[0][0]  ( .D(n12822), .CK(clk), .RN(n5811), .Q(
        \I_cache/cache[0][0] ), .QN(n2520) );
  DFFRX1 \I_cache/cache_reg[1][0]  ( .D(n12821), .CK(clk), .RN(n5811), .Q(
        \I_cache/cache[1][0] ), .QN(n769) );
  DFFRX1 \I_cache/cache_reg[2][0]  ( .D(n12820), .CK(clk), .RN(n5811), .Q(
        \I_cache/cache[2][0] ), .QN(n2521) );
  DFFRX1 \I_cache/cache_reg[3][0]  ( .D(n12819), .CK(clk), .RN(n5811), .Q(
        \I_cache/cache[3][0] ), .QN(n770) );
  DFFRX1 \I_cache/cache_reg[4][0]  ( .D(n12818), .CK(clk), .RN(n5811), .Q(
        \I_cache/cache[4][0] ), .QN(n2570) );
  DFFRX1 \I_cache/cache_reg[5][0]  ( .D(n12817), .CK(clk), .RN(n5811), .Q(
        \I_cache/cache[5][0] ), .QN(n799) );
  DFFRX1 \I_cache/cache_reg[6][0]  ( .D(n12816), .CK(clk), .RN(n5811), .Q(
        \I_cache/cache[6][0] ), .QN(n743) );
  DFFRX1 \I_cache/cache_reg[7][0]  ( .D(n12823), .CK(clk), .RN(n5812), .Q(
        \I_cache/cache[7][0] ), .QN(n2324) );
  DFFRX1 \I_cache/cache_reg[0][1]  ( .D(n12815), .CK(clk), .RN(n5812), .Q(
        \I_cache/cache[0][1] ), .QN(n1147) );
  DFFRX1 \I_cache/cache_reg[1][1]  ( .D(n12814), .CK(clk), .RN(n5812), .Q(
        \I_cache/cache[1][1] ), .QN(n2719) );
  DFFRX1 \I_cache/cache_reg[2][1]  ( .D(n12813), .CK(clk), .RN(n5812), .Q(
        \I_cache/cache[2][1] ), .QN(n1148) );
  DFFRX1 \I_cache/cache_reg[3][1]  ( .D(n12812), .CK(clk), .RN(n5812), .Q(
        \I_cache/cache[3][1] ), .QN(n2720) );
  DFFRX1 \I_cache/cache_reg[4][1]  ( .D(n12811), .CK(clk), .RN(n5812), .Q(
        \I_cache/cache[4][1] ), .QN(n1221) );
  DFFRX1 \I_cache/cache_reg[5][1]  ( .D(n12810), .CK(clk), .RN(n5812), .Q(
        \I_cache/cache[5][1] ), .QN(n2793) );
  DFFRX1 \I_cache/cache_reg[6][1]  ( .D(n12809), .CK(clk), .RN(n5812), .Q(
        \I_cache/cache[6][1] ), .QN(n1146) );
  DFFRX1 \I_cache/cache_reg[7][1]  ( .D(n12808), .CK(clk), .RN(n5812), .Q(
        \I_cache/cache[7][1] ), .QN(n2718) );
  DFFRX1 \I_cache/cache_reg[0][2]  ( .D(n12807), .CK(clk), .RN(n5812), .Q(
        \I_cache/cache[0][2] ), .QN(n1127) );
  DFFRX1 \I_cache/cache_reg[1][2]  ( .D(n12806), .CK(clk), .RN(n5812), .Q(
        \I_cache/cache[1][2] ), .QN(n2699) );
  DFFRX1 \I_cache/cache_reg[2][2]  ( .D(n12805), .CK(clk), .RN(n5812), .Q(
        \I_cache/cache[2][2] ), .QN(n1128) );
  DFFRX1 \I_cache/cache_reg[3][2]  ( .D(n12804), .CK(clk), .RN(n5813), .Q(
        \I_cache/cache[3][2] ), .QN(n2700) );
  DFFRX1 \I_cache/cache_reg[4][2]  ( .D(n12803), .CK(clk), .RN(n5813), .Q(
        \I_cache/cache[4][2] ), .QN(n2568) );
  DFFRX1 \I_cache/cache_reg[5][2]  ( .D(n12802), .CK(clk), .RN(n5813), .Q(
        \I_cache/cache[5][2] ), .QN(n797) );
  DFFRX1 \I_cache/cache_reg[6][2]  ( .D(n12801), .CK(clk), .RN(n5813), .Q(
        \I_cache/cache[6][2] ), .QN(n1126) );
  DFFRX1 \I_cache/cache_reg[7][2]  ( .D(n12800), .CK(clk), .RN(n5813), .Q(
        \I_cache/cache[7][2] ), .QN(n2698) );
  DFFRX1 \I_cache/cache_reg[0][3]  ( .D(n12799), .CK(clk), .RN(n5813), .Q(
        \I_cache/cache[0][3] ), .QN(n741) );
  DFFRX1 \I_cache/cache_reg[1][3]  ( .D(n12798), .CK(clk), .RN(n5813), .Q(
        \I_cache/cache[1][3] ), .QN(n2322) );
  DFFRX1 \I_cache/cache_reg[2][3]  ( .D(n12797), .CK(clk), .RN(n5813), .Q(
        \I_cache/cache[2][3] ), .QN(n742) );
  DFFRX1 \I_cache/cache_reg[3][3]  ( .D(n12796), .CK(clk), .RN(n5813), .Q(
        \I_cache/cache[3][3] ), .QN(n2323) );
  DFFRX1 \I_cache/cache_reg[4][3]  ( .D(n12795), .CK(clk), .RN(n5813), .Q(
        \I_cache/cache[4][3] ), .QN(n746) );
  DFFRX1 \I_cache/cache_reg[5][3]  ( .D(n12794), .CK(clk), .RN(n5813), .Q(
        \I_cache/cache[5][3] ), .QN(n2325) );
  DFFRX1 \I_cache/cache_reg[6][3]  ( .D(n12793), .CK(clk), .RN(n5813), .Q(
        \I_cache/cache[6][3] ), .QN(n740) );
  DFFRX1 \I_cache/cache_reg[7][3]  ( .D(n12792), .CK(clk), .RN(n5814), .Q(
        \I_cache/cache[7][3] ), .QN(n2321) );
  DFFRX1 \I_cache/cache_reg[0][4]  ( .D(n12791), .CK(clk), .RN(n5814), .Q(
        \I_cache/cache[0][4] ), .QN(n1105) );
  DFFRX1 \I_cache/cache_reg[1][4]  ( .D(n12790), .CK(clk), .RN(n5814), .Q(
        \I_cache/cache[1][4] ), .QN(n2677) );
  DFFRX1 \I_cache/cache_reg[2][4]  ( .D(n12789), .CK(clk), .RN(n5814), .Q(
        \I_cache/cache[2][4] ), .QN(n1106) );
  DFFRX1 \I_cache/cache_reg[3][4]  ( .D(n12788), .CK(clk), .RN(n5814), .Q(
        \I_cache/cache[3][4] ), .QN(n2678) );
  DFFRX1 \I_cache/cache_reg[4][4]  ( .D(n12787), .CK(clk), .RN(n5814), .Q(
        \I_cache/cache[4][4] ), .QN(n753) );
  DFFRX1 \I_cache/cache_reg[5][4]  ( .D(n12786), .CK(clk), .RN(n5814), .Q(
        \I_cache/cache[5][4] ), .QN(n2331) );
  DFFRX1 \I_cache/cache_reg[6][4]  ( .D(n12785), .CK(clk), .RN(n5814), .Q(
        \I_cache/cache[6][4] ), .QN(n2554) );
  DFFRX1 \I_cache/cache_reg[7][4]  ( .D(n12784), .CK(clk), .RN(n5814), .Q(
        \I_cache/cache[7][4] ), .QN(n783) );
  DFFRX1 \I_cache/cache_reg[0][5]  ( .D(n12783), .CK(clk), .RN(n5814), .Q(
        \I_cache/cache[0][5] ), .QN(n438) );
  DFFRX1 \I_cache/cache_reg[1][5]  ( .D(n12782), .CK(clk), .RN(n5814), .Q(
        \I_cache/cache[1][5] ), .QN(n2001) );
  DFFRX1 \I_cache/cache_reg[2][5]  ( .D(n12781), .CK(clk), .RN(n5814), .Q(
        \I_cache/cache[2][5] ), .QN(n2421) );
  DFFRX1 \I_cache/cache_reg[3][5]  ( .D(n12780), .CK(clk), .RN(n5815), .Q(
        \I_cache/cache[3][5] ), .QN(n444) );
  DFFRX1 \I_cache/cache_reg[4][5]  ( .D(n12779), .CK(clk), .RN(n5815), .Q(
        \I_cache/cache[4][5] ), .QN(n2526) );
  DFFRX1 \I_cache/cache_reg[6][5]  ( .D(n12777), .CK(clk), .RN(n5815), .Q(
        \I_cache/cache[6][5] ), .QN(n2420) );
  DFFRX1 \I_cache/cache_reg[0][6]  ( .D(n12775), .CK(clk), .RN(n5815), .Q(
        \I_cache/cache[0][6] ), .QN(n1066) );
  DFFRX1 \I_cache/cache_reg[1][6]  ( .D(n12774), .CK(clk), .RN(n5815), .Q(
        \I_cache/cache[1][6] ), .QN(n2638) );
  DFFRX1 \I_cache/cache_reg[2][6]  ( .D(n12773), .CK(clk), .RN(n5815), .Q(
        \I_cache/cache[2][6] ), .QN(n1064) );
  DFFRX1 \I_cache/cache_reg[3][6]  ( .D(n12772), .CK(clk), .RN(n5815), .Q(
        \I_cache/cache[3][6] ), .QN(n2636) );
  DFFRX1 \I_cache/cache_reg[4][6]  ( .D(n12771), .CK(clk), .RN(n5815), .Q(
        \I_cache/cache[4][6] ), .QN(n2536) );
  DFFRX1 \I_cache/cache_reg[5][6]  ( .D(n12770), .CK(clk), .RN(n5815), .Q(
        \I_cache/cache[5][6] ), .QN(n777) );
  DFFRX1 \I_cache/cache_reg[6][6]  ( .D(n12769), .CK(clk), .RN(n5815), .Q(
        \I_cache/cache[6][6] ), .QN(n1065) );
  DFFRX1 \I_cache/cache_reg[7][6]  ( .D(n12768), .CK(clk), .RN(n5816), .Q(
        \I_cache/cache[7][6] ), .QN(n2637) );
  DFFRX1 \I_cache/cache_reg[0][7]  ( .D(n12767), .CK(clk), .RN(n5816), .Q(
        \I_cache/cache[0][7] ), .QN(n994) );
  DFFRX1 \I_cache/cache_reg[1][7]  ( .D(n12766), .CK(clk), .RN(n5816), .Q(
        \I_cache/cache[1][7] ), .QN(n2546) );
  DFFRX1 \I_cache/cache_reg[2][7]  ( .D(n12765), .CK(clk), .RN(n5816), .Q(
        \I_cache/cache[2][7] ), .QN(n995) );
  DFFRX1 \I_cache/cache_reg[3][7]  ( .D(n12764), .CK(clk), .RN(n5816), .Q(
        \I_cache/cache[3][7] ), .QN(n2547) );
  DFFRX1 \I_cache/cache_reg[4][7]  ( .D(n12763), .CK(clk), .RN(n5816), .Q(
        \I_cache/cache[4][7] ), .QN(n996) );
  DFFRX1 \I_cache/cache_reg[5][7]  ( .D(n12762), .CK(clk), .RN(n5816), .Q(
        \I_cache/cache[5][7] ), .QN(n2548) );
  DFFRX1 \I_cache/cache_reg[6][7]  ( .D(n12761), .CK(clk), .RN(n5816), .Q(
        \I_cache/cache[6][7] ), .QN(n993) );
  DFFRX1 \I_cache/cache_reg[7][7]  ( .D(n12760), .CK(clk), .RN(n5816), .Q(
        \I_cache/cache[7][7] ), .QN(n2545) );
  DFFRX1 \I_cache/cache_reg[0][8]  ( .D(n12759), .CK(clk), .RN(n5816), .Q(
        \I_cache/cache[0][8] ), .QN(n1107) );
  DFFRX1 \I_cache/cache_reg[1][8]  ( .D(n12758), .CK(clk), .RN(n5816), .Q(
        \I_cache/cache[1][8] ), .QN(n2679) );
  DFFRX1 \I_cache/cache_reg[2][8]  ( .D(n12757), .CK(clk), .RN(n5816), .Q(
        \I_cache/cache[2][8] ), .QN(n1108) );
  DFFRX1 \I_cache/cache_reg[3][8]  ( .D(n12756), .CK(clk), .RN(n5817), .Q(
        \I_cache/cache[3][8] ), .QN(n2680) );
  DFFRX1 \I_cache/cache_reg[4][8]  ( .D(n12755), .CK(clk), .RN(n5817), .Q(
        \I_cache/cache[4][8] ), .QN(n1191) );
  DFFRX1 \I_cache/cache_reg[5][8]  ( .D(n12754), .CK(clk), .RN(n5817), .Q(
        \I_cache/cache[5][8] ), .QN(n2763) );
  DFFRX1 \I_cache/cache_reg[6][8]  ( .D(n12753), .CK(clk), .RN(n5817), .Q(
        \I_cache/cache[6][8] ), .QN(n1109) );
  DFFRX1 \I_cache/cache_reg[7][8]  ( .D(n12752), .CK(clk), .RN(n5817), .Q(
        \I_cache/cache[7][8] ), .QN(n2681) );
  DFFRX1 \I_cache/cache_reg[0][9]  ( .D(n12751), .CK(clk), .RN(n5817), .Q(
        \I_cache/cache[0][9] ), .QN(n1061) );
  DFFRX1 \I_cache/cache_reg[1][9]  ( .D(n12750), .CK(clk), .RN(n5817), .Q(
        \I_cache/cache[1][9] ), .QN(n2633) );
  DFFRX1 \I_cache/cache_reg[2][9]  ( .D(n12749), .CK(clk), .RN(n5817), .Q(
        \I_cache/cache[2][9] ), .QN(n1060) );
  DFFRX1 \I_cache/cache_reg[3][9]  ( .D(n12748), .CK(clk), .RN(n5817), .Q(
        \I_cache/cache[3][9] ), .QN(n2632) );
  DFFRX1 \I_cache/cache_reg[6][9]  ( .D(n12745), .CK(clk), .RN(n5817), .Q(
        \I_cache/cache[6][9] ), .QN(n1067) );
  DFFRX1 \I_cache/cache_reg[7][9]  ( .D(n12744), .CK(clk), .RN(n5818), .Q(
        \I_cache/cache[7][9] ), .QN(n2639) );
  DFFRX1 \I_cache/cache_reg[0][10]  ( .D(n12743), .CK(clk), .RN(n5818), .Q(
        \I_cache/cache[0][10] ), .QN(n918) );
  DFFRX1 \I_cache/cache_reg[1][10]  ( .D(n12742), .CK(clk), .RN(n5818), .Q(
        \I_cache/cache[1][10] ), .QN(n2435) );
  DFFRX1 \I_cache/cache_reg[2][10]  ( .D(n12741), .CK(clk), .RN(n5818), .Q(
        \I_cache/cache[2][10] ), .QN(n919) );
  DFFRX1 \I_cache/cache_reg[3][10]  ( .D(n12740), .CK(clk), .RN(n5818), .Q(
        \I_cache/cache[3][10] ), .QN(n2436) );
  DFFRX1 \I_cache/cache_reg[6][10]  ( .D(n12737), .CK(clk), .RN(n5818), .Q(
        \I_cache/cache[6][10] ), .QN(n1002) );
  DFFRX1 \I_cache/cache_reg[7][10]  ( .D(n12736), .CK(clk), .RN(n5818), .Q(
        \I_cache/cache[7][10] ), .QN(n2574) );
  DFFRX1 \I_cache/cache_reg[0][11]  ( .D(n12735), .CK(clk), .RN(n5818), .Q(
        \I_cache/cache[0][11] ), .QN(n1000) );
  DFFRX1 \I_cache/cache_reg[1][11]  ( .D(n12734), .CK(clk), .RN(n5818), .Q(
        \I_cache/cache[1][11] ), .QN(n2572) );
  DFFRX1 \I_cache/cache_reg[2][11]  ( .D(n12733), .CK(clk), .RN(n5818), .Q(
        \I_cache/cache[2][11] ), .QN(n1001) );
  DFFRX1 \I_cache/cache_reg[3][11]  ( .D(n12732), .CK(clk), .RN(n5819), .Q(
        \I_cache/cache[3][11] ), .QN(n2573) );
  DFFRX1 \I_cache/cache_reg[4][11]  ( .D(n12731), .CK(clk), .RN(n5819), .Q(
        \I_cache/cache[4][11] ), .QN(n1205) );
  DFFRX1 \I_cache/cache_reg[5][11]  ( .D(n12730), .CK(clk), .RN(n5819), .Q(
        \I_cache/cache[5][11] ), .QN(n2777) );
  DFFRX1 \I_cache/cache_reg[6][11]  ( .D(n12729), .CK(clk), .RN(n5819), .Q(
        \I_cache/cache[6][11] ), .QN(n999) );
  DFFRX1 \I_cache/cache_reg[7][11]  ( .D(n12728), .CK(clk), .RN(n5819), .Q(
        \I_cache/cache[7][11] ), .QN(n2571) );
  DFFRX1 \I_cache/cache_reg[0][12]  ( .D(n12727), .CK(clk), .RN(n5819), .Q(
        \I_cache/cache[0][12] ), .QN(n1034) );
  DFFRX1 \I_cache/cache_reg[1][12]  ( .D(n12726), .CK(clk), .RN(n5819), .Q(
        \I_cache/cache[1][12] ), .QN(n2606) );
  DFFRX1 \I_cache/cache_reg[3][12]  ( .D(n12724), .CK(clk), .RN(n5819), .Q(
        \I_cache/cache[3][12] ), .QN(n2607) );
  DFFRX1 \I_cache/cache_reg[4][12]  ( .D(n12723), .CK(clk), .RN(n5819), .Q(
        \I_cache/cache[4][12] ), .QN(n1051) );
  DFFRX1 \I_cache/cache_reg[6][12]  ( .D(n12721), .CK(clk), .RN(n5819), .Q(
        \I_cache/cache[6][12] ), .QN(n1036) );
  DFFRX1 \I_cache/cache_reg[7][12]  ( .D(n12720), .CK(clk), .RN(n5820), .Q(
        \I_cache/cache[7][12] ), .QN(n2608) );
  DFFRX1 \I_cache/cache_reg[0][13]  ( .D(n12719), .CK(clk), .RN(n5820), .Q(
        \I_cache/cache[0][13] ), .QN(n911) );
  DFFRX1 \I_cache/cache_reg[1][13]  ( .D(n12718), .CK(clk), .RN(n5820), .Q(
        \I_cache/cache[1][13] ), .QN(n2428) );
  DFFRX1 \I_cache/cache_reg[2][13]  ( .D(n12717), .CK(clk), .RN(n5820), .Q(
        \I_cache/cache[2][13] ), .QN(n912) );
  DFFRX1 \I_cache/cache_reg[3][13]  ( .D(n12716), .CK(clk), .RN(n5820), .Q(
        \I_cache/cache[3][13] ), .QN(n2429) );
  DFFRX1 \I_cache/cache_reg[4][13]  ( .D(n12715), .CK(clk), .RN(n5820), .Q(
        \I_cache/cache[4][13] ), .QN(n755) );
  DFFRX1 \I_cache/cache_reg[5][13]  ( .D(n12714), .CK(clk), .RN(n5820), .Q(
        \I_cache/cache[5][13] ), .QN(n2333) );
  DFFRX1 \I_cache/cache_reg[6][13]  ( .D(n12713), .CK(clk), .RN(n5820), .Q(
        \I_cache/cache[6][13] ), .QN(n908) );
  DFFRX1 \I_cache/cache_reg[7][13]  ( .D(n12712), .CK(clk), .RN(n5820), .Q(
        \I_cache/cache[7][13] ), .QN(n2425) );
  DFFRX1 \I_cache/cache_reg[0][14]  ( .D(n12711), .CK(clk), .RN(n5820), .Q(
        \I_cache/cache[0][14] ), .QN(n1023) );
  DFFRX1 \I_cache/cache_reg[1][14]  ( .D(n12710), .CK(clk), .RN(n5820), .Q(
        \I_cache/cache[1][14] ), .QN(n2595) );
  DFFRX1 \I_cache/cache_reg[2][14]  ( .D(n12709), .CK(clk), .RN(n5820), .Q(
        \I_cache/cache[2][14] ), .QN(n1024) );
  DFFRX1 \I_cache/cache_reg[3][14]  ( .D(n12708), .CK(clk), .RN(n5821), .Q(
        \I_cache/cache[3][14] ), .QN(n2596) );
  DFFRX1 \I_cache/cache_reg[4][14]  ( .D(n12707), .CK(clk), .RN(n5821), .Q(
        \I_cache/cache[4][14] ), .QN(n1202) );
  DFFRX1 \I_cache/cache_reg[5][14]  ( .D(n12706), .CK(clk), .RN(n5821), .Q(
        \I_cache/cache[5][14] ), .QN(n2774) );
  DFFRX1 \I_cache/cache_reg[6][14]  ( .D(n12705), .CK(clk), .RN(n5821), .Q(
        \I_cache/cache[6][14] ), .QN(n1025) );
  DFFRX1 \I_cache/cache_reg[7][14]  ( .D(n12704), .CK(clk), .RN(n5821), .Q(
        \I_cache/cache[7][14] ), .QN(n2597) );
  DFFRX1 \I_cache/cache_reg[0][15]  ( .D(n12703), .CK(clk), .RN(n5821), .Q(
        \I_cache/cache[0][15] ), .QN(n1238) );
  DFFRX1 \I_cache/cache_reg[1][15]  ( .D(n12702), .CK(clk), .RN(n5821), .Q(
        \I_cache/cache[1][15] ), .QN(n2843) );
  DFFRX1 \I_cache/cache_reg[2][15]  ( .D(n12701), .CK(clk), .RN(n5821), .Q(
        \I_cache/cache[2][15] ), .QN(n1496) );
  DFFRX1 \I_cache/cache_reg[3][15]  ( .D(n12700), .CK(clk), .RN(n5821), .Q(
        \I_cache/cache[3][15] ), .QN(n3109) );
  DFFRX1 \I_cache/cache_reg[4][15]  ( .D(n12699), .CK(clk), .RN(n5821), .Q(
        \I_cache/cache[4][15] ), .QN(n1580) );
  DFFRX1 \I_cache/cache_reg[5][15]  ( .D(n12698), .CK(clk), .RN(n5821), .Q(
        \I_cache/cache[5][15] ), .QN(n3193) );
  DFFRX1 \I_cache/cache_reg[6][15]  ( .D(n12697), .CK(clk), .RN(n5821), .Q(
        \I_cache/cache[6][15] ), .QN(n1495) );
  DFFRX1 \I_cache/cache_reg[7][15]  ( .D(n12696), .CK(clk), .RN(n5822), .Q(
        \I_cache/cache[7][15] ), .QN(n3108) );
  DFFRX1 \I_cache/cache_reg[0][32]  ( .D(n12567), .CK(clk), .RN(n5832), .Q(
        \I_cache/cache[0][32] ), .QN(n2523) );
  DFFRX1 \I_cache/cache_reg[1][32]  ( .D(n12566), .CK(clk), .RN(n5832), .Q(
        \I_cache/cache[1][32] ), .QN(n772) );
  DFFRX1 \I_cache/cache_reg[2][32]  ( .D(n12565), .CK(clk), .RN(n5832), .Q(
        \I_cache/cache[2][32] ), .QN(n2524) );
  DFFRX1 \I_cache/cache_reg[3][32]  ( .D(n12564), .CK(clk), .RN(n5833), .Q(
        \I_cache/cache[3][32] ), .QN(n773) );
  DFFRX1 \I_cache/cache_reg[4][32]  ( .D(n12563), .CK(clk), .RN(n5833), .Q(
        \I_cache/cache[4][32] ), .QN(n1199) );
  DFFRX1 \I_cache/cache_reg[5][32]  ( .D(n12562), .CK(clk), .RN(n5833), .Q(
        \I_cache/cache[5][32] ), .QN(n2771) );
  DFFRX1 \I_cache/cache_reg[6][32]  ( .D(n12561), .CK(clk), .RN(n5833), .Q(
        \I_cache/cache[6][32] ), .QN(n2522) );
  DFFRX1 \I_cache/cache_reg[7][32]  ( .D(n12560), .CK(clk), .RN(n5833), .Q(
        \I_cache/cache[7][32] ), .QN(n771) );
  DFFRX1 \I_cache/cache_reg[0][33]  ( .D(n12559), .CK(clk), .RN(n5833), .Q(
        \I_cache/cache[0][33] ), .QN(n1072) );
  DFFRX1 \I_cache/cache_reg[1][33]  ( .D(n12558), .CK(clk), .RN(n5833), .Q(
        \I_cache/cache[1][33] ), .QN(n2644) );
  DFFRX1 \I_cache/cache_reg[2][33]  ( .D(n12557), .CK(clk), .RN(n5833), .Q(
        \I_cache/cache[2][33] ), .QN(n1071) );
  DFFRX1 \I_cache/cache_reg[3][33]  ( .D(n12556), .CK(clk), .RN(n5833), .Q(
        \I_cache/cache[3][33] ), .QN(n2643) );
  DFFRX1 \I_cache/cache_reg[4][33]  ( .D(n12555), .CK(clk), .RN(n5833), .Q(
        \I_cache/cache[4][33] ), .QN(n2538) );
  DFFRX1 \I_cache/cache_reg[5][33]  ( .D(n12554), .CK(clk), .RN(n5833), .Q(
        \I_cache/cache[5][33] ), .QN(n779) );
  DFFRX1 \I_cache/cache_reg[6][33]  ( .D(n12553), .CK(clk), .RN(n5833), .Q(
        \I_cache/cache[6][33] ), .QN(n2532) );
  DFFRX1 \I_cache/cache_reg[7][33]  ( .D(n12552), .CK(clk), .RN(n5834), .Q(
        \I_cache/cache[7][33] ), .QN(n776) );
  DFFRX1 \I_cache/cache_reg[0][34]  ( .D(n12551), .CK(clk), .RN(n5834), .Q(
        \I_cache/cache[0][34] ), .QN(n1124) );
  DFFRX1 \I_cache/cache_reg[1][34]  ( .D(n12550), .CK(clk), .RN(n5834), .Q(
        \I_cache/cache[1][34] ), .QN(n2696) );
  DFFRX1 \I_cache/cache_reg[2][34]  ( .D(n12549), .CK(clk), .RN(n5834), .Q(
        \I_cache/cache[2][34] ), .QN(n1125) );
  DFFRX1 \I_cache/cache_reg[3][34]  ( .D(n12548), .CK(clk), .RN(n5834), .Q(
        \I_cache/cache[3][34] ), .QN(n2697) );
  DFFRX1 \I_cache/cache_reg[4][34]  ( .D(n12547), .CK(clk), .RN(n5834), .Q(
        \I_cache/cache[4][34] ), .QN(n2567) );
  DFFRX1 \I_cache/cache_reg[5][34]  ( .D(n12546), .CK(clk), .RN(n5834), .Q(
        \I_cache/cache[5][34] ), .QN(n796) );
  DFFRX1 \I_cache/cache_reg[6][34]  ( .D(n12545), .CK(clk), .RN(n5834), .Q(
        \I_cache/cache[6][34] ), .QN(n1123) );
  DFFRX1 \I_cache/cache_reg[7][34]  ( .D(n12544), .CK(clk), .RN(n5834), .Q(
        \I_cache/cache[7][34] ), .QN(n2695) );
  DFFRX1 \I_cache/cache_reg[0][35]  ( .D(n12543), .CK(clk), .RN(n5834), .Q(
        \I_cache/cache[0][35] ), .QN(n2517) );
  DFFRX1 \I_cache/cache_reg[1][35]  ( .D(n12542), .CK(clk), .RN(n5834), .Q(
        \I_cache/cache[1][35] ), .QN(n766) );
  DFFRX1 \I_cache/cache_reg[2][35]  ( .D(n12541), .CK(clk), .RN(n5834), .Q(
        \I_cache/cache[2][35] ), .QN(n2518) );
  DFFRX1 \I_cache/cache_reg[3][35]  ( .D(n12540), .CK(clk), .RN(n5835), .Q(
        \I_cache/cache[3][35] ), .QN(n767) );
  DFFRX1 \I_cache/cache_reg[4][35]  ( .D(n12539), .CK(clk), .RN(n5835), .Q(
        \I_cache/cache[4][35] ), .QN(n1194) );
  DFFRX1 \I_cache/cache_reg[5][35]  ( .D(n12538), .CK(clk), .RN(n5835), .Q(
        \I_cache/cache[5][35] ), .QN(n2766) );
  DFFRX1 \I_cache/cache_reg[6][35]  ( .D(n12537), .CK(clk), .RN(n5835), .Q(
        \I_cache/cache[6][35] ), .QN(n2516) );
  DFFRX1 \I_cache/cache_reg[7][35]  ( .D(n12536), .CK(clk), .RN(n5835), .Q(
        \I_cache/cache[7][35] ), .QN(n765) );
  DFFRX1 \I_cache/cache_reg[0][36]  ( .D(n12535), .CK(clk), .RN(n5835), .Q(
        \I_cache/cache[0][36] ), .QN(n1101) );
  DFFRX1 \I_cache/cache_reg[1][36]  ( .D(n12534), .CK(clk), .RN(n5835), .Q(
        \I_cache/cache[1][36] ), .QN(n2673) );
  DFFRX1 \I_cache/cache_reg[2][36]  ( .D(n12533), .CK(clk), .RN(n5835), .Q(
        \I_cache/cache[2][36] ), .QN(n2553) );
  DFFRX1 \I_cache/cache_reg[3][36]  ( .D(n12532), .CK(clk), .RN(n5835), .Q(
        \I_cache/cache[3][36] ), .QN(n782) );
  DFFRX1 \I_cache/cache_reg[4][36]  ( .D(n12531), .CK(clk), .RN(n5835), .Q(
        \I_cache/cache[4][36] ), .QN(n751) );
  DFFRX1 \I_cache/cache_reg[5][36]  ( .D(n12530), .CK(clk), .RN(n5835), .Q(
        \I_cache/cache[5][36] ), .QN(n2329) );
  DFFRX1 \I_cache/cache_reg[6][36]  ( .D(n12529), .CK(clk), .RN(n5835), .Q(
        \I_cache/cache[6][36] ), .QN(n2552) );
  DFFRX1 \I_cache/cache_reg[7][36]  ( .D(n12528), .CK(clk), .RN(n5836), .Q(
        \I_cache/cache[7][36] ), .QN(n781) );
  DFFRX1 \I_cache/cache_reg[0][37]  ( .D(n12527), .CK(clk), .RN(n5836), .Q(
        \I_cache/cache[0][37] ), .QN(n1136) );
  DFFRX1 \I_cache/cache_reg[1][37]  ( .D(n12526), .CK(clk), .RN(n5836), .Q(
        \I_cache/cache[1][37] ), .QN(n2708) );
  DFFRX1 \I_cache/cache_reg[2][37]  ( .D(n12525), .CK(clk), .RN(n5836), .Q(
        \I_cache/cache[2][37] ), .QN(n1137) );
  DFFRX1 \I_cache/cache_reg[3][37]  ( .D(n12524), .CK(clk), .RN(n5836), .Q(
        \I_cache/cache[3][37] ), .QN(n2709) );
  DFFRX1 \I_cache/cache_reg[4][37]  ( .D(n12523), .CK(clk), .RN(n5836), .Q(
        \I_cache/cache[4][37] ), .QN(n757) );
  DFFRX1 \I_cache/cache_reg[5][37]  ( .D(n12522), .CK(clk), .RN(n5836), .Q(
        \I_cache/cache[5][37] ), .QN(n2335) );
  DFFRX1 \I_cache/cache_reg[6][37]  ( .D(n12521), .CK(clk), .RN(n5836), .Q(
        \I_cache/cache[6][37] ), .QN(n1135) );
  DFFRX1 \I_cache/cache_reg[7][37]  ( .D(n12520), .CK(clk), .RN(n5836), .Q(
        \I_cache/cache[7][37] ), .QN(n2707) );
  DFFRX1 \I_cache/cache_reg[0][38]  ( .D(n12519), .CK(clk), .RN(n5836), .Q(
        \I_cache/cache[0][38] ), .QN(n1099) );
  DFFRX1 \I_cache/cache_reg[1][38]  ( .D(n12518), .CK(clk), .RN(n5836), .Q(
        \I_cache/cache[1][38] ), .QN(n2671) );
  DFFRX1 \I_cache/cache_reg[2][38]  ( .D(n12517), .CK(clk), .RN(n5836), .Q(
        \I_cache/cache[2][38] ), .QN(n1100) );
  DFFRX1 \I_cache/cache_reg[3][38]  ( .D(n12516), .CK(clk), .RN(n5837), .Q(
        \I_cache/cache[3][38] ), .QN(n2672) );
  DFFRX1 \I_cache/cache_reg[4][38]  ( .D(n12515), .CK(clk), .RN(n5837), .Q(
        \I_cache/cache[4][38] ), .QN(n1188) );
  DFFRX1 \I_cache/cache_reg[5][38]  ( .D(n12514), .CK(clk), .RN(n5837), .Q(
        \I_cache/cache[5][38] ), .QN(n2760) );
  DFFRX1 \I_cache/cache_reg[6][38]  ( .D(n12513), .CK(clk), .RN(n5837), .Q(
        \I_cache/cache[6][38] ), .QN(n1098) );
  DFFRX1 \I_cache/cache_reg[7][38]  ( .D(n12512), .CK(clk), .RN(n5837), .Q(
        \I_cache/cache[7][38] ), .QN(n2670) );
  DFFRX1 \I_cache/cache_reg[0][39]  ( .D(n12511), .CK(clk), .RN(n5837), .Q(
        \I_cache/cache[0][39] ), .QN(n1118) );
  DFFRX1 \I_cache/cache_reg[1][39]  ( .D(n12510), .CK(clk), .RN(n5837), .Q(
        \I_cache/cache[1][39] ), .QN(n2690) );
  DFFRX1 \I_cache/cache_reg[2][39]  ( .D(n12509), .CK(clk), .RN(n5837), .Q(
        \I_cache/cache[2][39] ), .QN(n1119) );
  DFFRX1 \I_cache/cache_reg[3][39]  ( .D(n12508), .CK(clk), .RN(n5837), .Q(
        \I_cache/cache[3][39] ), .QN(n2691) );
  DFFRX1 \I_cache/cache_reg[4][39]  ( .D(n12507), .CK(clk), .RN(n5837), .Q(
        \I_cache/cache[4][39] ), .QN(n1189) );
  DFFRX1 \I_cache/cache_reg[5][39]  ( .D(n12506), .CK(clk), .RN(n5837), .Q(
        \I_cache/cache[5][39] ), .QN(n2761) );
  DFFRX1 \I_cache/cache_reg[6][39]  ( .D(n12505), .CK(clk), .RN(n5837), .Q(
        \I_cache/cache[6][39] ), .QN(n1117) );
  DFFRX1 \I_cache/cache_reg[7][39]  ( .D(n12504), .CK(clk), .RN(n5838), .Q(
        \I_cache/cache[7][39] ), .QN(n2689) );
  DFFRX1 \I_cache/cache_reg[0][40]  ( .D(n12503), .CK(clk), .RN(n5838), .Q(
        \I_cache/cache[0][40] ), .QN(n1110) );
  DFFRX1 \I_cache/cache_reg[1][40]  ( .D(n12502), .CK(clk), .RN(n5838), .Q(
        \I_cache/cache[1][40] ), .QN(n2682) );
  DFFRX1 \I_cache/cache_reg[2][40]  ( .D(n12501), .CK(clk), .RN(n5838), .Q(
        \I_cache/cache[2][40] ), .QN(n1111) );
  DFFRX1 \I_cache/cache_reg[3][40]  ( .D(n12500), .CK(clk), .RN(n5838), .Q(
        \I_cache/cache[3][40] ), .QN(n2683) );
  DFFRX1 \I_cache/cache_reg[4][40]  ( .D(n12499), .CK(clk), .RN(n5838), .Q(
        \I_cache/cache[4][40] ), .QN(n1193) );
  DFFRX1 \I_cache/cache_reg[5][40]  ( .D(n12498), .CK(clk), .RN(n5838), .Q(
        \I_cache/cache[5][40] ), .QN(n2765) );
  DFFRX1 \I_cache/cache_reg[6][40]  ( .D(n12497), .CK(clk), .RN(n5838), .Q(
        \I_cache/cache[6][40] ), .QN(n1112) );
  DFFRX1 \I_cache/cache_reg[7][40]  ( .D(n12496), .CK(clk), .RN(n5838), .Q(
        \I_cache/cache[7][40] ), .QN(n2684) );
  DFFRX1 \I_cache/cache_reg[0][41]  ( .D(n12495), .CK(clk), .RN(n5838), .Q(
        \I_cache/cache[0][41] ), .QN(n1090) );
  DFFRX1 \I_cache/cache_reg[1][41]  ( .D(n12494), .CK(clk), .RN(n5838), .Q(
        \I_cache/cache[1][41] ), .QN(n2662) );
  DFFRX1 \I_cache/cache_reg[2][41]  ( .D(n12493), .CK(clk), .RN(n5838), .Q(
        \I_cache/cache[2][41] ), .QN(n1091) );
  DFFRX1 \I_cache/cache_reg[3][41]  ( .D(n12492), .CK(clk), .RN(n5839), .Q(
        \I_cache/cache[3][41] ), .QN(n2663) );
  DFFRX1 \I_cache/cache_reg[4][41]  ( .D(n12491), .CK(clk), .RN(n5839), .Q(
        \I_cache/cache[4][41] ), .QN(n750) );
  DFFRX1 \I_cache/cache_reg[5][41]  ( .D(n12490), .CK(clk), .RN(n5839), .Q(
        \I_cache/cache[5][41] ), .QN(n2328) );
  DFFRX1 \I_cache/cache_reg[6][41]  ( .D(n12489), .CK(clk), .RN(n5839), .Q(
        \I_cache/cache[6][41] ), .QN(n2803) );
  DFFRX1 \I_cache/cache_reg[7][41]  ( .D(n12488), .CK(clk), .RN(n5839), .Q(
        \I_cache/cache[7][41] ), .QN(n1223) );
  DFFRX1 \I_cache/cache_reg[0][42]  ( .D(n12487), .CK(clk), .RN(n5839), .Q(
        \I_cache/cache[0][42] ), .QN(n1130) );
  DFFRX1 \I_cache/cache_reg[1][42]  ( .D(n12486), .CK(clk), .RN(n5839), .Q(
        \I_cache/cache[1][42] ), .QN(n2702) );
  DFFRX1 \I_cache/cache_reg[2][42]  ( .D(n12485), .CK(clk), .RN(n5839), .Q(
        \I_cache/cache[2][42] ), .QN(n1131) );
  DFFRX1 \I_cache/cache_reg[3][42]  ( .D(n12484), .CK(clk), .RN(n5839), .Q(
        \I_cache/cache[3][42] ), .QN(n2703) );
  DFFRX1 \I_cache/cache_reg[4][42]  ( .D(n12483), .CK(clk), .RN(n5839), .Q(
        \I_cache/cache[4][42] ), .QN(n1195) );
  DFFRX1 \I_cache/cache_reg[5][42]  ( .D(n12482), .CK(clk), .RN(n5839), .Q(
        \I_cache/cache[5][42] ), .QN(n2767) );
  DFFRX1 \I_cache/cache_reg[6][42]  ( .D(n12481), .CK(clk), .RN(n5839), .Q(
        \I_cache/cache[6][42] ), .QN(n1129) );
  DFFRX1 \I_cache/cache_reg[7][42]  ( .D(n12480), .CK(clk), .RN(n5840), .Q(
        \I_cache/cache[7][42] ), .QN(n2701) );
  DFFRX1 \I_cache/cache_reg[0][43]  ( .D(n12479), .CK(clk), .RN(n5840), .Q(
        \I_cache/cache[0][43] ), .QN(n1153) );
  DFFRX1 \I_cache/cache_reg[1][43]  ( .D(n12478), .CK(clk), .RN(n5840), .Q(
        \I_cache/cache[1][43] ), .QN(n2725) );
  DFFRX1 \I_cache/cache_reg[2][43]  ( .D(n12477), .CK(clk), .RN(n5840), .Q(
        \I_cache/cache[2][43] ), .QN(n1154) );
  DFFRX1 \I_cache/cache_reg[3][43]  ( .D(n12476), .CK(clk), .RN(n5840), .Q(
        \I_cache/cache[3][43] ), .QN(n2726) );
  DFFRX1 \I_cache/cache_reg[4][43]  ( .D(n12475), .CK(clk), .RN(n5840), .Q(
        \I_cache/cache[4][43] ), .QN(n1197) );
  DFFRX1 \I_cache/cache_reg[5][43]  ( .D(n12474), .CK(clk), .RN(n5840), .Q(
        \I_cache/cache[5][43] ), .QN(n2769) );
  DFFRX1 \I_cache/cache_reg[6][43]  ( .D(n12473), .CK(clk), .RN(n5840), .Q(
        \I_cache/cache[6][43] ), .QN(n1152) );
  DFFRX1 \I_cache/cache_reg[7][43]  ( .D(n12472), .CK(clk), .RN(n5840), .Q(
        \I_cache/cache[7][43] ), .QN(n2724) );
  DFFRX1 \I_cache/cache_reg[0][44]  ( .D(n12471), .CK(clk), .RN(n5840), .Q(
        \I_cache/cache[0][44] ), .QN(n1039) );
  DFFRX1 \I_cache/cache_reg[1][44]  ( .D(n12470), .CK(clk), .RN(n5840), .Q(
        \I_cache/cache[1][44] ), .QN(n2611) );
  DFFRX1 \I_cache/cache_reg[2][44]  ( .D(n12469), .CK(clk), .RN(n5840), .Q(
        \I_cache/cache[2][44] ), .QN(n1040) );
  DFFRX1 \I_cache/cache_reg[3][44]  ( .D(n12468), .CK(clk), .RN(n5841), .Q(
        \I_cache/cache[3][44] ), .QN(n2612) );
  DFFRX1 \I_cache/cache_reg[4][44]  ( .D(n12467), .CK(clk), .RN(n5841), .Q(
        \I_cache/cache[4][44] ), .QN(n1204) );
  DFFRX1 \I_cache/cache_reg[6][44]  ( .D(n12465), .CK(clk), .RN(n5841), .Q(
        \I_cache/cache[6][44] ), .QN(n1041) );
  DFFRX1 \I_cache/cache_reg[0][45]  ( .D(n12463), .CK(clk), .RN(n5841), .Q(
        \I_cache/cache[0][45] ), .QN(n1093) );
  DFFRX1 \I_cache/cache_reg[1][45]  ( .D(n12462), .CK(clk), .RN(n5841), .Q(
        \I_cache/cache[1][45] ), .QN(n2665) );
  DFFRX1 \I_cache/cache_reg[2][45]  ( .D(n12461), .CK(clk), .RN(n5841), .Q(
        \I_cache/cache[2][45] ), .QN(n1094) );
  DFFRX1 \I_cache/cache_reg[3][45]  ( .D(n12460), .CK(clk), .RN(n5841), .Q(
        \I_cache/cache[3][45] ), .QN(n2666) );
  DFFRX1 \I_cache/cache_reg[4][45]  ( .D(n12459), .CK(clk), .RN(n5841), .Q(
        \I_cache/cache[4][45] ), .QN(n754) );
  DFFRX1 \I_cache/cache_reg[5][45]  ( .D(n12458), .CK(clk), .RN(n5841), .Q(
        \I_cache/cache[5][45] ), .QN(n2332) );
  DFFRX1 \I_cache/cache_reg[6][45]  ( .D(n12457), .CK(clk), .RN(n5841), .Q(
        \I_cache/cache[6][45] ), .QN(n1095) );
  DFFRX1 \I_cache/cache_reg[7][45]  ( .D(n12456), .CK(clk), .RN(n5842), .Q(
        \I_cache/cache[7][45] ), .QN(n2667) );
  DFFRX1 \I_cache/cache_reg[0][46]  ( .D(n12455), .CK(clk), .RN(n5842), .Q(
        \I_cache/cache[0][46] ), .QN(n1029) );
  DFFRX1 \I_cache/cache_reg[1][46]  ( .D(n12454), .CK(clk), .RN(n5842), .Q(
        \I_cache/cache[1][46] ), .QN(n2601) );
  DFFRX1 \I_cache/cache_reg[2][46]  ( .D(n12453), .CK(clk), .RN(n5842), .Q(
        \I_cache/cache[2][46] ), .QN(n1030) );
  DFFRX1 \I_cache/cache_reg[3][46]  ( .D(n12452), .CK(clk), .RN(n5842), .Q(
        \I_cache/cache[3][46] ), .QN(n2602) );
  DFFRX1 \I_cache/cache_reg[4][46]  ( .D(n12451), .CK(clk), .RN(n5842), .Q(
        \I_cache/cache[4][46] ), .QN(n1201) );
  DFFRX1 \I_cache/cache_reg[5][46]  ( .D(n12450), .CK(clk), .RN(n5842), .Q(
        \I_cache/cache[5][46] ), .QN(n2773) );
  DFFRX1 \I_cache/cache_reg[6][46]  ( .D(n12449), .CK(clk), .RN(n5842), .Q(
        \I_cache/cache[6][46] ), .QN(n1031) );
  DFFRX1 \I_cache/cache_reg[7][46]  ( .D(n12448), .CK(clk), .RN(n5842), .Q(
        \I_cache/cache[7][46] ), .QN(n2603) );
  DFFRX1 \I_cache/cache_reg[0][47]  ( .D(n12447), .CK(clk), .RN(n5842), .Q(
        \I_cache/cache[0][47] ), .QN(n1473) );
  DFFRX1 \I_cache/cache_reg[1][47]  ( .D(n12446), .CK(clk), .RN(n5842), .Q(
        \I_cache/cache[1][47] ), .QN(n3086) );
  DFFRX1 \I_cache/cache_reg[2][47]  ( .D(n12445), .CK(clk), .RN(n5842), .Q(
        \I_cache/cache[2][47] ), .QN(n1232) );
  DFFRX1 \I_cache/cache_reg[3][47]  ( .D(n12444), .CK(clk), .RN(n5843), .Q(
        \I_cache/cache[3][47] ), .QN(n2837) );
  DFFRX1 \I_cache/cache_reg[4][47]  ( .D(n12443), .CK(clk), .RN(n5843), .Q(
        \I_cache/cache[4][47] ), .QN(n1474) );
  DFFRX1 \I_cache/cache_reg[5][47]  ( .D(n12442), .CK(clk), .RN(n5843), .Q(
        \I_cache/cache[5][47] ), .QN(n3087) );
  DFFRX1 \I_cache/cache_reg[6][47]  ( .D(n12441), .CK(clk), .RN(n5843), .Q(
        \I_cache/cache[6][47] ), .QN(n2854) );
  DFFRX1 \I_cache/cache_reg[7][47]  ( .D(n12440), .CK(clk), .RN(n5843), .Q(
        \I_cache/cache[7][47] ), .QN(n847) );
  DFFRX1 \I_cache/cache_reg[0][65]  ( .D(n12303), .CK(clk), .RN(n5854), .Q(
        \I_cache/cache[0][65] ), .QN(n1138) );
  DFFRX1 \I_cache/cache_reg[1][65]  ( .D(n12302), .CK(clk), .RN(n5854), .Q(
        \I_cache/cache[1][65] ), .QN(n2710) );
  DFFRX1 \I_cache/cache_reg[2][65]  ( .D(n12301), .CK(clk), .RN(n5854), .Q(
        \I_cache/cache[2][65] ), .QN(n1139) );
  DFFRX1 \I_cache/cache_reg[3][65]  ( .D(n12300), .CK(clk), .RN(n5855), .Q(
        \I_cache/cache[3][65] ), .QN(n2711) );
  DFFRX1 \I_cache/cache_reg[4][65]  ( .D(n12299), .CK(clk), .RN(n5855), .Q(
        \I_cache/cache[4][65] ), .QN(n2569) );
  DFFRX1 \I_cache/cache_reg[5][65]  ( .D(n12298), .CK(clk), .RN(n5855), .Q(
        \I_cache/cache[5][65] ), .QN(n798) );
  DFFRX1 \I_cache/cache_reg[6][65]  ( .D(n12297), .CK(clk), .RN(n5855), .Q(
        \I_cache/cache[6][65] ), .QN(n2557) );
  DFFRX1 \I_cache/cache_reg[7][65]  ( .D(n12296), .CK(clk), .RN(n5855), .Q(
        \I_cache/cache[7][65] ), .QN(n786) );
  DFFRX1 \I_cache/cache_reg[0][66]  ( .D(n12295), .CK(clk), .RN(n5855), .Q(
        \I_cache/cache[0][66] ), .QN(n1121) );
  DFFRX1 \I_cache/cache_reg[1][66]  ( .D(n12294), .CK(clk), .RN(n5855), .Q(
        \I_cache/cache[1][66] ), .QN(n2693) );
  DFFRX1 \I_cache/cache_reg[2][66]  ( .D(n12293), .CK(clk), .RN(n5855), .Q(
        \I_cache/cache[2][66] ), .QN(n1122) );
  DFFRX1 \I_cache/cache_reg[3][66]  ( .D(n12292), .CK(clk), .RN(n5855), .Q(
        \I_cache/cache[3][66] ), .QN(n2694) );
  DFFRX1 \I_cache/cache_reg[4][66]  ( .D(n12291), .CK(clk), .RN(n5855), .Q(
        \I_cache/cache[4][66] ), .QN(n2566) );
  DFFRX1 \I_cache/cache_reg[5][66]  ( .D(n12290), .CK(clk), .RN(n5855), .Q(
        \I_cache/cache[5][66] ), .QN(n795) );
  DFFRX1 \I_cache/cache_reg[6][66]  ( .D(n12289), .CK(clk), .RN(n5855), .Q(
        \I_cache/cache[6][66] ), .QN(n1120) );
  DFFRX1 \I_cache/cache_reg[7][66]  ( .D(n12288), .CK(clk), .RN(n5856), .Q(
        \I_cache/cache[7][66] ), .QN(n2692) );
  DFFRX1 \I_cache/cache_reg[0][67]  ( .D(n12287), .CK(clk), .RN(n5856), .Q(
        \I_cache/cache[0][67] ), .QN(n1150) );
  DFFRX1 \I_cache/cache_reg[1][67]  ( .D(n12286), .CK(clk), .RN(n5856), .Q(
        \I_cache/cache[1][67] ), .QN(n2722) );
  DFFRX1 \I_cache/cache_reg[2][67]  ( .D(n12285), .CK(clk), .RN(n5856), .Q(
        \I_cache/cache[2][67] ), .QN(n1151) );
  DFFRX1 \I_cache/cache_reg[3][67]  ( .D(n12284), .CK(clk), .RN(n5856), .Q(
        \I_cache/cache[3][67] ), .QN(n2723) );
  DFFRX1 \I_cache/cache_reg[4][67]  ( .D(n12283), .CK(clk), .RN(n5856), .Q(
        \I_cache/cache[4][67] ), .QN(n1083) );
  DFFRX1 \I_cache/cache_reg[5][67]  ( .D(n12282), .CK(clk), .RN(n5856), .Q(
        \I_cache/cache[5][67] ), .QN(n2655) );
  DFFRX1 \I_cache/cache_reg[6][67]  ( .D(n12281), .CK(clk), .RN(n5856), .Q(
        \I_cache/cache[6][67] ), .QN(n1149) );
  DFFRX1 \I_cache/cache_reg[7][67]  ( .D(n12280), .CK(clk), .RN(n5856), .Q(
        \I_cache/cache[7][67] ), .QN(n2721) );
  DFFRX1 \I_cache/cache_reg[0][68]  ( .D(n12279), .CK(clk), .RN(n5856), .Q(
        \I_cache/cache[0][68] ), .QN(n714) );
  DFFRX1 \I_cache/cache_reg[1][68]  ( .D(n12278), .CK(clk), .RN(n5856), .Q(
        \I_cache/cache[1][68] ), .QN(n2314) );
  DFFRX1 \I_cache/cache_reg[2][68]  ( .D(n12277), .CK(clk), .RN(n5856), .Q(
        \I_cache/cache[2][68] ), .QN(n442) );
  DFFRX1 \I_cache/cache_reg[3][68]  ( .D(n12276), .CK(clk), .RN(n5857), .Q(
        \I_cache/cache[3][68] ), .QN(n2004) );
  DFFRX1 \I_cache/cache_reg[4][68]  ( .D(n12275), .CK(clk), .RN(n5857), .Q(
        \I_cache/cache[4][68] ), .QN(n2551) );
  DFFRX1 \I_cache/cache_reg[5][68]  ( .D(n12274), .CK(clk), .RN(n5857), .Q(
        \I_cache/cache[5][68] ), .QN(n780) );
  DFFRX1 \I_cache/cache_reg[6][68]  ( .D(n12273), .CK(clk), .RN(n5857), .Q(
        \I_cache/cache[6][68] ), .QN(n441) );
  DFFRX1 \I_cache/cache_reg[7][68]  ( .D(n12272), .CK(clk), .RN(n5857), .Q(
        \I_cache/cache[7][68] ), .QN(n2003) );
  DFFRX1 \I_cache/cache_reg[0][69]  ( .D(n12271), .CK(clk), .RN(n5857), .Q(
        \I_cache/cache[0][69] ), .QN(n1133) );
  DFFRX1 \I_cache/cache_reg[1][69]  ( .D(n12270), .CK(clk), .RN(n5857), .Q(
        \I_cache/cache[1][69] ), .QN(n2705) );
  DFFRX1 \I_cache/cache_reg[2][69]  ( .D(n12269), .CK(clk), .RN(n5857), .Q(
        \I_cache/cache[2][69] ), .QN(n1134) );
  DFFRX1 \I_cache/cache_reg[3][69]  ( .D(n12268), .CK(clk), .RN(n5857), .Q(
        \I_cache/cache[3][69] ), .QN(n2706) );
  DFFRX1 \I_cache/cache_reg[4][69]  ( .D(n12267), .CK(clk), .RN(n5857), .Q(
        \I_cache/cache[4][69] ), .QN(n756) );
  DFFRX1 \I_cache/cache_reg[5][69]  ( .D(n12266), .CK(clk), .RN(n5857), .Q(
        \I_cache/cache[5][69] ), .QN(n2334) );
  DFFRX1 \I_cache/cache_reg[6][69]  ( .D(n12265), .CK(clk), .RN(n5857), .Q(
        \I_cache/cache[6][69] ), .QN(n1132) );
  DFFRX1 \I_cache/cache_reg[7][69]  ( .D(n12264), .CK(clk), .RN(n5858), .Q(
        \I_cache/cache[7][69] ), .QN(n2704) );
  DFFRX1 \I_cache/cache_reg[0][70]  ( .D(n12263), .CK(clk), .RN(n5858), .Q(
        \I_cache/cache[0][70] ), .QN(n906) );
  DFFRX1 \I_cache/cache_reg[1][70]  ( .D(n12262), .CK(clk), .RN(n5858), .Q(
        \I_cache/cache[1][70] ), .QN(n2417) );
  DFFRX1 \I_cache/cache_reg[2][70]  ( .D(n12261), .CK(clk), .RN(n5858), .Q(
        \I_cache/cache[2][70] ), .QN(n2424) );
  DFFRX1 \I_cache/cache_reg[3][70]  ( .D(n12260), .CK(clk), .RN(n5858), .Q(
        \I_cache/cache[3][70] ), .QN(n447) );
  DFFRX1 \I_cache/cache_reg[4][70]  ( .D(n12259), .CK(clk), .RN(n5858), .Q(
        \I_cache/cache[4][70] ), .QN(n1044) );
  DFFRX1 \I_cache/cache_reg[5][70]  ( .D(n12258), .CK(clk), .RN(n5858), .Q(
        \I_cache/cache[5][70] ), .QN(n2616) );
  DFFRX1 \I_cache/cache_reg[6][70]  ( .D(n12257), .CK(clk), .RN(n5858), .Q(
        \I_cache/cache[6][70] ), .QN(n2423) );
  DFFRX1 \I_cache/cache_reg[7][70]  ( .D(n12256), .CK(clk), .RN(n5858), .Q(
        \I_cache/cache[7][70] ), .QN(n446) );
  DFFRX1 \I_cache/cache_reg[0][71]  ( .D(n12255), .CK(clk), .RN(n5858), .Q(
        \I_cache/cache[0][71] ), .QN(n1097) );
  DFFRX1 \I_cache/cache_reg[1][71]  ( .D(n12254), .CK(clk), .RN(n5858), .Q(
        \I_cache/cache[1][71] ), .QN(n2669) );
  DFFRX1 \I_cache/cache_reg[2][71]  ( .D(n12253), .CK(clk), .RN(n5858), .Q(
        \I_cache/cache[2][71] ), .QN(n909) );
  DFFRX1 \I_cache/cache_reg[3][71]  ( .D(n12252), .CK(clk), .RN(n5859), .Q(
        \I_cache/cache[3][71] ), .QN(n2426) );
  DFFRX1 \I_cache/cache_reg[4][71]  ( .D(n12251), .CK(clk), .RN(n5859), .Q(
        \I_cache/cache[4][71] ), .QN(n2565) );
  DFFRX1 \I_cache/cache_reg[5][71]  ( .D(n12250), .CK(clk), .RN(n5859), .Q(
        \I_cache/cache[5][71] ), .QN(n794) );
  DFFRX1 \I_cache/cache_reg[6][71]  ( .D(n12249), .CK(clk), .RN(n5859), .Q(
        \I_cache/cache[6][71] ), .QN(n1096) );
  DFFRX1 \I_cache/cache_reg[7][71]  ( .D(n12248), .CK(clk), .RN(n5859), .Q(
        \I_cache/cache[7][71] ), .QN(n2668) );
  DFFRX1 \I_cache/cache_reg[0][72]  ( .D(n12247), .CK(clk), .RN(n5859), .Q(
        \I_cache/cache[0][72] ), .QN(n924) );
  DFFRX1 \I_cache/cache_reg[1][72]  ( .D(n12246), .CK(clk), .RN(n5859), .Q(
        \I_cache/cache[1][72] ), .QN(n2438) );
  DFFRX1 \I_cache/cache_reg[2][72]  ( .D(n12245), .CK(clk), .RN(n5859), .Q(
        \I_cache/cache[2][72] ), .QN(n917) );
  DFFRX1 \I_cache/cache_reg[3][72]  ( .D(n12244), .CK(clk), .RN(n5859), .Q(
        \I_cache/cache[3][72] ), .QN(n2434) );
  DFFRX1 \I_cache/cache_reg[4][72]  ( .D(n12243), .CK(clk), .RN(n5859), .Q(
        \I_cache/cache[4][72] ), .QN(n1192) );
  DFFRX1 \I_cache/cache_reg[5][72]  ( .D(n12242), .CK(clk), .RN(n5859), .Q(
        \I_cache/cache[5][72] ), .QN(n2764) );
  DFFRX1 \I_cache/cache_reg[6][72]  ( .D(n12241), .CK(clk), .RN(n5859), .Q(
        \I_cache/cache[6][72] ), .QN(n2422) );
  DFFRX1 \I_cache/cache_reg[7][72]  ( .D(n12240), .CK(clk), .RN(n5860), .Q(
        \I_cache/cache[7][72] ), .QN(n445) );
  DFFRX1 \I_cache/cache_reg[1][73]  ( .D(n12238), .CK(clk), .RN(n5860), .Q(
        \I_cache/cache[1][73] ), .QN(n2660) );
  DFFRX1 \I_cache/cache_reg[2][73]  ( .D(n12237), .CK(clk), .RN(n5860), .Q(
        \I_cache/cache[2][73] ), .QN(n1089) );
  DFFRX1 \I_cache/cache_reg[3][73]  ( .D(n12236), .CK(clk), .RN(n5860), .Q(
        \I_cache/cache[3][73] ), .QN(n2661) );
  DFFRX1 \I_cache/cache_reg[4][73]  ( .D(n12235), .CK(clk), .RN(n5860), .Q(
        \I_cache/cache[4][73] ), .QN(n749) );
  DFFRX1 \I_cache/cache_reg[6][73]  ( .D(n12233), .CK(clk), .RN(n5860), .Q(
        \I_cache/cache[6][73] ), .QN(n1087) );
  DFFRX1 \I_cache/cache_reg[7][73]  ( .D(n12232), .CK(clk), .RN(n5860), .Q(
        \I_cache/cache[7][73] ), .QN(n2659) );
  DFFRX1 \I_cache/cache_reg[1][74]  ( .D(n12230), .CK(clk), .RN(n5860), .Q(
        \I_cache/cache[1][74] ), .QN(n2418) );
  DFFRX1 \I_cache/cache_reg[2][74]  ( .D(n12229), .CK(clk), .RN(n5860), .Q(
        \I_cache/cache[2][74] ), .QN(n916) );
  DFFRX1 \I_cache/cache_reg[3][74]  ( .D(n12228), .CK(clk), .RN(n5861), .Q(
        \I_cache/cache[3][74] ), .QN(n2433) );
  DFFRX1 \I_cache/cache_reg[4][74]  ( .D(n12227), .CK(clk), .RN(n5861), .Q(
        \I_cache/cache[4][74] ), .QN(n2506) );
  DFFRX1 \I_cache/cache_reg[6][74]  ( .D(n12225), .CK(clk), .RN(n5861), .Q(
        \I_cache/cache[6][74] ), .QN(n915) );
  DFFRX1 \I_cache/cache_reg[7][74]  ( .D(n12224), .CK(clk), .RN(n5861), .Q(
        \I_cache/cache[7][74] ), .QN(n2432) );
  DFFRX1 \I_cache/cache_reg[0][75]  ( .D(n12223), .CK(clk), .RN(n5861), .Q(
        \I_cache/cache[0][75] ), .QN(n1081) );
  DFFRX1 \I_cache/cache_reg[1][75]  ( .D(n12222), .CK(clk), .RN(n5861), .Q(
        \I_cache/cache[1][75] ), .QN(n2653) );
  DFFRX1 \I_cache/cache_reg[2][75]  ( .D(n12221), .CK(clk), .RN(n5861), .Q(
        \I_cache/cache[2][75] ), .QN(n1082) );
  DFFRX1 \I_cache/cache_reg[3][75]  ( .D(n12220), .CK(clk), .RN(n5861), .Q(
        \I_cache/cache[3][75] ), .QN(n2654) );
  DFFRX1 \I_cache/cache_reg[4][75]  ( .D(n12219), .CK(clk), .RN(n5861), .Q(
        \I_cache/cache[4][75] ), .QN(n1086) );
  DFFRX1 \I_cache/cache_reg[5][75]  ( .D(n12218), .CK(clk), .RN(n5861), .Q(
        \I_cache/cache[5][75] ), .QN(n2658) );
  DFFRX1 \I_cache/cache_reg[6][75]  ( .D(n12217), .CK(clk), .RN(n5861), .Q(
        \I_cache/cache[6][75] ), .QN(n1080) );
  DFFRX1 \I_cache/cache_reg[7][75]  ( .D(n12216), .CK(clk), .RN(n5862), .Q(
        \I_cache/cache[7][75] ), .QN(n2652) );
  DFFRX1 \I_cache/cache_reg[0][76]  ( .D(n12215), .CK(clk), .RN(n5862), .Q(
        \I_cache/cache[0][76] ), .QN(n1037) );
  DFFRX1 \I_cache/cache_reg[1][76]  ( .D(n12214), .CK(clk), .RN(n5862), .Q(
        \I_cache/cache[1][76] ), .QN(n2609) );
  DFFRX1 \I_cache/cache_reg[2][76]  ( .D(n12213), .CK(clk), .RN(n5862), .Q(
        \I_cache/cache[2][76] ), .QN(n1038) );
  DFFRX1 \I_cache/cache_reg[3][76]  ( .D(n12212), .CK(clk), .RN(n5862), .Q(
        \I_cache/cache[3][76] ), .QN(n2610) );
  DFFRX1 \I_cache/cache_reg[4][76]  ( .D(n12211), .CK(clk), .RN(n5862), .Q(
        \I_cache/cache[4][76] ), .QN(n1203) );
  DFFRX1 \I_cache/cache_reg[6][76]  ( .D(n12209), .CK(clk), .RN(n5862), .Q(
        \I_cache/cache[6][76] ), .QN(n1053) );
  DFFRX1 \I_cache/cache_reg[0][77]  ( .D(n12207), .CK(clk), .RN(n5862), .Q(
        \I_cache/cache[0][77] ), .QN(n913) );
  DFFRX1 \I_cache/cache_reg[1][77]  ( .D(n12206), .CK(clk), .RN(n5862), .Q(
        \I_cache/cache[1][77] ), .QN(n2430) );
  DFFRX1 \I_cache/cache_reg[2][77]  ( .D(n12205), .CK(clk), .RN(n5862), .Q(
        \I_cache/cache[2][77] ), .QN(n914) );
  DFFRX1 \I_cache/cache_reg[3][77]  ( .D(n12204), .CK(clk), .RN(n5863), .Q(
        \I_cache/cache[3][77] ), .QN(n2431) );
  DFFRX1 \I_cache/cache_reg[4][77]  ( .D(n12203), .CK(clk), .RN(n5863), .Q(
        \I_cache/cache[4][77] ), .QN(n1084) );
  DFFRX1 \I_cache/cache_reg[5][77]  ( .D(n12202), .CK(clk), .RN(n5863), .Q(
        \I_cache/cache[5][77] ), .QN(n2656) );
  DFFRX1 \I_cache/cache_reg[6][77]  ( .D(n12201), .CK(clk), .RN(n5863), .Q(
        \I_cache/cache[6][77] ), .QN(n1092) );
  DFFRX1 \I_cache/cache_reg[7][77]  ( .D(n12200), .CK(clk), .RN(n5863), .Q(
        \I_cache/cache[7][77] ), .QN(n2664) );
  DFFRX1 \I_cache/cache_reg[0][78]  ( .D(n12199), .CK(clk), .RN(n5863), .Q(
        \I_cache/cache[0][78] ), .QN(n1026) );
  DFFRX1 \I_cache/cache_reg[1][78]  ( .D(n12198), .CK(clk), .RN(n5863), .Q(
        \I_cache/cache[1][78] ), .QN(n2598) );
  DFFRX1 \I_cache/cache_reg[2][78]  ( .D(n12197), .CK(clk), .RN(n5863), .Q(
        \I_cache/cache[2][78] ), .QN(n1027) );
  DFFRX1 \I_cache/cache_reg[3][78]  ( .D(n12196), .CK(clk), .RN(n5863), .Q(
        \I_cache/cache[3][78] ), .QN(n2599) );
  DFFRX1 \I_cache/cache_reg[4][78]  ( .D(n12195), .CK(clk), .RN(n5863), .Q(
        \I_cache/cache[4][78] ), .QN(n1200) );
  DFFRX1 \I_cache/cache_reg[5][78]  ( .D(n12194), .CK(clk), .RN(n5863), .Q(
        \I_cache/cache[5][78] ), .QN(n2772) );
  DFFRX1 \I_cache/cache_reg[6][78]  ( .D(n12193), .CK(clk), .RN(n5863), .Q(
        \I_cache/cache[6][78] ), .QN(n1028) );
  DFFRX1 \I_cache/cache_reg[7][78]  ( .D(n12192), .CK(clk), .RN(n5864), .Q(
        \I_cache/cache[7][78] ), .QN(n2600) );
  DFFRX1 \I_cache/cache_reg[0][79]  ( .D(n12191), .CK(clk), .RN(n5864), .Q(
        \I_cache/cache[0][79] ), .QN(n949) );
  DFFRX1 \I_cache/cache_reg[1][79]  ( .D(n12190), .CK(clk), .RN(n5864), .Q(
        \I_cache/cache[1][79] ), .QN(n2474) );
  DFFRX1 \I_cache/cache_reg[2][79]  ( .D(n12189), .CK(clk), .RN(n5864), .Q(
        \I_cache/cache[2][79] ), .QN(n947) );
  DFFRX1 \I_cache/cache_reg[3][79]  ( .D(n12188), .CK(clk), .RN(n5864), .Q(
        \I_cache/cache[3][79] ), .QN(n2472) );
  DFFRX1 \I_cache/cache_reg[4][79]  ( .D(n12187), .CK(clk), .RN(n5864), .Q(
        \I_cache/cache[4][79] ), .QN(n2444) );
  DFFRX1 \I_cache/cache_reg[5][79]  ( .D(n12186), .CK(clk), .RN(n5864), .Q(
        \I_cache/cache[5][79] ), .QN(n469) );
  DFFRX1 \I_cache/cache_reg[6][79]  ( .D(n12185), .CK(clk), .RN(n5864), .Q(
        \I_cache/cache[6][79] ), .QN(n948) );
  DFFRX1 \I_cache/cache_reg[7][79]  ( .D(n12184), .CK(clk), .RN(n5864), .Q(
        \I_cache/cache[7][79] ), .QN(n2473) );
  DFFRX1 \I_cache/cache_reg[0][96]  ( .D(n12055), .CK(clk), .RN(n5875), .Q(
        \I_cache/cache[0][96] ), .QN(n1042) );
  DFFRX1 \I_cache/cache_reg[1][96]  ( .D(n12054), .CK(clk), .RN(n5875), .Q(
        \I_cache/cache[1][96] ), .QN(n2614) );
  DFFRX1 \I_cache/cache_reg[2][96]  ( .D(n12053), .CK(clk), .RN(n5875), .Q(
        \I_cache/cache[2][96] ), .QN(n1043) );
  DFFRX1 \I_cache/cache_reg[3][96]  ( .D(n12052), .CK(clk), .RN(n5875), .Q(
        \I_cache/cache[3][96] ), .QN(n2615) );
  DFFRX1 \I_cache/cache_reg[4][96]  ( .D(n12051), .CK(clk), .RN(n5875), .Q(
        \I_cache/cache[4][96] ), .QN(n1198) );
  DFFRX1 \I_cache/cache_reg[5][96]  ( .D(n12050), .CK(clk), .RN(n5875), .Q(
        \I_cache/cache[5][96] ), .QN(n2770) );
  DFFRX1 \I_cache/cache_reg[6][96]  ( .D(n12049), .CK(clk), .RN(n5875), .Q(
        \I_cache/cache[6][96] ), .QN(n2519) );
  DFFRX1 \I_cache/cache_reg[7][96]  ( .D(n12048), .CK(clk), .RN(n5876), .Q(
        \I_cache/cache[7][96] ), .QN(n768) );
  DFFRX1 \I_cache/cache_reg[0][97]  ( .D(n12047), .CK(clk), .RN(n5876), .Q(
        \I_cache/cache[0][97] ), .QN(n1141) );
  DFFRX1 \I_cache/cache_reg[1][97]  ( .D(n12046), .CK(clk), .RN(n5876), .Q(
        \I_cache/cache[1][97] ), .QN(n2713) );
  DFFRX1 \I_cache/cache_reg[2][97]  ( .D(n12045), .CK(clk), .RN(n5876), .Q(
        \I_cache/cache[2][97] ), .QN(n1142) );
  DFFRX1 \I_cache/cache_reg[3][97]  ( .D(n12044), .CK(clk), .RN(n5876), .Q(
        \I_cache/cache[3][97] ), .QN(n2714) );
  DFFRX1 \I_cache/cache_reg[4][97]  ( .D(n12043), .CK(clk), .RN(n5876), .Q(
        \I_cache/cache[4][97] ), .QN(n1222) );
  DFFRX1 \I_cache/cache_reg[6][97]  ( .D(n12041), .CK(clk), .RN(n5876), .Q(
        \I_cache/cache[6][97] ), .QN(n1140) );
  DFFRX1 \I_cache/cache_reg[0][98]  ( .D(n12039), .CK(clk), .RN(n5876), .Q(
        \I_cache/cache[0][98] ), .QN(n1070) );
  DFFRX1 \I_cache/cache_reg[1][98]  ( .D(n12038), .CK(clk), .RN(n5876), .Q(
        \I_cache/cache[1][98] ), .QN(n2642) );
  DFFRX1 \I_cache/cache_reg[2][98]  ( .D(n12037), .CK(clk), .RN(n5876), .Q(
        \I_cache/cache[2][98] ), .QN(n1068) );
  DFFRX1 \I_cache/cache_reg[3][98]  ( .D(n12036), .CK(clk), .RN(n5877), .Q(
        \I_cache/cache[3][98] ), .QN(n2640) );
  DFFRX1 \I_cache/cache_reg[4][98]  ( .D(n12035), .CK(clk), .RN(n5877), .Q(
        \I_cache/cache[4][98] ), .QN(n2537) );
  DFFRX1 \I_cache/cache_reg[5][98]  ( .D(n12034), .CK(clk), .RN(n5877), .Q(
        \I_cache/cache[5][98] ), .QN(n778) );
  DFFRX1 \I_cache/cache_reg[6][98]  ( .D(n12033), .CK(clk), .RN(n5877), .Q(
        \I_cache/cache[6][98] ), .QN(n1069) );
  DFFRX1 \I_cache/cache_reg[7][98]  ( .D(n12032), .CK(clk), .RN(n5877), .Q(
        \I_cache/cache[7][98] ), .QN(n2641) );
  DFFRX1 \I_cache/cache_reg[0][99]  ( .D(n12031), .CK(clk), .RN(n5877), .Q(
        \I_cache/cache[0][99] ), .QN(n738) );
  DFFRX1 \I_cache/cache_reg[1][99]  ( .D(n12030), .CK(clk), .RN(n5877), .Q(
        \I_cache/cache[1][99] ), .QN(n2319) );
  DFFRX1 \I_cache/cache_reg[2][99]  ( .D(n12029), .CK(clk), .RN(n5877), .Q(
        \I_cache/cache[2][99] ), .QN(n739) );
  DFFRX1 \I_cache/cache_reg[3][99]  ( .D(n12028), .CK(clk), .RN(n5877), .Q(
        \I_cache/cache[3][99] ), .QN(n2320) );
  DFFRX1 \I_cache/cache_reg[4][99]  ( .D(n12027), .CK(clk), .RN(n5877), .Q(
        \I_cache/cache[4][99] ), .QN(n736) );
  DFFRX1 \I_cache/cache_reg[5][99]  ( .D(n12026), .CK(clk), .RN(n5877), .Q(
        \I_cache/cache[5][99] ), .QN(n2317) );
  DFFRX1 \I_cache/cache_reg[6][99]  ( .D(n12025), .CK(clk), .RN(n5877), .Q(
        \I_cache/cache[6][99] ), .QN(n1934) );
  DFFRX1 \I_cache/cache_reg[7][99]  ( .D(n12024), .CK(clk), .RN(n5878), .Q(
        \I_cache/cache[7][99] ), .QN(n353) );
  DFFRX1 \I_cache/cache_reg[0][100]  ( .D(n12023), .CK(clk), .RN(n5878), .Q(
        \I_cache/cache[0][100] ), .QN(n1115) );
  DFFRX1 \I_cache/cache_reg[1][100]  ( .D(n12022), .CK(clk), .RN(n5878), .Q(
        \I_cache/cache[1][100] ), .QN(n2687) );
  DFFRX1 \I_cache/cache_reg[2][100]  ( .D(n12021), .CK(clk), .RN(n5878), .Q(
        \I_cache/cache[2][100] ), .QN(n1116) );
  DFFRX1 \I_cache/cache_reg[3][100]  ( .D(n12020), .CK(clk), .RN(n5878), .Q(
        \I_cache/cache[3][100] ), .QN(n2688) );
  DFFRX1 \I_cache/cache_reg[4][100]  ( .D(n12019), .CK(clk), .RN(n5878), .Q(
        \I_cache/cache[4][100] ), .QN(n752) );
  DFFRX1 \I_cache/cache_reg[5][100]  ( .D(n12018), .CK(clk), .RN(n5878), .Q(
        \I_cache/cache[5][100] ), .QN(n2330) );
  DFFRX1 \I_cache/cache_reg[6][100]  ( .D(n12017), .CK(clk), .RN(n5878), .Q(
        \I_cache/cache[6][100] ), .QN(n2556) );
  DFFRX1 \I_cache/cache_reg[7][100]  ( .D(n12016), .CK(clk), .RN(n5878), .Q(
        \I_cache/cache[7][100] ), .QN(n785) );
  DFFRX1 \I_cache/cache_reg[0][101]  ( .D(n12015), .CK(clk), .RN(n5878), .Q(
        \I_cache/cache[0][101] ), .QN(n1144) );
  DFFRX1 \I_cache/cache_reg[1][101]  ( .D(n12014), .CK(clk), .RN(n5878), .Q(
        \I_cache/cache[1][101] ), .QN(n2716) );
  DFFRX1 \I_cache/cache_reg[2][101]  ( .D(n12013), .CK(clk), .RN(n5878), .Q(
        \I_cache/cache[2][101] ), .QN(n1145) );
  DFFRX1 \I_cache/cache_reg[3][101]  ( .D(n12012), .CK(clk), .RN(n5879), .Q(
        \I_cache/cache[3][101] ), .QN(n2717) );
  DFFRX1 \I_cache/cache_reg[4][101]  ( .D(n12011), .CK(clk), .RN(n5879), .Q(
        \I_cache/cache[4][101] ), .QN(n737) );
  DFFRX1 \I_cache/cache_reg[5][101]  ( .D(n12010), .CK(clk), .RN(n5879), .Q(
        \I_cache/cache[5][101] ), .QN(n2318) );
  DFFRX1 \I_cache/cache_reg[6][101]  ( .D(n12009), .CK(clk), .RN(n5879), .Q(
        \I_cache/cache[6][101] ), .QN(n1143) );
  DFFRX1 \I_cache/cache_reg[7][101]  ( .D(n12008), .CK(clk), .RN(n5879), .Q(
        \I_cache/cache[7][101] ), .QN(n2715) );
  DFFRX1 \I_cache/cache_reg[0][102]  ( .D(n12007), .CK(clk), .RN(n5879), .Q(
        \I_cache/cache[0][102] ), .QN(n1103) );
  DFFRX1 \I_cache/cache_reg[1][102]  ( .D(n12006), .CK(clk), .RN(n5879), .Q(
        \I_cache/cache[1][102] ), .QN(n2675) );
  DFFRX1 \I_cache/cache_reg[2][102]  ( .D(n12005), .CK(clk), .RN(n5879), .Q(
        \I_cache/cache[2][102] ), .QN(n1104) );
  DFFRX1 \I_cache/cache_reg[3][102]  ( .D(n12004), .CK(clk), .RN(n5879), .Q(
        \I_cache/cache[3][102] ), .QN(n2676) );
  DFFRX1 \I_cache/cache_reg[4][102]  ( .D(n12003), .CK(clk), .RN(n5879), .Q(
        \I_cache/cache[4][102] ), .QN(n1190) );
  DFFRX1 \I_cache/cache_reg[5][102]  ( .D(n12002), .CK(clk), .RN(n5879), .Q(
        \I_cache/cache[5][102] ), .QN(n2762) );
  DFFRX1 \I_cache/cache_reg[6][102]  ( .D(n12001), .CK(clk), .RN(n5879), .Q(
        \I_cache/cache[6][102] ), .QN(n1102) );
  DFFRX1 \I_cache/cache_reg[7][102]  ( .D(n12000), .CK(clk), .RN(n5880), .Q(
        \I_cache/cache[7][102] ), .QN(n2674) );
  DFFRX1 \I_cache/cache_reg[0][103]  ( .D(n11999), .CK(clk), .RN(n5880), .Q(
        \I_cache/cache[0][103] ), .QN(n1078) );
  DFFRX1 \I_cache/cache_reg[1][103]  ( .D(n11998), .CK(clk), .RN(n5880), .Q(
        \I_cache/cache[1][103] ), .QN(n2650) );
  DFFRX1 \I_cache/cache_reg[2][103]  ( .D(n11997), .CK(clk), .RN(n5880), .Q(
        \I_cache/cache[2][103] ), .QN(n1079) );
  DFFRX1 \I_cache/cache_reg[3][103]  ( .D(n11996), .CK(clk), .RN(n5880), .Q(
        \I_cache/cache[3][103] ), .QN(n2651) );
  DFFRX1 \I_cache/cache_reg[4][103]  ( .D(n11995), .CK(clk), .RN(n5880), .Q(
        \I_cache/cache[4][103] ), .QN(n979) );
  DFFRX1 \I_cache/cache_reg[5][103]  ( .D(n11994), .CK(clk), .RN(n5880), .Q(
        \I_cache/cache[5][103] ), .QN(n2525) );
  DFFRX1 \I_cache/cache_reg[6][103]  ( .D(n11993), .CK(clk), .RN(n5880), .Q(
        \I_cache/cache[6][103] ), .QN(n1077) );
  DFFRX1 \I_cache/cache_reg[7][103]  ( .D(n11992), .CK(clk), .RN(n5880), .Q(
        \I_cache/cache[7][103] ), .QN(n2649) );
  DFFRX1 \I_cache/cache_reg[0][104]  ( .D(n11991), .CK(clk), .RN(n5880), .Q(
        \I_cache/cache[0][104] ), .QN(n1113) );
  DFFRX1 \I_cache/cache_reg[1][104]  ( .D(n11990), .CK(clk), .RN(n5880), .Q(
        \I_cache/cache[1][104] ), .QN(n2685) );
  DFFRX1 \I_cache/cache_reg[2][104]  ( .D(n11989), .CK(clk), .RN(n5880), .Q(
        \I_cache/cache[2][104] ), .QN(n1114) );
  DFFRX1 \I_cache/cache_reg[3][104]  ( .D(n11988), .CK(clk), .RN(n5881), .Q(
        \I_cache/cache[3][104] ), .QN(n2686) );
  DFFRX1 \I_cache/cache_reg[4][104]  ( .D(n11987), .CK(clk), .RN(n5881), .Q(
        \I_cache/cache[4][104] ), .QN(n1085) );
  DFFRX1 \I_cache/cache_reg[5][104]  ( .D(n11986), .CK(clk), .RN(n5881), .Q(
        \I_cache/cache[5][104] ), .QN(n2657) );
  DFFRX1 \I_cache/cache_reg[6][104]  ( .D(n11985), .CK(clk), .RN(n5881), .Q(
        \I_cache/cache[6][104] ), .QN(n2555) );
  DFFRX1 \I_cache/cache_reg[7][104]  ( .D(n11984), .CK(clk), .RN(n5881), .Q(
        \I_cache/cache[7][104] ), .QN(n784) );
  DFFRX1 \I_cache/cache_reg[1][105]  ( .D(n11982), .CK(clk), .RN(n5881), .Q(
        \I_cache/cache[1][105] ), .QN(n2648) );
  DFFRX1 \I_cache/cache_reg[2][105]  ( .D(n11981), .CK(clk), .RN(n5881), .Q(
        \I_cache/cache[2][105] ), .QN(n1075) );
  DFFRX1 \I_cache/cache_reg[3][105]  ( .D(n11980), .CK(clk), .RN(n5881), .Q(
        \I_cache/cache[3][105] ), .QN(n2647) );
  DFFRX1 \I_cache/cache_reg[4][105]  ( .D(n11979), .CK(clk), .RN(n5881), .Q(
        \I_cache/cache[4][105] ), .QN(n2507) );
  DFFRX1 \I_cache/cache_reg[6][105]  ( .D(n11977), .CK(clk), .RN(n5881), .Q(
        \I_cache/cache[6][105] ), .QN(n440) );
  DFFRX1 \I_cache/cache_reg[7][105]  ( .D(n11976), .CK(clk), .RN(n5882), .Q(
        \I_cache/cache[7][105] ), .QN(n2002) );
  DFFRX1 \I_cache/cache_reg[0][106]  ( .D(n11975), .CK(clk), .RN(n5882), .Q(
        \I_cache/cache[0][106] ), .QN(n991) );
  DFFRX1 \I_cache/cache_reg[1][106]  ( .D(n11974), .CK(clk), .RN(n5882), .Q(
        \I_cache/cache[1][106] ), .QN(n2543) );
  DFFRX1 \I_cache/cache_reg[2][106]  ( .D(n11973), .CK(clk), .RN(n5882), .Q(
        \I_cache/cache[2][106] ), .QN(n992) );
  DFFRX1 \I_cache/cache_reg[3][106]  ( .D(n11972), .CK(clk), .RN(n5882), .Q(
        \I_cache/cache[3][106] ), .QN(n2544) );
  DFFRX1 \I_cache/cache_reg[4][106]  ( .D(n11971), .CK(clk), .RN(n5882), .Q(
        \I_cache/cache[4][106] ), .QN(n1059) );
  DFFRX1 \I_cache/cache_reg[5][106]  ( .D(n11970), .CK(clk), .RN(n5882), .Q(
        \I_cache/cache[5][106] ), .QN(n2631) );
  DFFRX1 \I_cache/cache_reg[6][106]  ( .D(n11969), .CK(clk), .RN(n5882), .Q(
        \I_cache/cache[6][106] ), .QN(n990) );
  DFFRX1 \I_cache/cache_reg[7][106]  ( .D(n11968), .CK(clk), .RN(n5882), .Q(
        \I_cache/cache[7][106] ), .QN(n2542) );
  DFFRX1 \I_cache/cache_reg[0][107]  ( .D(n11967), .CK(clk), .RN(n5882), .Q(
        \I_cache/cache[0][107] ), .QN(n986) );
  DFFRX1 \I_cache/cache_reg[1][107]  ( .D(n11966), .CK(clk), .RN(n5882), .Q(
        \I_cache/cache[1][107] ), .QN(n2535) );
  DFFRX1 \I_cache/cache_reg[2][107]  ( .D(n11965), .CK(clk), .RN(n5882), .Q(
        \I_cache/cache[2][107] ), .QN(n984) );
  DFFRX1 \I_cache/cache_reg[3][107]  ( .D(n11964), .CK(clk), .RN(n5883), .Q(
        \I_cache/cache[3][107] ), .QN(n2533) );
  DFFRX1 \I_cache/cache_reg[4][107]  ( .D(n11963), .CK(clk), .RN(n5883), .Q(
        \I_cache/cache[4][107] ), .QN(n997) );
  DFFRX1 \I_cache/cache_reg[5][107]  ( .D(n11962), .CK(clk), .RN(n5883), .Q(
        \I_cache/cache[5][107] ), .QN(n2549) );
  DFFRX1 \I_cache/cache_reg[6][107]  ( .D(n11961), .CK(clk), .RN(n5883), .Q(
        \I_cache/cache[6][107] ), .QN(n985) );
  DFFRX1 \I_cache/cache_reg[7][107]  ( .D(n11960), .CK(clk), .RN(n5883), .Q(
        \I_cache/cache[7][107] ), .QN(n2534) );
  DFFRX1 \I_cache/cache_reg[0][108]  ( .D(n11959), .CK(clk), .RN(n5883), .Q(
        \I_cache/cache[0][108] ), .QN(n1032) );
  DFFRX1 \I_cache/cache_reg[1][108]  ( .D(n11958), .CK(clk), .RN(n5883), .Q(
        \I_cache/cache[1][108] ), .QN(n2604) );
  DFFRX1 \I_cache/cache_reg[2][108]  ( .D(n11957), .CK(clk), .RN(n5883), .Q(
        \I_cache/cache[2][108] ), .QN(n1033) );
  DFFRX1 \I_cache/cache_reg[3][108]  ( .D(n11956), .CK(clk), .RN(n5883), .Q(
        \I_cache/cache[3][108] ), .QN(n2605) );
  DFFRX1 \I_cache/cache_reg[4][108]  ( .D(n11955), .CK(clk), .RN(n5883), .Q(
        \I_cache/cache[4][108] ), .QN(n1050) );
  DFFRX1 \I_cache/cache_reg[6][108]  ( .D(n11953), .CK(clk), .RN(n5883), .Q(
        \I_cache/cache[6][108] ), .QN(n910) );
  DFFRX1 \I_cache/cache_reg[0][109]  ( .D(n11951), .CK(clk), .RN(n5884), .Q(
        \I_cache/cache[0][109] ), .QN(n1055) );
  DFFRX1 \I_cache/cache_reg[1][109]  ( .D(n11950), .CK(clk), .RN(n5884), .Q(
        \I_cache/cache[1][109] ), .QN(n2627) );
  DFFRX1 \I_cache/cache_reg[2][109]  ( .D(n11949), .CK(clk), .RN(n5884), .Q(
        \I_cache/cache[2][109] ), .QN(n1056) );
  DFFRX1 \I_cache/cache_reg[3][109]  ( .D(n11948), .CK(clk), .RN(n5884), .Q(
        \I_cache/cache[3][109] ), .QN(n2628) );
  DFFRX1 \I_cache/cache_reg[4][109]  ( .D(n11947), .CK(clk), .RN(n5884), .Q(
        \I_cache/cache[4][109] ), .QN(n1058) );
  DFFRX1 \I_cache/cache_reg[5][109]  ( .D(n11946), .CK(clk), .RN(n5884), .Q(
        \I_cache/cache[5][109] ), .QN(n2630) );
  DFFRX1 \I_cache/cache_reg[6][109]  ( .D(n11945), .CK(clk), .RN(n5884), .Q(
        \I_cache/cache[6][109] ), .QN(n1054) );
  DFFRX1 \I_cache/cache_reg[7][109]  ( .D(n11944), .CK(clk), .RN(n5884), .Q(
        \I_cache/cache[7][109] ), .QN(n2626) );
  DFFRX1 \I_cache/cache_reg[0][110]  ( .D(n11943), .CK(clk), .RN(n5884), .Q(
        \I_cache/cache[0][110] ), .QN(n1020) );
  DFFRX1 \I_cache/cache_reg[1][110]  ( .D(n11942), .CK(clk), .RN(n5884), .Q(
        \I_cache/cache[1][110] ), .QN(n2592) );
  DFFRX1 \I_cache/cache_reg[2][110]  ( .D(n11941), .CK(clk), .RN(n5884), .Q(
        \I_cache/cache[2][110] ), .QN(n1021) );
  DFFRX1 \I_cache/cache_reg[3][110]  ( .D(n11940), .CK(clk), .RN(n5885), .Q(
        \I_cache/cache[3][110] ), .QN(n2593) );
  DFFRX1 \I_cache/cache_reg[4][110]  ( .D(n11939), .CK(clk), .RN(n5885), .Q(
        \I_cache/cache[4][110] ), .QN(n983) );
  DFFRX1 \I_cache/cache_reg[5][110]  ( .D(n11938), .CK(clk), .RN(n5885), .Q(
        \I_cache/cache[5][110] ), .QN(n2531) );
  DFFRX1 \I_cache/cache_reg[6][110]  ( .D(n11937), .CK(clk), .RN(n5885), .Q(
        \I_cache/cache[6][110] ), .QN(n1022) );
  DFFRX1 \I_cache/cache_reg[7][110]  ( .D(n11936), .CK(clk), .RN(n5885), .Q(
        \I_cache/cache[7][110] ), .QN(n2594) );
  DFFRX1 \I_cache/cache_reg[0][111]  ( .D(n11935), .CK(clk), .RN(n5885), .Q(
        \I_cache/cache[0][111] ), .QN(n1488) );
  DFFRX1 \I_cache/cache_reg[1][111]  ( .D(n11934), .CK(clk), .RN(n5885), .Q(
        \I_cache/cache[1][111] ), .QN(n3101) );
  DFFRX1 \I_cache/cache_reg[2][111]  ( .D(n11933), .CK(clk), .RN(n5885), .Q(
        \I_cache/cache[2][111] ), .QN(n1489) );
  DFFRX1 \I_cache/cache_reg[3][111]  ( .D(n11932), .CK(clk), .RN(n5885), .Q(
        \I_cache/cache[3][111] ), .QN(n3102) );
  DFFRX1 \I_cache/cache_reg[4][111]  ( .D(n11931), .CK(clk), .RN(n5885), .Q(
        \I_cache/cache[4][111] ), .QN(n817) );
  DFFRX1 \I_cache/cache_reg[5][111]  ( .D(n11930), .CK(clk), .RN(n5885), .Q(
        \I_cache/cache[5][111] ), .QN(n2349) );
  DFFRX1 \I_cache/cache_reg[6][111]  ( .D(n11929), .CK(clk), .RN(n5885), .Q(
        \I_cache/cache[6][111] ), .QN(n2857) );
  DFFRX1 \I_cache/cache_reg[7][111]  ( .D(n11928), .CK(clk), .RN(n5886), .Q(
        \I_cache/cache[7][111] ), .QN(n848) );
  DFFRX1 \I_cache/cache_reg[0][153]  ( .D(n11599), .CK(clk), .RN(n5913), .Q(
        \I_cache/cache[0][153] ), .QN(n2336) );
  DFFRX1 \I_cache/cache_reg[1][153]  ( .D(n11598), .CK(clk), .RN(n5913), .Q(
        \I_cache/cache[1][153] ), .QN(n800) );
  DFFRX1 \I_cache/cache_reg[2][153]  ( .D(n11597), .CK(clk), .RN(n5913), .Q(
        \I_cache/cache[2][153] ), .QN(n2338) );
  DFFRX1 \I_cache/cache_reg[3][153]  ( .D(n11596), .CK(clk), .RN(n5913), .Q(
        \I_cache/cache[3][153] ), .QN(n802) );
  DFFRX1 \I_cache/cache_reg[4][153]  ( .D(n11595), .CK(clk), .RN(n5913), .Q(
        \I_cache/cache[4][153] ), .QN(n1220) );
  DFFRX1 \I_cache/cache_reg[5][153]  ( .D(n11594), .CK(clk), .RN(n5913), .Q(
        \I_cache/cache[5][153] ), .QN(n2792) );
  DFFRX1 \I_cache/cache_reg[6][153]  ( .D(n11593), .CK(clk), .RN(n5913), .Q(
        \I_cache/cache[6][153] ), .QN(n1052) );
  DFFRX1 \I_cache/cache_reg[7][153]  ( .D(n11592), .CK(clk), .RN(n5913), .Q(
        \I_cache/cache[7][153] ), .QN(n2624) );
  DFFRX1 \I_cache/cache_reg[4][128]  ( .D(n11795), .CK(clk), .RN(n5897), .Q(
        \I_cache/cache[4][128] ), .QN(n3285) );
  DFFRX1 \I_cache/cache_reg[4][139]  ( .D(n11707), .CK(clk), .RN(n5904), .Q(
        \I_cache/cache[4][139] ) );
  DFFRX1 \I_cache/cache_reg[4][131]  ( .D(n11771), .CK(clk), .RN(n5899), .Q(
        \I_cache/cache[4][131] ), .QN(n458) );
  DFFRX1 \I_cache/cache_reg[0][131]  ( .D(n11775), .CK(clk), .RN(n5898), .Q(
        \I_cache/cache[0][131] ), .QN(n457) );
  DFFRX1 \I_cache/cache_reg[5][151]  ( .D(n11610), .CK(clk), .RN(n5912), .Q(
        \I_cache/cache[5][151] ), .QN(n3213) );
  DFFRX1 \I_cache/cache_reg[6][132]  ( .D(n11761), .CK(clk), .RN(n5899), .Q(
        \I_cache/cache[6][132] ), .QN(n308) );
  DFFRX1 \I_cache/cache_reg[5][129]  ( .D(n11786), .CK(clk), .RN(n5897), .Q(
        \I_cache/cache[5][129] ), .QN(n356) );
  DFFRX1 \I_cache/cache_reg[2][131]  ( .D(n11773), .CK(clk), .RN(n5898), .Q(
        \I_cache/cache[2][131] ), .QN(n1962) );
  DFFRX1 \I_cache/cache_reg[1][132]  ( .D(n11766), .CK(clk), .RN(n5899), .Q(
        \I_cache/cache[1][132] ), .QN(n323) );
  DFFRX1 \I_cache/cache_reg[2][129]  ( .D(n11789), .CK(clk), .RN(n5897), .Q(
        \I_cache/cache[2][129] ), .QN(n3274) );
  DFFRX1 \I_cache/cache_reg[0][133]  ( .D(n11759), .CK(clk), .RN(n5900), .Q(
        \I_cache/cache[0][133] ), .QN(n1952) );
  DFFRX1 \I_cache/cache_reg[5][131]  ( .D(n11770), .CK(clk), .RN(n5899), .Q(
        \I_cache/cache[5][131] ), .QN(n2012) );
  DFFRX1 \I_cache/cache_reg[5][132]  ( .D(n11762), .CK(clk), .RN(n5899), .Q(
        \I_cache/cache[5][132] ), .QN(n1583) );
  DFFRX1 \I_cache/cache_reg[6][131]  ( .D(n11769), .CK(clk), .RN(n5899), .Q(
        \I_cache/cache[6][131] ), .QN(n2021) );
  DFFRX1 \I_cache/cache_reg[0][134]  ( .D(n11751), .CK(clk), .RN(n5900), .Q(
        \I_cache/cache[0][134] ), .QN(n1984) );
  DFFRX1 \I_cache/cache_reg[1][131]  ( .D(n11774), .CK(clk), .RN(n5898), .Q(
        \I_cache/cache[1][131] ), .QN(n2011) );
  DFFRX1 \I_cache/cache_reg[4][134]  ( .D(n11747), .CK(clk), .RN(n5901), .Q(
        \I_cache/cache[4][134] ), .QN(n3275) );
  DFFRX1 \I_cache/cache_reg[7][129]  ( .D(n11784), .CK(clk), .RN(n5897), .Q(
        \I_cache/cache[7][129] ), .QN(n359) );
  DFFRX1 \I_cache/cache_reg[0][146]  ( .D(n11655), .CK(clk), .RN(n5908), .Q(
        \I_cache/cache[0][146] ), .QN(n1981) );
  DFFRX1 \I_cache/cache_reg[4][130]  ( .D(n11779), .CK(clk), .RN(n5898), .Q(
        \I_cache/cache[4][130] ), .QN(n3280) );
  DFFRX1 \I_cache/cache_reg[3][132]  ( .D(n11764), .CK(clk), .RN(n5899), .Q(
        \I_cache/cache[3][132] ), .QN(n324) );
  DFFRX1 \I_cache/cache_reg[0][138]  ( .D(n11719), .CK(clk), .RN(n5903), .Q(
        \I_cache/cache[0][138] ), .QN(n1951) );
  DFFRX1 \I_cache/cache_reg[3][131]  ( .D(n11772), .CK(clk), .RN(n5898), .Q(
        \I_cache/cache[3][131] ), .QN(n390) );
  DFFRX1 \D_cache/cache_reg[2][129]  ( .D(\D_cache/n762 ), .CK(clk), .RN(n5794), .Q(\D_cache/cache[2][129] ), .QN(n1936) );
  DFFRX1 \D_cache/cache_reg[3][129]  ( .D(\D_cache/n761 ), .CK(clk), .RN(n5794), .Q(\D_cache/cache[3][129] ), .QN(n355) );
  DFFRX1 \D_cache/cache_reg[6][129]  ( .D(\D_cache/n758 ), .CK(clk), .RN(n5794), .Q(\D_cache/cache[6][129] ), .QN(n1898) );
  DFFRX1 \D_cache/cache_reg[7][129]  ( .D(\D_cache/n757 ), .CK(clk), .RN(n5794), .Q(\D_cache/cache[7][129] ) );
  DFFRX1 \D_cache/cache_reg[2][130]  ( .D(\D_cache/n754 ), .CK(clk), .RN(n5794), .Q(\D_cache/cache[2][130] ), .QN(n314) );
  DFFRX1 \D_cache/cache_reg[3][130]  ( .D(\D_cache/n753 ), .CK(clk), .RN(n5794), .Q(\D_cache/cache[3][130] ), .QN(n1889) );
  DFFRX1 \D_cache/cache_reg[5][130]  ( .D(\D_cache/n751 ), .CK(clk), .RN(n5795), .Q(\D_cache/cache[5][130] ), .QN(n3248) );
  DFFRX1 \D_cache/cache_reg[6][130]  ( .D(\D_cache/n750 ), .CK(clk), .RN(n5795), .Q(\D_cache/cache[6][130] ), .QN(n1894) );
  DFFRX1 \D_cache/cache_reg[7][130]  ( .D(\D_cache/n749 ), .CK(clk), .RN(n5795), .Q(\D_cache/cache[7][130] ), .QN(n1878) );
  DFFRX1 \D_cache/cache_reg[2][131]  ( .D(\D_cache/n746 ), .CK(clk), .RN(n5795), .Q(\D_cache/cache[2][131] ), .QN(n1935) );
  DFFRX1 \D_cache/cache_reg[3][131]  ( .D(\D_cache/n745 ), .CK(clk), .RN(n5795), .Q(\D_cache/cache[3][131] ), .QN(n354) );
  DFFRX1 \D_cache/cache_reg[5][131]  ( .D(\D_cache/n743 ), .CK(clk), .RN(n5795), .Q(\D_cache/cache[5][131] ), .QN(n2800) );
  DFFRX1 \D_cache/cache_reg[6][131]  ( .D(\D_cache/n742 ), .CK(clk), .RN(n5795), .Q(\D_cache/cache[6][131] ), .QN(n1900) );
  DFFRX1 \D_cache/cache_reg[7][132]  ( .D(\D_cache/n733 ), .CK(clk), .RN(n5796), .Q(\D_cache/cache[7][132] ), .QN(n406) );
  DFFRX1 \D_cache/cache_reg[3][133]  ( .D(\D_cache/n729 ), .CK(clk), .RN(n5796), .Q(\D_cache/cache[3][133] ), .QN(n2005) );
  DFFRX1 \D_cache/cache_reg[6][133]  ( .D(\D_cache/n726 ), .CK(clk), .RN(n5797), .Q(\D_cache/cache[6][133] ), .QN(n1963) );
  DFFRX1 \D_cache/cache_reg[7][133]  ( .D(\D_cache/n725 ), .CK(clk), .RN(n5797), .Q(\D_cache/cache[7][133] ), .QN(n391) );
  DFFRX1 \D_cache/cache_reg[3][134]  ( .D(\D_cache/n721 ), .CK(clk), .RN(n5797), .Q(\D_cache/cache[3][134] ), .QN(n2007) );
  DFFRX1 \D_cache/cache_reg[6][134]  ( .D(\D_cache/n718 ), .CK(clk), .RN(n5797), .Q(\D_cache/cache[6][134] ), .QN(n452) );
  DFFRX1 \D_cache/cache_reg[7][134]  ( .D(\D_cache/n717 ), .CK(clk), .RN(n5797), .Q(\D_cache/cache[7][134] ), .QN(n2008) );
  DFFRX1 \D_cache/cache_reg[7][135]  ( .D(\D_cache/n709 ), .CK(clk), .RN(n5798), .Q(\D_cache/cache[7][135] ), .QN(n3264) );
  DFFRX1 \D_cache/cache_reg[7][137]  ( .D(\D_cache/n693 ), .CK(clk), .RN(n5799), .Q(\D_cache/cache[7][137] ), .QN(n3263) );
  DFFRX1 \D_cache/cache_reg[2][138]  ( .D(\D_cache/n690 ), .CK(clk), .RN(n5800), .Q(\D_cache/cache[2][138] ), .QN(n2401) );
  DFFRX1 \D_cache/cache_reg[3][138]  ( .D(\D_cache/n689 ), .CK(clk), .RN(n5800), .Q(\D_cache/cache[3][138] ), .QN(n379) );
  DFFRX1 \D_cache/cache_reg[6][138]  ( .D(\D_cache/n686 ), .CK(clk), .RN(n5800), .Q(\D_cache/cache[6][138] ), .QN(n1945) );
  DFFRX1 \D_cache/cache_reg[7][138]  ( .D(\D_cache/n685 ), .CK(clk), .RN(n5800), .Q(\D_cache/cache[7][138] ), .QN(n367) );
  DFFRX1 \D_cache/cache_reg[1][139]  ( .D(\D_cache/n683 ), .CK(clk), .RN(n5800), .Q(\D_cache/cache[1][139] ), .QN(n321) );
  DFFRX1 \D_cache/cache_reg[2][139]  ( .D(\D_cache/n682 ), .CK(clk), .RN(n5800), .Q(\D_cache/cache[2][139] ), .QN(n1955) );
  DFFRX1 \D_cache/cache_reg[3][139]  ( .D(\D_cache/n681 ), .CK(clk), .RN(n5800), .Q(\D_cache/cache[3][139] ), .QN(n380) );
  DFFRX1 \D_cache/cache_reg[5][139]  ( .D(\D_cache/n679 ), .CK(clk), .RN(n5801), .Q(\D_cache/cache[5][139] ), .QN(n1991) );
  DFFRX1 \D_cache/cache_reg[6][139]  ( .D(\D_cache/n678 ), .CK(clk), .RN(n5801), .Q(\D_cache/cache[6][139] ), .QN(n1957) );
  DFFRX1 \D_cache/cache_reg[7][139]  ( .D(\D_cache/n677 ), .CK(clk), .RN(n5801), .Q(\D_cache/cache[7][139] ), .QN(n385) );
  DFFRX1 \D_cache/cache_reg[0][140]  ( .D(\D_cache/n676 ), .CK(clk), .RN(n5801), .Q(\D_cache/cache[0][140] ), .QN(n1884) );
  DFFRX1 \D_cache/cache_reg[1][140]  ( .D(\D_cache/n675 ), .CK(clk), .RN(n5801), .Q(\D_cache/cache[1][140] ), .QN(n253) );
  DFFRX1 \D_cache/cache_reg[2][140]  ( .D(\D_cache/n674 ), .CK(clk), .RN(n5801), .Q(\D_cache/cache[2][140] ), .QN(n1947) );
  DFFRX1 \D_cache/cache_reg[3][140]  ( .D(\D_cache/n673 ), .CK(clk), .RN(n5801), .Q(\D_cache/cache[3][140] ), .QN(n369) );
  DFFRX1 \D_cache/cache_reg[4][140]  ( .D(\D_cache/n672 ), .CK(clk), .RN(n5801), .Q(\D_cache/cache[4][140] ), .QN(n1883) );
  DFFRX1 \D_cache/cache_reg[5][140]  ( .D(\D_cache/n671 ), .CK(clk), .RN(n5801), .Q(\D_cache/cache[5][140] ), .QN(n317) );
  DFFRX1 \D_cache/cache_reg[6][140]  ( .D(\D_cache/n670 ), .CK(clk), .RN(n5801), .Q(\D_cache/cache[6][140] ), .QN(n1975) );
  DFFRX1 \D_cache/cache_reg[7][140]  ( .D(\D_cache/n669 ), .CK(clk), .RN(n5801), .Q(\D_cache/cache[7][140] ), .QN(n407) );
  DFFRX1 \D_cache/cache_reg[2][142]  ( .D(\D_cache/n658 ), .CK(clk), .RN(n5802), .Q(\D_cache/cache[2][142] ), .QN(n2439) );
  DFFRX1 \D_cache/cache_reg[3][142]  ( .D(\D_cache/n657 ), .CK(clk), .RN(n5802), .Q(\D_cache/cache[3][142] ), .QN(n463) );
  DFFRX1 \D_cache/cache_reg[6][142]  ( .D(\D_cache/n654 ), .CK(clk), .RN(n5803), .Q(\D_cache/cache[6][142] ), .QN(n2356) );
  DFFRX1 \D_cache/cache_reg[7][142]  ( .D(\D_cache/n653 ), .CK(clk), .RN(n5803), .Q(\D_cache/cache[7][142] ), .QN(n360) );
  DFFRX1 \D_cache/cache_reg[0][144]  ( .D(\D_cache/n644 ), .CK(clk), .RN(n5804), .Q(\D_cache/cache[0][144] ), .QN(n1885) );
  DFFRX1 \D_cache/cache_reg[1][144]  ( .D(\D_cache/n643 ), .CK(clk), .RN(n5804), .Q(\D_cache/cache[1][144] ), .QN(n318) );
  DFFRX1 \D_cache/cache_reg[2][144]  ( .D(\D_cache/n642 ), .CK(clk), .RN(n5804), .Q(\D_cache/cache[2][144] ) );
  DFFRX1 \D_cache/cache_reg[3][144]  ( .D(\D_cache/n641 ), .CK(clk), .RN(n5804), .Q(\D_cache/cache[3][144] ), .QN(n1896) );
  DFFRX1 \D_cache/cache_reg[4][144]  ( .D(\D_cache/n640 ), .CK(clk), .RN(n5804), .Q(\D_cache/cache[4][144] ), .QN(n1886) );
  DFFRX1 \D_cache/cache_reg[5][144]  ( .D(\D_cache/n639 ), .CK(clk), .RN(n5804), .Q(\D_cache/cache[5][144] ), .QN(n319) );
  DFFRX1 \D_cache/cache_reg[6][144]  ( .D(\D_cache/n638 ), .CK(clk), .RN(n5804), .Q(\D_cache/cache[6][144] ), .QN(n1899) );
  DFFRX1 \D_cache/cache_reg[3][146]  ( .D(\D_cache/n625 ), .CK(clk), .RN(n5805), .Q(\D_cache/cache[3][146] ), .QN(n1888) );
  DFFRX1 \D_cache/cache_reg[6][146]  ( .D(\D_cache/n622 ), .CK(clk), .RN(n5805), .Q(\D_cache/cache[6][146] ), .QN(n1961) );
  DFFRX1 \D_cache/cache_reg[7][146]  ( .D(\D_cache/n621 ), .CK(clk), .RN(n5805), .Q(\D_cache/cache[7][146] ), .QN(n389) );
  DFFRX1 \D_cache/cache_reg[2][152]  ( .D(\D_cache/n578 ), .CK(clk), .RN(n5809), .Q(\D_cache/cache[2][152] ), .QN(n1954) );
  DFFRX1 \D_cache/cache_reg[3][152]  ( .D(\D_cache/n577 ), .CK(clk), .RN(n5809), .Q(\D_cache/cache[3][152] ), .QN(n378) );
  DFFRX1 \D_cache/cache_reg[6][152]  ( .D(\D_cache/n574 ), .CK(clk), .RN(n5809), .Q(\D_cache/cache[6][152] ), .QN(n453) );
  DFFRX1 \D_cache/cache_reg[7][152]  ( .D(\D_cache/n573 ), .CK(clk), .RN(n5809), .Q(\D_cache/cache[7][152] ), .QN(n2009) );
  DFFRX1 \I_cache/cache_reg[2][133]  ( .D(n11757), .CK(clk), .RN(n5900), .Q(
        \I_cache/cache[2][133] ), .QN(n1939) );
  DFFRX1 \D_cache/cache_reg[1][142]  ( .D(\D_cache/n659 ), .CK(clk), .RN(n5802), .Q(\D_cache/cache[1][142] ), .QN(n1881) );
  DFFRX1 \I_cache/cache_reg[6][128]  ( .D(n11793), .CK(clk), .RN(n5897), .Q(
        \I_cache/cache[6][128] ), .QN(n1970) );
  DFFRX1 \I_cache/cache_reg[2][134]  ( .D(n11749), .CK(clk), .RN(n5900), .Q(
        \I_cache/cache[2][134] ), .QN(n1985) );
  DFFRX1 \I_cache/cache_reg[1][128]  ( .D(n11798), .CK(clk), .RN(n5896), .Q(
        \I_cache/cache[1][128] ), .QN(n399) );
  DFFRX1 \I_cache/cache_reg[5][130]  ( .D(n11778), .CK(clk), .RN(n5898), .Q(
        \I_cache/cache[5][130] ), .QN(n1624) );
  DFFRX1 \I_cache/cache_reg[4][146]  ( .D(n11651), .CK(clk), .RN(n5909), .Q(
        \I_cache/cache[4][146] ), .QN(n1950) );
  DFFRX1 \I_cache/cache_reg[2][145]  ( .D(n11661), .CK(clk), .RN(n5908), .Q(
        \I_cache/cache[2][145] ), .QN(n1949) );
  DFFRX1 \I_cache/cache_reg[4][150]  ( .D(n11619), .CK(clk), .RN(n5911), .Q(
        \I_cache/cache[4][150] ), .QN(n3286) );
  DFFRX1 \I_cache/cache_reg[3][129]  ( .D(n11788), .CK(clk), .RN(n5897), .Q(
        \I_cache/cache[3][129] ), .QN(n1618) );
  DFFRX1 \I_cache/cache_reg[6][139]  ( .D(n11705), .CK(clk), .RN(n5904), .Q(
        \I_cache/cache[6][139] ), .QN(n1897) );
  DFFRX1 \I_cache/cache_reg[0][130]  ( .D(n11783), .CK(clk), .RN(n5898), .Q(
        \I_cache/cache[0][130] ), .QN(n1976) );
  DFFRX1 \I_cache/cache_reg[2][138]  ( .D(n11717), .CK(clk), .RN(n5903), .Q(
        \I_cache/cache[2][138] ), .QN(n1953) );
  DFFRX1 \I_cache/cache_reg[7][131]  ( .D(n11768), .CK(clk), .RN(n5899), .Q(
        \I_cache/cache[7][131] ), .QN(n2026) );
  DFFRX1 \I_cache/cache_reg[0][148]  ( .D(n11639), .CK(clk), .RN(n5910), .Q(
        \I_cache/cache[0][148] ), .QN(n1968) );
  DFFRX1 \I_cache/cache_reg[1][139]  ( .D(n11710), .CK(clk), .RN(n5904), .Q(
        \I_cache/cache[1][139] ), .QN(n404) );
  DFFRX1 \I_cache/cache_reg[2][130]  ( .D(n11781), .CK(clk), .RN(n5898), .Q(
        \I_cache/cache[2][130] ), .QN(n1977) );
  DFFRX1 \I_cache/cache_reg[5][150]  ( .D(n11618), .CK(clk), .RN(n5911), .Q(
        \I_cache/cache[5][150] ), .QN(n1626) );
  DFFRX1 \I_cache/cache_reg[5][134]  ( .D(n11746), .CK(clk), .RN(n5901), .Q(
        \I_cache/cache[5][134] ), .QN(n1619) );
  DFFRX1 \I_cache/cache_reg[2][146]  ( .D(n11653), .CK(clk), .RN(n5908), .Q(
        \I_cache/cache[2][146] ), .QN(n1982) );
  DFFRX1 \I_cache/cache_reg[5][128]  ( .D(n11794), .CK(clk), .RN(n5897), .Q(
        \I_cache/cache[5][128] ), .QN(n1625) );
  DFFRX1 \I_cache/cache_reg[1][133]  ( .D(n11758), .CK(clk), .RN(n5900), .Q(
        \I_cache/cache[1][133] ), .QN(n376) );
  DFFRX1 \I_cache/cache_reg[4][148]  ( .D(n11635), .CK(clk), .RN(n5910), .Q(
        \I_cache/cache[4][148] ) );
  DFFRX1 \I_cache/cache_reg[6][130]  ( .D(n11777), .CK(clk), .RN(n5898), .Q(
        \I_cache/cache[6][130] ), .QN(n1978) );
  DFFRX1 \I_cache/cache_reg[1][130]  ( .D(n11782), .CK(clk), .RN(n5898), .Q(
        \I_cache/cache[1][130] ), .QN(n409) );
  DFFRX1 \I_cache/cache_reg[7][132]  ( .D(n11760), .CK(clk), .RN(n5899), .Q(
        \I_cache/cache[7][132] ), .QN(n1876) );
  DFFRX1 \I_cache/cache_reg[4][145]  ( .D(n11659), .CK(clk), .RN(n5908), .Q(
        \I_cache/cache[4][145] ), .QN(n1966) );
  DFFRX1 \I_cache/cache_reg[4][144]  ( .D(n11667), .CK(clk), .RN(n5907), .Q(
        \I_cache/cache[4][144] ) );
  DFFRX1 \I_cache/cache_reg[6][134]  ( .D(n11745), .CK(clk), .RN(n5901), .Q(
        \I_cache/cache[6][134] ), .QN(n1986) );
  DFFRX1 \I_cache/cache_reg[3][130]  ( .D(n11780), .CK(clk), .RN(n5898), .Q(
        \I_cache/cache[3][130] ), .QN(n410) );
  DFFRX1 \I_cache/cache_reg[0][150]  ( .D(n11623), .CK(clk), .RN(n5911), .Q(
        \I_cache/cache[0][150] ), .QN(n1979) );
  DFFRX1 \I_cache/cache_reg[1][134]  ( .D(n11750), .CK(clk), .RN(n5900), .Q(
        \I_cache/cache[1][134] ), .QN(n417) );
  DFFRX1 \I_cache/cache_reg[0][144]  ( .D(n11671), .CK(clk), .RN(n5907), .Q(
        \I_cache/cache[0][144] ), .QN(n1972) );
  DFFRX1 \I_cache/cache_reg[3][128]  ( .D(n11796), .CK(clk), .RN(n5897), .Q(
        \I_cache/cache[3][128] ), .QN(n400) );
  DFFRX1 \I_cache/cache_reg[1][138]  ( .D(n11718), .CK(clk), .RN(n5903), .Q(
        \I_cache/cache[1][138] ), .QN(n375) );
  DFFRX1 \I_cache/cache_reg[5][139]  ( .D(n11706), .CK(clk), .RN(n5904), .Q(
        \I_cache/cache[5][139] ), .QN(n3215) );
  DFFRX1 \I_cache/cache_reg[4][133]  ( .D(n11755), .CK(clk), .RN(n5900), .Q(
        \I_cache/cache[4][133] ), .QN(n3278) );
  DFFRX1 \I_cache/cache_reg[2][150]  ( .D(n11621), .CK(clk), .RN(n5911), .Q(
        \I_cache/cache[2][150] ), .QN(n1941) );
  DFFRX1 \I_cache/cache_reg[7][151]  ( .D(n11608), .CK(clk), .RN(n5912), .Q(
        \I_cache/cache[7][151] ), .QN(n408) );
  DFFRX1 \I_cache/cache_reg[3][133]  ( .D(n11756), .CK(clk), .RN(n5900), .Q(
        \I_cache/cache[3][133] ), .QN(n361) );
  DFFRX1 \I_cache/cache_reg[4][138]  ( .D(n11715), .CK(clk), .RN(n5903), .Q(
        \I_cache/cache[4][138] ), .QN(n3279) );
  DFFRX1 \I_cache/cache_reg[2][148]  ( .D(n11637), .CK(clk), .RN(n5910), .Q(
        \I_cache/cache[2][148] ), .QN(n1969) );
  DFFRX1 \I_cache/cache_reg[6][145]  ( .D(n11657), .CK(clk), .RN(n5908), .Q(
        \I_cache/cache[6][145] ), .QN(n1942) );
  DFFRX1 \I_cache/cache_reg[7][130]  ( .D(n11776), .CK(clk), .RN(n5898), .Q(
        \I_cache/cache[7][130] ), .QN(n411) );
  DFFRX1 \I_cache/cache_reg[6][150]  ( .D(n11617), .CK(clk), .RN(n5911), .Q(
        \I_cache/cache[6][150] ), .QN(n1980) );
  DFFRX1 \I_cache/cache_reg[1][150]  ( .D(n11622), .CK(clk), .RN(n5911), .Q(
        \I_cache/cache[1][150] ), .QN(n412) );
  DFFRX1 \I_cache/cache_reg[0][145]  ( .D(n11663), .CK(clk), .RN(n5908), .Q(
        \I_cache/cache[0][145] ), .QN(n3276) );
  DFFRX1 \I_cache/cache_reg[3][138]  ( .D(n11716), .CK(clk), .RN(n5903), .Q(
        \I_cache/cache[3][138] ), .QN(n377) );
  DFFRX1 \I_cache/cache_reg[3][134]  ( .D(n11748), .CK(clk), .RN(n5900), .Q(
        \I_cache/cache[3][134] ), .QN(n418) );
  DFFRX1 \I_cache/cache_reg[5][146]  ( .D(n11650), .CK(clk), .RN(n5909), .Q(
        \I_cache/cache[5][146] ), .QN(n372) );
  DFFRX1 \I_cache/cache_reg[3][139]  ( .D(n11708), .CK(clk), .RN(n5904), .Q(
        \I_cache/cache[3][139] ), .QN(n405) );
  DFFRX1 \I_cache/cache_reg[3][150]  ( .D(n11620), .CK(clk), .RN(n5911), .Q(
        \I_cache/cache[3][150] ), .QN(n363) );
  DFFRX1 \I_cache/cache_reg[2][144]  ( .D(n11669), .CK(clk), .RN(n5907), .Q(
        \I_cache/cache[2][144] ), .QN(n1973) );
  DFFRX1 \I_cache/cache_reg[4][137]  ( .D(n11723), .CK(clk), .RN(n5903), .Q(
        \I_cache/cache[4][137] ) );
  DFFRX1 \I_cache/cache_reg[6][146]  ( .D(n11649), .CK(clk), .RN(n5909), .Q(
        \I_cache/cache[6][146] ), .QN(n1983) );
  DFFRX1 \I_cache/cache_reg[1][146]  ( .D(n11654), .CK(clk), .RN(n5908), .Q(
        \I_cache/cache[1][146] ), .QN(n414) );
  DFFRX1 \I_cache/cache_reg[7][150]  ( .D(n11616), .CK(clk), .RN(n5911), .Q(
        \I_cache/cache[7][150] ), .QN(n413) );
  DFFRX1 \I_cache/cache_reg[5][133]  ( .D(n11754), .CK(clk), .RN(n5900), .Q(
        \I_cache/cache[5][133] ), .QN(n1622) );
  DFFRX1 \I_cache/cache_reg[3][145]  ( .D(n11660), .CK(clk), .RN(n5908), .Q(
        \I_cache/cache[3][145] ), .QN(n371) );
  DFFRX1 \I_cache/cache_reg[5][138]  ( .D(n11714), .CK(clk), .RN(n5903), .Q(
        \I_cache/cache[5][138] ), .QN(n1623) );
  DFFRX1 \I_cache/cache_reg[0][137]  ( .D(n11727), .CK(clk), .RN(n5902), .Q(
        \I_cache/cache[0][137] ), .QN(n1971) );
  DFFRX1 \I_cache/cache_reg[4][135]  ( .D(n11739), .CK(clk), .RN(n5901), .Q(
        \I_cache/cache[4][135] ) );
  DFFRX1 \I_cache/cache_reg[7][134]  ( .D(n11744), .CK(clk), .RN(n5901), .Q(
        \I_cache/cache[7][134] ), .QN(n419) );
  DFFRX1 \I_cache/cache_reg[5][144]  ( .D(n11666), .CK(clk), .RN(n5907), .Q(
        \I_cache/cache[5][144] ), .QN(n3214) );
  DFFRX1 \I_cache/cache_reg[7][128]  ( .D(n11792), .CK(clk), .RN(n5914), .Q(
        \I_cache/cache[7][128] ), .QN(n398) );
  DFFRX1 \I_cache/cache_reg[5][148]  ( .D(n11634), .CK(clk), .RN(n5910), .Q(
        \I_cache/cache[5][148] ), .QN(n3211) );
  DFFRX1 \I_cache/cache_reg[4][140]  ( .D(n11699), .CK(clk), .RN(n5905), .Q(
        \I_cache/cache[4][140] ) );
  DFFRX1 \I_cache/cache_reg[6][148]  ( .D(n11633), .CK(clk), .RN(n5910), .Q(
        \I_cache/cache[6][148] ), .QN(n425) );
  DFFRX1 \I_cache/cache_reg[3][146]  ( .D(n11652), .CK(clk), .RN(n5908), .Q(
        \I_cache/cache[3][146] ), .QN(n415) );
  DFFRX1 \I_cache/cache_reg[5][145]  ( .D(n11658), .CK(clk), .RN(n5908), .Q(
        \I_cache/cache[5][145] ), .QN(n394) );
  DFFRX1 \I_cache/cache_reg[2][137]  ( .D(n11725), .CK(clk), .RN(n5902), .Q(
        \I_cache/cache[2][137] ), .QN(n426) );
  DFFRX1 \I_cache/cache_reg[1][145]  ( .D(n11662), .CK(clk), .RN(n5908), .Q(
        \I_cache/cache[1][145] ), .QN(n1620) );
  DFFRX1 \I_cache/cache_reg[6][144]  ( .D(n11665), .CK(clk), .RN(n5907), .Q(
        \I_cache/cache[6][144] ), .QN(n427) );
  DFFRX1 \I_cache/cache_reg[0][142]  ( .D(n11687), .CK(clk), .RN(n5906), .Q(
        \I_cache/cache[0][142] ), .QN(n455) );
  DFFRX1 \I_cache/cache_reg[4][143]  ( .D(n11675), .CK(clk), .RN(n5907), .Q(
        \I_cache/cache[4][143] ), .QN(n3277) );
  DFFRX1 \I_cache/cache_reg[1][144]  ( .D(n11670), .CK(clk), .RN(n5907), .Q(
        \I_cache/cache[1][144] ), .QN(n402) );
  DFFRX1 \I_cache/cache_reg[4][136]  ( .D(n11731), .CK(clk), .RN(n5902), .Q(
        \I_cache/cache[4][136] ), .QN(n1630) );
  DFFRX1 \I_cache/cache_reg[0][135]  ( .D(n11743), .CK(clk), .RN(n5901), .Q(
        \I_cache/cache[0][135] ), .QN(n3283) );
  DFFRX1 \I_cache/cache_reg[0][140]  ( .D(n11703), .CK(clk), .RN(n5904), .Q(
        \I_cache/cache[0][140] ), .QN(n3281) );
  DFFRX1 \I_cache/cache_reg[4][132]  ( .D(n11763), .CK(clk), .RN(n5899), .Q(
        \I_cache/cache[4][132] ), .QN(n3222) );
  DFFRX1 \I_cache/cache_reg[4][147]  ( .D(n11643), .CK(clk), .RN(n5909), .Q(
        \I_cache/cache[4][147] ) );
  DFFRX1 \I_cache/cache_reg[3][144]  ( .D(n11668), .CK(clk), .RN(n5907), .Q(
        \I_cache/cache[3][144] ), .QN(n403) );
  DFFRX1 \I_cache/cache_reg[2][135]  ( .D(n11741), .CK(clk), .RN(n5901), .Q(
        \I_cache/cache[2][135] ), .QN(n3284) );
  DFFRX1 \I_cache/cache_reg[7][146]  ( .D(n11648), .CK(clk), .RN(n5909), .Q(
        \I_cache/cache[7][146] ), .QN(n416) );
  DFFRX1 \I_cache/cache_reg[2][140]  ( .D(n11701), .CK(clk), .RN(n5904), .Q(
        \I_cache/cache[2][140] ), .QN(n3282) );
  DFFRX1 \I_cache/cache_reg[2][142]  ( .D(n11685), .CK(clk), .RN(n5906), .Q(
        \I_cache/cache[2][142] ), .QN(n448) );
  DFFRX1 \I_cache/cache_reg[6][137]  ( .D(n11721), .CK(clk), .RN(n5903), .Q(
        \I_cache/cache[6][137] ), .QN(n428) );
  DFFRX1 \I_cache/cache_reg[5][136]  ( .D(n11730), .CK(clk), .RN(n5902), .Q(
        \I_cache/cache[5][136] ), .QN(n3293) );
  DFFRX1 \I_cache/cache_reg[1][137]  ( .D(n11726), .CK(clk), .RN(n5902), .Q(
        \I_cache/cache[1][137] ), .QN(n401) );
  DFFRX1 \I_cache/cache_reg[0][143]  ( .D(n11679), .CK(clk), .RN(n5906), .Q(
        \I_cache/cache[0][143] ), .QN(n456) );
  DFFRX1 \I_cache/cache_reg[0][136]  ( .D(n11735), .CK(clk), .RN(n5902), .Q(
        \I_cache/cache[0][136] ), .QN(n420) );
  DFFRX1 \i_MIPS/EX_MEM_reg[3]  ( .D(\i_MIPS/n524 ), .CK(clk), .RN(n5616), .Q(
        DCACHE_ren), .QN(\i_MIPS/n334 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[103]  ( .D(\i_MIPS/n482 ), .CK(clk), .RN(n5610), 
        .Q(\i_MIPS/ID_EX[103] ), .QN(n4639) );
  DFFRX1 \i_MIPS/ID_EX_reg[99]  ( .D(\i_MIPS/n486 ), .CK(clk), .RN(n5610), .Q(
        \i_MIPS/ID_EX[99] ), .QN(n4493) );
  DFFRX1 \i_MIPS/ID_EX_reg[96]  ( .D(\i_MIPS/n489 ), .CK(clk), .RN(n5611), .Q(
        \i_MIPS/ID_EX[96] ), .QN(n4649) );
  DFFRX1 \i_MIPS/ID_EX_reg[98]  ( .D(\i_MIPS/n487 ), .CK(clk), .RN(n5610), .Q(
        \i_MIPS/ID_EX[98] ), .QN(n4650) );
  DFFRX1 \i_MIPS/ID_EX_reg[94]  ( .D(\i_MIPS/n491 ), .CK(clk), .RN(n5611), .Q(
        \i_MIPS/ID_EX[94] ), .QN(n4647) );
  DFFRX1 \i_MIPS/ID_EX_reg[92]  ( .D(\i_MIPS/n493 ), .CK(clk), .RN(n5611), .Q(
        \i_MIPS/ID_EX[92] ), .QN(n4645) );
  DFFRX1 \i_MIPS/Register/register_reg[30][2]  ( .D(\i_MIPS/Register/n150 ), 
        .CK(clk), .RN(n5625), .Q(\i_MIPS/Register/register[30][2] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][3]  ( .D(\i_MIPS/Register/n151 ), 
        .CK(clk), .RN(n5625), .Q(\i_MIPS/Register/register[30][3] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][6]  ( .D(\i_MIPS/Register/n154 ), 
        .CK(clk), .RN(n5625), .Q(\i_MIPS/Register/register[30][6] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][7]  ( .D(\i_MIPS/Register/n155 ), 
        .CK(clk), .RN(n5626), .Q(\i_MIPS/Register/register[30][7] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][9]  ( .D(\i_MIPS/Register/n157 ), 
        .CK(clk), .RN(n5626), .Q(\i_MIPS/Register/register[30][9] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][13]  ( .D(\i_MIPS/Register/n161 ), 
        .CK(clk), .RN(n5626), .Q(\i_MIPS/Register/register[30][13] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][14]  ( .D(\i_MIPS/Register/n162 ), 
        .CK(clk), .RN(n5626), .Q(\i_MIPS/Register/register[30][14] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][16]  ( .D(\i_MIPS/Register/n164 ), 
        .CK(clk), .RN(n5626), .Q(\i_MIPS/Register/register[30][16] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][20]  ( .D(\i_MIPS/Register/n168 ), 
        .CK(clk), .RN(n5627), .Q(\i_MIPS/Register/register[30][20] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][21]  ( .D(\i_MIPS/Register/n169 ), 
        .CK(clk), .RN(n5627), .Q(\i_MIPS/Register/register[30][21] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][22]  ( .D(\i_MIPS/Register/n170 ), 
        .CK(clk), .RN(n5627), .Q(\i_MIPS/Register/register[30][22] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][23]  ( .D(\i_MIPS/Register/n171 ), 
        .CK(clk), .RN(n5627), .Q(\i_MIPS/Register/register[30][23] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][24]  ( .D(\i_MIPS/Register/n172 ), 
        .CK(clk), .RN(n5627), .Q(\i_MIPS/Register/register[30][24] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][25]  ( .D(\i_MIPS/Register/n173 ), 
        .CK(clk), .RN(n5627), .Q(\i_MIPS/Register/register[30][25] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][27]  ( .D(\i_MIPS/Register/n175 ), 
        .CK(clk), .RN(n5627), .Q(\i_MIPS/Register/register[30][27] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][28]  ( .D(\i_MIPS/Register/n176 ), 
        .CK(clk), .RN(n5627), .Q(\i_MIPS/Register/register[30][28] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][2]  ( .D(\i_MIPS/Register/n662 ), 
        .CK(clk), .RN(n5668), .Q(\i_MIPS/Register/register[14][2] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][3]  ( .D(\i_MIPS/Register/n663 ), 
        .CK(clk), .RN(n5668), .Q(\i_MIPS/Register/register[14][3] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][6]  ( .D(\i_MIPS/Register/n666 ), 
        .CK(clk), .RN(n5668), .Q(\i_MIPS/Register/register[14][6] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][7]  ( .D(\i_MIPS/Register/n667 ), 
        .CK(clk), .RN(n5668), .Q(\i_MIPS/Register/register[14][7] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][13]  ( .D(\i_MIPS/Register/n673 ), 
        .CK(clk), .RN(n5669), .Q(\i_MIPS/Register/register[14][13] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][14]  ( .D(\i_MIPS/Register/n674 ), 
        .CK(clk), .RN(n5669), .Q(\i_MIPS/Register/register[14][14] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][16]  ( .D(\i_MIPS/Register/n676 ), 
        .CK(clk), .RN(n5669), .Q(\i_MIPS/Register/register[14][16] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][20]  ( .D(\i_MIPS/Register/n680 ), 
        .CK(clk), .RN(n5669), .Q(\i_MIPS/Register/register[14][20] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][21]  ( .D(\i_MIPS/Register/n681 ), 
        .CK(clk), .RN(n5669), .Q(\i_MIPS/Register/register[14][21] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][22]  ( .D(\i_MIPS/Register/n682 ), 
        .CK(clk), .RN(n5669), .Q(\i_MIPS/Register/register[14][22] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][23]  ( .D(\i_MIPS/Register/n683 ), 
        .CK(clk), .RN(n5670), .Q(\i_MIPS/Register/register[14][23] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][24]  ( .D(\i_MIPS/Register/n684 ), 
        .CK(clk), .RN(n5670), .Q(\i_MIPS/Register/register[14][24] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][25]  ( .D(\i_MIPS/Register/n685 ), 
        .CK(clk), .RN(n5670), .Q(\i_MIPS/Register/register[14][25] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][27]  ( .D(\i_MIPS/Register/n687 ), 
        .CK(clk), .RN(n5670), .Q(\i_MIPS/Register/register[14][27] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][28]  ( .D(\i_MIPS/Register/n688 ), 
        .CK(clk), .RN(n5670), .Q(\i_MIPS/Register/register[14][28] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][3]  ( .D(\i_MIPS/Register/n407 ), 
        .CK(clk), .RN(n5647), .Q(\i_MIPS/Register/register[22][3] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][16]  ( .D(\i_MIPS/Register/n420 ), 
        .CK(clk), .RN(n5648), .Q(\i_MIPS/Register/register[22][16] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][20]  ( .D(\i_MIPS/Register/n424 ), 
        .CK(clk), .RN(n5648), .Q(\i_MIPS/Register/register[22][20] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][22]  ( .D(\i_MIPS/Register/n426 ), 
        .CK(clk), .RN(n5648), .Q(\i_MIPS/Register/register[22][22] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][23]  ( .D(\i_MIPS/Register/n427 ), 
        .CK(clk), .RN(n5648), .Q(\i_MIPS/Register/register[22][23] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][24]  ( .D(\i_MIPS/Register/n428 ), 
        .CK(clk), .RN(n5648), .Q(\i_MIPS/Register/register[22][24] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][3]  ( .D(\i_MIPS/Register/n919 ), 
        .CK(clk), .RN(n5689), .Q(\i_MIPS/Register/register[6][3] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][16]  ( .D(\i_MIPS/Register/n932 ), 
        .CK(clk), .RN(n5690), .Q(\i_MIPS/Register/register[6][16] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][20]  ( .D(\i_MIPS/Register/n936 ), 
        .CK(clk), .RN(n5691), .Q(\i_MIPS/Register/register[6][20] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][22]  ( .D(\i_MIPS/Register/n938 ), 
        .CK(clk), .RN(n5691), .Q(\i_MIPS/Register/register[6][22] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][23]  ( .D(\i_MIPS/Register/n939 ), 
        .CK(clk), .RN(n5691), .Q(\i_MIPS/Register/register[6][23] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][24]  ( .D(\i_MIPS/Register/n940 ), 
        .CK(clk), .RN(n5691), .Q(\i_MIPS/Register/register[6][24] ) );
  DFFRX1 \i_MIPS/Register/register_reg[29][2]  ( .D(\i_MIPS/Register/n182 ), 
        .CK(clk), .RN(n5628), .Q(\i_MIPS/Register/register[29][2] ), .QN(n571)
         );
  DFFRX1 \i_MIPS/Register/register_reg[29][3]  ( .D(\i_MIPS/Register/n183 ), 
        .CK(clk), .RN(n5628), .Q(\i_MIPS/Register/register[29][3] ), .QN(n580)
         );
  DFFRX1 \i_MIPS/Register/register_reg[29][4]  ( .D(\i_MIPS/Register/n184 ), 
        .CK(clk), .RN(n5628), .Q(\i_MIPS/Register/register[29][4] ), .QN(n340)
         );
  DFFRX1 \i_MIPS/Register/register_reg[29][5]  ( .D(\i_MIPS/Register/n185 ), 
        .CK(clk), .RN(n5628), .Q(\i_MIPS/Register/register[29][5] ), .QN(n551)
         );
  DFFRX1 \i_MIPS/Register/register_reg[29][6]  ( .D(\i_MIPS/Register/n186 ), 
        .CK(clk), .RN(n5628), .Q(\i_MIPS/Register/register[29][6] ), .QN(n660)
         );
  DFFRX1 \i_MIPS/Register/register_reg[29][7]  ( .D(\i_MIPS/Register/n187 ), 
        .CK(clk), .RN(n5628), .Q(\i_MIPS/Register/register[29][7] ), .QN(n523)
         );
  DFFRX1 \i_MIPS/Register/register_reg[29][8]  ( .D(\i_MIPS/Register/n188 ), 
        .CK(clk), .RN(n5628), .Q(\i_MIPS/Register/register[29][8] ), .QN(n565)
         );
  DFFRX1 \i_MIPS/Register/register_reg[29][9]  ( .D(\i_MIPS/Register/n189 ), 
        .CK(clk), .RN(n5628), .Q(\i_MIPS/Register/register[29][9] ), .QN(n563)
         );
  DFFRX1 \i_MIPS/Register/register_reg[29][10]  ( .D(\i_MIPS/Register/n190 ), 
        .CK(clk), .RN(n5628), .Q(\i_MIPS/Register/register[29][10] ), .QN(n343) );
  DFFRX1 \i_MIPS/Register/register_reg[29][11]  ( .D(\i_MIPS/Register/n191 ), 
        .CK(clk), .RN(n5629), .Q(\i_MIPS/Register/register[29][11] ), .QN(n342) );
  DFFRX1 \i_MIPS/Register/register_reg[29][12]  ( .D(\i_MIPS/Register/n192 ), 
        .CK(clk), .RN(n5629), .Q(\i_MIPS/Register/register[29][12] ), .QN(n350) );
  DFFRX1 \i_MIPS/Register/register_reg[29][13]  ( .D(\i_MIPS/Register/n193 ), 
        .CK(clk), .RN(n5629), .Q(\i_MIPS/Register/register[29][13] ), .QN(n567) );
  DFFRX1 \i_MIPS/Register/register_reg[29][14]  ( .D(\i_MIPS/Register/n194 ), 
        .CK(clk), .RN(n5629), .Q(\i_MIPS/Register/register[29][14] ), .QN(n349) );
  DFFRX1 \i_MIPS/Register/register_reg[29][15]  ( .D(\i_MIPS/Register/n195 ), 
        .CK(clk), .RN(n5629), .Q(\i_MIPS/Register/register[29][15] ), .QN(n524) );
  DFFRX1 \i_MIPS/Register/register_reg[29][16]  ( .D(\i_MIPS/Register/n196 ), 
        .CK(clk), .RN(n5629), .Q(\i_MIPS/Register/register[29][16] ), .QN(n261) );
  DFFRX1 \i_MIPS/Register/register_reg[29][17]  ( .D(\i_MIPS/Register/n197 ), 
        .CK(clk), .RN(n5629), .Q(\i_MIPS/Register/register[29][17] ), .QN(n487) );
  DFFRX1 \i_MIPS/Register/register_reg[29][18]  ( .D(\i_MIPS/Register/n198 ), 
        .CK(clk), .RN(n5629), .Q(\i_MIPS/Register/register[29][18] ), .QN(n437) );
  DFFRX1 \i_MIPS/Register/register_reg[29][20]  ( .D(\i_MIPS/Register/n200 ), 
        .CK(clk), .RN(n5629), .Q(\i_MIPS/Register/register[29][20] ), .QN(n255) );
  DFFRX1 \i_MIPS/Register/register_reg[29][21]  ( .D(\i_MIPS/Register/n201 ), 
        .CK(clk), .RN(n5629), .Q(\i_MIPS/Register/register[29][21] ), .QN(n263) );
  DFFRX1 \i_MIPS/Register/register_reg[29][22]  ( .D(\i_MIPS/Register/n202 ), 
        .CK(clk), .RN(n5629), .Q(\i_MIPS/Register/register[29][22] ), .QN(n433) );
  DFFRX1 \i_MIPS/Register/register_reg[29][23]  ( .D(\i_MIPS/Register/n203 ), 
        .CK(clk), .RN(n5630), .Q(\i_MIPS/Register/register[29][23] ), .QN(n258) );
  DFFRX1 \i_MIPS/Register/register_reg[29][24]  ( .D(\i_MIPS/Register/n204 ), 
        .CK(clk), .RN(n5630), .Q(\i_MIPS/Register/register[29][24] ), .QN(n578) );
  DFFRX1 \i_MIPS/Register/register_reg[29][25]  ( .D(\i_MIPS/Register/n205 ), 
        .CK(clk), .RN(n5630), .Q(\i_MIPS/Register/register[29][25] ), .QN(n256) );
  DFFRX1 \i_MIPS/Register/register_reg[29][26]  ( .D(\i_MIPS/Register/n206 ), 
        .CK(clk), .RN(n5630), .Q(\i_MIPS/Register/register[29][26] ), .QN(n265) );
  DFFRX1 \i_MIPS/Register/register_reg[29][27]  ( .D(\i_MIPS/Register/n207 ), 
        .CK(clk), .RN(n5630), .Q(\i_MIPS/Register/register[29][27] ), .QN(n667) );
  DFFRX1 \i_MIPS/Register/register_reg[29][28]  ( .D(\i_MIPS/Register/n208 ), 
        .CK(clk), .RN(n5630), .Q(\i_MIPS/Register/register[29][28] ), .QN(n579) );
  DFFRX1 \i_MIPS/Register/register_reg[29][29]  ( .D(\i_MIPS/Register/n209 ), 
        .CK(clk), .RN(n5630), .Q(\i_MIPS/Register/register[29][29] ), .QN(n337) );
  DFFRX1 \i_MIPS/Register/register_reg[29][31]  ( .D(\i_MIPS/Register/n211 ), 
        .CK(clk), .RN(n5630), .Q(\i_MIPS/Register/register[29][31] ), .QN(n657) );
  DFFRX1 \i_MIPS/Register/register_reg[28][24]  ( .D(\i_MIPS/Register/n236 ), 
        .CK(clk), .RN(n5632), .Q(\i_MIPS/Register/register[28][24] ), .QN(n599) );
  DFFRX1 \i_MIPS/Register/register_reg[27][2]  ( .D(\i_MIPS/Register/n246 ), 
        .CK(clk), .RN(n5633), .Q(\i_MIPS/Register/register[27][2] ), .QN(n570)
         );
  DFFRX1 \i_MIPS/Register/register_reg[27][3]  ( .D(\i_MIPS/Register/n247 ), 
        .CK(clk), .RN(n5633), .Q(\i_MIPS/Register/register[27][3] ), .QN(n503)
         );
  DFFRX1 \i_MIPS/Register/register_reg[27][4]  ( .D(\i_MIPS/Register/n248 ), 
        .CK(clk), .RN(n5633), .Q(\i_MIPS/Register/register[27][4] ), .QN(n588)
         );
  DFFRX1 \i_MIPS/Register/register_reg[27][5]  ( .D(\i_MIPS/Register/n249 ), 
        .CK(clk), .RN(n5633), .Q(\i_MIPS/Register/register[27][5] ), .QN(n514)
         );
  DFFRX1 \i_MIPS/Register/register_reg[27][6]  ( .D(\i_MIPS/Register/n250 ), 
        .CK(clk), .RN(n5633), .Q(\i_MIPS/Register/register[27][6] ), .QN(n527)
         );
  DFFRX1 \i_MIPS/Register/register_reg[27][7]  ( .D(\i_MIPS/Register/n251 ), 
        .CK(clk), .RN(n5634), .Q(\i_MIPS/Register/register[27][7] ), .QN(n531)
         );
  DFFRX1 \i_MIPS/Register/register_reg[27][9]  ( .D(\i_MIPS/Register/n253 ), 
        .CK(clk), .RN(n5634), .Q(\i_MIPS/Register/register[27][9] ), .QN(n556)
         );
  DFFRX1 \i_MIPS/Register/register_reg[27][10]  ( .D(\i_MIPS/Register/n254 ), 
        .CK(clk), .RN(n5634), .Q(\i_MIPS/Register/register[27][10] ), .QN(n506) );
  DFFRX1 \i_MIPS/Register/register_reg[27][11]  ( .D(\i_MIPS/Register/n255 ), 
        .CK(clk), .RN(n5634), .Q(\i_MIPS/Register/register[27][11] ), .QN(n490) );
  DFFRX1 \i_MIPS/Register/register_reg[27][12]  ( .D(\i_MIPS/Register/n256 ), 
        .CK(clk), .RN(n5634), .Q(\i_MIPS/Register/register[27][12] ), .QN(n535) );
  DFFRX1 \i_MIPS/Register/register_reg[27][13]  ( .D(\i_MIPS/Register/n257 ), 
        .CK(clk), .RN(n5634), .Q(\i_MIPS/Register/register[27][13] ), .QN(n554) );
  DFFRX1 \i_MIPS/Register/register_reg[27][14]  ( .D(\i_MIPS/Register/n258 ), 
        .CK(clk), .RN(n5634), .Q(\i_MIPS/Register/register[27][14] ), .QN(n649) );
  DFFRX1 \i_MIPS/Register/register_reg[27][16]  ( .D(\i_MIPS/Register/n260 ), 
        .CK(clk), .RN(n5634), .Q(\i_MIPS/Register/register[27][16] ), .QN(n505) );
  DFFRX1 \i_MIPS/Register/register_reg[27][18]  ( .D(\i_MIPS/Register/n262 ), 
        .CK(clk), .RN(n5634), .Q(\i_MIPS/Register/register[27][18] ), .QN(n533) );
  DFFRX1 \i_MIPS/Register/register_reg[27][20]  ( .D(\i_MIPS/Register/n264 ), 
        .CK(clk), .RN(n5635), .Q(\i_MIPS/Register/register[27][20] ), .QN(n557) );
  DFFRX1 \i_MIPS/Register/register_reg[27][21]  ( .D(\i_MIPS/Register/n265 ), 
        .CK(clk), .RN(n5635), .Q(\i_MIPS/Register/register[27][21] ), .QN(n529) );
  DFFRX1 \i_MIPS/Register/register_reg[27][22]  ( .D(\i_MIPS/Register/n266 ), 
        .CK(clk), .RN(n5635), .Q(\i_MIPS/Register/register[27][22] ), .QN(n587) );
  DFFRX1 \i_MIPS/Register/register_reg[27][23]  ( .D(\i_MIPS/Register/n267 ), 
        .CK(clk), .RN(n5635), .Q(\i_MIPS/Register/register[27][23] ), .QN(n501) );
  DFFRX1 \i_MIPS/Register/register_reg[27][24]  ( .D(\i_MIPS/Register/n268 ), 
        .CK(clk), .RN(n5635), .Q(\i_MIPS/Register/register[27][24] ), .QN(n539) );
  DFFRX1 \i_MIPS/Register/register_reg[27][25]  ( .D(\i_MIPS/Register/n269 ), 
        .CK(clk), .RN(n5635), .Q(\i_MIPS/Register/register[27][25] ), .QN(n497) );
  DFFRX1 \i_MIPS/Register/register_reg[27][26]  ( .D(\i_MIPS/Register/n270 ), 
        .CK(clk), .RN(n5635), .Q(\i_MIPS/Register/register[27][26] ), .QN(n590) );
  DFFRX1 \i_MIPS/Register/register_reg[27][27]  ( .D(\i_MIPS/Register/n271 ), 
        .CK(clk), .RN(n5635), .Q(\i_MIPS/Register/register[27][27] ), .QN(n647) );
  DFFRX1 \i_MIPS/Register/register_reg[27][28]  ( .D(\i_MIPS/Register/n272 ), 
        .CK(clk), .RN(n5635), .Q(\i_MIPS/Register/register[27][28] ), .QN(n486) );
  DFFRX1 \i_MIPS/Register/register_reg[27][29]  ( .D(\i_MIPS/Register/n273 ), 
        .CK(clk), .RN(n5635), .Q(\i_MIPS/Register/register[27][29] ), .QN(n351) );
  DFFRX1 \i_MIPS/Register/register_reg[25][2]  ( .D(\i_MIPS/Register/n310 ), 
        .CK(clk), .RN(n5638), .Q(\i_MIPS/Register/register[25][2] ), .QN(n480)
         );
  DFFRX1 \i_MIPS/Register/register_reg[25][3]  ( .D(\i_MIPS/Register/n311 ), 
        .CK(clk), .RN(n5639), .Q(\i_MIPS/Register/register[25][3] ), .QN(n653)
         );
  DFFRX1 \i_MIPS/Register/register_reg[25][4]  ( .D(\i_MIPS/Register/n312 ), 
        .CK(clk), .RN(n5639), .Q(\i_MIPS/Register/register[25][4] ), .QN(n482)
         );
  DFFRX1 \i_MIPS/Register/register_reg[25][5]  ( .D(\i_MIPS/Register/n313 ), 
        .CK(clk), .RN(n5639), .Q(\i_MIPS/Register/register[25][5] ), .QN(n655)
         );
  DFFRX1 \i_MIPS/Register/register_reg[25][6]  ( .D(\i_MIPS/Register/n314 ), 
        .CK(clk), .RN(n5639), .Q(\i_MIPS/Register/register[25][6] ), .QN(n515)
         );
  DFFRX1 \i_MIPS/Register/register_reg[25][7]  ( .D(\i_MIPS/Register/n315 ), 
        .CK(clk), .RN(n5639), .Q(\i_MIPS/Register/register[25][7] ), .QN(n520)
         );
  DFFRX1 \i_MIPS/Register/register_reg[25][8]  ( .D(\i_MIPS/Register/n316 ), 
        .CK(clk), .RN(n5639), .Q(\i_MIPS/Register/register[25][8] ), .QN(n212)
         );
  DFFRX1 \i_MIPS/Register/register_reg[25][9]  ( .D(\i_MIPS/Register/n317 ), 
        .CK(clk), .RN(n5639), .Q(\i_MIPS/Register/register[25][9] ), .QN(n210)
         );
  DFFRX1 \i_MIPS/Register/register_reg[25][10]  ( .D(\i_MIPS/Register/n318 ), 
        .CK(clk), .RN(n5639), .Q(\i_MIPS/Register/register[25][10] ), .QN(n491) );
  DFFRX1 \i_MIPS/Register/register_reg[25][11]  ( .D(\i_MIPS/Register/n319 ), 
        .CK(clk), .RN(n5639), .Q(\i_MIPS/Register/register[25][11] ), .QN(n519) );
  DFFRX1 \i_MIPS/Register/register_reg[25][12]  ( .D(\i_MIPS/Register/n320 ), 
        .CK(clk), .RN(n5639), .Q(\i_MIPS/Register/register[25][12] ), .QN(n208) );
  DFFRX1 \i_MIPS/Register/register_reg[25][13]  ( .D(\i_MIPS/Register/n321 ), 
        .CK(clk), .RN(n5639), .Q(\i_MIPS/Register/register[25][13] ), .QN(n206) );
  DFFRX1 \i_MIPS/Register/register_reg[25][14]  ( .D(\i_MIPS/Register/n322 ), 
        .CK(clk), .RN(n5639), .Q(\i_MIPS/Register/register[25][14] ), .QN(n218) );
  DFFRX1 \i_MIPS/Register/register_reg[25][15]  ( .D(\i_MIPS/Register/n323 ), 
        .CK(clk), .RN(n5640), .Q(\i_MIPS/Register/register[25][15] ), .QN(n517) );
  DFFRX1 \i_MIPS/Register/register_reg[25][16]  ( .D(\i_MIPS/Register/n324 ), 
        .CK(clk), .RN(n5640), .Q(\i_MIPS/Register/register[25][16] ), .QN(n511) );
  DFFRX1 \i_MIPS/Register/register_reg[25][17]  ( .D(\i_MIPS/Register/n325 ), 
        .CK(clk), .RN(n5640), .Q(\i_MIPS/Register/register[25][17] ), .QN(n348) );
  DFFRX1 \i_MIPS/Register/register_reg[25][18]  ( .D(\i_MIPS/Register/n326 ), 
        .CK(clk), .RN(n5640), .Q(\i_MIPS/Register/register[25][18] ), .QN(n347) );
  DFFRX1 \i_MIPS/Register/register_reg[25][20]  ( .D(\i_MIPS/Register/n328 ), 
        .CK(clk), .RN(n5640), .Q(\i_MIPS/Register/register[25][20] ), .QN(n550) );
  DFFRX1 \i_MIPS/Register/register_reg[25][21]  ( .D(\i_MIPS/Register/n329 ), 
        .CK(clk), .RN(n5640), .Q(\i_MIPS/Register/register[25][21] ), .QN(n545) );
  DFFRX1 \i_MIPS/Register/register_reg[25][22]  ( .D(\i_MIPS/Register/n330 ), 
        .CK(clk), .RN(n5640), .Q(\i_MIPS/Register/register[25][22] ), .QN(n334) );
  DFFRX1 \i_MIPS/Register/register_reg[25][23]  ( .D(\i_MIPS/Register/n331 ), 
        .CK(clk), .RN(n5640), .Q(\i_MIPS/Register/register[25][23] ), .QN(n549) );
  DFFRX1 \i_MIPS/Register/register_reg[25][24]  ( .D(\i_MIPS/Register/n332 ), 
        .CK(clk), .RN(n5640), .Q(\i_MIPS/Register/register[25][24] ), .QN(n560) );
  DFFRX1 \i_MIPS/Register/register_reg[25][25]  ( .D(\i_MIPS/Register/n333 ), 
        .CK(clk), .RN(n5640), .Q(\i_MIPS/Register/register[25][25] ), .QN(n547) );
  DFFRX1 \i_MIPS/Register/register_reg[25][26]  ( .D(\i_MIPS/Register/n334 ), 
        .CK(clk), .RN(n5640), .Q(\i_MIPS/Register/register[25][26] ), .QN(n483) );
  DFFRX1 \i_MIPS/Register/register_reg[25][27]  ( .D(\i_MIPS/Register/n335 ), 
        .CK(clk), .RN(n5641), .Q(\i_MIPS/Register/register[25][27] ), .QN(n652) );
  DFFRX1 \i_MIPS/Register/register_reg[25][28]  ( .D(\i_MIPS/Register/n336 ), 
        .CK(clk), .RN(n5641), .Q(\i_MIPS/Register/register[25][28] ), .QN(n485) );
  DFFRX1 \i_MIPS/Register/register_reg[25][29]  ( .D(\i_MIPS/Register/n337 ), 
        .CK(clk), .RN(n5641), .Q(\i_MIPS/Register/register[25][29] ), .QN(n217) );
  DFFRX1 \i_MIPS/Register/register_reg[25][31]  ( .D(\i_MIPS/Register/n339 ), 
        .CK(clk), .RN(n5641), .Q(\i_MIPS/Register/register[25][31] ), .QN(n650) );
  DFFRX1 \i_MIPS/Register/register_reg[24][3]  ( .D(\i_MIPS/Register/n343 ), 
        .CK(clk), .RN(n5641), .Q(\i_MIPS/Register/register[24][3] ), .QN(n620)
         );
  DFFRX1 \i_MIPS/Register/register_reg[24][24]  ( .D(\i_MIPS/Register/n364 ), 
        .CK(clk), .RN(n5643), .Q(\i_MIPS/Register/register[24][24] ), .QN(n612) );
  DFFRX1 \i_MIPS/Register/register_reg[15][2]  ( .D(\i_MIPS/Register/n630 ), 
        .CK(clk), .RN(n5665), .Q(\i_MIPS/Register/register[15][2] ), .QN(n572)
         );
  DFFRX1 \i_MIPS/Register/register_reg[15][3]  ( .D(\i_MIPS/Register/n631 ), 
        .CK(clk), .RN(n5665), .Q(\i_MIPS/Register/register[15][3] ), .QN(n585)
         );
  DFFRX1 \i_MIPS/Register/register_reg[15][4]  ( .D(\i_MIPS/Register/n632 ), 
        .CK(clk), .RN(n5665), .Q(\i_MIPS/Register/register[15][4] ), .QN(n339)
         );
  DFFRX1 \i_MIPS/Register/register_reg[15][5]  ( .D(\i_MIPS/Register/n633 ), 
        .CK(clk), .RN(n5665), .Q(\i_MIPS/Register/register[15][5] ), .QN(n669)
         );
  DFFRX1 \i_MIPS/Register/register_reg[15][6]  ( .D(\i_MIPS/Register/n634 ), 
        .CK(clk), .RN(n5665), .Q(\i_MIPS/Register/register[15][6] ), .QN(n220)
         );
  DFFRX1 \i_MIPS/Register/register_reg[15][7]  ( .D(\i_MIPS/Register/n635 ), 
        .CK(clk), .RN(n5666), .Q(\i_MIPS/Register/register[15][7] ), .QN(n664)
         );
  DFFRX1 \i_MIPS/Register/register_reg[15][10]  ( .D(\i_MIPS/Register/n638 ), 
        .CK(clk), .RN(n5666), .Q(\i_MIPS/Register/register[15][10] ), .QN(n288) );
  DFFRX1 \i_MIPS/Register/register_reg[15][11]  ( .D(\i_MIPS/Register/n639 ), 
        .CK(clk), .RN(n5666), .Q(\i_MIPS/Register/register[15][11] ), .QN(n596) );
  DFFRX1 \i_MIPS/Register/register_reg[15][13]  ( .D(\i_MIPS/Register/n641 ), 
        .CK(clk), .RN(n5666), .Q(\i_MIPS/Register/register[15][13] ), .QN(n311) );
  DFFRX1 \i_MIPS/Register/register_reg[15][14]  ( .D(\i_MIPS/Register/n642 ), 
        .CK(clk), .RN(n5666), .Q(\i_MIPS/Register/register[15][14] ), .QN(n326) );
  DFFRX1 \i_MIPS/Register/register_reg[15][16]  ( .D(\i_MIPS/Register/n644 ), 
        .CK(clk), .RN(n5666), .Q(\i_MIPS/Register/register[15][16] ), .QN(n593) );
  DFFRX1 \i_MIPS/Register/register_reg[15][20]  ( .D(\i_MIPS/Register/n648 ), 
        .CK(clk), .RN(n5667), .Q(\i_MIPS/Register/register[15][20] ), .QN(n592) );
  DFFRX1 \i_MIPS/Register/register_reg[15][21]  ( .D(\i_MIPS/Register/n649 ), 
        .CK(clk), .RN(n5667), .Q(\i_MIPS/Register/register[15][21] ), .QN(n666) );
  DFFRX1 \i_MIPS/Register/register_reg[15][22]  ( .D(\i_MIPS/Register/n650 ), 
        .CK(clk), .RN(n5667), .Q(\i_MIPS/Register/register[15][22] ), .QN(n216) );
  DFFRX1 \i_MIPS/Register/register_reg[15][23]  ( .D(\i_MIPS/Register/n651 ), 
        .CK(clk), .RN(n5667), .Q(\i_MIPS/Register/register[15][23] ), .QN(n575) );
  DFFRX1 \i_MIPS/Register/register_reg[15][24]  ( .D(\i_MIPS/Register/n652 ), 
        .CK(clk), .RN(n5667), .Q(\i_MIPS/Register/register[15][24] ), .QN(n581) );
  DFFRX1 \i_MIPS/Register/register_reg[15][25]  ( .D(\i_MIPS/Register/n653 ), 
        .CK(clk), .RN(n5667), .Q(\i_MIPS/Register/register[15][25] ), .QN(n569) );
  DFFRX1 \i_MIPS/Register/register_reg[15][26]  ( .D(\i_MIPS/Register/n654 ), 
        .CK(clk), .RN(n5667), .Q(\i_MIPS/Register/register[15][26] ), .QN(n594) );
  DFFRX1 \i_MIPS/Register/register_reg[15][27]  ( .D(\i_MIPS/Register/n655 ), 
        .CK(clk), .RN(n5667), .Q(\i_MIPS/Register/register[15][27] ), .QN(n576) );
  DFFRX1 \i_MIPS/Register/register_reg[15][28]  ( .D(\i_MIPS/Register/n656 ), 
        .CK(clk), .RN(n5667), .Q(\i_MIPS/Register/register[15][28] ), .QN(n583) );
  DFFRX1 \i_MIPS/Register/register_reg[15][29]  ( .D(\i_MIPS/Register/n657 ), 
        .CK(clk), .RN(n5667), .Q(\i_MIPS/Register/register[15][29] ), .QN(n325) );
  DFFRX1 \i_MIPS/Register/register_reg[13][2]  ( .D(\i_MIPS/Register/n694 ), 
        .CK(clk), .RN(n5670), .Q(\i_MIPS/Register/register[13][2] ), .QN(n574)
         );
  DFFRX1 \i_MIPS/Register/register_reg[13][3]  ( .D(\i_MIPS/Register/n695 ), 
        .CK(clk), .RN(n5671), .Q(\i_MIPS/Register/register[13][3] ), .QN(n586)
         );
  DFFRX1 \i_MIPS/Register/register_reg[13][4]  ( .D(\i_MIPS/Register/n696 ), 
        .CK(clk), .RN(n5671), .Q(\i_MIPS/Register/register[13][4] ), .QN(n341)
         );
  DFFRX1 \i_MIPS/Register/register_reg[13][5]  ( .D(\i_MIPS/Register/n697 ), 
        .CK(clk), .RN(n5671), .Q(\i_MIPS/Register/register[13][5] ), .QN(n526)
         );
  DFFRX1 \i_MIPS/Register/register_reg[13][6]  ( .D(\i_MIPS/Register/n698 ), 
        .CK(clk), .RN(n5671), .Q(\i_MIPS/Register/register[13][6] ), .QN(n661)
         );
  DFFRX1 \i_MIPS/Register/register_reg[13][7]  ( .D(\i_MIPS/Register/n699 ), 
        .CK(clk), .RN(n5671), .Q(\i_MIPS/Register/register[13][7] ), .QN(n493)
         );
  DFFRX1 \i_MIPS/Register/register_reg[13][8]  ( .D(\i_MIPS/Register/n700 ), 
        .CK(clk), .RN(n5671), .Q(\i_MIPS/Register/register[13][8] ), .QN(n566)
         );
  DFFRX1 \i_MIPS/Register/register_reg[13][9]  ( .D(\i_MIPS/Register/n701 ), 
        .CK(clk), .RN(n5671), .Q(\i_MIPS/Register/register[13][9] ), .QN(n564)
         );
  DFFRX1 \i_MIPS/Register/register_reg[13][10]  ( .D(\i_MIPS/Register/n702 ), 
        .CK(clk), .RN(n5671), .Q(\i_MIPS/Register/register[13][10] ), .QN(n344) );
  DFFRX1 \i_MIPS/Register/register_reg[13][11]  ( .D(\i_MIPS/Register/n703 ), 
        .CK(clk), .RN(n5671), .Q(\i_MIPS/Register/register[13][11] ), .QN(n597) );
  DFFRX1 \i_MIPS/Register/register_reg[13][12]  ( .D(\i_MIPS/Register/n704 ), 
        .CK(clk), .RN(n5671), .Q(\i_MIPS/Register/register[13][12] ), .QN(n663) );
  DFFRX1 \i_MIPS/Register/register_reg[13][13]  ( .D(\i_MIPS/Register/n705 ), 
        .CK(clk), .RN(n5671), .Q(\i_MIPS/Register/register[13][13] ), .QN(n568) );
  DFFRX1 \i_MIPS/Register/register_reg[13][14]  ( .D(\i_MIPS/Register/n706 ), 
        .CK(clk), .RN(n5671), .Q(\i_MIPS/Register/register[13][14] ), .QN(n338) );
  DFFRX1 \i_MIPS/Register/register_reg[13][15]  ( .D(\i_MIPS/Register/n707 ), 
        .CK(clk), .RN(n5672), .Q(\i_MIPS/Register/register[13][15] ), .QN(n525) );
  DFFRX1 \i_MIPS/Register/register_reg[13][16]  ( .D(\i_MIPS/Register/n708 ), 
        .CK(clk), .RN(n5672), .Q(\i_MIPS/Register/register[13][16] ), .QN(n262) );
  DFFRX1 \i_MIPS/Register/register_reg[13][17]  ( .D(\i_MIPS/Register/n709 ), 
        .CK(clk), .RN(n5672), .Q(\i_MIPS/Register/register[13][17] ), .QN(n488) );
  DFFRX1 \i_MIPS/Register/register_reg[13][18]  ( .D(\i_MIPS/Register/n710 ), 
        .CK(clk), .RN(n5672), .Q(\i_MIPS/Register/register[13][18] ), .QN(n435) );
  DFFRX1 \i_MIPS/Register/register_reg[13][20]  ( .D(\i_MIPS/Register/n712 ), 
        .CK(clk), .RN(n5672), .Q(\i_MIPS/Register/register[13][20] ), .QN(n260) );
  DFFRX1 \i_MIPS/Register/register_reg[13][21]  ( .D(\i_MIPS/Register/n713 ), 
        .CK(clk), .RN(n5672), .Q(\i_MIPS/Register/register[13][21] ), .QN(n264) );
  DFFRX1 \i_MIPS/Register/register_reg[13][22]  ( .D(\i_MIPS/Register/n714 ), 
        .CK(clk), .RN(n5672), .Q(\i_MIPS/Register/register[13][22] ), .QN(n434) );
  DFFRX1 \i_MIPS/Register/register_reg[13][23]  ( .D(\i_MIPS/Register/n715 ), 
        .CK(clk), .RN(n5672), .Q(\i_MIPS/Register/register[13][23] ), .QN(n259) );
  DFFRX1 \i_MIPS/Register/register_reg[13][24]  ( .D(\i_MIPS/Register/n716 ), 
        .CK(clk), .RN(n5672), .Q(\i_MIPS/Register/register[13][24] ), .QN(n582) );
  DFFRX1 \i_MIPS/Register/register_reg[13][25]  ( .D(\i_MIPS/Register/n717 ), 
        .CK(clk), .RN(n5672), .Q(\i_MIPS/Register/register[13][25] ), .QN(n257) );
  DFFRX1 \i_MIPS/Register/register_reg[13][26]  ( .D(\i_MIPS/Register/n718 ), 
        .CK(clk), .RN(n5672), .Q(\i_MIPS/Register/register[13][26] ), .QN(n266) );
  DFFRX1 \i_MIPS/Register/register_reg[13][27]  ( .D(\i_MIPS/Register/n719 ), 
        .CK(clk), .RN(n5673), .Q(\i_MIPS/Register/register[13][27] ), .QN(n577) );
  DFFRX1 \i_MIPS/Register/register_reg[13][28]  ( .D(\i_MIPS/Register/n720 ), 
        .CK(clk), .RN(n5673), .Q(\i_MIPS/Register/register[13][28] ), .QN(n584) );
  DFFRX1 \i_MIPS/Register/register_reg[13][29]  ( .D(\i_MIPS/Register/n721 ), 
        .CK(clk), .RN(n5673), .Q(\i_MIPS/Register/register[13][29] ), .QN(n336) );
  DFFRX1 \i_MIPS/Register/register_reg[13][31]  ( .D(\i_MIPS/Register/n723 ), 
        .CK(clk), .RN(n5673), .Q(\i_MIPS/Register/register[13][31] ), .QN(n659) );
  DFFRX1 \i_MIPS/Register/register_reg[12][24]  ( .D(\i_MIPS/Register/n748 ), 
        .CK(clk), .RN(n5675), .Q(\i_MIPS/Register/register[12][24] ), .QN(n639) );
  DFFRX1 \i_MIPS/Register/register_reg[11][2]  ( .D(\i_MIPS/Register/n758 ), 
        .CK(clk), .RN(n5676), .Q(\i_MIPS/Register/register[11][2] ), .QN(n573)
         );
  DFFRX1 \i_MIPS/Register/register_reg[11][3]  ( .D(\i_MIPS/Register/n759 ), 
        .CK(clk), .RN(n5676), .Q(\i_MIPS/Register/register[11][3] ), .QN(n504)
         );
  DFFRX1 \i_MIPS/Register/register_reg[11][4]  ( .D(\i_MIPS/Register/n760 ), 
        .CK(clk), .RN(n5676), .Q(\i_MIPS/Register/register[11][4] ), .QN(n591)
         );
  DFFRX1 \i_MIPS/Register/register_reg[11][5]  ( .D(\i_MIPS/Register/n761 ), 
        .CK(clk), .RN(n5676), .Q(\i_MIPS/Register/register[11][5] ), .QN(n542)
         );
  DFFRX1 \i_MIPS/Register/register_reg[11][6]  ( .D(\i_MIPS/Register/n762 ), 
        .CK(clk), .RN(n5676), .Q(\i_MIPS/Register/register[11][6] ), .QN(n528)
         );
  DFFRX1 \i_MIPS/Register/register_reg[11][7]  ( .D(\i_MIPS/Register/n763 ), 
        .CK(clk), .RN(n5676), .Q(\i_MIPS/Register/register[11][7] ), .QN(n532)
         );
  DFFRX1 \i_MIPS/Register/register_reg[11][9]  ( .D(\i_MIPS/Register/n765 ), 
        .CK(clk), .RN(n5676), .Q(\i_MIPS/Register/register[11][9] ), .QN(n496)
         );
  DFFRX1 \i_MIPS/Register/register_reg[11][10]  ( .D(\i_MIPS/Register/n766 ), 
        .CK(clk), .RN(n5676), .Q(\i_MIPS/Register/register[11][10] ), .QN(n507) );
  DFFRX1 \i_MIPS/Register/register_reg[11][11]  ( .D(\i_MIPS/Register/n767 ), 
        .CK(clk), .RN(n5677), .Q(\i_MIPS/Register/register[11][11] ), .QN(n509) );
  DFFRX1 \i_MIPS/Register/register_reg[11][12]  ( .D(\i_MIPS/Register/n768 ), 
        .CK(clk), .RN(n5677), .Q(\i_MIPS/Register/register[11][12] ), .QN(n536) );
  DFFRX1 \i_MIPS/Register/register_reg[11][13]  ( .D(\i_MIPS/Register/n769 ), 
        .CK(clk), .RN(n5677), .Q(\i_MIPS/Register/register[11][13] ), .QN(n555) );
  DFFRX1 \i_MIPS/Register/register_reg[11][14]  ( .D(\i_MIPS/Register/n770 ), 
        .CK(clk), .RN(n5677), .Q(\i_MIPS/Register/register[11][14] ), .QN(n498) );
  DFFRX1 \i_MIPS/Register/register_reg[11][16]  ( .D(\i_MIPS/Register/n772 ), 
        .CK(clk), .RN(n5677), .Q(\i_MIPS/Register/register[11][16] ), .QN(n508) );
  DFFRX1 \i_MIPS/Register/register_reg[11][18]  ( .D(\i_MIPS/Register/n774 ), 
        .CK(clk), .RN(n5677), .Q(\i_MIPS/Register/register[11][18] ), .QN(n534) );
  DFFRX1 \i_MIPS/Register/register_reg[11][20]  ( .D(\i_MIPS/Register/n776 ), 
        .CK(clk), .RN(n5677), .Q(\i_MIPS/Register/register[11][20] ), .QN(n553) );
  DFFRX1 \i_MIPS/Register/register_reg[11][21]  ( .D(\i_MIPS/Register/n777 ), 
        .CK(clk), .RN(n5677), .Q(\i_MIPS/Register/register[11][21] ), .QN(n530) );
  DFFRX1 \i_MIPS/Register/register_reg[11][22]  ( .D(\i_MIPS/Register/n778 ), 
        .CK(clk), .RN(n5677), .Q(\i_MIPS/Register/register[11][22] ), .QN(n589) );
  DFFRX1 \i_MIPS/Register/register_reg[11][23]  ( .D(\i_MIPS/Register/n779 ), 
        .CK(clk), .RN(n5678), .Q(\i_MIPS/Register/register[11][23] ), .QN(n502) );
  DFFRX1 \i_MIPS/Register/register_reg[11][24]  ( .D(\i_MIPS/Register/n780 ), 
        .CK(clk), .RN(n5678), .Q(\i_MIPS/Register/register[11][24] ), .QN(n540) );
  DFFRX1 \i_MIPS/Register/register_reg[11][25]  ( .D(\i_MIPS/Register/n781 ), 
        .CK(clk), .RN(n5678), .Q(\i_MIPS/Register/register[11][25] ), .QN(n552) );
  DFFRX1 \i_MIPS/Register/register_reg[11][26]  ( .D(\i_MIPS/Register/n782 ), 
        .CK(clk), .RN(n5678), .Q(\i_MIPS/Register/register[11][26] ), .QN(n595) );
  DFFRX1 \i_MIPS/Register/register_reg[11][27]  ( .D(\i_MIPS/Register/n783 ), 
        .CK(clk), .RN(n5678), .Q(\i_MIPS/Register/register[11][27] ), .QN(n541) );
  DFFRX1 \i_MIPS/Register/register_reg[11][28]  ( .D(\i_MIPS/Register/n784 ), 
        .CK(clk), .RN(n5678), .Q(\i_MIPS/Register/register[11][28] ), .QN(n668) );
  DFFRX1 \i_MIPS/Register/register_reg[11][29]  ( .D(\i_MIPS/Register/n785 ), 
        .CK(clk), .RN(n5678), .Q(\i_MIPS/Register/register[11][29] ), .QN(n345) );
  DFFRX1 \i_MIPS/Register/register_reg[9][2]  ( .D(\i_MIPS/Register/n822 ), 
        .CK(clk), .RN(n5681), .Q(\i_MIPS/Register/register[9][2] ), .QN(n481)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][3]  ( .D(\i_MIPS/Register/n823 ), 
        .CK(clk), .RN(n5681), .Q(\i_MIPS/Register/register[9][3] ), .QN(n562)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][4]  ( .D(\i_MIPS/Register/n824 ), 
        .CK(clk), .RN(n5681), .Q(\i_MIPS/Register/register[9][4] ), .QN(n484)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][5]  ( .D(\i_MIPS/Register/n825 ), 
        .CK(clk), .RN(n5681), .Q(\i_MIPS/Register/register[9][5] ), .QN(n656)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][6]  ( .D(\i_MIPS/Register/n826 ), 
        .CK(clk), .RN(n5681), .Q(\i_MIPS/Register/register[9][6] ), .QN(n516)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][7]  ( .D(\i_MIPS/Register/n827 ), 
        .CK(clk), .RN(n5682), .Q(\i_MIPS/Register/register[9][7] ), .QN(n522)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][8]  ( .D(\i_MIPS/Register/n828 ), 
        .CK(clk), .RN(n5682), .Q(\i_MIPS/Register/register[9][8] ), .QN(n213)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][9]  ( .D(\i_MIPS/Register/n829 ), 
        .CK(clk), .RN(n5682), .Q(\i_MIPS/Register/register[9][9] ), .QN(n211)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][10]  ( .D(\i_MIPS/Register/n830 ), 
        .CK(clk), .RN(n5682), .Q(\i_MIPS/Register/register[9][10] ), .QN(n492)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][11]  ( .D(\i_MIPS/Register/n831 ), 
        .CK(clk), .RN(n5682), .Q(\i_MIPS/Register/register[9][11] ), .QN(n521)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][12]  ( .D(\i_MIPS/Register/n832 ), 
        .CK(clk), .RN(n5682), .Q(\i_MIPS/Register/register[9][12] ), .QN(n209)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][13]  ( .D(\i_MIPS/Register/n833 ), 
        .CK(clk), .RN(n5682), .Q(\i_MIPS/Register/register[9][13] ), .QN(n207)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][14]  ( .D(\i_MIPS/Register/n834 ), 
        .CK(clk), .RN(n5682), .Q(\i_MIPS/Register/register[9][14] ), .QN(n219)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][15]  ( .D(\i_MIPS/Register/n835 ), 
        .CK(clk), .RN(n5682), .Q(\i_MIPS/Register/register[9][15] ), .QN(n518)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][16]  ( .D(\i_MIPS/Register/n836 ), 
        .CK(clk), .RN(n5682), .Q(\i_MIPS/Register/register[9][16] ), .QN(n512)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][17]  ( .D(\i_MIPS/Register/n837 ), 
        .CK(clk), .RN(n5682), .Q(\i_MIPS/Register/register[9][17] ), .QN(n558)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][18]  ( .D(\i_MIPS/Register/n838 ), 
        .CK(clk), .RN(n5682), .Q(\i_MIPS/Register/register[9][18] ), .QN(n333)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][20]  ( .D(\i_MIPS/Register/n840 ), 
        .CK(clk), .RN(n5683), .Q(\i_MIPS/Register/register[9][20] ), .QN(n648)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][21]  ( .D(\i_MIPS/Register/n841 ), 
        .CK(clk), .RN(n5683), .Q(\i_MIPS/Register/register[9][21] ), .QN(n546)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][22]  ( .D(\i_MIPS/Register/n842 ), 
        .CK(clk), .RN(n5683), .Q(\i_MIPS/Register/register[9][22] ), .QN(n335)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][23]  ( .D(\i_MIPS/Register/n843 ), 
        .CK(clk), .RN(n5683), .Q(\i_MIPS/Register/register[9][23] ), .QN(n510)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][24]  ( .D(\i_MIPS/Register/n844 ), 
        .CK(clk), .RN(n5683), .Q(\i_MIPS/Register/register[9][24] ), .QN(n561)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][25]  ( .D(\i_MIPS/Register/n845 ), 
        .CK(clk), .RN(n5683), .Q(\i_MIPS/Register/register[9][25] ), .QN(n548)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][26]  ( .D(\i_MIPS/Register/n846 ), 
        .CK(clk), .RN(n5683), .Q(\i_MIPS/Register/register[9][26] ), .QN(n692)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][27]  ( .D(\i_MIPS/Register/n847 ), 
        .CK(clk), .RN(n5683), .Q(\i_MIPS/Register/register[9][27] ), .QN(n654)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][28]  ( .D(\i_MIPS/Register/n848 ), 
        .CK(clk), .RN(n5683), .Q(\i_MIPS/Register/register[9][28] ), .QN(n559)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][29]  ( .D(\i_MIPS/Register/n849 ), 
        .CK(clk), .RN(n5683), .Q(\i_MIPS/Register/register[9][29] ), .QN(n205)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][31]  ( .D(\i_MIPS/Register/n851 ), 
        .CK(clk), .RN(n5684), .Q(\i_MIPS/Register/register[9][31] ), .QN(n651)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][3]  ( .D(\i_MIPS/Register/n855 ), 
        .CK(clk), .RN(n5684), .Q(\i_MIPS/Register/register[8][3] ), .QN(n621)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][24]  ( .D(\i_MIPS/Register/n876 ), 
        .CK(clk), .RN(n5686), .Q(\i_MIPS/Register/register[8][24] ), .QN(n613)
         );
  DFFRX1 \i_MIPS/Register/register_reg[23][2]  ( .D(\i_MIPS/Register/n374 ), 
        .CK(clk), .RN(n5644), .Q(\i_MIPS/Register/register[23][2] ), .QN(n2080) );
  DFFRX1 \i_MIPS/Register/register_reg[23][3]  ( .D(\i_MIPS/Register/n375 ), 
        .CK(clk), .RN(n5644), .Q(\i_MIPS/Register/register[23][3] ), .QN(n2094) );
  DFFRX1 \i_MIPS/Register/register_reg[23][4]  ( .D(\i_MIPS/Register/n376 ), 
        .CK(clk), .RN(n5644), .Q(\i_MIPS/Register/register[23][4] ), .QN(n1916) );
  DFFRX1 \i_MIPS/Register/register_reg[23][5]  ( .D(\i_MIPS/Register/n377 ), 
        .CK(clk), .RN(n5644), .Q(\i_MIPS/Register/register[23][5] ), .QN(n2197) );
  DFFRX1 \i_MIPS/Register/register_reg[23][6]  ( .D(\i_MIPS/Register/n378 ), 
        .CK(clk), .RN(n5644), .Q(\i_MIPS/Register/register[23][6] ), .QN(n724)
         );
  DFFRX1 \i_MIPS/Register/register_reg[23][7]  ( .D(\i_MIPS/Register/n379 ), 
        .CK(clk), .RN(n5644), .Q(\i_MIPS/Register/register[23][7] ), .QN(n2189) );
  DFFRX1 \i_MIPS/Register/register_reg[23][10]  ( .D(\i_MIPS/Register/n382 ), 
        .CK(clk), .RN(n5644), .Q(\i_MIPS/Register/register[23][10] ), .QN(
        n1919) );
  DFFRX1 \i_MIPS/Register/register_reg[23][11]  ( .D(\i_MIPS/Register/n383 ), 
        .CK(clk), .RN(n5645), .Q(\i_MIPS/Register/register[23][11] ), .QN(
        n1918) );
  DFFRX1 \i_MIPS/Register/register_reg[23][13]  ( .D(\i_MIPS/Register/n385 ), 
        .CK(clk), .RN(n5645), .Q(\i_MIPS/Register/register[23][13] ), .QN(
        n2074) );
  DFFRX1 \i_MIPS/Register/register_reg[23][14]  ( .D(\i_MIPS/Register/n386 ), 
        .CK(clk), .RN(n5645), .Q(\i_MIPS/Register/register[23][14] ), .QN(
        n1927) );
  DFFRX1 \i_MIPS/Register/register_reg[23][16]  ( .D(\i_MIPS/Register/n388 ), 
        .CK(clk), .RN(n5645), .Q(\i_MIPS/Register/register[23][16] ), .QN(
        n2106) );
  DFFRX1 \i_MIPS/Register/register_reg[23][18]  ( .D(\i_MIPS/Register/n390 ), 
        .CK(clk), .RN(n5645), .Q(\i_MIPS/Register/register[23][18] ), .QN(n726) );
  DFFRX1 \i_MIPS/Register/register_reg[23][20]  ( .D(\i_MIPS/Register/n392 ), 
        .CK(clk), .RN(n5645), .Q(\i_MIPS/Register/register[23][20] ), .QN(
        n2105) );
  DFFRX1 \i_MIPS/Register/register_reg[23][21]  ( .D(\i_MIPS/Register/n393 ), 
        .CK(clk), .RN(n5645), .Q(\i_MIPS/Register/register[23][21] ), .QN(
        n2193) );
  DFFRX1 \i_MIPS/Register/register_reg[23][22]  ( .D(\i_MIPS/Register/n394 ), 
        .CK(clk), .RN(n5645), .Q(\i_MIPS/Register/register[23][22] ), .QN(n717) );
  DFFRX1 \i_MIPS/Register/register_reg[23][23]  ( .D(\i_MIPS/Register/n395 ), 
        .CK(clk), .RN(n5646), .Q(\i_MIPS/Register/register[23][23] ), .QN(
        n2086) );
  DFFRX1 \i_MIPS/Register/register_reg[23][24]  ( .D(\i_MIPS/Register/n396 ), 
        .CK(clk), .RN(n5646), .Q(\i_MIPS/Register/register[23][24] ), .QN(
        n2090) );
  DFFRX1 \i_MIPS/Register/register_reg[23][25]  ( .D(\i_MIPS/Register/n397 ), 
        .CK(clk), .RN(n5646), .Q(\i_MIPS/Register/register[23][25] ), .QN(
        n2078) );
  DFFRX1 \i_MIPS/Register/register_reg[23][26]  ( .D(\i_MIPS/Register/n398 ), 
        .CK(clk), .RN(n5646), .Q(\i_MIPS/Register/register[23][26] ), .QN(
        n2107) );
  DFFRX1 \i_MIPS/Register/register_reg[23][27]  ( .D(\i_MIPS/Register/n399 ), 
        .CK(clk), .RN(n5646), .Q(\i_MIPS/Register/register[23][27] ), .QN(
        n2265) );
  DFFRX1 \i_MIPS/Register/register_reg[23][28]  ( .D(\i_MIPS/Register/n400 ), 
        .CK(clk), .RN(n5646), .Q(\i_MIPS/Register/register[23][28] ), .QN(
        n2092) );
  DFFRX1 \i_MIPS/Register/register_reg[23][29]  ( .D(\i_MIPS/Register/n401 ), 
        .CK(clk), .RN(n5646), .Q(\i_MIPS/Register/register[23][29] ), .QN(
        n1902) );
  DFFRX1 \i_MIPS/Register/register_reg[21][2]  ( .D(\i_MIPS/Register/n438 ), 
        .CK(clk), .RN(n5649), .Q(\i_MIPS/Register/register[21][2] ), .QN(n2082) );
  DFFRX1 \i_MIPS/Register/register_reg[21][3]  ( .D(\i_MIPS/Register/n439 ), 
        .CK(clk), .RN(n5649), .Q(\i_MIPS/Register/register[21][3] ), .QN(n2095) );
  DFFRX1 \i_MIPS/Register/register_reg[21][4]  ( .D(\i_MIPS/Register/n440 ), 
        .CK(clk), .RN(n5649), .Q(\i_MIPS/Register/register[21][4] ), .QN(n1921) );
  DFFRX1 \i_MIPS/Register/register_reg[21][5]  ( .D(\i_MIPS/Register/n441 ), 
        .CK(clk), .RN(n5649), .Q(\i_MIPS/Register/register[21][5] ), .QN(n2054) );
  DFFRX1 \i_MIPS/Register/register_reg[21][6]  ( .D(\i_MIPS/Register/n442 ), 
        .CK(clk), .RN(n5649), .Q(\i_MIPS/Register/register[21][6] ), .QN(n2184) );
  DFFRX1 \i_MIPS/Register/register_reg[21][7]  ( .D(\i_MIPS/Register/n443 ), 
        .CK(clk), .RN(n5650), .Q(\i_MIPS/Register/register[21][7] ), .QN(n2278) );
  DFFRX1 \i_MIPS/Register/register_reg[21][8]  ( .D(\i_MIPS/Register/n444 ), 
        .CK(clk), .RN(n5650), .Q(\i_MIPS/Register/register[21][8] ), .QN(n2071) );
  DFFRX1 \i_MIPS/Register/register_reg[21][9]  ( .D(\i_MIPS/Register/n445 ), 
        .CK(clk), .RN(n5650), .Q(\i_MIPS/Register/register[21][9] ), .QN(n2067) );
  DFFRX1 \i_MIPS/Register/register_reg[21][10]  ( .D(\i_MIPS/Register/n446 ), 
        .CK(clk), .RN(n5650), .Q(\i_MIPS/Register/register[21][10] ), .QN(
        n1924) );
  DFFRX1 \i_MIPS/Register/register_reg[21][11]  ( .D(\i_MIPS/Register/n447 ), 
        .CK(clk), .RN(n5650), .Q(\i_MIPS/Register/register[21][11] ), .QN(
        n1923) );
  DFFRX1 \i_MIPS/Register/register_reg[21][12]  ( .D(\i_MIPS/Register/n448 ), 
        .CK(clk), .RN(n5650), .Q(\i_MIPS/Register/register[21][12] ), .QN(
        n1932) );
  DFFRX1 \i_MIPS/Register/register_reg[21][13]  ( .D(\i_MIPS/Register/n449 ), 
        .CK(clk), .RN(n5650), .Q(\i_MIPS/Register/register[21][13] ), .QN(
        n2075) );
  DFFRX1 \i_MIPS/Register/register_reg[21][14]  ( .D(\i_MIPS/Register/n450 ), 
        .CK(clk), .RN(n5650), .Q(\i_MIPS/Register/register[21][14] ), .QN(
        n1931) );
  DFFRX1 \i_MIPS/Register/register_reg[21][15]  ( .D(\i_MIPS/Register/n451 ), 
        .CK(clk), .RN(n5650), .Q(\i_MIPS/Register/register[21][15] ), .QN(
        n2279) );
  DFFRX1 \i_MIPS/Register/register_reg[21][16]  ( .D(\i_MIPS/Register/n452 ), 
        .CK(clk), .RN(n5650), .Q(\i_MIPS/Register/register[21][16] ), .QN(
        n2243) );
  DFFRX1 \i_MIPS/Register/register_reg[21][17]  ( .D(\i_MIPS/Register/n453 ), 
        .CK(clk), .RN(n5650), .Q(\i_MIPS/Register/register[21][17] ), .QN(
        n2231) );
  DFFRX1 \i_MIPS/Register/register_reg[21][18]  ( .D(\i_MIPS/Register/n454 ), 
        .CK(clk), .RN(n5650), .Q(\i_MIPS/Register/register[21][18] ), .QN(
        n2000) );
  DFFRX1 \i_MIPS/Register/register_reg[21][20]  ( .D(\i_MIPS/Register/n456 ), 
        .CK(clk), .RN(n5651), .Q(\i_MIPS/Register/register[21][20] ), .QN(
        n2234) );
  DFFRX1 \i_MIPS/Register/register_reg[21][21]  ( .D(\i_MIPS/Register/n457 ), 
        .CK(clk), .RN(n5651), .Q(\i_MIPS/Register/register[21][21] ), .QN(
        n2276) );
  DFFRX1 \i_MIPS/Register/register_reg[21][22]  ( .D(\i_MIPS/Register/n458 ), 
        .CK(clk), .RN(n5651), .Q(\i_MIPS/Register/register[21][22] ), .QN(
        n1996) );
  DFFRX1 \i_MIPS/Register/register_reg[21][23]  ( .D(\i_MIPS/Register/n459 ), 
        .CK(clk), .RN(n5651), .Q(\i_MIPS/Register/register[21][23] ), .QN(
        n2240) );
  DFFRX1 \i_MIPS/Register/register_reg[21][24]  ( .D(\i_MIPS/Register/n460 ), 
        .CK(clk), .RN(n5651), .Q(\i_MIPS/Register/register[21][24] ), .QN(
        n2091) );
  DFFRX1 \i_MIPS/Register/register_reg[21][25]  ( .D(\i_MIPS/Register/n461 ), 
        .CK(clk), .RN(n5651), .Q(\i_MIPS/Register/register[21][25] ), .QN(
        n2238) );
  DFFRX1 \i_MIPS/Register/register_reg[21][26]  ( .D(\i_MIPS/Register/n462 ), 
        .CK(clk), .RN(n5651), .Q(\i_MIPS/Register/register[21][26] ), .QN(
        n2109) );
  DFFRX1 \i_MIPS/Register/register_reg[21][27]  ( .D(\i_MIPS/Register/n463 ), 
        .CK(clk), .RN(n5651), .Q(\i_MIPS/Register/register[21][27] ), .QN(
        n2195) );
  DFFRX1 \i_MIPS/Register/register_reg[21][28]  ( .D(\i_MIPS/Register/n464 ), 
        .CK(clk), .RN(n5651), .Q(\i_MIPS/Register/register[21][28] ), .QN(
        n2093) );
  DFFRX1 \i_MIPS/Register/register_reg[21][29]  ( .D(\i_MIPS/Register/n465 ), 
        .CK(clk), .RN(n5651), .Q(\i_MIPS/Register/register[21][29] ), .QN(
        n1914) );
  DFFRX1 \i_MIPS/Register/register_reg[21][31]  ( .D(\i_MIPS/Register/n467 ), 
        .CK(clk), .RN(n5652), .Q(\i_MIPS/Register/register[21][31] ), .QN(
        n2181) );
  DFFRX1 \i_MIPS/Register/register_reg[20][3]  ( .D(\i_MIPS/Register/n471 ), 
        .CK(clk), .RN(n5652), .Q(\i_MIPS/Register/register[20][3] ), .QN(n2121) );
  DFFRX1 \i_MIPS/Register/register_reg[20][16]  ( .D(\i_MIPS/Register/n484 ), 
        .CK(clk), .RN(n5653), .Q(\i_MIPS/Register/register[20][16] ), .QN(
        n1907) );
  DFFRX1 \i_MIPS/Register/register_reg[20][22]  ( .D(\i_MIPS/Register/n490 ), 
        .CK(clk), .RN(n5653), .Q(\i_MIPS/Register/register[20][22] ), .QN(
        n2120) );
  DFFRX1 \i_MIPS/Register/register_reg[20][23]  ( .D(\i_MIPS/Register/n491 ), 
        .CK(clk), .RN(n5654), .Q(\i_MIPS/Register/register[20][23] ), .QN(
        n1904) );
  DFFRX1 \i_MIPS/Register/register_reg[20][24]  ( .D(\i_MIPS/Register/n492 ), 
        .CK(clk), .RN(n5654), .Q(\i_MIPS/Register/register[20][24] ), .QN(
        n2119) );
  DFFRX1 \i_MIPS/Register/register_reg[19][2]  ( .D(\i_MIPS/Register/n502 ), 
        .CK(clk), .RN(n5654), .Q(\i_MIPS/Register/register[19][2] ), .QN(n2081) );
  DFFRX1 \i_MIPS/Register/register_reg[19][3]  ( .D(\i_MIPS/Register/n503 ), 
        .CK(clk), .RN(n5655), .Q(\i_MIPS/Register/register[19][3] ), .QN(n2255) );
  DFFRX1 \i_MIPS/Register/register_reg[19][4]  ( .D(\i_MIPS/Register/n504 ), 
        .CK(clk), .RN(n5655), .Q(\i_MIPS/Register/register[19][4] ), .QN(n2103) );
  DFFRX1 \i_MIPS/Register/register_reg[19][5]  ( .D(\i_MIPS/Register/n505 ), 
        .CK(clk), .RN(n5655), .Q(\i_MIPS/Register/register[19][5] ), .QN(n2267) );
  DFFRX1 \i_MIPS/Register/register_reg[19][6]  ( .D(\i_MIPS/Register/n506 ), 
        .CK(clk), .RN(n5655), .Q(\i_MIPS/Register/register[19][6] ), .QN(n2282) );
  DFFRX1 \i_MIPS/Register/register_reg[19][7]  ( .D(\i_MIPS/Register/n507 ), 
        .CK(clk), .RN(n5655), .Q(\i_MIPS/Register/register[19][7] ), .QN(n2286) );
  DFFRX1 \i_MIPS/Register/register_reg[19][8]  ( .D(\i_MIPS/Register/n508 ), 
        .CK(clk), .RN(n5655), .Q(\i_MIPS/Register/register[19][8] ), .QN(n2251) );
  DFFRX1 \i_MIPS/Register/register_reg[19][9]  ( .D(\i_MIPS/Register/n509 ), 
        .CK(clk), .RN(n5655), .Q(\i_MIPS/Register/register[19][9] ), .QN(n2059) );
  DFFRX1 \i_MIPS/Register/register_reg[19][10]  ( .D(\i_MIPS/Register/n510 ), 
        .CK(clk), .RN(n5655), .Q(\i_MIPS/Register/register[19][10] ), .QN(
        n2258) );
  DFFRX1 \i_MIPS/Register/register_reg[19][11]  ( .D(\i_MIPS/Register/n511 ), 
        .CK(clk), .RN(n5655), .Q(\i_MIPS/Register/register[19][11] ), .QN(
        n2235) );
  DFFRX1 \i_MIPS/Register/register_reg[19][12]  ( .D(\i_MIPS/Register/n512 ), 
        .CK(clk), .RN(n5655), .Q(\i_MIPS/Register/register[19][12] ), .QN(
        n2290) );
  DFFRX1 \i_MIPS/Register/register_reg[19][13]  ( .D(\i_MIPS/Register/n513 ), 
        .CK(clk), .RN(n5655), .Q(\i_MIPS/Register/register[19][13] ), .QN(
        n2057) );
  DFFRX1 \i_MIPS/Register/register_reg[19][14]  ( .D(\i_MIPS/Register/n514 ), 
        .CK(clk), .RN(n5655), .Q(\i_MIPS/Register/register[19][14] ), .QN(
        n2172) );
  DFFRX1 \i_MIPS/Register/register_reg[19][15]  ( .D(\i_MIPS/Register/n515 ), 
        .CK(clk), .RN(n5656), .Q(\i_MIPS/Register/register[19][15] ), .QN(
        n2292) );
  DFFRX1 \i_MIPS/Register/register_reg[19][16]  ( .D(\i_MIPS/Register/n516 ), 
        .CK(clk), .RN(n5656), .Q(\i_MIPS/Register/register[19][16] ), .QN(
        n2257) );
  DFFRX1 \i_MIPS/Register/register_reg[19][17]  ( .D(\i_MIPS/Register/n517 ), 
        .CK(clk), .RN(n5656), .Q(\i_MIPS/Register/register[19][17] ), .QN(
        n2246) );
  DFFRX1 \i_MIPS/Register/register_reg[19][18]  ( .D(\i_MIPS/Register/n518 ), 
        .CK(clk), .RN(n5656), .Q(\i_MIPS/Register/register[19][18] ), .QN(
        n2288) );
  DFFRX1 \i_MIPS/Register/register_reg[19][20]  ( .D(\i_MIPS/Register/n520 ), 
        .CK(clk), .RN(n5656), .Q(\i_MIPS/Register/register[19][20] ), .QN(
        n2060) );
  DFFRX1 \i_MIPS/Register/register_reg[19][21]  ( .D(\i_MIPS/Register/n521 ), 
        .CK(clk), .RN(n5656), .Q(\i_MIPS/Register/register[19][21] ), .QN(
        n2284) );
  DFFRX1 \i_MIPS/Register/register_reg[19][22]  ( .D(\i_MIPS/Register/n522 ), 
        .CK(clk), .RN(n5656), .Q(\i_MIPS/Register/register[19][22] ), .QN(
        n2102) );
  DFFRX1 \i_MIPS/Register/register_reg[19][23]  ( .D(\i_MIPS/Register/n523 ), 
        .CK(clk), .RN(n5656), .Q(\i_MIPS/Register/register[19][23] ), .QN(
        n2253) );
  DFFRX1 \i_MIPS/Register/register_reg[19][24]  ( .D(\i_MIPS/Register/n524 ), 
        .CK(clk), .RN(n5656), .Q(\i_MIPS/Register/register[19][24] ), .QN(
        n2294) );
  DFFRX1 \i_MIPS/Register/register_reg[19][25]  ( .D(\i_MIPS/Register/n525 ), 
        .CK(clk), .RN(n5656), .Q(\i_MIPS/Register/register[19][25] ), .QN(
        n2249) );
  DFFRX1 \i_MIPS/Register/register_reg[19][26]  ( .D(\i_MIPS/Register/n526 ), 
        .CK(clk), .RN(n5656), .Q(\i_MIPS/Register/register[19][26] ), .QN(
        n2108) );
  DFFRX1 \i_MIPS/Register/register_reg[19][27]  ( .D(\i_MIPS/Register/n527 ), 
        .CK(clk), .RN(n5657), .Q(\i_MIPS/Register/register[19][27] ), .QN(
        n2168) );
  DFFRX1 \i_MIPS/Register/register_reg[19][28]  ( .D(\i_MIPS/Register/n528 ), 
        .CK(clk), .RN(n5657), .Q(\i_MIPS/Register/register[19][28] ), .QN(
        n2053) );
  DFFRX1 \i_MIPS/Register/register_reg[19][29]  ( .D(\i_MIPS/Register/n529 ), 
        .CK(clk), .RN(n5657), .Q(\i_MIPS/Register/register[19][29] ), .QN(
        n1933) );
  DFFRX1 \i_MIPS/Register/register_reg[19][31]  ( .D(\i_MIPS/Register/n531 ), 
        .CK(clk), .RN(n5657), .Q(\i_MIPS/Register/register[19][31] ), .QN(
        n2298) );
  DFFRX1 \i_MIPS/Register/register_reg[17][2]  ( .D(\i_MIPS/Register/n566 ), 
        .CK(clk), .RN(n5660), .Q(\i_MIPS/Register/register[17][2] ), .QN(n2033) );
  DFFRX1 \i_MIPS/Register/register_reg[17][3]  ( .D(\i_MIPS/Register/n567 ), 
        .CK(clk), .RN(n5660), .Q(\i_MIPS/Register/register[17][3] ), .QN(n2176) );
  DFFRX1 \i_MIPS/Register/register_reg[17][4]  ( .D(\i_MIPS/Register/n568 ), 
        .CK(clk), .RN(n5660), .Q(\i_MIPS/Register/register[17][4] ), .QN(n2035) );
  DFFRX1 \i_MIPS/Register/register_reg[17][5]  ( .D(\i_MIPS/Register/n569 ), 
        .CK(clk), .RN(n5660), .Q(\i_MIPS/Register/register[17][5] ), .QN(n2178) );
  DFFRX1 \i_MIPS/Register/register_reg[17][6]  ( .D(\i_MIPS/Register/n570 ), 
        .CK(clk), .RN(n5660), .Q(\i_MIPS/Register/register[17][6] ), .QN(n2268) );
  DFFRX1 \i_MIPS/Register/register_reg[17][7]  ( .D(\i_MIPS/Register/n571 ), 
        .CK(clk), .RN(n5660), .Q(\i_MIPS/Register/register[17][7] ), .QN(n2273) );
  DFFRX1 \i_MIPS/Register/register_reg[17][8]  ( .D(\i_MIPS/Register/n572 ), 
        .CK(clk), .RN(n5660), .Q(\i_MIPS/Register/register[17][8] ), .QN(n2312) );
  DFFRX1 \i_MIPS/Register/register_reg[17][9]  ( .D(\i_MIPS/Register/n573 ), 
        .CK(clk), .RN(n5660), .Q(\i_MIPS/Register/register[17][9] ), .QN(n2310) );
  DFFRX1 \i_MIPS/Register/register_reg[17][10]  ( .D(\i_MIPS/Register/n574 ), 
        .CK(clk), .RN(n5660), .Q(\i_MIPS/Register/register[17][10] ), .QN(
        n2236) );
  DFFRX1 \i_MIPS/Register/register_reg[17][11]  ( .D(\i_MIPS/Register/n575 ), 
        .CK(clk), .RN(n5661), .Q(\i_MIPS/Register/register[17][11] ), .QN(
        n2272) );
  DFFRX1 \i_MIPS/Register/register_reg[17][12]  ( .D(\i_MIPS/Register/n576 ), 
        .CK(clk), .RN(n5661), .Q(\i_MIPS/Register/register[17][12] ), .QN(
        n2308) );
  DFFRX1 \i_MIPS/Register/register_reg[17][13]  ( .D(\i_MIPS/Register/n577 ), 
        .CK(clk), .RN(n5661), .Q(\i_MIPS/Register/register[17][13] ), .QN(
        n2306) );
  DFFRX1 \i_MIPS/Register/register_reg[17][14]  ( .D(\i_MIPS/Register/n578 ), 
        .CK(clk), .RN(n5661), .Q(\i_MIPS/Register/register[17][14] ), .QN(
        n2170) );
  DFFRX1 \i_MIPS/Register/register_reg[17][15]  ( .D(\i_MIPS/Register/n579 ), 
        .CK(clk), .RN(n5661), .Q(\i_MIPS/Register/register[17][15] ), .QN(
        n2270) );
  DFFRX1 \i_MIPS/Register/register_reg[17][16]  ( .D(\i_MIPS/Register/n580 ), 
        .CK(clk), .RN(n5661), .Q(\i_MIPS/Register/register[17][16] ), .QN(
        n2263) );
  DFFRX1 \i_MIPS/Register/register_reg[17][17]  ( .D(\i_MIPS/Register/n581 ), 
        .CK(clk), .RN(n5661), .Q(\i_MIPS/Register/register[17][17] ), .QN(
        n1930) );
  DFFRX1 \i_MIPS/Register/register_reg[17][18]  ( .D(\i_MIPS/Register/n582 ), 
        .CK(clk), .RN(n5661), .Q(\i_MIPS/Register/register[17][18] ), .QN(
        n1929) );
  DFFRX1 \i_MIPS/Register/register_reg[17][20]  ( .D(\i_MIPS/Register/n584 ), 
        .CK(clk), .RN(n5661), .Q(\i_MIPS/Register/register[17][20] ), .QN(
        n2305) );
  DFFRX1 \i_MIPS/Register/register_reg[17][21]  ( .D(\i_MIPS/Register/n585 ), 
        .CK(clk), .RN(n5661), .Q(\i_MIPS/Register/register[17][21] ), .QN(
        n2300) );
  DFFRX1 \i_MIPS/Register/register_reg[17][22]  ( .D(\i_MIPS/Register/n586 ), 
        .CK(clk), .RN(n5661), .Q(\i_MIPS/Register/register[17][22] ), .QN(
        n1911) );
  DFFRX1 \i_MIPS/Register/register_reg[17][23]  ( .D(\i_MIPS/Register/n587 ), 
        .CK(clk), .RN(n5662), .Q(\i_MIPS/Register/register[17][23] ), .QN(
        n2304) );
  DFFRX1 \i_MIPS/Register/register_reg[17][24]  ( .D(\i_MIPS/Register/n588 ), 
        .CK(clk), .RN(n5662), .Q(\i_MIPS/Register/register[17][24] ), .QN(
        n2063) );
  DFFRX1 \i_MIPS/Register/register_reg[17][25]  ( .D(\i_MIPS/Register/n589 ), 
        .CK(clk), .RN(n5662), .Q(\i_MIPS/Register/register[17][25] ), .QN(
        n2302) );
  DFFRX1 \i_MIPS/Register/register_reg[17][26]  ( .D(\i_MIPS/Register/n590 ), 
        .CK(clk), .RN(n5662), .Q(\i_MIPS/Register/register[17][26] ), .QN(
        n2036) );
  DFFRX1 \i_MIPS/Register/register_reg[17][27]  ( .D(\i_MIPS/Register/n591 ), 
        .CK(clk), .RN(n5662), .Q(\i_MIPS/Register/register[17][27] ), .QN(
        n2175) );
  DFFRX1 \i_MIPS/Register/register_reg[17][28]  ( .D(\i_MIPS/Register/n592 ), 
        .CK(clk), .RN(n5662), .Q(\i_MIPS/Register/register[17][28] ), .QN(
        n2052) );
  DFFRX1 \i_MIPS/Register/register_reg[17][29]  ( .D(\i_MIPS/Register/n593 ), 
        .CK(clk), .RN(n5662), .Q(\i_MIPS/Register/register[17][29] ), .QN(
        n2155) );
  DFFRX1 \i_MIPS/Register/register_reg[17][31]  ( .D(\i_MIPS/Register/n595 ), 
        .CK(clk), .RN(n5662), .Q(\i_MIPS/Register/register[17][31] ), .QN(
        n2173) );
  DFFRX1 \i_MIPS/Register/register_reg[16][2]  ( .D(\i_MIPS/Register/n598 ), 
        .CK(clk), .RN(n5662), .Q(\i_MIPS/Register/register[16][2] ), .QN(n2146) );
  DFFRX1 \i_MIPS/Register/register_reg[16][3]  ( .D(\i_MIPS/Register/n599 ), 
        .CK(clk), .RN(n5663), .Q(\i_MIPS/Register/register[16][3] ), .QN(n2140) );
  DFFRX1 \i_MIPS/Register/register_reg[16][16]  ( .D(\i_MIPS/Register/n612 ), 
        .CK(clk), .RN(n5664), .Q(\i_MIPS/Register/register[16][16] ), .QN(
        n2134) );
  DFFRX1 \i_MIPS/Register/register_reg[16][20]  ( .D(\i_MIPS/Register/n616 ), 
        .CK(clk), .RN(n5664), .Q(\i_MIPS/Register/register[16][20] ), .QN(
        n2142) );
  DFFRX1 \i_MIPS/Register/register_reg[16][21]  ( .D(\i_MIPS/Register/n617 ), 
        .CK(clk), .RN(n5664), .Q(\i_MIPS/Register/register[16][21] ), .QN(
        n2143) );
  DFFRX1 \i_MIPS/Register/register_reg[16][22]  ( .D(\i_MIPS/Register/n618 ), 
        .CK(clk), .RN(n5664), .Q(\i_MIPS/Register/register[16][22] ), .QN(
        n2138) );
  DFFRX1 \i_MIPS/Register/register_reg[16][23]  ( .D(\i_MIPS/Register/n619 ), 
        .CK(clk), .RN(n5664), .Q(\i_MIPS/Register/register[16][23] ), .QN(
        n2136) );
  DFFRX1 \i_MIPS/Register/register_reg[16][24]  ( .D(\i_MIPS/Register/n620 ), 
        .CK(clk), .RN(n5664), .Q(\i_MIPS/Register/register[16][24] ), .QN(
        n2132) );
  DFFRX1 \i_MIPS/Register/register_reg[7][2]  ( .D(\i_MIPS/Register/n886 ), 
        .CK(clk), .RN(n5686), .Q(\i_MIPS/Register/register[7][2] ), .QN(n2083)
         );
  DFFRX1 \i_MIPS/Register/register_reg[7][3]  ( .D(\i_MIPS/Register/n887 ), 
        .CK(clk), .RN(n5687), .Q(\i_MIPS/Register/register[7][3] ), .QN(n2100)
         );
  DFFRX1 \i_MIPS/Register/register_reg[7][4]  ( .D(\i_MIPS/Register/n888 ), 
        .CK(clk), .RN(n5687), .Q(\i_MIPS/Register/register[7][4] ), .QN(n1917)
         );
  DFFRX1 \i_MIPS/Register/register_reg[7][5]  ( .D(\i_MIPS/Register/n889 ), 
        .CK(clk), .RN(n5687), .Q(\i_MIPS/Register/register[7][5] ), .QN(n2198)
         );
  DFFRX1 \i_MIPS/Register/register_reg[7][6]  ( .D(\i_MIPS/Register/n890 ), 
        .CK(clk), .RN(n5687), .Q(\i_MIPS/Register/register[7][6] ), .QN(n725)
         );
  DFFRX1 \i_MIPS/Register/register_reg[7][7]  ( .D(\i_MIPS/Register/n891 ), 
        .CK(clk), .RN(n5687), .Q(\i_MIPS/Register/register[7][7] ), .QN(n2190)
         );
  DFFRX1 \i_MIPS/Register/register_reg[7][10]  ( .D(\i_MIPS/Register/n894 ), 
        .CK(clk), .RN(n5687), .Q(\i_MIPS/Register/register[7][10] ), .QN(n1920) );
  DFFRX1 \i_MIPS/Register/register_reg[7][11]  ( .D(\i_MIPS/Register/n895 ), 
        .CK(clk), .RN(n5687), .Q(\i_MIPS/Register/register[7][11] ), .QN(n2116) );
  DFFRX1 \i_MIPS/Register/register_reg[7][13]  ( .D(\i_MIPS/Register/n897 ), 
        .CK(clk), .RN(n5687), .Q(\i_MIPS/Register/register[7][13] ), .QN(n2076) );
  DFFRX1 \i_MIPS/Register/register_reg[7][14]  ( .D(\i_MIPS/Register/n898 ), 
        .CK(clk), .RN(n5687), .Q(\i_MIPS/Register/register[7][14] ), .QN(n1903) );
  DFFRX1 \i_MIPS/Register/register_reg[7][16]  ( .D(\i_MIPS/Register/n900 ), 
        .CK(clk), .RN(n5688), .Q(\i_MIPS/Register/register[7][16] ), .QN(n2112) );
  DFFRX1 \i_MIPS/Register/register_reg[7][18]  ( .D(\i_MIPS/Register/n902 ), 
        .CK(clk), .RN(n5688), .Q(\i_MIPS/Register/register[7][18] ), .QN(n715)
         );
  DFFRX1 \i_MIPS/Register/register_reg[7][20]  ( .D(\i_MIPS/Register/n904 ), 
        .CK(clk), .RN(n5688), .Q(\i_MIPS/Register/register[7][20] ), .QN(n2111) );
  DFFRX1 \i_MIPS/Register/register_reg[7][21]  ( .D(\i_MIPS/Register/n905 ), 
        .CK(clk), .RN(n5688), .Q(\i_MIPS/Register/register[7][21] ), .QN(n2194) );
  DFFRX1 \i_MIPS/Register/register_reg[7][22]  ( .D(\i_MIPS/Register/n906 ), 
        .CK(clk), .RN(n5688), .Q(\i_MIPS/Register/register[7][22] ), .QN(n718)
         );
  DFFRX1 \i_MIPS/Register/register_reg[7][23]  ( .D(\i_MIPS/Register/n907 ), 
        .CK(clk), .RN(n5688), .Q(\i_MIPS/Register/register[7][23] ), .QN(n2087) );
  DFFRX1 \i_MIPS/Register/register_reg[7][24]  ( .D(\i_MIPS/Register/n908 ), 
        .CK(clk), .RN(n5688), .Q(\i_MIPS/Register/register[7][24] ), .QN(n2096) );
  DFFRX1 \i_MIPS/Register/register_reg[7][25]  ( .D(\i_MIPS/Register/n909 ), 
        .CK(clk), .RN(n5688), .Q(\i_MIPS/Register/register[7][25] ), .QN(n2079) );
  DFFRX1 \i_MIPS/Register/register_reg[7][26]  ( .D(\i_MIPS/Register/n910 ), 
        .CK(clk), .RN(n5688), .Q(\i_MIPS/Register/register[7][26] ), .QN(n2113) );
  DFFRX1 \i_MIPS/Register/register_reg[7][27]  ( .D(\i_MIPS/Register/n911 ), 
        .CK(clk), .RN(n5689), .Q(\i_MIPS/Register/register[7][27] ), .QN(n2088) );
  DFFRX1 \i_MIPS/Register/register_reg[7][28]  ( .D(\i_MIPS/Register/n912 ), 
        .CK(clk), .RN(n5689), .Q(\i_MIPS/Register/register[7][28] ), .QN(n2098) );
  DFFRX1 \i_MIPS/Register/register_reg[7][29]  ( .D(\i_MIPS/Register/n913 ), 
        .CK(clk), .RN(n5689), .Q(\i_MIPS/Register/register[7][29] ), .QN(n1901) );
  DFFRX1 \i_MIPS/Register/register_reg[5][2]  ( .D(\i_MIPS/Register/n950 ), 
        .CK(clk), .RN(n5692), .Q(\i_MIPS/Register/register[5][2] ), .QN(n2085)
         );
  DFFRX1 \i_MIPS/Register/register_reg[5][3]  ( .D(\i_MIPS/Register/n951 ), 
        .CK(clk), .RN(n5692), .Q(\i_MIPS/Register/register[5][3] ), .QN(n2101)
         );
  DFFRX1 \i_MIPS/Register/register_reg[5][4]  ( .D(\i_MIPS/Register/n952 ), 
        .CK(clk), .RN(n5692), .Q(\i_MIPS/Register/register[5][4] ), .QN(n1922)
         );
  DFFRX1 \i_MIPS/Register/register_reg[5][5]  ( .D(\i_MIPS/Register/n953 ), 
        .CK(clk), .RN(n5692), .Q(\i_MIPS/Register/register[5][5] ), .QN(n2281)
         );
  DFFRX1 \i_MIPS/Register/register_reg[5][6]  ( .D(\i_MIPS/Register/n954 ), 
        .CK(clk), .RN(n5692), .Q(\i_MIPS/Register/register[5][6] ), .QN(n2185)
         );
  DFFRX1 \i_MIPS/Register/register_reg[5][7]  ( .D(\i_MIPS/Register/n955 ), 
        .CK(clk), .RN(n5692), .Q(\i_MIPS/Register/register[5][7] ), .QN(n2245)
         );
  DFFRX1 \i_MIPS/Register/register_reg[5][8]  ( .D(\i_MIPS/Register/n956 ), 
        .CK(clk), .RN(n5692), .Q(\i_MIPS/Register/register[5][8] ), .QN(n2073)
         );
  DFFRX1 \i_MIPS/Register/register_reg[5][9]  ( .D(\i_MIPS/Register/n957 ), 
        .CK(clk), .RN(n5692), .Q(\i_MIPS/Register/register[5][9] ), .QN(n2069)
         );
  DFFRX1 \i_MIPS/Register/register_reg[5][10]  ( .D(\i_MIPS/Register/n958 ), 
        .CK(clk), .RN(n5692), .Q(\i_MIPS/Register/register[5][10] ), .QN(n1925) );
  DFFRX1 \i_MIPS/Register/register_reg[5][11]  ( .D(\i_MIPS/Register/n959 ), 
        .CK(clk), .RN(n5693), .Q(\i_MIPS/Register/register[5][11] ), .QN(n2117) );
  DFFRX1 \i_MIPS/Register/register_reg[5][12]  ( .D(\i_MIPS/Register/n960 ), 
        .CK(clk), .RN(n5693), .Q(\i_MIPS/Register/register[5][12] ), .QN(n2188) );
  DFFRX1 \i_MIPS/Register/register_reg[5][13]  ( .D(\i_MIPS/Register/n961 ), 
        .CK(clk), .RN(n5693), .Q(\i_MIPS/Register/register[5][13] ), .QN(n2077) );
  DFFRX1 \i_MIPS/Register/register_reg[5][14]  ( .D(\i_MIPS/Register/n962 ), 
        .CK(clk), .RN(n5693), .Q(\i_MIPS/Register/register[5][14] ), .QN(n1915) );
  DFFRX1 \i_MIPS/Register/register_reg[5][15]  ( .D(\i_MIPS/Register/n963 ), 
        .CK(clk), .RN(n5693), .Q(\i_MIPS/Register/register[5][15] ), .QN(n2280) );
  DFFRX1 \i_MIPS/Register/register_reg[5][16]  ( .D(\i_MIPS/Register/n964 ), 
        .CK(clk), .RN(n5693), .Q(\i_MIPS/Register/register[5][16] ), .QN(n2244) );
  DFFRX1 \i_MIPS/Register/register_reg[5][17]  ( .D(\i_MIPS/Register/n965 ), 
        .CK(clk), .RN(n5693), .Q(\i_MIPS/Register/register[5][17] ), .QN(n2232) );
  DFFRX1 \i_MIPS/Register/register_reg[5][18]  ( .D(\i_MIPS/Register/n966 ), 
        .CK(clk), .RN(n5693), .Q(\i_MIPS/Register/register[5][18] ), .QN(n1998) );
  DFFRX1 \i_MIPS/Register/register_reg[5][20]  ( .D(\i_MIPS/Register/n968 ), 
        .CK(clk), .RN(n5693), .Q(\i_MIPS/Register/register[5][20] ), .QN(n2242) );
  DFFRX1 \i_MIPS/Register/register_reg[5][21]  ( .D(\i_MIPS/Register/n969 ), 
        .CK(clk), .RN(n5693), .Q(\i_MIPS/Register/register[5][21] ), .QN(n2277) );
  DFFRX1 \i_MIPS/Register/register_reg[5][22]  ( .D(\i_MIPS/Register/n970 ), 
        .CK(clk), .RN(n5693), .Q(\i_MIPS/Register/register[5][22] ), .QN(n1997) );
  DFFRX1 \i_MIPS/Register/register_reg[5][23]  ( .D(\i_MIPS/Register/n971 ), 
        .CK(clk), .RN(n5694), .Q(\i_MIPS/Register/register[5][23] ), .QN(n2241) );
  DFFRX1 \i_MIPS/Register/register_reg[5][24]  ( .D(\i_MIPS/Register/n972 ), 
        .CK(clk), .RN(n5694), .Q(\i_MIPS/Register/register[5][24] ), .QN(n2097) );
  DFFRX1 \i_MIPS/Register/register_reg[5][25]  ( .D(\i_MIPS/Register/n973 ), 
        .CK(clk), .RN(n5694), .Q(\i_MIPS/Register/register[5][25] ), .QN(n2239) );
  DFFRX1 \i_MIPS/Register/register_reg[5][26]  ( .D(\i_MIPS/Register/n974 ), 
        .CK(clk), .RN(n5694), .Q(\i_MIPS/Register/register[5][26] ), .QN(n2115) );
  DFFRX1 \i_MIPS/Register/register_reg[5][27]  ( .D(\i_MIPS/Register/n975 ), 
        .CK(clk), .RN(n5694), .Q(\i_MIPS/Register/register[5][27] ), .QN(n2089) );
  DFFRX1 \i_MIPS/Register/register_reg[5][28]  ( .D(\i_MIPS/Register/n976 ), 
        .CK(clk), .RN(n5694), .Q(\i_MIPS/Register/register[5][28] ), .QN(n2099) );
  DFFRX1 \i_MIPS/Register/register_reg[5][29]  ( .D(\i_MIPS/Register/n977 ), 
        .CK(clk), .RN(n5694), .Q(\i_MIPS/Register/register[5][29] ), .QN(n1913) );
  DFFRX1 \i_MIPS/Register/register_reg[5][31]  ( .D(\i_MIPS/Register/n979 ), 
        .CK(clk), .RN(n5694), .Q(\i_MIPS/Register/register[5][31] ), .QN(n2183) );
  DFFRX1 \i_MIPS/Register/register_reg[4][3]  ( .D(\i_MIPS/Register/n983 ), 
        .CK(clk), .RN(n5695), .Q(\i_MIPS/Register/register[4][3] ), .QN(n2162)
         );
  DFFRX1 \i_MIPS/Register/register_reg[4][16]  ( .D(\i_MIPS/Register/n996 ), 
        .CK(clk), .RN(n5696), .Q(\i_MIPS/Register/register[4][16] ), .QN(n1906) );
  DFFRX1 \i_MIPS/Register/register_reg[4][22]  ( .D(\i_MIPS/Register/n1002 ), 
        .CK(clk), .RN(n5696), .Q(\i_MIPS/Register/register[4][22] ), .QN(n2161) );
  DFFRX1 \i_MIPS/Register/register_reg[4][23]  ( .D(\i_MIPS/Register/n1003 ), 
        .CK(clk), .RN(n5696), .Q(\i_MIPS/Register/register[4][23] ), .QN(n1905) );
  DFFRX1 \i_MIPS/Register/register_reg[4][24]  ( .D(\i_MIPS/Register/n1004 ), 
        .CK(clk), .RN(n5696), .Q(\i_MIPS/Register/register[4][24] ), .QN(n2160) );
  DFFRX1 \i_MIPS/Register/register_reg[3][2]  ( .D(\i_MIPS/Register/n1014 ), 
        .CK(clk), .RN(n5697), .Q(\i_MIPS/Register/register[3][2] ), .QN(n2084)
         );
  DFFRX1 \i_MIPS/Register/register_reg[3][3]  ( .D(\i_MIPS/Register/n1015 ), 
        .CK(clk), .RN(n5697), .Q(\i_MIPS/Register/register[3][3] ), .QN(n2256)
         );
  DFFRX1 \i_MIPS/Register/register_reg[3][4]  ( .D(\i_MIPS/Register/n1016 ), 
        .CK(clk), .RN(n5697), .Q(\i_MIPS/Register/register[3][4] ), .QN(n2110)
         );
  DFFRX1 \i_MIPS/Register/register_reg[3][5]  ( .D(\i_MIPS/Register/n1017 ), 
        .CK(clk), .RN(n5697), .Q(\i_MIPS/Register/register[3][5] ), .QN(n2297)
         );
  DFFRX1 \i_MIPS/Register/register_reg[3][6]  ( .D(\i_MIPS/Register/n1018 ), 
        .CK(clk), .RN(n5697), .Q(\i_MIPS/Register/register[3][6] ), .QN(n2283)
         );
  DFFRX1 \i_MIPS/Register/register_reg[3][7]  ( .D(\i_MIPS/Register/n1019 ), 
        .CK(clk), .RN(n5698), .Q(\i_MIPS/Register/register[3][7] ), .QN(n2287)
         );
  DFFRX1 \i_MIPS/Register/register_reg[3][8]  ( .D(\i_MIPS/Register/n1020 ), 
        .CK(clk), .RN(n5698), .Q(\i_MIPS/Register/register[3][8] ), .QN(n2252)
         );
  DFFRX1 \i_MIPS/Register/register_reg[3][9]  ( .D(\i_MIPS/Register/n1021 ), 
        .CK(clk), .RN(n5698), .Q(\i_MIPS/Register/register[3][9] ), .QN(n2248)
         );
  DFFRX1 \i_MIPS/Register/register_reg[3][10]  ( .D(\i_MIPS/Register/n1022 ), 
        .CK(clk), .RN(n5698), .Q(\i_MIPS/Register/register[3][10] ), .QN(n2259) );
  DFFRX1 \i_MIPS/Register/register_reg[3][11]  ( .D(\i_MIPS/Register/n1023 ), 
        .CK(clk), .RN(n5698), .Q(\i_MIPS/Register/register[3][11] ), .QN(n2261) );
  DFFRX1 \i_MIPS/Register/register_reg[3][12]  ( .D(\i_MIPS/Register/n1024 ), 
        .CK(clk), .RN(n5698), .Q(\i_MIPS/Register/register[3][12] ), .QN(n2291) );
  DFFRX1 \i_MIPS/Register/register_reg[3][13]  ( .D(\i_MIPS/Register/n1025 ), 
        .CK(clk), .RN(n5698), .Q(\i_MIPS/Register/register[3][13] ), .QN(n2058) );
  DFFRX1 \i_MIPS/Register/register_reg[3][14]  ( .D(\i_MIPS/Register/n1026 ), 
        .CK(clk), .RN(n5698), .Q(\i_MIPS/Register/register[3][14] ), .QN(n2250) );
  DFFRX1 \i_MIPS/Register/register_reg[3][15]  ( .D(\i_MIPS/Register/n1027 ), 
        .CK(clk), .RN(n5698), .Q(\i_MIPS/Register/register[3][15] ), .QN(n2293) );
  DFFRX1 \i_MIPS/Register/register_reg[3][16]  ( .D(\i_MIPS/Register/n1028 ), 
        .CK(clk), .RN(n5698), .Q(\i_MIPS/Register/register[3][16] ), .QN(n2260) );
  DFFRX1 \i_MIPS/Register/register_reg[3][17]  ( .D(\i_MIPS/Register/n1029 ), 
        .CK(clk), .RN(n5698), .Q(\i_MIPS/Register/register[3][17] ), .QN(n2247) );
  DFFRX1 \i_MIPS/Register/register_reg[3][18]  ( .D(\i_MIPS/Register/n1030 ), 
        .CK(clk), .RN(n5698), .Q(\i_MIPS/Register/register[3][18] ), .QN(n2289) );
  DFFRX1 \i_MIPS/Register/register_reg[3][20]  ( .D(\i_MIPS/Register/n1032 ), 
        .CK(clk), .RN(n5699), .Q(\i_MIPS/Register/register[3][20] ), .QN(n2056) );
  DFFRX1 \i_MIPS/Register/register_reg[3][21]  ( .D(\i_MIPS/Register/n1033 ), 
        .CK(clk), .RN(n5699), .Q(\i_MIPS/Register/register[3][21] ), .QN(n2285) );
  DFFRX1 \i_MIPS/Register/register_reg[3][22]  ( .D(\i_MIPS/Register/n1034 ), 
        .CK(clk), .RN(n5699), .Q(\i_MIPS/Register/register[3][22] ), .QN(n2104) );
  DFFRX1 \i_MIPS/Register/register_reg[3][23]  ( .D(\i_MIPS/Register/n1035 ), 
        .CK(clk), .RN(n5699), .Q(\i_MIPS/Register/register[3][23] ), .QN(n2254) );
  DFFRX1 \i_MIPS/Register/register_reg[3][24]  ( .D(\i_MIPS/Register/n1036 ), 
        .CK(clk), .RN(n5699), .Q(\i_MIPS/Register/register[3][24] ), .QN(n2295) );
  DFFRX1 \i_MIPS/Register/register_reg[3][25]  ( .D(\i_MIPS/Register/n1037 ), 
        .CK(clk), .RN(n5699), .Q(\i_MIPS/Register/register[3][25] ), .QN(n2055) );
  DFFRX1 \i_MIPS/Register/register_reg[3][26]  ( .D(\i_MIPS/Register/n1038 ), 
        .CK(clk), .RN(n5699), .Q(\i_MIPS/Register/register[3][26] ), .QN(n2114) );
  DFFRX1 \i_MIPS/Register/register_reg[3][27]  ( .D(\i_MIPS/Register/n1039 ), 
        .CK(clk), .RN(n5699), .Q(\i_MIPS/Register/register[3][27] ), .QN(n2296) );
  DFFRX1 \i_MIPS/Register/register_reg[3][28]  ( .D(\i_MIPS/Register/n1040 ), 
        .CK(clk), .RN(n5699), .Q(\i_MIPS/Register/register[3][28] ), .QN(n2196) );
  DFFRX1 \i_MIPS/Register/register_reg[3][29]  ( .D(\i_MIPS/Register/n1041 ), 
        .CK(clk), .RN(n5699), .Q(\i_MIPS/Register/register[3][29] ), .QN(n1926) );
  DFFRX1 \i_MIPS/Register/register_reg[3][31]  ( .D(\i_MIPS/Register/n1043 ), 
        .CK(clk), .RN(n5700), .Q(\i_MIPS/Register/register[3][31] ), .QN(n2299) );
  DFFRX1 \i_MIPS/Register/register_reg[1][2]  ( .D(\i_MIPS/Register/n1078 ), 
        .CK(clk), .RN(n5702), .Q(\i_MIPS/Register/register[1][2] ), .QN(n2034)
         );
  DFFRX1 \i_MIPS/Register/register_reg[1][3]  ( .D(\i_MIPS/Register/n1079 ), 
        .CK(clk), .RN(n5703), .Q(\i_MIPS/Register/register[1][3] ), .QN(n2065)
         );
  DFFRX1 \i_MIPS/Register/register_reg[1][4]  ( .D(\i_MIPS/Register/n1080 ), 
        .CK(clk), .RN(n5703), .Q(\i_MIPS/Register/register[1][4] ), .QN(n2037)
         );
  DFFRX1 \i_MIPS/Register/register_reg[1][5]  ( .D(\i_MIPS/Register/n1081 ), 
        .CK(clk), .RN(n5703), .Q(\i_MIPS/Register/register[1][5] ), .QN(n2179)
         );
  DFFRX1 \i_MIPS/Register/register_reg[1][6]  ( .D(\i_MIPS/Register/n1082 ), 
        .CK(clk), .RN(n5703), .Q(\i_MIPS/Register/register[1][6] ), .QN(n2269)
         );
  DFFRX1 \i_MIPS/Register/register_reg[1][7]  ( .D(\i_MIPS/Register/n1083 ), 
        .CK(clk), .RN(n5703), .Q(\i_MIPS/Register/register[1][7] ), .QN(n2275)
         );
  DFFRX1 \i_MIPS/Register/register_reg[1][8]  ( .D(\i_MIPS/Register/n1084 ), 
        .CK(clk), .RN(n5703), .Q(\i_MIPS/Register/register[1][8] ), .QN(n2313)
         );
  DFFRX1 \i_MIPS/Register/register_reg[1][9]  ( .D(\i_MIPS/Register/n1085 ), 
        .CK(clk), .RN(n5703), .Q(\i_MIPS/Register/register[1][9] ), .QN(n2311)
         );
  DFFRX1 \i_MIPS/Register/register_reg[1][10]  ( .D(\i_MIPS/Register/n1086 ), 
        .CK(clk), .RN(n5703), .Q(\i_MIPS/Register/register[1][10] ), .QN(n2237) );
  DFFRX1 \i_MIPS/Register/register_reg[1][11]  ( .D(\i_MIPS/Register/n1087 ), 
        .CK(clk), .RN(n5703), .Q(\i_MIPS/Register/register[1][11] ), .QN(n2274) );
  DFFRX1 \i_MIPS/Register/register_reg[1][12]  ( .D(\i_MIPS/Register/n1088 ), 
        .CK(clk), .RN(n5703), .Q(\i_MIPS/Register/register[1][12] ), .QN(n2309) );
  DFFRX1 \i_MIPS/Register/register_reg[1][13]  ( .D(\i_MIPS/Register/n1089 ), 
        .CK(clk), .RN(n5703), .Q(\i_MIPS/Register/register[1][13] ), .QN(n2307) );
  DFFRX1 \i_MIPS/Register/register_reg[1][14]  ( .D(\i_MIPS/Register/n1090 ), 
        .CK(clk), .RN(n5703), .Q(\i_MIPS/Register/register[1][14] ), .QN(n2171) );
  DFFRX1 \i_MIPS/Register/register_reg[1][15]  ( .D(\i_MIPS/Register/n1091 ), 
        .CK(clk), .RN(n5704), .Q(\i_MIPS/Register/register[1][15] ), .QN(n2271) );
  DFFRX1 \i_MIPS/Register/register_reg[1][16]  ( .D(\i_MIPS/Register/n1092 ), 
        .CK(clk), .RN(n5704), .Q(\i_MIPS/Register/register[1][16] ), .QN(n2264) );
  DFFRX1 \i_MIPS/Register/register_reg[1][17]  ( .D(\i_MIPS/Register/n1093 ), 
        .CK(clk), .RN(n5704), .Q(\i_MIPS/Register/register[1][17] ), .QN(n2061) );
  DFFRX1 \i_MIPS/Register/register_reg[1][18]  ( .D(\i_MIPS/Register/n1094 ), 
        .CK(clk), .RN(n5704), .Q(\i_MIPS/Register/register[1][18] ), .QN(n1910) );
  DFFRX1 \i_MIPS/Register/register_reg[1][20]  ( .D(\i_MIPS/Register/n1096 ), 
        .CK(clk), .RN(n5704), .Q(\i_MIPS/Register/register[1][20] ), .QN(n2169) );
  DFFRX1 \i_MIPS/Register/register_reg[1][21]  ( .D(\i_MIPS/Register/n1097 ), 
        .CK(clk), .RN(n5704), .Q(\i_MIPS/Register/register[1][21] ), .QN(n2301) );
  DFFRX1 \i_MIPS/Register/register_reg[1][22]  ( .D(\i_MIPS/Register/n1098 ), 
        .CK(clk), .RN(n5704), .Q(\i_MIPS/Register/register[1][22] ), .QN(n1912) );
  DFFRX1 \i_MIPS/Register/register_reg[1][23]  ( .D(\i_MIPS/Register/n1099 ), 
        .CK(clk), .RN(n5704), .Q(\i_MIPS/Register/register[1][23] ), .QN(n2262) );
  DFFRX1 \i_MIPS/Register/register_reg[1][24]  ( .D(\i_MIPS/Register/n1100 ), 
        .CK(clk), .RN(n5704), .Q(\i_MIPS/Register/register[1][24] ), .QN(n2064) );
  DFFRX1 \i_MIPS/Register/register_reg[1][25]  ( .D(\i_MIPS/Register/n1101 ), 
        .CK(clk), .RN(n5704), .Q(\i_MIPS/Register/register[1][25] ), .QN(n2303) );
  DFFRX1 \i_MIPS/Register/register_reg[1][26]  ( .D(\i_MIPS/Register/n1102 ), 
        .CK(clk), .RN(n5704), .Q(\i_MIPS/Register/register[1][26] ), .QN(n2221) );
  DFFRX1 \i_MIPS/Register/register_reg[1][27]  ( .D(\i_MIPS/Register/n1103 ), 
        .CK(clk), .RN(n5705), .Q(\i_MIPS/Register/register[1][27] ), .QN(n2177) );
  DFFRX1 \i_MIPS/Register/register_reg[1][28]  ( .D(\i_MIPS/Register/n1104 ), 
        .CK(clk), .RN(n5705), .Q(\i_MIPS/Register/register[1][28] ), .QN(n2062) );
  DFFRX1 \i_MIPS/Register/register_reg[1][29]  ( .D(\i_MIPS/Register/n1105 ), 
        .CK(clk), .RN(n5705), .Q(\i_MIPS/Register/register[1][29] ), .QN(n2038) );
  DFFRX1 \i_MIPS/Register/register_reg[1][31]  ( .D(\i_MIPS/Register/n1107 ), 
        .CK(clk), .RN(n5705), .Q(\i_MIPS/Register/register[1][31] ), .QN(n2174) );
  DFFRX1 \i_MIPS/Register/register_reg[0][2]  ( .D(\i_MIPS/Register/n1110 ), 
        .CK(clk), .RN(n5705), .Q(\i_MIPS/Register/register[0][2] ), .QN(n2147)
         );
  DFFRX1 \i_MIPS/Register/register_reg[0][3]  ( .D(\i_MIPS/Register/n1111 ), 
        .CK(clk), .RN(n5705), .Q(\i_MIPS/Register/register[0][3] ), .QN(n2141)
         );
  DFFRX1 \i_MIPS/Register/register_reg[0][16]  ( .D(\i_MIPS/Register/n1124 ), 
        .CK(clk), .RN(n5706), .Q(\i_MIPS/Register/register[0][16] ), .QN(n2135) );
  DFFRX1 \i_MIPS/Register/register_reg[0][20]  ( .D(\i_MIPS/Register/n1128 ), 
        .CK(clk), .RN(n5707), .Q(\i_MIPS/Register/register[0][20] ), .QN(n2144) );
  DFFRX1 \i_MIPS/Register/register_reg[0][21]  ( .D(\i_MIPS/Register/n1129 ), 
        .CK(clk), .RN(n5707), .Q(\i_MIPS/Register/register[0][21] ), .QN(n2145) );
  DFFRX1 \i_MIPS/Register/register_reg[0][22]  ( .D(\i_MIPS/Register/n1130 ), 
        .CK(clk), .RN(n5707), .Q(\i_MIPS/Register/register[0][22] ), .QN(n2139) );
  DFFRX1 \i_MIPS/Register/register_reg[0][23]  ( .D(\i_MIPS/Register/n1131 ), 
        .CK(clk), .RN(n5707), .Q(\i_MIPS/Register/register[0][23] ), .QN(n2137) );
  DFFRX1 \i_MIPS/Register/register_reg[0][24]  ( .D(\i_MIPS/Register/n1132 ), 
        .CK(clk), .RN(n5707), .Q(\i_MIPS/Register/register[0][24] ), .QN(n2133) );
  DFFRX1 \i_MIPS/Register/register_reg[26][3]  ( .D(\i_MIPS/Register/n279 ), 
        .CK(clk), .RN(n5636), .Q(\i_MIPS/Register/register[26][3] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][16]  ( .D(\i_MIPS/Register/n292 ), 
        .CK(clk), .RN(n5637), .Q(\i_MIPS/Register/register[26][16] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][3]  ( .D(\i_MIPS/Register/n791 ), 
        .CK(clk), .RN(n5679), .Q(\i_MIPS/Register/register[10][3] ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[0]  ( .D(\i_MIPS/n563 ), .CK(clk), .RN(n5619), .Q(
        \i_MIPS/EX_MEM_0 ), .QN(\i_MIPS/n373 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[35]  ( .D(\i_MIPS/n536 ), .CK(clk), .RN(n5617), .Q(
        \i_MIPS/ALUin1[26] ), .QN(\i_MIPS/n345 ) );
  DFFRX2 \i_MIPS/EX_MEM_reg[1]  ( .D(\i_MIPS/n526 ), .CK(clk), .RN(n5616), .Q(
        \i_MIPS/EX_MEM_1 ), .QN(\i_MIPS/n336 ) );
  DFFRX2 \i_MIPS/EX_MEM_reg[72]  ( .D(\i_MIPS/n474 ), .CK(clk), .RN(n5609), 
        .Q(\i_MIPS/Reg_W[3] ), .QN(n4716) );
  DFFRX2 \i_MIPS/EX_MEM_reg[69]  ( .D(\i_MIPS/n477 ), .CK(clk), .RN(n5610), 
        .Q(\i_MIPS/Reg_W[0] ), .QN(n287) );
  DFFRX2 \i_MIPS/EX_MEM_reg[70]  ( .D(\i_MIPS/n476 ), .CK(clk), .RN(n5610), 
        .Q(\i_MIPS/Reg_W[1] ), .QN(n229) );
  DFFRX2 \i_MIPS/EX_MEM_reg[71]  ( .D(\i_MIPS/n475 ), .CK(clk), .RN(n5609), 
        .Q(\i_MIPS/Reg_W[2] ), .QN(n4705) );
  DFFRX1 \I_cache/cache_reg[3][137]  ( .D(n11724), .CK(clk), .RN(n5902), .Q(
        \I_cache/cache[3][137] ), .QN(n3268) );
  DFFRX1 \I_cache/cache_reg[4][142]  ( .D(n11683), .CK(clk), .RN(n5906), .Q(
        \I_cache/cache[4][142] ), .QN(n4497) );
  DFFRHQX8 \i_MIPS/PC/PC_o_reg[4]  ( .D(\i_MIPS/PC/n38 ), .CK(clk), .RN(n5620), 
        .Q(n4502) );
  DFFRX1 \I_cache/cache_reg[5][137]  ( .D(n11722), .CK(clk), .RN(n5903), .Q(
        \I_cache/cache[5][137] ), .QN(n3210) );
  DFFRX1 \I_cache/cache_reg[4][141]  ( .D(n11691), .CK(clk), .RN(n5905), .Q(
        \I_cache/cache[4][141] ), .QN(n1600) );
  DFFRX1 \I_cache/cache_reg[2][143]  ( .D(n11677), .CK(clk), .RN(n5906), .Q(
        \I_cache/cache[2][143] ), .QN(n1611) );
  DFFRX1 \I_cache/cache_reg[4][149]  ( .D(n11627), .CK(clk), .RN(n5911), .Q(
        \I_cache/cache[4][149] ) );
  DFFRX1 \I_cache/cache_reg[4][152]  ( .D(n11603), .CK(clk), .RN(n5913), .Q(
        \I_cache/cache[4][152] ) );
  DFFRX1 \I_cache/cache_reg[6][133]  ( .D(n11753), .CK(clk), .RN(n5900), .Q(
        \I_cache/cache[6][133] ), .QN(n1940) );
  DFFRX1 \I_cache/cache_reg[6][138]  ( .D(n11713), .CK(clk), .RN(n5903), .Q(
        \I_cache/cache[6][138] ), .QN(n1944) );
  DFFRX1 \I_cache/cache_reg[7][145]  ( .D(n11656), .CK(clk), .RN(n5908), .Q(
        \I_cache/cache[7][145] ), .QN(n364) );
  DFFRX1 \I_cache/cache_reg[1][148]  ( .D(n11638), .CK(clk), .RN(n5910), .Q(
        \I_cache/cache[1][148] ), .QN(n396) );
  DFFRX1 \I_cache/cache_reg[3][148]  ( .D(n11636), .CK(clk), .RN(n5910), .Q(
        \I_cache/cache[3][148] ), .QN(n397) );
  DFFRX1 \I_cache/cache_reg[0][132]  ( .D(n11767), .CK(clk), .RN(n5899), .Q(
        \I_cache/cache[0][132] ), .QN(n3200) );
  DFFRX1 \I_cache/cache_reg[2][132]  ( .D(n11765), .CK(clk), .RN(n5899), .Q(
        \I_cache/cache[2][132] ), .QN(n3201) );
  DFFRX1 \I_cache/cache_reg[7][133]  ( .D(n11752), .CK(clk), .RN(n5900), .Q(
        \I_cache/cache[7][133] ), .QN(n362) );
  DFFRHQX8 \i_MIPS/EX_MEM_reg[10]  ( .D(\i_MIPS/n464 ), .CK(clk), .RN(n5609), 
        .Q(net138398) );
  DFFRX1 \I_cache/cache_reg[0][128]  ( .D(n11799), .CK(clk), .RN(n5896), .Q(
        \I_cache/cache[0][128] ), .QN(n3228) );
  DFFRX1 \I_cache/cache_reg[2][128]  ( .D(n11797), .CK(clk), .RN(n5896), .Q(
        \I_cache/cache[2][128] ), .QN(n3229) );
  DFFRX1 \I_cache/cache_reg[0][129]  ( .D(n11791), .CK(clk), .RN(n5897), .Q(
        \I_cache/cache[0][129] ), .QN(n3225) );
  DFFRX1 \I_cache/cache_reg[1][135]  ( .D(n11742), .CK(clk), .RN(n5901), .Q(
        \I_cache/cache[1][135] ), .QN(n1593) );
  DFFRX1 \I_cache/cache_reg[3][135]  ( .D(n11740), .CK(clk), .RN(n5901), .Q(
        \I_cache/cache[3][135] ), .QN(n1594) );
  DFFRX1 \I_cache/cache_reg[5][135]  ( .D(n11738), .CK(clk), .RN(n5901), .Q(
        \I_cache/cache[5][135] ), .QN(n3209) );
  DFFRX1 \I_cache/cache_reg[6][135]  ( .D(n11737), .CK(clk), .RN(n5901), .Q(
        \I_cache/cache[6][135] ), .QN(n1606) );
  DFFRX1 \I_cache/cache_reg[2][136]  ( .D(n11733), .CK(clk), .RN(n5902), .Q(
        \I_cache/cache[2][136] ), .QN(n3236) );
  DFFRX1 \I_cache/cache_reg[3][136]  ( .D(n11732), .CK(clk), .RN(n5902), .Q(
        \I_cache/cache[3][136] ), .QN(n1598) );
  DFFRX1 \I_cache/cache_reg[6][136]  ( .D(n11729), .CK(clk), .RN(n5902), .Q(
        \I_cache/cache[6][136] ), .QN(n1607) );
  DFFRX1 \I_cache/cache_reg[0][139]  ( .D(n11711), .CK(clk), .RN(n5904), .Q(
        \I_cache/cache[0][139] ), .QN(n3234) );
  DFFRX1 \I_cache/cache_reg[1][140]  ( .D(n11702), .CK(clk), .RN(n5904), .Q(
        \I_cache/cache[1][140] ), .QN(n1591) );
  DFFRX1 \I_cache/cache_reg[3][140]  ( .D(n11700), .CK(clk), .RN(n5904), .Q(
        \I_cache/cache[3][140] ), .QN(n1592) );
  DFFRX1 \I_cache/cache_reg[5][140]  ( .D(n11698), .CK(clk), .RN(n5905), .Q(
        \I_cache/cache[5][140] ), .QN(n3208) );
  DFFRX1 \I_cache/cache_reg[6][140]  ( .D(n11697), .CK(clk), .RN(n5905), .Q(
        \I_cache/cache[6][140] ), .QN(n1605) );
  DFFRX1 \I_cache/cache_reg[0][141]  ( .D(n11695), .CK(clk), .RN(n5905), .Q(
        \I_cache/cache[0][141] ), .QN(n3223) );
  DFFRX1 \I_cache/cache_reg[1][141]  ( .D(n11694), .CK(clk), .RN(n5905), .Q(
        \I_cache/cache[1][141] ), .QN(n1584) );
  DFFRX1 \I_cache/cache_reg[2][141]  ( .D(n11693), .CK(clk), .RN(n5905), .Q(
        \I_cache/cache[2][141] ), .QN(n3224) );
  DFFRX1 \I_cache/cache_reg[3][141]  ( .D(n11692), .CK(clk), .RN(n5905), .Q(
        \I_cache/cache[3][141] ), .QN(n1585) );
  DFFRX1 \I_cache/cache_reg[6][141]  ( .D(n11689), .CK(clk), .RN(n5905), .Q(
        \I_cache/cache[6][141] ), .QN(n3237) );
  DFFRX1 \I_cache/cache_reg[7][141]  ( .D(n11688), .CK(clk), .RN(n5905), .Q(
        \I_cache/cache[7][141] ), .QN(n1599) );
  DFFRX1 \I_cache/cache_reg[5][142]  ( .D(n11682), .CK(clk), .RN(n5906), .Q(
        \I_cache/cache[5][142] ), .QN(n3205) );
  DFFRX1 \I_cache/cache_reg[1][143]  ( .D(n11678), .CK(clk), .RN(n5906), .Q(
        \I_cache/cache[1][143] ), .QN(n3241) );
  DFFRX1 \I_cache/cache_reg[3][143]  ( .D(n11676), .CK(clk), .RN(n5906), .Q(
        \I_cache/cache[3][143] ), .QN(n3242) );
  DFFRX1 \I_cache/cache_reg[6][143]  ( .D(n11673), .CK(clk), .RN(n5907), .Q(
        \I_cache/cache[6][143] ), .QN(n1612) );
  DFFRX1 \I_cache/cache_reg[0][147]  ( .D(n11647), .CK(clk), .RN(n5909), .Q(
        \I_cache/cache[0][147] ), .QN(n3232) );
  DFFRX1 \I_cache/cache_reg[1][147]  ( .D(n11646), .CK(clk), .RN(n5909), .Q(
        \I_cache/cache[1][147] ), .QN(n1595) );
  DFFRX1 \I_cache/cache_reg[2][147]  ( .D(n11645), .CK(clk), .RN(n5909), .Q(
        \I_cache/cache[2][147] ), .QN(n3233) );
  DFFRX1 \I_cache/cache_reg[3][147]  ( .D(n11644), .CK(clk), .RN(n5909), .Q(
        \I_cache/cache[3][147] ), .QN(n1596) );
  DFFRX1 \I_cache/cache_reg[5][147]  ( .D(n11642), .CK(clk), .RN(n5909), .Q(
        \I_cache/cache[5][147] ), .QN(n3216) );
  DFFRX1 \I_cache/cache_reg[6][147]  ( .D(n11641), .CK(clk), .RN(n5909), .Q(
        \I_cache/cache[6][147] ), .QN(n3235) );
  DFFRX1 \I_cache/cache_reg[7][147]  ( .D(n11640), .CK(clk), .RN(n5909), .Q(
        \I_cache/cache[7][147] ), .QN(n1597) );
  DFFRX1 \I_cache/cache_reg[0][149]  ( .D(n11631), .CK(clk), .RN(n5910), .Q(
        \I_cache/cache[0][149] ), .QN(n3226) );
  DFFRX1 \I_cache/cache_reg[1][149]  ( .D(n11630), .CK(clk), .RN(n5910), .Q(
        \I_cache/cache[1][149] ), .QN(n1587) );
  DFFRX1 \I_cache/cache_reg[2][149]  ( .D(n11629), .CK(clk), .RN(n5910), .Q(
        \I_cache/cache[2][149] ), .QN(n3227) );
  DFFRX1 \I_cache/cache_reg[3][149]  ( .D(n11628), .CK(clk), .RN(n5910), .Q(
        \I_cache/cache[3][149] ), .QN(n1588) );
  DFFRX1 \I_cache/cache_reg[5][149]  ( .D(n11626), .CK(clk), .RN(n5911), .Q(
        \I_cache/cache[5][149] ), .QN(n3217) );
  DFFRX1 \I_cache/cache_reg[6][149]  ( .D(n11625), .CK(clk), .RN(n5911), .Q(
        \I_cache/cache[6][149] ), .QN(n1601) );
  DFFRX1 \I_cache/cache_reg[0][151]  ( .D(n11615), .CK(clk), .RN(n5912), .Q(
        \I_cache/cache[0][151] ), .QN(n1603) );
  DFFRX1 \I_cache/cache_reg[2][151]  ( .D(n11613), .CK(clk), .RN(n5912), .Q(
        \I_cache/cache[2][151] ), .QN(n1604) );
  DFFRX1 \I_cache/cache_reg[0][152]  ( .D(n11607), .CK(clk), .RN(n5912), .Q(
        \I_cache/cache[0][152] ), .QN(n3230) );
  DFFRX1 \I_cache/cache_reg[1][152]  ( .D(n11606), .CK(clk), .RN(n5912), .Q(
        \I_cache/cache[1][152] ), .QN(n1589) );
  DFFRX1 \I_cache/cache_reg[2][152]  ( .D(n11605), .CK(clk), .RN(n5912), .Q(
        \I_cache/cache[2][152] ), .QN(n3231) );
  DFFRX1 \I_cache/cache_reg[3][152]  ( .D(n11604), .CK(clk), .RN(n5912), .Q(
        \I_cache/cache[3][152] ), .QN(n1590) );
  DFFRX1 \I_cache/cache_reg[5][152]  ( .D(n11602), .CK(clk), .RN(n5913), .Q(
        \I_cache/cache[5][152] ), .QN(n3212) );
  DFFRX1 \I_cache/cache_reg[6][152]  ( .D(n11601), .CK(clk), .RN(n5913), .Q(
        \I_cache/cache[6][152] ), .QN(n1602) );
  DFFRX1 \I_cache/cache_reg[4][154]  ( .D(n11587), .CK(clk), .RN(n5914), .Q(
        \I_cache/cache[4][154] ), .QN(n3207) );
  DFFRX1 \I_cache/cache_reg[7][135]  ( .D(n11736), .CK(clk), .RN(n5901), .Q(
        \I_cache/cache[7][135] ), .QN(n3272) );
  DFFRX1 \I_cache/cache_reg[7][136]  ( .D(n11728), .CK(clk), .RN(n5902), .Q(
        \I_cache/cache[7][136] ), .QN(n3273) );
  DFFRX1 \I_cache/cache_reg[7][137]  ( .D(n11720), .CK(clk), .RN(n5903), .Q(
        \I_cache/cache[7][137] ), .QN(n3271) );
  DFFRX1 \I_cache/cache_reg[7][140]  ( .D(n11696), .CK(clk), .RN(n5905), .Q(
        \I_cache/cache[7][140] ), .QN(n3269) );
  DFFRX1 \I_cache/cache_reg[5][141]  ( .D(n11690), .CK(clk), .RN(n5905), .Q(
        \I_cache/cache[5][141] ), .QN(n3260) );
  DFFRX1 \I_cache/cache_reg[6][142]  ( .D(n11681), .CK(clk), .RN(n5906), .Q(
        \I_cache/cache[6][142] ), .QN(n1627) );
  DFFRX1 \I_cache/cache_reg[5][143]  ( .D(n11674), .CK(clk), .RN(n5907), .Q(
        \I_cache/cache[5][143] ), .QN(n1621) );
  DFFRX1 \I_cache/cache_reg[7][143]  ( .D(n11672), .CK(clk), .RN(n5907), .Q(
        \I_cache/cache[7][143] ), .QN(n3294) );
  DFFRX1 \I_cache/cache_reg[7][144]  ( .D(n11664), .CK(clk), .RN(n5907), .Q(
        \I_cache/cache[7][144] ), .QN(n3270) );
  DFFRX1 \I_cache/cache_reg[7][148]  ( .D(n11632), .CK(clk), .RN(n5910), .Q(
        \I_cache/cache[7][148] ), .QN(n3266) );
  DFFRX1 \I_cache/cache_reg[7][149]  ( .D(n11624), .CK(clk), .RN(n5911), .Q(
        \I_cache/cache[7][149] ), .QN(n3265) );
  DFFRX1 \I_cache/cache_reg[7][152]  ( .D(n11600), .CK(clk), .RN(n5913), .Q(
        \I_cache/cache[7][152] ), .QN(n3267) );
  DFFRX1 \I_cache/cache_reg[0][154]  ( .D(n11591), .CK(clk), .RN(n5914), .Q(
        \I_cache/cache[0][154] ), .QN(n3298) );
  DFFRX1 \I_cache/cache_reg[1][154]  ( .D(n11590), .CK(clk), .RN(n5914), .Q(
        \I_cache/cache[1][154] ), .QN(n1633) );
  DFFRX1 \I_cache/cache_reg[2][154]  ( .D(n11589), .CK(clk), .RN(n5914), .Q(
        \I_cache/cache[2][154] ), .QN(n3299) );
  DFFRX1 \I_cache/cache_reg[3][154]  ( .D(n11588), .CK(clk), .RN(n5914), .Q(
        \I_cache/cache[3][154] ), .QN(n1634) );
  DFFRX1 \I_cache/cache_reg[6][154]  ( .D(n11585), .CK(clk), .RN(n5914), .Q(
        \I_cache/cache[6][154] ), .QN(n3300) );
  DFFRX1 \I_cache/cache_reg[7][154]  ( .D(n11584), .CK(clk), .RN(n5914), .Q(
        \I_cache/cache[7][154] ), .QN(n1635) );
  DFFRX1 \I_cache/cache_reg[4][151]  ( .D(n11611), .CK(clk), .RN(n5912), .Q(
        \I_cache/cache[4][151] ) );
  DFFRX1 \I_cache/cache_reg[5][154]  ( .D(n11586), .CK(clk), .RN(n5914), .Q(
        \I_cache/cache[5][154] ) );
  DFFRX1 \i_MIPS/ID_EX_reg[86]  ( .D(\i_MIPS/n499 ), .CK(clk), .RN(n5611), .Q(
        \i_MIPS/ID_EX[86] ), .QN(n4709) );
  DFFRX1 \I_cache/cache_reg[7][138]  ( .D(n11712), .CK(clk), .RN(n5903), .Q(
        \I_cache/cache[7][138] ), .QN(n366) );
  DFFRX1 \I_cache/cache_reg[1][129]  ( .D(n11790), .CK(clk), .RN(n5897), .Q(
        \I_cache/cache[1][129] ), .QN(n1586) );
  DFFRX1 \I_cache/cache_reg[4][129]  ( .D(n11787), .CK(clk), .RN(n5897), .Q(
        \I_cache/cache[4][129] ), .QN(n3220) );
  DFFRX1 \I_cache/cache_reg[6][129]  ( .D(n11785), .CK(clk), .RN(n5897), .Q(
        \I_cache/cache[6][129] ), .QN(n3221) );
  DFFRX1 \I_cache/cache_reg[1][136]  ( .D(n11734), .CK(clk), .RN(n5902), .Q(
        \I_cache/cache[1][136] ), .QN(n3219) );
  DFFRX1 \I_cache/cache_reg[1][142]  ( .D(n11686), .CK(clk), .RN(n5906), .Q(
        \I_cache/cache[1][142] ), .QN(n3240) );
  DFFRX1 \I_cache/cache_reg[3][142]  ( .D(n11684), .CK(clk), .RN(n5906), .Q(
        \I_cache/cache[3][142] ), .QN(n3243) );
  DFFRX4 \i_MIPS/ID_EX_reg[9]  ( .D(\i_MIPS/n562 ), .CK(clk), .RN(n5619), .Q(
        \i_MIPS/ALUin1[0] ), .QN(\i_MIPS/n371 ) );
  DFFRX4 \i_MIPS/PC/PC_o_reg[3]  ( .D(\i_MIPS/PC/n37 ), .CK(clk), .RN(n5620), 
        .Q(ICACHE_addr[1]), .QN(\i_MIPS/PC/n5 ) );
  DFFRX4 \i_MIPS/ID_EX_reg[107]  ( .D(\i_MIPS/n520 ), .CK(clk), .RN(n5615), 
        .Q(\i_MIPS/ID_EX[107] ), .QN(\i_MIPS/n327 ) );
  DFFRHQX8 \i_MIPS/ID_EX_reg[8]  ( .D(\i_MIPS/n470 ), .CK(clk), .RN(n5609), 
        .Q(n4428) );
  DFFRHQX8 \i_MIPS/PC/PC_o_reg[5]  ( .D(\i_MIPS/PC/n39 ), .CK(clk), .RN(n5620), 
        .Q(n4425) );
  DFFRHQX8 \i_MIPS/PC/PC_o_reg[6]  ( .D(\i_MIPS/PC/n40 ), .CK(clk), .RN(n5620), 
        .Q(n4423) );
  DFFRHQX8 \i_MIPS/ID_EX_reg[6]  ( .D(\i_MIPS/n472 ), .CK(clk), .RN(n5609), 
        .Q(n4413) );
  DFFRX4 \i_MIPS/ID_EX_reg[10]  ( .D(\i_MIPS/n561 ), .CK(clk), .RN(n5619), .Q(
        \i_MIPS/ALUin1[1] ), .QN(\i_MIPS/n370 ) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[16]  ( .D(\i_MIPS/PC/n50 ), .CK(clk), .RN(n5621), 
        .Q(ICACHE_addr[14]), .QN(\i_MIPS/PC/n18 ) );
  DFFRX4 \i_MIPS/ID_EX_reg[11]  ( .D(\i_MIPS/n560 ), .CK(clk), .RN(n5619), .Q(
        \i_MIPS/ALUin1[2] ), .QN(\i_MIPS/n369 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[58]  ( .D(\i_MIPS/n403 ), .CK(clk), .RN(n5603), .Q(
        n3489), .QN(\i_MIPS/n275 ) );
  DFFRX4 \i_MIPS/ID_EX_reg[87]  ( .D(\i_MIPS/n498 ), .CK(clk), .RN(n5611), .Q(
        \i_MIPS/ID_EX[87] ), .QN(n4713) );
  DFFRX4 \i_MIPS/IF_ID_reg[50]  ( .D(\i_MIPS/N73 ), .CK(clk), .RN(n5614), .Q(
        \i_MIPS/IR_ID[18] ), .QN(\i_MIPS/n316 ) );
  DFFRX4 \i_MIPS/ID_EX_reg[41]  ( .D(\i_MIPS/n437 ), .CK(clk), .RN(n5606), .Q(
        \i_MIPS/ID_EX[41] ), .QN(\i_MIPS/n309 ) );
  DFFRX4 \i_MIPS/PC/PC_o_reg[2]  ( .D(\i_MIPS/PC/n36 ), .CK(clk), .RN(n5620), 
        .Q(ICACHE_addr[0]), .QN(\i_MIPS/PC/n4 ) );
  DFFRX4 \i_MIPS/IF_ID_reg[49]  ( .D(\i_MIPS/N72 ), .CK(clk), .RN(n5614), .Q(
        \i_MIPS/IR_ID[17] ), .QN(\i_MIPS/n314 ) );
  DFFRX4 \i_MIPS/ID_EX_reg[45]  ( .D(\i_MIPS/n429 ), .CK(clk), .RN(n5606), .Q(
        n3487), .QN(\i_MIPS/n301 ) );
  DFFRX4 \i_MIPS/IF_ID_reg[56]  ( .D(\i_MIPS/N79 ), .CK(clk), .RN(n5615), .Q(
        \i_MIPS/IR_ID[24] ), .QN(\i_MIPS/n231 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[92]  ( .D(\i_MIPS/N115 ), .CK(clk), .RN(n5596), .Q(
        \i_MIPS/IF_ID[92] ), .QN(\i_MIPS/n174 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[112]  ( .D(\i_MIPS/n514 ), .CK(clk), .RN(n5614), 
        .Q(\i_MIPS/ID_EX[112] ), .QN(\i_MIPS/n315 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[83]  ( .D(\i_MIPS/N106 ), .CK(clk), .RN(n5597), .Q(
        \i_MIPS/IF_ID[83] ), .QN(\i_MIPS/n165 ) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[17]  ( .D(\i_MIPS/PC/n51 ), .CK(clk), .RN(n5621), 
        .Q(ICACHE_addr[15]), .QN(\i_MIPS/PC/n19 ) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[24]  ( .D(\i_MIPS/PC/n58 ), .CK(clk), .RN(n5622), 
        .Q(ICACHE_addr[22]), .QN(\i_MIPS/PC/n26 ) );
  DFFRX4 \i_MIPS/ID_EX_reg[108]  ( .D(\i_MIPS/n521 ), .CK(clk), .RN(n5616), 
        .Q(\i_MIPS/ID_EX[108] ), .QN(\i_MIPS/n329 ) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[29]  ( .D(n11543), .CK(clk), .RN(n5622), .Q(
        ICACHE_addr[27]), .QN(\i_MIPS/PC/n31 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[96]  ( .D(\i_MIPS/N119 ), .CK(clk), .RN(n5596), .Q(
        \i_MIPS/IF_ID[96] ), .QN(\i_MIPS/n178 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[102]  ( .D(\i_MIPS/n483 ), .CK(clk), .RN(n5610), 
        .Q(\i_MIPS/ID_EX[102] ) );
  DFFRX2 \i_MIPS/IF_ID_reg[94]  ( .D(\i_MIPS/N117 ), .CK(clk), .RN(n5596), .Q(
        \i_MIPS/IF_ID[94] ), .QN(\i_MIPS/n176 ) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[26]  ( .D(\i_MIPS/PC/n60 ), .CK(clk), .RN(n5622), 
        .Q(ICACHE_addr[24]), .QN(\i_MIPS/PC/n28 ) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[19]  ( .D(\i_MIPS/PC/n53 ), .CK(clk), .RN(n5621), 
        .Q(ICACHE_addr[17]), .QN(\i_MIPS/PC/n21 ) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[23]  ( .D(\i_MIPS/PC/n57 ), .CK(clk), .RN(n5622), 
        .Q(ICACHE_addr[21]), .QN(\i_MIPS/PC/n25 ) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[7]  ( .D(\i_MIPS/PC/n41 ), .CK(clk), .RN(n5620), 
        .Q(ICACHE_addr[5]), .QN(\i_MIPS/PC/n9 ) );
  DFFRX4 \i_MIPS/PC/PC_o_reg[0]  ( .D(\i_MIPS/PC/n34 ), .CK(clk), .RN(n5620), 
        .Q(\i_MIPS/BranchAddr[0] ), .QN(n3502) );
  DFFRX2 \i_MIPS/IF_ID_reg[89]  ( .D(\i_MIPS/N112 ), .CK(clk), .RN(n5596), .Q(
        \i_MIPS/IF_ID[89] ), .QN(\i_MIPS/n171 ) );
  DFFRX4 \i_MIPS/IF_ID_reg[52]  ( .D(\i_MIPS/N75 ), .CK(clk), .RN(n5615), .Q(
        \i_MIPS/IR_ID[20] ), .QN(\i_MIPS/n320 ) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[28]  ( .D(\i_MIPS/PC/n62 ), .CK(clk), .RN(n5622), 
        .Q(ICACHE_addr[26]), .QN(\i_MIPS/PC/n30 ) );
  DFFRHQX8 \i_MIPS/EX_MEM_reg[11]  ( .D(\i_MIPS/n463 ), .CK(clk), .RN(n5608), 
        .Q(n3839) );
  DFFRX2 \i_MIPS/ID_EX_reg[63]  ( .D(\i_MIPS/n393 ), .CK(clk), .RN(n5603), .Q(
        n4498), .QN(\i_MIPS/n265 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[50]  ( .D(\i_MIPS/n419 ), .CK(clk), .RN(n5605), .Q(
        \i_MIPS/ID_EX[50] ), .QN(\i_MIPS/n291 ) );
  DFFRX4 \i_MIPS/ID_EX_reg[42]  ( .D(\i_MIPS/n435 ), .CK(clk), .RN(n5606), 
        .QN(\i_MIPS/n307 ) );
  DFFRHQX8 \i_MIPS/EX_MEM_reg[9]  ( .D(\i_MIPS/n465 ), .CK(clk), .RN(n5609), 
        .Q(n3751) );
  DFFRX4 \i_MIPS/ID_EX_reg[37]  ( .D(\i_MIPS/n534 ), .CK(clk), .RN(n5617), .Q(
        \i_MIPS/ALUin1[28] ), .QN(\i_MIPS/n343 ) );
  DFFRX4 \i_MIPS/ID_EX_reg[109]  ( .D(\i_MIPS/n522 ), .CK(clk), .RN(n5616), 
        .QN(\i_MIPS/n331 ) );
  DFFRX4 \i_MIPS/ID_EX_reg[110]  ( .D(\i_MIPS/n523 ), .CK(clk), .RN(n5616), 
        .QN(\i_MIPS/n333 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[27]  ( .D(\i_MIPS/n447 ), .CK(clk), .RN(n5607), 
        .Q(n12948), .QN(n2315) );
  DFFRHQX4 \i_MIPS/PC/PC_o_reg[10]  ( .D(\i_MIPS/PC/n44 ), .CK(clk), .RN(n5620), .Q(n3649) );
  DFFRHQX4 \i_MIPS/PC/PC_o_reg[8]  ( .D(\i_MIPS/PC/n42 ), .CK(clk), .RN(n5620), 
        .Q(n3647) );
  DFFRHQX4 \i_MIPS/PC/PC_o_reg[9]  ( .D(\i_MIPS/PC/n43 ), .CK(clk), .RN(n5620), 
        .Q(n3645) );
  DFFRX4 \i_MIPS/ID_EX_reg[52]  ( .D(\i_MIPS/n415 ), .CK(clk), .RN(n5604), .Q(
        n3633), .QN(\i_MIPS/n287 ) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[31]  ( .D(n11544), .CK(clk), .RN(n5622), .Q(
        ICACHE_addr[29]), .QN(\i_MIPS/PC/n33 ) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[20]  ( .D(\i_MIPS/PC/n54 ), .CK(clk), .RN(n5621), 
        .Q(ICACHE_addr[18]), .QN(\i_MIPS/PC/n22 ) );
  DFFRHQX8 \i_MIPS/ID_EX_reg[79]  ( .D(\i_MIPS/n506 ), .CK(clk), .RN(n5612), 
        .Q(n3524) );
  DFFRX1 \i_MIPS/EX_MEM_reg[28]  ( .D(\i_MIPS/n446 ), .CK(clk), .RN(n5607), 
        .Q(n12947), .QN(n5) );
  DFFRX1 \i_MIPS/IF_ID_reg[62]  ( .D(\i_MIPS/N85 ), .CK(clk), .RN(n5616), .Q(
        \i_MIPS/IR_ID[30] ), .QN(\i_MIPS/n330 ) );
  DFFRHQX2 \i_MIPS/ID_EX_reg[47]  ( .D(\i_MIPS/n425 ), .CK(clk), .RN(n5605), 
        .Q(n3791) );
  DFFRX1 \i_MIPS/IF_ID_reg[61]  ( .D(\i_MIPS/N84 ), .CK(clk), .RN(n5616), .Q(
        \i_MIPS/IR_ID[29] ), .QN(\i_MIPS/n328 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[59]  ( .D(\i_MIPS/N82 ), .CK(clk), .RN(n5615), .Q(
        \i_MIPS/IR_ID[27] ), .QN(\i_MIPS/n324 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[11]  ( .D(\i_MIPS/N34 ), .CK(clk), .RN(n5600), .QN(
        \i_MIPS/n191 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[13]  ( .D(\i_MIPS/N36 ), .CK(clk), .RN(n5600), .QN(
        \i_MIPS/n193 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[25]  ( .D(\i_MIPS/N48 ), .CK(clk), .RN(n5599), .QN(
        \i_MIPS/n205 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[71]  ( .D(\i_MIPS/n377 ), .CK(clk), .RN(n5601), .Q(
        n3501), .QN(\i_MIPS/n249 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[65]  ( .D(\i_MIPS/n389 ), .CK(clk), .RN(n5602), .Q(
        n3499), .QN(\i_MIPS/n261 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[61]  ( .D(\i_MIPS/n397 ), .CK(clk), .RN(n5603), .Q(
        n3498), .QN(\i_MIPS/n269 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[57]  ( .D(\i_MIPS/n405 ), .CK(clk), .RN(n5604), .Q(
        n3497), .QN(\i_MIPS/n277 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[48]  ( .D(\i_MIPS/n423 ), .CK(clk), .RN(n5605), .Q(
        n3496), .QN(\i_MIPS/n295 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[64]  ( .D(\i_MIPS/n391 ), .CK(clk), .RN(n5602), .Q(
        n3495), .QN(\i_MIPS/n263 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[54]  ( .D(\i_MIPS/n411 ), .CK(clk), .RN(n5604), .Q(
        n3494), .QN(\i_MIPS/n283 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[62]  ( .D(\i_MIPS/n395 ), .CK(clk), .RN(n5603), .Q(
        n3492), .QN(\i_MIPS/n267 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[44]  ( .D(\i_MIPS/n431 ), .CK(clk), .RN(n5606), .Q(
        n3491), .QN(\i_MIPS/n303 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[60]  ( .D(\i_MIPS/n399 ), .CK(clk), .RN(n5603), .Q(
        n3490), .QN(\i_MIPS/n271 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[46]  ( .D(\i_MIPS/n427 ), .CK(clk), .RN(n5605), .Q(
        n3486), .QN(\i_MIPS/n299 ) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[11]  ( .D(\i_MIPS/PC/n45 ), .CK(clk), .RN(n5621), 
        .Q(ICACHE_addr[9]), .QN(\i_MIPS/PC/n13 ) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[13]  ( .D(\i_MIPS/PC/n47 ), .CK(clk), .RN(n5621), 
        .Q(ICACHE_addr[11]), .QN(\i_MIPS/PC/n15 ) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[14]  ( .D(\i_MIPS/PC/n48 ), .CK(clk), .RN(n5621), 
        .Q(ICACHE_addr[12]), .QN(\i_MIPS/PC/n16 ) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[15]  ( .D(\i_MIPS/PC/n49 ), .CK(clk), .RN(n5621), 
        .Q(ICACHE_addr[13]), .QN(\i_MIPS/PC/n17 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[24]  ( .D(\i_MIPS/n450 ), .CK(clk), .RN(n5607), 
        .Q(n12951), .QN(n4746) );
  DFFRX1 \i_MIPS/EX_MEM_reg[34]  ( .D(\i_MIPS/n440 ), .CK(clk), .RN(n5607), 
        .Q(n12941), .QN(n4492) );
  DFFRX1 \i_MIPS/ID_EX_reg[114]  ( .D(\i_MIPS/n516 ), .CK(clk), .RN(n5614), 
        .Q(\i_MIPS/ID_EX[114] ), .QN(\i_MIPS/n319 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[105]  ( .D(\i_MIPS/n518 ), .CK(clk), .RN(n5615), 
        .Q(\i_MIPS/ID_EX[105] ), .QN(\i_MIPS/n323 ) );
  DFFRX1 \I_cache/cache_reg[7][142]  ( .D(n11680), .CK(clk), .RN(n5906), .Q(
        \I_cache/cache[7][142] ), .QN(n3309) );
  DFFRX1 \I_cache/cache_reg[6][151]  ( .D(n11609), .CK(clk), .RN(n5912), .Q(
        \I_cache/cache[6][151] ), .QN(n3308) );
  DFFRX1 \I_cache/cache_reg[2][139]  ( .D(n11709), .CK(clk), .RN(n5904), .Q(
        \I_cache/cache[2][139] ), .QN(n3307) );
  DFFRX1 \I_cache/cache_reg[3][151]  ( .D(n11612), .CK(clk), .RN(n5912), .Q(
        \I_cache/cache[3][151] ), .QN(n3306) );
  DFFRX1 \I_cache/cache_reg[1][151]  ( .D(n11614), .CK(clk), .RN(n5912), .Q(
        \I_cache/cache[1][151] ), .QN(n3305) );
  DFFRX1 \i_MIPS/EX_MEM_reg[29]  ( .D(\i_MIPS/n445 ), .CK(clk), .RN(n5607), 
        .Q(n12946), .QN(n4385) );
  DFFRX1 \i_MIPS/EX_MEM_reg[26]  ( .D(\i_MIPS/n448 ), .CK(clk), .RN(n5607), 
        .Q(n12949), .QN(n4756) );
  DFFRX1 \i_MIPS/EX_MEM_reg[25]  ( .D(\i_MIPS/n449 ), .CK(clk), .RN(n5607), 
        .Q(n12950), .QN(n3256) );
  DFFRX1 \i_MIPS/EX_MEM_reg[12]  ( .D(\i_MIPS/n462 ), .CK(clk), .RN(n5608), 
        .Q(n12963), .QN(n3255) );
  DFFRX1 \i_MIPS/EX_MEM_reg[20]  ( .D(\i_MIPS/n454 ), .CK(clk), .RN(n5608), 
        .Q(n12955), .QN(n3254) );
  DFFRX1 \i_MIPS/EX_MEM_reg[16]  ( .D(\i_MIPS/n458 ), .CK(clk), .RN(n5608), 
        .Q(n12959), .QN(n3253) );
  DFFRX1 \i_MIPS/EX_MEM_reg[14]  ( .D(\i_MIPS/n460 ), .CK(clk), .RN(n5608), 
        .Q(n12961), .QN(n3252) );
  DFFRX1 \i_MIPS/EX_MEM_reg[32]  ( .D(\i_MIPS/n442 ), .CK(clk), .RN(n5607), 
        .Q(n12943), .QN(n3251) );
  DFFRX1 \i_MIPS/EX_MEM_reg[35]  ( .D(\i_MIPS/n439 ), .CK(clk), .RN(n5606), 
        .Q(n12940), .QN(n3246) );
  DFFRX1 \i_MIPS/EX_MEM_reg[15]  ( .D(\i_MIPS/n459 ), .CK(clk), .RN(n5608), 
        .Q(n12960), .QN(n3245) );
  DFFRX2 \i_MIPS/ID_EX_reg[36]  ( .D(\i_MIPS/n535 ), .CK(clk), .RN(n5617), .Q(
        \i_MIPS/ALUin1[27] ), .QN(\i_MIPS/n344 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[18]  ( .D(\i_MIPS/n456 ), .CK(clk), .RN(n5608), 
        .Q(n12957), .QN(n285) );
  DFFRX1 \i_MIPS/EX_MEM_reg[13]  ( .D(\i_MIPS/n461 ), .CK(clk), .RN(n5608), 
        .Q(n12962), .QN(n3244) );
  DFFRX1 \i_MIPS/EX_MEM_reg[19]  ( .D(\i_MIPS/n455 ), .CK(clk), .RN(n5608), 
        .Q(n12956), .QN(n283) );
  DFFRX2 \i_MIPS/ID_EX_reg[30]  ( .D(\i_MIPS/n541 ), .CK(clk), .RN(n5618), .Q(
        \i_MIPS/ALUin1[21] ), .QN(\i_MIPS/n350 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[8]  ( .D(\i_MIPS/n466 ), .CK(clk), .RN(n5609), .Q(
        n12964), .QN(n3238) );
  DFFRX1 \i_MIPS/ID_EX_reg[113]  ( .D(\i_MIPS/n515 ), .CK(clk), .RN(n5614), 
        .Q(\i_MIPS/ID_EX[113] ), .QN(\i_MIPS/n317 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[111]  ( .D(\i_MIPS/n513 ), .CK(clk), .RN(n5614), 
        .Q(\i_MIPS/ID_EX[111] ), .QN(\i_MIPS/n313 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[21]  ( .D(\i_MIPS/n453 ), .CK(clk), .RN(n5608), 
        .Q(n12954), .QN(n3199) );
  DFFRX2 \i_MIPS/ID_EX_reg[16]  ( .D(\i_MIPS/n555 ), .CK(clk), .RN(n5619), .Q(
        \i_MIPS/ALUin1[7] ), .QN(\i_MIPS/n364 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[20]  ( .D(\i_MIPS/n551 ), .CK(clk), .RN(n5618), .Q(
        \i_MIPS/ALUin1[11] ), .QN(\i_MIPS/n360 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[39]  ( .D(\i_MIPS/n532 ), .CK(clk), .RN(n5617), .Q(
        \i_MIPS/ALUin1[30] ), .QN(\i_MIPS/n341 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[22]  ( .D(\i_MIPS/n549 ), .CK(clk), .RN(n5618), .Q(
        \i_MIPS/ALUin1[13] ), .QN(\i_MIPS/n358 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[28]  ( .D(\i_MIPS/n543 ), .CK(clk), .RN(n5618), .Q(
        \i_MIPS/ALUin1[19] ), .QN(\i_MIPS/n352 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[34]  ( .D(\i_MIPS/n537 ), .CK(clk), .RN(n5617), .Q(
        \i_MIPS/ALUin1[25] ), .QN(\i_MIPS/n346 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[32]  ( .D(\i_MIPS/n539 ), .CK(clk), .RN(n5617), .Q(
        \i_MIPS/ALUin1[23] ), .QN(\i_MIPS/n348 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[55]  ( .D(\i_MIPS/n409 ), .CK(clk), .RN(n5604), .Q(
        \i_MIPS/ID_EX[55] ), .QN(\i_MIPS/n281 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[115]  ( .D(\i_MIPS/n517 ), .CK(clk), .RN(n5615), 
        .Q(\i_MIPS/ID_EX[115] ), .QN(\i_MIPS/n321 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[31]  ( .D(\i_MIPS/n540 ), .CK(clk), .RN(n5618), .Q(
        \i_MIPS/ALUin1[22] ), .QN(\i_MIPS/n349 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[26]  ( .D(\i_MIPS/n545 ), .CK(clk), .RN(n5618), .Q(
        \i_MIPS/ALUin1[17] ), .QN(\i_MIPS/n354 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[33]  ( .D(\i_MIPS/n538 ), .CK(clk), .RN(n5617), .Q(
        \i_MIPS/ALUin1[24] ), .QN(\i_MIPS/n347 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[21]  ( .D(\i_MIPS/n550 ), .CK(clk), .RN(n5618), .Q(
        \i_MIPS/ALUin1[12] ), .QN(\i_MIPS/n359 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[29]  ( .D(\i_MIPS/n542 ), .CK(clk), .RN(n5618), .Q(
        \i_MIPS/ALUin1[20] ), .QN(\i_MIPS/n351 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[40]  ( .D(\i_MIPS/n531 ), .CK(clk), .RN(n5617), .Q(
        \i_MIPS/ALU/N303 ), .QN(\i_MIPS/n340 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[38]  ( .D(\i_MIPS/n533 ), .CK(clk), .RN(n5617), .Q(
        \i_MIPS/ALUin1[29] ), .QN(\i_MIPS/n342 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[27]  ( .D(\i_MIPS/n544 ), .CK(clk), .RN(n5618), .Q(
        \i_MIPS/ALUin1[18] ), .QN(\i_MIPS/n353 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[4]  ( .D(\i_MIPS/n479 ), .CK(clk), .RN(n5610), 
        .QN(\i_MIPS/n310 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[60]  ( .D(\i_MIPS/N83 ), .CK(clk), .RN(n5616), .Q(
        \i_MIPS/IR_ID[28] ), .QN(\i_MIPS/n326 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[58]  ( .D(\i_MIPS/N81 ), .CK(clk), .RN(n5615), .Q(
        \i_MIPS/IR_ID[26] ), .QN(\i_MIPS/n322 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[63]  ( .D(\i_MIPS/N86 ), .CK(clk), .RN(n5616), .Q(
        \i_MIPS/IR_ID[31] ), .QN(\i_MIPS/n332 ) );
  DFFRX2 \i_MIPS/EX_MEM_reg[73]  ( .D(\i_MIPS/n473 ), .CK(clk), .RN(n5609), 
        .Q(\i_MIPS/Reg_W[4] ), .QN(n4715) );
  DFFRX2 \i_MIPS/ID_EX_reg[19]  ( .D(\i_MIPS/n552 ), .CK(clk), .RN(n5619), .Q(
        \i_MIPS/ALUin1[10] ), .QN(\i_MIPS/n361 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[17]  ( .D(\i_MIPS/n554 ), .CK(clk), .RN(n5619), .Q(
        \i_MIPS/ALUin1[8] ), .QN(\i_MIPS/n363 ) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[12]  ( .D(\i_MIPS/PC/n46 ), .CK(clk), .RN(n5621), 
        .Q(ICACHE_addr[10]), .QN(\i_MIPS/PC/n14 ) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[18]  ( .D(\i_MIPS/PC/n52 ), .CK(clk), .RN(n5621), 
        .Q(ICACHE_addr[16]), .QN(\i_MIPS/PC/n20 ) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[21]  ( .D(\i_MIPS/PC/n55 ), .CK(clk), .RN(n5621), 
        .Q(ICACHE_addr[19]), .QN(\i_MIPS/PC/n23 ) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[22]  ( .D(\i_MIPS/PC/n56 ), .CK(clk), .RN(n5621), 
        .Q(ICACHE_addr[20]), .QN(\i_MIPS/PC/n24 ) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[25]  ( .D(\i_MIPS/PC/n59 ), .CK(clk), .RN(n5622), 
        .Q(ICACHE_addr[23]), .QN(\i_MIPS/PC/n27 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[106]  ( .D(\i_MIPS/n519 ), .CK(clk), .RN(n5615), 
        .Q(\i_MIPS/ID_EX[106] ), .QN(\i_MIPS/n325 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[91]  ( .D(\i_MIPS/n494 ), .CK(clk), .RN(n5611), .Q(
        \i_MIPS/ID_EX[91] ), .QN(n4642) );
  DFFRX1 \i_MIPS/EX_MEM_reg[33]  ( .D(\i_MIPS/n441 ), .CK(clk), .RN(n5607), 
        .Q(n12942), .QN(n4395) );
  DFFRX1 \i_MIPS/EX_MEM_reg[31]  ( .D(\i_MIPS/n443 ), .CK(clk), .RN(n5607), 
        .Q(n12944), .QN(n4393) );
  DFFRX1 \i_MIPS/EX_MEM_reg[68]  ( .D(\i_MIPS/n374 ), .CK(clk), .RN(n5601), 
        .Q(n12966), .QN(\i_MIPS/n246 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[37]  ( .D(\i_MIPS/n436 ), .CK(clk), .RN(n5606), 
        .Q(n12997), .QN(\i_MIPS/n308 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[38]  ( .D(\i_MIPS/n434 ), .CK(clk), .RN(n5606), 
        .Q(n12996), .QN(\i_MIPS/n306 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[39]  ( .D(\i_MIPS/n432 ), .CK(clk), .RN(n5606), 
        .Q(n12995), .QN(\i_MIPS/n304 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[40]  ( .D(\i_MIPS/n430 ), .CK(clk), .RN(n5606), 
        .Q(n12994), .QN(\i_MIPS/n302 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[41]  ( .D(\i_MIPS/n428 ), .CK(clk), .RN(n5606), 
        .Q(n12993), .QN(\i_MIPS/n300 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[42]  ( .D(\i_MIPS/n426 ), .CK(clk), .RN(n5605), 
        .Q(n12992), .QN(\i_MIPS/n298 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[43]  ( .D(\i_MIPS/n424 ), .CK(clk), .RN(n5605), 
        .Q(n12991), .QN(\i_MIPS/n296 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[44]  ( .D(\i_MIPS/n422 ), .CK(clk), .RN(n5605), 
        .Q(n12990), .QN(\i_MIPS/n294 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[47]  ( .D(\i_MIPS/n416 ), .CK(clk), .RN(n5605), 
        .Q(n12987), .QN(\i_MIPS/n288 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[56]  ( .D(\i_MIPS/n398 ), .CK(clk), .RN(n5603), 
        .Q(n12978), .QN(\i_MIPS/n270 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[58]  ( .D(\i_MIPS/n394 ), .CK(clk), .RN(n5603), 
        .Q(n12976), .QN(\i_MIPS/n266 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[59]  ( .D(\i_MIPS/n392 ), .CK(clk), .RN(n5603), 
        .Q(n12975), .QN(\i_MIPS/n264 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[60]  ( .D(\i_MIPS/n390 ), .CK(clk), .RN(n5602), 
        .Q(n12974), .QN(\i_MIPS/n262 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[62]  ( .D(\i_MIPS/n386 ), .CK(clk), .RN(n5602), 
        .Q(n12972), .QN(\i_MIPS/n258 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[65]  ( .D(\i_MIPS/n380 ), .CK(clk), .RN(n5602), 
        .Q(n12969), .QN(\i_MIPS/n252 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[45]  ( .D(\i_MIPS/n420 ), .CK(clk), .RN(n5605), 
        .Q(n12989), .QN(\i_MIPS/n292 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[46]  ( .D(\i_MIPS/n418 ), .CK(clk), .RN(n5605), 
        .Q(n12988), .QN(\i_MIPS/n290 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[48]  ( .D(\i_MIPS/n414 ), .CK(clk), .RN(n5604), 
        .Q(n12986), .QN(\i_MIPS/n286 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[49]  ( .D(\i_MIPS/n412 ), .CK(clk), .RN(n5604), 
        .Q(n12985), .QN(\i_MIPS/n284 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[50]  ( .D(\i_MIPS/n410 ), .CK(clk), .RN(n5604), 
        .Q(n12984), .QN(\i_MIPS/n282 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[53]  ( .D(\i_MIPS/n404 ), .CK(clk), .RN(n5604), 
        .Q(n12981), .QN(\i_MIPS/n276 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[54]  ( .D(\i_MIPS/n402 ), .CK(clk), .RN(n5603), 
        .Q(n12980), .QN(\i_MIPS/n274 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[55]  ( .D(\i_MIPS/n400 ), .CK(clk), .RN(n5603), 
        .Q(n12979), .QN(\i_MIPS/n272 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[57]  ( .D(\i_MIPS/n396 ), .CK(clk), .RN(n5603), 
        .Q(n12977), .QN(\i_MIPS/n268 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[61]  ( .D(\i_MIPS/n388 ), .CK(clk), .RN(n5602), 
        .Q(n12973), .QN(\i_MIPS/n260 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[63]  ( .D(\i_MIPS/n384 ), .CK(clk), .RN(n5602), 
        .Q(n12971), .QN(\i_MIPS/n256 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[64]  ( .D(\i_MIPS/n382 ), .CK(clk), .RN(n5602), 
        .Q(n12970), .QN(\i_MIPS/n254 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[66]  ( .D(\i_MIPS/n378 ), .CK(clk), .RN(n5601), 
        .Q(n12968), .QN(\i_MIPS/n250 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[51]  ( .D(\i_MIPS/n408 ), .CK(clk), .RN(n5604), 
        .Q(n12983), .QN(\i_MIPS/n280 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[52]  ( .D(\i_MIPS/n406 ), .CK(clk), .RN(n5604), 
        .Q(n12982), .QN(\i_MIPS/n278 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[67]  ( .D(\i_MIPS/n376 ), .CK(clk), .RN(n5601), 
        .Q(n12967), .QN(\i_MIPS/n248 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[89]  ( .D(\i_MIPS/n496 ), .CK(clk), .RN(n5611), .Q(
        \i_MIPS/ID_EX[89] ), .QN(n4643) );
  DFFRX1 \i_MIPS/ID_EX_reg[90]  ( .D(\i_MIPS/n495 ), .CK(clk), .RN(n5611), .Q(
        \i_MIPS/ID_EX[90] ), .QN(n4644) );
  DFFRX1 \i_MIPS/ID_EX_reg[93]  ( .D(\i_MIPS/n492 ), .CK(clk), .RN(n5611), .Q(
        \i_MIPS/ID_EX[93] ), .QN(n4646) );
  DFFRX1 \i_MIPS/ID_EX_reg[97]  ( .D(\i_MIPS/n488 ), .CK(clk), .RN(n5611), .Q(
        \i_MIPS/ID_EX[97] ), .QN(n4648) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[1]  ( .D(\i_MIPS/PC/n35 ), .CK(clk), .RN(n5620), 
        .Q(\i_MIPS/PC_o[1] ), .QN(\i_MIPS/PC/n3 ) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[30]  ( .D(n11542), .CK(clk), .RN(n5622), .Q(
        ICACHE_addr[28]), .QN(\i_MIPS/PC/n32 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[87]  ( .D(\i_MIPS/N110 ), .CK(clk), .RN(n5596), .Q(
        \i_MIPS/IF_ID[87] ), .QN(\i_MIPS/n169 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[75]  ( .D(\i_MIPS/N98 ), .CK(clk), .RN(n5597), .Q(
        \i_MIPS/IF_ID[75] ), .QN(\i_MIPS/n244 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[95]  ( .D(\i_MIPS/N118 ), .CK(clk), .RN(n5596), .Q(
        \i_MIPS/IF_ID[95] ), .QN(\i_MIPS/n177 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[101]  ( .D(\i_MIPS/n484 ), .CK(clk), .RN(n5610), 
        .Q(\i_MIPS/ID_EX[101] ) );
  DFFRX1 \i_MIPS/ID_EX_reg[104]  ( .D(\i_MIPS/n481 ), .CK(clk), .RN(n5610), 
        .Q(\i_MIPS/ID_EX[104] ) );
  DFFRX2 \i_MIPS/ID_EX_reg[95]  ( .D(\i_MIPS/n490 ), .CK(clk), .RN(n5611), .Q(
        \i_MIPS/ID_EX[95] ) );
  DFFRX1 \D_cache/cache_reg[7][18]  ( .D(\D_cache/n1645 ), .CK(clk), .RN(n5720), .Q(\D_cache/cache[7][18] ) );
  DFFRX1 \D_cache/cache_reg[5][128]  ( .D(\D_cache/n767 ), .CK(clk), .RN(n5793), .Q(\D_cache/cache[5][128] ) );
  DFFRX1 \D_cache/cache_reg[4][128]  ( .D(\D_cache/n768 ), .CK(clk), .RN(n5793), .Q(\D_cache/cache[4][128] ) );
  DFFRX1 \D_cache/cache_reg[7][131]  ( .D(\D_cache/n741 ), .CK(clk), .RN(n5795), .Q(\D_cache/cache[7][131] ) );
  DFFRX1 \D_cache/cache_reg[3][136]  ( .D(\D_cache/n705 ), .CK(clk), .RN(n5798), .Q(\D_cache/cache[3][136] ) );
  DFFRX1 \D_cache/cache_reg[2][136]  ( .D(\D_cache/n706 ), .CK(clk), .RN(n5798), .Q(\D_cache/cache[2][136] ) );
  DFFRHQX4 \i_MIPS/ID_EX_reg[74]  ( .D(\i_MIPS/n511 ), .CK(clk), .RN(n5612), 
        .Q(n3768) );
  DFFRX2 \i_MIPS/ID_EX_reg[51]  ( .D(\i_MIPS/n417 ), .CK(clk), .RN(n5605), .Q(
        n3743), .QN(\i_MIPS/n289 ) );
  DFFRX1 \D_cache/cache_reg[7][144]  ( .D(\D_cache/n637 ), .CK(clk), .RN(n5804), .Q(\D_cache/cache[7][144] ) );
  DFFRX1 \D_cache/cache_reg[7][128]  ( .D(\D_cache/n765 ), .CK(clk), .RN(n5810), .Q(\D_cache/cache[7][128] ) );
  DFFRHQX2 \i_MIPS/ID_EX_reg[76]  ( .D(\i_MIPS/n509 ), .CK(clk), .RN(n5612), 
        .Q(n3708) );
  DFFRHQX2 \i_MIPS/ID_EX_reg[77]  ( .D(\i_MIPS/n508 ), .CK(clk), .RN(n5612), 
        .Q(n3700) );
  DFFRX1 \D_cache/cache_reg[5][148]  ( .D(\D_cache/n607 ), .CK(clk), .RN(n5807), .Q(\D_cache/cache[5][148] ) );
  DFFRX2 \i_MIPS/ID_EX_reg[84]  ( .D(\i_MIPS/n501 ), .CK(clk), .RN(n5612), .Q(
        \i_MIPS/ID_EX[84] ), .QN(n4712) );
  DFFRX1 \I_cache/cache_reg[7][139]  ( .D(n11704), .CK(clk), .RN(n5904), .Q(
        \I_cache/cache[7][139] ) );
  DFFRX1 \i_MIPS/ID_EX_reg[53]  ( .D(\i_MIPS/n413 ), .CK(clk), .RN(n5604), .Q(
        n3493), .QN(\i_MIPS/n285 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[59]  ( .D(\i_MIPS/n401 ), .CK(clk), .RN(n5603), .Q(
        n3500), .QN(\i_MIPS/n273 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[49]  ( .D(\i_MIPS/n421 ), .CK(clk), .RN(n5605), .Q(
        \i_MIPS/ID_EX[49] ), .QN(\i_MIPS/n293 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[43]  ( .D(\i_MIPS/n433 ), .CK(clk), .RN(n5606), .Q(
        n3506), .QN(\i_MIPS/n305 ) );
  DFFRX4 \i_MIPS/ID_EX_reg[85]  ( .D(\i_MIPS/n500 ), .CK(clk), .RN(n5612), .Q(
        \i_MIPS/ID_EX[85] ), .QN(n4708) );
  DFFRX4 \i_MIPS/ID_EX_reg[88]  ( .D(\i_MIPS/n497 ), .CK(clk), .RN(n5611), .Q(
        \i_MIPS/ID_EX[88] ), .QN(n3310) );
  DFFRX4 \i_MIPS/ID_EX_reg[100]  ( .D(\i_MIPS/n485 ), .CK(clk), .RN(n5610), 
        .Q(\i_MIPS/ID_EX[100] ) );
  DFFRX2 \i_MIPS/IF_ID_reg[64]  ( .D(\i_MIPS/N87 ), .CK(clk), .RN(n5601), .Q(
        \i_MIPS/IF_ID[64] ), .QN(\i_MIPS/n233 ) );
  DFFRHQX8 \i_MIPS/ID_EX_reg[23]  ( .D(\i_MIPS/n548 ), .CK(clk), .RN(n5618), 
        .Q(n3827) );
  DFFRX4 \i_MIPS/ID_EX_reg[25]  ( .D(\i_MIPS/n546 ), .CK(clk), .RN(n5618), .Q(
        \i_MIPS/ALUin1[16] ), .QN(\i_MIPS/n355 ) );
  DFFRX4 \i_MIPS/ID_EX_reg[12]  ( .D(\i_MIPS/n559 ), .CK(clk), .RN(n5619), .Q(
        \i_MIPS/ALUin1[3] ), .QN(\i_MIPS/n368 ) );
  DFFRX4 \i_MIPS/EX_MEM_reg[7]  ( .D(\i_MIPS/n467 ), .CK(clk), .RN(n5609), .Q(
        n12965), .QN(n4047) );
  DFFRX4 \i_MIPS/ID_EX_reg[56]  ( .D(\i_MIPS/n407 ), .CK(clk), .RN(n5604), .Q(
        \i_MIPS/ID_EX[56] ), .QN(\i_MIPS/n279 ) );
  DFFRX4 \i_MIPS/IF_ID_reg[53]  ( .D(\i_MIPS/N76 ), .CK(clk), .RN(n5615), .Q(
        \i_MIPS/IR_ID[21] ), .QN(\i_MIPS/n228 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[66]  ( .D(\i_MIPS/n387 ), .CK(clk), .RN(n5602), .Q(
        n3488), .QN(\i_MIPS/n259 ) );
  DFFRX2 \D_cache/cache_reg[0][5]  ( .D(\D_cache/n1756 ), .CK(clk), .RN(n5711), 
        .Q(\D_cache/cache[0][5] ), .QN(n1365) );
  DFFRX2 \i_MIPS/IF_ID_reg[41]  ( .D(\i_MIPS/N64 ), .CK(clk), .RN(n5613), .QN(
        \i_MIPS/n221 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[27]  ( .D(\i_MIPS/N50 ), .CK(clk), .RN(n5599), .QN(
        \i_MIPS/n207 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[97]  ( .D(\i_MIPS/N120 ), .CK(clk), .RN(n5601), .Q(
        \i_MIPS/IF_ID[97] ), .QN(\i_MIPS/n179 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[21]  ( .D(\i_MIPS/N44 ), .CK(clk), .RN(n5599), .QN(
        \i_MIPS/n201 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[7]  ( .D(\i_MIPS/N30 ), .CK(clk), .RN(n5600), .QN(
        \i_MIPS/n187 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[42]  ( .D(\i_MIPS/N65 ), .CK(clk), .RN(n5613), .QN(
        \i_MIPS/n222 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[35]  ( .D(\i_MIPS/N58 ), .CK(clk), .RN(n5613), .Q(
        \i_MIPS/Sign_Extend_ID[3] ), .QN(\i_MIPS/n215 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[33]  ( .D(\i_MIPS/N56 ), .CK(clk), .RN(n5613), .Q(
        \i_MIPS/Sign_Extend_ID[1] ), .QN(\i_MIPS/n213 ) );
  DFFRX4 \i_MIPS/PC/PC_o_reg[27]  ( .D(\i_MIPS/PC/n61 ), .CK(clk), .RN(n5622), 
        .Q(ICACHE_addr[25]), .QN(\i_MIPS/PC/n29 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[1]  ( .D(\i_MIPS/N24 ), .CK(clk), .RN(n5601), .Q(
        \i_MIPS/IF_ID_1 ), .QN(\i_MIPS/n181 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[81]  ( .D(\i_MIPS/N104 ), .CK(clk), .RN(n5597), .Q(
        \i_MIPS/IF_ID[81] ), .QN(\i_MIPS/n163 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[16]  ( .D(\i_MIPS/N39 ), .CK(clk), .RN(n5599), .QN(
        \i_MIPS/n196 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[68]  ( .D(\i_MIPS/N91 ), .CK(clk), .RN(n5598), .Q(
        \i_MIPS/IF_ID[68] ), .QN(\i_MIPS/n237 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[71]  ( .D(\i_MIPS/N94 ), .CK(clk), .RN(n5598), .Q(
        \i_MIPS/IF_ID[71] ), .QN(\i_MIPS/n240 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[72]  ( .D(\i_MIPS/N95 ), .CK(clk), .RN(n5598), .Q(
        \i_MIPS/IF_ID[72] ), .QN(\i_MIPS/n241 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[6]  ( .D(\i_MIPS/N29 ), .CK(clk), .RN(n5600), .QN(
        \i_MIPS/n186 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[76]  ( .D(\i_MIPS/N99 ), .CK(clk), .RN(n5597), .Q(
        \i_MIPS/IF_ID[76] ), .QN(\i_MIPS/n245 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[91]  ( .D(\i_MIPS/N114 ), .CK(clk), .RN(n5596), .Q(
        \i_MIPS/IF_ID[91] ), .QN(\i_MIPS/n173 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[2]  ( .D(\i_MIPS/N25 ), .CK(clk), .RN(n5601), .Q(
        \i_MIPS/IF_ID_2 ), .QN(\i_MIPS/n182 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[67]  ( .D(\i_MIPS/N90 ), .CK(clk), .RN(n5598), .Q(
        \i_MIPS/IF_ID[67] ), .QN(\i_MIPS/n236 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[44]  ( .D(\i_MIPS/N67 ), .CK(clk), .RN(n5614), .QN(
        \i_MIPS/n224 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[79]  ( .D(\i_MIPS/N102 ), .CK(clk), .RN(n5597), .Q(
        \i_MIPS/IF_ID[79] ), .QN(\i_MIPS/n161 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[77]  ( .D(\i_MIPS/N100 ), .CK(clk), .RN(n5597), .Q(
        \i_MIPS/IF_ID[77] ), .QN(\i_MIPS/n159 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[22]  ( .D(\i_MIPS/N45 ), .CK(clk), .RN(n5599), .QN(
        \i_MIPS/n202 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[19]  ( .D(\i_MIPS/N42 ), .CK(clk), .RN(n5599), .QN(
        \i_MIPS/n199 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[24]  ( .D(\i_MIPS/N47 ), .CK(clk), .RN(n5599), .QN(
        \i_MIPS/n204 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[46]  ( .D(\i_MIPS/N69 ), .CK(clk), .RN(n5614), .QN(
        \i_MIPS/n226 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[36]  ( .D(\i_MIPS/N59 ), .CK(clk), .RN(n5613), .Q(
        \i_MIPS/Sign_Extend_ID[4] ), .QN(\i_MIPS/n216 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[90]  ( .D(\i_MIPS/N113 ), .CK(clk), .RN(n5596), .Q(
        \i_MIPS/IF_ID[90] ), .QN(\i_MIPS/n172 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[45]  ( .D(\i_MIPS/N68 ), .CK(clk), .RN(n5614), .QN(
        \i_MIPS/n225 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[37]  ( .D(\i_MIPS/N60 ), .CK(clk), .RN(n5613), .Q(
        \i_MIPS/Sign_Extend_ID[5] ), .QN(\i_MIPS/n217 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[39]  ( .D(\i_MIPS/N62 ), .CK(clk), .RN(n5613), .QN(
        \i_MIPS/n219 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[34]  ( .D(\i_MIPS/N57 ), .CK(clk), .RN(n5613), .Q(
        \i_MIPS/Sign_Extend_ID[2] ), .QN(\i_MIPS/n214 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[31]  ( .D(\i_MIPS/N54 ), .CK(clk), .RN(n5596), .QN(
        \i_MIPS/n211 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[17]  ( .D(\i_MIPS/N40 ), .CK(clk), .RN(n5599), .QN(
        \i_MIPS/n197 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[15]  ( .D(\i_MIPS/N38 ), .CK(clk), .RN(n5600), .QN(
        \i_MIPS/n195 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[88]  ( .D(\i_MIPS/N111 ), .CK(clk), .RN(n5596), .Q(
        \i_MIPS/IF_ID[88] ), .QN(\i_MIPS/n170 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[70]  ( .D(\i_MIPS/N93 ), .CK(clk), .RN(n5598), .Q(
        \i_MIPS/IF_ID[70] ), .QN(\i_MIPS/n239 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[0]  ( .D(\i_MIPS/N23 ), .CK(clk), .RN(n5601), .QN(
        \i_MIPS/n180 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[74]  ( .D(\i_MIPS/N97 ), .CK(clk), .RN(n5597), .Q(
        \i_MIPS/IF_ID[74] ), .QN(\i_MIPS/n243 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[73]  ( .D(\i_MIPS/N96 ), .CK(clk), .RN(n5598), .Q(
        \i_MIPS/IF_ID[73] ), .QN(\i_MIPS/n242 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[32]  ( .D(\i_MIPS/N55 ), .CK(clk), .RN(n5617), .Q(
        \i_MIPS/Sign_Extend_ID[0] ), .QN(\i_MIPS/n212 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[18]  ( .D(\i_MIPS/N41 ), .CK(clk), .RN(n5599), .QN(
        \i_MIPS/n198 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[23]  ( .D(\i_MIPS/N46 ), .CK(clk), .RN(n5599), .QN(
        \i_MIPS/n203 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[66]  ( .D(\i_MIPS/N89 ), .CK(clk), .RN(n5598), .Q(
        \i_MIPS/IF_ID[66] ), .QN(\i_MIPS/n235 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[10]  ( .D(\i_MIPS/N33 ), .CK(clk), .RN(n5600), .QN(
        \i_MIPS/n190 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[9]  ( .D(\i_MIPS/N32 ), .CK(clk), .RN(n5600), .QN(
        \i_MIPS/n189 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[8]  ( .D(\i_MIPS/N31 ), .CK(clk), .RN(n5600), .Q(
        n171), .QN(\i_MIPS/n188 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[69]  ( .D(\i_MIPS/N92 ), .CK(clk), .RN(n5598), .Q(
        \i_MIPS/IF_ID[69] ), .QN(\i_MIPS/n238 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[3]  ( .D(\i_MIPS/N26 ), .CK(clk), .RN(n5601), .QN(
        \i_MIPS/n183 ) );
  DFFRX2 \I_cache/cache_reg[7][97]  ( .D(n12040), .CK(clk), .RN(n5876), .Q(
        \I_cache/cache[7][97] ), .QN(n2712) );
  DFFRX2 \i_MIPS/IF_ID_reg[43]  ( .D(\i_MIPS/N66 ), .CK(clk), .RN(n5613), .QN(
        \i_MIPS/n223 ) );
  DFFRX2 \I_cache/cache_reg[7][31]  ( .D(n12568), .CK(clk), .RN(n5832), .Q(
        \I_cache/cache[7][31] ), .QN(n2583) );
  DFFRX2 \I_cache/cache_reg[5][25]  ( .D(n12618), .CK(clk), .RN(n5828), .Q(
        \I_cache/cache[5][25] ), .QN(n3469) );
  DFFRX2 \I_cache/cache_reg[5][108]  ( .D(n11954), .CK(clk), .RN(n5883), .Q(
        \I_cache/cache[5][108] ), .QN(n2622) );
  DFFRX2 \i_MIPS/IF_ID_reg[14]  ( .D(\i_MIPS/N37 ), .CK(clk), .RN(n5600), .QN(
        \i_MIPS/n194 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[12]  ( .D(\i_MIPS/N35 ), .CK(clk), .RN(n5600), .QN(
        \i_MIPS/n192 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[26]  ( .D(\i_MIPS/N49 ), .CK(clk), .RN(n5599), .QN(
        \i_MIPS/n206 ) );
  DFFRX2 \I_cache/cache_reg[3][80]  ( .D(n12180), .CK(clk), .RN(n5865), .Q(
        \I_cache/cache[3][80] ), .QN(n3443) );
  DFFRX2 \I_cache/cache_reg[7][5]  ( .D(n12776), .CK(clk), .RN(n5815), .Q(
        \I_cache/cache[7][5] ), .QN(n443) );
  DFFRX2 \I_cache/cache_reg[7][82]  ( .D(n12160), .CK(clk), .RN(n5866), .Q(
        \I_cache/cache[7][82] ), .QN(n3381) );
  DFFRX2 \I_cache/cache_reg[5][44]  ( .D(n12466), .CK(clk), .RN(n5841), .Q(
        \I_cache/cache[5][44] ), .QN(n2776) );
  DFFRX2 \I_cache/cache_reg[5][105]  ( .D(n11978), .CK(clk), .RN(n5881), .Q(
        \I_cache/cache[5][105] ), .QN(n745) );
  DFFRX2 \I_cache/cache_reg[5][12]  ( .D(n12722), .CK(clk), .RN(n5819), .Q(
        \I_cache/cache[5][12] ), .QN(n2623) );
  DFFRX2 \I_cache/cache_reg[3][16]  ( .D(n12692), .CK(clk), .RN(n5822), .Q(
        \I_cache/cache[3][16] ), .QN(n3386) );
  DFFRX2 \I_cache/cache_reg[5][73]  ( .D(n12234), .CK(clk), .RN(n5860), .Q(
        \I_cache/cache[5][73] ), .QN(n2327) );
  DFFRX2 \i_MIPS/IF_ID_reg[38]  ( .D(\i_MIPS/N61 ), .CK(clk), .RN(n5613), .Q(
        \i_MIPS/Sign_Extend_ID[6] ), .QN(\i_MIPS/n218 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[84]  ( .D(\i_MIPS/N107 ), .CK(clk), .RN(n5597), .Q(
        \i_MIPS/IF_ID[84] ), .QN(\i_MIPS/n166 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[80]  ( .D(\i_MIPS/N103 ), .CK(clk), .RN(n5597), .Q(
        \i_MIPS/IF_ID[80] ), .QN(\i_MIPS/n162 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[47]  ( .D(\i_MIPS/N70 ), .CK(clk), .RN(n5614), .Q(
        \i_MIPS/Sign_Extend_ID[31] ), .QN(\i_MIPS/n227 ) );
  DFFRX2 \I_cache/cache_reg[5][121]  ( .D(n11850), .CK(clk), .RN(n5892), .Q(
        \I_cache/cache[5][121] ), .QN(n3470) );
  DFFRX2 \I_cache/cache_reg[5][10]  ( .D(n12738), .CK(clk), .RN(n5818), .Q(
        \I_cache/cache[5][10] ), .QN(n2768) );
  DFFRX2 \I_cache/cache_reg[7][48]  ( .D(n12432), .CK(clk), .RN(n5844), .Q(
        \I_cache/cache[7][48] ), .QN(n3393) );
  DFFRX2 \I_cache/cache_reg[3][50]  ( .D(n12420), .CK(clk), .RN(n5845), .Q(
        \I_cache/cache[3][50] ), .QN(n3383) );
  DFFRX2 \I_cache/cache_reg[7][112]  ( .D(n11920), .CK(clk), .RN(n5886), .Q(
        \I_cache/cache[7][112] ), .QN(n3390) );
  DFFRX2 \I_cache/cache_reg[3][114]  ( .D(n11908), .CK(clk), .RN(n5887), .Q(
        \I_cache/cache[3][114] ), .QN(n3377) );
  DFFRX2 \I_cache/cache_reg[5][76]  ( .D(n12210), .CK(clk), .RN(n5862), .Q(
        \I_cache/cache[5][76] ), .QN(n2775) );
  DFFRX2 \I_cache/cache_reg[5][90]  ( .D(n12098), .CK(clk), .RN(n5871), .Q(
        \I_cache/cache[5][90] ), .QN(n2620) );
  DFFRX2 \I_cache/cache_reg[4][64]  ( .D(n12307), .CK(clk), .RN(n5854), .Q(
        \I_cache/cache[4][64] ), .QN(n1795) );
  DFFRX2 \I_cache/cache_reg[5][9]  ( .D(n12746), .CK(clk), .RN(n5817), .Q(
        \I_cache/cache[5][9] ), .QN(n2326) );
  DFFRX2 \I_cache/cache_reg[5][74]  ( .D(n12226), .CK(clk), .RN(n5861), .Q(
        \I_cache/cache[5][74] ), .QN(n744) );
  DFFRX2 \i_MIPS/IF_ID_reg[28]  ( .D(\i_MIPS/N51 ), .CK(clk), .RN(n5598), .Q(
        \i_MIPS/IF_ID_28 ), .QN(\i_MIPS/n208 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[30]  ( .D(\i_MIPS/N53 ), .CK(clk), .RN(n5598), .QN(
        \i_MIPS/n210 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[65]  ( .D(\i_MIPS/N88 ), .CK(clk), .RN(n5598), .Q(
        \i_MIPS/IF_ID[65] ), .QN(\i_MIPS/n234 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[29]  ( .D(\i_MIPS/N52 ), .CK(clk), .RN(n5598), .QN(
        \i_MIPS/n209 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[20]  ( .D(\i_MIPS/N43 ), .CK(clk), .RN(n5599), .QN(
        \i_MIPS/n200 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[4]  ( .D(\i_MIPS/N27 ), .CK(clk), .RN(n5600), .QN(
        \i_MIPS/n184 ) );
  DFFRX2 \I_cache/cache_reg[5][97]  ( .D(n12042), .CK(clk), .RN(n5876), .Q(
        \I_cache/cache[5][97] ), .QN(n2794) );
  DFFRX2 \I_cache/cache_reg[5][31]  ( .D(n12570), .CK(clk), .RN(n5832), .Q(
        \I_cache/cache[5][31] ), .QN(n2619) );
  DFFRX2 \I_cache/cache_reg[7][80]  ( .D(n12176), .CK(clk), .RN(n5865), .Q(
        \I_cache/cache[7][80] ), .QN(n3444) );
  DFFRX2 \I_cache/cache_reg[1][82]  ( .D(n12166), .CK(clk), .RN(n5866), .Q(
        \I_cache/cache[1][82] ), .QN(n3379) );
  DFFRX2 \I_cache/cache_reg[5][5]  ( .D(n12778), .CK(clk), .RN(n5815), .Q(
        \I_cache/cache[5][5] ), .QN(n774) );
  DFFRX2 \I_cache/cache_reg[4][10]  ( .D(n12739), .CK(clk), .RN(n5818), .Q(
        \I_cache/cache[4][10] ), .QN(n1196) );
  DFFRX2 \I_cache/cache_reg[4][16]  ( .D(n12691), .CK(clk), .RN(n5822), .Q(
        \I_cache/cache[4][16] ), .QN(n1731) );
  DFFRX2 \I_cache/cache_reg[7][25]  ( .D(n12616), .CK(clk), .RN(n5828), .Q(
        \I_cache/cache[7][25] ), .QN(n3450) );
  DFFRX2 \I_cache/cache_reg[7][108]  ( .D(n11952), .CK(clk), .RN(n5884), .Q(
        \I_cache/cache[7][108] ), .QN(n2427) );
  DFFRX2 \I_cache/cache_reg[3][48]  ( .D(n12436), .CK(clk), .RN(n5843), .Q(
        \I_cache/cache[3][48] ), .QN(n3392) );
  DFFRX2 \I_cache/cache_reg[2][12]  ( .D(n12725), .CK(clk), .RN(n5819), .Q(
        \I_cache/cache[2][12] ), .QN(n1035) );
  DFFRX2 \I_cache/cache_reg[7][50]  ( .D(n12416), .CK(clk), .RN(n5845), .Q(
        \I_cache/cache[7][50] ), .QN(n3384) );
  DFFRX2 \I_cache/cache_reg[5][64]  ( .D(n12306), .CK(clk), .RN(n5854), .Q(
        \I_cache/cache[5][64] ), .QN(n3479) );
  DFFRX2 \I_cache/cache_reg[1][112]  ( .D(n11926), .CK(clk), .RN(n5886), .Q(
        \I_cache/cache[1][112] ), .QN(n3388) );
  DFFRX2 \I_cache/cache_reg[4][114]  ( .D(n11907), .CK(clk), .RN(n5887), .Q(
        \I_cache/cache[4][114] ), .QN(n1728) );
  DFFRX2 \I_cache/cache_reg[7][44]  ( .D(n12464), .CK(clk), .RN(n5841), .Q(
        \I_cache/cache[7][44] ), .QN(n2613) );
  DFFRX2 \I_cache/cache_reg[7][121]  ( .D(n11848), .CK(clk), .RN(n5892), .Q(
        \I_cache/cache[7][121] ), .QN(n3453) );
  DFFRX2 \I_cache/cache_reg[4][90]  ( .D(n12099), .CK(clk), .RN(n5871), .Q(
        \I_cache/cache[4][90] ), .QN(n1048) );
  DFFRX2 \I_cache/cache_reg[7][76]  ( .D(n12208), .CK(clk), .RN(n5862), .Q(
        \I_cache/cache[7][76] ), .QN(n2625) );
  DFFRX2 \I_cache/cache_reg[4][9]  ( .D(n12747), .CK(clk), .RN(n5817), .Q(
        \I_cache/cache[4][9] ), .QN(n747) );
  DFFRX2 \I_cache/cache_reg[0][105]  ( .D(n11983), .CK(clk), .RN(n5881), .Q(
        \I_cache/cache[0][105] ), .QN(n1076) );
  DFFRX2 \I_cache/cache_reg[0][73]  ( .D(n12239), .CK(clk), .RN(n5860), .Q(
        \I_cache/cache[0][73] ), .QN(n1088) );
  DFFRX2 \I_cache/cache_reg[0][74]  ( .D(n12231), .CK(clk), .RN(n5860), .Q(
        \I_cache/cache[0][74] ), .QN(n907) );
  MX2X1 U2 ( .A(\I_cache/cache[4][9] ), .B(n9645), .S0(n5327), .Y(n12747) );
  MX2X1 U3 ( .A(\I_cache/cache[4][90] ), .B(n9711), .S0(n5327), .Y(n12099) );
  MX2X1 U4 ( .A(\I_cache/cache[7][121] ), .B(n10119), .S0(n5366), .Y(n11848)
         );
  MX2X1 U5 ( .A(\I_cache/cache[4][114] ), .B(n10041), .S0(n5324), .Y(n11907)
         );
  MX2X1 U6 ( .A(\I_cache/cache[1][112] ), .B(n10070), .S0(n5108), .Y(n11926)
         );
  MX2X1 U7 ( .A(\I_cache/cache[5][64] ), .B(n9683), .S0(n5279), .Y(n12306) );
  MX2X1 U8 ( .A(\I_cache/cache[7][50] ), .B(n10036), .S0(n5371), .Y(n12416) );
  MX2X1 U9 ( .A(\I_cache/cache[2][12] ), .B(n10085), .S0(n5240), .Y(n12725) );
  MX2X1 U10 ( .A(\I_cache/cache[3][48] ), .B(n10065), .S0(n5195), .Y(n12436)
         );
  MX2X1 U11 ( .A(\I_cache/cache[7][108] ), .B(n10095), .S0(n5366), .Y(n11952)
         );
  MX2X1 U12 ( .A(\I_cache/cache[4][16] ), .B(n10060), .S0(n5324), .Y(n12691)
         );
  MX2X1 U13 ( .A(\I_cache/cache[4][10] ), .B(n9659), .S0(n5327), .Y(n12739) );
  MX2X1 U14 ( .A(\I_cache/cache[5][5] ), .B(n9541), .S0(n5285), .Y(n12778) );
  MX2X1 U15 ( .A(\I_cache/cache[1][82] ), .B(n10046), .S0(n5108), .Y(n12166)
         );
  MX2X1 U16 ( .A(\I_cache/cache[7][80] ), .B(n10075), .S0(n5371), .Y(n12176)
         );
  MX2X1 U17 ( .A(\I_cache/cache[5][31] ), .B(n11035), .S0(n5278), .Y(n12570)
         );
  MX2X1 U18 ( .A(\I_cache/cache[5][97] ), .B(n9361), .S0(n5284), .Y(n12042) );
  OR2X2 U19 ( .A(n4558), .B(net110243), .Y(n3543) );
  OAI2BB2X1 U20 ( .B0(\i_MIPS/n191 ), .B1(net110217), .A0N(n11075), .A1N(n176), 
        .Y(\i_MIPS/N34 ) );
  INVX16 U21 ( .A(n1817), .Y(mem_addr_D[10]) );
  INVX16 U22 ( .A(n1822), .Y(mem_addr_D[15]) );
  INVX16 U23 ( .A(n1824), .Y(mem_addr_D[17]) );
  INVX16 U24 ( .A(n1809), .Y(mem_addr_D[23]) );
  MXI2X1 U25 ( .A(n10536), .B(n10535), .S0(n5494), .Y(n10537) );
  AOI222X4 U26 ( .A0(n5480), .A1(n11472), .B0(mem_rdata_D[85]), .B1(n116), 
        .C0(n12976), .C1(n5477), .Y(n10536) );
  BUFX4 U27 ( .A(n10537), .Y(n4272) );
  AO22X4 U28 ( .A0(mem_rdata_I[10]), .A1(n114), .B0(n5469), .B1(n11240), .Y(
        n9669) );
  MX2X1 U29 ( .A(\I_cache/cache[5][74] ), .B(n9673), .S0(n5281), .Y(n12226) );
  MX2X1 U30 ( .A(\I_cache/cache[5][9] ), .B(n9645), .S0(n5282), .Y(n12746) );
  MX2X1 U31 ( .A(\I_cache/cache[4][64] ), .B(n9683), .S0(n5327), .Y(n12307) );
  MX2X1 U32 ( .A(\I_cache/cache[5][90] ), .B(n9711), .S0(n5283), .Y(n12098) );
  MX2X1 U33 ( .A(\I_cache/cache[5][76] ), .B(n10100), .S0(n5277), .Y(n12210)
         );
  MX2X1 U34 ( .A(\I_cache/cache[3][114] ), .B(n10041), .S0(n5195), .Y(n11908)
         );
  MX2X1 U35 ( .A(\I_cache/cache[7][112] ), .B(n10070), .S0(n5371), .Y(n11920)
         );
  MX2X1 U36 ( .A(\I_cache/cache[3][50] ), .B(n10036), .S0(n5195), .Y(n12420)
         );
  MX2X1 U37 ( .A(\I_cache/cache[7][48] ), .B(n10065), .S0(n5371), .Y(n12432)
         );
  MX2X1 U38 ( .A(\I_cache/cache[5][10] ), .B(n9659), .S0(n5279), .Y(n12738) );
  MX2X1 U39 ( .A(\I_cache/cache[5][121] ), .B(n10119), .S0(n5277), .Y(n11850)
         );
  MX2X1 U40 ( .A(\I_cache/cache[5][73] ), .B(n9640), .S0(n5285), .Y(n12234) );
  MX2X1 U41 ( .A(\I_cache/cache[3][16] ), .B(n10060), .S0(n5195), .Y(n12692)
         );
  MX2X1 U42 ( .A(\I_cache/cache[5][12] ), .B(n10085), .S0(n5277), .Y(n12722)
         );
  MX2X1 U43 ( .A(\I_cache/cache[5][105] ), .B(n9650), .S0(n5285), .Y(n11978)
         );
  MX2X1 U44 ( .A(\I_cache/cache[5][44] ), .B(n10090), .S0(n5277), .Y(n12466)
         );
  MX2X1 U45 ( .A(\I_cache/cache[7][82] ), .B(n10046), .S0(n5371), .Y(n12160)
         );
  MX2X1 U46 ( .A(\I_cache/cache[7][5] ), .B(n9541), .S0(n5373), .Y(n12776) );
  MX2X1 U47 ( .A(\I_cache/cache[3][80] ), .B(n10075), .S0(n5195), .Y(n12180)
         );
  OAI2BB2X1 U48 ( .B0(\i_MIPS/n205 ), .B1(net110225), .A0N(n10343), .A1N(n175), 
        .Y(\i_MIPS/N48 ) );
  MX2X1 U49 ( .A(\I_cache/cache[5][108] ), .B(n10095), .S0(n5277), .Y(n11954)
         );
  MX2X1 U50 ( .A(\I_cache/cache[5][25] ), .B(n10109), .S0(n5277), .Y(n12618)
         );
  MX2X1 U51 ( .A(\I_cache/cache[7][31] ), .B(n11035), .S0(n5368), .Y(n12568)
         );
  MX2X1 U52 ( .A(\I_cache/cache[7][97] ), .B(n9361), .S0(n5368), .Y(n12040) );
  AND4X8 U53 ( .A(n10254), .B(net110227), .C(n10389), .D(n10253), .Y(n3726) );
  INVX16 U54 ( .A(n10386), .Y(n10254) );
  OAI222X2 U55 ( .A0(\i_MIPS/PC/n23 ), .A1(net110213), .B0(n4533), .B1(
        net110241), .C0(n11027), .C1(net110247), .Y(n11033) );
  OAI222X2 U56 ( .A0(\i_MIPS/PC/n18 ), .A1(net110215), .B0(n4535), .B1(
        net110241), .C0(net110249), .C1(n10928), .Y(n10933) );
  OAI222X2 U57 ( .A0(\i_MIPS/PC/n25 ), .A1(net110213), .B0(n4557), .B1(
        net110241), .C0(n10967), .C1(net110247), .Y(n10973) );
  CLKINVX16 U58 ( .A(net110253), .Y(net110247) );
  AOI2BB2X2 U59 ( .B0(\i_MIPS/IF_ID[88] ), .B1(n147), .A0N(net110191), .A1N(
        \i_MIPS/n203 ), .Y(n10971) );
  AOI2BB2X2 U60 ( .B0(\i_MIPS/IF_ID[81] ), .B1(n150), .A0N(net110191), .A1N(
        \i_MIPS/n196 ), .Y(n10931) );
  AO22X1 U61 ( .A0(n3647), .A1(mem_read_I), .B0(n4795), .B1(n11365), .Y(n12837) );
  AOI2BB2X4 U62 ( .B0(\i_MIPS/IF_ID[86] ), .B1(n149), .A0N(net110191), .A1N(
        \i_MIPS/n201 ), .Y(n11031) );
  NAND3BX1 U63 ( .AN(n3731), .B(net114031), .C(net98881), .Y(n10863) );
  INVXL U64 ( .A(n11373), .Y(n4322) );
  INVX4 U65 ( .A(n10908), .Y(n10919) );
  OAI2BB2X1 U66 ( .B0(\i_MIPS/n185 ), .B1(net110217), .A0N(n11050), .A1N(n173), 
        .Y(\i_MIPS/N28 ) );
  BUFX16 U67 ( .A(n11201), .Y(n5474) );
  OAI2BB2X1 U68 ( .B0(\i_MIPS/n193 ), .B1(net110217), .A0N(n11085), .A1N(n174), 
        .Y(\i_MIPS/N36 ) );
  NAND3BX4 U69 ( .AN(n10341), .B(n10340), .C(n10339), .Y(\i_MIPS/PC/n59 ) );
  AOI2BB2X2 U70 ( .B0(\i_MIPS/IF_ID[90] ), .B1(n147), .A0N(net110189), .A1N(
        \i_MIPS/n205 ), .Y(n10339) );
  NAND3BX4 U71 ( .AN(n10947), .B(n10946), .C(n10945), .Y(\i_MIPS/PC/n52 ) );
  AOI2BB2X2 U72 ( .B0(\i_MIPS/IF_ID[83] ), .B1(n147), .A0N(net110191), .A1N(
        \i_MIPS/n198 ), .Y(n10945) );
  NAND3BX4 U73 ( .AN(n11082), .B(n11081), .C(n11080), .Y(\i_MIPS/PC/n45 ) );
  AOI2BB2X2 U74 ( .B0(\i_MIPS/IF_ID[76] ), .B1(n148), .A0N(net110191), .A1N(
        \i_MIPS/n191 ), .Y(n11080) );
  AOI221X2 U75 ( .A0(n4924), .A1(n7098), .B0(n3289), .B1(n9258), .C0(n4800), 
        .Y(n7118) );
  AND2X4 U76 ( .A(n4170), .B(n7193), .Y(n3289) );
  INVX4 U77 ( .A(n6062), .Y(n10623) );
  CLKBUFX16 U78 ( .A(net100093), .Y(net112607) );
  CLKINVX1 U79 ( .A(net99078), .Y(net102900) );
  INVX3 U80 ( .A(n4796), .Y(n4348) );
  INVX12 U81 ( .A(n3999), .Y(mem_wdata_I[116]) );
  AO22X4 U82 ( .A0(net113455), .A1(n11425), .B0(net113461), .B1(n11394), .Y(
        n7410) );
  INVX4 U83 ( .A(net100044), .Y(n4084) );
  CLKBUFX20 U84 ( .A(net100093), .Y(n3709) );
  NAND4X6 U85 ( .A(n4091), .B(n4092), .C(n4093), .D(n4094), .Y(n4090) );
  NAND3BX1 U86 ( .AN(n8254), .B(n8927), .C(n8923), .Y(n8255) );
  CLKINVX3 U87 ( .A(n8923), .Y(n8281) );
  OAI211X2 U88 ( .A0(n8927), .A1(n8332), .B0(n8331), .C0(n8330), .Y(n8427) );
  NAND3X6 U89 ( .A(n3712), .B(n3713), .C(net103392), .Y(n4135) );
  CLKINVX8 U90 ( .A(net99087), .Y(net102745) );
  NAND4X8 U91 ( .A(n3689), .B(n8826), .C(n8825), .D(n8824), .Y(net99087) );
  INVX6 U92 ( .A(n10895), .Y(n10901) );
  OAI2BB2X1 U93 ( .B0(\i_MIPS/n220 ), .B1(net110227), .A0N(n174), .A1N(n10895), 
        .Y(\i_MIPS/N63 ) );
  NAND4X8 U94 ( .A(n9687), .B(n9686), .C(n9685), .D(n9684), .Y(n10895) );
  INVX3 U95 ( .A(net99313), .Y(net104705) );
  CLKINVX1 U96 ( .A(n7859), .Y(n84) );
  NAND2X1 U97 ( .A(n4518), .B(n7777), .Y(n7859) );
  INVX6 U98 ( .A(net99267), .Y(net104525) );
  MXI2X2 U99 ( .A(n8066), .B(n8065), .S0(n5587), .Y(n3853) );
  NAND4X4 U100 ( .A(n4102), .B(n4101), .C(n4104), .D(n4103), .Y(n4088) );
  BUFX8 U101 ( .A(n6231), .Y(n4320) );
  OA22X2 U102 ( .A0(net112483), .A1(n933), .B0(net112359), .B1(n2457), .Y(
        n8391) );
  INVX1 U103 ( .A(n6046), .Y(n10638) );
  NAND2X2 U104 ( .A(n10638), .B(n10639), .Y(n6047) );
  NAND2X2 U105 ( .A(n12957), .B(n6144), .Y(n3758) );
  CLKAND2X2 U106 ( .A(n10883), .B(n10882), .Y(n4510) );
  CLKINVX6 U107 ( .A(n10883), .Y(n10272) );
  NAND4X6 U108 ( .A(n9562), .B(n9564), .C(n9563), .D(n9565), .Y(n3631) );
  OAI211X2 U109 ( .A0(n9000), .A1(n9275), .B0(n8999), .C0(n4501), .Y(n9012) );
  INVX8 U110 ( .A(n7957), .Y(n8073) );
  INVX4 U111 ( .A(n6060), .Y(n10624) );
  OAI2BB1X4 U112 ( .A0N(n4517), .A1N(n4707), .B0(n7476), .Y(n8274) );
  INVX3 U113 ( .A(n6567), .Y(n6568) );
  BUFX4 U114 ( .A(n6568), .Y(n161) );
  INVX8 U115 ( .A(net98929), .Y(net104831) );
  OA22X1 U116 ( .A0(\i_MIPS/n356 ), .A1(n4826), .B0(\i_MIPS/n355 ), .B1(n4818), 
        .Y(n7870) );
  CLKINVX16 U117 ( .A(n4827), .Y(n4826) );
  NOR4BX2 U118 ( .AN(n7979), .B(n7976), .C(n7977), .D(n7978), .Y(n7985) );
  OAI222X2 U119 ( .A0(n7969), .A1(n9007), .B0(n141), .B1(n9269), .C0(n9287), 
        .C1(n8534), .Y(n7977) );
  BUFX16 U120 ( .A(n5319), .Y(n5318) );
  AND2X2 U121 ( .A(n8914), .B(n3636), .Y(n48) );
  BUFX8 U122 ( .A(n4470), .Y(n3636) );
  AND2X4 U123 ( .A(n8916), .B(n8915), .Y(n47) );
  BUFX6 U124 ( .A(net99307), .Y(n2) );
  OAI221X2 U125 ( .A0(n7869), .A1(n7365), .B0(n4802), .B1(n7364), .C0(n7789), 
        .Y(n3) );
  MX2X6 U126 ( .A(n6764), .B(n6777), .S0(n5590), .Y(n7364) );
  OAI221X1 U127 ( .A0(n7869), .A1(n7365), .B0(n4802), .B1(n7364), .C0(n7789), 
        .Y(n8535) );
  OR2X2 U128 ( .A(n7672), .B(net102087), .Y(n3629) );
  AND3X6 U129 ( .A(n6296), .B(n6295), .C(n6294), .Y(n6297) );
  INVX4 U130 ( .A(n6056), .Y(n10627) );
  NAND4X4 U131 ( .A(n6076), .B(n6075), .C(n6074), .D(n6073), .Y(n6112) );
  OA21X2 U132 ( .A0(n9615), .A1(n5453), .B0(n9614), .Y(n9622) );
  CLKBUFX6 U133 ( .A(n3631), .Y(n5453) );
  CLKINVX1 U134 ( .A(n10247), .Y(n10221) );
  NAND3X6 U135 ( .A(n4404), .B(n4405), .C(n4406), .Y(n10260) );
  NOR4X8 U136 ( .A(n4118), .B(n4116), .C(n4115), .D(n4117), .Y(net102397) );
  NAND2X4 U137 ( .A(n3203), .B(net98932), .Y(n4114) );
  NAND4X4 U138 ( .A(n8270), .B(n8269), .C(n8268), .D(n8267), .Y(n8278) );
  NAND3X6 U139 ( .A(n4167), .B(n4166), .C(n9210), .Y(n3861) );
  NAND2X4 U140 ( .A(n4605), .B(n10731), .Y(net102183) );
  INVX3 U141 ( .A(n6088), .Y(n10653) );
  OAI221X1 U142 ( .A0(net112655), .A1(n254), .B0(net112589), .B1(n204), .C0(
        n6087), .Y(n6088) );
  NAND4X8 U143 ( .A(n6099), .B(n6096), .C(n6097), .D(n6098), .Y(n6111) );
  NAND2X4 U144 ( .A(n10656), .B(n10655), .Y(n6095) );
  AND2X1 U145 ( .A(n9002), .B(n4470), .Y(n3786) );
  AND3X4 U146 ( .A(n4471), .B(n6263), .C(n6447), .Y(n4470) );
  AND2X8 U147 ( .A(net134117), .B(net99734), .Y(n4532) );
  NAND4X6 U148 ( .A(n4098), .B(n4097), .C(n4096), .D(n4095), .Y(n4089) );
  CLKBUFX8 U149 ( .A(net110229), .Y(net110213) );
  BUFX16 U150 ( .A(net112143), .Y(net112139) );
  XNOR2X4 U151 ( .A(n6068), .B(n4), .Y(n6069) );
  CLKINVX20 U152 ( .A(DCACHE_addr[17]), .Y(n4) );
  AND3X6 U153 ( .A(n4496), .B(n6208), .C(\i_MIPS/ALU_Control/n20 ), .Y(n4495)
         );
  NAND2BX1 U154 ( .AN(\i_MIPS/ALUOp[1] ), .B(n4413), .Y(n6208) );
  XNOR2X4 U155 ( .A(n6063), .B(n5), .Y(n6070) );
  NAND2X8 U156 ( .A(n10621), .B(n10620), .Y(n6068) );
  INVX8 U157 ( .A(n11186), .Y(n6) );
  INVX12 U158 ( .A(n11185), .Y(n11186) );
  BUFX12 U159 ( .A(n4514), .Y(n5473) );
  INVX2 U160 ( .A(n10568), .Y(n8995) );
  OAI222X2 U161 ( .A0(\i_MIPS/PC/n29 ), .A1(net110215), .B0(n4530), .B1(
        net110241), .C0(n10369), .C1(n3602), .Y(n10374) );
  AOI222X1 U162 ( .A0(n5480), .A1(n11473), .B0(mem_rdata_D[86]), .B1(n116), 
        .C0(n12975), .C1(n5477), .Y(n10548) );
  BUFX12 U163 ( .A(n11205), .Y(n5480) );
  INVX20 U164 ( .A(n4130), .Y(net110241) );
  NAND3BX2 U165 ( .AN(n10313), .B(n10910), .C(n10912), .Y(n10883) );
  AND3X6 U166 ( .A(n10912), .B(n10911), .C(n10910), .Y(n10914) );
  OR2X2 U167 ( .A(n4542), .B(net110243), .Y(n3655) );
  OA22X2 U168 ( .A0(n11030), .A1(net140280), .B0(net98430), .B1(n11029), .Y(
        n11032) );
  OA22X2 U169 ( .A0(n10338), .A1(net140280), .B0(net98430), .B1(n10342), .Y(
        n10340) );
  OA22X2 U170 ( .A0(n10371), .A1(net140280), .B0(net98430), .B1(n10380), .Y(
        n10373) );
  NAND3X4 U171 ( .A(n3763), .B(n3764), .C(n3765), .Y(n11116) );
  OR2X2 U172 ( .A(n4560), .B(net110243), .Y(n3764) );
  CLKINVX12 U173 ( .A(n9569), .Y(n9553) );
  NOR4X1 U174 ( .A(n9566), .B(n9568), .C(n9569), .D(n5984), .Y(n6037) );
  NOR4X2 U175 ( .A(n9567), .B(n9568), .C(n9569), .D(n9566), .Y(n9590) );
  AO22X2 U176 ( .A0(net113447), .A1(n11456), .B0(net102346), .B1(n11487), .Y(
        n7409) );
  CLKMX2X4 U177 ( .A(n7140), .B(n7139), .S0(n5588), .Y(net105824) );
  NOR2X1 U178 ( .A(n6032), .B(n6035), .Y(n29) );
  NAND4X1 U179 ( .A(n4696), .B(n9582), .C(n4042), .D(n4694), .Y(n6032) );
  CLKBUFX3 U180 ( .A(n4966), .Y(n4968) );
  AO22XL U181 ( .A0(n4973), .A1(n215), .B0(n4966), .B1(n716), .Y(n7677) );
  INVX6 U182 ( .A(net99384), .Y(net103708) );
  NOR2X4 U183 ( .A(n3562), .B(n9016), .Y(n4410) );
  NAND2X6 U184 ( .A(n3533), .B(n9020), .Y(net99971) );
  BUFX4 U185 ( .A(net112505), .Y(net112459) );
  NAND4X4 U186 ( .A(n9240), .B(n9239), .C(n9238), .D(n9237), .Y(n11512) );
  OAI221X4 U187 ( .A0(net112663), .A1(n2047), .B0(net112561), .B1(n707), .C0(
        n6135), .Y(n6136) );
  BUFX16 U188 ( .A(net112589), .Y(net112561) );
  BUFX8 U189 ( .A(n4691), .Y(n4828) );
  CLKAND2X2 U190 ( .A(n4815), .B(\i_MIPS/n356 ), .Y(n4600) );
  INVX3 U191 ( .A(n8253), .Y(n8328) );
  NAND2X6 U192 ( .A(n10624), .B(n10623), .Y(n6063) );
  BUFX16 U193 ( .A(net111979), .Y(net111915) );
  NAND2X2 U194 ( .A(n6565), .B(\i_MIPS/n344 ), .Y(n8646) );
  INVX8 U195 ( .A(n103), .Y(n6565) );
  INVX6 U196 ( .A(n9184), .Y(n9180) );
  AO22X1 U197 ( .A0(net113447), .A1(n11462), .B0(net102346), .B1(n11493), .Y(
        n7157) );
  AOI222X4 U198 ( .A0(n5474), .A1(n11493), .B0(mem_rdata_D[107]), .B1(n117), 
        .C0(n12986), .C1(n5473), .Y(n10778) );
  NAND4X2 U199 ( .A(n7156), .B(n7155), .C(n7154), .D(n7153), .Y(n11493) );
  OA22X2 U200 ( .A0(\i_MIPS/Register/register[6][10] ), .A1(n4936), .B0(
        \i_MIPS/Register/register[14][10] ), .B1(n4930), .Y(n7249) );
  BUFX2 U201 ( .A(net102300), .Y(net113169) );
  MXI2XL U202 ( .A(\i_MIPS/n356 ), .B(n4536), .S0(n5510), .Y(\i_MIPS/n547 ) );
  CLKBUFX3 U203 ( .A(n11139), .Y(n5409) );
  INVX16 U204 ( .A(n5460), .Y(n5456) );
  BUFX20 U205 ( .A(n3848), .Y(n5460) );
  NAND2BX2 U206 ( .AN(n5454), .B(n11299), .Y(n9629) );
  NAND2X6 U207 ( .A(n11188), .B(n6), .Y(net139669) );
  AO22X1 U208 ( .A0(\i_MIPS/IF_ID[67] ), .A1(n11186), .B0(\i_MIPS/IF_ID_2 ), 
        .B1(n11185), .Y(n11187) );
  INVX3 U209 ( .A(n7788), .Y(n7790) );
  OAI2BB2X4 U210 ( .B0(n7783), .B1(n7867), .A0N(n7785), .A1N(n7784), .Y(n7788)
         );
  INVX6 U211 ( .A(n3548), .Y(n4020) );
  NAND2X4 U212 ( .A(n4515), .B(n4801), .Y(n8513) );
  AOI33X2 U213 ( .A0(n7803), .A1(n7802), .A2(n9258), .B0(n7801), .B1(n7800), 
        .B2(n9258), .Y(n7804) );
  AO22X2 U214 ( .A0(n4809), .A1(\i_MIPS/ALUin1[1] ), .B0(n4814), .B1(
        \i_MIPS/ALUin1[0] ), .Y(n7693) );
  CLKBUFX12 U215 ( .A(n4631), .Y(n4809) );
  INVX4 U216 ( .A(net99461), .Y(net105426) );
  MX2X1 U217 ( .A(\D_cache/cache[0][5] ), .B(n10754), .S0(net112645), .Y(
        \D_cache/n1756 ) );
  MX2X1 U218 ( .A(\D_cache/cache[1][5] ), .B(n10754), .S0(net112543), .Y(
        \D_cache/n1755 ) );
  MX2X1 U219 ( .A(\D_cache/cache[7][5] ), .B(n10754), .S0(net111883), .Y(
        \D_cache/n1749 ) );
  MX2X1 U220 ( .A(\D_cache/cache[6][5] ), .B(n10754), .S0(net112009), .Y(
        \D_cache/n1750 ) );
  MX2X1 U221 ( .A(\D_cache/cache[5][5] ), .B(n10754), .S0(net112131), .Y(
        \D_cache/n1751 ) );
  MX2X1 U222 ( .A(\D_cache/cache[4][5] ), .B(n10754), .S0(net112211), .Y(
        \D_cache/n1752 ) );
  MX2X1 U223 ( .A(\D_cache/cache[3][5] ), .B(n10754), .S0(net112295), .Y(
        \D_cache/n1753 ) );
  MX2X1 U224 ( .A(\D_cache/cache[2][5] ), .B(n10754), .S0(net112419), .Y(
        \D_cache/n1754 ) );
  NAND2X2 U225 ( .A(n10751), .B(n10750), .Y(net140444) );
  INVX6 U226 ( .A(net99605), .Y(net103391) );
  CLKINVX8 U227 ( .A(n6235), .Y(n6233) );
  AO22X2 U228 ( .A0(net113447), .A1(n11479), .B0(net102346), .B1(n11510), .Y(
        n9060) );
  BUFX16 U229 ( .A(n11103), .Y(n4724) );
  BUFX6 U230 ( .A(n5187), .Y(n5164) );
  BUFX16 U231 ( .A(n5144), .Y(n5187) );
  BUFX16 U232 ( .A(net99330), .Y(n152) );
  NAND2X6 U233 ( .A(n3315), .B(net99316), .Y(n3663) );
  NOR2BX4 U234 ( .AN(n4815), .B(\i_MIPS/n341 ), .Y(n4682) );
  BUFX12 U235 ( .A(n4627), .Y(n4815) );
  NAND2X6 U236 ( .A(net98973), .B(net98974), .Y(n4119) );
  NAND2X8 U237 ( .A(n4641), .B(n3826), .Y(n4419) );
  NAND2X8 U238 ( .A(n6230), .B(\i_MIPS/n362 ), .Y(n7180) );
  AND2X6 U239 ( .A(net134133), .B(net99293), .Y(n4560) );
  OA22X1 U240 ( .A0(net112061), .A1(n1512), .B0(net111937), .B1(n3125), .Y(
        n7726) );
  AND3X4 U241 ( .A(\i_MIPS/ID_EX[78] ), .B(\i_MIPS/ID_EX[73] ), .C(
        \i_MIPS/ID_EX[75] ), .Y(n4714) );
  MX2X4 U242 ( .A(\i_MIPS/ID_EX[75] ), .B(n4641), .S0(n3768), .Y(n6211) );
  NAND2X6 U243 ( .A(n10635), .B(n10634), .Y(n6042) );
  NAND3X4 U244 ( .A(n43), .B(n44), .C(net106110), .Y(net99576) );
  OAI222X4 U245 ( .A0(n8538), .A1(n7544), .B0(n8659), .B1(n7359), .C0(n8817), 
        .C1(n7353), .Y(n7372) );
  OAI221X4 U246 ( .A0(n8540), .A1(n8539), .B0(n8538), .B1(n8537), .C0(n4501), 
        .Y(n8550) );
  OA22X1 U247 ( .A0(n8726), .A1(n9006), .B0(n8538), .B1(n8729), .Y(n6266) );
  BUFX12 U248 ( .A(n4692), .Y(n4822) );
  CLKBUFX8 U249 ( .A(n4692), .Y(n4823) );
  CLKBUFX12 U250 ( .A(n4692), .Y(n4821) );
  BUFX16 U251 ( .A(n4692), .Y(n4820) );
  CLKAND2X4 U252 ( .A(n3524), .B(\i_MIPS/ID_EX[80] ), .Y(n4691) );
  CLKINVX6 U253 ( .A(n41), .Y(n42) );
  INVX16 U254 ( .A(net113081), .Y(net113075) );
  CLKXOR2X1 U255 ( .A(n6293), .B(\i_MIPS/IR_ID[22] ), .Y(n6294) );
  NAND3X6 U256 ( .A(n61), .B(n62), .C(n63), .Y(n64) );
  INVX4 U257 ( .A(n10312), .Y(n63) );
  NAND2X8 U258 ( .A(n64), .B(n10311), .Y(n10315) );
  AND3X6 U259 ( .A(n10316), .B(n10935), .C(n4590), .Y(n3635) );
  OA22X4 U260 ( .A0(n5248), .A1(n3224), .B0(n5203), .B1(n1585), .Y(n4466) );
  AO22X4 U261 ( .A0(net113455), .A1(n11424), .B0(net113461), .B1(n11393), .Y(
        n8779) );
  BUFX4 U262 ( .A(net102372), .Y(net113461) );
  MX2X1 U263 ( .A(n3486), .B(net99064), .S0(n5510), .Y(\i_MIPS/n427 ) );
  INVX6 U264 ( .A(n5376), .Y(n3617) );
  CLKBUFX4 U265 ( .A(n5449), .Y(n5420) );
  NAND2X6 U266 ( .A(\i_MIPS/ALUin1[13] ), .B(n6351), .Y(n6936) );
  CLKMX2X12 U267 ( .A(\i_MIPS/n283 ), .B(n4709), .S0(n3826), .Y(n6351) );
  CLKAND2X3 U268 ( .A(n6464), .B(n6473), .Y(n6468) );
  INVX8 U269 ( .A(n6636), .Y(n8249) );
  NAND2X4 U270 ( .A(n6583), .B(\i_MIPS/n348 ), .Y(n8891) );
  INVX3 U271 ( .A(n10942), .Y(n3846) );
  INVX8 U272 ( .A(n10212), .Y(n10872) );
  NAND4X6 U273 ( .A(n7891), .B(n7889), .C(n7890), .D(n7888), .Y(net99290) );
  NOR4BX4 U274 ( .AN(n3612), .B(n7883), .C(n7882), .D(n7881), .Y(n7889) );
  AOI2BB1X4 U275 ( .A0N(\i_MIPS/n347 ), .A1N(n4818), .B0(n4666), .Y(n6950) );
  OAI222X4 U276 ( .A0(n7869), .A1(n7868), .B0(n7867), .B1(n7866), .C0(n7865), 
        .C1(n4797), .Y(n7873) );
  NAND3X2 U277 ( .A(n31), .B(n32), .C(n6953), .Y(n7865) );
  BUFX20 U278 ( .A(net138398), .Y(n3671) );
  AO22X1 U279 ( .A0(net113455), .A1(n11433), .B0(net113461), .B1(n11402), .Y(
        n6394) );
  NAND4X2 U280 ( .A(net105008), .B(net105009), .C(net105010), .D(net105011), 
        .Y(net98089) );
  NAND4X8 U281 ( .A(net99845), .B(n10257), .C(n10256), .D(n4494), .Y(n10813)
         );
  NAND3X2 U282 ( .A(net99849), .B(net98881), .C(\i_MIPS/IF_ID[64] ), .Y(n79)
         );
  INVX3 U283 ( .A(n8432), .Y(n6651) );
  AOI2BB2X4 U284 ( .B0(net113039), .B1(net99078), .A0N(net102087), .A1N(n3614), 
        .Y(n3613) );
  OAI211XL U285 ( .A0(n6668), .A1(n9275), .B0(n6667), .C0(n4501), .Y(n6681) );
  NAND2X4 U286 ( .A(n6666), .B(n9170), .Y(n6661) );
  NAND2X6 U287 ( .A(n4654), .B(n4583), .Y(n9223) );
  MXI2X2 U288 ( .A(n8761), .B(n8760), .S0(n5587), .Y(n3614) );
  OAI2BB2X4 U289 ( .B0(\i_MIPS/n176 ), .B1(net110227), .A0N(n174), .A1N(n4543), 
        .Y(\i_MIPS/N117 ) );
  NAND2X1 U290 ( .A(n9364), .B(ICACHE_addr[15]), .Y(n9365) );
  NAND3BX4 U291 ( .AN(n10949), .B(n10487), .C(n10325), .Y(n10318) );
  NAND4X2 U292 ( .A(n10099), .B(n10098), .C(n10097), .D(n10096), .Y(n11274) );
  BUFX12 U293 ( .A(n3722), .Y(net112161) );
  INVX3 U294 ( .A(net99110), .Y(net105151) );
  INVX8 U295 ( .A(net112121), .Y(n3722) );
  CLKINVX2 U296 ( .A(n3754), .Y(n3836) );
  CLKINVX2 U297 ( .A(n3836), .Y(n3808) );
  OAI2BB1X2 U298 ( .A0N(n7547), .A1N(n7546), .B0(n3670), .Y(n7456) );
  AO21X2 U299 ( .A0(n8806), .A1(n8823), .B0(n8812), .Y(n8716) );
  AND3X8 U300 ( .A(n4599), .B(n10499), .C(n10498), .Y(n10502) );
  CLKXOR2X2 U301 ( .A(n9363), .B(ICACHE_addr[20]), .Y(n10959) );
  NAND2X2 U302 ( .A(n10317), .B(net113551), .Y(n10323) );
  INVX4 U303 ( .A(n10959), .Y(n10317) );
  NAND4X6 U304 ( .A(n5960), .B(n5959), .C(n5958), .D(n5957), .Y(n3565) );
  AOI211X2 U305 ( .A0(n3590), .A1(n11233), .B0(n11050), .C0(n4549), .Y(n9623)
         );
  CLKINVX2 U306 ( .A(n151), .Y(n10886) );
  OAI221X2 U307 ( .A0(net105425), .A1(net112709), .B0(net105426), .B1(
        net112723), .C0(net105427), .Y(net99064) );
  AO21X2 U308 ( .A0(net100038), .A1(net100039), .B0(net113077), .Y(net100035)
         );
  NAND2X2 U309 ( .A(n11095), .B(n11093), .Y(n10907) );
  INVX6 U310 ( .A(n11093), .Y(n11099) );
  NAND3X4 U311 ( .A(n3531), .B(n8069), .C(n8252), .Y(n3532) );
  CLKINVX3 U312 ( .A(n3772), .Y(n3531) );
  NAND3BX4 U313 ( .AN(n9015), .B(n9258), .C(n9016), .Y(n9021) );
  NAND2X8 U314 ( .A(\i_MIPS/ALUin1[18] ), .B(n161), .Y(n8516) );
  INVX6 U315 ( .A(net106977), .Y(net98970) );
  NAND2X4 U316 ( .A(n6592), .B(\i_MIPS/n347 ), .Y(n9156) );
  INVX8 U317 ( .A(n10306), .Y(n10211) );
  OAI2BB2X1 U318 ( .B0(\i_MIPS/n164 ), .B1(net110217), .A0N(n173), .A1N(n11111), .Y(\i_MIPS/N105 ) );
  INVX2 U319 ( .A(n11112), .Y(n11111) );
  NAND2X6 U320 ( .A(\i_MIPS/ALUin1[22] ), .B(n6582), .Y(n8922) );
  INVX12 U321 ( .A(n6585), .Y(n6582) );
  NAND3X4 U322 ( .A(n8934), .B(n8932), .C(n74), .Y(n10568) );
  INVX4 U323 ( .A(n73), .Y(n74) );
  CLKINVX12 U324 ( .A(n9284), .Y(n9130) );
  OAI221X2 U325 ( .A0(n7869), .A1(n7286), .B0(n4802), .B1(n8083), .C0(n7789), 
        .Y(n8084) );
  CLKINVX8 U326 ( .A(\i_MIPS/ID_EX[80] ), .Y(n9272) );
  INVX4 U327 ( .A(n7285), .Y(n7875) );
  NAND2X4 U328 ( .A(n4802), .B(n5589), .Y(n7285) );
  BUFX20 U329 ( .A(net138398), .Y(n3672) );
  NAND4X4 U330 ( .A(n8684), .B(n8683), .C(n8682), .D(n8681), .Y(n11478) );
  BUFX6 U331 ( .A(net112599), .Y(net112587) );
  AND2X8 U332 ( .A(n3613), .B(net99450), .Y(n4134) );
  NAND4X4 U333 ( .A(n8854), .B(n8853), .C(n8852), .D(n8851), .Y(n11392) );
  NAND2X4 U334 ( .A(n6252), .B(n6251), .Y(n3597) );
  NAND2X1 U335 ( .A(n7545), .B(n7454), .Y(n3668) );
  NAND2X4 U336 ( .A(n6571), .B(\i_MIPS/n355 ), .Y(n8150) );
  INVX3 U337 ( .A(n8150), .Y(n8146) );
  OAI2BB1X4 U338 ( .A0N(net99637), .A1N(net99638), .B0(net114085), .Y(
        net103220) );
  NAND4X4 U339 ( .A(n8585), .B(n8584), .C(n8583), .D(n8582), .Y(n11440) );
  CLKMX2X4 U340 ( .A(\i_MIPS/n279 ), .B(n3310), .S0(n3826), .Y(n6613) );
  MX2X2 U341 ( .A(\i_MIPS/n279 ), .B(n3310), .S0(n3826), .Y(n167) );
  NAND4X6 U342 ( .A(n4081), .B(n4079), .C(n4080), .D(n4082), .Y(n4072) );
  AOI222X1 U343 ( .A0(n5475), .A1(n11488), .B0(mem_rdata_D[101]), .B1(n116), 
        .C0(n12992), .C1(n5473), .Y(n10753) );
  NAND4X4 U344 ( .A(n7330), .B(n7329), .C(n7328), .D(n7327), .Y(n11488) );
  INVX3 U345 ( .A(n6044), .Y(n10639) );
  OAI221X2 U346 ( .A0(net112651), .A1(n280), .B0(net112593), .B1(n1231), .C0(
        n6043), .Y(n6044) );
  INVX20 U347 ( .A(net113532), .Y(net108204) );
  BUFX20 U348 ( .A(n3751), .Y(net113540) );
  BUFX12 U349 ( .A(net130594), .Y(net109801) );
  CLKAND2X8 U350 ( .A(n10161), .B(n4589), .Y(net130594) );
  INVX3 U351 ( .A(n6779), .Y(n6436) );
  CLKMX2X4 U352 ( .A(n9141), .B(n4799), .S0(n6433), .Y(n6434) );
  OAI221X4 U353 ( .A0(\i_MIPS/ALUin1[13] ), .A1(n4810), .B0(
        \i_MIPS/ALUin1[12] ), .B1(n4803), .C0(n6261), .Y(n6431) );
  AOI2BB2X2 U354 ( .B0(n4796), .B1(n11366), .A0N(n3646), .A1N(n4324), .Y(n3865) );
  OR2X8 U355 ( .A(n10939), .B(n10938), .Y(n4157) );
  MX2X2 U356 ( .A(n6777), .B(n7365), .S0(n5589), .Y(n6778) );
  OA22X4 U357 ( .A0(n7869), .A1(n6777), .B0(n6424), .B1(n4797), .Y(n6425) );
  OAI221X4 U358 ( .A0(\i_MIPS/n346 ), .A1(n4810), .B0(\i_MIPS/n347 ), .B1(
        n4803), .C0(n6259), .Y(n6777) );
  OR2X6 U359 ( .A(n8527), .B(n8526), .Y(n55) );
  NAND2X6 U360 ( .A(n6633), .B(n6632), .Y(n6932) );
  NAND2X6 U361 ( .A(n4436), .B(n4435), .Y(n4437) );
  INVX12 U362 ( .A(n5593), .Y(n4199) );
  INVX8 U363 ( .A(n3577), .Y(n4158) );
  NAND3X8 U364 ( .A(n6643), .B(n6644), .C(n3850), .Y(n6646) );
  INVX3 U365 ( .A(n6634), .Y(n6635) );
  INVX3 U366 ( .A(n8913), .Y(n8915) );
  CLKAND2X8 U367 ( .A(n4813), .B(\i_MIPS/ALUin1[29] ), .Y(n4673) );
  BUFX20 U368 ( .A(n4627), .Y(n4813) );
  NAND3X8 U369 ( .A(n4438), .B(n4439), .C(n9169), .Y(n6664) );
  BUFX8 U370 ( .A(n3839), .Y(net113533) );
  NAND4X8 U371 ( .A(n6159), .B(n6157), .C(n6156), .D(n6158), .Y(n6168) );
  NAND2X4 U372 ( .A(n1608), .B(n3295), .Y(n6144) );
  NOR4X6 U373 ( .A(n6112), .B(n6111), .C(n6109), .D(n6110), .Y(n6171) );
  CLKAND2X12 U374 ( .A(n7183), .B(n7193), .Y(n4617) );
  INVX8 U375 ( .A(n4320), .Y(n6244) );
  NAND2X8 U376 ( .A(n6237), .B(\i_MIPS/n366 ), .Y(n7458) );
  INVX12 U377 ( .A(n7458), .Y(n7287) );
  AOI2BB1X4 U378 ( .A0N(n4007), .A1N(n6769), .B0(n6605), .Y(n6226) );
  NAND2X8 U379 ( .A(n6581), .B(\i_MIPS/n350 ), .Y(n8067) );
  INVX12 U380 ( .A(n6584), .Y(n6581) );
  AND2X4 U381 ( .A(\i_MIPS/ALU_Control/n15 ), .B(\i_MIPS/ALUOp[1] ), .Y(n6210)
         );
  OAI221X4 U382 ( .A0(n8548), .A1(n8886), .B0(n8547), .B1(n8546), .C0(n8545), 
        .Y(n8549) );
  NAND2X6 U383 ( .A(n9130), .B(n4707), .Y(n8886) );
  CLKMX2X2 U384 ( .A(n9280), .B(n9279), .S0(n8544), .Y(n8545) );
  MX2X6 U385 ( .A(\i_MIPS/n285 ), .B(n4708), .S0(n5594), .Y(n6249) );
  NAND2X8 U386 ( .A(n6250), .B(\i_MIPS/ALUin1[12] ), .Y(n6598) );
  AND4X2 U387 ( .A(\i_MIPS/n323 ), .B(\i_MIPS/ALUOp[1] ), .C(
        \i_MIPS/ALU_Control/n11 ), .D(\i_MIPS/ID_EX[106] ), .Y(
        \i_MIPS/ALU_Control/n10 ) );
  CLKINVX6 U388 ( .A(\i_MIPS/ALU_Control/n10 ), .Y(n6220) );
  NAND2X2 U389 ( .A(n3727), .B(n6660), .Y(n3746) );
  NAND2XL U390 ( .A(n3593), .B(net100866), .Y(net98449) );
  NAND2X2 U391 ( .A(n8822), .B(n3787), .Y(n7101) );
  NAND2X6 U392 ( .A(\i_MIPS/ALUin1[7] ), .B(n6239), .Y(n7461) );
  NAND2X8 U393 ( .A(n7461), .B(n6771), .Y(n7181) );
  NAND2X2 U394 ( .A(n7090), .B(n7461), .Y(n6845) );
  NAND2X6 U395 ( .A(n8923), .B(n8922), .Y(n3640) );
  AND3X6 U396 ( .A(n10254), .B(net110227), .C(n10865), .Y(n10246) );
  MX2X8 U397 ( .A(\i_MIPS/n257 ), .B(n4493), .S0(n3826), .Y(n6587) );
  NAND2X2 U398 ( .A(n4550), .B(n8647), .Y(n9153) );
  CLKINVX4 U399 ( .A(n10913), .Y(n10311) );
  OAI2BB1X4 U400 ( .A0N(n11075), .A1N(n11073), .B0(n10265), .Y(n10266) );
  INVX4 U401 ( .A(n5459), .Y(n5458) );
  CLKBUFX8 U402 ( .A(n3848), .Y(n5459) );
  NAND2X6 U403 ( .A(n10671), .B(n10670), .Y(n6139) );
  OAI221X4 U404 ( .A0(net112231), .A1(n1227), .B0(net112137), .B1(n2806), .C0(
        n6137), .Y(n6138) );
  BUFX8 U405 ( .A(n4514), .Y(n5472) );
  INVX20 U406 ( .A(n5460), .Y(n5457) );
  NAND4X6 U407 ( .A(n6006), .B(n6005), .C(n6004), .D(n6003), .Y(n11365) );
  OA22X4 U408 ( .A0(n5249), .A1(n3274), .B0(n5204), .B1(n1618), .Y(n6005) );
  NAND4X8 U409 ( .A(n10055), .B(n10054), .C(n10053), .D(n10052), .Y(n11093) );
  INVX8 U410 ( .A(n4501), .Y(n8089) );
  INVX20 U411 ( .A(n8726), .Y(n8821) );
  CLKINVX1 U412 ( .A(n8643), .Y(n6616) );
  INVX6 U413 ( .A(n7042), .Y(n7708) );
  NAND2XL U414 ( .A(\i_MIPS/ID_EX[100] ), .B(n3826), .Y(n102) );
  MX2X1 U415 ( .A(\i_MIPS/n301 ), .B(n6216), .S0(n3826), .Y(n3790) );
  INVXL U416 ( .A(n3826), .Y(n100) );
  MXI2X1 U417 ( .A(\i_MIPS/n301 ), .B(n6216), .S0(n3826), .Y(n3720) );
  MXI2X6 U418 ( .A(\i_MIPS/ID_EX[50] ), .B(n4802), .S0(n3826), .Y(n6230) );
  NOR3X4 U419 ( .A(n7796), .B(n7797), .C(n3557), .Y(n7805) );
  AOI22X4 U420 ( .A0(n6930), .A1(n1224), .B0(n1224), .B1(n6934), .Y(n6640) );
  NAND4X1 U421 ( .A(n4662), .B(n9548), .C(n4665), .D(n4695), .Y(n9336) );
  INVX16 U422 ( .A(n11361), .Y(n4794) );
  OAI221X1 U423 ( .A0(n7867), .A1(n6764), .B0(n7285), .B1(n7365), .C0(n6425), 
        .Y(n6426) );
  AND4X4 U424 ( .A(n10255), .B(net99855), .C(net110227), .D(n10254), .Y(n4509)
         );
  NAND4X6 U425 ( .A(n4696), .B(n9582), .C(n4042), .D(n4694), .Y(n9583) );
  NAND2BX4 U426 ( .AN(n5457), .B(n11231), .Y(n9601) );
  NAND4X8 U427 ( .A(n9602), .B(n9601), .C(n9600), .D(n9599), .Y(n11044) );
  XOR3X1 U428 ( .A(n10207), .B(n10870), .C(n10212), .Y(n10866) );
  CLKINVX1 U429 ( .A(n11329), .Y(n9615) );
  NAND2X8 U430 ( .A(n11050), .B(n11053), .Y(n11059) );
  NAND4X2 U431 ( .A(n9511), .B(n9510), .C(n9509), .D(n9508), .Y(n11329) );
  NAND2X2 U432 ( .A(n3313), .B(net99974), .Y(n4111) );
  INVX4 U433 ( .A(n7033), .Y(n7032) );
  AOI22X4 U434 ( .A0(net99609), .A1(net113041), .B0(net102300), .B1(n7089), 
        .Y(n3313) );
  NAND4X8 U435 ( .A(n3733), .B(n7049), .C(n7048), .D(n7047), .Y(net99609) );
  NAND4X6 U436 ( .A(n9555), .B(n9554), .C(n3964), .D(n9553), .Y(n9561) );
  AND2X4 U437 ( .A(n3532), .B(n8095), .Y(n3318) );
  OAI31X2 U438 ( .A0(n3772), .A1(n7955), .A2(n7954), .B0(n8095), .Y(n3859) );
  BUFX4 U439 ( .A(n4904), .Y(n4907) );
  CLKBUFX8 U440 ( .A(n4479), .Y(n4904) );
  OA22X1 U441 ( .A0(\i_MIPS/Register/register[22][16] ), .A1(n4913), .B0(
        \i_MIPS/Register/register[30][16] ), .B1(n4907), .Y(n8184) );
  BUFX8 U442 ( .A(n10577), .Y(n4308) );
  MXI2X2 U443 ( .A(n10576), .B(n10575), .S0(n5493), .Y(n10577) );
  NAND2X8 U444 ( .A(n3811), .B(n7950), .Y(n9165) );
  AND3X6 U445 ( .A(n9165), .B(n9168), .C(n2802), .Y(n9176) );
  OAI221X4 U446 ( .A0(n7975), .A1(n9004), .B0(n7974), .B1(n8537), .C0(n7973), 
        .Y(n7976) );
  INVXL U447 ( .A(n7970), .Y(n7975) );
  INVX6 U448 ( .A(n9577), .Y(n9548) );
  NAND3BX2 U449 ( .AN(n9577), .B(n4665), .C(n4662), .Y(n6035) );
  XOR3X2 U450 ( .A(n11050), .B(n11062), .C(n11053), .Y(n11052) );
  NAND3BX4 U451 ( .AN(n7092), .B(n7180), .C(n3766), .Y(n4170) );
  INVX8 U452 ( .A(n10205), .Y(n10269) );
  INVX8 U453 ( .A(n11073), .Y(n11079) );
  CLKINVX12 U454 ( .A(n8729), .Y(n8822) );
  NAND2X8 U455 ( .A(n8148), .B(n4577), .Y(n8729) );
  NAND2X6 U456 ( .A(n6260), .B(n7968), .Y(n8148) );
  INVX6 U457 ( .A(net98952), .Y(net106419) );
  MXI2X4 U458 ( .A(n7783), .B(n7791), .S0(n5590), .Y(n4517) );
  CLKINVX1 U459 ( .A(n7791), .Y(n7108) );
  MXI2X2 U460 ( .A(n4683), .B(n7791), .S0(n3787), .Y(n3666) );
  AND2X6 U461 ( .A(n3218), .B(net100035), .Y(n4086) );
  OAI211X4 U462 ( .A0(n9137), .A1(n8444), .B0(n8443), .C0(n8442), .Y(n8445) );
  NAND4X2 U463 ( .A(n4743), .B(n8440), .C(n9259), .D(n9156), .Y(n8443) );
  INVX12 U464 ( .A(n6664), .Y(n9015) );
  NAND2X4 U465 ( .A(n3757), .B(n3758), .Y(n6159) );
  MXI2X2 U466 ( .A(n10563), .B(n10562), .S0(n5493), .Y(n10564) );
  BUFX8 U467 ( .A(n10564), .Y(n4309) );
  CLKINVX16 U468 ( .A(n4509), .Y(n172) );
  NAND2X6 U469 ( .A(n8152), .B(n8143), .Y(n7704) );
  OR2X2 U470 ( .A(net100082), .B(n1990), .Y(n3798) );
  NAND3X6 U471 ( .A(n3798), .B(n3799), .C(n6057), .Y(n6058) );
  MXI2X2 U472 ( .A(n10551), .B(n10550), .S0(n5493), .Y(n10552) );
  BUFX8 U473 ( .A(n10552), .Y(n4310) );
  NAND3X4 U474 ( .A(n3542), .B(n3543), .C(n3544), .Y(n10892) );
  NAND3BX4 U475 ( .AN(n10892), .B(n10891), .C(n10890), .Y(\i_MIPS/PC/n43 ) );
  INVX20 U476 ( .A(net110205), .Y(net140280) );
  BUFX4 U477 ( .A(n10962), .Y(n153) );
  OAI221X2 U478 ( .A0(n7867), .A1(n7365), .B0(n4797), .B1(n6777), .C0(n7476), 
        .Y(n8910) );
  AND2X4 U479 ( .A(\i_MIPS/ID_EX[80] ), .B(n3525), .Y(n4692) );
  AND3X4 U480 ( .A(n4663), .B(n9547), .C(n4695), .Y(n9565) );
  INVX4 U481 ( .A(n10314), .Y(n61) );
  NAND2BX4 U482 ( .AN(n5453), .B(n11331), .Y(n9627) );
  NAND2X6 U483 ( .A(n4175), .B(n4177), .Y(n37) );
  OR2X6 U484 ( .A(net110251), .B(n10285), .Y(n4177) );
  NAND2X6 U485 ( .A(n38), .B(n4176), .Y(n10288) );
  NAND3X2 U486 ( .A(n89), .B(n90), .C(n91), .Y(n8277) );
  OAI221X2 U487 ( .A0(n4798), .A1(n8716), .B0(n4552), .B1(n9262), .C0(n8805), 
        .Y(n8721) );
  NOR4X6 U488 ( .A(n9586), .B(n9585), .C(n9584), .D(n9583), .Y(n9587) );
  INVX8 U489 ( .A(n10884), .Y(n10889) );
  INVX12 U490 ( .A(n10813), .Y(n11188) );
  OR2X4 U491 ( .A(n10814), .B(n10813), .Y(n4192) );
  NAND2X6 U492 ( .A(n10629), .B(n3621), .Y(n4167) );
  NAND2X4 U493 ( .A(n80), .B(net98880), .Y(n10257) );
  NAND2X8 U494 ( .A(n4210), .B(n3748), .Y(n6071) );
  AOI222X4 U495 ( .A0(net109791), .A1(n11398), .B0(mem_rdata_D[9]), .B1(n116), 
        .C0(n12988), .C1(net109801), .Y(n10772) );
  NAND2X6 U496 ( .A(n10882), .B(n10893), .Y(n10267) );
  NAND2X4 U497 ( .A(n10874), .B(n10873), .Y(n10882) );
  OA22X2 U498 ( .A0(n5337), .A1(n1188), .B0(n5293), .B1(n2760), .Y(n9443) );
  OR2X8 U499 ( .A(n7118), .B(n7117), .Y(n3805) );
  OA22X2 U500 ( .A0(\i_MIPS/n360 ), .A1(n4811), .B0(\i_MIPS/n359 ), .B1(n4805), 
        .Y(n6255) );
  INVX12 U501 ( .A(n4822), .Y(n4817) );
  CLKINVX2 U502 ( .A(net110257), .Y(n3610) );
  NAND4X4 U503 ( .A(n7400), .B(n7399), .C(n7398), .D(n7397), .Y(n11394) );
  OA22X2 U504 ( .A0(net112467), .A1(n932), .B0(net112343), .B1(n2456), .Y(
        n7321) );
  OAI221X2 U505 ( .A0(\i_MIPS/n362 ), .A1(n4825), .B0(\i_MIPS/n361 ), .B1(
        n4817), .C0(n6255), .Y(n8142) );
  INVX16 U506 ( .A(n4808), .Y(n4803) );
  OR2X4 U507 ( .A(\i_MIPS/n346 ), .B(n4803), .Y(n4197) );
  OAI221X2 U508 ( .A0(\i_MIPS/n363 ), .A1(n4810), .B0(\i_MIPS/n362 ), .B1(
        n4803), .C0(n6357), .Y(n8088) );
  OR2X2 U509 ( .A(net98430), .B(n10270), .Y(n76) );
  NAND2X4 U510 ( .A(n8249), .B(n4523), .Y(n8889) );
  NAND2X8 U511 ( .A(n6574), .B(\i_MIPS/n354 ), .Y(n7777) );
  CLKBUFX4 U512 ( .A(n5274), .Y(n5246) );
  INVX4 U513 ( .A(n10313), .Y(n62) );
  INVX4 U514 ( .A(n11069), .Y(n3628) );
  NOR3X6 U515 ( .A(n24), .B(n25), .C(n26), .Y(n7208) );
  AND2X8 U516 ( .A(n7189), .B(n7865), .Y(n25) );
  NAND2X2 U517 ( .A(n8822), .B(n5589), .Y(n7102) );
  OR2X2 U518 ( .A(n4548), .B(n8337), .Y(n4432) );
  OR2X6 U519 ( .A(n8337), .B(n8336), .Y(n4433) );
  OR2X8 U520 ( .A(n4089), .B(n4090), .Y(n4031) );
  NAND2X2 U521 ( .A(n9258), .B(n8338), .Y(n8337) );
  XOR3X2 U522 ( .A(net111409), .B(n10500), .C(n10384), .Y(n10391) );
  NAND2X8 U523 ( .A(n10292), .B(n155), .Y(n10950) );
  AOI211X2 U524 ( .A0(n4564), .A1(n10379), .B0(n10492), .C0(n10378), .Y(n10383) );
  NAND4X8 U525 ( .A(n6023), .B(n6022), .C(n6021), .D(n6020), .Y(n11370) );
  BUFX20 U526 ( .A(n3631), .Y(n5452) );
  NAND3BX4 U527 ( .AN(n10279), .B(n10278), .C(n11084), .Y(n10280) );
  INVX6 U528 ( .A(n10277), .Y(n11084) );
  NAND3BX2 U529 ( .AN(n10298), .B(n10276), .C(n10277), .Y(n10281) );
  NAND2X6 U530 ( .A(n4553), .B(n4801), .Y(n7850) );
  BUFX16 U531 ( .A(n8644), .Y(n4801) );
  OR2X2 U532 ( .A(n4526), .B(net110241), .Y(n3569) );
  NAND2X8 U533 ( .A(n6245), .B(\i_MIPS/ALUin1[11] ), .Y(n7107) );
  INVX8 U534 ( .A(n6246), .Y(n6245) );
  AND3X6 U535 ( .A(n3726), .B(n10255), .C(net99855), .Y(n3725) );
  OR2X2 U536 ( .A(n4561), .B(net110241), .Y(n4405) );
  NAND2X2 U537 ( .A(n12965), .B(DCACHE_addr[1]), .Y(n10152) );
  CLKINVX6 U538 ( .A(n12964), .Y(n4318) );
  INVX6 U539 ( .A(n10487), .Y(n11012) );
  NAND2BX4 U540 ( .AN(n5458), .B(n11236), .Y(n9837) );
  NAND4X6 U541 ( .A(n9973), .B(n9972), .C(n9971), .D(n9970), .Y(n11083) );
  NAND2BX4 U542 ( .AN(n5452), .B(n11337), .Y(n9973) );
  AOI21X4 U543 ( .A0(n10300), .A1(n10299), .B0(n10298), .Y(n4590) );
  INVX6 U544 ( .A(n10264), .Y(n10298) );
  OAI2BB2X2 U545 ( .B0(\i_MIPS/n168 ), .B1(net110219), .A0N(n175), .A1N(n11026), .Y(\i_MIPS/N109 ) );
  INVX3 U546 ( .A(n11027), .Y(n11026) );
  NAND2X8 U547 ( .A(n6243), .B(\i_MIPS/n363 ), .Y(n7179) );
  NAND2X8 U548 ( .A(n7179), .B(n7180), .Y(n6224) );
  OR2X4 U549 ( .A(n4537), .B(net110243), .Y(n4176) );
  OR2X4 U550 ( .A(n9336), .B(n9339), .Y(n3301) );
  NOR3X6 U551 ( .A(n9337), .B(n3301), .C(n9338), .Y(n9340) );
  AO22X4 U552 ( .A0(mem_rdata_I[73]), .A1(n115), .B0(n5469), .B1(n11303), .Y(
        n9635) );
  NAND2X4 U553 ( .A(n11118), .B(n155), .Y(n11015) );
  BUFX4 U554 ( .A(n5313), .Y(n5305) );
  BUFX8 U555 ( .A(n5290), .Y(n5313) );
  OAI2BB2X2 U556 ( .B0(\i_MIPS/n177 ), .B1(net110227), .A0N(n10708), .A1N(n176), .Y(\i_MIPS/N118 ) );
  BUFX20 U557 ( .A(net110259), .Y(net110255) );
  INVX8 U558 ( .A(n6930), .Y(n6639) );
  NAND2X8 U559 ( .A(n7096), .B(n7186), .Y(n6930) );
  CLKINVX2 U560 ( .A(n3696), .Y(n7707) );
  NAND3X8 U561 ( .A(ICACHE_addr[18]), .B(ICACHE_addr[17]), .C(n9362), .Y(
        n10291) );
  INVX8 U562 ( .A(n10289), .Y(n9362) );
  CLKINVX12 U563 ( .A(n10200), .Y(n10361) );
  NAND3X8 U564 ( .A(ICACHE_addr[22]), .B(ICACHE_addr[21]), .C(n10201), .Y(
        n10200) );
  INVX20 U565 ( .A(n4423), .Y(n4424) );
  OR2X8 U566 ( .A(n10697), .B(\i_MIPS/PC/n31 ), .Y(n10714) );
  OAI2BB1X1 U567 ( .A0N(net111405), .A1N(n10719), .B0(n10718), .Y(n10720) );
  OR2X4 U568 ( .A(n10336), .B(net110251), .Y(n4417) );
  NAND3X2 U569 ( .A(n4416), .B(n4415), .C(n4417), .Y(n10341) );
  OR2X1 U570 ( .A(net98501), .B(net110243), .Y(n3653) );
  NOR4X2 U571 ( .A(n7346), .B(n7345), .C(n7344), .D(n7343), .Y(n7347) );
  CLKBUFX3 U572 ( .A(n9308), .Y(n4975) );
  INVX4 U573 ( .A(n6514), .Y(n9308) );
  CLKINVX20 U574 ( .A(n5595), .Y(n5594) );
  INVX16 U575 ( .A(n4743), .Y(n8655) );
  OR2X1 U576 ( .A(n8075), .B(n7961), .Y(n7) );
  OR2X2 U577 ( .A(n8527), .B(n7), .Y(n4440) );
  NAND2X6 U578 ( .A(n4440), .B(n3724), .Y(n7981) );
  OR2X2 U579 ( .A(n6677), .B(n9171), .Y(n8) );
  OR2X2 U580 ( .A(n11224), .B(n6676), .Y(n9) );
  OR2X1 U581 ( .A(n9137), .B(n8439), .Y(n10) );
  NAND3X4 U582 ( .A(n8), .B(n9), .C(n10), .Y(n6678) );
  NAND2X2 U583 ( .A(n9258), .B(n6661), .Y(n6677) );
  NAND2X1 U584 ( .A(\i_MIPS/ALUin1[28] ), .B(n6617), .Y(n9171) );
  NAND2X4 U585 ( .A(n6617), .B(\i_MIPS/n343 ), .Y(n11224) );
  NAND2X8 U586 ( .A(n5589), .B(n9140), .Y(n9137) );
  OAI221X4 U587 ( .A0(\i_MIPS/ALUin1[22] ), .A1(n4825), .B0(
        \i_MIPS/ALUin1[23] ), .B1(n4817), .C0(n6675), .Y(n8439) );
  CLKAND2X8 U588 ( .A(n8067), .B(n7956), .Y(n11) );
  AND3X8 U589 ( .A(n4555), .B(n11), .C(n8520), .Y(n4523) );
  NAND2X4 U590 ( .A(n6582), .B(\i_MIPS/n349 ), .Y(n7956) );
  NAND2X8 U591 ( .A(n6580), .B(\i_MIPS/n351 ), .Y(n8520) );
  CLKAND2X12 U592 ( .A(n7025), .B(n7030), .Y(n4555) );
  NAND2X2 U593 ( .A(\i_MIPS/ID_EX[78] ), .B(n3769), .Y(n12) );
  INVX1 U594 ( .A(n6214), .Y(n13) );
  AND2X4 U595 ( .A(n12), .B(n13), .Y(n6207) );
  CLKINVX2 U596 ( .A(n3768), .Y(n3769) );
  NAND2X6 U597 ( .A(n3755), .B(n3800), .Y(n6214) );
  NOR3X2 U598 ( .A(n8976), .B(n8978), .C(n8977), .Y(n14) );
  NOR2X4 U599 ( .A(n8979), .B(n15), .Y(n8980) );
  INVX3 U600 ( .A(n14), .Y(n15) );
  AO22XL U601 ( .A0(n4974), .A1(n581), .B0(n4967), .B1(n2096), .Y(n8979) );
  NAND4BX4 U602 ( .AN(n8983), .B(n8982), .C(n8981), .D(n8980), .Y(n8994) );
  OR2X8 U603 ( .A(n9949), .B(n5452), .Y(n16) );
  OR2X6 U604 ( .A(n9948), .B(n5457), .Y(n17) );
  NAND3X8 U605 ( .A(n16), .B(n17), .C(n9947), .Y(net99146) );
  INVX6 U606 ( .A(n11341), .Y(n9949) );
  INVX3 U607 ( .A(n11245), .Y(n9948) );
  BUFX20 U608 ( .A(net99146), .Y(net113551) );
  NAND2X4 U609 ( .A(n11025), .B(net99146), .Y(n10952) );
  OR2X4 U610 ( .A(n7270), .B(n7544), .Y(n18) );
  OR2X1 U611 ( .A(n8659), .B(n7459), .Y(n19) );
  OR2X6 U612 ( .A(n8817), .B(n7269), .Y(n20) );
  NAND3X6 U613 ( .A(n18), .B(n19), .C(n20), .Y(n7293) );
  INVX1 U614 ( .A(n8083), .Y(n7270) );
  INVX6 U615 ( .A(n4470), .Y(n8659) );
  INVX8 U616 ( .A(n7293), .Y(n3701) );
  NOR3X2 U617 ( .A(n8985), .B(n8987), .C(n8986), .Y(n21) );
  NOR2X4 U618 ( .A(n8988), .B(n22), .Y(n8989) );
  INVX3 U619 ( .A(n21), .Y(n22) );
  AO22XL U620 ( .A0(n4974), .A1(n242), .B0(n4967), .B1(n2090), .Y(n8988) );
  NAND4BX4 U621 ( .AN(n8992), .B(n8991), .C(n8990), .D(n8989), .Y(n8993) );
  OR3X4 U622 ( .A(n3696), .B(n4800), .C(n7706), .Y(n23) );
  NAND2X4 U623 ( .A(n23), .B(n7705), .Y(n7717) );
  OA21X1 U624 ( .A0(n9259), .A1(n4800), .B0(n7714), .Y(n7705) );
  CLKAND2X2 U625 ( .A(n8263), .B(n8819), .Y(n24) );
  AND2X4 U626 ( .A(n7188), .B(n7866), .Y(n26) );
  CLKINVX8 U627 ( .A(n157), .Y(n7189) );
  CLKINVX8 U628 ( .A(n158), .Y(n7188) );
  OA21X4 U629 ( .A0(n9061), .A1(n9060), .B0(net102344), .Y(n27) );
  NAND2X6 U630 ( .A(n27), .B(net112607), .Y(net99970) );
  AO22X2 U631 ( .A0(net113455), .A1(n11448), .B0(net113463), .B1(n11417), .Y(
        n9061) );
  CLKINVX12 U632 ( .A(net100096), .Y(net102344) );
  OR3X8 U633 ( .A(n6626), .B(n6625), .C(n6624), .Y(n28) );
  NAND2X6 U634 ( .A(n28), .B(n7852), .Y(n3642) );
  INVX8 U635 ( .A(n8144), .Y(n6624) );
  NAND2X8 U636 ( .A(n161), .B(\i_MIPS/n353 ), .Y(n7852) );
  OR2X8 U637 ( .A(n3642), .B(n7858), .Y(n7957) );
  NOR3X4 U638 ( .A(n6034), .B(n30), .C(n6033), .Y(n6036) );
  INVX4 U639 ( .A(n29), .Y(n30) );
  NAND2X1 U640 ( .A(n4613), .B(n4695), .Y(n6034) );
  NAND2X2 U641 ( .A(n4616), .B(n9579), .Y(n6033) );
  OR2X1 U642 ( .A(\i_MIPS/n350 ), .B(n4824), .Y(n31) );
  OR2X1 U643 ( .A(\i_MIPS/n351 ), .B(n4817), .Y(n32) );
  OA21X1 U644 ( .A0(\i_MIPS/n352 ), .A1(n4812), .B0(n7871), .Y(n6953) );
  NOR3X2 U645 ( .A(n8692), .B(n8694), .C(n8693), .Y(n33) );
  NOR2X4 U646 ( .A(n8695), .B(n34), .Y(n8696) );
  INVX3 U647 ( .A(n33), .Y(n34) );
  AO22XL U648 ( .A0(n4974), .A1(n576), .B0(n4967), .B1(n2088), .Y(n8695) );
  AO22X1 U649 ( .A0(n4977), .A1(n541), .B0(n9309), .B1(n2296), .Y(n8694) );
  NAND4BX4 U650 ( .AN(n8699), .B(n8698), .C(n8697), .D(n8696), .Y(n8710) );
  OA21X4 U651 ( .A0(n6938), .A1(n6937), .B0(n6935), .Y(n35) );
  NAND2X6 U652 ( .A(n35), .B(n6936), .Y(n3664) );
  NAND2X6 U653 ( .A(n7095), .B(n1613), .Y(n6935) );
  OAI2BB1X4 U654 ( .A0N(n3664), .A1N(n7025), .B0(n7024), .Y(n7035) );
  NAND2X4 U655 ( .A(n4555), .B(n3664), .Y(n8156) );
  AND2X4 U656 ( .A(n6600), .B(n6599), .Y(n36) );
  CLKAND2X12 U657 ( .A(n4617), .B(n36), .Y(n6611) );
  INVX1 U658 ( .A(n6601), .Y(n6600) );
  CLKINVX6 U659 ( .A(n37), .Y(n38) );
  NOR2X8 U660 ( .A(n10493), .B(n10490), .Y(n39) );
  NOR3X8 U661 ( .A(n10332), .B(n40), .C(n10489), .Y(n10333) );
  INVX8 U662 ( .A(n39), .Y(n40) );
  NAND2X4 U663 ( .A(n4508), .B(n10331), .Y(n10493) );
  NAND2X8 U664 ( .A(n10952), .B(n10950), .Y(n10490) );
  INVX3 U665 ( .A(n10494), .Y(n10332) );
  NAND2X8 U666 ( .A(n10324), .B(n10323), .Y(n10489) );
  NAND2X8 U667 ( .A(n10487), .B(n10333), .Y(n10379) );
  NAND3X4 U668 ( .A(n6297), .B(n6300), .C(n6299), .Y(n41) );
  NAND2X8 U669 ( .A(n42), .B(n6298), .Y(net104563) );
  XOR2X1 U670 ( .A(n6291), .B(\i_MIPS/IR_ID[24] ), .Y(n6300) );
  CLKXOR2X1 U671 ( .A(n10129), .B(\i_MIPS/IR_ID[25] ), .Y(n6299) );
  OR2X6 U672 ( .A(net104831), .B(net104563), .Y(n3630) );
  OR2X6 U673 ( .A(net104525), .B(net104563), .Y(net139682) );
  NAND2X6 U674 ( .A(net104563), .B(n6301), .Y(n6303) );
  NAND2X8 U675 ( .A(net113075), .B(net104563), .Y(net102087) );
  OR2X2 U676 ( .A(net106108), .B(net112709), .Y(n43) );
  OR2X4 U677 ( .A(net106109), .B(net112723), .Y(n44) );
  MX2X1 U678 ( .A(n6926), .B(n6925), .S0(net108963), .Y(net106108) );
  CLKBUFX12 U679 ( .A(net112725), .Y(net112723) );
  AO21X2 U680 ( .A0(net99581), .A1(net99582), .B0(net112727), .Y(net106110) );
  AND2X2 U681 ( .A(\i_MIPS/ID_EX[103] ), .B(n5516), .Y(n45) );
  OR2XL U682 ( .A(n45), .B(n4499), .Y(\i_MIPS/n482 ) );
  AND2X4 U683 ( .A(\i_MIPS/Sign_Extend_ID[31] ), .B(n5511), .Y(n4499) );
  AND2XL U684 ( .A(n4800), .B(n8929), .Y(n46) );
  NOR3X2 U685 ( .A(n46), .B(n47), .C(n48), .Y(n8917) );
  BUFX20 U686 ( .A(n3723), .Y(n4800) );
  CLKINVX8 U687 ( .A(n8901), .Y(n8914) );
  NOR2X8 U688 ( .A(n3550), .B(n6628), .Y(n49) );
  NOR2X8 U689 ( .A(n3549), .B(n50), .Y(n3548) );
  INVX8 U690 ( .A(n49), .Y(n50) );
  NOR2X6 U691 ( .A(n8900), .B(n8899), .Y(n3549) );
  INVX16 U692 ( .A(n8897), .Y(n6628) );
  OR2X1 U693 ( .A(n4520), .B(n7851), .Y(n51) );
  OR2X8 U694 ( .A(n7850), .B(n7851), .Y(n52) );
  NAND3X6 U695 ( .A(n51), .B(n52), .C(n7849), .Y(n7855) );
  OA21X1 U696 ( .A0(n7848), .A1(n8151), .B0(n7847), .Y(n7849) );
  INVX8 U697 ( .A(n7855), .Y(n7854) );
  OR2X2 U698 ( .A(n6866), .B(n6867), .Y(n53) );
  OR2X8 U699 ( .A(n6865), .B(n6864), .Y(n54) );
  NAND3X6 U700 ( .A(n53), .B(n54), .C(n6863), .Y(net99062) );
  AND2XL U701 ( .A(n6850), .B(n3747), .Y(n6864) );
  INVX4 U702 ( .A(net99062), .Y(net106271) );
  OR2X1 U703 ( .A(n8525), .B(n4596), .Y(n56) );
  NAND3X6 U704 ( .A(n55), .B(n56), .C(n8524), .Y(n8554) );
  NAND2X2 U705 ( .A(n8249), .B(n4555), .Y(n8526) );
  INVX6 U706 ( .A(n8071), .Y(n8525) );
  CLKAND2X2 U707 ( .A(n7957), .B(n7853), .Y(n4596) );
  NAND3BX4 U708 ( .AN(n8528), .B(n4928), .C(n8554), .Y(n8559) );
  INVX4 U709 ( .A(n8554), .Y(n8555) );
  NOR3X2 U710 ( .A(n8495), .B(n8497), .C(n8496), .Y(n57) );
  NOR2X4 U711 ( .A(n8498), .B(n58), .Y(n8499) );
  INVX3 U712 ( .A(n57), .Y(n58) );
  AO22XL U713 ( .A0(n4973), .A1(n569), .B0(n4966), .B1(n2079), .Y(n8498) );
  AO22X1 U714 ( .A0(n5001), .A1(n548), .B0(n4997), .B1(n2303), .Y(n8495) );
  NAND4BX4 U715 ( .AN(n8502), .B(n8501), .C(n8500), .D(n8499), .Y(net103393)
         );
  NAND3X6 U716 ( .A(n6024), .B(n6025), .C(n6027), .Y(n59) );
  NAND2X8 U717 ( .A(n60), .B(n6026), .Y(n11369) );
  INVX8 U718 ( .A(n59), .Y(n60) );
  CLKINVX6 U719 ( .A(n10911), .Y(n10313) );
  NAND2X8 U720 ( .A(n3635), .B(n10315), .Y(n10487) );
  OR2X4 U721 ( .A(net104023), .B(net112709), .Y(n65) );
  OR2X8 U722 ( .A(net104024), .B(net112721), .Y(n66) );
  NAND3X8 U723 ( .A(n65), .B(n66), .C(net104025), .Y(net99424) );
  INVX20 U724 ( .A(net130301), .Y(net112709) );
  CLKINVX8 U725 ( .A(net99430), .Y(net104024) );
  BUFX16 U726 ( .A(net99424), .Y(n3732) );
  NOR3X2 U727 ( .A(n8504), .B(n8505), .C(n8506), .Y(n67) );
  NOR2X4 U728 ( .A(n8507), .B(n68), .Y(n8508) );
  INVX3 U729 ( .A(n67), .Y(n68) );
  AO22XL U730 ( .A0(n4973), .A1(n240), .B0(n4966), .B1(n2078), .Y(n8507) );
  AO22X1 U731 ( .A0(n4979), .A1(n497), .B0(n9309), .B1(n2249), .Y(n8506) );
  AO22X1 U732 ( .A0(n5001), .A1(n547), .B0(n4997), .B1(n2302), .Y(n8504) );
  NAND4BX4 U733 ( .AN(n8511), .B(n8510), .C(n8509), .D(n8508), .Y(net103394)
         );
  NAND3X6 U734 ( .A(n69), .B(n70), .C(n71), .Y(n72) );
  NAND2X8 U735 ( .A(n72), .B(n6241), .Y(n8896) );
  CLKINVX2 U736 ( .A(n3754), .Y(n69) );
  INVX3 U737 ( .A(n7453), .Y(n70) );
  INVX3 U738 ( .A(n3668), .Y(n71) );
  NAND2X2 U739 ( .A(n8712), .B(n7354), .Y(n7453) );
  AOI211X4 U740 ( .A0(n3665), .A1(n7452), .B0(n6240), .C0(n6455), .Y(n6241) );
  NAND2X2 U741 ( .A(n7463), .B(n8896), .Y(n6848) );
  CLKINVX12 U742 ( .A(n8896), .Y(n7095) );
  NAND2X4 U743 ( .A(n4606), .B(n8896), .Y(n6643) );
  NAND2X2 U744 ( .A(n4606), .B(n8896), .Y(n108) );
  NAND2X4 U745 ( .A(n8933), .B(n164), .Y(n73) );
  INVX3 U746 ( .A(n8935), .Y(n164) );
  OR2X4 U747 ( .A(n10271), .B(net140280), .Y(n75) );
  AND2X2 U748 ( .A(n75), .B(n76), .Y(n10259) );
  INVX6 U749 ( .A(n10273), .Y(n10271) );
  NAND2X2 U750 ( .A(n9955), .B(n9956), .Y(n77) );
  NAND3X6 U751 ( .A(n9957), .B(n9958), .C(n78), .Y(n11305) );
  INVX3 U752 ( .A(n77), .Y(n78) );
  AO22X4 U753 ( .A0(mem_rdata_I[75]), .A1(n113), .B0(n5468), .B1(n11305), .Y(
        n9959) );
  NAND2BX2 U754 ( .AN(n5454), .B(n11305), .Y(n9972) );
  INVX3 U755 ( .A(n79), .Y(n80) );
  INVX12 U756 ( .A(n3731), .Y(net99849) );
  OR2X6 U757 ( .A(net105577), .B(net112709), .Y(n81) );
  OR2X8 U758 ( .A(net105578), .B(net112723), .Y(n82) );
  NAND3X8 U759 ( .A(n81), .B(n82), .C(net105579), .Y(net99330) );
  MX2X1 U760 ( .A(n7268), .B(n7267), .S0(net108963), .Y(net105577) );
  CLKINVX8 U761 ( .A(net99336), .Y(net105578) );
  NAND3X4 U762 ( .A(n83), .B(n84), .C(n85), .Y(n86) );
  NAND2X6 U763 ( .A(n86), .B(n4596), .Y(n7779) );
  INVX2 U764 ( .A(n8527), .Y(n83) );
  INVX3 U765 ( .A(n7778), .Y(n85) );
  NAND2X4 U766 ( .A(n7779), .B(n7802), .Y(n7806) );
  INVX4 U767 ( .A(n7779), .Y(n7780) );
  NAND2X6 U768 ( .A(net102413), .B(net137470), .Y(n87) );
  NAND2X8 U769 ( .A(n88), .B(net137471), .Y(net99654) );
  INVX12 U770 ( .A(n87), .Y(n88) );
  OR2X4 U771 ( .A(n9082), .B(net112707), .Y(net137470) );
  NAND2X8 U772 ( .A(n3528), .B(n3621), .Y(net137471) );
  OR2XL U773 ( .A(n4517), .B(n8537), .Y(n89) );
  OR2X1 U774 ( .A(n9128), .B(n141), .Y(n90) );
  OR2XL U775 ( .A(n8273), .B(n8805), .Y(n91) );
  INVX12 U776 ( .A(n139), .Y(n141) );
  INVX16 U777 ( .A(n3723), .Y(n8805) );
  NOR4X6 U778 ( .A(n8279), .B(n8276), .C(n8277), .D(n8278), .Y(n8285) );
  OR2X1 U779 ( .A(net112655), .B(n1884), .Y(n92) );
  OR2X2 U780 ( .A(net112587), .B(n253), .Y(n93) );
  NAND3X6 U781 ( .A(n92), .B(n93), .C(n6064), .Y(n6065) );
  BUFX20 U782 ( .A(net112695), .Y(net112655) );
  INVX8 U783 ( .A(n6065), .Y(n10621) );
  OR2X6 U784 ( .A(net104351), .B(net112709), .Y(n94) );
  OR2X8 U785 ( .A(net104352), .B(net112721), .Y(n95) );
  NAND3X8 U786 ( .A(n94), .B(n95), .C(net104353), .Y(n3856) );
  CLKINVX8 U787 ( .A(net99290), .Y(net104352) );
  CLKBUFX20 U788 ( .A(net112725), .Y(net112721) );
  NOR2X8 U789 ( .A(net99849), .B(net99664), .Y(n96) );
  INVX6 U790 ( .A(net99932), .Y(n97) );
  NOR2X8 U791 ( .A(n96), .B(n97), .Y(n3795) );
  NAND2X8 U792 ( .A(\i_MIPS/IF_ID[64] ), .B(\i_MIPS/IF_ID[97] ), .Y(net99664)
         );
  OR2X4 U793 ( .A(n8527), .B(n8889), .Y(n98) );
  OR2X2 U794 ( .A(n8251), .B(n3767), .Y(n99) );
  NAND3X6 U795 ( .A(n98), .B(n99), .C(n8250), .Y(n8256) );
  CLKINVX1 U796 ( .A(n7956), .Y(n8251) );
  CLKINVX6 U797 ( .A(n8256), .Y(n8257) );
  NAND3BX4 U798 ( .AN(n8273), .B(n4927), .C(n8256), .Y(n8287) );
  NAND2X2 U799 ( .A(\i_MIPS/ID_EX[68] ), .B(n100), .Y(n101) );
  NAND2X4 U800 ( .A(n101), .B(n102), .Y(n103) );
  CLKINVX20 U801 ( .A(n5595), .Y(n3826) );
  INVX6 U802 ( .A(n6565), .Y(n6615) );
  NAND2XL U803 ( .A(n8327), .B(n8328), .Y(n104) );
  NAND2X4 U804 ( .A(n105), .B(n4801), .Y(n8923) );
  INVX3 U805 ( .A(n104), .Y(n105) );
  CLKINVX12 U806 ( .A(n8515), .Y(n8327) );
  NAND2X6 U807 ( .A(n3206), .B(n9155), .Y(n106) );
  NAND2X8 U808 ( .A(n107), .B(n4743), .Y(n9158) );
  CLKINVX8 U809 ( .A(n106), .Y(n107) );
  BUFX16 U810 ( .A(n9154), .Y(n4743) );
  CLKINVX4 U811 ( .A(n9153), .Y(n9155) );
  AND2X4 U812 ( .A(n9156), .B(n9157), .Y(n3206) );
  INVX1 U813 ( .A(n8895), .Y(n109) );
  NAND2X2 U814 ( .A(n108), .B(n109), .Y(n8899) );
  OR2X6 U815 ( .A(n9295), .B(n9296), .Y(n110) );
  OR2X6 U816 ( .A(n9293), .B(n9294), .Y(n111) );
  NAND3X6 U817 ( .A(n110), .B(n111), .C(n9292), .Y(n10637) );
  NOR3X4 U818 ( .A(n3572), .B(n3573), .C(n4800), .Y(n9295) );
  AND2X1 U819 ( .A(n9257), .B(n9256), .Y(n9296) );
  AND4X6 U820 ( .A(n9291), .B(n9290), .C(n9289), .D(n9288), .Y(n9292) );
  BUFX16 U821 ( .A(n10637), .Y(n4727) );
  INVX4 U822 ( .A(n8930), .Y(n8928) );
  OR2X2 U823 ( .A(n10732), .B(n10719), .Y(n3570) );
  INVX6 U824 ( .A(n10153), .Y(n10147) );
  NAND2X2 U825 ( .A(DCACHE_addr[1]), .B(n4047), .Y(n10153) );
  OR2X4 U826 ( .A(net112651), .B(n2416), .Y(n3715) );
  BUFX20 U827 ( .A(net112697), .Y(net112651) );
  NOR3BX4 U828 ( .AN(n10717), .B(n10712), .C(n10702), .Y(n10706) );
  AOI2BB2X2 U829 ( .B0(\i_MIPS/IF_ID[65] ), .B1(n11186), .A0N(n11186), .A1N(
        \i_MIPS/n180 ), .Y(n10814) );
  OAI22X1 U830 ( .A0(net110241), .A1(net98901), .B0(net110213), .B1(
        \i_MIPS/PC/n3 ), .Y(n10834) );
  OA22X4 U831 ( .A0(n10970), .A1(net140281), .B0(net98430), .B1(n10969), .Y(
        n10972) );
  CLKXOR2X4 U832 ( .A(n10320), .B(ICACHE_addr[21]), .Y(n10969) );
  AOI2BB1X2 U833 ( .A0N(n10272), .A1N(n10308), .B0(n10909), .Y(n10275) );
  CLKINVX4 U834 ( .A(n10909), .Y(n10916) );
  AND4X6 U835 ( .A(n10730), .B(n10729), .C(n10728), .D(n10727), .Y(n4444) );
  NAND4X1 U836 ( .A(n10726), .B(n10722), .C(n10717), .D(n10723), .Y(n10730) );
  NAND2X2 U837 ( .A(net111405), .B(n10698), .Y(n10718) );
  INVX3 U838 ( .A(n11162), .Y(n112) );
  INVX12 U839 ( .A(n112), .Y(n113) );
  INVX12 U840 ( .A(n112), .Y(n114) );
  INVX12 U841 ( .A(n112), .Y(n115) );
  AOI21XL U842 ( .A0(n9572), .A1(n9344), .B0(n11358), .Y(n11162) );
  NAND2X8 U843 ( .A(n3795), .B(net99933), .Y(n10386) );
  OR2X8 U844 ( .A(n10942), .B(net110251), .Y(n4214) );
  BUFX20 U845 ( .A(net98391), .Y(n116) );
  BUFX20 U846 ( .A(net98391), .Y(n117) );
  AND2X4 U847 ( .A(n10138), .B(mem_ready_D), .Y(net98391) );
  MX2X1 U848 ( .A(\D_cache/cache[4][140] ), .B(n10622), .S0(net112197), .Y(
        \D_cache/n672 ) );
  MX2X1 U849 ( .A(\D_cache/cache[6][140] ), .B(n10622), .S0(net111995), .Y(
        \D_cache/n670 ) );
  MX2X1 U850 ( .A(\D_cache/cache[1][140] ), .B(n10622), .S0(net112533), .Y(
        \D_cache/n675 ) );
  MX2X1 U851 ( .A(\D_cache/cache[0][140] ), .B(n10622), .S0(net112635), .Y(
        \D_cache/n676 ) );
  MX2X1 U852 ( .A(\D_cache/cache[3][140] ), .B(n10622), .S0(net112285), .Y(
        \D_cache/n673 ) );
  MX2X1 U853 ( .A(\D_cache/cache[2][140] ), .B(n10622), .S0(net112409), .Y(
        \D_cache/n674 ) );
  AO22X4 U854 ( .A0(n5062), .A1(n12951), .B0(n5060), .B1(n11529), .Y(n10622)
         );
  MX2X1 U855 ( .A(\D_cache/cache[3][146] ), .B(n10669), .S0(net112277), .Y(
        \D_cache/n625 ) );
  MX2X1 U856 ( .A(\D_cache/cache[1][146] ), .B(n10669), .S0(net112535), .Y(
        \D_cache/n627 ) );
  MX2X1 U857 ( .A(\D_cache/cache[0][146] ), .B(n10669), .S0(net112637), .Y(
        \D_cache/n628 ) );
  MX2X1 U858 ( .A(\D_cache/cache[2][146] ), .B(n10669), .S0(net112411), .Y(
        \D_cache/n626 ) );
  MX2X1 U859 ( .A(\D_cache/cache[4][146] ), .B(n10669), .S0(net112211), .Y(
        \D_cache/n624 ) );
  MX2X1 U860 ( .A(\D_cache/cache[7][146] ), .B(n10669), .S0(net111881), .Y(
        \D_cache/n621 ) );
  AO22X4 U861 ( .A0(n5063), .A1(n12945), .B0(n5061), .B1(n11535), .Y(n10669)
         );
  BUFX12 U862 ( .A(n10633), .Y(n118) );
  AO22X1 U863 ( .A0(n5062), .A1(DCACHE_addr[5]), .B0(n5060), .B1(n11518), .Y(
        n10633) );
  BUFX8 U864 ( .A(n10662), .Y(n119) );
  AO22X1 U865 ( .A0(n5063), .A1(n12941), .B0(n5061), .B1(n11539), .Y(n10662)
         );
  BUFX8 U866 ( .A(n10646), .Y(n120) );
  AO22X1 U867 ( .A0(n5062), .A1(n12942), .B0(n5060), .B1(n11538), .Y(n10646)
         );
  BUFX12 U868 ( .A(n10659), .Y(n121) );
  AO22X1 U869 ( .A0(n5063), .A1(n12946), .B0(n5061), .B1(n11534), .Y(n10659)
         );
  BUFX8 U870 ( .A(n10643), .Y(n122) );
  AO22X1 U871 ( .A0(n5062), .A1(n12944), .B0(n5060), .B1(n11536), .Y(n10643)
         );
  BUFX8 U872 ( .A(n10665), .Y(n123) );
  AO22X1 U873 ( .A0(n5063), .A1(n12958), .B0(n5061), .B1(n11523), .Y(n10665)
         );
  BUFX8 U874 ( .A(n10628), .Y(n124) );
  AO22X1 U875 ( .A0(n5062), .A1(DCACHE_addr[16]), .B0(n5060), .B1(n3832), .Y(
        n10628) );
  BUFX8 U876 ( .A(n10674), .Y(n125) );
  AO22X1 U877 ( .A0(n5063), .A1(DCACHE_addr[18]), .B0(n5061), .B1(n11530), .Y(
        n10674) );
  BUFX8 U878 ( .A(n10631), .Y(n126) );
  AO22X1 U879 ( .A0(n5062), .A1(DCACHE_addr[29]), .B0(n5060), .B1(n11541), .Y(
        n10631) );
  OAI22X2 U880 ( .A0(n10703), .A1(n10717), .B0(n10701), .B1(n10700), .Y(n10707) );
  BUFX8 U881 ( .A(n10663), .Y(n127) );
  AO22X1 U882 ( .A0(n5063), .A1(DCACHE_addr[11]), .B0(n5061), .B1(n11524), .Y(
        n10663) );
  BUFX8 U883 ( .A(n10625), .Y(n128) );
  AO22X1 U884 ( .A0(n5062), .A1(DCACHE_addr[21]), .B0(n5060), .B1(n11533), .Y(
        n10625) );
  BUFX8 U885 ( .A(n10667), .Y(n129) );
  AO22X1 U886 ( .A0(n5063), .A1(n12953), .B0(n5061), .B1(n11528), .Y(n10667)
         );
  BUFX8 U887 ( .A(n10649), .Y(n130) );
  AO22X1 U888 ( .A0(n5062), .A1(DCACHE_addr[12]), .B0(n5060), .B1(n11525), .Y(
        n10649) );
  BUFX8 U889 ( .A(n10676), .Y(n131) );
  AO22X1 U890 ( .A0(n5063), .A1(DCACHE_addr[7]), .B0(n5061), .B1(n11520), .Y(
        n10676) );
  BUFX8 U891 ( .A(n10640), .Y(n132) );
  AO22X1 U892 ( .A0(n5062), .A1(DCACHE_addr[28]), .B0(n5060), .B1(n11540), .Y(
        n10640) );
  CLKINVX8 U893 ( .A(n10677), .Y(n133) );
  INVX12 U894 ( .A(n133), .Y(n134) );
  BUFX4 U895 ( .A(n4626), .Y(n135) );
  BUFX8 U896 ( .A(n10652), .Y(n136) );
  AO22X1 U897 ( .A0(n5062), .A1(DCACHE_addr[14]), .B0(n5060), .B1(n11527), .Y(
        n10652) );
  BUFX8 U898 ( .A(n10680), .Y(n137) );
  AO22X1 U899 ( .A0(n5063), .A1(DCACHE_addr[6]), .B0(n5061), .B1(n11519), .Y(
        n10680) );
  XOR3X1 U900 ( .A(n10885), .B(n156), .C(n10884), .Y(n10887) );
  BUFX6 U901 ( .A(n4510), .Y(n156) );
  NAND2X6 U902 ( .A(net99850), .B(n4145), .Y(net99855) );
  CLKBUFX16 U903 ( .A(n12836), .Y(mem_addr_I[10]) );
  INVX3 U904 ( .A(n3885), .Y(n12836) );
  INVX16 U905 ( .A(n8536), .Y(n139) );
  INVX12 U906 ( .A(n139), .Y(n140) );
  BUFX8 U907 ( .A(n10636), .Y(n142) );
  AO22X1 U908 ( .A0(n5062), .A1(DCACHE_addr[13]), .B0(n5060), .B1(n11526), .Y(
        n10636) );
  BUFX8 U909 ( .A(n10672), .Y(n143) );
  AO22X1 U910 ( .A0(n5063), .A1(DCACHE_addr[20]), .B0(n5061), .B1(n11532), .Y(
        n10672) );
  NAND2X8 U911 ( .A(net114031), .B(n10387), .Y(n10255) );
  BUFX16 U912 ( .A(net98880), .Y(net114031) );
  BUFX8 U913 ( .A(n10654), .Y(n144) );
  AO22X1 U914 ( .A0(n5062), .A1(DCACHE_addr[25]), .B0(n5060), .B1(n11537), .Y(
        n10654) );
  BUFX8 U915 ( .A(n10657), .Y(n145) );
  AO22X1 U916 ( .A0(n5063), .A1(DCACHE_addr[9]), .B0(n5061), .B1(n11522), .Y(
        n10657) );
  CLKINVX1 U917 ( .A(n10719), .Y(n10713) );
  BUFX8 U918 ( .A(net99080), .Y(n181) );
  OA22X2 U919 ( .A0(net112245), .A1(n1371), .B0(net112163), .B1(n2984), .Y(
        n7236) );
  CLKBUFX12 U920 ( .A(net112165), .Y(net112163) );
  NAND4BX2 U921 ( .AN(n10834), .B(n10833), .C(n10832), .D(n10831), .Y(
        \i_MIPS/PC/n35 ) );
  CLKINVX12 U922 ( .A(n4327), .Y(mem_addr_I[14]) );
  NOR2X2 U923 ( .A(n4330), .B(n4331), .Y(n4327) );
  CLKINVX12 U924 ( .A(net130509), .Y(n146) );
  INVX16 U925 ( .A(n146), .Y(n147) );
  INVX16 U926 ( .A(n146), .Y(n148) );
  INVX12 U927 ( .A(n146), .Y(n149) );
  INVX12 U928 ( .A(n146), .Y(n150) );
  CLKAND2X12 U929 ( .A(n11188), .B(n11186), .Y(net130509) );
  NAND3X6 U930 ( .A(n3615), .B(n3616), .C(net107043), .Y(net98988) );
  AO21X2 U931 ( .A0(net98992), .A1(net98993), .B0(net112727), .Y(net107043) );
  OAI222X2 U932 ( .A0(\i_MIPS/PC/n24 ), .A1(net110215), .B0(n4528), .B1(
        net110241), .C0(n10957), .C1(net110247), .Y(n10963) );
  INVX8 U933 ( .A(n8523), .Y(n8522) );
  AND3X8 U934 ( .A(n3539), .B(n3540), .C(net104526), .Y(n3316) );
  NAND3X4 U935 ( .A(net139681), .B(net139682), .C(net104564), .Y(net99991) );
  NAND2X6 U936 ( .A(n6585), .B(\i_MIPS/n349 ), .Y(n7971) );
  MXI2X6 U937 ( .A(n4498), .B(\i_MIPS/ID_EX[95] ), .S0(n3771), .Y(n6585) );
  CLKAND2X2 U938 ( .A(n9258), .B(n9263), .Y(n3573) );
  INVX6 U939 ( .A(n4411), .Y(n8645) );
  NAND2BX4 U940 ( .AN(n8253), .B(n4412), .Y(n4411) );
  INVX20 U941 ( .A(net102087), .Y(net102300) );
  CLKBUFX4 U942 ( .A(net102300), .Y(net113167) );
  AOI22X4 U943 ( .A0(net113041), .A1(net99336), .B0(net113169), .B1(net105666), 
        .Y(n3315) );
  AOI2BB1X2 U944 ( .A0N(n4618), .A1N(n156), .B0(n10894), .Y(n10896) );
  MXI2X6 U945 ( .A(n3633), .B(\i_MIPS/ID_EX[84] ), .S0(n5594), .Y(n6246) );
  INVXL U946 ( .A(n8512), .Y(n8529) );
  NAND2X6 U947 ( .A(n8512), .B(n8080), .Y(n7954) );
  AO22X4 U948 ( .A0(net113457), .A1(n11446), .B0(net113463), .B1(n11415), .Y(
        n8402) );
  BUFX20 U949 ( .A(net100093), .Y(net112609) );
  AND3X8 U950 ( .A(n8257), .B(n8258), .C(n4926), .Y(n8279) );
  BUFX6 U951 ( .A(net100099), .Y(n182) );
  AO22X2 U952 ( .A0(net113455), .A1(n11423), .B0(net113461), .B1(n11392), .Y(
        n8864) );
  NAND2X6 U953 ( .A(net99363), .B(net99364), .Y(n4122) );
  AO21X4 U954 ( .A0(net99969), .A1(net99970), .B0(net112731), .Y(net102413) );
  BUFX4 U955 ( .A(n10887), .Y(n151) );
  CLKINVX6 U956 ( .A(n10957), .Y(n10956) );
  NAND3X2 U957 ( .A(n4213), .B(n4212), .C(n4214), .Y(n10947) );
  OAI2BB2X2 U958 ( .B0(\i_MIPS/n165 ), .B1(net110221), .A0N(n175), .A1N(n3846), 
        .Y(\i_MIPS/N106 ) );
  AND3XL U959 ( .A(n9554), .B(n4685), .C(n4651), .Y(n9334) );
  AOI211X2 U960 ( .A0(n167), .A1(\i_MIPS/n356 ), .B0(n6612), .C0(n6947), .Y(
        n6572) );
  MX2X8 U961 ( .A(\i_MIPS/n281 ), .B(n4713), .S0(n5594), .Y(n6612) );
  NAND4X6 U962 ( .A(n5960), .B(n5959), .C(n5958), .D(n5957), .Y(n11388) );
  CLKINVX12 U963 ( .A(n9567), .Y(n9554) );
  OAI222X2 U964 ( .A0(n6766), .A1(n158), .B0(n6765), .B1(n157), .C0(n8726), 
        .C1(n8910), .Y(n6784) );
  NOR4X8 U965 ( .A(n7115), .B(n7114), .C(n7113), .D(n7112), .Y(n7116) );
  AO22X4 U966 ( .A0(n7189), .A1(n7103), .B0(n7188), .B1(n7783), .Y(n7115) );
  OA22X2 U967 ( .A0(n10960), .A1(net140281), .B0(net98430), .B1(n10959), .Y(
        n10962) );
  OAI221X1 U968 ( .A0(\i_MIPS/ALUin1[18] ), .A1(n4810), .B0(
        \i_MIPS/ALUin1[19] ), .B1(n4803), .C0(n7792), .Y(n8272) );
  AOI2BB1X4 U969 ( .A0N(\i_MIPS/ALUin1[16] ), .A1N(n4826), .B0(n4612), .Y(
        n7792) );
  CLKINVX12 U970 ( .A(n9574), .Y(n9556) );
  NOR4X4 U971 ( .A(n9576), .B(n9575), .C(n9574), .D(n9573), .Y(n9588) );
  NOR4X8 U972 ( .A(n4072), .B(n4074), .C(n4075), .D(n4073), .Y(n4071) );
  XOR2X4 U973 ( .A(n11373), .B(ICACHE_addr[14]), .Y(n9568) );
  AOI2BB2X4 U974 ( .B0(n4681), .B1(\I_cache/cache[4][144] ), .A0N(n5286), 
        .A1N(n3214), .Y(n5955) );
  INVX4 U975 ( .A(net112609), .Y(net113919) );
  NOR2X2 U976 ( .A(n11001), .B(net110247), .Y(n4431) );
  AOI2BB2X2 U977 ( .B0(\i_MIPS/IF_ID[93] ), .B1(n150), .A0N(n10391), .A1N(
        net110251), .Y(n10392) );
  AOI2BB2X1 U978 ( .B0(\i_MIPS/IF_ID[68] ), .B1(n150), .A0N(net110191), .A1N(
        \i_MIPS/n183 ), .Y(n11004) );
  AOI2BB2X1 U979 ( .B0(\i_MIPS/IF_ID[82] ), .B1(n148), .A0N(net110189), .A1N(
        \i_MIPS/n197 ), .Y(n11114) );
  AOI2BB2X1 U980 ( .B0(\i_MIPS/IF_ID[72] ), .B1(n150), .A0N(net110189), .A1N(
        \i_MIPS/n187 ), .Y(n10867) );
  AOI2BB2X1 U981 ( .B0(\i_MIPS/IF_ID[78] ), .B1(n149), .A0N(net110191), .A1N(
        \i_MIPS/n193 ), .Y(n11090) );
  AOI2BB2X1 U982 ( .B0(\i_MIPS/IF_ID[80] ), .B1(n147), .A0N(net110189), .A1N(
        \i_MIPS/n195 ), .Y(n11100) );
  AOI2BB2X1 U983 ( .B0(\i_MIPS/IF_ID[91] ), .B1(n149), .A0N(net110189), .A1N(
        \i_MIPS/n206 ), .Y(n10358) );
  AOI2BB2X1 U984 ( .B0(\i_MIPS/IF_ID[89] ), .B1(n148), .A0N(net110189), .A1N(
        \i_MIPS/n204 ), .Y(n4138) );
  AOI2BB2X1 U985 ( .B0(\i_MIPS/IF_ID[85] ), .B1(n148), .A0N(net110191), .A1N(
        \i_MIPS/n200 ), .Y(n11021) );
  INVX4 U986 ( .A(n6213), .Y(n6218) );
  CLKINVX4 U987 ( .A(n6214), .Y(n6217) );
  CLKINVX12 U988 ( .A(n9573), .Y(n9557) );
  NAND3BX4 U989 ( .AN(n9571), .B(n4024), .C(n4018), .Y(n9576) );
  BUFX6 U990 ( .A(n11219), .Y(n154) );
  NAND2XL U991 ( .A(n11360), .B(n11515), .Y(n11219) );
  OAI221X4 U992 ( .A0(n9949), .A1(n5452), .B0(n9948), .B1(n5457), .C0(n9947), 
        .Y(n155) );
  CLKINVX12 U993 ( .A(net111405), .Y(n168) );
  INVX20 U994 ( .A(net113551), .Y(net98564) );
  OAI222X2 U995 ( .A0(n3650), .A1(net110215), .B0(n4540), .B1(net110243), .C0(
        n10899), .C1(net110249), .Y(n10904) );
  NAND3X2 U996 ( .A(n3569), .B(n3570), .C(n3571), .Y(n10711) );
  NAND2X2 U997 ( .A(net99850), .B(\i_MIPS/n233 ), .Y(net99845) );
  AOI32X2 U998 ( .A0(n10310), .A1(n10305), .A2(n10304), .B0(n10310), .B1(
        n10303), .Y(n10316) );
  OR2X2 U999 ( .A(net110251), .B(n10247), .Y(n4406) );
  NAND3BX2 U1000 ( .AN(n10726), .B(n10725), .C(n10724), .Y(n10727) );
  CLKINVX1 U1001 ( .A(n10712), .Y(n10726) );
  AOI2BB2X2 U1002 ( .B0(\i_MIPS/IF_ID[77] ), .B1(n147), .A0N(net110189), .A1N(
        \i_MIPS/n192 ), .Y(n10258) );
  NAND3BX2 U1003 ( .AN(n3693), .B(n3637), .C(n9620), .Y(n9453) );
  AOI2BB2X2 U1004 ( .B0(\i_MIPS/IF_ID[87] ), .B1(n150), .A0N(net110191), .A1N(
        \i_MIPS/n202 ), .Y(n10961) );
  NAND2X2 U1005 ( .A(n10381), .B(net113551), .Y(n10488) );
  INVX6 U1006 ( .A(n10380), .Y(n10381) );
  INVX6 U1007 ( .A(n10377), .Y(n10492) );
  NAND2X2 U1008 ( .A(n10364), .B(n155), .Y(n10377) );
  NAND3BX2 U1009 ( .AN(n10374), .B(n10373), .C(n10372), .Y(\i_MIPS/PC/n61 ) );
  NAND3BX2 U1010 ( .AN(n11033), .B(n11032), .C(n11031), .Y(\i_MIPS/PC/n55 ) );
  NAND2X6 U1011 ( .A(n4426), .B(n4427), .Y(n6567) );
  NAND2X2 U1012 ( .A(\i_MIPS/n273 ), .B(n4199), .Y(n4426) );
  NAND4X6 U1013 ( .A(n4461), .B(n4462), .C(n5955), .D(n5954), .Y(n11380) );
  NAND3X4 U1014 ( .A(n10246), .B(n10255), .C(net99855), .Y(net98436) );
  NAND3BX2 U1015 ( .AN(n10711), .B(n10710), .C(n10709), .Y(n11542) );
  NAND4X6 U1016 ( .A(n4453), .B(n4454), .C(n5950), .D(n5949), .Y(n11376) );
  AOI2BB2X4 U1017 ( .B0(n4681), .B1(\I_cache/cache[4][140] ), .A0N(n5286), 
        .A1N(n3208), .Y(n5950) );
  NAND4X6 U1018 ( .A(n4465), .B(n4466), .C(n5986), .D(n5985), .Y(n11377) );
  XOR2X4 U1019 ( .A(n11387), .B(ICACHE_addr[28]), .Y(n9567) );
  NAND4X8 U1020 ( .A(n4468), .B(n4469), .C(n5966), .D(n5965), .Y(n11387) );
  NAND3BX4 U1021 ( .AN(n10260), .B(n10259), .C(n10258), .Y(\i_MIPS/PC/n46 ) );
  OA22X4 U1022 ( .A0(net112465), .A1(n1370), .B0(net112341), .B1(n2983), .Y(
        n7237) );
  CLKBUFX4 U1023 ( .A(net112503), .Y(net112465) );
  OA22X4 U1024 ( .A0(n5248), .A1(n1977), .B0(n5203), .B1(n410), .Y(n6001) );
  BUFX16 U1025 ( .A(n5274), .Y(n5248) );
  XOR2X2 U1026 ( .A(n9453), .B(ICACHE_addr[5]), .Y(n10871) );
  INVX2 U1027 ( .A(n9453), .Y(n9451) );
  NAND2BX4 U1028 ( .AN(n5452), .B(n11336), .Y(n9677) );
  OA22X4 U1029 ( .A0(n5428), .A1(n3221), .B0(n5384), .B1(n359), .Y(n6003) );
  BUFX8 U1030 ( .A(n5408), .Y(n5384) );
  OR2X4 U1031 ( .A(net112139), .B(n1991), .Y(n3799) );
  OAI2BB2X1 U1032 ( .B0(\i_MIPS/n244 ), .B1(net110221), .A0N(n176), .A1N(
        n10898), .Y(\i_MIPS/N98 ) );
  CLKINVX2 U1033 ( .A(n10899), .Y(n10898) );
  OAI2BB2X4 U1034 ( .B0(net112019), .B1(n1862), .A0N(net111873), .A1N(
        \D_cache/cache[7][128] ), .Y(n3829) );
  NAND4X2 U1035 ( .A(n7822), .B(n7821), .C(n7820), .D(n7819), .Y(n11501) );
  OA22XL U1036 ( .A0(net112465), .A1(n956), .B0(net112351), .B1(n2481), .Y(
        n7821) );
  NAND2X8 U1037 ( .A(n7950), .B(n4515), .Y(n8253) );
  INVX4 U1038 ( .A(n7952), .Y(n7950) );
  INVX6 U1039 ( .A(n10888), .Y(n10885) );
  CLKAND2X12 U1040 ( .A(n10889), .B(n10888), .Y(n4618) );
  CLKXOR2X2 U1041 ( .A(n9431), .B(n3645), .Y(n10888) );
  INVX4 U1042 ( .A(n9281), .Y(n9282) );
  OAI221X4 U1043 ( .A0(\i_MIPS/ALUin1[23] ), .A1(n4824), .B0(
        \i_MIPS/ALUin1[24] ), .B1(n4816), .C0(n8347), .Y(n9281) );
  INVX8 U1044 ( .A(n11481), .Y(n10686) );
  NAND4X4 U1045 ( .A(n9244), .B(n9243), .C(n9242), .D(n9241), .Y(n11481) );
  NAND4X4 U1046 ( .A(n7238), .B(n7237), .C(n7236), .D(n7235), .Y(n11399) );
  CLKINVX8 U1047 ( .A(n8898), .Y(n6630) );
  NOR2X6 U1048 ( .A(n3767), .B(n8898), .Y(n3550) );
  NAND2X4 U1049 ( .A(n7956), .B(n8891), .Y(n8898) );
  NAND3X8 U1050 ( .A(n3804), .B(n3805), .C(n7116), .Y(net99039) );
  NAND2X2 U1051 ( .A(\i_MIPS/ALUin1[20] ), .B(n6580), .Y(n8512) );
  INVX3 U1052 ( .A(n6578), .Y(n6580) );
  OAI21X1 U1053 ( .A0(n10936), .A1(n10935), .B0(n10934), .Y(n10938) );
  NAND2X4 U1054 ( .A(net98564), .B(n11113), .Y(n10934) );
  NAND2X4 U1055 ( .A(\i_MIPS/ALUin1[26] ), .B(n6587), .Y(n8334) );
  AND2X8 U1056 ( .A(n7187), .B(n7100), .Y(n1224) );
  INVX8 U1057 ( .A(n6432), .Y(n6423) );
  CLKMX2X8 U1058 ( .A(\i_MIPS/n309 ), .B(n3800), .S0(n3826), .Y(n6432) );
  CLKAND2X12 U1059 ( .A(n7029), .B(n7709), .Y(n4553) );
  NAND2X4 U1060 ( .A(n167), .B(\i_MIPS/n356 ), .Y(n7709) );
  NAND2X6 U1061 ( .A(n3202), .B(n10666), .Y(n6152) );
  INVX8 U1062 ( .A(n6151), .Y(n10666) );
  AND3X8 U1063 ( .A(n4181), .B(n4182), .C(n6149), .Y(n3202) );
  CLKMX2X6 U1064 ( .A(\i_MIPS/n259 ), .B(n4650), .S0(n3826), .Y(n6586) );
  CLKMX2X6 U1065 ( .A(\i_MIPS/n321 ), .B(n3310), .S0(\i_MIPS/ID_EX_5 ), .Y(
        n10129) );
  AOI21X2 U1066 ( .A0(n4713), .A1(n3827), .B0(n3310), .Y(n6621) );
  NAND2X6 U1067 ( .A(n4159), .B(n4160), .Y(n6589) );
  INVX8 U1068 ( .A(n10379), .Y(n10366) );
  NAND2X8 U1069 ( .A(n4564), .B(n10379), .Y(n10352) );
  INVX6 U1070 ( .A(n6351), .Y(n6350) );
  BUFX20 U1071 ( .A(n5232), .Y(n5203) );
  INVX20 U1072 ( .A(n4318), .Y(DCACHE_addr[1]) );
  AOI22X4 U1073 ( .A0(net99639), .A1(net113039), .B0(net102300), .B1(n8581), 
        .Y(n3312) );
  OA22X4 U1074 ( .A0(net112493), .A1(n461), .B0(net112353), .B1(n2015), .Y(
        n9243) );
  OA22X2 U1075 ( .A0(net112493), .A1(n1421), .B0(net112369), .B1(n3034), .Y(
        n9097) );
  OA22X2 U1076 ( .A0(net112493), .A1(n1262), .B0(net112369), .B1(n2873), .Y(
        n9093) );
  OA22X2 U1077 ( .A0(net112493), .A1(n1362), .B0(net112369), .B1(n2975), .Y(
        n9089) );
  OA22X2 U1078 ( .A0(net112493), .A1(n1265), .B0(net112369), .B1(n2876), .Y(
        n9085) );
  BUFX16 U1079 ( .A(net112497), .Y(net112493) );
  BUFX8 U1080 ( .A(n7101), .Y(n157) );
  INVX20 U1081 ( .A(n9225), .Y(n9118) );
  NAND2X2 U1082 ( .A(n4653), .B(n4583), .Y(n9225) );
  BUFX8 U1083 ( .A(n7877), .Y(n159) );
  NAND2X2 U1084 ( .A(n6567), .B(\i_MIPS/n353 ), .Y(n7877) );
  NAND3BX4 U1085 ( .AN(n6641), .B(n6928), .C(n6640), .Y(n8894) );
  AND3X8 U1086 ( .A(n4607), .B(n6642), .C(n6928), .Y(n4606) );
  INVX8 U1087 ( .A(n6931), .Y(n6928) );
  INVX16 U1088 ( .A(n8153), .Y(n8527) );
  NAND2X6 U1089 ( .A(n10302), .B(n10301), .Y(n10915) );
  NAND2X4 U1090 ( .A(n11085), .B(n11083), .Y(n10301) );
  CLKAND2X4 U1091 ( .A(n4927), .B(n3574), .Y(n3572) );
  NOR3X4 U1092 ( .A(n10707), .B(n10706), .C(n162), .Y(n10708) );
  BUFX6 U1093 ( .A(n7102), .Y(n158) );
  OAI33X2 U1094 ( .A0(n9182), .A1(n4592), .A2(n9262), .B0(n9180), .B1(n4592), 
        .B2(n3600), .Y(n9187) );
  INVX4 U1095 ( .A(n160), .Y(n9620) );
  INVX12 U1096 ( .A(n7093), .Y(n6934) );
  NAND2X8 U1097 ( .A(n6847), .B(n6850), .Y(n7093) );
  INVX8 U1098 ( .A(n10210), .Y(n3598) );
  NAND2X8 U1099 ( .A(n11059), .B(n11047), .Y(n10210) );
  CLKINVX4 U1100 ( .A(n10493), .Y(n10495) );
  AO21X2 U1101 ( .A0(n10304), .A1(n10305), .B0(n10303), .Y(n10909) );
  INVX4 U1102 ( .A(n10266), .Y(n10304) );
  INVX3 U1103 ( .A(n10928), .Y(n10927) );
  OAI211X2 U1104 ( .A0(n10926), .A1(n10925), .B0(n10924), .C0(n10923), .Y(
        n10928) );
  CLKBUFX8 U1105 ( .A(net100082), .Y(net112263) );
  BUFX6 U1106 ( .A(net100082), .Y(net112265) );
  CLKBUFX2 U1107 ( .A(net112265), .Y(net112221) );
  INVX4 U1108 ( .A(net112265), .Y(net112217) );
  INVX3 U1109 ( .A(net112221), .Y(net112213) );
  INVX8 U1110 ( .A(net112221), .Y(net112211) );
  NAND2X4 U1111 ( .A(n8252), .B(n9165), .Y(n8280) );
  INVX6 U1112 ( .A(n7954), .Y(n8252) );
  AOI33X2 U1113 ( .A0(n3318), .A1(n7980), .A2(n9258), .B0(n7964), .B1(n9258), 
        .B2(n3859), .Y(n7987) );
  NAND2X2 U1114 ( .A(\i_MIPS/EX_MEM_1 ), .B(n10146), .Y(net102120) );
  INVX8 U1115 ( .A(n10152), .Y(n10146) );
  CLKINVX4 U1116 ( .A(n9182), .Y(n9183) );
  OAI2BB1X4 U1117 ( .A0N(n9261), .A1N(n9257), .B0(n9256), .Y(n9182) );
  AO21X4 U1118 ( .A0(net99037), .A1(net99038), .B0(net112727), .Y(net105737)
         );
  AO21X4 U1119 ( .A0(net99037), .A1(net99038), .B0(net113077), .Y(net99019) );
  NAND2X6 U1120 ( .A(n10310), .B(n10309), .Y(n10913) );
  INVX4 U1121 ( .A(n10915), .Y(n10310) );
  MXI2X2 U1122 ( .A(n4708), .B(\i_MIPS/n224 ), .S0(n5510), .Y(\i_MIPS/n500 )
         );
  NAND2X6 U1123 ( .A(n7875), .B(\i_MIPS/n340 ), .Y(n7789) );
  INVX6 U1124 ( .A(n6641), .Y(n6642) );
  NAND2X4 U1125 ( .A(n6936), .B(n8250), .Y(n6641) );
  AOI2BB1XL U1126 ( .A0N(n10918), .A1N(n10908), .B0(n10922), .Y(n10926) );
  NAND2X6 U1127 ( .A(n11099), .B(n11098), .Y(n10908) );
  OAI211X2 U1128 ( .A0(n3892), .A1(n3603), .B0(n7458), .C0(n7457), .Y(n7460)
         );
  NAND3X8 U1129 ( .A(ICACHE_addr[16]), .B(ICACHE_addr[15]), .C(n9364), .Y(
        n10289) );
  OA22X4 U1130 ( .A0(n5450), .A1(n1970), .B0(n5378), .B1(n398), .Y(n5961) );
  CLKBUFX8 U1131 ( .A(n5405), .Y(n5378) );
  AOI221X2 U1132 ( .A0(net112217), .A1(\D_cache/cache[4][128] ), .B0(net112121), .B1(\D_cache/cache[5][128] ), .C0(n3829), .Y(n3828) );
  NAND3BX4 U1133 ( .AN(n8525), .B(n7852), .C(n6635), .Y(n6636) );
  NAND2X4 U1134 ( .A(n10304), .B(n10268), .Y(n10308) );
  CLKINVX6 U1135 ( .A(n10267), .Y(n10268) );
  NAND3X4 U1136 ( .A(n4208), .B(n4209), .C(n1224), .Y(n6247) );
  AND3X4 U1137 ( .A(n6933), .B(n1224), .C(n6934), .Y(n1613) );
  BUFX3 U1138 ( .A(n9427), .Y(n160) );
  OAI211X2 U1139 ( .A0(n10220), .A1(n10219), .B0(n10218), .C0(n10217), .Y(
        n10247) );
  OAI2BB2X1 U1140 ( .B0(\i_MIPS/n169 ), .B1(net110219), .A0N(n175), .A1N(
        n10956), .Y(\i_MIPS/N110 ) );
  NAND2XL U1141 ( .A(n9558), .B(n4005), .Y(n9427) );
  NAND4X2 U1142 ( .A(n9558), .B(n3637), .C(ICACHE_addr[5]), .D(n3645), .Y(
        n9332) );
  INVX6 U1143 ( .A(n9607), .Y(n9558) );
  INVX8 U1144 ( .A(n10877), .Y(n10874) );
  OA22X4 U1145 ( .A0(n10878), .A1(net140281), .B0(net98430), .B1(n10877), .Y(
        n10880) );
  XOR2X4 U1146 ( .A(n9452), .B(n3647), .Y(n10877) );
  INVX2 U1147 ( .A(n9578), .Y(n9547) );
  XOR2X4 U1148 ( .A(n11366), .B(n3645), .Y(n9578) );
  XOR3X2 U1149 ( .A(net111405), .B(n11025), .C(n11024), .Y(n11027) );
  NAND3BX4 U1150 ( .AN(n10963), .B(n10961), .C(n153), .Y(\i_MIPS/PC/n56 ) );
  NAND2X6 U1151 ( .A(n11079), .B(n11078), .Y(n10205) );
  XOR2X4 U1152 ( .A(n11377), .B(ICACHE_addr[18]), .Y(n9577) );
  INVX8 U1153 ( .A(n10320), .Y(n10201) );
  NAND3X6 U1154 ( .A(ICACHE_addr[20]), .B(ICACHE_addr[19]), .C(n10198), .Y(
        n10320) );
  XOR2X4 U1155 ( .A(n10714), .B(ICACHE_addr[28]), .Y(n10719) );
  XOR2X4 U1156 ( .A(n11365), .B(n3648), .Y(n4695) );
  CLKXOR2X4 U1157 ( .A(n10375), .B(ICACHE_addr[25]), .Y(n10380) );
  INVX8 U1158 ( .A(n10725), .Y(n10723) );
  OAI22X1 U1159 ( .A0(n10704), .A1(n10703), .B0(n10718), .B1(n10702), .Y(
        n10705) );
  NAND2X6 U1160 ( .A(n10702), .B(n10718), .Y(n10703) );
  INVXL U1161 ( .A(n10702), .Y(n10700) );
  BUFX3 U1162 ( .A(n10705), .Y(n162) );
  OA22X4 U1163 ( .A0(n10723), .A1(n10722), .B0(n10725), .B1(n10724), .Y(n10728) );
  NAND2X2 U1164 ( .A(n10713), .B(n168), .Y(n10722) );
  NAND2X2 U1165 ( .A(n10343), .B(net113551), .Y(n10344) );
  INVX6 U1166 ( .A(n10342), .Y(n10343) );
  XOR2X4 U1167 ( .A(n10719), .B(net111405), .Y(n10702) );
  NOR2X4 U1168 ( .A(n9551), .B(n3852), .Y(n9563) );
  NAND3X6 U1169 ( .A(n6450), .B(n6451), .C(n8802), .Y(n6236) );
  NAND2X6 U1170 ( .A(n3640), .B(n3641), .Y(n8924) );
  INVX1 U1171 ( .A(n8926), .Y(n3641) );
  NAND2X6 U1172 ( .A(n4132), .B(n4133), .Y(n4095) );
  INVX4 U1173 ( .A(n3601), .Y(n8823) );
  NAND2X4 U1174 ( .A(n9139), .B(n3787), .Y(n9286) );
  CLKBUFX3 U1175 ( .A(net112517), .Y(net112503) );
  NAND2X2 U1176 ( .A(n6778), .B(n4707), .Y(n8913) );
  NAND3X6 U1177 ( .A(n3534), .B(n3535), .C(n9172), .Y(n9177) );
  AND3X2 U1178 ( .A(n9171), .B(n9170), .C(n9169), .Y(n9172) );
  NAND2X4 U1179 ( .A(n9271), .B(n3787), .Y(n8539) );
  AND2X6 U1180 ( .A(n6246), .B(\i_MIPS/n360 ), .Y(n3704) );
  NAND2X4 U1181 ( .A(n9259), .B(n6669), .Y(n6656) );
  INVX3 U1182 ( .A(n7981), .Y(n7982) );
  INVX1 U1183 ( .A(n7863), .Y(n9287) );
  INVX3 U1184 ( .A(n4628), .Y(n4958) );
  CLKINVX1 U1185 ( .A(n7869), .Y(n8348) );
  BUFX4 U1186 ( .A(net112505), .Y(net112463) );
  BUFX12 U1187 ( .A(net100084), .Y(net112517) );
  NAND3BX2 U1188 ( .AN(n10130), .B(n10129), .C(n10132), .Y(n6200) );
  INVX2 U1189 ( .A(n7473), .Y(n8724) );
  MX2X1 U1190 ( .A(n9124), .B(n9123), .S0(n5587), .Y(n9125) );
  CLKINVX3 U1191 ( .A(net99039), .Y(net105736) );
  NAND3X6 U1192 ( .A(ICACHE_addr[14]), .B(ICACHE_addr[13]), .C(n9366), .Y(
        n10290) );
  AND2X2 U1193 ( .A(net109795), .B(n11390), .Y(n4178) );
  NAND4X2 U1194 ( .A(n6388), .B(n6387), .C(n6386), .D(n6385), .Y(n11464) );
  OA22X1 U1195 ( .A0(net112665), .A1(n2377), .B0(net112575), .B1(n873), .Y(
        n7242) );
  OA22X2 U1196 ( .A0(net112245), .A1(n2397), .B0(net112161), .B1(n892), .Y(
        n7240) );
  NAND4X2 U1197 ( .A(n8858), .B(n8857), .C(n8856), .D(n8855), .Y(n11454) );
  BUFX4 U1198 ( .A(net112519), .Y(net112497) );
  AO22X1 U1199 ( .A0(net113455), .A1(n11426), .B0(net113461), .B1(n11395), .Y(
        n7332) );
  INVX3 U1200 ( .A(n7711), .Y(n7713) );
  OR2X4 U1201 ( .A(n11112), .B(net110247), .Y(n3765) );
  NAND4X6 U1202 ( .A(n9629), .B(n9628), .C(n9627), .D(n9626), .Y(n10212) );
  NAND2X6 U1203 ( .A(n10648), .B(n10647), .Y(n6081) );
  NAND2X2 U1204 ( .A(n6846), .B(n7463), .Y(n7094) );
  NAND3X2 U1205 ( .A(n6936), .B(n7024), .C(n7031), .Y(n6472) );
  NAND2X4 U1206 ( .A(n4642), .B(n3771), .Y(n4427) );
  INVX4 U1207 ( .A(n6238), .Y(n6232) );
  INVX16 U1208 ( .A(n6243), .Y(n6228) );
  INVX1 U1209 ( .A(n4704), .Y(n3742) );
  NAND2X2 U1210 ( .A(n4809), .B(\i_MIPS/ALUin1[18] ), .Y(n7871) );
  NOR2X6 U1211 ( .A(\i_MIPS/n362 ), .B(n6230), .Y(n3817) );
  NAND2X4 U1212 ( .A(n6570), .B(\i_MIPS/n356 ), .Y(n7030) );
  CLKINVX8 U1213 ( .A(n6613), .Y(n6570) );
  AND2X8 U1214 ( .A(n7846), .B(n159), .Y(n4515) );
  NAND2X4 U1215 ( .A(n6578), .B(\i_MIPS/n351 ), .Y(n8543) );
  BUFX4 U1216 ( .A(n9311), .Y(n4982) );
  NAND2X4 U1217 ( .A(net99089), .B(net99090), .Y(n4078) );
  INVX3 U1218 ( .A(n4886), .Y(n4885) );
  BUFX12 U1219 ( .A(n4631), .Y(n4808) );
  CLKINVX1 U1220 ( .A(n9014), .Y(n9163) );
  AND2X4 U1221 ( .A(n4691), .B(\i_MIPS/ALUin1[25] ), .Y(n4666) );
  NAND2X6 U1222 ( .A(n4418), .B(n4419), .Y(n6237) );
  BUFX4 U1223 ( .A(net100084), .Y(net112515) );
  CLKINVX1 U1224 ( .A(n4413), .Y(n4414) );
  NAND2X6 U1225 ( .A(\i_MIPS/ALUin1[18] ), .B(n6567), .Y(n7853) );
  NAND2X2 U1226 ( .A(n4821), .B(\i_MIPS/ALUin1[7] ), .Y(n7281) );
  NAND2X4 U1227 ( .A(n3661), .B(n3662), .Y(n9611) );
  NAND2X6 U1228 ( .A(n4728), .B(\i_MIPS/PC/n4 ), .Y(n3662) );
  OAI22X2 U1229 ( .A0(n7610), .A1(n4802), .B0(n7611), .B1(n7869), .Y(n7613) );
  CLKINVX6 U1230 ( .A(n7028), .Y(n7710) );
  NAND2X6 U1231 ( .A(n4508), .B(n11010), .Y(n10322) );
  BUFX12 U1232 ( .A(n4889), .Y(n4891) );
  NAND2X4 U1233 ( .A(n10661), .B(n10660), .Y(n3718) );
  CLKINVX6 U1234 ( .A(net112511), .Y(n3560) );
  OAI221XL U1235 ( .A0(\i_MIPS/Register/register[2][3] ), .A1(n4921), .B0(
        \i_MIPS/Register/register[10][3] ), .B1(n4917), .C0(n8746), .Y(n8749)
         );
  AO22X1 U1236 ( .A0(n4898), .A1(n332), .B0(n4893), .B1(n1909), .Y(n8567) );
  NAND4BX2 U1237 ( .AN(n7773), .B(n7772), .C(n7771), .D(n7770), .Y(n7774) );
  NAND3X2 U1238 ( .A(n3841), .B(n3842), .C(n6367), .Y(n6371) );
  AOI221X1 U1239 ( .A0(n9259), .A1(n6349), .B0(n4636), .B1(n9258), .C0(n4800), 
        .Y(n6374) );
  AND2X6 U1240 ( .A(n3599), .B(n8342), .Y(n3579) );
  AND2X2 U1241 ( .A(n9283), .B(n9282), .Y(n4634) );
  INVX1 U1242 ( .A(n3529), .Y(n7457) );
  CLKMX2X3 U1243 ( .A(\i_MIPS/n340 ), .B(\i_MIPS/n341 ), .S0(n4809), .Y(n7874)
         );
  AO22X2 U1244 ( .A0(n9312), .A1(n341), .B0(n4981), .B1(n1922), .Y(n7413) );
  INVX3 U1245 ( .A(n7876), .Y(n8350) );
  NAND2X6 U1246 ( .A(n7200), .B(n3787), .Y(n8814) );
  OAI22X2 U1247 ( .A0(n5428), .A1(n308), .B0(n5384), .B1(n1876), .Y(n4449) );
  BUFX8 U1248 ( .A(n11139), .Y(n5407) );
  AND2X4 U1249 ( .A(n10161), .B(n10146), .Y(n4514) );
  INVX16 U1250 ( .A(n4813), .Y(n4812) );
  INVX12 U1251 ( .A(n3700), .Y(n6216) );
  INVX4 U1252 ( .A(n3708), .Y(n6209) );
  NAND2X4 U1253 ( .A(n6566), .B(\i_MIPS/n354 ), .Y(n7846) );
  NAND2X4 U1254 ( .A(n4507), .B(n10326), .Y(n10498) );
  CLKINVX3 U1255 ( .A(net102088), .Y(net113081) );
  BUFX6 U1256 ( .A(net102371), .Y(net113457) );
  BUFX4 U1257 ( .A(n5314), .Y(n5302) );
  CLKAND2X8 U1258 ( .A(n4152), .B(n4153), .Y(n5995) );
  OA22X1 U1259 ( .A0(net112245), .A1(n2384), .B0(net112161), .B1(n879), .Y(
        n7497) );
  NOR2X2 U1260 ( .A(n4206), .B(n4207), .Y(n6113) );
  INVX3 U1261 ( .A(n4211), .Y(n3678) );
  AOI2BB2X2 U1262 ( .B0(net111873), .B1(\D_cache/cache[7][131] ), .A0N(
        net112037), .A1N(n1900), .Y(n6117) );
  INVX4 U1263 ( .A(n6092), .Y(n10656) );
  AOI22X2 U1264 ( .A0(n3813), .A1(\D_cache/cache[2][136] ), .B0(n3814), .B1(
        \D_cache/cache[3][136] ), .Y(n6038) );
  INVX3 U1265 ( .A(net112301), .Y(n3814) );
  INVX3 U1266 ( .A(n6041), .Y(n10634) );
  INVX6 U1267 ( .A(n6085), .Y(n10650) );
  CLKMX2X2 U1268 ( .A(n4799), .B(n9141), .S0(n7179), .Y(n6780) );
  NOR4X2 U1269 ( .A(n6681), .B(n6680), .C(n6679), .D(n6678), .Y(n6682) );
  NAND3X6 U1270 ( .A(ICACHE_addr[10]), .B(ICACHE_addr[9]), .C(n10202), .Y(
        n10263) );
  NAND4BX1 U1271 ( .AN(n8128), .B(n8127), .C(n8126), .D(n8125), .Y(n8139) );
  OAI221XL U1272 ( .A0(\i_MIPS/Register/register[2][21] ), .A1(n4946), .B0(
        \i_MIPS/Register/register[10][21] ), .B1(n4939), .C0(n8120), .Y(n8128)
         );
  NAND4X4 U1273 ( .A(n7985), .B(n7987), .C(n7984), .D(n7986), .Y(net99407) );
  NAND2X6 U1274 ( .A(n8818), .B(n4707), .Y(n7544) );
  AND3X6 U1275 ( .A(n3781), .B(n3782), .C(n8813), .Y(n3689) );
  BUFX16 U1276 ( .A(net110259), .Y(net110257) );
  NAND3X6 U1277 ( .A(n3629), .B(n3630), .C(n7671), .Y(net104829) );
  OA22X1 U1278 ( .A0(net112237), .A1(n946), .B0(net112155), .B1(n2471), .Y(
        n8678) );
  OA22X2 U1279 ( .A0(net112667), .A1(n2408), .B0(net112565), .B1(n902), .Y(
        n8291) );
  OA22X2 U1280 ( .A0(net112673), .A1(n2376), .B0(net112575), .B1(n872), .Y(
        n7144) );
  OA22X2 U1281 ( .A0(net112245), .A1(n2396), .B0(net112161), .B1(n891), .Y(
        n7142) );
  OA22XL U1282 ( .A0(net112233), .A1(n936), .B0(net112165), .B1(n2461), .Y(
        n6794) );
  NAND4X2 U1283 ( .A(net105020), .B(net105021), .C(net105022), .D(net105023), 
        .Y(net98121) );
  NAND4X4 U1284 ( .A(n8688), .B(n8687), .C(n8686), .D(n8685), .Y(n11509) );
  OA22X2 U1285 ( .A0(net112075), .A1(n2399), .B0(net111951), .B1(n894), .Y(
        n8685) );
  OA22X2 U1286 ( .A0(net112667), .A1(n2409), .B0(net112565), .B1(n903), .Y(
        n8400) );
  AOI2BB2X1 U1287 ( .B0(net111873), .B1(\D_cache/cache[7][18] ), .A0N(
        net112065), .A1N(n2316), .Y(n7924) );
  NAND4X2 U1288 ( .A(n8206), .B(n8205), .C(n8204), .D(n8203), .Y(n11498) );
  OA22XL U1289 ( .A0(net112673), .A1(n804), .B0(net112575), .B1(n2351), .Y(
        n6975) );
  AO22XL U1290 ( .A0(net113455), .A1(n11430), .B0(net113461), .B1(n11399), .Y(
        n7248) );
  NAND2XL U1291 ( .A(DCACHE_addr[1]), .B(\i_MIPS/n336 ), .Y(net100103) );
  CLKMX2X2 U1292 ( .A(n9081), .B(n9080), .S0(net108959), .Y(n9082) );
  INVX1 U1293 ( .A(net112721), .Y(n3621) );
  AO22XL U1294 ( .A0(net113455), .A1(n11451), .B0(net113461), .B1(n11420), .Y(
        n9100) );
  INVX3 U1295 ( .A(n9275), .Y(n8820) );
  INVX3 U1296 ( .A(n10215), .Y(n11074) );
  INVX2 U1297 ( .A(n10920), .Y(n11094) );
  NAND2X4 U1298 ( .A(n10582), .B(n10581), .Y(n4445) );
  INVXL U1299 ( .A(n4518), .Y(n3697) );
  OAI221X1 U1300 ( .A0(n4519), .A1(n8886), .B0(n9275), .B1(n8439), .C0(n4501), 
        .Y(n8446) );
  NOR4X1 U1301 ( .A(n7302), .B(n7301), .C(n7300), .D(n7299), .Y(n7313) );
  OA22X2 U1302 ( .A0(net112237), .A1(n2369), .B0(net112153), .B1(n373), .Y(
        n6532) );
  INVX12 U1303 ( .A(net109181), .Y(net113605) );
  OA22X1 U1304 ( .A0(net112245), .A1(n2382), .B0(net112161), .B1(n877), .Y(
        n7394) );
  OA22X1 U1305 ( .A0(net112245), .A1(n2386), .B0(net112161), .B1(n881), .Y(
        n7485) );
  OA22X1 U1306 ( .A0(net112233), .A1(n2412), .B0(net112151), .B1(n904), .Y(
        n8192) );
  OA22X1 U1307 ( .A0(net112485), .A1(n2359), .B0(net112361), .B1(n856), .Y(
        n8584) );
  OA22X1 U1308 ( .A0(net112233), .A1(n2411), .B0(net112151), .B1(n383), .Y(
        n8103) );
  NAND4X2 U1309 ( .A(n8388), .B(n8387), .C(n8386), .D(n8385), .Y(n11446) );
  NAND4X4 U1310 ( .A(n9252), .B(n9251), .C(n9250), .D(n9249), .Y(n11450) );
  OA22XL U1311 ( .A0(net112673), .A1(n1958), .B0(net112571), .B1(n386), .Y(
        n9252) );
  OA22X2 U1312 ( .A0(net112083), .A1(n1948), .B0(net111959), .B1(n370), .Y(
        n9249) );
  OA22X1 U1313 ( .A0(net112237), .A1(n2363), .B0(net112153), .B1(n860), .Y(
        n6278) );
  OA22X2 U1314 ( .A0(net112473), .A1(n2358), .B0(net112349), .B1(n855), .Y(
        n7728) );
  OA22X1 U1315 ( .A0(net112663), .A1(n953), .B0(net112561), .B1(n2478), .Y(
        n7818) );
  OA22X2 U1316 ( .A0(net112075), .A1(n2403), .B0(net111951), .B1(n897), .Y(
        n8681) );
  OA22X2 U1317 ( .A0(net112487), .A1(n2405), .B0(net112363), .B1(n899), .Y(
        n8683) );
  OA22X1 U1318 ( .A0(net112245), .A1(n2368), .B0(net112153), .B1(n865), .Y(
        n6540) );
  OA22X1 U1319 ( .A0(net112077), .A1(n2357), .B0(net111953), .B1(n854), .Y(
        n8774) );
  OA22X1 U1320 ( .A0(net112245), .A1(n2380), .B0(net112161), .B1(n876), .Y(
        n7328) );
  OA22X2 U1321 ( .A0(net112233), .A1(n2410), .B0(net112151), .B1(n382), .Y(
        n8022) );
  INVX6 U1322 ( .A(net113605), .Y(net113916) );
  AND2XL U1323 ( .A(n3613), .B(net99450), .Y(n4556) );
  MXI2X1 U1324 ( .A(n7755), .B(n7754), .S0(n5588), .Y(n3840) );
  INVX3 U1325 ( .A(net99583), .Y(net106109) );
  AND2XL U1326 ( .A(net98973), .B(net98974), .Y(n4538) );
  OR2X4 U1327 ( .A(n11077), .B(net110247), .Y(n3606) );
  INVX4 U1328 ( .A(n10698), .Y(n10699) );
  INVX6 U1329 ( .A(n10900), .Y(n10897) );
  OR2X2 U1330 ( .A(n151), .B(net110249), .Y(n3544) );
  AND2XL U1331 ( .A(net99814), .B(net99815), .Y(n4537) );
  NAND2X1 U1332 ( .A(\i_MIPS/IF_ID[66] ), .B(n147), .Y(n10833) );
  INVXL U1333 ( .A(net104829), .Y(net98901) );
  INVX4 U1334 ( .A(n11063), .Y(n11069) );
  INVX16 U1335 ( .A(n4130), .Y(net110243) );
  XOR3X2 U1336 ( .A(net111409), .B(n11016), .C(n11020), .Y(n11018) );
  XOR3X2 U1337 ( .A(net111405), .B(n11110), .C(n11109), .Y(n11112) );
  NAND2BX2 U1338 ( .AN(n11108), .B(n11107), .Y(n11109) );
  BUFX4 U1339 ( .A(net110231), .Y(net110217) );
  NAND2BX1 U1340 ( .AN(n5461), .B(n11274), .Y(n10101) );
  OAI2BB2XL U1341 ( .B0(\i_MIPS/n241 ), .B1(net110219), .A0N(n173), .A1N(n9630), .Y(\i_MIPS/N95 ) );
  NAND2X4 U1342 ( .A(n6642), .B(n6932), .Y(n8890) );
  INVX4 U1343 ( .A(n8332), .Y(n8329) );
  INVX3 U1344 ( .A(n6593), .Y(n6614) );
  NAND2X6 U1345 ( .A(n7355), .B(n7271), .Y(n7452) );
  NAND2X6 U1346 ( .A(\i_MIPS/ALUin1[1] ), .B(n7619), .Y(n6451) );
  CLKINVX1 U1347 ( .A(n8891), .Y(n6637) );
  CLKINVX1 U1348 ( .A(n8250), .Y(n8893) );
  AND2X4 U1349 ( .A(n4658), .B(n4653), .Y(n4619) );
  AND2X2 U1350 ( .A(\i_MIPS/n231 ), .B(\i_MIPS/n230 ), .Y(n4581) );
  NAND2X6 U1351 ( .A(n7107), .B(n6598), .Y(n6601) );
  INVX1 U1352 ( .A(n8894), .Y(n8895) );
  INVX4 U1353 ( .A(n6658), .Y(n6659) );
  AND4X4 U1354 ( .A(n4516), .B(n8329), .C(n6614), .D(n8327), .Y(n4412) );
  AND2X2 U1355 ( .A(n8252), .B(n8331), .Y(n2802) );
  INVX4 U1356 ( .A(n6596), .Y(n9168) );
  CLKINVX6 U1357 ( .A(n7798), .Y(n6575) );
  INVX6 U1358 ( .A(n4099), .Y(n4131) );
  NAND2X1 U1359 ( .A(net134109), .B(net99019), .Y(n4085) );
  CLKAND2X8 U1360 ( .A(\i_MIPS/IR_ID[23] ), .B(\i_MIPS/n231 ), .Y(n4655) );
  AND2X4 U1361 ( .A(\i_MIPS/n229 ), .B(\i_MIPS/n228 ), .Y(n4583) );
  NAND2X4 U1362 ( .A(\i_MIPS/n299 ), .B(n3770), .Y(n4418) );
  NAND3X4 U1363 ( .A(n3752), .B(n3671), .C(net113533), .Y(net134088) );
  AOI211X1 U1364 ( .A0(n6456), .A1(n3796), .B0(n3792), .C0(n6455), .Y(n6457)
         );
  INVX4 U1365 ( .A(n9549), .Y(n9580) );
  AND2X2 U1366 ( .A(n7562), .B(n7477), .Y(n4522) );
  NAND2X4 U1367 ( .A(n7099), .B(n6638), .Y(n6931) );
  INVX3 U1368 ( .A(n7958), .Y(n6619) );
  INVX4 U1369 ( .A(n10208), .Y(n10307) );
  CLKAND2X8 U1370 ( .A(\i_MIPS/IR_ID[22] ), .B(\i_MIPS/n228 ), .Y(n4500) );
  AND2X4 U1371 ( .A(\i_MIPS/IR_ID[24] ), .B(\i_MIPS/n230 ), .Y(n4653) );
  NAND2X2 U1372 ( .A(n10653), .B(n1637), .Y(n6090) );
  NAND2X2 U1373 ( .A(n283), .B(n3778), .Y(n3779) );
  NAND2X2 U1374 ( .A(n12956), .B(n6081), .Y(n3780) );
  NAND2X4 U1375 ( .A(n3734), .B(n10664), .Y(n6148) );
  NAND2X2 U1376 ( .A(n12953), .B(n6152), .Y(n3683) );
  NAND2X2 U1377 ( .A(n4752), .B(n3681), .Y(n3682) );
  INVX3 U1378 ( .A(n6152), .Y(n3681) );
  NAND2X4 U1379 ( .A(n1632), .B(n3297), .Y(n6126) );
  NAND2X2 U1380 ( .A(n2437), .B(n10673), .Y(n6134) );
  INVX8 U1381 ( .A(n9335), .Y(n9582) );
  OAI221XL U1382 ( .A0(\i_MIPS/Register/register[2][19] ), .A1(n4922), .B0(
        \i_MIPS/Register/register[10][19] ), .B1(n4915), .C0(n7756), .Y(n7764)
         );
  OAI221XL U1383 ( .A0(\i_MIPS/Register/register[18][19] ), .A1(n4922), .B0(
        \i_MIPS/Register/register[26][19] ), .B1(n4916), .C0(n7765), .Y(n7773)
         );
  AND2X2 U1384 ( .A(n4821), .B(\i_MIPS/n354 ), .Y(n4612) );
  CLKAND2X3 U1385 ( .A(n4814), .B(\i_MIPS/n355 ), .Y(n4597) );
  NAND2X1 U1386 ( .A(n4828), .B(\i_MIPS/n353 ), .Y(n7022) );
  MX2X6 U1387 ( .A(\i_MIPS/n303 ), .B(n6209), .S0(n5594), .Y(n6238) );
  NOR2BX2 U1388 ( .AN(n4815), .B(\i_MIPS/n354 ), .Y(n4690) );
  NOR3X4 U1389 ( .A(n3843), .B(n3844), .C(n3845), .Y(n6367) );
  AND2X2 U1390 ( .A(n6365), .B(n3636), .Y(n3844) );
  NAND2X1 U1391 ( .A(n7279), .B(n6944), .Y(n3841) );
  NOR2BX1 U1392 ( .AN(n4809), .B(\i_MIPS/n340 ), .Y(n4683) );
  CLKMX2X2 U1393 ( .A(n6852), .B(n6851), .S0(n5590), .Y(n7610) );
  OA22X2 U1394 ( .A0(n8659), .A1(n7183), .B0(n8728), .B1(n8438), .Y(n6860) );
  OAI2BB1X1 U1395 ( .A0N(n6848), .A1N(n6847), .B0(n6846), .Y(n6849) );
  INVX3 U1396 ( .A(n7103), .Y(n7784) );
  INVX3 U1397 ( .A(n7462), .Y(n6240) );
  NAND2X2 U1398 ( .A(n8645), .B(n8646), .Y(n9173) );
  CLKBUFX3 U1399 ( .A(n4991), .Y(n4989) );
  OA22X1 U1400 ( .A0(\i_MIPS/Register/register[6][28] ), .A1(n4914), .B0(
        \i_MIPS/Register/register[14][28] ), .B1(n4908), .Y(n9028) );
  NAND4X1 U1401 ( .A(n9027), .B(n9026), .C(n9025), .D(n9024), .Y(n9032) );
  NAND2X4 U1402 ( .A(\i_MIPS/ALUin1[6] ), .B(n3821), .Y(n7545) );
  NAND2X2 U1403 ( .A(n3198), .B(net100013), .Y(n4076) );
  NAND2X6 U1404 ( .A(n6233), .B(\i_MIPS/ALUin1[2] ), .Y(n8802) );
  INVX4 U1405 ( .A(n3759), .Y(n8803) );
  CLKBUFX3 U1406 ( .A(n4991), .Y(n4990) );
  CLKBUFX3 U1407 ( .A(n4933), .Y(n4936) );
  AND2X4 U1408 ( .A(\i_MIPS/IR_ID[18] ), .B(\i_MIPS/n318 ), .Y(n4656) );
  CLKMX2X4 U1409 ( .A(n8888), .B(n8533), .S0(n5589), .Y(n9005) );
  AND2X4 U1410 ( .A(n9003), .B(n9130), .Y(n3784) );
  AND2X2 U1411 ( .A(n4800), .B(n9018), .Y(n3785) );
  NAND2X4 U1412 ( .A(n4655), .B(n4583), .Y(n9224) );
  NAND2X4 U1413 ( .A(\i_MIPS/ALUin1[5] ), .B(n6237), .Y(n7454) );
  AND2X2 U1414 ( .A(mem_ready_D), .B(n11514), .Y(n4669) );
  AND2X2 U1415 ( .A(n3238), .B(n4047), .Y(n4589) );
  BUFX4 U1416 ( .A(net100087), .Y(net112599) );
  INVX6 U1417 ( .A(n10139), .Y(n10161) );
  BUFX12 U1418 ( .A(net112705), .Y(net112701) );
  INVX3 U1419 ( .A(n6509), .Y(n9313) );
  NAND2X4 U1420 ( .A(n10147), .B(\i_MIPS/EX_MEM_1 ), .Y(net102121) );
  NAND2X2 U1421 ( .A(n4589), .B(\i_MIPS/EX_MEM_1 ), .Y(net102094) );
  NAND2X1 U1422 ( .A(n352), .B(\i_MIPS/EX_MEM_1 ), .Y(net102095) );
  NAND2X6 U1423 ( .A(DCACHE_ren), .B(n11389), .Y(net100096) );
  BUFX6 U1424 ( .A(n4450), .Y(n5365) );
  BUFX8 U1425 ( .A(n11138), .Y(n5276) );
  NAND2X1 U1426 ( .A(n4648), .B(n3826), .Y(n4160) );
  NAND2X2 U1427 ( .A(\i_MIPS/n261 ), .B(n4158), .Y(n4159) );
  AOI2BB1X1 U1428 ( .A0N(n6466), .A1N(n7187), .B0(n6465), .Y(n6467) );
  CLKINVX1 U1429 ( .A(n7025), .Y(n6463) );
  NAND2X2 U1430 ( .A(n7777), .B(n8143), .Y(n6634) );
  AND4X6 U1431 ( .A(\i_MIPS/ID_EX[108] ), .B(\i_MIPS/n333 ), .C(\i_MIPS/n331 ), 
        .D(n4413), .Y(\i_MIPS/ALU_Control/n11 ) );
  INVX3 U1432 ( .A(n10314), .Y(n10912) );
  OAI211X1 U1433 ( .A0(n8349), .A1(n7880), .B0(n7879), .C0(n4501), .Y(n7881)
         );
  CLKMX2X2 U1434 ( .A(n9280), .B(n9279), .S0(n7878), .Y(n7879) );
  AO22X2 U1435 ( .A0(n9271), .A1(n7876), .B0(n4568), .B1(n9267), .Y(n7882) );
  INVX3 U1436 ( .A(n7885), .Y(n7886) );
  INVX6 U1437 ( .A(n6566), .Y(n6574) );
  NAND2X4 U1438 ( .A(n6573), .B(\i_MIPS/n355 ), .Y(n8143) );
  INVX4 U1439 ( .A(n6589), .Y(n6592) );
  INVX4 U1440 ( .A(n6586), .Y(n6591) );
  AO21X2 U1441 ( .A0(\i_MIPS/ID_EX[80] ), .A1(\i_MIPS/ALU/N303 ), .B0(n6356), 
        .Y(n7286) );
  AND3X4 U1442 ( .A(n10307), .B(n10306), .C(n3598), .Y(n10312) );
  INVX4 U1443 ( .A(n4869), .Y(n4867) );
  INVX4 U1444 ( .A(n4888), .Y(n4884) );
  INVX4 U1445 ( .A(n4878), .Y(n4876) );
  XOR2X1 U1446 ( .A(n10132), .B(\i_MIPS/IR_ID[23] ), .Y(n6296) );
  XOR2X1 U1447 ( .A(n6292), .B(\i_MIPS/IR_ID[21] ), .Y(n6295) );
  NAND4X1 U1448 ( .A(n6290), .B(n6289), .C(n6288), .D(n6287), .Y(n6304) );
  AND4X6 U1449 ( .A(n8327), .B(n7950), .C(n4515), .D(n4801), .Y(n3772) );
  NAND2X2 U1450 ( .A(\i_MIPS/ALUin1[21] ), .B(n6581), .Y(n8080) );
  CLKINVX1 U1451 ( .A(n7279), .Y(n8087) );
  INVX6 U1452 ( .A(n4870), .Y(n4866) );
  INVX6 U1453 ( .A(n4847), .Y(n4842) );
  INVX6 U1454 ( .A(n4878), .Y(n4875) );
  INVX6 U1455 ( .A(n4887), .Y(n4883) );
  INVX4 U1456 ( .A(n4888), .Y(n4881) );
  INVX4 U1457 ( .A(n4879), .Y(n4873) );
  INVX4 U1458 ( .A(n4872), .Y(n4864) );
  NAND4X4 U1459 ( .A(n4472), .B(n4473), .C(n5951), .D(n4474), .Y(n9572) );
  AOI2BB2X2 U1460 ( .B0(n4675), .B1(\I_cache/cache[5][154] ), .A0N(n5357), 
        .A1N(n3207), .Y(n5951) );
  OR2X1 U1461 ( .A(net112145), .B(n2023), .Y(n4220) );
  OR2X6 U1462 ( .A(net112659), .B(n1879), .Y(n4211) );
  BUFX4 U1463 ( .A(net112509), .Y(net112427) );
  AO22X1 U1464 ( .A0(n4971), .A1(n326), .B0(n4965), .B1(n1903), .Y(n6911) );
  AO22X1 U1465 ( .A0(n4991), .A1(n338), .B0(n4984), .B1(n1915), .Y(n6909) );
  AO22X1 U1466 ( .A0(n4971), .A1(n232), .B0(n4965), .B1(n1927), .Y(n6920) );
  AO22X1 U1467 ( .A0(n4991), .A1(n349), .B0(n4984), .B1(n1931), .Y(n6918) );
  INVX3 U1468 ( .A(n8156), .Y(n8155) );
  NAND3BX1 U1469 ( .AN(n4615), .B(n8141), .C(n8140), .Y(n8533) );
  AOI2BB1X1 U1470 ( .A0N(\i_MIPS/ALUin1[16] ), .A1N(n4806), .B0(n4600), .Y(
        n8140) );
  NAND2X4 U1471 ( .A(\i_MIPS/ALUin1[3] ), .B(n6238), .Y(n8712) );
  NAND2X6 U1472 ( .A(n6939), .B(n6947), .Y(n7025) );
  NAND2X2 U1473 ( .A(n3827), .B(n6612), .Y(n7024) );
  NAND2X4 U1474 ( .A(n6350), .B(\i_MIPS/n358 ), .Y(n6632) );
  NAND2X2 U1475 ( .A(n6351), .B(\i_MIPS/n358 ), .Y(n6603) );
  NAND2X1 U1476 ( .A(\i_MIPS/ALUin1[13] ), .B(n6350), .Y(n6609) );
  NAND2X2 U1477 ( .A(n7183), .B(n7184), .Y(n7191) );
  CLKMX2X2 U1478 ( .A(n8272), .B(n7793), .S0(n5589), .Y(n8665) );
  CLKINVX1 U1479 ( .A(n8262), .Y(n7793) );
  INVX3 U1480 ( .A(n7787), .Y(n8641) );
  AOI21X2 U1481 ( .A0(n6845), .A1(n7179), .B0(n6844), .Y(n4570) );
  CLKINVX1 U1482 ( .A(n6849), .Y(n3627) );
  NAND2X4 U1483 ( .A(n6229), .B(\i_MIPS/n362 ), .Y(n6850) );
  INVX3 U1484 ( .A(n6230), .Y(n6229) );
  INVX3 U1485 ( .A(n6462), .Y(n3747) );
  INVX3 U1486 ( .A(n3817), .Y(n7183) );
  AOI221X1 U1487 ( .A0(n4924), .A1(n6849), .B0(n4570), .B1(n9258), .C0(n4800), 
        .Y(n6865) );
  NAND2X4 U1488 ( .A(n6245), .B(\i_MIPS/n360 ), .Y(n7100) );
  OA22X1 U1489 ( .A0(\i_MIPS/ALUin1[8] ), .A1(n4811), .B0(\i_MIPS/ALUin1[7] ), 
        .B1(n4804), .Y(n7472) );
  INVX3 U1490 ( .A(n7456), .Y(n7464) );
  INVX3 U1491 ( .A(n4820), .Y(n4819) );
  OAI222XL U1492 ( .A0(n9007), .A1(n6673), .B0(n6672), .B1(n8805), .C0(n8086), 
        .C1(n9004), .Y(n6680) );
  CLKINVX1 U1493 ( .A(n6656), .Y(n6653) );
  CLKINVX1 U1494 ( .A(n7802), .Y(n7786) );
  CLKMX2X2 U1495 ( .A(n9280), .B(n9279), .S0(n8519), .Y(n7782) );
  NOR4X1 U1496 ( .A(n7839), .B(n7838), .C(n7837), .D(n7836), .Y(n7840) );
  AO22X1 U1497 ( .A0(n9312), .A1(n289), .B0(n4985), .B1(n1859), .Y(n7837) );
  AO22X1 U1498 ( .A0(n5000), .A1(n234), .B0(n4996), .B1(n1832), .Y(n7836) );
  OAI221XL U1499 ( .A0(\i_MIPS/Register/register[2][19] ), .A1(n4946), .B0(
        \i_MIPS/Register/register[10][19] ), .B1(n4939), .C0(n7826), .Y(n7834)
         );
  NOR4X1 U1500 ( .A(n7830), .B(n7829), .C(n7828), .D(n7827), .Y(n7831) );
  AO22X1 U1501 ( .A0(n9312), .A1(n236), .B0(n4985), .B1(n1861), .Y(n7828) );
  AO22X1 U1502 ( .A0(n5000), .A1(n235), .B0(n4996), .B1(n1833), .Y(n7827) );
  AO22X1 U1503 ( .A0(n4978), .A1(n290), .B0(n4976), .B1(n1860), .Y(n7829) );
  OA22X1 U1504 ( .A0(\i_MIPS/Register/register[22][20] ), .A1(n4938), .B0(
        \i_MIPS/Register/register[30][20] ), .B1(n4931), .Y(n8609) );
  OA22X1 U1505 ( .A0(\i_MIPS/Register/register[6][20] ), .A1(n4938), .B0(
        \i_MIPS/Register/register[14][20] ), .B1(n4931), .Y(n8600) );
  OAI221XL U1506 ( .A0(\i_MIPS/Register/register[2][24] ), .A1(n4947), .B0(
        \i_MIPS/Register/register[10][24] ), .B1(n4940), .C0(n8975), .Y(n8983)
         );
  OA22X1 U1507 ( .A0(\i_MIPS/Register/register[6][24] ), .A1(n4938), .B0(
        \i_MIPS/Register/register[14][24] ), .B1(n4932), .Y(n8975) );
  OAI221XL U1508 ( .A0(\i_MIPS/Register/register[18][24] ), .A1(n4944), .B0(
        \i_MIPS/Register/register[26][24] ), .B1(n4939), .C0(n8984), .Y(n8992)
         );
  OA22X1 U1509 ( .A0(\i_MIPS/Register/register[22][24] ), .A1(n4938), .B0(
        \i_MIPS/Register/register[30][24] ), .B1(n4932), .Y(n8984) );
  OA22X1 U1510 ( .A0(\i_MIPS/Register/register[6][30] ), .A1(n4938), .B0(
        \i_MIPS/Register/register[14][30] ), .B1(n4932), .Y(n9297) );
  BUFX4 U1511 ( .A(n4924), .Y(n4926) );
  NAND2X1 U1512 ( .A(n7475), .B(n4707), .Y(n8275) );
  AO22X1 U1513 ( .A0(n4898), .A1(n431), .B0(n4894), .B1(n1994), .Y(n9120) );
  AO22X1 U1514 ( .A0(n4896), .A1(n430), .B0(n4894), .B1(n1993), .Y(n9107) );
  AO22X1 U1515 ( .A0(n4991), .A1(n342), .B0(n4981), .B1(n1923), .Y(n7170) );
  AO22X1 U1516 ( .A0(n4972), .A1(n233), .B0(n4965), .B1(n1918), .Y(n7172) );
  CLKMX2X2 U1517 ( .A(n9280), .B(n9279), .S0(n7972), .Y(n7973) );
  OAI221XL U1518 ( .A0(\i_MIPS/Register/register[18][28] ), .A1(n4921), .B0(
        \i_MIPS/Register/register[26][28] ), .B1(n4917), .C0(n9037), .Y(n9040)
         );
  NOR2BX1 U1519 ( .AN(n4809), .B(\i_MIPS/n371 ), .Y(n4684) );
  INVX6 U1520 ( .A(n4807), .Y(n4806) );
  INVX3 U1521 ( .A(n3892), .Y(n7272) );
  NAND2X4 U1522 ( .A(\i_MIPS/ALUin1[4] ), .B(n3790), .Y(n7354) );
  AO22X1 U1523 ( .A0(n4896), .A1(n436), .B0(n4892), .B1(n1999), .Y(n6984) );
  OAI221XL U1524 ( .A0(\i_MIPS/Register/register[2][14] ), .A1(n4920), .B0(
        \i_MIPS/Register/register[10][14] ), .B1(n4916), .C0(n6982), .Y(n6985)
         );
  NAND3X4 U1525 ( .A(n4150), .B(n4151), .C(n7789), .Y(n7969) );
  NAND2X6 U1526 ( .A(n4707), .B(n7974), .Y(n4151) );
  NAND2X2 U1527 ( .A(n7460), .B(n7459), .Y(n7548) );
  NAND2X4 U1528 ( .A(n3823), .B(\i_MIPS/n365 ), .Y(n7546) );
  NAND2X1 U1529 ( .A(n4827), .B(\i_MIPS/n358 ), .Y(n8141) );
  NAND2X4 U1530 ( .A(net99814), .B(net99815), .Y(n4112) );
  CLKINVX1 U1531 ( .A(n10375), .Y(n10486) );
  OAI221XL U1532 ( .A0(\i_MIPS/Register/register[18][29] ), .A1(n4920), .B0(
        \i_MIPS/Register/register[26][29] ), .B1(n4915), .C0(n6737), .Y(n6740)
         );
  OAI221XL U1533 ( .A0(\i_MIPS/Register/register[2][29] ), .A1(n4920), .B0(
        \i_MIPS/Register/register[10][29] ), .B1(n4915), .C0(n6728), .Y(n6731)
         );
  NAND4X1 U1534 ( .A(n8939), .B(n8938), .C(n8937), .D(n8936), .Y(n8944) );
  CLKINVX1 U1535 ( .A(n8800), .Y(n8801) );
  INVX4 U1536 ( .A(n11104), .Y(n10935) );
  NAND2X2 U1537 ( .A(n4686), .B(n4652), .Y(n6514) );
  NAND2X2 U1538 ( .A(n6591), .B(\i_MIPS/n346 ), .Y(n8431) );
  NAND2X1 U1539 ( .A(\i_MIPS/ALUin1[26] ), .B(n6594), .Y(n8346) );
  CLKMX2X2 U1540 ( .A(n9280), .B(n9279), .S0(n8352), .Y(n8353) );
  CLKMX2X2 U1541 ( .A(n9280), .B(n9279), .S0(n9163), .Y(n8999) );
  BUFX6 U1542 ( .A(n4451), .Y(n5275) );
  INVX6 U1543 ( .A(n3693), .Y(n3676) );
  BUFX8 U1544 ( .A(n11137), .Y(n5189) );
  BUFX4 U1545 ( .A(net134103), .Y(net112385) );
  BUFX4 U1546 ( .A(net112705), .Y(net112693) );
  NAND3BX2 U1547 ( .AN(n3671), .B(n3752), .C(net113533), .Y(net100082) );
  AO22X1 U1548 ( .A0(n4977), .A1(n345), .B0(n4976), .B1(n1926), .Y(n6689) );
  AO22X1 U1549 ( .A0(n4991), .A1(n336), .B0(n4984), .B1(n1913), .Y(n6688) );
  AO22X1 U1550 ( .A0(n4971), .A1(n325), .B0(n4965), .B1(n1901), .Y(n6690) );
  AO22X1 U1551 ( .A0(n4977), .A1(n351), .B0(n4976), .B1(n1933), .Y(n6698) );
  AO22X1 U1552 ( .A0(n4991), .A1(n337), .B0(n4984), .B1(n1914), .Y(n6697) );
  AO22X1 U1553 ( .A0(n4971), .A1(n231), .B0(n4965), .B1(n1902), .Y(n6699) );
  OA22X1 U1554 ( .A0(\i_MIPS/Register/register[22][26] ), .A1(n4934), .B0(
        \i_MIPS/Register/register[30][26] ), .B1(n4931), .Y(n8412) );
  OA22X1 U1555 ( .A0(\i_MIPS/Register/register[6][26] ), .A1(n4938), .B0(
        \i_MIPS/Register/register[14][26] ), .B1(n4931), .Y(n8403) );
  NOR4X1 U1556 ( .A(n8407), .B(n8406), .C(n8405), .D(n8404), .Y(n8408) );
  OA22X1 U1557 ( .A0(\i_MIPS/Register/register[22][28] ), .A1(n4938), .B0(
        \i_MIPS/Register/register[30][28] ), .B1(n4932), .Y(n9071) );
  OA22X1 U1558 ( .A0(\i_MIPS/Register/register[6][28] ), .A1(n4938), .B0(
        \i_MIPS/Register/register[14][28] ), .B1(n4932), .Y(n9062) );
  BUFX4 U1559 ( .A(n5407), .Y(n5404) );
  BUFX6 U1560 ( .A(n5451), .Y(n5449) );
  CLKBUFX3 U1561 ( .A(n5231), .Y(n5225) );
  CLKINVX1 U1562 ( .A(n11220), .Y(n11222) );
  AND2X2 U1563 ( .A(n11220), .B(n9256), .Y(n4591) );
  NAND2X2 U1564 ( .A(\i_MIPS/ALUin1[25] ), .B(n6586), .Y(n8432) );
  NOR2BX2 U1565 ( .AN(n4813), .B(\i_MIPS/n369 ), .Y(n4674) );
  NAND2X6 U1566 ( .A(n11065), .B(n11063), .Y(n10206) );
  INVX3 U1567 ( .A(n10308), .Y(n10309) );
  OAI2BB1X2 U1568 ( .A0N(net98564), .A1N(n10944), .B0(n10934), .Y(n11010) );
  BUFX6 U1569 ( .A(n11181), .Y(n4728) );
  AOI222XL U1570 ( .A0(n4800), .A1(n9181), .B0(n4799), .B1(n9145), .C0(n9144), 
        .C1(n3636), .Y(n9146) );
  INVX4 U1571 ( .A(n7365), .Y(n9010) );
  INVX3 U1572 ( .A(n4797), .Y(n7785) );
  NAND2X4 U1573 ( .A(n6586), .B(\i_MIPS/n346 ), .Y(n8426) );
  INVX3 U1574 ( .A(n6590), .Y(n8331) );
  CLKAND2X3 U1575 ( .A(n8920), .B(n8905), .Y(n4516) );
  INVX4 U1576 ( .A(n8280), .Y(n8927) );
  NAND2X1 U1577 ( .A(n6853), .B(n4707), .Y(n8438) );
  CLKMX2X2 U1578 ( .A(n7611), .B(n7279), .S0(n5590), .Y(n6853) );
  INVX1 U1579 ( .A(n10330), .Y(n10331) );
  NAND2X2 U1580 ( .A(n10935), .B(n11105), .Y(n10494) );
  INVX3 U1581 ( .A(n9258), .Y(n3600) );
  CLKINVX1 U1582 ( .A(n8074), .Y(n3555) );
  OAI211X1 U1583 ( .A0(n8073), .A1(n8072), .B0(n8520), .C0(n8071), .Y(n8074)
         );
  INVX12 U1584 ( .A(net102120), .Y(net102346) );
  NAND4X1 U1585 ( .A(net101970), .B(net101971), .C(\i_MIPS/n213 ), .D(
        net101973), .Y(net99933) );
  NAND4X1 U1586 ( .A(n7297), .B(n7296), .C(n7295), .D(n7294), .Y(n7302) );
  OAI221XL U1587 ( .A0(\i_MIPS/Register/register[2][8] ), .A1(n4920), .B0(
        \i_MIPS/Register/register[10][8] ), .B1(n4915), .C0(n6807), .Y(n6810)
         );
  OAI221XL U1588 ( .A0(\i_MIPS/Register/register[18][8] ), .A1(n4920), .B0(
        \i_MIPS/Register/register[26][8] ), .B1(n4915), .C0(n6816), .Y(n6819)
         );
  OAI221XL U1589 ( .A0(\i_MIPS/Register/register[18][9] ), .A1(n4920), .B0(
        \i_MIPS/Register/register[26][9] ), .B1(n4915), .C0(n6899), .Y(n6902)
         );
  OAI221XL U1590 ( .A0(\i_MIPS/Register/register[2][9] ), .A1(n4920), .B0(
        \i_MIPS/Register/register[10][9] ), .B1(n4915), .C0(n6890), .Y(n6893)
         );
  CLKINVX1 U1591 ( .A(\i_MIPS/ID_EX[81] ), .Y(n5592) );
  BUFX2 U1592 ( .A(n5409), .Y(n5395) );
  OR2X4 U1593 ( .A(n11359), .B(n4565), .Y(n11228) );
  INVX3 U1594 ( .A(n9346), .Y(n4565) );
  AOI2BB2X2 U1595 ( .B0(n4680), .B1(\I_cache/cache[4][147] ), .A0N(n5318), 
        .A1N(n3216), .Y(n5968) );
  OA22X2 U1596 ( .A0(net112245), .A1(n2383), .B0(net112161), .B1(n878), .Y(
        n7489) );
  BUFX4 U1597 ( .A(net111947), .Y(net111953) );
  CLKBUFX3 U1598 ( .A(net112085), .Y(net112077) );
  BUFX12 U1599 ( .A(net112587), .Y(net112565) );
  INVX3 U1600 ( .A(n6138), .Y(n10670) );
  OA22X2 U1601 ( .A0(net112041), .A1(n1946), .B0(net111915), .B1(n368), .Y(
        n6137) );
  INVX3 U1602 ( .A(n6136), .Y(n10671) );
  INVX3 U1603 ( .A(n3750), .Y(n3735) );
  INVX3 U1604 ( .A(n6154), .Y(n10668) );
  OAI221X1 U1605 ( .A0(net112231), .A1(n2042), .B0(net112139), .B1(n315), .C0(
        n6153), .Y(n6154) );
  INVX3 U1606 ( .A(n6101), .Y(n10645) );
  OAI221X1 U1607 ( .A0(net112657), .A1(n2050), .B0(net112563), .B1(n709), .C0(
        n6100), .Y(n6101) );
  INVX3 U1608 ( .A(n6163), .Y(n10660) );
  OA22X2 U1609 ( .A0(net112101), .A1(n422), .B0(net111983), .B1(n3262), .Y(
        n6045) );
  INVX3 U1610 ( .A(n6053), .Y(n10630) );
  AND3X4 U1611 ( .A(n3715), .B(n3716), .C(n6051), .Y(n3311) );
  OR2X2 U1612 ( .A(net112593), .B(n1614), .Y(n3716) );
  NOR4X1 U1613 ( .A(n8750), .B(n8749), .C(n8748), .D(n8747), .Y(n8761) );
  NOR4X1 U1614 ( .A(n7909), .B(n7908), .C(n7907), .D(n7906), .Y(n7910) );
  CLKINVX4 U1615 ( .A(net107168), .Y(net99935) );
  AO21X2 U1616 ( .A0(n10185), .A1(n10184), .B0(net113077), .Y(net104564) );
  INVX6 U1617 ( .A(net107011), .Y(net98973) );
  NOR4X1 U1618 ( .A(n7510), .B(n7509), .C(n7508), .D(n7507), .Y(n7521) );
  AO21X2 U1619 ( .A0(net99108), .A1(net99109), .B0(net113077), .Y(net99090) );
  NAND3BX1 U1620 ( .AN(\i_MIPS/ID_EX[83] ), .B(n8149), .C(n8148), .Y(n8165) );
  CLKINVX1 U1621 ( .A(n8163), .Y(n8147) );
  CLKINVX1 U1622 ( .A(n8158), .Y(n8154) );
  NAND2X4 U1623 ( .A(n6244), .B(\i_MIPS/n361 ), .Y(n7187) );
  NAND2X6 U1624 ( .A(\i_MIPS/ALUin1[10] ), .B(n4320), .Y(n7186) );
  AND2X2 U1625 ( .A(n7200), .B(n4593), .Y(n3578) );
  NAND2X1 U1626 ( .A(n9271), .B(n9270), .Y(n9290) );
  OAI222X1 U1627 ( .A0(n8724), .A1(n8660), .B0(n8659), .B1(n9169), .C0(n8658), 
        .C1(n8657), .Y(n8663) );
  CLKINVX1 U1628 ( .A(n3816), .Y(n8657) );
  INVX6 U1629 ( .A(n8537), .Y(n9139) );
  CLKMX2X2 U1630 ( .A(n9141), .B(n4799), .S0(n9166), .Y(n8652) );
  INVX3 U1631 ( .A(n9007), .Y(n9267) );
  CLKMX2X2 U1632 ( .A(n9141), .B(n4799), .S0(n3704), .Y(n7112) );
  AO22X1 U1633 ( .A0(n7464), .A1(n9259), .B0(n9258), .B1(n7465), .Y(n7470) );
  NAND4BX1 U1634 ( .AN(n7341), .B(n7340), .C(n7339), .D(n7338), .Y(n7352) );
  NOR4X1 U1635 ( .A(n7337), .B(n7336), .C(n7335), .D(n7334), .Y(n7338) );
  NAND4BX1 U1636 ( .AN(n7350), .B(n7349), .C(n7348), .D(n7347), .Y(n7351) );
  OA22X1 U1637 ( .A0(\i_MIPS/Register/register[22][25] ), .A1(n4938), .B0(
        \i_MIPS/Register/register[30][25] ), .B1(n4931), .Y(n8503) );
  OA22X1 U1638 ( .A0(\i_MIPS/Register/register[6][25] ), .A1(n4934), .B0(
        \i_MIPS/Register/register[14][25] ), .B1(n4931), .Y(n8494) );
  AOI32X1 U1639 ( .A0(n8261), .A1(n8260), .A2(n4577), .B0(n8259), .B1(n3636), 
        .Y(n8270) );
  NAND2X1 U1640 ( .A(n8263), .B(n8262), .Y(n8269) );
  BUFX6 U1641 ( .A(n4924), .Y(n4927) );
  CLKMX2X2 U1642 ( .A(n9141), .B(n4799), .S0(n3529), .Y(n7368) );
  OAI221X1 U1643 ( .A0(n4798), .A1(n7357), .B0(n7358), .B1(n9262), .C0(n8805), 
        .Y(n7362) );
  OAI221X1 U1644 ( .A0(\i_MIPS/ALUin1[11] ), .A1(n4825), .B0(
        \i_MIPS/ALUin1[10] ), .B1(n4817), .C0(n6430), .Y(n7353) );
  AO22X1 U1645 ( .A0(net113457), .A1(n11442), .B0(net113463), .B1(n11411), .Y(
        n8026) );
  CLKMX2X2 U1646 ( .A(n4799), .B(n9141), .S0(n7562), .Y(n7563) );
  OAI221X1 U1647 ( .A0(n4798), .A1(n7548), .B0(n7549), .B1(n9262), .C0(n8805), 
        .Y(n7553) );
  CLKINVX1 U1648 ( .A(n10276), .Y(n10278) );
  AND2X2 U1649 ( .A(net111405), .B(n10969), .Y(n4610) );
  CLKINVX4 U1650 ( .A(net103795), .Y(net99363) );
  NOR4X1 U1651 ( .A(n8246), .B(n8245), .C(n8244), .D(n8243), .Y(n8247) );
  CLKXOR2X2 U1652 ( .A(n10363), .B(net111405), .Y(n10348) );
  NAND3X2 U1653 ( .A(ICACHE_addr[26]), .B(ICACHE_addr[25]), .C(n10486), .Y(
        n10697) );
  INVX8 U1654 ( .A(net98436), .Y(net110259) );
  CLKMX2X2 U1655 ( .A(n7430), .B(n7429), .S0(net108963), .Y(net105284) );
  NAND4BX1 U1656 ( .AN(n7428), .B(n7427), .C(n7426), .D(n7425), .Y(n7429) );
  NOR4X1 U1657 ( .A(n7686), .B(n7685), .C(n7684), .D(n7683), .Y(n7687) );
  OAI221XL U1658 ( .A0(\i_MIPS/Register/register[2][17] ), .A1(n4946), .B0(
        \i_MIPS/Register/register[10][17] ), .B1(n4484), .C0(n7673), .Y(n7681)
         );
  MXI2X1 U1659 ( .A(n8846), .B(n8845), .S0(n5587), .Y(n3594) );
  NAND2X2 U1660 ( .A(net140444), .B(net140445), .Y(net100866) );
  INVX6 U1661 ( .A(n10294), .Y(n9366) );
  MXI2X1 U1662 ( .A(n8190), .B(n8189), .S0(n5587), .Y(n3554) );
  NOR4X1 U1663 ( .A(n8179), .B(n8178), .C(n8177), .D(n8176), .Y(n8190) );
  INVX3 U1664 ( .A(n8359), .Y(n8340) );
  NAND2X1 U1665 ( .A(net102300), .B(net106801), .Y(net98965) );
  CLKMX2X2 U1666 ( .A(n6564), .B(n6563), .S0(\i_MIPS/IR_ID[25] ), .Y(net106801) );
  CLKMX2X4 U1667 ( .A(\i_MIPS/n313 ), .B(n4712), .S0(\i_MIPS/ID_EX_5 ), .Y(
        n6292) );
  CLKMX2X4 U1668 ( .A(\i_MIPS/n319 ), .B(n4713), .S0(\i_MIPS/ID_EX_5 ), .Y(
        n6291) );
  NOR4X1 U1669 ( .A(n8381), .B(n8380), .C(n8379), .D(n8378), .Y(n8382) );
  OAI2BB1X2 U1670 ( .A0N(n10409), .A1N(n10408), .B0(net113083), .Y(net99712)
         );
  NAND4X4 U1671 ( .A(n4467), .B(n5983), .C(n5982), .D(n5981), .Y(n11372) );
  OA22X2 U1672 ( .A0(n5162), .A1(n420), .B0(n5119), .B1(n3219), .Y(n4467) );
  INVX3 U1673 ( .A(n6019), .Y(n4446) );
  NAND4X6 U1674 ( .A(n5964), .B(n5963), .C(n5962), .D(n5961), .Y(n11364) );
  OA22X2 U1675 ( .A0(n5157), .A1(n3228), .B0(n5119), .B1(n399), .Y(n5964) );
  OA22X2 U1676 ( .A0(n5164), .A1(n2336), .B0(n5123), .B1(n800), .Y(n4491) );
  OA22X2 U1677 ( .A0(n5250), .A1(n2338), .B0(n5205), .B1(n802), .Y(n9331) );
  BUFX2 U1678 ( .A(n5406), .Y(n5377) );
  CLKBUFX3 U1679 ( .A(n5275), .Y(n5245) );
  BUFX4 U1680 ( .A(n5318), .Y(n5286) );
  CLKBUFX3 U1681 ( .A(n5143), .Y(n5112) );
  NAND4X2 U1682 ( .A(n10135), .B(n10134), .C(n4489), .D(n4490), .Y(n4488) );
  OA22X1 U1683 ( .A0(net112241), .A1(n2337), .B0(net112159), .B1(n801), .Y(
        n4489) );
  OA22X1 U1684 ( .A0(net112673), .A1(n3239), .B0(net112571), .B1(n1610), .Y(
        n10135) );
  OA22X2 U1685 ( .A0(net112489), .A1(n2339), .B0(net112353), .B1(n803), .Y(
        n10134) );
  AND2X2 U1686 ( .A(n117), .B(n11168), .Y(n4576) );
  CLKBUFX6 U1687 ( .A(n4576), .Y(n5063) );
  CLKBUFX3 U1688 ( .A(n10681), .Y(n5061) );
  CLKBUFX6 U1689 ( .A(n4576), .Y(n5062) );
  NAND4X1 U1690 ( .A(n8392), .B(n8391), .C(n8390), .D(n8389), .Y(n11415) );
  OA22X1 U1691 ( .A0(net112667), .A1(n2407), .B0(net112565), .B1(n901), .Y(
        n8392) );
  OA22X1 U1692 ( .A0(net112071), .A1(n2440), .B0(net111947), .B1(n464), .Y(
        n8389) );
  OA22X1 U1693 ( .A0(net112235), .A1(n2443), .B0(net112153), .B1(n468), .Y(
        n8390) );
  NAND4X2 U1694 ( .A(n8109), .B(n8108), .C(n8107), .D(n8106), .Y(n11410) );
  OA22X1 U1695 ( .A0(net112233), .A1(n2413), .B0(net112151), .B1(n384), .Y(
        n8107) );
  NAND4X2 U1696 ( .A(n7919), .B(n7918), .C(n7917), .D(n7916), .Y(n11407) );
  OA22X1 U1697 ( .A0(net112663), .A1(n960), .B0(net112561), .B1(n2485), .Y(
        n7919) );
  OA22X1 U1698 ( .A0(net112493), .A1(n2447), .B0(net112351), .B1(n472), .Y(
        n7918) );
  NAND4X1 U1699 ( .A(n7058), .B(n7057), .C(n7056), .D(n7055), .Y(n11404) );
  OA22X1 U1700 ( .A0(net112673), .A1(n2371), .B0(net112575), .B1(n867), .Y(
        n7058) );
  NAND4X1 U1701 ( .A(n7148), .B(n7147), .C(n7146), .D(n7145), .Y(n11400) );
  OA22X1 U1702 ( .A0(net112051), .A1(n2445), .B0(net111927), .B1(n470), .Y(
        n7145) );
  OA22X1 U1703 ( .A0(net112665), .A1(n934), .B0(net112575), .B1(n2459), .Y(
        n7148) );
  NAND4X1 U1704 ( .A(n6272), .B(n6271), .C(n6270), .D(n6269), .Y(n11432) );
  OA22X1 U1705 ( .A0(net112237), .A1(n2366), .B0(net112153), .B1(n863), .Y(
        n6270) );
  OA22X1 U1706 ( .A0(net112673), .A1(n459), .B0(net112571), .B1(n2013), .Y(
        n9244) );
  OA22X1 U1707 ( .A0(net112241), .A1(n462), .B0(net112159), .B1(n2016), .Y(
        n9242) );
  OA22X1 U1708 ( .A0(net112083), .A1(n460), .B0(net111959), .B1(n2014), .Y(
        n9241) );
  OA22X1 U1709 ( .A0(net112667), .A1(n2406), .B0(net112565), .B1(n900), .Y(
        n8396) );
  NAND4X2 U1710 ( .A(n7923), .B(n7922), .C(n7921), .D(n7920), .Y(n11469) );
  NAND4X1 U1711 ( .A(n6879), .B(n6878), .C(n6877), .D(n6876), .Y(n11460) );
  NAND4X2 U1712 ( .A(n7326), .B(n7325), .C(n7324), .D(n7323), .Y(n11457) );
  OA22X1 U1713 ( .A0(net112239), .A1(n2387), .B0(net112161), .B1(n882), .Y(
        n7324) );
  NAND4X1 U1714 ( .A(n7404), .B(n7403), .C(n7402), .D(n7401), .Y(n11456) );
  OA22X1 U1715 ( .A0(net112239), .A1(n2388), .B0(net112161), .B1(n883), .Y(
        n7402) );
  OA22X1 U1716 ( .A0(net112665), .A1(n966), .B0(net112565), .B1(n2491), .Y(
        n8597) );
  OA22X1 U1717 ( .A0(net112485), .A1(n965), .B0(net112361), .B1(n2490), .Y(
        n8596) );
  OA22X1 U1718 ( .A0(net112663), .A1(n957), .B0(net112561), .B1(n2482), .Y(
        n7822) );
  OA22X1 U1719 ( .A0(net112063), .A1(n937), .B0(net111939), .B1(n2462), .Y(
        n7819) );
  NAND4X2 U1720 ( .A(n7733), .B(n7732), .C(n7731), .D(n7730), .Y(n11499) );
  NAND4X1 U1721 ( .A(n6284), .B(n6283), .C(n6282), .D(n6281), .Y(n11494) );
  OA22X1 U1722 ( .A0(net112245), .A1(n2364), .B0(net112155), .B1(n861), .Y(
        n6282) );
  OA22X1 U1723 ( .A0(net112673), .A1(n2374), .B0(net112575), .B1(n870), .Y(
        n7156) );
  OA22X2 U1724 ( .A0(net112245), .A1(n2391), .B0(net112161), .B1(n886), .Y(
        n7154) );
  BUFX4 U1725 ( .A(net112143), .Y(net112147) );
  BUFX4 U1726 ( .A(net111961), .Y(net111941) );
  BUFX4 U1727 ( .A(net112509), .Y(net112429) );
  BUFX4 U1728 ( .A(net99406), .Y(net114113) );
  AO22X2 U1729 ( .A0(net113445), .A1(n11467), .B0(net102346), .B1(n11498), .Y(
        n8207) );
  AO22X2 U1730 ( .A0(net113457), .A1(n11436), .B0(net113463), .B1(n11405), .Y(
        n8208) );
  NAND2X1 U1731 ( .A(n12954), .B(net113089), .Y(n10448) );
  AO22X1 U1732 ( .A0(net113457), .A1(net98153), .B0(net113463), .B1(net98185), 
        .Y(net105006) );
  OA22X1 U1733 ( .A0(\i_MIPS/Register/register[22][31] ), .A1(n4938), .B0(
        \i_MIPS/Register/register[30][31] ), .B1(n4932), .Y(n9199) );
  OA22X1 U1734 ( .A0(\i_MIPS/Register/register[6][31] ), .A1(n4938), .B0(
        \i_MIPS/Register/register[14][31] ), .B1(n4932), .Y(n9190) );
  NOR3X1 U1735 ( .A(\i_MIPS/Reg_W[0] ), .B(\i_MIPS/Reg_W[2] ), .C(n229), .Y(
        \i_MIPS/Register/n115 ) );
  NOR3X1 U1736 ( .A(\i_MIPS/Reg_W[1] ), .B(\i_MIPS/Reg_W[2] ), .C(n287), .Y(
        \i_MIPS/Register/n117 ) );
  NOR3X1 U1737 ( .A(n287), .B(\i_MIPS/Reg_W[2] ), .C(n229), .Y(
        \i_MIPS/Register/n113 ) );
  NOR3X1 U1738 ( .A(n287), .B(\i_MIPS/Reg_W[1] ), .C(n4705), .Y(
        \i_MIPS/Register/n109 ) );
  NOR3X1 U1739 ( .A(n229), .B(\i_MIPS/Reg_W[0] ), .C(n4705), .Y(
        \i_MIPS/Register/n107 ) );
  BUFX2 U1740 ( .A(n5274), .Y(n5247) );
  CLKBUFX3 U1741 ( .A(n5187), .Y(n5156) );
  BUFX6 U1742 ( .A(n5471), .Y(n5469) );
  CLKINVX8 U1743 ( .A(n3685), .Y(n3686) );
  INVX4 U1744 ( .A(n6448), .Y(n3685) );
  CLKINVX1 U1745 ( .A(n8902), .Y(n6629) );
  CLKINVX1 U1746 ( .A(n8334), .Y(n6650) );
  NAND2X4 U1747 ( .A(n3530), .B(n282), .Y(n6447) );
  AOI211X1 U1748 ( .A0(n6491), .A1(n8068), .B0(n6490), .C0(n7961), .Y(n6493)
         );
  AO22X1 U1749 ( .A0(n7621), .A1(n9259), .B0(n286), .B1(n9258), .Y(n7624) );
  MXI2X2 U1750 ( .A(n7269), .B(n6856), .S0(n5590), .Y(n4598) );
  CLKINVX1 U1751 ( .A(n6855), .Y(n6856) );
  NOR3X1 U1752 ( .A(\i_MIPS/Reg_W[1] ), .B(\i_MIPS/Reg_W[2] ), .C(
        \i_MIPS/Reg_W[0] ), .Y(\i_MIPS/Register/n119 ) );
  NOR3X1 U1753 ( .A(\i_MIPS/Reg_W[0] ), .B(\i_MIPS/Reg_W[1] ), .C(n4705), .Y(
        \i_MIPS/Register/n111 ) );
  CLKAND2X3 U1754 ( .A(net98564), .B(n11151), .Y(n4609) );
  CLKINVX1 U1755 ( .A(n11049), .Y(n11062) );
  NAND2X2 U1756 ( .A(n10905), .B(n10906), .Y(n11107) );
  NAND2X4 U1757 ( .A(n10917), .B(n10907), .Y(n11105) );
  NAND2X2 U1758 ( .A(ICACHE_addr[1]), .B(ICACHE_addr[0]), .Y(n9607) );
  XOR2X4 U1759 ( .A(net102183), .B(n3861), .Y(n3731) );
  INVX1 U1760 ( .A(n7364), .Y(n8538) );
  NAND2X1 U1761 ( .A(n6254), .B(n6253), .Y(n3596) );
  CLKMX2X2 U1762 ( .A(n6431), .B(n6765), .S0(n5589), .Y(n7366) );
  CLKMX2X2 U1763 ( .A(n4799), .B(n9141), .S0(n6602), .Y(n6264) );
  INVX3 U1764 ( .A(n8449), .Y(n8450) );
  NAND3X4 U1765 ( .A(ICACHE_addr[24]), .B(ICACHE_addr[23]), .C(n10361), .Y(
        n10375) );
  INVX6 U1766 ( .A(n10291), .Y(n10198) );
  CLKAND2X3 U1767 ( .A(net98564), .B(n11029), .Y(n4608) );
  CLKINVX4 U1768 ( .A(net104271), .Y(net99386) );
  NAND2BX2 U1769 ( .AN(n10951), .B(n10950), .Y(n11024) );
  INVX8 U1770 ( .A(n10290), .Y(n9364) );
  INVX8 U1771 ( .A(n10204), .Y(n10202) );
  NOR4X1 U1772 ( .A(n7381), .B(n7380), .C(n7379), .D(n7378), .Y(n7392) );
  AO21X2 U1773 ( .A0(net100048), .A1(net100049), .B0(net113077), .Y(net100042)
         );
  AO21X2 U1774 ( .A0(net99977), .A1(net99978), .B0(net113077), .Y(net99974) );
  CLKBUFX3 U1775 ( .A(n5592), .Y(n5591) );
  NAND4X1 U1776 ( .A(n9360), .B(n9359), .C(n9358), .D(n9357), .Y(n11231) );
  NAND4X1 U1777 ( .A(n9462), .B(n9461), .C(n9460), .D(n9459), .Y(n11234) );
  NAND4X1 U1778 ( .A(n9440), .B(n9439), .C(n9438), .D(n9437), .Y(n11236) );
  NAND4X2 U1779 ( .A(n9829), .B(n9828), .C(n9827), .D(n9826), .Y(n11237) );
  NAND4X1 U1780 ( .A(n9425), .B(n9424), .C(n9423), .D(n9422), .Y(n11238) );
  NAND4X1 U1781 ( .A(n9963), .B(n9962), .C(n9961), .D(n9960), .Y(n11241) );
  OA22X1 U1782 ( .A0(n5444), .A1(n910), .B0(n5398), .B1(n2427), .Y(n10091) );
  NAND4X1 U1783 ( .A(n9381), .B(n9380), .C(n9379), .D(n9378), .Y(n11243) );
  NAND4X1 U1784 ( .A(n9526), .B(n9525), .C(n9524), .D(n9523), .Y(n11265) );
  OA22X1 U1785 ( .A0(n5254), .A1(n442), .B0(n5208), .B1(n2004), .Y(n9471) );
  OA22X1 U1786 ( .A0(n5253), .A1(n2424), .B0(n5207), .B1(n447), .Y(n9449) );
  OAI22XL U1787 ( .A0(n5167), .A1(n906), .B0(n5123), .B1(n2417), .Y(n4475) );
  OA22X1 U1788 ( .A0(n5432), .A1(n2423), .B0(n5388), .B1(n446), .Y(n9447) );
  OA22X1 U1789 ( .A0(n5262), .A1(n909), .B0(n5216), .B1(n2426), .Y(n9818) );
  OA22X1 U1790 ( .A0(n5252), .A1(n917), .B0(n5206), .B1(n2434), .Y(n9415) );
  OA22X1 U1791 ( .A0(n5431), .A1(n2422), .B0(n5387), .B1(n445), .Y(n9413) );
  OA22X1 U1792 ( .A0(n5165), .A1(n913), .B0(n5121), .B1(n2430), .Y(n9386) );
  OA22X1 U1793 ( .A0(n5251), .A1(n914), .B0(n5205), .B1(n2431), .Y(n9385) );
  NAND4X1 U1794 ( .A(n9531), .B(n9530), .C(n9529), .D(n9528), .Y(n11299) );
  NAND4X1 U1795 ( .A(n9445), .B(n9444), .C(n9443), .D(n9442), .Y(n11300) );
  NAND4X1 U1796 ( .A(n9411), .B(n9410), .C(n9409), .D(n9408), .Y(n11302) );
  NAND4X1 U1797 ( .A(n10089), .B(n10088), .C(n10087), .D(n10086), .Y(n11306)
         );
  NAND4X1 U1798 ( .A(n9355), .B(n9354), .C(n9353), .D(n9352), .Y(n11327) );
  NAND4X1 U1799 ( .A(n9457), .B(n9456), .C(n9455), .D(n9454), .Y(n11330) );
  OA22X1 U1800 ( .A0(n5256), .A1(n2421), .B0(n5210), .B1(n444), .Y(n9540) );
  OAI22XL U1801 ( .A0(n5170), .A1(n438), .B0(n5126), .B1(n2001), .Y(n4486) );
  NAND4X1 U1802 ( .A(n9435), .B(n9434), .C(n9433), .D(n9432), .Y(n11332) );
  NAND4X1 U1803 ( .A(n9420), .B(n9419), .C(n9418), .D(n9417), .Y(n11334) );
  OA22X2 U1804 ( .A0(n5333), .A1(n3220), .B0(n5290), .B1(n356), .Y(n6004) );
  OA22X2 U1805 ( .A0(n5163), .A1(n3225), .B0(n5120), .B1(n1586), .Y(n6006) );
  NAND4X4 U1806 ( .A(n6002), .B(n6001), .C(n6000), .D(n5999), .Y(n11366) );
  OA22X2 U1807 ( .A0(n5332), .A1(n3280), .B0(n5289), .B1(n1624), .Y(n6000) );
  OA22X2 U1808 ( .A0(n5162), .A1(n1976), .B0(n5119), .B1(n409), .Y(n6002) );
  OA22X2 U1809 ( .A0(n3611), .A1(n1978), .B0(n5383), .B1(n411), .Y(n5999) );
  NAND4X4 U1810 ( .A(n5998), .B(n5997), .C(n5996), .D(n5995), .Y(n11367) );
  OA22X2 U1811 ( .A0(n5248), .A1(n1962), .B0(n5203), .B1(n390), .Y(n5997) );
  OA22X2 U1812 ( .A0(n5332), .A1(n1600), .B0(n5289), .B1(n3260), .Y(n5986) );
  OA22X2 U1813 ( .A0(n5162), .A1(n3223), .B0(n5119), .B1(n1584), .Y(n4465) );
  OA22X2 U1814 ( .A0(n3611), .A1(n3237), .B0(n5383), .B1(n1599), .Y(n5985) );
  NAND4X4 U1815 ( .A(n5994), .B(n5993), .C(n5992), .D(n5991), .Y(n11378) );
  OA22X2 U1816 ( .A0(n5332), .A1(n4497), .B0(n5289), .B1(n3205), .Y(n5992) );
  OA22X2 U1817 ( .A0(n3611), .A1(n1627), .B0(n5383), .B1(n3309), .Y(n5991) );
  NAND4X4 U1818 ( .A(n5990), .B(n5989), .C(n5988), .D(n5987), .Y(n11379) );
  OA22X2 U1819 ( .A0(n5332), .A1(n3277), .B0(n5289), .B1(n1621), .Y(n5988) );
  NAND4X4 U1820 ( .A(n6014), .B(n6013), .C(n6012), .D(n6011), .Y(n11381) );
  NAND4X4 U1821 ( .A(n6018), .B(n6017), .C(n6016), .D(n6015), .Y(n11382) );
  NAND4X4 U1822 ( .A(n5976), .B(n5975), .C(n5974), .D(n5973), .Y(n11385) );
  AOI2BB2X2 U1823 ( .B0(n4698), .B1(\I_cache/cache[4][149] ), .A0N(n5317), 
        .A1N(n3217), .Y(n5974) );
  NAND4X2 U1824 ( .A(n7640), .B(n7639), .C(n7638), .D(n7637), .Y(n11391) );
  OA22X1 U1825 ( .A0(net112673), .A1(n925), .B0(net112571), .B1(n2448), .Y(
        n7640) );
  OA22X1 U1826 ( .A0(net112059), .A1(n926), .B0(net111935), .B1(n2449), .Y(
        n7637) );
  OA22X1 U1827 ( .A0(net112239), .A1(n2381), .B0(net112161), .B1(n374), .Y(
        n7398) );
  NAND4X2 U1828 ( .A(n7322), .B(n7321), .C(n7320), .D(n7319), .Y(n11395) );
  OA22X2 U1829 ( .A0(net112239), .A1(n2379), .B0(net112161), .B1(n875), .Y(
        n7320) );
  OA22X1 U1830 ( .A0(net112245), .A1(n2360), .B0(net112153), .B1(n857), .Y(
        n6274) );
  OA22X1 U1831 ( .A0(net112245), .A1(n2361), .B0(net112153), .B1(n858), .Y(
        n6382) );
  CLKINVX1 U1832 ( .A(n11404), .Y(n10192) );
  OA22X1 U1833 ( .A0(net112663), .A1(n959), .B0(net112561), .B1(n2484), .Y(
        n7814) );
  OA22X1 U1834 ( .A0(net112459), .A1(n958), .B0(net112351), .B1(n2483), .Y(
        n7813) );
  NAND4X2 U1835 ( .A(n9051), .B(n9050), .C(n9049), .D(n9048), .Y(n11417) );
  OA22X1 U1836 ( .A0(net112245), .A1(n2365), .B0(net112153), .B1(n862), .Y(
        n6528) );
  NAND4X2 U1837 ( .A(n7721), .B(n7720), .C(n7719), .D(n7718), .Y(n11437) );
  OA22X1 U1838 ( .A0(net112473), .A1(n951), .B0(net112349), .B1(n2476), .Y(
        n7720) );
  OA22X1 U1839 ( .A0(net112679), .A1(n2378), .B0(net112575), .B1(n874), .Y(
        n6971) );
  OA22X1 U1840 ( .A0(net112245), .A1(n2394), .B0(net112161), .B1(n889), .Y(
        n6969) );
  OA22X1 U1841 ( .A0(net112665), .A1(n2372), .B0(net112575), .B1(n868), .Y(
        n7062) );
  OA22X2 U1842 ( .A0(net112245), .A1(n2390), .B0(net112163), .B1(n885), .Y(
        n7060) );
  NAND4X2 U1843 ( .A(n8593), .B(n8592), .C(n8591), .D(n8590), .Y(n11471) );
  NAND4X2 U1844 ( .A(n8113), .B(n8112), .C(n8111), .D(n8110), .Y(n11472) );
  NAND4X2 U1845 ( .A(n8299), .B(n8298), .C(n8297), .D(n8296), .Y(n11474) );
  NAND4X2 U1846 ( .A(n9055), .B(n9054), .C(n9053), .D(n9052), .Y(n11479) );
  NAND4X2 U1847 ( .A(n7648), .B(n7647), .C(n7646), .D(n7645), .Y(n11484) );
  OA22X1 U1848 ( .A0(net112473), .A1(n931), .B0(net112349), .B1(n2455), .Y(
        n7647) );
  NAND4X2 U1849 ( .A(n7408), .B(n7407), .C(n7406), .D(n7405), .Y(n11487) );
  OA22X1 U1850 ( .A0(net112057), .A1(n950), .B0(net111933), .B1(n2475), .Y(
        n7405) );
  OA22X1 U1851 ( .A0(net112245), .A1(n2385), .B0(net112161), .B1(n880), .Y(
        n7406) );
  NAND4X2 U1852 ( .A(n7246), .B(n7245), .C(n7244), .D(n7243), .Y(n11492) );
  OA22X2 U1853 ( .A0(net112671), .A1(n2375), .B0(net112575), .B1(n871), .Y(
        n7246) );
  OA22X2 U1854 ( .A0(net112245), .A1(n2392), .B0(net112161), .B1(n887), .Y(
        n7244) );
  NAND4X2 U1855 ( .A(n6392), .B(n6391), .C(n6390), .D(n6389), .Y(n11495) );
  OA22X1 U1856 ( .A0(net112245), .A1(n2362), .B0(net112153), .B1(n859), .Y(
        n6390) );
  NAND4X2 U1857 ( .A(n8117), .B(n8116), .C(n8115), .D(n8114), .Y(n11503) );
  NAND4X2 U1858 ( .A(n8303), .B(n8302), .C(n8301), .D(n8300), .Y(n11505) );
  OA22X1 U1859 ( .A0(net112235), .A1(n943), .B0(net112153), .B1(n2468), .Y(
        n8301) );
  NAND4X2 U1860 ( .A(n8491), .B(n8490), .C(n8489), .D(n8488), .Y(n11507) );
  OA22X1 U1861 ( .A0(net112667), .A1(n941), .B0(net112565), .B1(n2466), .Y(
        n8491) );
  OA22X1 U1862 ( .A0(net112235), .A1(n940), .B0(net112153), .B1(n2465), .Y(
        n8489) );
  OA22X1 U1863 ( .A0(net112671), .A1(n935), .B0(net112569), .B1(n2460), .Y(
        n9059) );
  NAND4X2 U1864 ( .A(n9098), .B(n9097), .C(n9096), .D(n9095), .Y(n11513) );
  NAND2X1 U1865 ( .A(net113605), .B(n4784), .Y(n11516) );
  NAND3BX1 U1866 ( .AN(n11515), .B(n11548), .C(n11514), .Y(n4784) );
  NAND2X6 U1867 ( .A(n10627), .B(n10626), .Y(n3832) );
  INVX3 U1868 ( .A(n6058), .Y(n10626) );
  NAND2X2 U1869 ( .A(n10642), .B(n10641), .Y(n11536) );
  CLKMX2X2 U1870 ( .A(n8884), .B(n8883), .S0(net108959), .Y(net102744) );
  CLKMX2X2 U1871 ( .A(n7949), .B(n7948), .S0(net108963), .Y(net104351) );
  CLKMX2X2 U1872 ( .A(n6193), .B(n6192), .S0(net108959), .Y(net107236) );
  BUFX4 U1873 ( .A(net99607), .Y(n4029) );
  INVX4 U1874 ( .A(net99609), .Y(net105930) );
  NOR3X6 U1875 ( .A(n3618), .B(n3619), .C(n3620), .Y(n6959) );
  AOI211X1 U1876 ( .A0(n9140), .A1(n8145), .B0(n6781), .C0(n6780), .Y(n6782)
         );
  INVX3 U1877 ( .A(n3834), .Y(net99639) );
  AO21X2 U1878 ( .A0(n10184), .A1(n10185), .B0(net112729), .Y(net104526) );
  CLKMX2X2 U1879 ( .A(n8799), .B(n8798), .S0(net108959), .Y(net102899) );
  OR2X1 U1880 ( .A(net107041), .B(net112709), .Y(n3615) );
  CLKMX2X2 U1881 ( .A(n8325), .B(n8324), .S0(net108959), .Y(net103707) );
  CLKMX2X2 U1882 ( .A(n7450), .B(n7449), .S0(net108963), .Y(net105150) );
  AND3X6 U1883 ( .A(n3793), .B(n3794), .C(n9325), .Y(n3314) );
  OR2X4 U1884 ( .A(n9326), .B(net112709), .Y(n3793) );
  CLKINVX1 U1885 ( .A(n10299), .Y(n10296) );
  CLKINVX1 U1886 ( .A(n10270), .Y(n10274) );
  CLKINVX1 U1887 ( .A(n10871), .Y(n10207) );
  NAND4X1 U1888 ( .A(n9739), .B(n9738), .C(n9737), .D(n9736), .Y(n10249) );
  OR2X2 U1889 ( .A(net105735), .B(net112709), .Y(n3802) );
  INVX4 U1890 ( .A(net99407), .Y(net104184) );
  INVX3 U1891 ( .A(\i_MIPS/n307 ), .Y(n10837) );
  CLKMX2X2 U1892 ( .A(n7609), .B(n7608), .S0(net108963), .Y(net104868) );
  CLKMX2X2 U1893 ( .A(n8046), .B(n8045), .S0(net108959), .Y(net104183) );
  NAND4BX1 U1894 ( .AN(n8044), .B(n8043), .C(n8042), .D(n8041), .Y(n8045) );
  CLKINVX1 U1895 ( .A(n10244), .Y(n10245) );
  CLKINVX1 U1896 ( .A(n10249), .Y(n11040) );
  OR2X4 U1897 ( .A(n11146), .B(net110247), .Y(n3654) );
  AND2X4 U1898 ( .A(n10704), .B(n10717), .Y(n4544) );
  INVX3 U1899 ( .A(net140280), .Y(net140278) );
  INVX3 U1900 ( .A(n10906), .Y(n10930) );
  AND2X2 U1901 ( .A(n3553), .B(net99541), .Y(n4535) );
  INVX6 U1902 ( .A(n3815), .Y(n4434) );
  NAND3X4 U1903 ( .A(n3701), .B(n7291), .C(n7292), .Y(net99461) );
  CLKMX2X4 U1904 ( .A(\i_MIPS/n317 ), .B(n6199), .S0(\i_MIPS/ID_EX_5 ), .Y(
        n10132) );
  CLKINVX1 U1905 ( .A(\i_MIPS/ID_EX[86] ), .Y(n6199) );
  CLKINVX1 U1906 ( .A(n6293), .Y(n10131) );
  INVX1 U1907 ( .A(n6292), .Y(n10133) );
  AO22X2 U1908 ( .A0(n115), .A1(ICACHE_addr[13]), .B0(n5463), .B1(n11372), .Y(
        n10980) );
  CLKINVX1 U1909 ( .A(n10982), .Y(n3509) );
  CLKINVX1 U1910 ( .A(n10975), .Y(n3513) );
  AO22X2 U1911 ( .A0(n115), .A1(ICACHE_addr[15]), .B0(n5463), .B1(n11374), .Y(
        n10989) );
  AO22X2 U1912 ( .A0(n113), .A1(ICACHE_addr[9]), .B0(n5463), .B1(n11368), .Y(
        n10986) );
  CLKINVX1 U1913 ( .A(n10979), .Y(n3511) );
  INVX3 U1914 ( .A(n5318), .Y(n4675) );
  AO22X2 U1915 ( .A0(mem_rdata_I[0]), .A1(n113), .B0(n5465), .B1(n11230), .Y(
        n9507) );
  AO22X2 U1916 ( .A0(mem_rdata_I[37]), .A1(n115), .B0(n5465), .B1(n11267), .Y(
        n9537) );
  AO22X2 U1917 ( .A0(mem_rdata_I[69]), .A1(n114), .B0(n5465), .B1(n11299), .Y(
        n9532) );
  AO22X2 U1918 ( .A0(mem_rdata_I[64]), .A1(n114), .B0(n5465), .B1(n11294), .Y(
        n9502) );
  AO22X2 U1919 ( .A0(mem_rdata_I[111]), .A1(n113), .B0(n5466), .B1(n11341), 
        .Y(n9351) );
  BUFX2 U1920 ( .A(n5406), .Y(n5376) );
  AO22X2 U1921 ( .A0(mem_rdata_I[96]), .A1(n114), .B0(n5465), .B1(n11326), .Y(
        n9497) );
  AOI222X1 U1922 ( .A0(net109795), .A1(n11420), .B0(mem_rdata_D[31]), .B1(n117), .C0(net109805), .C1(n12966), .Y(n11210) );
  CLKBUFX3 U1923 ( .A(n10470), .Y(n4305) );
  AOI222X1 U1924 ( .A0(net109791), .A1(n11416), .B0(mem_rdata_D[27]), .B1(n116), .C0(n12970), .C1(net109801), .Y(n10469) );
  BUFX6 U1925 ( .A(n10603), .Y(n4314) );
  CLKBUFX3 U1926 ( .A(n10457), .Y(n4315) );
  AOI222X1 U1927 ( .A0(net109791), .A1(n11405), .B0(mem_rdata_D[16]), .B1(n117), .C0(n12981), .C1(net109801), .Y(n10456) );
  CLKINVX1 U1928 ( .A(n11403), .Y(n10441) );
  CLKBUFX8 U1929 ( .A(n10773), .Y(n4316) );
  MXI2X1 U1930 ( .A(n10772), .B(n10771), .S0(n5490), .Y(n10773) );
  CLKBUFX3 U1931 ( .A(n10515), .Y(n4317) );
  AOI222X1 U1932 ( .A0(net109791), .A1(n11393), .B0(mem_rdata_D[3]), .B1(n117), 
        .C0(n12994), .C1(net109801), .Y(n10514) );
  AOI222X1 U1933 ( .A0(net109795), .A1(n11392), .B0(mem_rdata_D[2]), .B1(n116), 
        .C0(n12995), .C1(net109805), .Y(n11176) );
  MXI2X2 U1934 ( .A(n10858), .B(n10857), .S0(n5498), .Y(n10859) );
  NOR3X1 U1935 ( .A(n4178), .B(n4179), .C(n4180), .Y(n10858) );
  BUFX4 U1936 ( .A(n11216), .Y(n4245) );
  BUFX4 U1937 ( .A(n10694), .Y(n4283) );
  CLKBUFX3 U1938 ( .A(n10485), .Y(n4284) );
  CLKBUFX3 U1939 ( .A(n10406), .Y(n4285) );
  BUFX4 U1940 ( .A(n10473), .Y(n4286) );
  BUFX4 U1941 ( .A(n10422), .Y(n4287) );
  BUFX4 U1942 ( .A(n10434), .Y(n4288) );
  BUFX4 U1943 ( .A(n10580), .Y(n4289) );
  BUFX4 U1944 ( .A(n10567), .Y(n4290) );
  BUFX4 U1945 ( .A(n10555), .Y(n4291) );
  BUFX4 U1946 ( .A(n10543), .Y(n4292) );
  CLKBUFX3 U1947 ( .A(n10531), .Y(n4293) );
  BUFX4 U1948 ( .A(n10183), .Y(n4294) );
  CLKBUFX3 U1949 ( .A(n10619), .Y(n4295) );
  CLKBUFX3 U1950 ( .A(n10460), .Y(n4296) );
  BUFX4 U1951 ( .A(n10197), .Y(n4297) );
  CLKBUFX3 U1952 ( .A(n10446), .Y(n4298) );
  AOI222X1 U1953 ( .A0(n5486), .A1(n11434), .B0(mem_rdata_D[46]), .B1(n116), 
        .C0(n12983), .C1(n5482), .Y(n10445) );
  CLKBUFX3 U1954 ( .A(n10812), .Y(n4241) );
  BUFX4 U1955 ( .A(n10788), .Y(n4244) );
  CLKBUFX3 U1956 ( .A(n10776), .Y(n4299) );
  BUFX4 U1957 ( .A(n10828), .Y(n4242) );
  BUFX4 U1958 ( .A(n10749), .Y(n4300) );
  CLKBUFX3 U1959 ( .A(n10171), .Y(n4282) );
  AOI222X1 U1960 ( .A0(n5486), .A1(net98153), .B0(mem_rdata_D[38]), .B1(n116), 
        .C0(n12991), .C1(n5482), .Y(n10170) );
  BUFX4 U1961 ( .A(n10763), .Y(n4301) );
  CLKBUFX3 U1962 ( .A(n10164), .Y(n4251) );
  BUFX4 U1963 ( .A(n10518), .Y(n4302) );
  BUFX4 U1964 ( .A(n11180), .Y(n4246) );
  BUFX4 U1965 ( .A(n10849), .Y(n4243) );
  CLKBUFX3 U1966 ( .A(n10479), .Y(n4267) );
  AOI222X1 U1967 ( .A0(n5479), .A1(n11480), .B0(mem_rdata_D[93]), .B1(n116), 
        .C0(n12968), .C1(n5476), .Y(n10478) );
  CLKBUFX3 U1968 ( .A(n10467), .Y(n4268) );
  AOI222X1 U1969 ( .A0(n5479), .A1(n11478), .B0(mem_rdata_D[91]), .B1(n117), 
        .C0(n12970), .C1(n5476), .Y(n10466) );
  INVX3 U1970 ( .A(n3566), .Y(n10549) );
  CLKMX2X2 U1971 ( .A(n10547), .B(n10548), .S0(n3567), .Y(n3566) );
  MXI2X1 U1972 ( .A(n10176), .B(n10175), .S0(n5497), .Y(n10177) );
  INVX8 U1973 ( .A(net111915), .Y(net111873) );
  AOI222X1 U1974 ( .A0(n5480), .A1(n11468), .B0(mem_rdata_D[81]), .B1(n117), 
        .C0(n12980), .C1(n5477), .Y(n10599) );
  BUFX4 U1975 ( .A(n10806), .Y(n4236) );
  MXI2X1 U1976 ( .A(n10805), .B(n10804), .S0(n5489), .Y(n10806) );
  BUFX4 U1977 ( .A(n10782), .Y(n4239) );
  MXI2X1 U1978 ( .A(n10781), .B(n10780), .S0(n5490), .Y(n10782) );
  AOI222X1 U1979 ( .A0(n5480), .A1(n11461), .B0(mem_rdata_D[74]), .B1(n116), 
        .C0(n12987), .C1(n5477), .Y(n10587) );
  BUFX4 U1980 ( .A(n10822), .Y(n4237) );
  MXI2X1 U1981 ( .A(n10821), .B(n10820), .S0(n5489), .Y(n10822) );
  CLKBUFX3 U1982 ( .A(n11174), .Y(n4240) );
  AOI222X1 U1983 ( .A0(n5481), .A1(n11454), .B0(mem_rdata_D[66]), .B1(n116), 
        .C0(n12995), .C1(n5478), .Y(n11173) );
  BUFX4 U1984 ( .A(n10843), .Y(n4238) );
  MXI2X1 U1985 ( .A(n10842), .B(n10841), .S0(n5489), .Y(n10843) );
  AOI222X1 U1986 ( .A0(n5481), .A1(n11452), .B0(mem_rdata_D[64]), .B1(n116), 
        .C0(n12997), .C1(n5478), .Y(n10855) );
  CLKBUFX6 U1987 ( .A(n10685), .Y(n4253) );
  CLKBUFX3 U1988 ( .A(n10464), .Y(n4256) );
  AOI222X1 U1989 ( .A0(n5474), .A1(n11509), .B0(mem_rdata_D[123]), .B1(n116), 
        .C0(n12970), .C1(n5472), .Y(n10463) );
  MXI2X1 U1990 ( .A(n10412), .B(n10411), .S0(n5496), .Y(n10413) );
  BUFX6 U1991 ( .A(n10571), .Y(n4258) );
  AOI222X1 U1992 ( .A0(n5475), .A1(n11506), .B0(mem_rdata_D[120]), .B1(n117), 
        .C0(n12973), .C1(n5473), .Y(n10570) );
  CLKBUFX6 U1993 ( .A(n10546), .Y(n4260) );
  BUFX6 U1994 ( .A(n10610), .Y(n4262) );
  AOI222X1 U1995 ( .A0(n5475), .A1(n11500), .B0(mem_rdata_D[114]), .B1(n117), 
        .C0(n12979), .C1(n5473), .Y(n10609) );
  CLKBUFX3 U1996 ( .A(n10451), .Y(n4263) );
  AOI222X1 U1997 ( .A0(n5474), .A1(n11496), .B0(mem_rdata_D[110]), .B1(n117), 
        .C0(n12983), .C1(n5472), .Y(n10436) );
  AOI222X1 U1998 ( .A0(n5475), .A1(n11491), .B0(mem_rdata_D[105]), .B1(n117), 
        .C0(n12988), .C1(n5473), .Y(n10766) );
  AOI222X1 U1999 ( .A0(n5474), .A1(n11490), .B0(mem_rdata_D[104]), .B1(n117), 
        .C0(n12989), .C1(n5473), .Y(n10818) );
  INVX6 U2000 ( .A(net112143), .Y(net112123) );
  BUFX4 U2001 ( .A(n10740), .Y(n4265) );
  MXI2X1 U2002 ( .A(n10739), .B(n10738), .S0(n5491), .Y(n10740) );
  AOI222X1 U2003 ( .A0(n5474), .A1(n11486), .B0(mem_rdata_D[99]), .B1(n116), 
        .C0(n12994), .C1(n5472), .Y(n10141) );
  MXI2X1 U2004 ( .A(n11170), .B(n11169), .S0(n5492), .Y(n11171) );
  OR2X6 U2005 ( .A(net106564), .B(net112723), .Y(n3690) );
  NAND3X6 U2006 ( .A(n3728), .B(n3729), .C(n8423), .Y(net99624) );
  OR2X4 U2007 ( .A(n8425), .B(net112707), .Y(n3728) );
  AO21X2 U2008 ( .A0(n9932), .A1(n9931), .B0(net112731), .Y(n9210) );
  AO22X2 U2009 ( .A0(mem_rdata_I[22]), .A1(n113), .B0(n5466), .B1(n11252), .Y(
        n9853) );
  INVX3 U2010 ( .A(n5329), .Y(n4678) );
  AO22X2 U2011 ( .A0(mem_rdata_I[54]), .A1(n115), .B0(n5466), .B1(n11284), .Y(
        n9858) );
  AO22X2 U2012 ( .A0(mem_rdata_I[32]), .A1(n115), .B0(n5469), .B1(n11262), .Y(
        n9683) );
  INVX3 U2013 ( .A(n5331), .Y(n4676) );
  AO22X2 U2014 ( .A0(mem_rdata_I[86]), .A1(n115), .B0(n5466), .B1(n11316), .Y(
        n9848) );
  AO22X2 U2015 ( .A0(mem_rdata_I[122]), .A1(n115), .B0(n5465), .B1(n11352), 
        .Y(n9696) );
  AO22X2 U2016 ( .A0(mem_rdata_I[117]), .A1(n114), .B0(n5466), .B1(n11347), 
        .Y(n9863) );
  AO22X2 U2017 ( .A0(mem_rdata_I[112]), .A1(n113), .B0(n5469), .B1(n11342), 
        .Y(n10060) );
  INVX3 U2018 ( .A(n5514), .Y(n5506) );
  NAND3BX1 U2019 ( .AN(n10269), .B(n10214), .C(n10215), .Y(n10218) );
  NAND3BX1 U2020 ( .AN(n10919), .B(n10918), .C(n10920), .Y(n10924) );
  CLKINVX1 U2021 ( .A(n11098), .Y(n11095) );
  CLKINVX1 U2022 ( .A(n11113), .Y(n11110) );
  CLKINVX1 U2023 ( .A(n11151), .Y(n11118) );
  AND4X4 U2024 ( .A(n7703), .B(n7702), .C(n7701), .D(n7700), .Y(n3797) );
  NAND2X2 U2025 ( .A(n4564), .B(n10499), .Y(n10365) );
  XOR2X2 U2026 ( .A(n10200), .B(ICACHE_addr[23]), .Y(n10342) );
  BUFX12 U2027 ( .A(net98375), .Y(net113592) );
  AOI33X1 U2028 ( .A0(\i_MIPS/Hazard_detection/n7 ), .A1(n5944), .A2(n5943), 
        .B0(\i_MIPS/Hazard_detection/n4 ), .B1(n5942), .B2(n5941), .Y(n6173)
         );
  INVX3 U2029 ( .A(n5514), .Y(n5508) );
  INVX16 U2030 ( .A(n5591), .Y(n5589) );
  INVX3 U2031 ( .A(n5512), .Y(n5511) );
  INVX3 U2032 ( .A(n5515), .Y(n5507) );
  INVX12 U2033 ( .A(n4047), .Y(DCACHE_addr[0]) );
  INVX16 U2034 ( .A(n3518), .Y(DCACHE_addr[2]) );
  CLKINVX1 U2035 ( .A(net113541), .Y(n3518) );
  CLKBUFX3 U2036 ( .A(net113540), .Y(net113541) );
  INVX12 U2037 ( .A(n3889), .Y(mem_wdata_I[4]) );
  NAND2BX1 U2038 ( .AN(n11361), .B(n11234), .Y(n3889) );
  INVX12 U2039 ( .A(n3890), .Y(mem_wdata_I[5]) );
  NAND2BX1 U2040 ( .AN(n11361), .B(n11235), .Y(n3890) );
  INVX12 U2041 ( .A(n3891), .Y(mem_wdata_I[6]) );
  NAND2BX1 U2042 ( .AN(n11361), .B(n11236), .Y(n3891) );
  INVX12 U2043 ( .A(n3893), .Y(mem_wdata_I[7]) );
  NAND2BX1 U2044 ( .AN(n11361), .B(n11237), .Y(n3893) );
  INVX16 U2045 ( .A(n3998), .Y(mem_wdata_I[109]) );
  CLKINVX12 U2046 ( .A(n4008), .Y(mem_wdata_I[112]) );
  INVX12 U2047 ( .A(n3996), .Y(mem_wdata_I[120]) );
  OR2X1 U2048 ( .A(n11361), .B(n3997), .Y(n3996) );
  CLKINVX12 U2049 ( .A(n4022), .Y(mem_wdata_I[121]) );
  CLKINVX12 U2050 ( .A(n4001), .Y(mem_wdata_I[123]) );
  INVX12 U2051 ( .A(n4011), .Y(mem_wdata_I[126]) );
  NAND2BX1 U2052 ( .AN(n11361), .B(n11356), .Y(n4011) );
  INVX12 U2053 ( .A(n3865), .Y(mem_addr_I[9]) );
  AOI2BB2X1 U2054 ( .B0(n4794), .B1(n11367), .A0N(n3650), .A1N(n4349), .Y(
        n3885) );
  INVX12 U2055 ( .A(n1829), .Y(mem_addr_I[12]) );
  NOR2X1 U2056 ( .A(n4328), .B(n11361), .Y(n4330) );
  NOR2X1 U2057 ( .A(n4329), .B(\i_MIPS/PC/n16 ), .Y(n4331) );
  BUFX12 U2058 ( .A(n12835), .Y(mem_addr_I[17]) );
  INVX12 U2059 ( .A(n1828), .Y(mem_addr_I[29]) );
  INVX12 U2060 ( .A(n4719), .Y(mem_addr_I[30]) );
  CLKINVX1 U2061 ( .A(n12824), .Y(n4719) );
  INVX12 U2062 ( .A(n1830), .Y(mem_addr_I[31]) );
  BUFX16 U2063 ( .A(n11546), .Y(mem_read_I) );
  INVX12 U2064 ( .A(n3855), .Y(mem_wdata_D[1]) );
  NAND2BX1 U2065 ( .AN(net113725), .B(n11391), .Y(n3855) );
  INVX12 U2066 ( .A(n3857), .Y(mem_wdata_D[3]) );
  OR2X1 U2067 ( .A(net113725), .B(n10513), .Y(n3857) );
  INVX12 U2068 ( .A(n3858), .Y(mem_wdata_D[9]) );
  OR2X1 U2069 ( .A(net113725), .B(n10771), .Y(n3858) );
  INVX12 U2070 ( .A(n3860), .Y(mem_wdata_D[11]) );
  OR2X1 U2071 ( .A(net113605), .B(n10783), .Y(n3860) );
  INVX12 U2072 ( .A(n3862), .Y(mem_wdata_D[12]) );
  NAND2BX1 U2073 ( .AN(net113725), .B(n11401), .Y(n3862) );
  INVX12 U2074 ( .A(n3864), .Y(mem_wdata_D[14]) );
  NAND2BX1 U2075 ( .AN(net113725), .B(n11403), .Y(n3864) );
  INVX12 U2076 ( .A(n3867), .Y(mem_wdata_D[15]) );
  OR2X1 U2077 ( .A(net113725), .B(n10192), .Y(n3867) );
  INVX12 U2078 ( .A(n3868), .Y(mem_wdata_D[16]) );
  OR2X1 U2079 ( .A(net113725), .B(n10455), .Y(n3868) );
  INVX12 U2080 ( .A(n3869), .Y(mem_wdata_D[17]) );
  OR2X1 U2081 ( .A(net113725), .B(n10601), .Y(n3869) );
  INVX12 U2082 ( .A(n3870), .Y(mem_wdata_D[18]) );
  OR2X1 U2083 ( .A(net113725), .B(n10614), .Y(n3870) );
  INVX12 U2084 ( .A(n3871), .Y(mem_wdata_D[20]) );
  OR2X1 U2085 ( .A(net113725), .B(n10526), .Y(n3871) );
  INVX12 U2086 ( .A(n3883), .Y(mem_wdata_D[21]) );
  OR2X1 U2087 ( .A(net113725), .B(n10538), .Y(n3883) );
  INVX12 U2088 ( .A(n3884), .Y(mem_wdata_D[22]) );
  OR2X1 U2089 ( .A(net113725), .B(n10550), .Y(n3884) );
  INVX12 U2090 ( .A(n4003), .Y(mem_wdata_D[23]) );
  OR2X1 U2091 ( .A(net113725), .B(n10562), .Y(n4003) );
  INVX12 U2092 ( .A(n4004), .Y(mem_wdata_D[24]) );
  OR2X1 U2093 ( .A(net113725), .B(n10575), .Y(n4004) );
  INVX12 U2094 ( .A(n4006), .Y(mem_wdata_D[25]) );
  OR2X1 U2095 ( .A(net113725), .B(n10429), .Y(n4006) );
  INVX12 U2096 ( .A(n4010), .Y(mem_wdata_D[26]) );
  OR2X1 U2097 ( .A(net113725), .B(n10417), .Y(n4010) );
  INVX12 U2098 ( .A(n4012), .Y(mem_wdata_D[27]) );
  OR2X1 U2099 ( .A(net113725), .B(n10468), .Y(n4012) );
  INVX12 U2100 ( .A(n4015), .Y(mem_wdata_D[30]) );
  OR2X1 U2101 ( .A(net113725), .B(n10689), .Y(n4015) );
  INVX12 U2102 ( .A(n4016), .Y(mem_wdata_D[31]) );
  OR2X1 U2103 ( .A(net113725), .B(n11209), .Y(n4016) );
  INVX12 U2104 ( .A(n4017), .Y(mem_wdata_D[33]) );
  OR2X1 U2105 ( .A(net113725), .B(n10847), .Y(n4017) );
  INVX12 U2106 ( .A(n4021), .Y(mem_wdata_D[34]) );
  OR2X1 U2107 ( .A(net113725), .B(n11178), .Y(n4021) );
  INVX12 U2108 ( .A(n4023), .Y(mem_wdata_D[35]) );
  OR2X1 U2109 ( .A(net113725), .B(n10516), .Y(n4023) );
  INVX12 U2110 ( .A(n4032), .Y(mem_wdata_D[37]) );
  OR2X1 U2111 ( .A(net113725), .B(n10761), .Y(n4032) );
  INVX12 U2112 ( .A(n4033), .Y(mem_wdata_D[38]) );
  OR2X1 U2113 ( .A(net113725), .B(net100023), .Y(n4033) );
  INVX12 U2114 ( .A(n4034), .Y(mem_wdata_D[39]) );
  NAND2BX1 U2115 ( .AN(net113725), .B(n11427), .Y(n4034) );
  INVX12 U2116 ( .A(n4037), .Y(mem_wdata_D[40]) );
  OR2X1 U2117 ( .A(net113725), .B(n10826), .Y(n4037) );
  INVX12 U2118 ( .A(n4041), .Y(mem_wdata_D[41]) );
  INVX12 U2119 ( .A(n4048), .Y(mem_wdata_D[42]) );
  OR2X1 U2120 ( .A(net113725), .B(n10592), .Y(n4048) );
  INVX12 U2121 ( .A(n4052), .Y(mem_wdata_D[43]) );
  OR2X1 U2122 ( .A(net113725), .B(n10786), .Y(n4052) );
  INVX12 U2123 ( .A(n4056), .Y(mem_wdata_D[44]) );
  OR2X1 U2124 ( .A(net113725), .B(n10798), .Y(n4056) );
  INVX12 U2125 ( .A(n4038), .Y(mem_wdata_D[55]) );
  OR2X1 U2126 ( .A(net113725), .B(n10565), .Y(n4038) );
  INVX12 U2127 ( .A(n4043), .Y(mem_wdata_D[56]) );
  OR2X1 U2128 ( .A(net113725), .B(n10578), .Y(n4043) );
  INVX12 U2129 ( .A(n4049), .Y(mem_wdata_D[57]) );
  OR2X1 U2130 ( .A(net113725), .B(n10432), .Y(n4049) );
  INVX12 U2131 ( .A(n4053), .Y(mem_wdata_D[60]) );
  OR2X1 U2132 ( .A(net113725), .B(n10404), .Y(n4053) );
  INVX12 U2133 ( .A(n4036), .Y(mem_wdata_D[63]) );
  OR2X1 U2134 ( .A(net113725), .B(n11214), .Y(n4036) );
  INVX12 U2135 ( .A(n4040), .Y(mem_wdata_D[64]) );
  OR2X1 U2136 ( .A(net113725), .B(n10854), .Y(n4040) );
  INVX12 U2137 ( .A(n4045), .Y(mem_wdata_D[65]) );
  OR2X1 U2138 ( .A(net113725), .B(n10841), .Y(n4045) );
  INVX12 U2139 ( .A(n4051), .Y(mem_wdata_D[66]) );
  OR2X1 U2140 ( .A(net113725), .B(n11172), .Y(n4051) );
  INVX12 U2141 ( .A(n4055), .Y(mem_wdata_D[67]) );
  INVX12 U2142 ( .A(n4060), .Y(mem_wdata_D[68]) );
  OR2X1 U2143 ( .A(net113725), .B(n10148), .Y(n4060) );
  INVX12 U2144 ( .A(n4064), .Y(mem_wdata_D[69]) );
  OR2X1 U2145 ( .A(net113725), .B(n10755), .Y(n4064) );
  INVX12 U2146 ( .A(n4035), .Y(mem_wdata_D[70]) );
  OR2X1 U2147 ( .A(net113725), .B(net100029), .Y(n4035) );
  INVX12 U2148 ( .A(n4057), .Y(mem_wdata_D[72]) );
  OR2X1 U2149 ( .A(net113725), .B(n10820), .Y(n4057) );
  INVX12 U2150 ( .A(n4039), .Y(mem_wdata_D[73]) );
  OR2X1 U2151 ( .A(net113725), .B(n10768), .Y(n4039) );
  INVX12 U2152 ( .A(n4044), .Y(mem_wdata_D[74]) );
  OR2X1 U2153 ( .A(net113725), .B(n10586), .Y(n4044) );
  INVX12 U2154 ( .A(n4050), .Y(mem_wdata_D[75]) );
  OR2X1 U2155 ( .A(net113725), .B(n10780), .Y(n4050) );
  INVX12 U2156 ( .A(n1831), .Y(mem_wdata_D[76]) );
  INVX12 U2157 ( .A(n4054), .Y(mem_wdata_D[77]) );
  OR2X1 U2158 ( .A(net113725), .B(n10804), .Y(n4054) );
  INVX12 U2159 ( .A(n4058), .Y(mem_wdata_D[78]) );
  NAND2BX1 U2160 ( .AN(net113725), .B(n11465), .Y(n4058) );
  INVX12 U2161 ( .A(n4062), .Y(mem_wdata_D[80]) );
  OR2X1 U2162 ( .A(net113725), .B(n10452), .Y(n4062) );
  INVX12 U2163 ( .A(n4068), .Y(mem_wdata_D[82]) );
  OR2X1 U2164 ( .A(net113725), .B(n10611), .Y(n4068) );
  INVX12 U2165 ( .A(n4069), .Y(mem_wdata_D[89]) );
  OR2X1 U2166 ( .A(net113725), .B(n10426), .Y(n4069) );
  INVX12 U2167 ( .A(n4061), .Y(mem_wdata_D[90]) );
  OR2X1 U2168 ( .A(net113725), .B(n10414), .Y(n4061) );
  INVX12 U2169 ( .A(n1890), .Y(mem_wdata_D[93]) );
  INVX12 U2170 ( .A(n4065), .Y(mem_wdata_D[94]) );
  OR2X1 U2171 ( .A(net113725), .B(n10686), .Y(n4065) );
  INVX12 U2172 ( .A(n1844), .Y(mem_wdata_D[95]) );
  INVX12 U2173 ( .A(n1846), .Y(mem_wdata_D[96]) );
  INVX12 U2174 ( .A(n1847), .Y(mem_wdata_D[101]) );
  INVX12 U2175 ( .A(n1845), .Y(mem_wdata_D[102]) );
  INVX12 U2176 ( .A(n1848), .Y(mem_wdata_D[103]) );
  INVX12 U2177 ( .A(n4070), .Y(mem_wdata_D[115]) );
  OR2X1 U2178 ( .A(net113725), .B(n10172), .Y(n4070) );
  INVX12 U2179 ( .A(n1814), .Y(mem_addr_D[7]) );
  INVX12 U2180 ( .A(n1815), .Y(mem_addr_D[8]) );
  INVX12 U2181 ( .A(n1816), .Y(mem_addr_D[9]) );
  INVX12 U2182 ( .A(n1818), .Y(mem_addr_D[11]) );
  INVX12 U2183 ( .A(n1819), .Y(mem_addr_D[12]) );
  INVX12 U2184 ( .A(n1820), .Y(mem_addr_D[13]) );
  INVX12 U2185 ( .A(n1821), .Y(mem_addr_D[14]) );
  INVX12 U2186 ( .A(n1823), .Y(mem_addr_D[16]) );
  INVX12 U2187 ( .A(n1825), .Y(mem_addr_D[19]) );
  INVX12 U2188 ( .A(n1826), .Y(mem_addr_D[20]) );
  INVX12 U2189 ( .A(n1827), .Y(mem_addr_D[21]) );
  OAI2BB2XL U2190 ( .B0(\i_MIPS/n228 ), .B1(net110227), .A0N(n174), .A1N(
        n10968), .Y(\i_MIPS/N76 ) );
  NAND3BX2 U2191 ( .AN(n11102), .B(n11101), .C(n11100), .Y(\i_MIPS/PC/n49 ) );
  OA22X2 U2192 ( .A0(n11099), .A1(net140281), .B0(net98430), .B1(n11098), .Y(
        n11101) );
  NAND3X2 U2193 ( .A(n4172), .B(n4173), .C(n4174), .Y(n11102) );
  OA22X2 U2194 ( .A0(n10300), .A1(net140280), .B0(net98430), .B1(n10299), .Y(
        n10287) );
  NAND3BX2 U2195 ( .AN(n11092), .B(n11091), .C(n11090), .Y(\i_MIPS/PC/n47 ) );
  NAND3X2 U2196 ( .A(n4189), .B(n4190), .C(n4191), .Y(n11092) );
  AO22X1 U2197 ( .A0(n175), .A1(n10249), .B0(net113592), .B1(
        \i_MIPS/IR_ID[27] ), .Y(\i_MIPS/N82 ) );
  AO22X1 U2198 ( .A0(n174), .A1(n11164), .B0(net113592), .B1(
        \i_MIPS/IR_ID[29] ), .Y(\i_MIPS/N84 ) );
  NAND3BX2 U2199 ( .AN(n11023), .B(n11022), .C(n11021), .Y(\i_MIPS/PC/n54 ) );
  AOI2BB2X2 U2200 ( .B0(\i_MIPS/IF_ID[74] ), .B1(n150), .A0N(net110189), .A1N(
        \i_MIPS/n189 ), .Y(n10890) );
  AOI22X2 U2201 ( .A0(\i_MIPS/IF_ID[73] ), .A1(n149), .B0(net130576), .B1(n171), .Y(n10879) );
  OAI222X1 U2202 ( .A0(n3648), .A1(net110215), .B0(n4541), .B1(net110243), 
        .C0(n10876), .C1(net110249), .Y(n10881) );
  AOI2BB2X2 U2203 ( .B0(\i_MIPS/IF_ID[75] ), .B1(n148), .A0N(net110191), .A1N(
        \i_MIPS/n190 ), .Y(n10902) );
  NAND3X2 U2204 ( .A(n3536), .B(n3537), .C(n3538), .Y(n10394) );
  NAND3BX2 U2205 ( .AN(n10869), .B(n10868), .C(n10867), .Y(\i_MIPS/PC/n41 ) );
  OAI2BB2XL U2206 ( .B0(\i_MIPS/n173 ), .B1(net110225), .A0N(n10354), .A1N(
        n176), .Y(\i_MIPS/N114 ) );
  CLKINVX1 U2207 ( .A(n10355), .Y(n10354) );
  MXI2X1 U2208 ( .A(\i_MIPS/n329 ), .B(\i_MIPS/n328 ), .S0(n5504), .Y(
        \i_MIPS/n521 ) );
  NAND3BX2 U2209 ( .AN(n4136), .B(n4137), .C(n4138), .Y(\i_MIPS/PC/n58 ) );
  NAND3BX2 U2210 ( .AN(n11116), .B(n11115), .C(n11114), .Y(\i_MIPS/PC/n51 ) );
  NAND2X1 U2211 ( .A(n10708), .B(net110253), .Y(n10710) );
  AOI2BB2X1 U2212 ( .B0(\i_MIPS/IF_ID[95] ), .B1(n149), .A0N(net110189), .A1N(
        \i_MIPS/n210 ), .Y(n10709) );
  OAI2BB1X1 U2213 ( .A0N(net110251), .A1N(net98430), .B0(\i_MIPS/PC_o[1] ), 
        .Y(n10831) );
  MXI2X1 U2214 ( .A(\i_MIPS/n294 ), .B(\i_MIPS/n295 ), .S0(n5502), .Y(
        \i_MIPS/n422 ) );
  MXI2X1 U2215 ( .A(\i_MIPS/n302 ), .B(\i_MIPS/n303 ), .S0(n5505), .Y(
        \i_MIPS/n430 ) );
  OA22X2 U2216 ( .A0(n11069), .A1(net140281), .B0(net98430), .B1(n11068), .Y(
        n11071) );
  OR3X2 U2217 ( .A(n4431), .B(n4430), .C(n4429), .Y(n11006) );
  CLKMX2X2 U2218 ( .A(\I_cache/cache[5][142] ), .B(n11034), .S0(n5279), .Y(
        n11682) );
  NAND3X2 U2219 ( .A(n4183), .B(n4184), .C(n4185), .Y(n11199) );
  CLKMX2X2 U2220 ( .A(\D_cache/cache[4][73] ), .B(n4299), .S0(net112213), .Y(
        \D_cache/n1208 ) );
  CLKMX2X2 U2221 ( .A(\D_cache/cache[4][69] ), .B(n4301), .S0(net112213), .Y(
        \D_cache/n1240 ) );
  CLKMX2X2 U2222 ( .A(\D_cache/cache[4][41] ), .B(n4278), .S0(net112213), .Y(
        \D_cache/n1464 ) );
  CLKMX2X2 U2223 ( .A(\D_cache/cache[4][9] ), .B(n10767), .S0(net112213), .Y(
        \D_cache/n1720 ) );
  AO21X1 U2224 ( .A0(n5515), .A1(\i_MIPS/ID_EX_3 ), .B0(n4588), .Y(
        \i_MIPS/n525 ) );
  NAND2X1 U2225 ( .A(n4664), .B(n4494), .Y(n4700) );
  OAI2BB2X2 U2226 ( .B0(\i_MIPS/n167 ), .B1(net110219), .A0N(n175), .A1N(
        n11017), .Y(\i_MIPS/N108 ) );
  OAI2BB2XL U2227 ( .B0(\i_MIPS/n240 ), .B1(net110219), .A0N(n173), .A1N(
        n11066), .Y(\i_MIPS/N94 ) );
  CLKINVX1 U2228 ( .A(n11077), .Y(n11076) );
  OAI2BB2XL U2229 ( .B0(\i_MIPS/n159 ), .B1(net110225), .A0N(n10221), .A1N(
        n174), .Y(\i_MIPS/N100 ) );
  OAI2BB2X1 U2230 ( .B0(\i_MIPS/n160 ), .B1(net110217), .A0N(n173), .A1N(
        n11086), .Y(\i_MIPS/N101 ) );
  CLKINVX1 U2231 ( .A(n11097), .Y(n11096) );
  OAI2BB2XL U2232 ( .B0(\i_MIPS/n163 ), .B1(net110221), .A0N(n10927), .A1N(
        n173), .Y(\i_MIPS/N104 ) );
  OAI2BB2XL U2233 ( .B0(\i_MIPS/n170 ), .B1(net110219), .A0N(n175), .A1N(
        n10966), .Y(\i_MIPS/N111 ) );
  CLKINVX1 U2234 ( .A(n10967), .Y(n10966) );
  OAI2BB2XL U2235 ( .B0(\i_MIPS/n184 ), .B1(net110217), .A0N(n3515), .A1N(n176), .Y(\i_MIPS/N27 ) );
  OAI2BB2XL U2236 ( .B0(\i_MIPS/n202 ), .B1(net110217), .A0N(n10317), .A1N(
        n174), .Y(\i_MIPS/N45 ) );
  MXI2X1 U2237 ( .A(\i_MIPS/Pred_2bit/n1 ), .B(n10864), .S0(n4494), .Y(
        \i_MIPS/Pred_2bit/n8 ) );
  CLKMX2X2 U2238 ( .A(n4699), .B(\i_MIPS/Pred_2bit/current_state[0] ), .S0(
        n4664), .Y(n10864) );
  OAI2BB2XL U2239 ( .B0(\i_MIPS/n223 ), .B1(net110215), .A0N(n176), .A1N(
        n11083), .Y(\i_MIPS/N66 ) );
  OAI2BB2XL U2240 ( .B0(\i_MIPS/n218 ), .B1(net110227), .A0N(n176), .A1N(
        n10873), .Y(\i_MIPS/N61 ) );
  AOI2BB2X1 U2241 ( .B0(\i_MIPS/IF_ID[92] ), .B1(n150), .A0N(net110189), .A1N(
        \i_MIPS/n207 ), .Y(n10372) );
  NAND2X6 U2242 ( .A(n3721), .B(n6423), .Y(n8713) );
  CLKINVX6 U2243 ( .A(net102651), .Y(n4140) );
  AOI222X1 U2244 ( .A0(n5475), .A1(n11489), .B0(mem_rdata_D[103]), .B1(n117), 
        .C0(n12990), .C1(n5472), .Y(n10739) );
  BUFX6 U2245 ( .A(net99104), .Y(n178) );
  NAND2X4 U2246 ( .A(n3204), .B(net99042), .Y(n4113) );
  INVX2 U2247 ( .A(n4442), .Y(n163) );
  INVX3 U2248 ( .A(n8655), .Y(n4442) );
  NAND4X6 U2249 ( .A(n8285), .B(n8287), .C(n8284), .D(n8286), .Y(net99384) );
  AOI222XL U2250 ( .A0(n5487), .A1(n11441), .B0(mem_rdata_D[53]), .B1(n117), 
        .C0(n12976), .C1(n5483), .Y(n10542) );
  AO21X2 U2251 ( .A0(net99428), .A1(net99429), .B0(net113075), .Y(net99410) );
  OA22X1 U2252 ( .A0(net112681), .A1(n2370), .B0(net112575), .B1(n866), .Y(
        n7066) );
  CLKBUFX6 U2253 ( .A(net112703), .Y(net112681) );
  OA22X2 U2254 ( .A0(net112467), .A1(n1364), .B0(net112343), .B1(n2977), .Y(
        n7329) );
  NOR4X2 U2255 ( .A(n8372), .B(n8371), .C(n8370), .D(n8369), .Y(n8383) );
  AO22X1 U2256 ( .A0(net113445), .A1(n11470), .B0(net102346), .B1(n11501), .Y(
        n7823) );
  INVX1 U2257 ( .A(n11233), .Y(n9612) );
  MXI2X1 U2258 ( .A(\i_MIPS/n262 ), .B(\i_MIPS/n263 ), .S0(n5509), .Y(
        \i_MIPS/n390 ) );
  MX2X6 U2259 ( .A(\i_MIPS/n263 ), .B(n4649), .S0(n3771), .Y(n6588) );
  NAND2X6 U2260 ( .A(\i_MIPS/ALUin1[23] ), .B(n6583), .Y(n8925) );
  INVX3 U2261 ( .A(n11512), .Y(n10683) );
  OAI22X4 U2262 ( .A0(n10683), .A1(net102120), .B0(n10686), .B1(net102121), 
        .Y(n4602) );
  CLKINVX1 U2263 ( .A(n7109), .Y(n165) );
  AO22XL U2264 ( .A0(n174), .A1(n10244), .B0(net113592), .B1(
        \i_MIPS/IR_ID[26] ), .Y(\i_MIPS/N81 ) );
  OA22X1 U2265 ( .A0(n5178), .A1(n1473), .B0(n5134), .B1(n3086), .Y(n9940) );
  AO22XL U2266 ( .A0(n174), .A1(n10248), .B0(net113592), .B1(
        \i_MIPS/IR_ID[28] ), .Y(\i_MIPS/N83 ) );
  OAI2BB1X2 U2267 ( .A0N(net111405), .A1N(n10363), .B0(n10362), .Y(n10382) );
  INVX12 U2268 ( .A(n4828), .Y(n4825) );
  NAND2X1 U2269 ( .A(n4828), .B(\i_MIPS/n354 ), .Y(n8531) );
  NAND2X1 U2270 ( .A(n4828), .B(\i_MIPS/ALUin1[8] ), .Y(n7280) );
  OA21X2 U2271 ( .A0(\i_MIPS/ALUin1[19] ), .A1(n4818), .B0(n7022), .Y(n6670)
         );
  NAND3BX1 U2272 ( .AN(n4612), .B(n7022), .C(n7021), .Y(n7106) );
  AOI2BB1X2 U2273 ( .A0N(n8281), .A1N(n8280), .B0(n8332), .Y(n8283) );
  AO22X2 U2274 ( .A0(net113455), .A1(n11428), .B0(net113461), .B1(n11397), .Y(
        n6802) );
  AO22XL U2275 ( .A0(n175), .A1(n10958), .B0(net113592), .B1(net108963), .Y(
        \i_MIPS/N75 ) );
  MX2X2 U2276 ( .A(n6763), .B(n6762), .S0(net108963), .Y(net106418) );
  CLKBUFX12 U2277 ( .A(net101983), .Y(net112729) );
  AO21X2 U2278 ( .A0(net99536), .A1(net99537), .B0(net113075), .Y(net99693) );
  OAI211X2 U2279 ( .A0(n6802), .A1(n6801), .B0(net113437), .C0(n3709), .Y(
        net98951) );
  CLKMX2X12 U2280 ( .A(\i_MIPS/n267 ), .B(n4647), .S0(n3771), .Y(n6584) );
  NAND2X2 U2281 ( .A(n7781), .B(n8543), .Y(n7952) );
  INVX8 U2282 ( .A(n9263), .Y(n9179) );
  CLKINVX1 U2283 ( .A(n3520), .Y(n166) );
  NAND2X4 U2284 ( .A(net99270), .B(net134118), .Y(n3710) );
  INVX6 U2285 ( .A(n4801), .Y(n9174) );
  INVX4 U2286 ( .A(n10407), .Y(n8424) );
  NAND2X4 U2287 ( .A(n4099), .B(net99624), .Y(n4132) );
  INVX6 U2288 ( .A(net99624), .Y(n4100) );
  AO22X2 U2289 ( .A0(net113457), .A1(n11427), .B0(net113463), .B1(n11396), .Y(
        n7501) );
  NAND2X6 U2290 ( .A(n7200), .B(n3787), .Y(n3638) );
  INVX6 U2291 ( .A(n3562), .Y(n9019) );
  OA22X1 U2292 ( .A0(net112681), .A1(n2373), .B0(net112575), .B1(n869), .Y(
        n7054) );
  OA22X1 U2293 ( .A0(net112681), .A1(n923), .B0(net112565), .B1(n2450), .Y(
        n6276) );
  INVX3 U2294 ( .A(net99016), .Y(net107237) );
  OA22X2 U2295 ( .A0(n8726), .A1(n7695), .B0(n8728), .B1(n7699), .Y(n7617) );
  OA22X2 U2296 ( .A0(n8726), .A1(n8725), .B0(n8724), .B1(n9275), .Y(n8740) );
  AND3X2 U2297 ( .A(n7035), .B(n3508), .C(n4924), .Y(n7046) );
  BUFX16 U2298 ( .A(n9259), .Y(n4924) );
  CLKAND2X3 U2299 ( .A(n7111), .B(n8261), .Y(n7044) );
  OAI221X2 U2300 ( .A0(\i_MIPS/n364 ), .A1(n4810), .B0(\i_MIPS/n363 ), .B1(
        n4803), .C0(n6256), .Y(n8542) );
  NAND2X4 U2301 ( .A(n3783), .B(n9009), .Y(n9011) );
  OAI221X4 U2302 ( .A0(n9275), .A1(n8997), .B0(n8887), .B1(n8886), .C0(n4501), 
        .Y(n8935) );
  CLKMX2X2 U2303 ( .A(n7866), .B(n7868), .S0(n5590), .Y(n7559) );
  CLKMX2X4 U2304 ( .A(n7868), .B(n7863), .S0(n5590), .Y(n7198) );
  OAI221X1 U2305 ( .A0(n7560), .A1(n7867), .B0(n4797), .B1(n7868), .C0(n7476), 
        .Y(n7197) );
  OAI221X4 U2306 ( .A0(\i_MIPS/n342 ), .A1(n4825), .B0(\i_MIPS/n343 ), .B1(
        n4817), .C0(n6951), .Y(n7868) );
  AOI2BB2X2 U2307 ( .B0(n4927), .B1(n3627), .A0N(n4570), .A1N(n4798), .Y(n6866) );
  CLKXOR2X8 U2308 ( .A(n10941), .B(n10944), .Y(n169) );
  OA22X1 U2309 ( .A0(n5434), .A1(n1934), .B0(n5395), .B1(n353), .Y(n9513) );
  OA22X1 U2310 ( .A0(n5441), .A1(n948), .B0(n5395), .B1(n2473), .Y(n9941) );
  OA22X1 U2311 ( .A0(net112679), .A1(n1535), .B0(net112573), .B1(n3148), .Y(
        n7499) );
  OAI221X4 U2312 ( .A0(\i_MIPS/ALUin1[19] ), .A1(n4810), .B0(
        \i_MIPS/ALUin1[20] ), .B1(n4803), .C0(n8532), .Y(n8888) );
  NAND2X4 U2313 ( .A(\i_MIPS/ALUin1[19] ), .B(n6569), .Y(n8517) );
  NAND2X6 U2314 ( .A(\i_MIPS/ALUin1[19] ), .B(n6577), .Y(n8524) );
  XOR2X4 U2315 ( .A(n169), .B(n168), .Y(n10942) );
  OAI222X2 U2316 ( .A0(n8659), .A1(n7042), .B0(n9129), .B1(n7561), .C0(n284), 
        .C1(n8805), .Y(n7043) );
  NOR3X8 U2317 ( .A(n8168), .B(n8170), .C(n8169), .Y(n3547) );
  NOR2BX2 U2318 ( .AN(n9580), .B(n9581), .Y(n4616) );
  OAI211X2 U2319 ( .A0(n8927), .A1(n8332), .B0(n8331), .C0(n8330), .Y(n170) );
  INVX12 U2320 ( .A(n6510), .Y(n9312) );
  CLKBUFX2 U2321 ( .A(n9312), .Y(n4992) );
  NAND2X4 U2322 ( .A(n4659), .B(n4652), .Y(n6510) );
  INVX3 U2323 ( .A(n6927), .Y(n6929) );
  INVX4 U2324 ( .A(n4863), .Y(n4855) );
  INVX4 U2325 ( .A(n4860), .Y(n4857) );
  INVX6 U2326 ( .A(n4862), .Y(n4856) );
  INVX3 U2327 ( .A(n4859), .Y(n4858) );
  MXI2XL U2328 ( .A(\i_MIPS/n304 ), .B(\i_MIPS/n305 ), .S0(n5504), .Y(
        \i_MIPS/n432 ) );
  BUFX8 U2329 ( .A(n5407), .Y(n5406) );
  INVX3 U2330 ( .A(n8889), .Y(n8892) );
  NAND2X8 U2331 ( .A(n7853), .B(n8524), .Y(n8072) );
  CLKINVX20 U2332 ( .A(n172), .Y(n173) );
  CLKINVX20 U2333 ( .A(n172), .Y(n174) );
  CLKINVX20 U2334 ( .A(n172), .Y(n175) );
  CLKINVX20 U2335 ( .A(n172), .Y(n176) );
  OR2X6 U2336 ( .A(n7794), .B(n7795), .Y(n3557) );
  NAND4X6 U2337 ( .A(\i_MIPS/ALUOp[1] ), .B(n4414), .C(n6209), .D(n6216), .Y(
        n6213) );
  CLKINVX1 U2338 ( .A(n6424), .Y(n6765) );
  OAI221X4 U2339 ( .A0(\i_MIPS/n352 ), .A1(n4826), .B0(\i_MIPS/n353 ), .B1(
        n4817), .C0(n6262), .Y(n6424) );
  NAND4X6 U2340 ( .A(n3749), .B(n8363), .C(n8362), .D(n8361), .Y(n10407) );
  CLKBUFX3 U2341 ( .A(net112377), .Y(net112349) );
  BUFX12 U2342 ( .A(net112383), .Y(net112377) );
  NOR2X6 U2343 ( .A(n9019), .B(n9018), .Y(n4409) );
  CLKINVX8 U2344 ( .A(n3561), .Y(n3562) );
  BUFX12 U2345 ( .A(n6445), .Y(n4067) );
  OA22XL U2346 ( .A0(net112081), .A1(n1235), .B0(net111957), .B1(n2840), .Y(
        n9095) );
  OA22XL U2347 ( .A0(net112081), .A1(n2446), .B0(net111957), .B1(n471), .Y(
        n9056) );
  BUFX4 U2348 ( .A(net112085), .Y(net112081) );
  BUFX8 U2349 ( .A(n4706), .Y(n177) );
  INVXL U2350 ( .A(n9309), .Y(n179) );
  CLKINVX1 U2351 ( .A(n4976), .Y(n180) );
  INVX8 U2352 ( .A(n6513), .Y(n9309) );
  BUFX16 U2353 ( .A(n9309), .Y(n4976) );
  NAND2X2 U2354 ( .A(n4686), .B(n4582), .Y(n6513) );
  INVX6 U2355 ( .A(n4836), .Y(n4835) );
  INVX4 U2356 ( .A(n4840), .Y(n4832) );
  INVX4 U2357 ( .A(n4839), .Y(n4833) );
  INVX4 U2358 ( .A(n4837), .Y(n4834) );
  CLKINVX1 U2359 ( .A(n7035), .Y(n7026) );
  NOR3BX2 U2360 ( .AN(\i_MIPS/Register/n120 ), .B(\i_MIPS/Reg_W[3] ), .C(
        \i_MIPS/Reg_W[4] ), .Y(\i_MIPS/Register/n140 ) );
  NOR2BX2 U2361 ( .AN(\i_MIPS/EX_MEM_0 ), .B(\i_MIPS/EX_MEM_74 ), .Y(
        \i_MIPS/Register/n120 ) );
  AOI2BB1X2 U2362 ( .A0N(n9140), .A1N(n7200), .B0(n8911), .Y(n6435) );
  CLKINVX12 U2363 ( .A(n8736), .Y(n7200) );
  AO22X2 U2364 ( .A0(n8916), .A1(n4569), .B0(n9140), .B1(n8343), .Y(n7883) );
  INVX20 U2365 ( .A(n140), .Y(n9140) );
  NOR4X4 U2366 ( .A(n8358), .B(n8357), .C(n8356), .D(n8355), .Y(n8362) );
  NAND2X8 U2367 ( .A(n9140), .B(n3787), .Y(n9275) );
  BUFX16 U2368 ( .A(n11140), .Y(n5451) );
  BUFX8 U2369 ( .A(n5448), .Y(n5429) );
  INVX4 U2370 ( .A(n5515), .Y(n5503) );
  INVX3 U2371 ( .A(n5514), .Y(n5504) );
  INVX4 U2372 ( .A(n5513), .Y(n5509) );
  BUFX6 U2373 ( .A(n5364), .Y(n5363) );
  BUFX4 U2374 ( .A(n5362), .Y(n5330) );
  CLKBUFX3 U2375 ( .A(n5275), .Y(n5272) );
  BUFX16 U2376 ( .A(n5275), .Y(n5274) );
  BUFX12 U2377 ( .A(n11136), .Y(n5144) );
  CLKBUFX4 U2378 ( .A(net112377), .Y(net112353) );
  CLKBUFX8 U2379 ( .A(net111979), .Y(net111955) );
  BUFX4 U2380 ( .A(net112271), .Y(net112229) );
  BUFX12 U2381 ( .A(net112257), .Y(net112237) );
  BUFX8 U2382 ( .A(n5448), .Y(n5428) );
  BUFX12 U2383 ( .A(n5364), .Y(n5362) );
  BUFX4 U2384 ( .A(n5363), .Y(n5357) );
  CLKBUFX3 U2385 ( .A(net112085), .Y(net112083) );
  CLKBUFX2 U2386 ( .A(net111983), .Y(net111961) );
  CLKBUFX8 U2387 ( .A(n3750), .Y(net111957) );
  BUFX8 U2388 ( .A(n5231), .Y(n5229) );
  CLKBUFX3 U2389 ( .A(n5319), .Y(n5317) );
  BUFX3 U2390 ( .A(net112105), .Y(net112101) );
  BUFX4 U2391 ( .A(net112087), .Y(net112071) );
  CLKBUFX3 U2392 ( .A(net112089), .Y(net112061) );
  INVX6 U2393 ( .A(n3730), .Y(net100079) );
  BUFX12 U2394 ( .A(net112231), .Y(net112241) );
  INVX4 U2395 ( .A(n5512), .Y(n5505) );
  INVX3 U2396 ( .A(n5513), .Y(n5502) );
  INVX4 U2397 ( .A(n5512), .Y(n5510) );
  BUFX6 U2398 ( .A(n5144), .Y(n5188) );
  BUFX4 U2399 ( .A(net112385), .Y(n3688) );
  CLKBUFX3 U2400 ( .A(net112377), .Y(net112337) );
  BUFX16 U2401 ( .A(n11135), .Y(n5143) );
  BUFX4 U2402 ( .A(net112089), .Y(net112063) );
  CLKBUFX4 U2403 ( .A(net112503), .Y(net112471) );
  CLKBUFX3 U2404 ( .A(net112379), .Y(net112303) );
  CLKBUFX2 U2405 ( .A(net112383), .Y(net112331) );
  BUFX6 U2406 ( .A(net112187), .Y(net112169) );
  CLKBUFX6 U2407 ( .A(n5464), .Y(n5468) );
  BUFX8 U2408 ( .A(n5451), .Y(n5450) );
  CLKBUFX2 U2409 ( .A(n5231), .Y(n5230) );
  BUFX4 U2410 ( .A(net112107), .Y(net112087) );
  CLKBUFX3 U2411 ( .A(net112497), .Y(net112491) );
  CLKBUFX3 U2412 ( .A(net112499), .Y(net112483) );
  CLKBUFX3 U2413 ( .A(net112499), .Y(net112487) );
  CLKBUFX8 U2414 ( .A(net111983), .Y(net111965) );
  CLKBUFX4 U2415 ( .A(net111979), .Y(net111905) );
  BUFX16 U2416 ( .A(net112145), .Y(net112159) );
  INVX1 U2417 ( .A(net109181), .Y(net113667) );
  CLKBUFX8 U2418 ( .A(net112271), .Y(net112245) );
  CLKBUFX8 U2419 ( .A(net112231), .Y(net112239) );
  BUFX16 U2420 ( .A(net112105), .Y(net112095) );
  CLKBUFX8 U2421 ( .A(net112107), .Y(net112089) );
  BUFX6 U2422 ( .A(net112095), .Y(net112041) );
  BUFX16 U2423 ( .A(net134103), .Y(net112383) );
  BUFX4 U2424 ( .A(net134103), .Y(net112381) );
  BUFX6 U2425 ( .A(net112383), .Y(net112329) );
  BUFX4 U2426 ( .A(net112381), .Y(net112339) );
  INVX3 U2427 ( .A(net113605), .Y(net113608) );
  CLKBUFX3 U2428 ( .A(n5143), .Y(n5116) );
  CLKBUFX2 U2429 ( .A(n5432), .Y(n5439) );
  CLKBUFX3 U2430 ( .A(n5384), .Y(n5388) );
  CLKBUFX3 U2431 ( .A(n5409), .Y(n5398) );
  BUFX4 U2432 ( .A(n5274), .Y(n5244) );
  BUFX12 U2433 ( .A(net111983), .Y(n3750) );
  CLKBUFX8 U2434 ( .A(net134103), .Y(net112379) );
  CLKBUFX8 U2435 ( .A(net112169), .Y(net112165) );
  CLKBUFX6 U2436 ( .A(net112259), .Y(net112233) );
  CLKBUFX8 U2437 ( .A(net112257), .Y(net112235) );
  BUFX4 U2438 ( .A(n5407), .Y(n5405) );
  BUFX6 U2439 ( .A(n5408), .Y(n5383) );
  BUFX6 U2440 ( .A(net111979), .Y(net111969) );
  CLKBUFX3 U2441 ( .A(n3750), .Y(net111949) );
  BUFX6 U2442 ( .A(net112383), .Y(net112301) );
  INVX3 U2443 ( .A(net113605), .Y(net113607) );
  CLKBUFX3 U2444 ( .A(n5188), .Y(n5159) );
  CLKBUFX3 U2445 ( .A(n5188), .Y(n5158) );
  BUFX16 U2446 ( .A(n5189), .Y(n5232) );
  BUFX8 U2447 ( .A(n5232), .Y(n5204) );
  BUFX4 U2448 ( .A(n5274), .Y(n5243) );
  BUFX3 U2449 ( .A(net112105), .Y(net112091) );
  CLKBUFX4 U2450 ( .A(net112105), .Y(net112093) );
  CLKBUFX3 U2451 ( .A(net112379), .Y(net112341) );
  CLKBUFX3 U2452 ( .A(net112379), .Y(net112345) );
  CLKBUFX3 U2453 ( .A(net112379), .Y(net112343) );
  CLKINVX4 U2454 ( .A(n11361), .Y(n4795) );
  CLKBUFX3 U2455 ( .A(n9310), .Y(n4980) );
  INVX16 U2456 ( .A(net109181), .Y(net113725) );
  INVX3 U2457 ( .A(net113605), .Y(net113606) );
  BUFX3 U2458 ( .A(net112695), .Y(net112657) );
  BUFX8 U2459 ( .A(net112703), .Y(net112679) );
  BUFX8 U2460 ( .A(net112687), .Y(net112667) );
  BUFX2 U2461 ( .A(n5319), .Y(n5288) );
  BUFX6 U2462 ( .A(n5408), .Y(n5385) );
  BUFX3 U2463 ( .A(net112269), .Y(net112257) );
  BUFX6 U2464 ( .A(n5143), .Y(n5119) );
  CLKBUFX8 U2465 ( .A(n5143), .Y(n5120) );
  CLKINVX3 U2466 ( .A(net112081), .Y(net112003) );
  CLKINVX3 U2467 ( .A(net112019), .Y(net112005) );
  CLKBUFX3 U2468 ( .A(net111963), .Y(net111945) );
  CLKINVX3 U2469 ( .A(net111905), .Y(net111871) );
  BUFX6 U2470 ( .A(n4964), .Y(n4967) );
  CLKBUFX2 U2471 ( .A(n4995), .Y(n4994) );
  BUFX4 U2472 ( .A(n4994), .Y(n4998) );
  OR3X2 U2473 ( .A(n4751), .B(mem_ready_D), .C(n4750), .Y(n186) );
  BUFX4 U2474 ( .A(n5471), .Y(n5470) );
  BUFX6 U2475 ( .A(n4999), .Y(n5002) );
  BUFX8 U2476 ( .A(net112583), .Y(net112577) );
  BUFX4 U2477 ( .A(net112187), .Y(net112145) );
  CLKBUFX2 U2478 ( .A(n5189), .Y(n5201) );
  BUFX8 U2479 ( .A(n5451), .Y(n3611) );
  BUFX6 U2480 ( .A(n5361), .Y(n5334) );
  CLKINVX3 U2481 ( .A(net112459), .Y(net112411) );
  CLKINVX3 U2482 ( .A(net112425), .Y(net112415) );
  CLKINVX3 U2483 ( .A(net112083), .Y(net111993) );
  BUFX4 U2484 ( .A(net111967), .Y(net111929) );
  CLKBUFX8 U2485 ( .A(n4918), .Y(n4916) );
  NAND2X4 U2486 ( .A(n4660), .B(n4657), .Y(n4484) );
  NAND2X2 U2487 ( .A(n9932), .B(n9931), .Y(n9126) );
  AND2XL U2488 ( .A(n10696), .B(n10695), .Y(n1834) );
  BUFX4 U2489 ( .A(n4481), .Y(n4921) );
  INVX6 U2490 ( .A(n4846), .Y(n4843) );
  INVX3 U2491 ( .A(n4845), .Y(n4844) );
  INVX4 U2492 ( .A(n4852), .Y(n4851) );
  BUFX16 U2493 ( .A(n4900), .Y(n4902) );
  BUFX4 U2494 ( .A(n9116), .Y(n4898) );
  CLKBUFX3 U2495 ( .A(n9116), .Y(n4896) );
  AND2XL U2496 ( .A(n10750), .B(n10751), .Y(n222) );
  AND2XL U2497 ( .A(net99428), .B(net99429), .Y(n223) );
  BUFX4 U2498 ( .A(n5464), .Y(n5467) );
  BUFX4 U2499 ( .A(net112705), .Y(net112697) );
  CLKBUFX6 U2500 ( .A(net112687), .Y(net112671) );
  BUFX16 U2501 ( .A(net112601), .Y(net112583) );
  BUFX16 U2502 ( .A(net112583), .Y(net112575) );
  CLKBUFX3 U2503 ( .A(n11135), .Y(n5142) );
  INVX3 U2504 ( .A(n5362), .Y(n4681) );
  INVX3 U2505 ( .A(n5332), .Y(n4679) );
  CLKINVX3 U2506 ( .A(net112301), .Y(net112293) );
  CLKINVX3 U2507 ( .A(net112301), .Y(net112295) );
  CLKINVX3 U2508 ( .A(net112349), .Y(net112281) );
  BUFX4 U2509 ( .A(n4890), .Y(n4893) );
  BUFX4 U2510 ( .A(n4890), .Y(n4894) );
  CLKINVX1 U2511 ( .A(n11361), .Y(n11547) );
  INVX12 U2512 ( .A(n11361), .Y(n4796) );
  BUFX4 U2513 ( .A(n11156), .Y(n5463) );
  INVX4 U2514 ( .A(n4628), .Y(n4957) );
  BUFX4 U2515 ( .A(n4909), .Y(n4911) );
  AND2XL U2516 ( .A(net98992), .B(net98993), .Y(n1849) );
  AND2XL U2517 ( .A(net99014), .B(net99015), .Y(n1857) );
  AND2XL U2518 ( .A(net98950), .B(net98951), .Y(n1838) );
  AND2XL U2519 ( .A(n10830), .B(n10829), .Y(n1841) );
  AND2XL U2520 ( .A(net99502), .B(net99503), .Y(n1858) );
  AND2XL U2521 ( .A(net99969), .B(net99970), .Y(n1850) );
  AND2XL U2522 ( .A(net99603), .B(net99604), .Y(n1855) );
  AND2XL U2523 ( .A(net99359), .B(net99360), .Y(n1836) );
  AND2XL U2524 ( .A(net99383), .B(net99382), .Y(n1835) );
  AND2XL U2525 ( .A(net114113), .B(net99405), .Y(n1851) );
  AND2XL U2526 ( .A(n10185), .B(n10184), .Y(n1837) );
  AND2XL U2527 ( .A(net99311), .B(net99312), .Y(n1852) );
  AND2XL U2528 ( .A(net99977), .B(net99978), .Y(n1853) );
  AND2XL U2529 ( .A(net99581), .B(net99582), .Y(n1856) );
  AND2XL U2530 ( .A(net99060), .B(net99061), .Y(n1843) );
  AND2XL U2531 ( .A(net99108), .B(net99109), .Y(n1839) );
  AND2XL U2532 ( .A(net100019), .B(net100020), .Y(n1840) );
  AND2XL U2533 ( .A(net100103), .B(net100104), .Y(n1842) );
  AND2XL U2534 ( .A(net99637), .B(net99638), .Y(n1995) );
  BUFX4 U2535 ( .A(n4918), .Y(n4917) );
  AND2XL U2536 ( .A(net99037), .B(net99038), .Y(n4573) );
  NOR2X1 U2537 ( .A(\i_MIPS/PC/n4 ), .B(ICACHE_addr[1]), .Y(n4693) );
  BUFX4 U2538 ( .A(n9311), .Y(n4981) );
  BUFX6 U2539 ( .A(n4993), .Y(n4997) );
  CLKBUFX2 U2540 ( .A(net98432), .Y(net110233) );
  BUFX4 U2541 ( .A(n9117), .Y(n4900) );
  BUFX4 U2542 ( .A(n4899), .Y(n4901) );
  CLKBUFX2 U2543 ( .A(net130301), .Y(net112713) );
  INVX1 U2544 ( .A(net104563), .Y(net102036) );
  BUFX4 U2545 ( .A(n9310), .Y(n4977) );
  INVX1 U2546 ( .A(n6515), .Y(n9307) );
  BUFX4 U2547 ( .A(n9307), .Y(n4966) );
  BUFX4 U2548 ( .A(n4964), .Y(n4965) );
  AND2XL U2549 ( .A(net98967), .B(net98968), .Y(n1854) );
  BUFX6 U2550 ( .A(n4999), .Y(n5000) );
  BUFX6 U2551 ( .A(n4999), .Y(n5001) );
  AND3X1 U2552 ( .A(n3755), .B(n4641), .C(n3768), .Y(n282) );
  CLKBUFX4 U2553 ( .A(net112701), .Y(net112687) );
  BUFX8 U2554 ( .A(net112691), .Y(net112665) );
  BUFX16 U2555 ( .A(net112589), .Y(net112563) );
  BUFX12 U2556 ( .A(net112585), .Y(net112569) );
  BUFX16 U2557 ( .A(net100081), .Y(net112187) );
  INVX3 U2558 ( .A(n5329), .Y(n4698) );
  INVX3 U2559 ( .A(n5363), .Y(n4680) );
  CLKINVX1 U2560 ( .A(n5330), .Y(n4677) );
  CLKINVX3 U2561 ( .A(net112229), .Y(net112197) );
  CLKINVX3 U2562 ( .A(net112229), .Y(net112195) );
  CLKBUFX2 U2563 ( .A(net112329), .Y(net112361) );
  CLKBUFX3 U2564 ( .A(net112381), .Y(net112335) );
  CLKBUFX3 U2565 ( .A(net112379), .Y(net112347) );
  BUFX16 U2566 ( .A(net112515), .Y(net112509) );
  CLKBUFX3 U2567 ( .A(net112499), .Y(net112473) );
  BUFX6 U2568 ( .A(\i_MIPS/IR_ID[20] ), .Y(net108963) );
  AND2XL U2569 ( .A(n7031), .B(n7030), .Y(n284) );
  BUFX6 U2570 ( .A(n4944), .Y(n4946) );
  AND2X2 U2571 ( .A(\i_MIPS/ALUin1[0] ), .B(n6423), .Y(n286) );
  BUFX16 U2572 ( .A(n12952), .Y(DCACHE_addr[16]) );
  CLKINVX1 U2573 ( .A(n7180), .Y(n7091) );
  INVX4 U2574 ( .A(n4960), .Y(n4959) );
  INVX4 U2575 ( .A(n4693), .Y(n5461) );
  AND2X2 U2576 ( .A(ICACHE_addr[1]), .B(\i_MIPS/PC/n4 ), .Y(n312) );
  NAND2X6 U2577 ( .A(n11229), .B(n11358), .Y(n11361) );
  AND2X2 U2578 ( .A(n12965), .B(n3238), .Y(n352) );
  NOR2X8 U2579 ( .A(n3824), .B(n3825), .Y(n432) );
  NAND2BX1 U2580 ( .AN(n10974), .B(n11359), .Y(n11156) );
  BUFX4 U2581 ( .A(net102344), .Y(net113439) );
  CLKBUFX6 U2582 ( .A(net102344), .Y(net113437) );
  INVX6 U2583 ( .A(n4452), .Y(n9279) );
  AND3X4 U2584 ( .A(n4067), .B(n6660), .C(n4585), .Y(n4452) );
  NAND2X1 U2585 ( .A(n4500), .B(n4653), .Y(n4485) );
  BUFX16 U2586 ( .A(net109185), .Y(net109181) );
  CLKINVX1 U2587 ( .A(n9226), .Y(n9117) );
  INVX6 U2588 ( .A(net102121), .Y(net102345) );
  CLKBUFX8 U2589 ( .A(net102345), .Y(net113447) );
  AND3X4 U2590 ( .A(n4164), .B(n4165), .C(n6142), .Y(n1608) );
  AND3X8 U2591 ( .A(n4223), .B(n4224), .C(n6117), .Y(n1609) );
  BUFX12 U2592 ( .A(net98564), .Y(net111409) );
  INVX4 U2593 ( .A(n4629), .Y(n4949) );
  INVX3 U2594 ( .A(n4951), .Y(n4948) );
  BUFX16 U2595 ( .A(net98396), .Y(net109791) );
  CLKBUFX3 U2596 ( .A(n4620), .Y(n4870) );
  BUFX6 U2597 ( .A(n4993), .Y(n4996) );
  AND3X8 U2598 ( .A(n4204), .B(n4205), .C(n6124), .Y(n1632) );
  BUFX4 U2599 ( .A(n9312), .Y(n4991) );
  CLKINVX1 U2600 ( .A(n6508), .Y(n9314) );
  XNOR2X4 U2601 ( .A(\i_MIPS/n325 ), .B(\i_MIPS/n327 ), .Y(n1636) );
  AND2XL U2602 ( .A(net99334), .B(net99335), .Y(n4571) );
  AND3X8 U2603 ( .A(n4186), .B(n4187), .C(n6089), .Y(n1637) );
  CLKINVX1 U2604 ( .A(net102094), .Y(net102372) );
  CLKBUFX3 U2605 ( .A(net102372), .Y(net113463) );
  CLKINVX1 U2606 ( .A(n9224), .Y(n9115) );
  BUFX3 U2607 ( .A(net112601), .Y(net112593) );
  BUFX16 U2608 ( .A(net112599), .Y(net112589) );
  INVX16 U2609 ( .A(net110257), .Y(net110249) );
  CLKINVX1 U2610 ( .A(n11168), .Y(n11213) );
  INVX20 U2611 ( .A(net112143), .Y(net112121) );
  CLKINVX3 U2612 ( .A(n5266), .Y(n5237) );
  CLKINVX3 U2613 ( .A(n5177), .Y(n5153) );
  CLKBUFX3 U2614 ( .A(n5226), .Y(n5216) );
  CLKINVX3 U2615 ( .A(n5201), .Y(n5198) );
  CLKBUFX3 U2616 ( .A(n5362), .Y(n5331) );
  CLKINVX3 U2617 ( .A(net112239), .Y(net112199) );
  CLKINVX3 U2618 ( .A(net112237), .Y(net112201) );
  CLKBUFX2 U2619 ( .A(net111979), .Y(net111977) );
  INVX8 U2620 ( .A(n3822), .Y(net134103) );
  CLKBUFX3 U2621 ( .A(n5143), .Y(n5114) );
  NAND2X1 U2622 ( .A(n4796), .B(n11354), .Y(n1803) );
  NAND2X1 U2623 ( .A(net113606), .B(n11504), .Y(n1804) );
  NAND2X1 U2624 ( .A(net113916), .B(n11505), .Y(n1805) );
  NAND2X1 U2625 ( .A(net113607), .B(n11512), .Y(n1806) );
  NAND2X1 U2626 ( .A(net113916), .B(n11513), .Y(n1807) );
  AOI22X1 U2627 ( .A0(DCACHE_addr[16]), .A1(mem_read_D), .B0(net109181), .B1(
        n3832), .Y(n1808) );
  AOI22X1 U2628 ( .A0(DCACHE_addr[21]), .A1(mem_read_D), .B0(net113608), .B1(
        n11533), .Y(n1809) );
  AOI22X1 U2629 ( .A0(n12946), .A1(mem_read_D), .B0(net109179), .B1(n11534), 
        .Y(n1810) );
  AOI22X1 U2630 ( .A0(n12945), .A1(mem_read_D), .B0(net113606), .B1(n11535), 
        .Y(n1811) );
  AOI22X1 U2631 ( .A0(n12944), .A1(mem_read_D), .B0(net113607), .B1(n11536), 
        .Y(n1812) );
  AOI22X1 U2632 ( .A0(DCACHE_addr[25]), .A1(mem_read_D), .B0(net113983), .B1(
        n11537), .Y(n1813) );
  AOI22X1 U2633 ( .A0(DCACHE_addr[5]), .A1(mem_read_D), .B0(net113607), .B1(
        n11518), .Y(n1814) );
  AOI22X1 U2634 ( .A0(DCACHE_addr[6]), .A1(mem_read_D), .B0(net113916), .B1(
        n11519), .Y(n1815) );
  AOI22X1 U2635 ( .A0(DCACHE_addr[7]), .A1(mem_read_D), .B0(net113606), .B1(
        n11520), .Y(n1816) );
  AOI22X1 U2636 ( .A0(DCACHE_addr[8]), .A1(mem_read_D), .B0(net113608), .B1(
        n11521), .Y(n1817) );
  AOI22X1 U2637 ( .A0(DCACHE_addr[9]), .A1(mem_read_D), .B0(net113916), .B1(
        n11522), .Y(n1818) );
  AOI22X1 U2638 ( .A0(n12958), .A1(mem_read_D), .B0(net113606), .B1(n11523), 
        .Y(n1819) );
  AOI22X1 U2639 ( .A0(DCACHE_addr[11]), .A1(mem_read_D), .B0(net113607), .B1(
        n11524), .Y(n1820) );
  AOI22X1 U2640 ( .A0(DCACHE_addr[12]), .A1(mem_read_D), .B0(net113607), .B1(
        n11525), .Y(n1821) );
  AOI22X1 U2641 ( .A0(DCACHE_addr[13]), .A1(mem_read_D), .B0(net113608), .B1(
        n11526), .Y(n1822) );
  AOI22X1 U2642 ( .A0(DCACHE_addr[14]), .A1(mem_read_D), .B0(net113606), .B1(
        n11527), .Y(n1823) );
  AOI22X1 U2643 ( .A0(n12953), .A1(mem_read_D), .B0(net113608), .B1(n11528), 
        .Y(n1824) );
  AOI22X1 U2644 ( .A0(n12951), .A1(mem_read_D), .B0(net109181), .B1(n11529), 
        .Y(n1825) );
  AOI22X1 U2645 ( .A0(DCACHE_addr[18]), .A1(mem_read_D), .B0(net109181), .B1(
        n11530), .Y(n1826) );
  AOI22X1 U2646 ( .A0(n12949), .A1(mem_read_D), .B0(net109181), .B1(n11531), 
        .Y(n1827) );
  INVX3 U2647 ( .A(n11083), .Y(n11089) );
  CLKINVX1 U2648 ( .A(n9156), .Y(n8430) );
  AOI22X1 U2649 ( .A0(ICACHE_addr[27]), .A1(mem_read_I), .B0(n11547), .B1(
        n11386), .Y(n1828) );
  AOI22X1 U2650 ( .A0(ICACHE_addr[10]), .A1(mem_read_I), .B0(n4796), .B1(
        n11369), .Y(n1829) );
  AOI22X1 U2651 ( .A0(ICACHE_addr[29]), .A1(mem_read_I), .B0(n11547), .B1(
        n3565), .Y(n1830) );
  NAND2X1 U2652 ( .A(net113607), .B(n11463), .Y(n1831) );
  CLKINVX1 U2653 ( .A(n11195), .Y(n3515) );
  NAND2X1 U2654 ( .A(net113607), .B(n11482), .Y(n1844) );
  NAND2X1 U2655 ( .A(net113606), .B(net98089), .Y(n1845) );
  NAND2X1 U2656 ( .A(net113607), .B(n11483), .Y(n1846) );
  NAND2X1 U2657 ( .A(net113606), .B(n11488), .Y(n1847) );
  NAND2X1 U2658 ( .A(net113606), .B(n11489), .Y(n1848) );
  INVX8 U2659 ( .A(n6260), .Y(n9133) );
  NAND2X4 U2660 ( .A(\i_MIPS/ALUin1[8] ), .B(n6243), .Y(n6846) );
  INVX8 U2661 ( .A(n4067), .Y(n4471) );
  NAND2X4 U2662 ( .A(n3719), .B(\i_MIPS/n367 ), .Y(n7355) );
  NAND2X1 U2663 ( .A(net113607), .B(n11480), .Y(n1890) );
  AND2X2 U2664 ( .A(n4797), .B(\i_MIPS/n340 ), .Y(n1891) );
  AND2X2 U2665 ( .A(n8648), .B(n8647), .Y(n1987) );
  OR3X2 U2666 ( .A(n9262), .B(n4594), .C(n8661), .Y(n2017) );
  INVX3 U2667 ( .A(net113592), .Y(net98432) );
  AND3X2 U2668 ( .A(n4148), .B(n4149), .C(n6131), .Y(n2437) );
  BUFX4 U2669 ( .A(n4941), .Y(n4939) );
  CLKBUFX3 U2670 ( .A(n4630), .Y(n4956) );
  MXI2X2 U2671 ( .A(n10855), .B(n10854), .S0(n5496), .Y(n10856) );
  MXI2X2 U2672 ( .A(n10852), .B(n10851), .S0(n5494), .Y(n10853) );
  MXI2X2 U2673 ( .A(n10799), .B(n10798), .S0(n5490), .Y(n10800) );
  MXI2X2 U2674 ( .A(n10599), .B(n10598), .S0(n5492), .Y(n10600) );
  MXI2X2 U2675 ( .A(n10587), .B(n10586), .S0(n5492), .Y(n10588) );
  MXI2X2 U2676 ( .A(n10533), .B(n10532), .S0(n5494), .Y(n10534) );
  MXI2X2 U2677 ( .A(n10187), .B(n10186), .S0(n5497), .Y(n10188) );
  INVX3 U2678 ( .A(n8069), .Y(n7955) );
  NAND2X6 U2679 ( .A(n4154), .B(n7950), .Y(n8069) );
  OR2X4 U2680 ( .A(\i_MIPS/n369 ), .B(n6233), .Y(n3197) );
  CLKBUFX3 U2681 ( .A(n4482), .Y(n4943) );
  BUFX4 U2682 ( .A(n4943), .Y(n4944) );
  AOI22X2 U2683 ( .A0(net113041), .A1(net98472), .B0(net102300), .B1(n7589), 
        .Y(n3198) );
  AND2X2 U2684 ( .A(n4658), .B(n4654), .Y(n4625) );
  AOI22X2 U2685 ( .A0(net113041), .A1(net98952), .B0(net102300), .B1(n6823), 
        .Y(n3203) );
  AOI22X2 U2686 ( .A0(net113041), .A1(net99062), .B0(net102300), .B1(n6906), 
        .Y(n3204) );
  AND4X2 U2687 ( .A(n287), .B(n229), .C(\i_MIPS/forward_unit/n25 ), .D(n4705), 
        .Y(\i_MIPS/forward_unit/n10 ) );
  INVX3 U2688 ( .A(\i_MIPS/forward_unit/n10 ), .Y(n6302) );
  AOI22X2 U2689 ( .A0(net99461), .A1(net113041), .B0(net102300), .B1(n7314), 
        .Y(n3218) );
  NAND3X1 U2690 ( .A(n8078), .B(n8079), .C(n9258), .Y(n3247) );
  AND2X4 U2691 ( .A(n9558), .B(n9572), .Y(n3257) );
  AND3X2 U2692 ( .A(n4548), .B(n9258), .C(n8344), .Y(n3259) );
  INVX3 U2693 ( .A(n6511), .Y(n9311) );
  BUFX4 U2694 ( .A(n4479), .Y(n4903) );
  BUFX4 U2695 ( .A(n4904), .Y(n4906) );
  AND2X2 U2696 ( .A(n8167), .B(n8165), .Y(n3290) );
  AND3X4 U2697 ( .A(n6143), .B(n4169), .C(n4168), .Y(n3295) );
  BUFX12 U2698 ( .A(n4969), .Y(n4973) );
  NAND2X2 U2699 ( .A(\i_MIPS/ALUin1[16] ), .B(n6571), .Y(n8144) );
  AND2X4 U2700 ( .A(n4687), .B(n4581), .Y(n4622) );
  AND3X4 U2701 ( .A(n4221), .B(n4222), .C(n6125), .Y(n3297) );
  BUFX4 U2702 ( .A(n9117), .Y(n4899) );
  XOR2X1 U2703 ( .A(n9365), .B(ICACHE_addr[16]), .Y(n10944) );
  BUFX8 U2704 ( .A(n4691), .Y(n4827) );
  CLKBUFX8 U2705 ( .A(n11201), .Y(n5475) );
  AND2X6 U2706 ( .A(n8718), .B(n7359), .Y(n3302) );
  AND2X2 U2707 ( .A(n4687), .B(n4654), .Y(n4624) );
  INVX3 U2708 ( .A(n11024), .Y(n10954) );
  AND2X2 U2709 ( .A(n4658), .B(n4655), .Y(n4621) );
  NAND2X1 U2710 ( .A(n4669), .B(n4783), .Y(n10681) );
  CLKINVX1 U2711 ( .A(net102095), .Y(net102371) );
  BUFX4 U2712 ( .A(net102371), .Y(net113455) );
  AND3X4 U2713 ( .A(n4202), .B(n4203), .C(n6116), .Y(n3303) );
  AND2X4 U2714 ( .A(net102565), .B(net140423), .Y(n3304) );
  CLKBUFX3 U2715 ( .A(n9115), .Y(n4890) );
  AND2X2 U2716 ( .A(n4652), .B(n4584), .Y(n4629) );
  AND2X2 U2717 ( .A(n4657), .B(n4584), .Y(n4628) );
  AND3X8 U2718 ( .A(n3802), .B(n3803), .C(net105737), .Y(n3317) );
  CLKBUFX8 U2719 ( .A(net100087), .Y(net112601) );
  CLKAND2X6 U2720 ( .A(n8559), .B(n8557), .Y(n3319) );
  BUFX12 U2721 ( .A(n4627), .Y(n4814) );
  NAND2X2 U2722 ( .A(\i_MIPS/ALUin1[23] ), .B(n6588), .Y(n8897) );
  OAI211X2 U2723 ( .A0(n8690), .A1(n8689), .B0(net102344), .C0(n3709), .Y(
        net99537) );
  NAND2X4 U2724 ( .A(n4500), .B(n4655), .Y(n4483) );
  BUFX2 U2725 ( .A(n4483), .Y(n4910) );
  INVX3 U2726 ( .A(n9223), .Y(n9116) );
  NAND4X4 U2727 ( .A(n6031), .B(n6030), .C(n6029), .D(n6028), .Y(n11374) );
  NAND3X2 U2728 ( .A(n8514), .B(n8516), .C(n8513), .Y(n3320) );
  BUFX4 U2729 ( .A(n9313), .Y(n4995) );
  BUFX4 U2730 ( .A(n4995), .Y(n4993) );
  CLKBUFX3 U2731 ( .A(net112705), .Y(net112703) );
  AND2X2 U2732 ( .A(n4658), .B(n4581), .Y(n4620) );
  CLKBUFX3 U2733 ( .A(n4620), .Y(n4869) );
  CLKBUFX3 U2734 ( .A(n4620), .Y(n4872) );
  BUFX4 U2735 ( .A(n9314), .Y(n4999) );
  CLKINVX1 U2736 ( .A(n8717), .Y(n8734) );
  NAND2X2 U2737 ( .A(n6238), .B(\i_MIPS/n368 ), .Y(n8717) );
  BUFX4 U2738 ( .A(net112187), .Y(net112137) );
  AND2X2 U2739 ( .A(n11168), .B(mem_ready_D), .Y(n3321) );
  INVX3 U2740 ( .A(net99447), .Y(net105285) );
  NAND4X4 U2741 ( .A(n3797), .B(n7715), .C(n7716), .D(n7717), .Y(net99313) );
  BUFX8 U2742 ( .A(net112515), .Y(net112511) );
  INVX3 U2743 ( .A(n6094), .Y(n10655) );
  INVX16 U2744 ( .A(n4492), .Y(DCACHE_addr[27]) );
  INVX16 U2745 ( .A(n4746), .Y(DCACHE_addr[17]) );
  CLKBUFX3 U2746 ( .A(n5143), .Y(n5113) );
  CLKBUFX3 U2747 ( .A(n5406), .Y(n5375) );
  CLKBUFX3 U2748 ( .A(n5187), .Y(n5155) );
  INVX3 U2749 ( .A(n3791), .Y(n3820) );
  BUFX4 U2750 ( .A(n3753), .Y(net112269) );
  BUFX2 U2751 ( .A(n3753), .Y(net112271) );
  OR2X2 U2752 ( .A(net112231), .B(n2795), .Y(n4168) );
  BUFX4 U2753 ( .A(net110217), .Y(net110225) );
  AO21X2 U2754 ( .A0(net99382), .A1(net99383), .B0(net113075), .Y(net99364) );
  CLKBUFX8 U2755 ( .A(net112377), .Y(net112351) );
  CLKXOR2X1 U2756 ( .A(n9621), .B(n3637), .Y(n11068) );
  NAND2X4 U2757 ( .A(n4802), .B(n5592), .Y(n7869) );
  NAND2X1 U2758 ( .A(n3671), .B(net113087), .Y(net100038) );
  CLKINVX1 U2759 ( .A(n11390), .Y(n10857) );
  NAND2X1 U2760 ( .A(n12960), .B(net113087), .Y(net99334) );
  CLKAND2X12 U2761 ( .A(net113606), .B(n11484), .Y(mem_wdata_D[97]) );
  CLKAND2X12 U2762 ( .A(net113606), .B(n11458), .Y(mem_wdata_D[71]) );
  CLKAND2X12 U2763 ( .A(DCACHE_addr[2]), .B(n11516), .Y(mem_addr_D[4]) );
  CLKAND2X12 U2764 ( .A(n3672), .B(n11516), .Y(mem_addr_D[5]) );
  BUFX12 U2765 ( .A(net138398), .Y(net113537) );
  NAND2X2 U2766 ( .A(\i_MIPS/n334 ), .B(\i_MIPS/n310 ), .Y(n11168) );
  OA22X2 U2767 ( .A0(n11058), .A1(net140280), .B0(net98430), .B1(n11057), .Y(
        n11055) );
  XOR2X1 U2768 ( .A(n160), .B(n3692), .Y(n11057) );
  AO22X2 U2769 ( .A0(n115), .A1(ICACHE_addr[22]), .B0(n5463), .B1(n11381), .Y(
        n10990) );
  AO22X2 U2770 ( .A0(n113), .A1(ICACHE_addr[17]), .B0(n5463), .B1(n11376), .Y(
        n11157) );
  BUFX12 U2771 ( .A(net109185), .Y(net109179) );
  AO21X2 U2772 ( .A0(net99502), .A1(net99503), .B0(net113079), .Y(net99475) );
  NAND2X1 U2773 ( .A(n12941), .B(net113087), .Y(net99502) );
  NAND2X1 U2774 ( .A(n9156), .B(n8902), .Y(n8929) );
  NAND2X1 U2775 ( .A(\i_MIPS/ALUin1[24] ), .B(n6589), .Y(n8902) );
  CLKINVX1 U2776 ( .A(n284), .Y(n3508) );
  AO21X2 U2777 ( .A0(net99581), .A1(net99582), .B0(net113077), .Y(net99815) );
  NAND2X1 U2778 ( .A(n12956), .B(net113087), .Y(net99581) );
  NAND2X1 U2779 ( .A(n12942), .B(\i_MIPS/n336 ), .Y(net99969) );
  INVX3 U2780 ( .A(net112671), .Y(net112643) );
  CLKINVX1 U2781 ( .A(net98449), .Y(n3849) );
  NAND2X1 U2782 ( .A(n12958), .B(net113087), .Y(net99014) );
  NAND2X1 U2783 ( .A(n11223), .B(\i_MIPS/n341 ), .Y(n9277) );
  INVX3 U2784 ( .A(n3509), .Y(n3510) );
  INVX3 U2785 ( .A(n3511), .Y(n3512) );
  AO22X2 U2786 ( .A0(n115), .A1(ICACHE_addr[25]), .B0(n5463), .B1(n11384), .Y(
        n10983) );
  AO22X2 U2787 ( .A0(n114), .A1(n3647), .B0(n5463), .B1(n11365), .Y(n10995) );
  INVX3 U2788 ( .A(n3513), .Y(n3514) );
  AO22X2 U2789 ( .A0(n114), .A1(ICACHE_addr[12]), .B0(n5463), .B1(n3639), .Y(
        n10981) );
  AO22X2 U2790 ( .A0(n115), .A1(ICACHE_addr[5]), .B0(n5463), .B1(n11364), .Y(
        n10978) );
  AO22X2 U2791 ( .A0(n114), .A1(ICACHE_addr[23]), .B0(n5463), .B1(n11382), .Y(
        n10992) );
  AO22X2 U2792 ( .A0(n114), .A1(ICACHE_addr[27]), .B0(n5463), .B1(n11386), .Y(
        n10991) );
  CLKINVX1 U2793 ( .A(n5493), .Y(n3567) );
  CLKINVX1 U2794 ( .A(n11350), .Y(n3997) );
  CLKINVX1 U2795 ( .A(n11346), .Y(n4000) );
  AO22X2 U2796 ( .A0(mem_rdata_I[116]), .A1(n113), .B0(n5468), .B1(n11346), 
        .Y(n10007) );
  CLKMX2X2 U2797 ( .A(\D_cache/cache[0][14] ), .B(n10437), .S0(net112627), .Y(
        \D_cache/n1684 ) );
  CLKINVX1 U2798 ( .A(n3515), .Y(n3516) );
  BUFX16 U2799 ( .A(n12947), .Y(DCACHE_addr[21]) );
  NAND2X1 U2800 ( .A(DCACHE_addr[29]), .B(\i_MIPS/n336 ), .Y(n9932) );
  BUFX16 U2801 ( .A(n12939), .Y(DCACHE_addr[29]) );
  INVX3 U2802 ( .A(n5420), .Y(n5418) );
  CLKAND2X12 U2803 ( .A(n3692), .B(n11362), .Y(mem_addr_I[5]) );
  CLKAND2X12 U2804 ( .A(net113916), .B(n11436), .Y(mem_wdata_D[48]) );
  CLKAND2X12 U2805 ( .A(net113916), .B(n11471), .Y(mem_wdata_D[84]) );
  CLKAND2X12 U2806 ( .A(net109183), .B(n11390), .Y(mem_wdata_D[0]) );
  CLKAND2X12 U2807 ( .A(n4794), .B(n11230), .Y(mem_wdata_I[0]) );
  CLKAND2X12 U2808 ( .A(n4795), .B(n11281), .Y(mem_wdata_I[51]) );
  CLKAND2X12 U2809 ( .A(n4796), .B(n11278), .Y(mem_wdata_I[48]) );
  CLKAND2X12 U2810 ( .A(n4794), .B(n11280), .Y(mem_wdata_I[50]) );
  CLKAND2X12 U2811 ( .A(net109183), .B(net98185), .Y(mem_wdata_D[6]) );
  CLKAND2X12 U2812 ( .A(net109183), .B(n11399), .Y(mem_wdata_D[10]) );
  CLKAND2X12 U2813 ( .A(net109183), .B(n11417), .Y(mem_wdata_D[28]) );
  CLKAND2X12 U2814 ( .A(net109183), .B(n11402), .Y(mem_wdata_D[13]) );
  CLKAND2X12 U2815 ( .A(net109183), .B(n11425), .Y(mem_wdata_D[36]) );
  CLKAND2X12 U2816 ( .A(net109183), .B(n11421), .Y(mem_wdata_D[32]) );
  CLKAND2X12 U2817 ( .A(net109183), .B(n11397), .Y(mem_wdata_D[8]) );
  CLKBUFX3 U2818 ( .A(net109185), .Y(net109183) );
  CLKAND2X12 U2819 ( .A(n4794), .B(n11355), .Y(mem_wdata_I[125]) );
  INVX12 U2820 ( .A(n1803), .Y(mem_wdata_I[124]) );
  CLKAND2X12 U2821 ( .A(n4794), .B(n11331), .Y(mem_wdata_I[101]) );
  CLKAND2X12 U2822 ( .A(net113916), .B(n11503), .Y(mem_wdata_D[117]) );
  CLKAND2X12 U2823 ( .A(net113916), .B(n11507), .Y(mem_wdata_D[121]) );
  INVX3 U2824 ( .A(n5421), .Y(n5417) );
  MXI2X2 U2825 ( .A(n10445), .B(n10444), .S0(n5495), .Y(n10446) );
  MXI2X1 U2826 ( .A(n10456), .B(n10455), .S0(n5495), .Y(n10457) );
  MXI2X1 U2827 ( .A(n10469), .B(n10468), .S0(n5495), .Y(n10470) );
  MXI2X1 U2828 ( .A(n10475), .B(n10474), .S0(n5495), .Y(n10476) );
  MXI2X1 U2829 ( .A(n10466), .B(n10465), .S0(n5495), .Y(n10467) );
  MXI2X1 U2830 ( .A(n10453), .B(n10452), .S0(n5495), .Y(n10454) );
  MXI2X1 U2831 ( .A(n10459), .B(n10458), .S0(n5495), .Y(n10460) );
  MXI2X1 U2832 ( .A(n10463), .B(n10462), .S0(n5495), .Y(n10464) );
  MXI2X1 U2833 ( .A(n10472), .B(n10471), .S0(n5495), .Y(n10473) );
  MXI2X1 U2834 ( .A(n10478), .B(n10477), .S0(n5495), .Y(n10479) );
  CLKAND2X12 U2835 ( .A(n3637), .B(n11362), .Y(mem_addr_I[6]) );
  CLKAND2X12 U2836 ( .A(net109181), .B(n11472), .Y(mem_wdata_D[85]) );
  CLKAND2X12 U2837 ( .A(n4005), .B(n11362), .Y(mem_addr_I[4]) );
  NAND2X1 U2838 ( .A(n11361), .B(n11363), .Y(n11362) );
  CLKAND2X12 U2839 ( .A(net113608), .B(n11446), .Y(mem_wdata_D[58]) );
  BUFX12 U2840 ( .A(n11547), .Y(mem_write_I) );
  INVX3 U2841 ( .A(net100087), .Y(net112541) );
  INVX3 U2842 ( .A(net111949), .Y(net111877) );
  CLKAND2X12 U2843 ( .A(DCACHE_addr[4]), .B(n11516), .Y(mem_addr_D[6]) );
  INVX16 U2844 ( .A(net108204), .Y(DCACHE_addr[4]) );
  NAND2BX4 U2845 ( .AN(n5452), .B(n11327), .Y(n9602) );
  CLKBUFX2 U2846 ( .A(net104352), .Y(n3520) );
  NAND3X4 U2847 ( .A(n8426), .B(n4516), .C(n170), .Y(n8336) );
  NAND2X4 U2848 ( .A(net103061), .B(n3809), .Y(n3521) );
  NAND2X6 U2849 ( .A(n3522), .B(n3810), .Y(net99531) );
  INVX6 U2850 ( .A(n3521), .Y(n3522) );
  OR2X4 U2851 ( .A(net103059), .B(net112707), .Y(n3809) );
  NAND3X1 U2852 ( .A(n3585), .B(n3586), .C(net104185), .Y(n3523) );
  INVX4 U2853 ( .A(n3524), .Y(n3525) );
  NOR3BX4 U2854 ( .AN(n3708), .B(n3526), .C(n4413), .Y(n6215) );
  NAND2X1 U2855 ( .A(n8334), .B(n8333), .Y(n8344) );
  INVX4 U2856 ( .A(n10964), .Y(n10321) );
  CLKBUFX3 U2857 ( .A(n5201), .Y(n5205) );
  NAND4X4 U2858 ( .A(n8740), .B(n8741), .C(n8739), .D(n8738), .Y(net99078) );
  AND2X8 U2859 ( .A(n4419), .B(n4418), .Y(n3788) );
  INVX16 U2860 ( .A(net100095), .Y(net100093) );
  INVX3 U2861 ( .A(n6250), .Y(n3527) );
  INVX12 U2862 ( .A(n6249), .Y(n6250) );
  OA22X1 U2863 ( .A0(n5264), .A1(n1232), .B0(n5219), .B1(n2837), .Y(n9939) );
  XOR2X4 U2864 ( .A(net98915), .B(net104829), .Y(n4075) );
  AND2X8 U2865 ( .A(n3872), .B(net99410), .Y(n4533) );
  AO22X1 U2866 ( .A0(n113), .A1(ICACHE_addr[14]), .B0(n5463), .B1(n11373), .Y(
        n10982) );
  AND3XL U2867 ( .A(n3964), .B(n9553), .C(n9555), .Y(n9342) );
  NAND2X4 U2868 ( .A(n3533), .B(n9020), .Y(n3528) );
  AND2X2 U2869 ( .A(n6366), .B(n3599), .Y(n3843) );
  OA22X4 U2870 ( .A0(net112449), .A1(n1935), .B0(net112325), .B1(n354), .Y(
        n6116) );
  AND2X8 U2871 ( .A(n3789), .B(\i_MIPS/n367 ), .Y(n3529) );
  NAND2X1 U2872 ( .A(n4793), .B(n9328), .Y(n10974) );
  AO22XL U2873 ( .A0(ICACHE_addr[28]), .A1(mem_read_I), .B0(n4794), .B1(n11387), .Y(n12824) );
  AO22X1 U2874 ( .A0(n115), .A1(ICACHE_addr[28]), .B0(n5463), .B1(n11387), .Y(
        n10979) );
  INVX2 U2875 ( .A(n9001), .Y(n9003) );
  NAND2X4 U2876 ( .A(n4508), .B(n10297), .Y(n10949) );
  INVX3 U2877 ( .A(n11011), .Y(n10297) );
  OA22X2 U2878 ( .A0(n5430), .A1(n908), .B0(n5386), .B1(n2425), .Y(n9368) );
  NAND2X6 U2879 ( .A(n4157), .B(n10937), .Y(n10941) );
  NAND3X6 U2880 ( .A(n4026), .B(n6140), .C(n6141), .Y(n6169) );
  OR2X2 U2881 ( .A(net112693), .B(n2018), .Y(n4204) );
  AND2X4 U2882 ( .A(n6231), .B(\i_MIPS/n361 ), .Y(n3773) );
  AND3X8 U2883 ( .A(n9022), .B(n9021), .C(n9023), .Y(n3533) );
  INVX3 U2884 ( .A(n8521), .Y(n6618) );
  NAND2X6 U2885 ( .A(\i_MIPS/ALUin1[20] ), .B(n6578), .Y(n8521) );
  NAND2X6 U2886 ( .A(n4194), .B(n4195), .Y(n6578) );
  OA22X1 U2887 ( .A0(\i_MIPS/n362 ), .A1(n4811), .B0(\i_MIPS/n361 ), .B1(n4805), .Y(n6949) );
  OA22X2 U2888 ( .A0(\i_MIPS/n368 ), .A1(n4812), .B0(\i_MIPS/n367 ), .B1(n4805), .Y(n6257) );
  NAND2X6 U2889 ( .A(n3832), .B(n1877), .Y(n4210) );
  OAI221X1 U2890 ( .A0(\i_MIPS/Register/register[18][10] ), .A1(n4945), .B0(
        \i_MIPS/Register/register[26][10] ), .B1(n4942), .C0(n7258), .Y(n7266)
         );
  INVX12 U2891 ( .A(n7704), .Y(n6626) );
  AO22XL U2892 ( .A0(ICACHE_addr[25]), .A1(mem_read_I), .B0(n4796), .B1(n11384), .Y(n12825) );
  CLKINVX3 U2893 ( .A(n5380), .Y(n5368) );
  INVX1 U2894 ( .A(n8649), .Y(n8651) );
  AO22X1 U2895 ( .A0(n9312), .A1(n551), .B0(n4981), .B1(n2054), .Y(n7344) );
  INVX4 U2896 ( .A(n10263), .Y(n10261) );
  INVX3 U2897 ( .A(n3693), .Y(n3692) );
  CLKXOR2X2 U2898 ( .A(n10199), .B(ICACHE_addr[24]), .Y(n10363) );
  NAND2X2 U2899 ( .A(n10361), .B(ICACHE_addr[23]), .Y(n10199) );
  AND2X2 U2900 ( .A(n4555), .B(n8143), .Y(n4518) );
  CLKINVX3 U2901 ( .A(n10487), .Y(n3609) );
  CLKINVX2 U2902 ( .A(n4424), .Y(n3637) );
  CLKAND2X3 U2903 ( .A(n8431), .B(n8333), .Y(n4550) );
  OAI211X2 U2904 ( .A0(n8208), .A1(n8207), .B0(net113439), .C0(net112609), .Y(
        n10447) );
  CLKBUFX2 U2905 ( .A(net112517), .Y(net112505) );
  CLKBUFX2 U2906 ( .A(net112509), .Y(net112425) );
  CLKBUFX8 U2907 ( .A(net112507), .Y(net112453) );
  INVX3 U2908 ( .A(n10328), .Y(n4505) );
  MX2X2 U2909 ( .A(n6851), .B(n7611), .S0(n5590), .Y(n8083) );
  INVX4 U2910 ( .A(n6213), .Y(n3530) );
  CLKINVX3 U2911 ( .A(n3772), .Y(n8070) );
  MX2XL U2912 ( .A(DCACHE_addr[2]), .B(net99447), .S0(n5508), .Y(\i_MIPS/n465 ) );
  OAI221X1 U2913 ( .A0(n4798), .A1(n8806), .B0(n8807), .B1(n3746), .C0(n8805), 
        .Y(n8810) );
  NOR4X4 U2914 ( .A(n8445), .B(n8447), .C(n8446), .D(n8448), .Y(n8453) );
  OA21X4 U2915 ( .A0(n10321), .A1(n4610), .B0(n10324), .Y(net99765) );
  CLKINVX2 U2916 ( .A(n7854), .Y(n3698) );
  CLKINVX8 U2917 ( .A(n6242), .Y(n6239) );
  OAI21X4 U2918 ( .A0(n8527), .A1(n8075), .B0(n8521), .Y(n3556) );
  OAI221XL U2919 ( .A0(\i_MIPS/ID_EX[73] ), .A1(n4434), .B0(\i_MIPS/ID_EX[41] ), .B1(n3826), .C0(\i_MIPS/n371 ), .Y(n4441) );
  NAND2X6 U2920 ( .A(n6584), .B(\i_MIPS/n350 ), .Y(n8095) );
  CLKINVX12 U2921 ( .A(n6660), .Y(n6444) );
  INVXL U2922 ( .A(n3658), .Y(n3659) );
  INVX4 U2923 ( .A(net99432), .Y(n3658) );
  BUFX8 U2924 ( .A(n8821), .Y(n3599) );
  AND3X8 U2925 ( .A(n3686), .B(n4171), .C(n4067), .Y(n4587) );
  OAI221X2 U2926 ( .A0(net107236), .A1(net112707), .B0(net107237), .B1(
        net112723), .C0(net107238), .Y(net99009) );
  OA22X2 U2927 ( .A0(n8726), .A1(n8434), .B0(n4519), .B1(n141), .Y(n6859) );
  AND2X4 U2928 ( .A(n6235), .B(\i_MIPS/n369 ), .Y(n3759) );
  NAND4X4 U2929 ( .A(n4457), .B(n4458), .C(n5968), .D(n5967), .Y(n11383) );
  AO22X2 U2930 ( .A0(n113), .A1(ICACHE_addr[16]), .B0(n5463), .B1(n3564), .Y(
        n10976) );
  OR2X2 U2931 ( .A(net112663), .B(n2796), .Y(n4181) );
  NAND2BX2 U2932 ( .AN(net112561), .B(\D_cache/cache[1][138] ), .Y(n4182) );
  BUFX16 U2933 ( .A(net112691), .Y(net112663) );
  MXI2X1 U2934 ( .A(n10769), .B(n10768), .S0(n5490), .Y(n10770) );
  AOI222X4 U2935 ( .A0(n5480), .A1(n11460), .B0(mem_rdata_D[73]), .B1(n116), 
        .C0(n12988), .C1(n5477), .Y(n10769) );
  NAND2X2 U2936 ( .A(\i_MIPS/n275 ), .B(n4199), .Y(n4200) );
  INVX6 U2937 ( .A(n4199), .Y(n3577) );
  NAND2X2 U2938 ( .A(\i_MIPS/ID_EX[49] ), .B(n4199), .Y(n4435) );
  NAND2X6 U2939 ( .A(n4217), .B(n4218), .Y(n6571) );
  NAND2X4 U2940 ( .A(\i_MIPS/n277 ), .B(n3770), .Y(n4217) );
  CLKBUFX3 U2941 ( .A(n5408), .Y(n5403) );
  BUFX8 U2942 ( .A(n11139), .Y(n5408) );
  OA22X2 U2943 ( .A0(n8730), .A1(n8729), .B0(n8728), .B1(n8727), .Y(n8739) );
  MX2X1 U2944 ( .A(n7451), .B(n7106), .S0(n5589), .Y(n8730) );
  NAND4X1 U2945 ( .A(n3692), .B(n4005), .C(n3647), .D(n3649), .Y(n9333) );
  OR2X8 U2946 ( .A(net104184), .B(net112721), .Y(n3586) );
  NAND2X2 U2947 ( .A(n4616), .B(n4694), .Y(n9338) );
  INVX16 U2948 ( .A(n5593), .Y(n3770) );
  INVX4 U2949 ( .A(n9017), .Y(n3561) );
  OA22X2 U2950 ( .A0(net112511), .A1(n449), .B0(net112379), .B1(n3291), .Y(
        n6131) );
  AOI221X1 U2951 ( .A0(n9259), .A1(n3558), .B0(n7185), .B1(n9258), .C0(n4800), 
        .Y(n7210) );
  NAND3X6 U2952 ( .A(net98965), .B(net98966), .C(net98964), .Y(n4128) );
  CLKINVX6 U2953 ( .A(n10948), .Y(n10293) );
  INVX16 U2954 ( .A(n4425), .Y(n9428) );
  NAND3X8 U2955 ( .A(net99476), .B(net99477), .C(net99475), .Y(n4129) );
  NAND3X8 U2956 ( .A(n3690), .B(n3691), .C(net106566), .Y(net99464) );
  OA21X4 U2957 ( .A0(n3559), .A1(n4609), .B0(n11015), .Y(n11016) );
  OR2X6 U2958 ( .A(n9176), .B(n9175), .Y(n3534) );
  OR2X8 U2959 ( .A(n9174), .B(n9173), .Y(n3535) );
  OR2X2 U2960 ( .A(n3552), .B(net110241), .Y(n3536) );
  OR2X4 U2961 ( .A(n10732), .B(n10390), .Y(n3537) );
  OR2X1 U2962 ( .A(\i_MIPS/PC/n30 ), .B(net110213), .Y(n3538) );
  OR2X8 U2963 ( .A(n9333), .B(n9332), .Y(n10204) );
  NAND2X6 U2964 ( .A(n4809), .B(\i_MIPS/ALUin1[13] ), .Y(n6359) );
  MX2XL U2965 ( .A(n3489), .B(n2), .S0(n5509), .Y(\i_MIPS/n403 ) );
  CLKAND2X3 U2966 ( .A(n7199), .B(n8818), .Y(n3580) );
  AND2X6 U2967 ( .A(n3727), .B(n6660), .Y(n3587) );
  NAND2X8 U2968 ( .A(n6444), .B(n3727), .Y(n9264) );
  INVX1 U2969 ( .A(n10866), .Y(n9630) );
  NAND2BX2 U2970 ( .AN(n9624), .B(n10206), .Y(n9625) );
  OR2X6 U2971 ( .A(net104524), .B(net112709), .Y(n3539) );
  OR2X6 U2972 ( .A(net104525), .B(net112721), .Y(n3540) );
  CLKMX2X2 U2973 ( .A(n7845), .B(n7844), .S0(net108963), .Y(net104524) );
  NOR2X1 U2974 ( .A(\i_MIPS/PC/n9 ), .B(net110215), .Y(n3541) );
  NOR2X1 U2975 ( .A(n4329), .B(\i_MIPS/PC/n9 ), .Y(n4345) );
  OR2X1 U2976 ( .A(n10872), .B(n10871), .Y(n4155) );
  OA22X2 U2977 ( .A0(n10872), .A1(net140280), .B0(net98430), .B1(n10871), .Y(
        n10868) );
  NAND3BX2 U2978 ( .AN(n3541), .B(n3655), .C(n3656), .Y(n10869) );
  OR2X1 U2979 ( .A(n3646), .B(net110215), .Y(n3542) );
  INVX1 U2980 ( .A(n11188), .Y(n3545) );
  CLKINVX1 U2981 ( .A(n3545), .Y(n3546) );
  NAND3BX4 U2982 ( .AN(n3672), .B(net113540), .C(net113532), .Y(net100081) );
  OR2X2 U2983 ( .A(net112137), .B(n2797), .Y(n4169) );
  MXI2X1 U2984 ( .A(n10684), .B(n10683), .S0(n5491), .Y(n10685) );
  AOI222X1 U2985 ( .A0(n5475), .A1(n11512), .B0(mem_rdata_D[126]), .B1(n116), 
        .C0(n12967), .C1(n5473), .Y(n10684) );
  OA22X2 U2986 ( .A0(n4519), .A1(n9004), .B0(n141), .B1(n8433), .Y(n7701) );
  OA22X2 U2987 ( .A0(n8087), .A1(n8534), .B0(n8086), .B1(n141), .Y(n8092) );
  MX2X1 U2988 ( .A(\I_cache/cache[6][41] ), .B(n9635), .S0(n5418), .Y(n12489)
         );
  AND3X4 U2989 ( .A(n4162), .B(n4163), .C(n6145), .Y(n3734) );
  OR2X1 U2990 ( .A(net112663), .B(n3196), .Y(n4162) );
  INVX2 U2991 ( .A(n9174), .Y(n3831) );
  OAI222X4 U2992 ( .A0(n4517), .A1(n7544), .B0(n8659), .B1(n7461), .C0(n8817), 
        .C1(n7451), .Y(n7483) );
  INVXL U2993 ( .A(n4527), .Y(n3551) );
  CLKINVX1 U2994 ( .A(n3551), .Y(n3552) );
  AND2X2 U2995 ( .A(\i_MIPS/n312 ), .B(\i_MIPS/n314 ), .Y(n4584) );
  CLKMX2X2 U2996 ( .A(n8994), .B(n8993), .S0(net108959), .Y(n8996) );
  INVX3 U2997 ( .A(n4629), .Y(n4950) );
  INVX16 U2998 ( .A(n3827), .Y(n6947) );
  NAND2X6 U2999 ( .A(n10897), .B(n10895), .Y(n10265) );
  INVX3 U3000 ( .A(n11146), .Y(n11119) );
  NAND2BXL U3001 ( .AN(n5456), .B(n11256), .Y(n9713) );
  NOR2X4 U3002 ( .A(n3556), .B(n3555), .Y(n3699) );
  AOI2BB1X4 U3003 ( .A0N(\i_MIPS/n359 ), .A1N(n4812), .B0(n6360), .Y(n6361) );
  INVX6 U3004 ( .A(n6359), .Y(n6360) );
  OR2X2 U3005 ( .A(net112229), .B(n2019), .Y(n4223) );
  NAND2X8 U3006 ( .A(n3304), .B(net140424), .Y(net99354) );
  OR2X2 U3007 ( .A(net112663), .B(n2798), .Y(n4164) );
  NAND2X6 U3008 ( .A(net99504), .B(net113039), .Y(net99477) );
  NAND4BX2 U3009 ( .AN(n7439), .B(n7438), .C(n7437), .D(n7436), .Y(n7450) );
  OA22X4 U3010 ( .A0(n3547), .A1(net104563), .B0(net102087), .B1(n3554), .Y(
        n3553) );
  OR2X4 U3011 ( .A(n8996), .B(net112707), .Y(net140423) );
  CLKINVX4 U3012 ( .A(n7191), .Y(n7185) );
  NAND2X8 U3013 ( .A(n4443), .B(n8432), .Y(n8359) );
  NAND3X6 U3014 ( .A(n4442), .B(n9156), .C(n8431), .Y(n4443) );
  INVX4 U3015 ( .A(n7192), .Y(n3558) );
  CLKINVX6 U3016 ( .A(n7190), .Y(n7192) );
  BUFX4 U3017 ( .A(net112509), .Y(net112443) );
  NAND3X6 U3018 ( .A(n4106), .B(n4105), .C(n4121), .Y(n4087) );
  AOI2BB2X4 U3019 ( .B0(n3560), .B1(\D_cache/cache[2][148] ), .A0N(net112385), 
        .A1N(n1895), .Y(n6087) );
  AND3X4 U3020 ( .A(n8919), .B(n8918), .C(n8917), .Y(n8933) );
  INVX12 U3021 ( .A(n4437), .Y(n6243) );
  OR2X8 U3022 ( .A(net103391), .B(net112721), .Y(n3713) );
  MXI2X1 U3023 ( .A(n10570), .B(n10569), .S0(n5493), .Y(n10571) );
  NOR2X8 U3024 ( .A(n11014), .B(n3833), .Y(n3559) );
  INVX20 U3025 ( .A(n3559), .Y(n11117) );
  NAND4BBX4 U3026 ( .AN(n8332), .BN(n8253), .C(n8327), .D(n4801), .Y(n8330) );
  MXI2X1 U3027 ( .A(n10560), .B(n10559), .S0(n5493), .Y(n10561) );
  AOI222X4 U3028 ( .A0(n5480), .A1(n11474), .B0(mem_rdata_D[87]), .B1(n117), 
        .C0(n12974), .C1(n5477), .Y(n10560) );
  OA22X4 U3029 ( .A0(net112449), .A1(n1936), .B0(net112325), .B1(n355), .Y(
        n6119) );
  AOI2BB2X4 U3030 ( .B0(n3560), .B1(\D_cache/cache[2][144] ), .A0N(net112381), 
        .A1N(n1896), .Y(n6059) );
  CLKAND2X4 U3031 ( .A(net112609), .B(n11389), .Y(n4778) );
  INVX3 U3032 ( .A(n8656), .Y(n8664) );
  NOR2X4 U3033 ( .A(n4188), .B(n8662), .Y(n8669) );
  AND3X6 U3034 ( .A(net108204), .B(net113540), .C(n3672), .Y(n3822) );
  AND3X8 U3035 ( .A(n3751), .B(n3671), .C(net113532), .Y(n3730) );
  BUFX20 U3036 ( .A(n3839), .Y(net113532) );
  BUFX4 U3037 ( .A(net113047), .Y(net113041) );
  NAND3X4 U3038 ( .A(n4567), .B(n6444), .C(n6263), .Y(n6260) );
  NAND2X8 U3039 ( .A(n8260), .B(n4578), .Y(n8537) );
  NAND4BX2 U3040 ( .AN(n7448), .B(n7447), .C(n7446), .D(n7445), .Y(n7449) );
  NAND2BX1 U3041 ( .AN(n5452), .B(n11338), .Y(n10104) );
  NAND2BX2 U3042 ( .AN(n5452), .B(n11332), .Y(n9838) );
  NAND2BX2 U3043 ( .AN(n5452), .B(n11340), .Y(n10001) );
  NAND2BX2 U3044 ( .AN(n5452), .B(n11334), .Y(n9685) );
  CLKINVX6 U3045 ( .A(n3751), .Y(n3752) );
  OAI31X2 U3046 ( .A0(n8655), .A1(n8430), .A2(n9153), .B0(n4563), .Y(n9017) );
  NAND2X1 U3047 ( .A(n9451), .B(ICACHE_addr[5]), .Y(n9452) );
  BUFX4 U3048 ( .A(n4934), .Y(n4937) );
  NAND3BX2 U3049 ( .AN(n11056), .B(n11055), .C(n11054), .Y(\i_MIPS/PC/n39 ) );
  NAND3BX2 U3050 ( .AN(n11199), .B(n11198), .C(n11197), .Y(\i_MIPS/PC/n38 ) );
  INVXL U3051 ( .A(n11375), .Y(n3563) );
  CLKINVX1 U3052 ( .A(n3563), .Y(n3564) );
  AND2X1 U3053 ( .A(net134107), .B(net100042), .Y(n4562) );
  AOI211X2 U3054 ( .A0(n9140), .A1(n8541), .B0(n7369), .C0(n7368), .Y(n7370)
         );
  BUFX6 U3055 ( .A(n5232), .Y(n5228) );
  CLKBUFX4 U3056 ( .A(n5232), .Y(n5227) );
  INVX1 U3057 ( .A(n9571), .Y(n5956) );
  BUFX16 U3058 ( .A(n5276), .Y(n5316) );
  XOR2X4 U3059 ( .A(n6126), .B(n4756), .Y(n6127) );
  OAI22X2 U3060 ( .A0(n5163), .A1(n3200), .B0(n5120), .B1(n323), .Y(n4447) );
  BUFX8 U3061 ( .A(n5187), .Y(n5163) );
  AO21X4 U3062 ( .A0(n10387), .A1(net98880), .B0(n10386), .Y(n3568) );
  NOR2X4 U3063 ( .A(n3568), .B(net113592), .Y(n10388) );
  OR2X1 U3064 ( .A(\i_MIPS/PC/n32 ), .B(net110213), .Y(n3571) );
  OAI211X2 U3065 ( .A0(n11225), .A1(n9160), .B0(n9158), .C0(n9159), .Y(n3574)
         );
  INVX4 U3066 ( .A(n9327), .Y(n10387) );
  MXI2X2 U3067 ( .A(n10170), .B(net100023), .S0(n5497), .Y(n10171) );
  NAND2BX1 U3068 ( .AN(n9345), .B(n9346), .Y(n9344) );
  NAND4X4 U3069 ( .A(n9343), .B(n9342), .C(n9341), .D(n9340), .Y(n9346) );
  INVX16 U3070 ( .A(net99850), .Y(net98880) );
  NAND3X6 U3071 ( .A(n3673), .B(n4423), .C(n4005), .Y(n11139) );
  BUFX8 U3072 ( .A(net114092), .Y(net109185) );
  OR2X2 U3073 ( .A(net112663), .B(n2799), .Y(n4161) );
  MXI2X1 U3074 ( .A(n10190), .B(n10189), .S0(n5497), .Y(n10191) );
  AOI222X4 U3075 ( .A0(n5479), .A1(n11466), .B0(mem_rdata_D[79]), .B1(n117), 
        .C0(n12982), .C1(n5476), .Y(n10190) );
  OAI22X2 U3076 ( .A0(net112499), .A1(n313), .B0(net112319), .B1(n1888), .Y(
        n3738) );
  MX2X1 U3077 ( .A(\D_cache/cache[7][53] ), .B(n4272), .S0(net111877), .Y(
        \D_cache/n1365 ) );
  CLKBUFX3 U3078 ( .A(n5449), .Y(n5424) );
  CLKBUFX2 U3079 ( .A(n6450), .Y(n3575) );
  NAND4BX2 U3080 ( .AN(n8708), .B(n8707), .C(n8706), .D(n8705), .Y(n8709) );
  NOR4X2 U3081 ( .A(n8704), .B(n8703), .C(n8702), .D(n8701), .Y(n8705) );
  AO22XL U3082 ( .A0(n4974), .A1(n188), .B0(n4967), .B1(n2265), .Y(n8704) );
  AO22X1 U3083 ( .A0(n9310), .A1(n647), .B0(n4976), .B1(n2168), .Y(n8703) );
  MXI2X1 U3084 ( .A(n10396), .B(n10395), .S0(n5497), .Y(n10397) );
  AOI222X4 U3085 ( .A0(n5474), .A1(n11510), .B0(mem_rdata_D[124]), .B1(n116), 
        .C0(n12969), .C1(n5472), .Y(n10396) );
  MXI2X1 U3086 ( .A(n10609), .B(n10608), .S0(n5492), .Y(n10610) );
  OAI31X2 U3087 ( .A0(n6212), .A1(\i_MIPS/ID_EX[73] ), .A2(n6211), .B0(n6210), 
        .Y(n6448) );
  NAND2X6 U3088 ( .A(n4131), .B(n4100), .Y(n4133) );
  OA22X1 U3089 ( .A0(net112463), .A1(n1233), .B0(net112339), .B1(n2838), .Y(
        n7061) );
  INVX1 U3090 ( .A(n7200), .Y(n3576) );
  BUFX2 U3091 ( .A(n9116), .Y(n4897) );
  NAND3BX2 U3092 ( .AN(n11072), .B(n11071), .C(n11070), .Y(\i_MIPS/PC/n40 ) );
  NAND3X8 U3093 ( .A(n9557), .B(n9556), .C(n3257), .Y(n9559) );
  CLKINVX3 U3094 ( .A(n5424), .Y(n5412) );
  AND3X2 U3095 ( .A(n4640), .B(n9570), .C(n4661), .Y(n9343) );
  OA22X2 U3096 ( .A0(n10930), .A1(net140281), .B0(net98430), .B1(n10929), .Y(
        n10932) );
  BUFX4 U3097 ( .A(n4487), .Y(n4938) );
  MX2X1 U3098 ( .A(n6855), .B(n6852), .S0(n5589), .Y(n7290) );
  MXI2X1 U3099 ( .A(n10481), .B(n10480), .S0(n5495), .Y(n10482) );
  BUFX4 U3100 ( .A(n10482), .Y(n4304) );
  AOI222X4 U3101 ( .A0(net109791), .A1(n11418), .B0(mem_rdata_D[29]), .B1(n116), .C0(n12968), .C1(net109801), .Y(n10481) );
  AO22XL U3102 ( .A0(n9118), .A1(n513), .B0(n4901), .B1(n2266), .Y(n6319) );
  BUFX4 U3103 ( .A(n4483), .Y(n4909) );
  BUFX4 U3104 ( .A(n4918), .Y(n4915) );
  OA22X1 U3105 ( .A0(\i_MIPS/Register/register[22][12] ), .A1(n4909), .B0(
        \i_MIPS/Register/register[30][12] ), .B1(n4906), .Y(n6318) );
  NOR4X1 U3106 ( .A(n7744), .B(n7743), .C(n7742), .D(n7741), .Y(n7755) );
  NOR3X4 U3107 ( .A(n3578), .B(n3579), .C(n3580), .Y(n7201) );
  AND2X2 U3108 ( .A(n7206), .B(n7205), .Y(n3581) );
  AND2X2 U3109 ( .A(n7204), .B(n3636), .Y(n3582) );
  NOR3X4 U3110 ( .A(n3581), .B(n3582), .C(n7203), .Y(n7207) );
  INVX3 U3111 ( .A(n7197), .Y(n8342) );
  CLKINVX1 U3112 ( .A(n8345), .Y(n7199) );
  CLKINVX12 U3113 ( .A(n8728), .Y(n8818) );
  NAND2X8 U3114 ( .A(n3711), .B(n7207), .Y(net99336) );
  AOI22X4 U3115 ( .A0(net113041), .A1(net99039), .B0(net102300), .B1(net105824), .Y(net134109) );
  OAI221X4 U3116 ( .A0(n141), .A1(n8909), .B0(n8911), .B1(n8886), .C0(n4501), 
        .Y(n8170) );
  NAND2X8 U3117 ( .A(n3626), .B(n8517), .Y(n8523) );
  NAND2X2 U3118 ( .A(n3259), .B(n8336), .Y(n8335) );
  CLKINVX12 U3119 ( .A(n9428), .Y(n3673) );
  AOI2BB2X4 U3120 ( .B0(net113167), .B1(n8672), .A0N(net103060), .A1N(
        net104563), .Y(n3583) );
  NAND3XL U3121 ( .A(n3809), .B(n3810), .C(net103061), .Y(n3584) );
  OAI221X2 U3122 ( .A0(net104704), .A1(net112709), .B0(net104705), .B1(
        net112721), .C0(net104706), .Y(net99307) );
  OAI221X2 U3123 ( .A0(\i_MIPS/n349 ), .A1(n4824), .B0(\i_MIPS/n350 ), .B1(
        n4816), .C0(n7023), .Y(n7103) );
  NAND3BXL U3124 ( .AN(n4707), .B(n8912), .C(n9130), .Y(n8918) );
  NAND2X8 U3125 ( .A(n9130), .B(n8348), .Y(n8660) );
  AOI222X1 U3126 ( .A0(n9133), .A1(\i_MIPS/ALU/N303 ), .B0(n9271), .B1(n9132), 
        .C0(n9131), .C1(n9130), .Y(n9134) );
  AND3X8 U3127 ( .A(n6767), .B(n8823), .C(n8717), .Y(n3892) );
  BUFX3 U3128 ( .A(n5450), .Y(n5422) );
  OAI221X1 U3129 ( .A0(\i_MIPS/Register/register[18][4] ), .A1(n4945), .B0(
        \i_MIPS/Register/register[26][4] ), .B1(n4940), .C0(n7420), .Y(n7428)
         );
  NAND2X2 U3130 ( .A(n4724), .B(n10917), .Y(n10920) );
  NAND2BX2 U3131 ( .AN(n5458), .B(n11242), .Y(n10102) );
  AND3X4 U3132 ( .A(n4614), .B(n9556), .C(n9334), .Y(n9341) );
  NAND2X8 U3133 ( .A(n3623), .B(n6936), .Y(n8153) );
  NOR4X2 U3134 ( .A(n7415), .B(n7414), .C(n7413), .D(n7412), .Y(n7416) );
  OA22X2 U3135 ( .A0(\i_MIPS/Register/register[6][4] ), .A1(n4936), .B0(
        \i_MIPS/Register/register[14][4] ), .B1(n4930), .Y(n7411) );
  MX2X1 U3136 ( .A(n9280), .B(n9279), .S0(n3601), .Y(n8824) );
  OR2X4 U3137 ( .A(net104183), .B(net112709), .Y(n3585) );
  NAND3X6 U3138 ( .A(n3585), .B(n3586), .C(net104185), .Y(net99401) );
  AO21X2 U3139 ( .A0(net99406), .A1(net99405), .B0(net112729), .Y(net104185)
         );
  OAI222X2 U3140 ( .A0(n8659), .A1(n8517), .B0(n8727), .B1(n8437), .C0(n7786), 
        .C1(n8805), .Y(n7795) );
  OAI222X2 U3141 ( .A0(n8641), .A1(n9004), .B0(n8725), .B1(n9007), .C0(n141), 
        .C1(n8665), .Y(n7794) );
  INVX12 U3142 ( .A(net110255), .Y(n3602) );
  NAND2X6 U3143 ( .A(n10629), .B(net113039), .Y(n10731) );
  INVXL U3144 ( .A(n10629), .Y(n9211) );
  NAND2X2 U3145 ( .A(n8922), .B(n8332), .Y(n8921) );
  XOR2X4 U3146 ( .A(net99464), .B(n4129), .Y(n4118) );
  AO21X4 U3147 ( .A0(n6452), .A1(n8804), .B0(n7273), .Y(n6460) );
  CLKINVX1 U3148 ( .A(n6453), .Y(n6452) );
  NAND2BX4 U3149 ( .AN(n6478), .B(n3632), .Y(n6470) );
  NOR4X4 U3150 ( .A(n7046), .B(n7045), .C(n7044), .D(n7043), .Y(n7047) );
  INVX20 U3151 ( .A(n3587), .Y(n9262) );
  BUFX6 U3152 ( .A(n9259), .Y(n4925) );
  INVXL U3153 ( .A(n8802), .Y(n8715) );
  NAND2X6 U3154 ( .A(n4727), .B(n3621), .Y(n3794) );
  NOR2BX4 U3155 ( .AN(\i_MIPS/IR_ID[21] ), .B(\i_MIPS/n229 ), .Y(n4658) );
  CLKINVX1 U3156 ( .A(n11018), .Y(n11017) );
  NAND3X8 U3157 ( .A(n4196), .B(n4197), .C(n6355), .Y(n7611) );
  NAND2X2 U3158 ( .A(n8266), .B(n8265), .Y(n8267) );
  INVX1 U3159 ( .A(n8546), .Y(n8266) );
  NAND2X4 U3160 ( .A(n6588), .B(\i_MIPS/n348 ), .Y(n8920) );
  OAI221X2 U3161 ( .A0(\i_MIPS/n348 ), .A1(n4811), .B0(\i_MIPS/n349 ), .B1(
        n4803), .C0(n6950), .Y(n7866) );
  INVXL U3162 ( .A(n11383), .Y(n3588) );
  CLKINVX1 U3163 ( .A(n3588), .Y(n3589) );
  INVX1 U3164 ( .A(n5456), .Y(n3590) );
  NAND4X2 U3165 ( .A(n8174), .B(n8173), .C(n8172), .D(n8171), .Y(n8179) );
  AOI21X2 U3166 ( .A0(\i_MIPS/n281 ), .A1(n3827), .B0(\i_MIPS/n279 ), .Y(n6620) );
  CLKAND2X12 U3167 ( .A(\i_MIPS/IR_ID[16] ), .B(\i_MIPS/n314 ), .Y(n4659) );
  BUFX4 U3168 ( .A(n9310), .Y(n4978) );
  CLKMX2X2 U3169 ( .A(net103393), .B(net103394), .S0(net108959), .Y(net103390)
         );
  BUFX4 U3170 ( .A(n4943), .Y(n4947) );
  NAND2X1 U3171 ( .A(n9160), .B(n11224), .Y(n9018) );
  INVX3 U3172 ( .A(n6655), .Y(n6617) );
  MXI2X4 U3173 ( .A(\i_MIPS/ID_EX[69] ), .B(\i_MIPS/ID_EX[101] ), .S0(n3771), 
        .Y(n6655) );
  BUFX8 U3174 ( .A(n5451), .Y(n5448) );
  AOI2BB1X4 U3175 ( .A0N(n6234), .A1N(\i_MIPS/ALUin1[1] ), .B0(\i_MIPS/n371 ), 
        .Y(n3721) );
  AOI33X2 U3176 ( .A0(n9258), .A1(n7034), .A2(n7033), .B0(n9258), .B1(n3508), 
        .B2(n7032), .Y(n7048) );
  INVX1 U3177 ( .A(n7200), .Y(n3591) );
  INVX8 U3178 ( .A(n4809), .Y(n3592) );
  OA22X4 U3179 ( .A0(net104563), .A1(net102745), .B0(net102087), .B1(n3594), 
        .Y(n3593) );
  NAND2XL U3180 ( .A(n6944), .B(n7365), .Y(n3595) );
  AND3X4 U3181 ( .A(n3595), .B(n3596), .C(n3597), .Y(n6268) );
  INVX3 U3182 ( .A(n6368), .Y(n6944) );
  NAND2X4 U3183 ( .A(\i_MIPS/n269 ), .B(n4158), .Y(n4194) );
  NAND4X6 U3184 ( .A(n6959), .B(n6958), .C(n6957), .D(n6956), .Y(net99583) );
  AO22X2 U3185 ( .A0(n9271), .A1(n8343), .B0(n8342), .B1(n9267), .Y(n8358) );
  AOI32XL U3186 ( .A0(n3636), .A1(\i_MIPS/ALUin1[30] ), .A2(n9268), .B0(n9267), 
        .B1(n9266), .Y(n9291) );
  AND2X4 U3187 ( .A(n6233), .B(\i_MIPS/n369 ), .Y(n3601) );
  OAI221X4 U3188 ( .A0(n4798), .A1(n7274), .B0(n4551), .B1(n9262), .C0(n8805), 
        .Y(n7277) );
  OAI221X2 U3189 ( .A0(net102899), .A1(net112707), .B0(net102900), .B1(
        net112721), .C0(net102901), .Y(net100099) );
  NOR2X2 U3190 ( .A(n8664), .B(n2017), .Y(n8662) );
  OAI2BB1X4 U3191 ( .A0N(n7548), .A1N(n7562), .B0(n7550), .Y(n7465) );
  NAND3X8 U3192 ( .A(n7459), .B(n7550), .C(n3302), .Y(n6769) );
  NAND2X6 U3193 ( .A(\i_MIPS/ALUin1[6] ), .B(n3823), .Y(n7550) );
  MXI2X1 U3194 ( .A(n10415), .B(n10414), .S0(n5496), .Y(n10416) );
  AOI222X4 U3195 ( .A0(n5479), .A1(n11477), .B0(mem_rdata_D[90]), .B1(n117), 
        .C0(n12971), .C1(n5476), .Y(n10415) );
  BUFX4 U3196 ( .A(n4910), .Y(n4914) );
  INVXL U3197 ( .A(n3302), .Y(n3603) );
  OR2X1 U3198 ( .A(\i_MIPS/PC/n13 ), .B(net110213), .Y(n3604) );
  OR2X1 U3199 ( .A(n4539), .B(net110243), .Y(n3605) );
  NAND3X2 U3200 ( .A(n3605), .B(n3604), .C(n3606), .Y(n11082) );
  AND2XL U3201 ( .A(net134109), .B(net99019), .Y(n4539) );
  OR2X2 U3202 ( .A(n4536), .B(net110241), .Y(n4173) );
  NAND3BX2 U3203 ( .AN(n10360), .B(n10359), .C(n10358), .Y(\i_MIPS/PC/n60 ) );
  NAND3BX2 U3204 ( .AN(n10973), .B(n10972), .C(n10971), .Y(\i_MIPS/PC/n57 ) );
  INVXL U3205 ( .A(n8713), .Y(n3607) );
  CLKINVX1 U3206 ( .A(n3607), .Y(n3608) );
  INVX4 U3207 ( .A(n6610), .Y(n6607) );
  INVX4 U3208 ( .A(n6250), .Y(n3643) );
  NAND2X4 U3209 ( .A(n6250), .B(\i_MIPS/n359 ), .Y(n6633) );
  AOI2BB1X2 U3210 ( .A0N(n9284), .A1N(n7963), .B0(n8089), .Y(n7979) );
  AOI2BB1X4 U3211 ( .A0N(n3808), .A1N(n7453), .B0(n3740), .Y(n7455) );
  CLKINVX1 U3212 ( .A(n7547), .Y(n7549) );
  CLKINVX8 U3213 ( .A(net99504), .Y(net106564) );
  MX2XL U3214 ( .A(n3496), .B(n178), .S0(n5511), .Y(\i_MIPS/n423 ) );
  MX2XL U3215 ( .A(\i_MIPS/EX_MEM[6] ), .B(net98929), .S0(n5508), .Y(
        \i_MIPS/n468 ) );
  OAI221X2 U3216 ( .A0(ICACHE_addr[0]), .A1(net98430), .B0(n11191), .B1(n3610), 
        .C0(n11190), .Y(\i_MIPS/PC/n36 ) );
  CLKMX2X3 U3217 ( .A(n8710), .B(n8709), .S0(net108959), .Y(net103059) );
  NAND3X8 U3218 ( .A(n4504), .B(n4505), .C(n4506), .Y(n4507) );
  CLKINVX8 U3219 ( .A(n10329), .Y(n4504) );
  OAI2BB1X4 U3220 ( .A0N(n3831), .A1N(n7029), .B0(n7028), .Y(n7033) );
  NAND2X6 U3221 ( .A(n3827), .B(n6939), .Y(n7028) );
  NAND2X6 U3222 ( .A(n10499), .B(n10378), .Y(n10497) );
  CLKBUFX2 U3223 ( .A(n5316), .Y(n5291) );
  CLKINVX3 U3224 ( .A(n5157), .Y(n5150) );
  INVX3 U3225 ( .A(n9552), .Y(n9570) );
  OA22X2 U3226 ( .A0(\i_MIPS/n365 ), .A1(n4811), .B0(\i_MIPS/n364 ), .B1(n4804), .Y(n7039) );
  INVX20 U3227 ( .A(n4814), .Y(n4811) );
  INVX20 U3228 ( .A(n4808), .Y(n4804) );
  OA22XL U3229 ( .A0(n5429), .A1(n1052), .B0(n5385), .B1(n2624), .Y(n9329) );
  AOI22XL U3230 ( .A0(n4800), .A1(n7862), .B0(n7861), .B1(n3636), .Y(n3612) );
  NAND2X1 U3231 ( .A(n4728), .B(\i_MIPS/PC/n4 ), .Y(n11042) );
  NAND2X4 U3232 ( .A(n4727), .B(net113039), .Y(n10581) );
  CLKINVX8 U3233 ( .A(n9566), .Y(n9555) );
  CLKINVX16 U3234 ( .A(net139669), .Y(net130576) );
  BUFX2 U3235 ( .A(n5188), .Y(n5157) );
  OR2X4 U3236 ( .A(net107042), .B(net112723), .Y(n3616) );
  INVX2 U3237 ( .A(net98994), .Y(net107042) );
  OAI222X4 U3238 ( .A0(n8154), .A1(n8805), .B0(n8659), .B1(n8151), .C0(n8887), 
        .C1(n9004), .Y(n8169) );
  CLKINVX3 U3239 ( .A(n5156), .Y(n5151) );
  BUFX4 U3240 ( .A(n5464), .Y(n5466) );
  AOI2BB1X2 U3241 ( .A0N(n7095), .A1N(n7094), .B0(n7093), .Y(n7097) );
  INVX3 U3242 ( .A(n7801), .Y(n7803) );
  BUFX20 U3243 ( .A(n4502), .Y(n4005) );
  AOI2BB2X4 U3244 ( .B0(n3617), .B1(\I_cache/cache[7][139] ), .A0N(n5420), 
        .A1N(n1897), .Y(n5952) );
  INVX2 U3245 ( .A(net99932), .Y(n4146) );
  INVX20 U3246 ( .A(net110205), .Y(net140281) );
  NAND3X4 U3247 ( .A(net98898), .B(net98900), .C(net98899), .Y(n4127) );
  CLKBUFX3 U3248 ( .A(n5143), .Y(n5115) );
  XNOR2X1 U3249 ( .A(n6292), .B(\i_MIPS/IR_ID[16] ), .Y(n4702) );
  INVX16 U3250 ( .A(net110255), .Y(net110251) );
  BUFX4 U3251 ( .A(n5464), .Y(n5465) );
  AO22X4 U3252 ( .A0(n7192), .A1(n9259), .B0(n9258), .B1(n7191), .Y(n7206) );
  CLKINVX3 U3253 ( .A(n5136), .Y(n5108) );
  OR2X4 U3254 ( .A(n11194), .B(net110249), .Y(n4185) );
  CLKINVX3 U3255 ( .A(n5217), .Y(n5196) );
  OR2XL U3256 ( .A(n7825), .B(net102087), .Y(net139681) );
  CLKMX2X4 U3257 ( .A(n7775), .B(n7774), .S0(n5588), .Y(n7825) );
  AND2X4 U3258 ( .A(n4687), .B(n4655), .Y(n4623) );
  AOI2BB2X2 U3259 ( .B0(\i_MIPS/IF_ID[94] ), .B1(n148), .A0N(net110189), .A1N(
        \i_MIPS/n209 ), .Y(n10505) );
  AOI2BB2X2 U3260 ( .B0(\i_MIPS/IF_ID[71] ), .B1(n147), .A0N(net110191), .A1N(
        \i_MIPS/n186 ), .Y(n11070) );
  AOI2BB2X2 U3261 ( .B0(\i_MIPS/IF_ID[69] ), .B1(n148), .A0N(net110191), .A1N(
        \i_MIPS/n184 ), .Y(n11197) );
  AO22X1 U3262 ( .A0(net110227), .A1(n10002), .B0(\i_MIPS/ID_EX_5 ), .B1(n5514), .Y(\i_MIPS/n478 ) );
  AOI22X1 U3263 ( .A0(\i_MIPS/ALUin1[20] ), .A1(n4815), .B0(
        \i_MIPS/ALUin1[19] ), .B1(n4809), .Y(n7023) );
  OA22XL U3264 ( .A0(\i_MIPS/ALUin1[26] ), .A1(n4811), .B0(\i_MIPS/ALUin1[27] ), .B1(n4804), .Y(n8640) );
  OA22XL U3265 ( .A0(\i_MIPS/ALUin1[25] ), .A1(n4811), .B0(\i_MIPS/ALUin1[26] ), .B1(n4804), .Y(n8347) );
  OA22XL U3266 ( .A0(\i_MIPS/ALUin1[7] ), .A1(n4811), .B0(\i_MIPS/ALUin1[6] ), 
        .B1(n4804), .Y(n7556) );
  OA22X1 U3267 ( .A0(\i_MIPS/n358 ), .A1(n4812), .B0(n6947), .B1(n4804), .Y(
        n6948) );
  OA22XL U3268 ( .A0(\i_MIPS/ALUin1[21] ), .A1(n4811), .B0(\i_MIPS/ALUin1[22] ), .B1(n4804), .Y(n7965) );
  OA22X1 U3269 ( .A0(\i_MIPS/ALUin1[22] ), .A1(n4811), .B0(\i_MIPS/ALUin1[23] ), .B1(n4804), .Y(n8271) );
  INVXL U3270 ( .A(n11364), .Y(n4343) );
  INVXL U3271 ( .A(n8098), .Y(n7696) );
  OR2X8 U3272 ( .A(n11097), .B(net110247), .Y(n4174) );
  NOR3X6 U3273 ( .A(n3784), .B(n3785), .C(n3786), .Y(n9009) );
  BUFX2 U3274 ( .A(n5229), .Y(n5202) );
  NAND2X8 U3275 ( .A(net101969), .B(n4145), .Y(net99932) );
  NAND4X6 U3276 ( .A(n4463), .B(n4464), .C(n5952), .D(n5953), .Y(n11375) );
  CLKINVX12 U3277 ( .A(net98429), .Y(net110205) );
  MX2XL U3278 ( .A(n10837), .B(net98915), .S0(n5508), .Y(\i_MIPS/n435 ) );
  CLKAND2X2 U3279 ( .A(n6944), .B(n7863), .Y(n3618) );
  AND2X8 U3280 ( .A(n6943), .B(n6942), .Y(n3619) );
  AND2X2 U3281 ( .A(n6941), .B(n6940), .Y(n3620) );
  OAI2BB1X2 U3282 ( .A0N(n4813), .A1N(\i_MIPS/ALU/N303 ), .B0(n9274), .Y(n7863) );
  NAND2XL U3283 ( .A(n7024), .B(n7025), .Y(n6943) );
  OAI222X1 U3284 ( .A0(n9004), .A1(n8911), .B0(n8728), .B1(n8913), .C0(n6779), 
        .C1(n8736), .Y(n6781) );
  NAND4X8 U3285 ( .A(n9606), .B(n9605), .C(n9604), .D(n9603), .Y(n9678) );
  INVX4 U3286 ( .A(n6234), .Y(n7619) );
  NAND2BX4 U3287 ( .AN(n5457), .B(n11243), .Y(n10053) );
  NAND2BX2 U3288 ( .AN(n5457), .B(n11244), .Y(n9999) );
  NAND4BX2 U3289 ( .AN(n8873), .B(n8872), .C(n8871), .D(n8870), .Y(n8884) );
  NAND4X2 U3290 ( .A(n3530), .B(n6217), .C(n4641), .D(n3769), .Y(n6219) );
  NAND2X6 U3291 ( .A(\i_MIPS/ALUin1[9] ), .B(n6230), .Y(n7096) );
  AOI211X2 U3292 ( .A0(n8822), .A1(n7290), .B0(n7289), .C0(n7288), .Y(n7291)
         );
  OAI222X2 U3293 ( .A0(n8814), .A1(n7628), .B0(n7561), .B1(n8085), .C0(n8726), 
        .C1(n8084), .Y(n7289) );
  AO22X2 U3294 ( .A0(n114), .A1(ICACHE_addr[19]), .B0(n5463), .B1(n11378), .Y(
        n11034) );
  NAND3BX4 U3295 ( .AN(n10735), .B(n10734), .C(n10733), .Y(n11544) );
  AND3X4 U3296 ( .A(n4143), .B(n4142), .C(net110227), .Y(n3622) );
  AND2X8 U3297 ( .A(n3622), .B(n4144), .Y(n4130) );
  OA21X4 U3298 ( .A0(n6938), .A1(n6937), .B0(n6935), .Y(n3623) );
  BUFX20 U3299 ( .A(net110233), .Y(net110227) );
  AOI2BB1X2 U3300 ( .A0N(net99849), .A1N(net99664), .B0(n4146), .Y(n4143) );
  OR2X2 U3301 ( .A(net106565), .B(net112707), .Y(n3691) );
  NAND3BX2 U3302 ( .AN(n6604), .B(n6603), .C(n6602), .Y(n3624) );
  NAND3X6 U3303 ( .A(n3320), .B(n7781), .C(n3625), .Y(n3626) );
  INVX2 U3304 ( .A(n8518), .Y(n3625) );
  AOI21X4 U3305 ( .A0(n9165), .A1(n2802), .B0(n9167), .Y(n6597) );
  INVX4 U3306 ( .A(n11044), .Y(n11003) );
  OA22X4 U3307 ( .A0(net112427), .A1(n1937), .B0(n3688), .B1(n357), .Y(n6091)
         );
  OA22X2 U3308 ( .A0(n8659), .A1(n7028), .B0(n9285), .B1(n7561), .Y(n6958) );
  OAI2BB2X4 U3309 ( .B0(n3628), .B1(n11065), .A0N(n9623), .A1N(n9622), .Y(
        n10209) );
  MX2X1 U3310 ( .A(\I_cache/cache[4][139] ), .B(n10976), .S0(n4676), .Y(n11707) );
  BUFX20 U3311 ( .A(net111409), .Y(net111405) );
  CLKINVX1 U3312 ( .A(n3666), .Y(n8666) );
  OR2X4 U3313 ( .A(n10914), .B(n10913), .Y(n4408) );
  OAI222X4 U3314 ( .A0(n7974), .A1(n7544), .B0(n8659), .B1(n7550), .C0(n8817), 
        .C1(n7543), .Y(n7568) );
  CLKAND2X12 U3315 ( .A(n6364), .B(n6363), .Y(n3845) );
  OA21X4 U3316 ( .A0(n8893), .A1(n4523), .B0(n8890), .Y(n6645) );
  AO21X4 U3317 ( .A0(n4823), .A1(\i_MIPS/ALU/N303 ), .B0(n6356), .Y(n7279) );
  NAND2X4 U3318 ( .A(n8818), .B(n7785), .Y(n6368) );
  INVX6 U3319 ( .A(n7559), .Y(n7974) );
  NAND2X6 U3320 ( .A(n6232), .B(\i_MIPS/n368 ), .Y(n8711) );
  CLKINVX3 U3321 ( .A(n10369), .Y(n10368) );
  OR2XL U3322 ( .A(n4503), .B(net110215), .Y(n4183) );
  NAND3X4 U3323 ( .A(n4503), .B(n3676), .C(n4424), .Y(n4451) );
  AND2X8 U3324 ( .A(net134093), .B(net99671), .Y(n4527) );
  BUFX2 U3325 ( .A(n5451), .Y(n5421) );
  INVX6 U3326 ( .A(n9255), .Y(n10582) );
  OAI221X4 U3327 ( .A0(n9254), .A1(net102087), .B0(net113075), .B1(n10696), 
        .C0(n9253), .Y(n9255) );
  OA22X4 U3328 ( .A0(net112499), .A1(n1938), .B0(n3688), .B1(n358), .Y(n6077)
         );
  CLKINVX1 U3329 ( .A(n6240), .Y(n3632) );
  NAND2X6 U3330 ( .A(n6239), .B(\i_MIPS/n364 ), .Y(n7462) );
  AOI31X4 U3331 ( .A0(n6479), .A1(n6846), .A2(n3747), .B0(n6478), .Y(n6480) );
  OAI2BB1X2 U3332 ( .A0N(n6463), .A1N(n7031), .B0(n7030), .Y(n6474) );
  CLKINVX3 U3333 ( .A(n5221), .Y(n5197) );
  OAI2BB1X2 U3334 ( .A0N(n7357), .A1N(n7457), .B0(n7359), .Y(n7274) );
  CLKINVX1 U3335 ( .A(n6599), .Y(n6225) );
  CLKINVX8 U3336 ( .A(net103630), .Y(net99711) );
  NAND2X6 U3337 ( .A(n9133), .B(n7698), .Y(n9007) );
  CLKBUFX2 U3338 ( .A(n7477), .Y(n3634) );
  OAI221X2 U3339 ( .A0(net102744), .A1(net112707), .B0(net102745), .B1(
        net112721), .C0(net102746), .Y(net99080) );
  OAI221X1 U3340 ( .A0(n4798), .A1(n7465), .B0(n7464), .B1(n9262), .C0(n8805), 
        .Y(n7467) );
  CLKINVX1 U3341 ( .A(n10488), .Y(n10491) );
  XOR3X2 U3342 ( .A(n11065), .B(n11064), .C(n11063), .Y(n11067) );
  AOI2BB1X2 U3343 ( .A0N(n11062), .A1N(n11061), .B0(n11060), .Y(n11064) );
  AOI21X1 U3344 ( .A0(n8804), .A1(n8803), .B0(n8715), .Y(n4552) );
  AOI2BB1X4 U3345 ( .A0N(n8893), .A1N(n8249), .B0(n6637), .Y(n6644) );
  NAND2X2 U3346 ( .A(n4659), .B(n4657), .Y(n6508) );
  NAND2X2 U3347 ( .A(n4659), .B(n4656), .Y(n6511) );
  NOR2X2 U3348 ( .A(n3697), .B(n8527), .Y(n3696) );
  CLKBUFX4 U3349 ( .A(n4480), .Y(n4930) );
  OA22X1 U3350 ( .A0(\i_MIPS/Register/register[6][17] ), .A1(n4937), .B0(
        \i_MIPS/Register/register[14][17] ), .B1(n4930), .Y(n7673) );
  AOI22X4 U3351 ( .A0(net113039), .A1(net99605), .B0(net102300), .B1(net103479), .Y(net134117) );
  AOI22X4 U3352 ( .A0(net113039), .A1(net99290), .B0(net102300), .B1(net104440), .Y(net134118) );
  CLKBUFX4 U3353 ( .A(net102036), .Y(net113039) );
  NAND2X8 U3354 ( .A(n8260), .B(\i_MIPS/ID_EX[83] ), .Y(n8728) );
  CLKMX2X2 U3355 ( .A(n8354), .B(n7967), .S0(n5590), .Y(n9269) );
  OAI221X4 U3356 ( .A0(\i_MIPS/ALUin1[19] ), .A1(n4824), .B0(
        \i_MIPS/ALUin1[20] ), .B1(n4817), .C0(n7965), .Y(n8354) );
  CLKBUFX3 U3357 ( .A(n5142), .Y(n5125) );
  MX2XL U3358 ( .A(n4498), .B(n3523), .S0(n5507), .Y(\i_MIPS/n393 ) );
  INVX12 U3359 ( .A(n9280), .Y(n9141) );
  CLKINVX1 U3360 ( .A(n11087), .Y(n11086) );
  NAND2X8 U3361 ( .A(n11196), .B(n3516), .Y(n11048) );
  CLKINVX8 U3362 ( .A(n9678), .Y(n11196) );
  OAI211X2 U3363 ( .A0(n9137), .A1(n8354), .B0(n8353), .C0(n4501), .Y(n8355)
         );
  MX2X1 U3364 ( .A(n7966), .B(n7872), .S0(n5590), .Y(n8343) );
  NAND3BX2 U3365 ( .AN(n4690), .B(n7871), .C(n7870), .Y(n7966) );
  OR2X2 U3366 ( .A(n9212), .B(net112707), .Y(n4166) );
  INVX20 U3367 ( .A(n4827), .Y(n4824) );
  CLKINVX1 U3368 ( .A(n4328), .Y(n3639) );
  NAND4X6 U3369 ( .A(n4455), .B(n4456), .C(n5980), .D(n5979), .Y(n11371) );
  INVX3 U3370 ( .A(n9152), .Y(n9157) );
  OA22X4 U3371 ( .A0(n9284), .A1(n8085), .B0(n9007), .B1(n8084), .Y(n8093) );
  INVX6 U3372 ( .A(n4425), .Y(n3693) );
  NAND2X1 U3373 ( .A(n8921), .B(n8920), .Y(n8926) );
  NAND2X2 U3374 ( .A(\i_MIPS/ALUin1[30] ), .B(n11223), .Y(n9256) );
  NAND4BX4 U3375 ( .AN(n6422), .B(n3706), .C(n6444), .D(n4585), .Y(n6440) );
  NAND3BX1 U3376 ( .AN(n9151), .B(n4591), .C(n9160), .Y(n6443) );
  NAND2X4 U3377 ( .A(n6234), .B(\i_MIPS/n370 ), .Y(n7626) );
  MX2X1 U3378 ( .A(n9280), .B(n9279), .S0(n3773), .Y(n7202) );
  NOR2X2 U3379 ( .A(n4556), .B(net110241), .Y(n4430) );
  OR2X2 U3380 ( .A(n4562), .B(net110241), .Y(n4184) );
  OR2X2 U3381 ( .A(n4538), .B(net110241), .Y(n4190) );
  AOI2BB2XL U3382 ( .B0(\i_MIPS/BranchAddr[0] ), .B1(net113592), .A0N(n4546), 
        .A1N(net110241), .Y(n10816) );
  NAND2X4 U3383 ( .A(n7953), .B(n8514), .Y(n4154) );
  OAI2BB1X1 U3384 ( .A0N(n9277), .A1N(n9179), .B0(n9260), .Y(n3657) );
  NAND2X1 U3385 ( .A(n10699), .B(n168), .Y(n10701) );
  NAND2X1 U3386 ( .A(n10500), .B(n168), .Y(n10704) );
  INVX2 U3387 ( .A(n10327), .Y(n4506) );
  NAND2X1 U3388 ( .A(n10965), .B(net113551), .Y(n10324) );
  NAND3BX4 U3389 ( .AN(n10723), .B(n10721), .C(n10724), .Y(n10729) );
  AOI2BB1X2 U3390 ( .A0N(n3609), .A1N(n10949), .B0(n10948), .Y(n10951) );
  AOI2BB1XL U3391 ( .A0N(n10211), .A1N(n10210), .B0(n10209), .Y(n9624) );
  XOR2X4 U3392 ( .A(n3644), .B(n3658), .Y(n4097) );
  NAND2X6 U3393 ( .A(n3312), .B(net99634), .Y(n3644) );
  CLKINVX1 U3394 ( .A(n3645), .Y(n3646) );
  CLKINVX1 U3395 ( .A(n3647), .Y(n3648) );
  CLKINVX1 U3396 ( .A(n3649), .Y(n3650) );
  OR2X2 U3397 ( .A(n4534), .B(net110241), .Y(n4421) );
  AO22XL U3398 ( .A0(ICACHE_addr[16]), .A1(mem_read_I), .B0(n4796), .B1(n3564), 
        .Y(n12834) );
  AO22X2 U3399 ( .A0(n4551), .A1(n9259), .B0(n9258), .B1(n7274), .Y(n7276) );
  INVXL U3400 ( .A(net106564), .Y(n3651) );
  OR2X1 U3401 ( .A(\i_MIPS/PC/n21 ), .B(net110213), .Y(n3652) );
  NAND3X2 U3402 ( .A(n3653), .B(n3652), .C(n3654), .Y(n11155) );
  INVXL U3403 ( .A(net99991), .Y(net98501) );
  OAI221X4 U3404 ( .A0(\i_MIPS/n367 ), .A1(n4824), .B0(\i_MIPS/n366 ), .B1(
        n4816), .C0(n7039), .Y(n7474) );
  NOR3BX4 U3405 ( .AN(n4617), .B(n6226), .C(n6225), .Y(n6227) );
  NAND3BX1 U3406 ( .AN(n4588), .B(n11200), .C(n9810), .Y(\i_MIPS/n470 ) );
  AO21X4 U3407 ( .A0(n6651), .A1(n8333), .B0(n6650), .Y(n8661) );
  OR2X4 U3408 ( .A(n7095), .B(n6927), .Y(n4209) );
  AND2X8 U3409 ( .A(n6645), .B(n8894), .Y(n3850) );
  NOR4X2 U3410 ( .A(n8953), .B(n8952), .C(n8951), .D(n8950), .Y(n8954) );
  NAND4X2 U3411 ( .A(n8948), .B(n8947), .C(n8946), .D(n8945), .Y(n8953) );
  OA22XL U3412 ( .A0(\i_MIPS/Register/register[3][28] ), .A1(n4868), .B0(
        \i_MIPS/Register/register[11][28] ), .B1(n4858), .Y(n9025) );
  OA22X2 U3413 ( .A0(\i_MIPS/Register/register[19][28] ), .A1(n4868), .B0(
        \i_MIPS/Register/register[27][28] ), .B1(n4858), .Y(n9034) );
  OA22XL U3414 ( .A0(\i_MIPS/Register/register[19][24] ), .A1(n4868), .B0(
        \i_MIPS/Register/register[27][24] ), .B1(n4858), .Y(n8946) );
  NAND2X4 U3415 ( .A(n6246), .B(\i_MIPS/ALUin1[11] ), .Y(n7099) );
  OR2X4 U3416 ( .A(n10866), .B(net110249), .Y(n3656) );
  BUFX4 U3417 ( .A(net110229), .Y(net110215) );
  AOI33X2 U3418 ( .A0(n9258), .A1(n7714), .A2(n7713), .B0(n9258), .B1(n7712), 
        .B2(n7711), .Y(n7715) );
  CLKXOR2X2 U3419 ( .A(n9430), .B(n3649), .Y(n10900) );
  AO22X2 U3420 ( .A0(n115), .A1(n3649), .B0(n5463), .B1(n11367), .Y(n10994) );
  XOR2X1 U3421 ( .A(n10289), .B(ICACHE_addr[17]), .Y(n11151) );
  AND2XL U3422 ( .A(net134118), .B(net99270), .Y(n4559) );
  INVX1 U3423 ( .A(n6443), .Y(n6446) );
  INVX1 U3424 ( .A(n11223), .Y(n9268) );
  OA22X1 U3425 ( .A0(\i_MIPS/Register/register[5][7] ), .A1(n4849), .B0(
        \i_MIPS/Register/register[13][7] ), .B1(n4841), .Y(n7504) );
  INVX8 U3426 ( .A(n4853), .Y(n4849) );
  NAND2X2 U3427 ( .A(n10885), .B(n10884), .Y(n10893) );
  NAND4X6 U3428 ( .A(n6685), .B(n6684), .C(n6683), .D(n6682), .Y(net99504) );
  CLKMX2X2 U3429 ( .A(n9141), .B(n4799), .S0(n7287), .Y(n7288) );
  AND2X8 U3430 ( .A(n3593), .B(net100866), .Y(n3695) );
  AOI222X4 U3431 ( .A0(n7624), .A1(n7623), .B0(n4598), .B1(n8822), .C0(n8820), 
        .C1(n7693), .Y(n7630) );
  NAND2X4 U3432 ( .A(n4587), .B(\i_MIPS/ID_EX[83] ), .Y(n9284) );
  CLKXOR2X1 U3433 ( .A(net111405), .B(n10959), .Y(n3660) );
  XOR2X4 U3434 ( .A(n10955), .B(n3660), .Y(n10957) );
  NAND2X2 U3435 ( .A(n11044), .B(n11043), .Y(n3661) );
  CLKINVX1 U3436 ( .A(n11002), .Y(n11043) );
  OA22XL U3437 ( .A0(\i_MIPS/Register/register[3][24] ), .A1(n4868), .B0(
        \i_MIPS/Register/register[11][24] ), .B1(n4858), .Y(n8937) );
  NOR4X2 U3438 ( .A(n8944), .B(n8943), .C(n8942), .D(n8941), .Y(n8955) );
  CLKBUFX2 U3439 ( .A(n4622), .Y(n4836) );
  BUFX8 U3440 ( .A(net101981), .Y(net112725) );
  XNOR2X4 U3441 ( .A(n3663), .B(n152), .Y(n4080) );
  NAND2X1 U3442 ( .A(n4828), .B(n6947), .Y(n7104) );
  OAI211X4 U3443 ( .A0(\i_MIPS/ALUin1[15] ), .A1(n4818), .B0(n7104), .C0(n6671), .Y(n7697) );
  INVX20 U3444 ( .A(n4821), .Y(n4818) );
  OAI2BB1X4 U3445 ( .A0N(net98970), .A1N(net98971), .B0(net113041), .Y(
        net98966) );
  BUFX8 U3446 ( .A(n5362), .Y(n5329) );
  OA22X2 U3447 ( .A0(n10901), .A1(net140280), .B0(net98430), .B1(n10900), .Y(
        n10903) );
  OA22X2 U3448 ( .A0(n3289), .A1(n3600), .B0(n9262), .B1(n7098), .Y(n7119) );
  CLKINVX8 U3449 ( .A(n7968), .Y(n8260) );
  OAI32X4 U3450 ( .A0(n6934), .A1(n6931), .A2(n6930), .B0(n1224), .B1(n6931), 
        .Y(n6937) );
  NAND3BX4 U3451 ( .AN(n8360), .B(n8359), .C(n4928), .Y(n8361) );
  INVXL U3452 ( .A(n3316), .Y(n3705) );
  AOI2BB2X2 U3453 ( .B0(n9258), .B1(n9179), .A0N(n9262), .A1N(n3574), .Y(n9293) );
  CLKAND2X12 U3454 ( .A(n7545), .B(n7454), .Y(n3665) );
  NAND3X6 U3455 ( .A(n8164), .B(n8166), .C(n3290), .Y(n8168) );
  CLKINVX3 U3456 ( .A(n3638), .Y(n7615) );
  OAI222X2 U3457 ( .A0(n8726), .A1(n3), .B0(n3638), .B1(n7367), .C0(n8729), 
        .C1(n7366), .Y(n7369) );
  NAND4X2 U3458 ( .A(n8376), .B(n8375), .C(n8374), .D(n8373), .Y(n8381) );
  INVX2 U3459 ( .A(n10944), .Y(n10940) );
  NAND2X4 U3460 ( .A(n10940), .B(net113551), .Y(n11013) );
  AND2X8 U3461 ( .A(n11015), .B(n11013), .Y(n4508) );
  INVXL U3462 ( .A(n3547), .Y(n3667) );
  INVXL U3463 ( .A(n7545), .Y(n3669) );
  CLKINVX1 U3464 ( .A(n3669), .Y(n3670) );
  INVX12 U3465 ( .A(n6612), .Y(n6939) );
  NAND2X6 U3466 ( .A(n6612), .B(n6947), .Y(n7029) );
  CLKINVX3 U3467 ( .A(n5112), .Y(n5111) );
  MX2XL U3468 ( .A(\i_MIPS/ID_EX[49] ), .B(net98946), .S0(n5510), .Y(
        \i_MIPS/n421 ) );
  CLKAND2X3 U3469 ( .A(n4802), .B(n7698), .Y(n4577) );
  NAND2X8 U3470 ( .A(n4200), .B(n4201), .Y(n6566) );
  NAND2X4 U3471 ( .A(n4644), .B(n3771), .Y(n4201) );
  NAND2X6 U3472 ( .A(\i_MIPS/ALUin1[17] ), .B(n6566), .Y(n7856) );
  OAI221X2 U3473 ( .A0(net106418), .A1(net112709), .B0(net106419), .B1(
        net112723), .C0(net106420), .Y(net98946) );
  MXI2X4 U3474 ( .A(n3820), .B(n3525), .S0(n3826), .Y(n3823) );
  AOI2BB2X4 U3475 ( .B0(net111873), .B1(\D_cache/cache[7][129] ), .A0N(
        net112037), .A1N(n1898), .Y(n6121) );
  NAND2X6 U3476 ( .A(n3677), .B(n10675), .Y(n6115) );
  INVX6 U3477 ( .A(n6114), .Y(n10675) );
  BUFX12 U3478 ( .A(net111967), .Y(net111931) );
  INVXL U3479 ( .A(n7619), .Y(n3674) );
  CLKINVX1 U3480 ( .A(n3674), .Y(n3675) );
  OR2X4 U3481 ( .A(net112147), .B(n1988), .Y(n4222) );
  OA22X4 U3482 ( .A0(net112037), .A1(n2356), .B0(net111965), .B1(n360), .Y(
        n6125) );
  NAND2X6 U3483 ( .A(n4604), .B(n10157), .Y(n10145) );
  CLKMX2X2 U3484 ( .A(\D_cache/cache[2][26] ), .B(n4257), .S0(net112401), .Y(
        \D_cache/n1586 ) );
  NAND2X8 U3485 ( .A(n3682), .B(n3683), .Y(n6157) );
  AOI2BB2X2 U3486 ( .B0(n3813), .B1(\D_cache/cache[2][133] ), .A0N(net112379), 
        .A1N(n2005), .Y(n6145) );
  INVX2 U3487 ( .A(net112427), .Y(n3813) );
  BUFX12 U3488 ( .A(net112585), .Y(net112571) );
  AOI211X4 U3489 ( .A0(n6476), .A1(n6638), .B0(n6475), .C0(n6474), .Y(n6481)
         );
  AOI222X1 U3490 ( .A0(n5474), .A1(n11484), .B0(mem_rdata_D[97]), .B1(n116), 
        .C0(n12996), .C1(n5473), .Y(n10839) );
  AO22X4 U3491 ( .A0(net113445), .A1(n11453), .B0(net102346), .B1(n11484), .Y(
        n7649) );
  NAND2X1 U3492 ( .A(n8712), .B(n3836), .Y(n7356) );
  NOR3X4 U3493 ( .A(n3678), .B(n3679), .C(n3680), .Y(n3677) );
  NOR2X2 U3494 ( .A(net112583), .B(n1892), .Y(n3679) );
  OAI22X2 U3495 ( .A0(net112449), .A1(n314), .B0(net112325), .B1(n1889), .Y(
        n3680) );
  OAI221X2 U3496 ( .A0(net103218), .A1(net112707), .B0(n3834), .B1(net112721), 
        .C0(net103220), .Y(net99432) );
  OAI222X2 U3497 ( .A0(n9005), .A1(n141), .B0(n9007), .B1(n8535), .C0(n9010), 
        .C1(n8534), .Y(n8551) );
  NAND3BX2 U3498 ( .AN(n7968), .B(n4577), .C(n3787), .Y(n8534) );
  NAND2BX1 U3499 ( .AN(net112137), .B(\D_cache/cache[5][148] ), .Y(n4187) );
  CLKMX2X4 U3500 ( .A(n7474), .B(n7473), .S0(n5590), .Y(n7475) );
  AND2XL U3501 ( .A(n4605), .B(n10731), .Y(n4525) );
  NAND2X6 U3502 ( .A(n10627), .B(n3687), .Y(n3748) );
  NOR2X6 U3503 ( .A(n6058), .B(n1877), .Y(n3687) );
  OR2X8 U3504 ( .A(n8424), .B(net112721), .Y(n3729) );
  AOI2BB1X2 U3505 ( .A0N(\i_MIPS/n368 ), .A1N(n3592), .B0(n4674), .Y(n7038) );
  CLKBUFX8 U3506 ( .A(net112381), .Y(net112333) );
  BUFX16 U3507 ( .A(net112383), .Y(net112325) );
  NAND2X4 U3508 ( .A(n4686), .B(n4656), .Y(n6515) );
  NAND2X4 U3509 ( .A(n4686), .B(n4657), .Y(n6512) );
  AO22X1 U3510 ( .A0(n4979), .A1(n552), .B0(n9309), .B1(n2055), .Y(n8497) );
  BUFX3 U3511 ( .A(n9310), .Y(n4979) );
  NAND3X8 U3512 ( .A(n8713), .B(n3197), .C(n8714), .Y(n6767) );
  OR3X8 U3513 ( .A(n4409), .B(n4410), .C(n9262), .Y(n9020) );
  NAND2X1 U3514 ( .A(n4814), .B(\i_MIPS/ALUin1[1] ), .Y(n6946) );
  CLKINVX1 U3515 ( .A(n8819), .Y(n8349) );
  CLKMX2X2 U3516 ( .A(n7557), .B(n8819), .S0(n5589), .Y(n7558) );
  CLKMX2X2 U3517 ( .A(n6705), .B(n6704), .S0(net108963), .Y(net106565) );
  AO21X2 U3518 ( .A0(net99502), .A1(net99503), .B0(net112727), .Y(net106566)
         );
  MX2X2 U3519 ( .A(n9043), .B(n9042), .S0(n5587), .Y(net102500) );
  OA22X1 U3520 ( .A0(\i_MIPS/Register/register[17][24] ), .A1(n4835), .B0(
        \i_MIPS/Register/register[25][24] ), .B1(n4830), .Y(n8948) );
  OA22X1 U3521 ( .A0(\i_MIPS/Register/register[1][24] ), .A1(n4835), .B0(
        \i_MIPS/Register/register[9][24] ), .B1(n4829), .Y(n8939) );
  OA22X2 U3522 ( .A0(\i_MIPS/Register/register[17][28] ), .A1(n4835), .B0(
        \i_MIPS/Register/register[25][28] ), .B1(n4830), .Y(n9036) );
  OA22X4 U3523 ( .A0(n5250), .A1(n1939), .B0(n5227), .B1(n361), .Y(n6026) );
  OA22X4 U3524 ( .A0(n5429), .A1(n1940), .B0(n5385), .B1(n362), .Y(n6024) );
  AOI2BB1X4 U3525 ( .A0N(n8326), .A1N(n8914), .B0(n6593), .Y(n6595) );
  INVX4 U3526 ( .A(n8435), .Y(n8326) );
  INVXL U3527 ( .A(net104184), .Y(n3694) );
  XOR2X4 U3528 ( .A(n3695), .B(n181), .Y(n4092) );
  NAND2X6 U3529 ( .A(n7850), .B(n4520), .Y(n8163) );
  MX2X1 U3530 ( .A(\I_cache/cache[2][142] ), .B(n11034), .S0(n5234), .Y(n11685) );
  OA22X4 U3531 ( .A0(\i_MIPS/n344 ), .A1(n4811), .B0(\i_MIPS/n345 ), .B1(n4805), .Y(n6951) );
  NOR2X4 U3532 ( .A(net111967), .B(n1878), .Y(n4207) );
  CLKBUFX8 U3533 ( .A(n4905), .Y(n4908) );
  OA22XL U3534 ( .A0(\i_MIPS/Register/register[22][28] ), .A1(n4914), .B0(
        \i_MIPS/Register/register[30][28] ), .B1(n4908), .Y(n9037) );
  OA22X1 U3535 ( .A0(\i_MIPS/Register/register[22][24] ), .A1(n4914), .B0(
        \i_MIPS/Register/register[30][24] ), .B1(n4908), .Y(n8949) );
  OA22XL U3536 ( .A0(\i_MIPS/Register/register[6][24] ), .A1(n4914), .B0(
        \i_MIPS/Register/register[14][24] ), .B1(n4908), .Y(n8940) );
  AND2X4 U3537 ( .A(n4827), .B(\i_MIPS/ALUin1[26] ), .Y(n4671) );
  XOR2X4 U3538 ( .A(n6054), .B(n12939), .Y(n6072) );
  OA22X4 U3539 ( .A0(n5333), .A1(n3275), .B0(n5290), .B1(n1619), .Y(n6021) );
  CLKMX2X2 U3540 ( .A(n9141), .B(n4799), .S0(n8734), .Y(n8735) );
  CLKINVX6 U3541 ( .A(n6605), .Y(n6606) );
  INVX6 U3542 ( .A(n6078), .Y(n10648) );
  AO22X1 U3543 ( .A0(n114), .A1(ICACHE_addr[21]), .B0(n5463), .B1(n11380), .Y(
        n10975) );
  OR2X2 U3544 ( .A(net112147), .B(n2800), .Y(n4224) );
  CLKINVX20 U3545 ( .A(n3770), .Y(n3771) );
  NAND2X8 U3546 ( .A(n10651), .B(n10650), .Y(n6086) );
  NAND4X2 U3547 ( .A(n8258), .B(n8921), .C(n8255), .D(n9258), .Y(n8286) );
  MX2XL U3548 ( .A(n10508), .B(net99464), .S0(n5509), .Y(\i_MIPS/n379 ) );
  NAND2X4 U3549 ( .A(\i_MIPS/ALUin1[17] ), .B(n6574), .Y(n7847) );
  AO22XL U3550 ( .A0(ICACHE_addr[21]), .A1(mem_read_I), .B0(n4796), .B1(n11380), .Y(n12829) );
  MX2X1 U3551 ( .A(\i_MIPS/n249 ), .B(n4639), .S0(n3826), .Y(n11223) );
  NAND2X6 U3552 ( .A(n7626), .B(n6427), .Y(n6450) );
  XOR2X4 U3553 ( .A(net99991), .B(n3316), .Y(n4105) );
  OR2X4 U3554 ( .A(net112561), .B(n2415), .Y(n4165) );
  MXI2X4 U3555 ( .A(n10766), .B(n10765), .S0(n5490), .Y(n10767) );
  NAND2X6 U3556 ( .A(n10679), .B(n10678), .Y(n6123) );
  OR2XL U3557 ( .A(n9211), .B(net112721), .Y(n3702) );
  AOI222X2 U3558 ( .A0(n5488), .A1(n11432), .B0(mem_rdata_D[44]), .B1(n117), 
        .C0(n12985), .C1(n5484), .Y(n10799) );
  BUFX20 U3559 ( .A(n4575), .Y(n5484) );
  CLKINVX8 U3560 ( .A(net106078), .Y(net99814) );
  AND3X8 U3561 ( .A(n8558), .B(n8560), .C(n3319), .Y(n3834) );
  NAND2X6 U3562 ( .A(n4140), .B(n4141), .Y(n4125) );
  NAND3BX4 U3563 ( .AN(n10394), .B(n10392), .C(n10393), .Y(\i_MIPS/PC/n62 ) );
  NAND2X2 U3564 ( .A(net111409), .B(n10342), .Y(n10362) );
  OA22X2 U3565 ( .A0(n10889), .A1(net140280), .B0(net98430), .B1(n10888), .Y(
        n10891) );
  NAND2X6 U3566 ( .A(net99935), .B(net99936), .Y(n4120) );
  OAI221X2 U3567 ( .A0(n4798), .A1(n6347), .B0(n6248), .B1(n9262), .C0(n8805), 
        .Y(n6253) );
  CLKAND2X8 U3568 ( .A(n5956), .B(n9557), .Y(n4614) );
  INVXL U3569 ( .A(net104024), .Y(n3703) );
  NAND2BX2 U3570 ( .AN(n8526), .B(n8520), .Y(n8075) );
  AND2X6 U3571 ( .A(\i_MIPS/IR_ID[21] ), .B(\i_MIPS/n229 ), .Y(n4687) );
  NAND2X8 U3572 ( .A(n11003), .B(n11002), .Y(n11045) );
  AOI2BB1XL U3573 ( .A0N(\i_MIPS/ALUin1[15] ), .A1N(n4826), .B0(n4615), .Y(
        n6261) );
  INVXL U3574 ( .A(n4471), .Y(n3706) );
  OR2XL U3575 ( .A(n7270), .B(n8729), .Y(n3842) );
  INVXL U3576 ( .A(n3704), .Y(n3707) );
  CLKBUFX2 U3577 ( .A(n7454), .Y(n3796) );
  OAI2BB2X4 U3578 ( .B0(net102087), .B1(n3835), .A0N(net113041), .A1N(net99384), .Y(net103795) );
  MXI2X1 U3579 ( .A(n8248), .B(n8247), .S0(n5587), .Y(n3835) );
  NAND3BX4 U3580 ( .AN(n10922), .B(n10921), .C(n11094), .Y(n10923) );
  XNOR2X4 U3581 ( .A(n3710), .B(n3856), .Y(n4106) );
  NAND2X8 U3582 ( .A(n6232), .B(\i_MIPS/ALUin1[3] ), .Y(n8718) );
  OA22X1 U3583 ( .A0(net112041), .A1(n1234), .B0(net111917), .B1(n2839), .Y(
        n6273) );
  OA21X4 U3584 ( .A0(n7210), .A1(n7209), .B0(n7208), .Y(n3711) );
  AND2XL U3585 ( .A(n7187), .B(n7186), .Y(n7209) );
  OA22XL U3586 ( .A0(\i_MIPS/Register/register[6][3] ), .A1(n4914), .B0(
        \i_MIPS/Register/register[14][3] ), .B1(n4908), .Y(n8746) );
  OR2X2 U3587 ( .A(net103390), .B(net112707), .Y(n3712) );
  OA21X4 U3588 ( .A0(n8493), .A1(n8492), .B0(net113439), .Y(n3714) );
  NAND2X2 U3589 ( .A(n3714), .B(n3709), .Y(net99604) );
  AO22X4 U3590 ( .A0(net113445), .A1(n11476), .B0(net102346), .B1(n11507), .Y(
        n8492) );
  AO21X4 U3591 ( .A0(net99603), .A1(net99604), .B0(net113075), .Y(net99734) );
  OAI2BB1X4 U3592 ( .A0N(n10750), .A1N(n10751), .B0(net114085), .Y(net102746)
         );
  NAND2X2 U3593 ( .A(\i_MIPS/ALUin1[15] ), .B(n6613), .Y(n7031) );
  XOR2X4 U3594 ( .A(n3718), .B(DCACHE_addr[27]), .Y(n6167) );
  MXI2X4 U3595 ( .A(\i_MIPS/n301 ), .B(n6216), .S0(n3826), .Y(n3719) );
  OAI222X1 U3596 ( .A0(n8733), .A1(n8814), .B0(n7561), .B1(n8275), .C0(n8726), 
        .C1(n8274), .Y(n7479) );
  OA22X2 U3597 ( .A0(net111409), .A1(net140281), .B0(net98430), .B1(n11113), 
        .Y(n11115) );
  OA22X2 U3598 ( .A0(net112665), .A1(n927), .B0(net112563), .B1(n2451), .Y(
        n7927) );
  OA22X2 U3599 ( .A0(net112665), .A1(n928), .B0(net112563), .B1(n2452), .Y(
        n8024) );
  NAND2X2 U3600 ( .A(n8714), .B(n3608), .Y(n8806) );
  MX2XL U3601 ( .A(n12949), .B(n3703), .S0(n5507), .Y(\i_MIPS/n448 ) );
  INVXL U3602 ( .A(n3801), .Y(n6456) );
  OAI221X2 U3603 ( .A0(net112663), .A1(n2040), .B0(net112561), .B1(n702), .C0(
        n6164), .Y(n6165) );
  OA22X2 U3604 ( .A0(net112453), .A1(n1629), .B0(net112329), .B1(n3292), .Y(
        n6164) );
  NOR4X4 U3605 ( .A(n8550), .B(n8551), .C(n8552), .D(n8549), .Y(n8558) );
  NAND2XL U3606 ( .A(n10661), .B(n10660), .Y(n11539) );
  INVX6 U3607 ( .A(n6161), .Y(n10661) );
  CLKMX2X6 U3608 ( .A(n8533), .B(n8540), .S0(n5589), .Y(n8909) );
  NOR4X8 U3609 ( .A(n5984), .B(n9561), .C(n9560), .D(n9559), .Y(n9562) );
  INVX6 U3610 ( .A(n6133), .Y(n10673) );
  OAI221X4 U3611 ( .A0(net112229), .A1(n1225), .B0(net112147), .B1(n2804), 
        .C0(n6132), .Y(n6133) );
  NAND2X4 U3612 ( .A(n10632), .B(n3828), .Y(n6050) );
  INVX6 U3613 ( .A(n6049), .Y(n10632) );
  MX2X1 U3614 ( .A(n7106), .B(n7784), .S0(n5590), .Y(n7471) );
  OAI221X2 U3615 ( .A0(\i_MIPS/Register/register[2][0] ), .A1(n4944), .B0(
        \i_MIPS/Register/register[10][0] ), .B1(n4942), .C0(n6503), .Y(n6506)
         );
  AOI222X1 U3616 ( .A0(n5488), .A1(n11433), .B0(mem_rdata_D[45]), .B1(n116), 
        .C0(n12984), .C1(n5484), .Y(n10811) );
  NAND4X2 U3617 ( .A(n6380), .B(n6379), .C(n6378), .D(n6377), .Y(n11433) );
  CLKAND2X3 U3618 ( .A(n11360), .B(n135), .Y(n6172) );
  NAND2X2 U3619 ( .A(n5594), .B(\i_MIPS/ID_EX[81] ), .Y(n4436) );
  CLKBUFX8 U3620 ( .A(net112599), .Y(net112585) );
  NOR4X2 U3621 ( .A(n6986), .B(n6985), .C(n6984), .D(n6983), .Y(n6997) );
  INVX6 U3622 ( .A(n6080), .Y(n10647) );
  OAI221X2 U3623 ( .A0(net112655), .A1(n2041), .B0(net112587), .B1(n279), .C0(
        n6077), .Y(n6078) );
  NAND2X2 U3624 ( .A(n5593), .B(n4643), .Y(n4218) );
  OA22XL U3625 ( .A0(\i_MIPS/n355 ), .A1(n4826), .B0(\i_MIPS/n356 ), .B1(n4818), .Y(n6352) );
  NAND2BX2 U3626 ( .AN(net112583), .B(\D_cache/cache[1][141] ), .Y(n4149) );
  OA22X2 U3627 ( .A0(net112431), .A1(n450), .B0(net112379), .B1(n2006), .Y(
        n6135) );
  CLKINVX3 U3628 ( .A(n5443), .Y(n5415) );
  CLKBUFX3 U3629 ( .A(n5449), .Y(n5425) );
  CLKBUFX4 U3630 ( .A(n5404), .Y(n5381) );
  AND4X4 U3631 ( .A(n6444), .B(n6447), .C(n3686), .D(n4067), .Y(n3723) );
  INVX16 U3632 ( .A(n4495), .Y(n6660) );
  AND2XL U3633 ( .A(n3313), .B(net99974), .Y(n4536) );
  OR2X4 U3634 ( .A(n9174), .B(n9173), .Y(n4439) );
  CLKBUFX3 U3635 ( .A(n5404), .Y(n5380) );
  OAI221X2 U3636 ( .A0(net112265), .A1(n1616), .B0(net112143), .B1(n281), .C0(
        n6093), .Y(n6094) );
  OAI221X2 U3637 ( .A0(net105150), .A1(net112709), .B0(net105151), .B1(
        net112723), .C0(net105152), .Y(net99104) );
  OR2X4 U3638 ( .A(net112563), .B(n1989), .Y(n4203) );
  OR2X2 U3639 ( .A(net112693), .B(n2020), .Y(n4202) );
  NAND3BX2 U3640 ( .AN(n3731), .B(net98881), .C(net126164), .Y(n9327) );
  MX2X1 U3641 ( .A(n4799), .B(n9141), .S0(n7029), .Y(n6955) );
  AND3X2 U3642 ( .A(n8516), .B(n8515), .C(n8514), .Y(n8518) );
  CLKBUFX4 U3643 ( .A(net112107), .Y(net112085) );
  AOI2BB1X1 U3644 ( .A0N(n3576), .A1N(n7555), .B0(n6955), .Y(n6956) );
  NAND2XL U3645 ( .A(n4598), .B(n7200), .Y(n6858) );
  INVX20 U3646 ( .A(n7050), .Y(n3733) );
  CLKBUFX2 U3647 ( .A(n5403), .Y(n5399) );
  CLKBUFX2 U3648 ( .A(n5395), .Y(n5400) );
  INVX4 U3649 ( .A(n10295), .Y(n10300) );
  CLKINVX3 U3650 ( .A(net112335), .Y(net112283) );
  NAND2X8 U3651 ( .A(n3779), .B(n3780), .Y(n6099) );
  NAND3BX2 U3652 ( .AN(n7860), .B(n4924), .C(n7885), .Y(n7890) );
  INVX1 U3653 ( .A(n7706), .Y(n7857) );
  OA22X4 U3654 ( .A0(n5333), .A1(n3222), .B0(n5290), .B1(n1583), .Y(n6019) );
  OAI221X4 U3655 ( .A0(\i_MIPS/Register/register[18][3] ), .A1(n4921), .B0(
        \i_MIPS/Register/register[26][3] ), .B1(n4917), .C0(n8755), .Y(n8758)
         );
  INVX4 U3656 ( .A(n7090), .Y(n7182) );
  MX2XL U3657 ( .A(n3497), .B(net99555), .S0(n5506), .Y(\i_MIPS/n405 ) );
  OAI211X2 U3658 ( .A0(n8515), .A1(n8513), .B0(n8516), .C0(n8514), .Y(n7801)
         );
  NAND3BX2 U3659 ( .AN(n7962), .B(n4928), .C(n7981), .Y(n7986) );
  AO22X2 U3660 ( .A0(mem_rdata_I[30]), .A1(n113), .B0(n5466), .B1(n11260), .Y(
        n9798) );
  AO22X2 U3661 ( .A0(mem_rdata_I[62]), .A1(n113), .B0(n5466), .B1(n11292), .Y(
        n9803) );
  AO22X2 U3662 ( .A0(mem_rdata_I[94]), .A1(n113), .B0(n5466), .B1(n11324), .Y(
        n9793) );
  AO22X2 U3663 ( .A0(mem_rdata_I[71]), .A1(n115), .B0(n5466), .B1(n11301), .Y(
        n9815) );
  AO22X2 U3664 ( .A0(mem_rdata_I[7]), .A1(n113), .B0(n5466), .B1(n11237), .Y(
        n9830) );
  AO22X2 U3665 ( .A0(mem_rdata_I[118]), .A1(n113), .B0(n5466), .B1(n11348), 
        .Y(n9843) );
  CLKBUFX2 U3666 ( .A(n3767), .Y(n3724) );
  AND3XL U3667 ( .A(n6446), .B(n3706), .C(n6444), .Y(n6498) );
  NAND4BX4 U3668 ( .AN(n8283), .B(n8922), .C(n9258), .D(n8282), .Y(n8284) );
  AO22X4 U3669 ( .A0(net113457), .A1(n11441), .B0(net113463), .B1(n11410), .Y(
        n8119) );
  INVX20 U3670 ( .A(n3725), .Y(net98430) );
  AOI222X2 U3671 ( .A0(n5486), .A1(n11436), .B0(mem_rdata_D[48]), .B1(n117), 
        .C0(n12981), .C1(n5482), .Y(n10459) );
  NAND4X4 U3672 ( .A(n8194), .B(n8193), .C(n8192), .D(n8191), .Y(n11436) );
  AND3X8 U3673 ( .A(n6447), .B(n4471), .C(n3686), .Y(n3727) );
  MX2X1 U3674 ( .A(n8422), .B(n8421), .S0(net108959), .Y(n8425) );
  AOI21X4 U3675 ( .A0(n9287), .A1(n7875), .B0(n7873), .Y(n4569) );
  OAI2BB1X4 U3676 ( .A0N(n8163), .A1N(n8150), .B0(n8151), .Y(n7711) );
  CLKBUFX4 U3677 ( .A(n4480), .Y(n4931) );
  OA22X1 U3678 ( .A0(n5346), .A1(n979), .B0(n5302), .B1(n2525), .Y(n9827) );
  NAND2XL U3679 ( .A(n11168), .B(net100095), .Y(n4626) );
  NAND2X6 U3680 ( .A(n6570), .B(\i_MIPS/ALUin1[15] ), .Y(n7042) );
  AOI2BB1X1 U3681 ( .A0N(\i_MIPS/n356 ), .A1N(n4806), .B0(n4689), .Y(n7040) );
  OAI221X4 U3682 ( .A0(\i_MIPS/n359 ), .A1(n4824), .B0(\i_MIPS/n358 ), .B1(
        n4816), .C0(n7040), .Y(n8262) );
  OA22X4 U3683 ( .A0(n7869), .A1(n7474), .B0(n8262), .B1(n4797), .Y(n7041) );
  NOR2BX4 U3684 ( .AN(n4814), .B(n6947), .Y(n4689) );
  AO22X1 U3685 ( .A0(n8527), .A1(n9259), .B0(n9258), .B1(n4801), .Y(n6941) );
  NAND2X1 U3686 ( .A(n8897), .B(n8891), .Y(n8282) );
  OAI211X2 U3687 ( .A0(n8893), .A1(n8892), .B0(n8891), .C0(n8890), .Y(n8900)
         );
  BUFX8 U3688 ( .A(n4982), .Y(n4986) );
  AND2XL U3689 ( .A(net99935), .B(net99936), .Y(n4561) );
  AOI2BB2X4 U3690 ( .B0(n3735), .B1(\D_cache/cache[7][144] ), .A0N(net112091), 
        .A1N(n1899), .Y(n6061) );
  INVX12 U3691 ( .A(n7096), .Y(n6462) );
  OA22XL U3692 ( .A0(n5444), .A1(n1053), .B0(n5398), .B1(n2625), .Y(n10096) );
  AND4X4 U3693 ( .A(n6440), .B(n6439), .C(n6438), .D(n6437), .Y(n6441) );
  NAND2BX2 U3694 ( .AN(n8815), .B(n7615), .Y(n3782) );
  INVX8 U3695 ( .A(n8539), .Y(n8263) );
  NOR3BX4 U3696 ( .AN(n4161), .B(n3737), .C(n3738), .Y(n3736) );
  NOR2X2 U3697 ( .A(net112561), .B(n1893), .Y(n3737) );
  OR2X2 U3698 ( .A(n3611), .B(n2021), .Y(n4152) );
  NAND2X8 U3699 ( .A(n4754), .B(n3760), .Y(n3761) );
  AOI222X2 U3700 ( .A0(n5475), .A1(n11503), .B0(mem_rdata_D[117]), .B1(n117), 
        .C0(n12976), .C1(n5473), .Y(n10533) );
  AND2XL U3701 ( .A(n3707), .B(n165), .Y(n7120) );
  OAI31X4 U3702 ( .A0(n6227), .A1(n3704), .A2(n3773), .B0(n165), .Y(n6347) );
  INVX1 U3703 ( .A(n7100), .Y(n6465) );
  NAND3BX4 U3704 ( .AN(n8529), .B(n8070), .C(n8069), .Y(n8078) );
  OAI221X2 U3705 ( .A0(net112651), .A1(n2043), .B0(net112575), .B1(n703), .C0(
        n6038), .Y(n6039) );
  CLKBUFX2 U3706 ( .A(net112593), .Y(net112555) );
  INVXL U3707 ( .A(n7452), .Y(n3739) );
  INVX3 U3708 ( .A(n3739), .Y(n3740) );
  INVX1 U3709 ( .A(n8812), .Y(n3741) );
  INVX1 U3710 ( .A(n3197), .Y(n8812) );
  NAND2X8 U3711 ( .A(n4500), .B(n4654), .Y(n4479) );
  CLKMX2X2 U3712 ( .A(n4799), .B(n9141), .S0(n3634), .Y(n7478) );
  MX2XL U3713 ( .A(n3671), .B(net99461), .S0(n5509), .Y(\i_MIPS/n464 ) );
  MXI2X4 U3714 ( .A(n3743), .B(n3742), .S0(n5594), .Y(n6231) );
  MX2XL U3715 ( .A(n12958), .B(net99016), .S0(n5510), .Y(\i_MIPS/n457 ) );
  AO22X2 U3716 ( .A0(n6248), .A1(n9259), .B0(n9258), .B1(n6347), .Y(n6252) );
  CLKINVX3 U3717 ( .A(n6348), .Y(n6248) );
  AO22X4 U3718 ( .A0(net113041), .A1(net98994), .B0(net102300), .B1(n6415), 
        .Y(net107011) );
  NAND3BX4 U3719 ( .AN(n4503), .B(n3673), .C(n4424), .Y(n11137) );
  OA22X4 U3720 ( .A0(n5249), .A1(n1941), .B0(n5204), .B1(n363), .Y(n6009) );
  OAI221X4 U3721 ( .A0(n8730), .A1(n3591), .B0(n8724), .B1(n8539), .C0(n7110), 
        .Y(n7114) );
  AOI222X2 U3722 ( .A0(n9140), .A1(n7787), .B0(n7109), .B1(n3636), .C0(n8821), 
        .C1(n4547), .Y(n7110) );
  OAI221X2 U3723 ( .A0(net100082), .A1(n322), .B0(net112145), .B1(n3248), .C0(
        n6113), .Y(n6114) );
  BUFX20 U3724 ( .A(net100079), .Y(net111979) );
  MX2X2 U3725 ( .A(n7283), .B(n7693), .S0(n5590), .Y(n7284) );
  OAI221X4 U3726 ( .A0(\i_MIPS/n369 ), .A1(n4825), .B0(\i_MIPS/n368 ), .B1(
        n4817), .C0(n6358), .Y(n7283) );
  MX2XL U3727 ( .A(n3498), .B(n3659), .S0(n5508), .Y(\i_MIPS/n397 ) );
  OAI221X2 U3728 ( .A0(\i_MIPS/n347 ), .A1(n4825), .B0(\i_MIPS/n348 ), .B1(
        n4818), .C0(n6354), .Y(n6851) );
  OAI221X4 U3729 ( .A0(n4517), .A1(n8729), .B0(n3576), .B1(n7471), .C0(n4501), 
        .Y(n7050) );
  NAND2BX4 U3730 ( .AN(n5458), .B(n11238), .Y(n9684) );
  NAND3X4 U3731 ( .A(n4503), .B(n4423), .C(n9428), .Y(n4450) );
  NAND2BX4 U3732 ( .AN(n5456), .B(n11240), .Y(n9675) );
  AO22XL U3733 ( .A0(ICACHE_addr[23]), .A1(mem_read_I), .B0(n4796), .B1(n11382), .Y(n12827) );
  OR3X4 U3734 ( .A(n9581), .B(n9550), .C(n9549), .Y(n3852) );
  AOI32X2 U3735 ( .A0(n7615), .A1(\i_MIPS/ALUin1[1] ), .A2(n4809), .B0(n7614), 
        .B1(\i_MIPS/ALUin1[1] ), .Y(n7616) );
  OA22X4 U3736 ( .A0(n5428), .A1(n1942), .B0(n5384), .B1(n364), .Y(n6011) );
  BUFX4 U3737 ( .A(n5384), .Y(n5387) );
  AO22XL U3738 ( .A0(ICACHE_addr[22]), .A1(mem_read_I), .B0(n4796), .B1(n11381), .Y(n12828) );
  NAND2X4 U3739 ( .A(\i_MIPS/ALUin1[27] ), .B(n6615), .Y(n9169) );
  CLKAND2X2 U3740 ( .A(n9169), .B(n8646), .Y(n4594) );
  CLKINVX1 U3741 ( .A(n3792), .Y(n3744) );
  NAND2X8 U3742 ( .A(n3788), .B(\i_MIPS/n366 ), .Y(n7271) );
  NAND2X8 U3743 ( .A(n3761), .B(n3762), .Y(n6156) );
  OA22X2 U3744 ( .A0(net112511), .A1(n451), .B0(net112379), .B1(n2007), .Y(
        n6142) );
  AOI221XL U3745 ( .A0(net112213), .A1(\D_cache/cache[4][128] ), .B0(net112123), .B1(\D_cache/cache[5][128] ), .C0(n3829), .Y(n3745) );
  OAI221X1 U3746 ( .A0(\i_MIPS/Register/register[18][0] ), .A1(n4944), .B0(
        \i_MIPS/Register/register[26][0] ), .B1(n4942), .C0(n6520), .Y(n6523)
         );
  OA22X2 U3747 ( .A0(\i_MIPS/Register/register[22][0] ), .A1(n4935), .B0(
        \i_MIPS/Register/register[30][0] ), .B1(n4929), .Y(n6520) );
  NAND2X1 U3748 ( .A(n4660), .B(n4582), .Y(n4482) );
  AND2X8 U3749 ( .A(\i_MIPS/n316 ), .B(\i_MIPS/n318 ), .Y(n4582) );
  CLKAND2X6 U3750 ( .A(n4663), .B(n9547), .Y(n4613) );
  CLKAND2X12 U3751 ( .A(n4470), .B(n6660), .Y(n4632) );
  NOR4X4 U3752 ( .A(n8878), .B(n8877), .C(n8876), .D(n8875), .Y(n8879) );
  NAND2X4 U3753 ( .A(n6619), .B(n6630), .Y(n6649) );
  OAI211X4 U3754 ( .A0(n6618), .A1(n8071), .B0(n8520), .C0(n8067), .Y(n7958)
         );
  OA22X2 U3755 ( .A0(net112041), .A1(n452), .B0(net111915), .B1(n2008), .Y(
        n6143) );
  NAND3BX1 U3756 ( .AN(n4413), .B(n6209), .C(n6216), .Y(n6212) );
  NAND2BX1 U3757 ( .AN(net113725), .B(n11455), .Y(n4055) );
  INVX12 U3758 ( .A(n9550), .Y(n9579) );
  OAI2BB2X1 U3759 ( .B0(\i_MIPS/n174 ), .B1(net110215), .A0N(n174), .A1N(
        n10368), .Y(\i_MIPS/N115 ) );
  OAI31X4 U3760 ( .A0(\i_MIPS/ALUin1[30] ), .A1(n11223), .A2(n11222), .B0(
        n11221), .Y(n11582) );
  NAND2X1 U3761 ( .A(n3575), .B(n6451), .Y(n8804) );
  AND3X8 U3762 ( .A(n4433), .B(n8335), .C(n4432), .Y(n3749) );
  OAI222X2 U3763 ( .A0(n8142), .A1(n4797), .B0(n7867), .B1(n8542), .C0(n4707), 
        .C1(n8541), .Y(n9001) );
  MX2X6 U3764 ( .A(n6776), .B(n4684), .S0(n5590), .Y(n8541) );
  AO21XL U3765 ( .A0(\i_MIPS/ID_EX[88] ), .A1(n5517), .B0(n4499), .Y(
        \i_MIPS/n497 ) );
  INVX20 U3766 ( .A(n9262), .Y(n9259) );
  XNOR2X1 U3767 ( .A(n6293), .B(\i_MIPS/IR_ID[17] ), .Y(n4703) );
  AOI2BB1X4 U3768 ( .A0N(\i_MIPS/n365 ), .A1N(n4819), .B0(n4667), .Y(n6256) );
  INVX8 U3769 ( .A(n7546), .Y(n6455) );
  OA22X4 U3770 ( .A0(net112443), .A1(n1943), .B0(n3688), .B1(n365), .Y(n6082)
         );
  OA22X4 U3771 ( .A0(n5429), .A1(n1944), .B0(n5385), .B1(n366), .Y(n6028) );
  BUFX16 U3772 ( .A(n4723), .Y(n3815) );
  AND2X8 U3773 ( .A(n3524), .B(n9272), .Y(n4627) );
  NAND3BX4 U3774 ( .AN(n3672), .B(n3752), .C(net113533), .Y(n3753) );
  BUFX12 U3775 ( .A(net134088), .Y(net112105) );
  CLKBUFX6 U3776 ( .A(net134088), .Y(net112107) );
  INVX3 U3777 ( .A(n10391), .Y(n10385) );
  AND3X8 U3778 ( .A(n6236), .B(n8711), .C(n8803), .Y(n3754) );
  AND2XL U3779 ( .A(n11075), .B(n11073), .Y(n4521) );
  OA22X1 U3780 ( .A0(n7628), .A1(n8817), .B0(n7627), .B1(n7626), .Y(n7629) );
  INVX1 U3781 ( .A(n6108), .Y(n10641) );
  OAI22X4 U3782 ( .A0(n11582), .A1(n11581), .B0(n4591), .B1(n11582), .Y(n11583) );
  INVX12 U3783 ( .A(n3686), .Y(n6263) );
  NAND2X4 U3784 ( .A(n285), .B(n3756), .Y(n3757) );
  INVX3 U3785 ( .A(n6144), .Y(n3756) );
  INVX6 U3786 ( .A(n6083), .Y(n10651) );
  NAND3BX4 U3787 ( .AN(n4503), .B(n4423), .C(n9428), .Y(n11138) );
  CLKBUFX4 U3788 ( .A(net100084), .Y(net112519) );
  OA22X2 U3789 ( .A0(net112477), .A1(n929), .B0(net112353), .B1(n2453), .Y(
        n7926) );
  OA22X4 U3790 ( .A0(net112089), .A1(n1945), .B0(net111915), .B1(n367), .Y(
        n6150) );
  BUFX16 U3791 ( .A(net112705), .Y(net112695) );
  NAND2X4 U3792 ( .A(n12945), .B(n6155), .Y(n3762) );
  INVX3 U3793 ( .A(n6155), .Y(n3760) );
  OR2XL U3794 ( .A(\i_MIPS/PC/n19 ), .B(net110213), .Y(n3763) );
  NOR2X8 U3795 ( .A(n6447), .B(n4067), .Y(n4567) );
  OAI221X4 U3796 ( .A0(n9137), .A1(n9136), .B0(n9135), .B1(n9275), .C0(n9134), 
        .Y(n9189) );
  OAI221X4 U3797 ( .A0(\i_MIPS/ALUin1[20] ), .A1(n4824), .B0(
        \i_MIPS/ALUin1[21] ), .B1(n4816), .C0(n8271), .Y(n8642) );
  AO22X2 U3798 ( .A0(mem_rdata_I[28]), .A1(n114), .B0(n5465), .B1(n11258), .Y(
        n9774) );
  AO22X2 U3799 ( .A0(mem_rdata_I[60]), .A1(n114), .B0(n5467), .B1(n11290), .Y(
        n9779) );
  AO22X2 U3800 ( .A0(mem_rdata_I[126]), .A1(n114), .B0(n5467), .B1(n11356), 
        .Y(n9788) );
  AO22X2 U3801 ( .A0(mem_rdata_I[27]), .A1(n114), .B0(n5467), .B1(n11257), .Y(
        n9730) );
  AO22X2 U3802 ( .A0(mem_rdata_I[59]), .A1(n113), .B0(n5467), .B1(n11289), .Y(
        n9735) );
  BUFX4 U3803 ( .A(net112505), .Y(net112461) );
  BUFX4 U3804 ( .A(net112505), .Y(net112457) );
  NAND4X4 U3805 ( .A(n6967), .B(n6966), .C(n6965), .D(n6964), .Y(n11403) );
  NAND3BX1 U3806 ( .AN(n9335), .B(n4697), .C(n4696), .Y(n9339) );
  AOI2BB1XL U3807 ( .A0N(n10214), .A1N(n10205), .B0(n4521), .Y(n10220) );
  AO21X4 U3808 ( .A0(n9168), .A1(n9167), .B0(n9166), .Y(n9175) );
  CLKINVX6 U3809 ( .A(n6588), .Y(n6583) );
  CLKINVX3 U3810 ( .A(net112497), .Y(net112403) );
  OR2XL U3811 ( .A(n6244), .B(\i_MIPS/ALUin1[10] ), .Y(n3766) );
  OAI221X2 U3812 ( .A0(net112659), .A1(n1882), .B0(net112583), .B1(n316), .C0(
        n6119), .Y(n6120) );
  OA21X4 U3813 ( .A0(n6650), .A1(n6418), .B0(n8333), .Y(n6420) );
  NAND2X4 U3814 ( .A(n6594), .B(\i_MIPS/n345 ), .Y(n8333) );
  AOI2BB1X4 U3815 ( .A0N(n6652), .A1N(n6420), .B0(n6419), .Y(n6421) );
  INVX1 U3816 ( .A(n8647), .Y(n6419) );
  BUFX8 U3817 ( .A(net112583), .Y(net112573) );
  AO22X4 U3818 ( .A0(net113445), .A1(n11472), .B0(net102346), .B1(n11503), .Y(
        n8118) );
  BUFX4 U3819 ( .A(net112517), .Y(net112431) );
  OA21X4 U3820 ( .A0(n9010), .A1(n9286), .B0(n9008), .Y(n3783) );
  AOI2BB1X4 U3821 ( .A0N(\i_MIPS/n343 ), .A1N(n4806), .B0(n4673), .Y(n6223) );
  NOR2X8 U3822 ( .A(n7960), .B(n6631), .Y(n3767) );
  NAND2X2 U3823 ( .A(\i_MIPS/ALUin1[21] ), .B(n6584), .Y(n8068) );
  INVX4 U3824 ( .A(n8068), .Y(n6631) );
  INVX3 U3825 ( .A(n7286), .Y(n7612) );
  MX2XL U3826 ( .A(n3499), .B(net99354), .S0(n5510), .Y(\i_MIPS/n389 ) );
  CLKBUFX2 U3827 ( .A(n5363), .Y(n5328) );
  OAI221X4 U3828 ( .A0(net112697), .A1(n1226), .B0(net112585), .B1(n2805), 
        .C0(n6048), .Y(n6049) );
  NAND2X6 U3829 ( .A(n8260), .B(n7698), .Y(n8437) );
  INVX12 U3830 ( .A(n4722), .Y(n5593) );
  MX2XL U3831 ( .A(n3490), .B(n3705), .S0(n5507), .Y(\i_MIPS/n399 ) );
  OA22X4 U3832 ( .A0(\i_MIPS/n349 ), .A1(n4812), .B0(\i_MIPS/n350 ), .B1(n4805), .Y(n6354) );
  BUFX12 U3833 ( .A(net100079), .Y(net111983) );
  AOI222X2 U3834 ( .A0(n4554), .A1(n7365), .B0(n7363), .B1(n7362), .C0(n7361), 
        .C1(n7360), .Y(n7371) );
  INVX4 U3835 ( .A(n6426), .Y(n8149) );
  NAND2X4 U3836 ( .A(n4583), .B(n4581), .Y(n9226) );
  AOI221X2 U3837 ( .A0(net112217), .A1(\D_cache/cache[4][145] ), .B0(net112123), .B1(\D_cache/cache[5][145] ), .C0(n3775), .Y(n3774) );
  OAI22X1 U3838 ( .A0(net112041), .A1(n3288), .B0(net111917), .B1(n439), .Y(
        n3775) );
  BUFX20 U3839 ( .A(net112259), .Y(net112231) );
  MX2X8 U3840 ( .A(\i_MIPS/n271 ), .B(n4645), .S0(n3771), .Y(n6577) );
  INVXL U3841 ( .A(n3311), .Y(n3776) );
  CLKINVX1 U3842 ( .A(n3776), .Y(n3777) );
  NAND3BX2 U3843 ( .AN(n4689), .B(n6359), .C(n6352), .Y(n6855) );
  OAI221X4 U3844 ( .A0(\i_MIPS/ALUin1[12] ), .A1(n4825), .B0(
        \i_MIPS/ALUin1[11] ), .B1(n4817), .C0(n6854), .Y(n7269) );
  OAI211X4 U3845 ( .A0(n7650), .A1(n7649), .B0(net113439), .C0(net112607), .Y(
        n10829) );
  NAND4X2 U3846 ( .A(n8367), .B(n8366), .C(n8365), .D(n8364), .Y(n8372) );
  OAI221X4 U3847 ( .A0(\i_MIPS/Register/register[2][26] ), .A1(n4923), .B0(
        \i_MIPS/Register/register[10][26] ), .B1(n4917), .C0(n8368), .Y(n8371)
         );
  CLKMX2X6 U3848 ( .A(n3820), .B(n3525), .S0(n3815), .Y(n3821) );
  INVX4 U3849 ( .A(n6081), .Y(n3778) );
  NAND2XL U3850 ( .A(n3677), .B(n10675), .Y(n11520) );
  OA22X2 U3851 ( .A0(net112073), .A1(n930), .B0(net111949), .B1(n2454), .Y(
        n8582) );
  CLKMX2X6 U3852 ( .A(\i_MIPS/n295 ), .B(n177), .S0(n3815), .Y(n6242) );
  AO21X2 U3853 ( .A0(net99288), .A1(net99289), .B0(net113077), .Y(net99270) );
  NAND2XL U3854 ( .A(net99288), .B(net99289), .Y(n10607) );
  OAI211X4 U3855 ( .A0(n7929), .A1(n7928), .B0(net113439), .C0(net112609), .Y(
        net99289) );
  OA21X4 U3856 ( .A0(n6421), .A1(n6443), .B0(n11583), .Y(n6422) );
  NAND2X2 U3857 ( .A(n11110), .B(net113551), .Y(n10937) );
  MXI2X4 U3858 ( .A(n7543), .B(n7196), .S0(n5589), .Y(n4593) );
  OAI221X4 U3859 ( .A0(\i_MIPS/ALUin1[11] ), .A1(n4810), .B0(
        \i_MIPS/ALUin1[10] ), .B1(n4803), .C0(n7195), .Y(n7543) );
  OA21X2 U3860 ( .A0(\i_MIPS/ALUin1[12] ), .A1(n4818), .B0(n8141), .Y(n7195)
         );
  MX2XL U3861 ( .A(n3491), .B(n182), .S0(n5509), .Y(\i_MIPS/n431 ) );
  AOI31X2 U3862 ( .A0(n6471), .A1(n3670), .A2(n7463), .B0(n6470), .Y(n6482) );
  NAND2X4 U3863 ( .A(\i_MIPS/ALUin1[7] ), .B(n6242), .Y(n7463) );
  NAND2X4 U3864 ( .A(n4659), .B(n4582), .Y(n6509) );
  OA22XL U3865 ( .A0(\i_MIPS/Register/register[1][27] ), .A1(n4834), .B0(
        \i_MIPS/Register/register[9][27] ), .B1(n4829), .Y(n8623) );
  OA22XL U3866 ( .A0(\i_MIPS/Register/register[1][25] ), .A1(n4834), .B0(
        \i_MIPS/Register/register[9][25] ), .B1(n4830), .Y(n8459) );
  OA22XL U3867 ( .A0(\i_MIPS/Register/register[17][25] ), .A1(n4834), .B0(
        \i_MIPS/Register/register[25][25] ), .B1(n4829), .Y(n8468) );
  OA22XL U3868 ( .A0(\i_MIPS/Register/register[1][26] ), .A1(n4834), .B0(
        \i_MIPS/Register/register[9][26] ), .B1(n4831), .Y(n8367) );
  OA22XL U3869 ( .A0(\i_MIPS/Register/register[17][26] ), .A1(n4834), .B0(
        \i_MIPS/Register/register[25][26] ), .B1(n4830), .Y(n8376) );
  CLKBUFX2 U3870 ( .A(n4622), .Y(n4838) );
  CLKINVX12 U3871 ( .A(n4687), .Y(n3824) );
  CLKBUFX3 U3872 ( .A(n4622), .Y(n4837) );
  OR2X8 U3873 ( .A(n9166), .B(n6616), .Y(n4438) );
  CLKINVX20 U3874 ( .A(n4792), .Y(mem_addr_D[31]) );
  INVX3 U3875 ( .A(n4772), .Y(n4792) );
  AOI211X4 U3876 ( .A0(n7480), .A1(n8822), .B0(n7479), .C0(n7478), .Y(n7481)
         );
  INVX1 U3877 ( .A(n7471), .Y(n7480) );
  OAI211X2 U3878 ( .A0(n8026), .A1(n8025), .B0(net113439), .C0(n3709), .Y(
        net99406) );
  NAND4X4 U3879 ( .A(n8400), .B(n8399), .C(n8398), .D(n8397), .Y(n11508) );
  OR2X2 U3880 ( .A(net112263), .B(n2022), .Y(n4186) );
  CLKINVX8 U3881 ( .A(net113083), .Y(net113077) );
  AO22X4 U3882 ( .A0(net113447), .A1(n11454), .B0(net102346), .B1(n11485), .Y(
        n8863) );
  OR2X1 U3883 ( .A(n8817), .B(n8816), .Y(n3781) );
  NAND2X8 U3884 ( .A(n7200), .B(n5589), .Y(n8817) );
  CLKAND2X8 U3885 ( .A(net98881), .B(net99849), .Y(net131142) );
  NAND4X4 U3886 ( .A(n6268), .B(n6267), .C(n6266), .D(n6265), .Y(net99016) );
  MX2X1 U3887 ( .A(DCACHE_addr[13]), .B(net99609), .S0(n5506), .Y(
        \i_MIPS/n454 ) );
  OAI221X2 U3888 ( .A0(net112263), .A1(n1883), .B0(net112137), .B1(n317), .C0(
        n6066), .Y(n6067) );
  NAND2X4 U3889 ( .A(n3821), .B(\i_MIPS/n365 ), .Y(n7562) );
  CLKINVX1 U3890 ( .A(n9171), .Y(n9002) );
  OA22X4 U3891 ( .A0(net112503), .A1(n1947), .B0(net112377), .B1(n369), .Y(
        n6064) );
  INVX20 U3892 ( .A(n3787), .Y(n5590) );
  AOI222X1 U3893 ( .A0(n5474), .A1(n11498), .B0(mem_rdata_D[112]), .B1(n117), 
        .C0(n12981), .C1(n5472), .Y(n10450) );
  AO22XL U3894 ( .A0(n4969), .A1(n184), .B0(n4966), .B1(n203), .Y(n7839) );
  BUFX4 U3895 ( .A(n7864), .Y(n4797) );
  OA22X4 U3896 ( .A0(n7869), .A1(n7283), .B0(n8098), .B1(n4797), .Y(n6362) );
  INVX6 U3897 ( .A(n6067), .Y(n10620) );
  MX2X4 U3898 ( .A(\i_MIPS/n301 ), .B(n6216), .S0(n3815), .Y(n3789) );
  AOI222XL U3899 ( .A0(n5480), .A1(n11471), .B0(mem_rdata_D[84]), .B1(n117), 
        .C0(n12977), .C1(n5477), .Y(n10524) );
  AO21X2 U3900 ( .A0(net99637), .A1(net99638), .B0(net113075), .Y(net99634) );
  OAI221X2 U3901 ( .A0(\i_MIPS/ID_EX[73] ), .A1(n4434), .B0(\i_MIPS/ID_EX[41] ), .B1(n5594), .C0(\i_MIPS/n371 ), .Y(n6427) );
  AND2XL U3902 ( .A(n3788), .B(\i_MIPS/n366 ), .Y(n3792) );
  MX2XL U3903 ( .A(\i_MIPS/ID_EX[55] ), .B(net99576), .S0(n5506), .Y(
        \i_MIPS/n409 ) );
  AO22X4 U3904 ( .A0(net113447), .A1(n11465), .B0(net102346), .B1(n11496), .Y(
        n6976) );
  AOI222X4 U3905 ( .A0(n9139), .A1(n8083), .B0(n4800), .B1(n8082), .C0(n8081), 
        .C1(n3636), .Y(n8094) );
  OAI211XL U3906 ( .A0(\i_MIPS/ID_EX[80] ), .A1(n8732), .B0(n7281), .C0(n7280), 
        .Y(n7282) );
  AOI222X1 U3907 ( .A0(n5486), .A1(n11448), .B0(mem_rdata_D[60]), .B1(n117), 
        .C0(n12969), .C1(n5482), .Y(n10405) );
  OAI2BB2X2 U3908 ( .B0(\i_MIPS/n175 ), .B1(net110227), .A0N(n174), .A1N(
        n10385), .Y(\i_MIPS/N116 ) );
  AOI222X2 U3909 ( .A0(n8723), .A1(n3636), .B0(n8722), .B1(n8721), .C0(n8720), 
        .C1(n8719), .Y(n8741) );
  NAND2X2 U3910 ( .A(n10704), .B(n10701), .Y(n10712) );
  NAND3BX4 U3911 ( .AN(n7568), .B(n7567), .C(n7566), .Y(net98472) );
  AOI222X2 U3912 ( .A0(n4554), .A1(n7863), .B0(n7554), .B1(n7553), .C0(n7552), 
        .C1(n7551), .Y(n7567) );
  NAND2XL U3913 ( .A(n3719), .B(\i_MIPS/n367 ), .Y(n3801) );
  OA22X1 U3914 ( .A0(net112061), .A1(n1236), .B0(net111937), .B1(n2841), .Y(
        n7718) );
  AO21X4 U3915 ( .A0(net98950), .A1(net98951), .B0(net112727), .Y(net106420)
         );
  AO21X4 U3916 ( .A0(net98950), .A1(net98951), .B0(net113077), .Y(net98932) );
  NAND4X2 U3917 ( .A(n6800), .B(n6799), .C(n6798), .D(n6797), .Y(n11490) );
  OR2X8 U3918 ( .A(n8995), .B(net112721), .Y(net140424) );
  INVX3 U3919 ( .A(n9265), .Y(n9266) );
  AO21X2 U3920 ( .A0(n7785), .A1(n7874), .B0(n1891), .Y(n9265) );
  BUFX20 U3921 ( .A(n4513), .Y(n5477) );
  INVX1 U3922 ( .A(n8431), .Y(n8339) );
  INVX1 U3923 ( .A(n8803), .Y(n6449) );
  OAI31X2 U3924 ( .A0(n6460), .A1(n6459), .A2(n6458), .B0(n6457), .Y(n6471) );
  OA22X2 U3925 ( .A0(net112097), .A1(n453), .B0(net111983), .B1(n2009), .Y(
        n6052) );
  OAI211X2 U3926 ( .A0(n8599), .A1(n8598), .B0(net102344), .C0(n3709), .Y(
        net99638) );
  OA22X4 U3927 ( .A0(n4636), .A1(n3600), .B0(n9262), .B1(n6349), .Y(n6375) );
  MXI2X2 U3928 ( .A(\i_MIPS/ID_EX[72] ), .B(\i_MIPS/ID_EX[104] ), .S0(n3771), 
        .Y(n9142) );
  MXI2X2 U3929 ( .A(\i_MIPS/ID_EX[70] ), .B(\i_MIPS/ID_EX[102] ), .S0(n3771), 
        .Y(n6658) );
  NAND2X2 U3930 ( .A(n4646), .B(n3771), .Y(n4195) );
  CLKMX2X2 U3931 ( .A(\D_cache/cache[4][107] ), .B(n10785), .S0(net112213), 
        .Y(\D_cache/n936 ) );
  NAND3BX4 U3932 ( .AN(n3672), .B(net108204), .C(net113540), .Y(net100087) );
  OAI221X4 U3933 ( .A0(net112231), .A1(n2801), .B0(net112137), .B1(n735), .C0(
        n6150), .Y(n6151) );
  INVX6 U3934 ( .A(n6120), .Y(n10679) );
  OR2X8 U3935 ( .A(net105736), .B(net112723), .Y(n3803) );
  OR2X8 U3936 ( .A(n7120), .B(n7119), .Y(n3804) );
  AND2XL U3937 ( .A(n7100), .B(n7099), .Y(n7117) );
  OR2X2 U3938 ( .A(net105284), .B(net112709), .Y(n3806) );
  OR2X6 U3939 ( .A(net105285), .B(net112723), .Y(n3807) );
  NAND3X6 U3940 ( .A(n3806), .B(n3807), .C(net105286), .Y(net100044) );
  CLKMX2X2 U3941 ( .A(n3487), .B(net100044), .S0(n5509), .Y(\i_MIPS/n429 ) );
  AOI222X1 U3942 ( .A0(n5487), .A1(n11429), .B0(mem_rdata_D[41]), .B1(n116), 
        .C0(n12988), .C1(n5483), .Y(n10775) );
  BUFX20 U3943 ( .A(n4575), .Y(n5483) );
  CLKAND2X12 U3944 ( .A(n10161), .B(n352), .Y(n4575) );
  AOI2BB1X1 U3945 ( .A0N(n6462), .A1N(n6847), .B0(n6461), .Y(n6469) );
  MX2X1 U3946 ( .A(n3636), .B(n7625), .S0(n3675), .Y(n7614) );
  BUFX20 U3947 ( .A(n5276), .Y(n5319) );
  OAI211X2 U3948 ( .A0(n8305), .A1(n8304), .B0(net113439), .C0(n3709), .Y(
        net99383) );
  AOI2BB1X4 U3949 ( .A0N(n10293), .A1N(n10490), .B0(n10327), .Y(n10319) );
  OR2X8 U3950 ( .A(net103060), .B(net112721), .Y(n3810) );
  OA21X4 U3951 ( .A0(n4515), .A1(n7951), .B0(n6579), .Y(n3811) );
  NAND2X2 U3952 ( .A(n8516), .B(n8517), .Y(n7951) );
  OAI211X2 U3953 ( .A0(n8864), .A1(n8863), .B0(net113439), .C0(net112609), .Y(
        n10750) );
  AO21X4 U3954 ( .A0(n10408), .A1(n10409), .B0(net112729), .Y(n8423) );
  OR2X8 U3955 ( .A(n4088), .B(n4087), .Y(n3812) );
  AND4X4 U3956 ( .A(n7463), .B(n3747), .C(n6846), .D(n7186), .Y(n4607) );
  OAI22X2 U3957 ( .A0(n9287), .A1(n9286), .B0(n9285), .B1(n9284), .Y(n4635) );
  AND2X1 U3958 ( .A(n6603), .B(n6609), .Y(n6376) );
  MX2X1 U3959 ( .A(n9141), .B(n4799), .S0(n7091), .Y(n6861) );
  BUFX20 U3960 ( .A(n5189), .Y(n5231) );
  BUFX3 U3961 ( .A(n4910), .Y(n4912) );
  OA22X2 U3962 ( .A0(net112465), .A1(n454), .B0(net112353), .B1(n2010), .Y(
        n9251) );
  NOR2X4 U3963 ( .A(n9262), .B(n1987), .Y(n3816) );
  INVXL U3964 ( .A(n4728), .Y(n3818) );
  CLKINVX1 U3965 ( .A(n3818), .Y(n3819) );
  INVX12 U3966 ( .A(n4823), .Y(n4816) );
  INVXL U3967 ( .A(n6472), .Y(n6476) );
  XOR2X4 U3968 ( .A(n2315), .B(n6139), .Y(n6140) );
  NAND2XL U3969 ( .A(n10624), .B(n10623), .Y(n11533) );
  OA22X4 U3970 ( .A0(n5249), .A1(n1949), .B0(n5204), .B1(n371), .Y(n6013) );
  OA22X4 U3971 ( .A0(n5163), .A1(n3276), .B0(n5120), .B1(n1620), .Y(n6014) );
  XOR2X4 U3972 ( .A(n11368), .B(\i_MIPS/PC/n13 ), .Y(n4696) );
  OA22X4 U3973 ( .A0(n5333), .A1(n1950), .B0(n5290), .B1(n372), .Y(n6016) );
  OAI211X2 U3974 ( .A0(n7618), .A1(n3638), .B0(n7616), .C0(n7617), .Y(n7632)
         );
  BUFX8 U3975 ( .A(net112105), .Y(net112097) );
  BUFX8 U3976 ( .A(n4450), .Y(n5364) );
  CLKINVX20 U3977 ( .A(n4653), .Y(n3825) );
  OAI221X2 U3978 ( .A0(net112237), .A1(n2044), .B0(net112137), .B1(n704), .C0(
        n6040), .Y(n6041) );
  NAND2X8 U3979 ( .A(net99711), .B(net99712), .Y(n4099) );
  NAND3X2 U3980 ( .A(\i_MIPS/ALU_Control/n11 ), .B(\i_MIPS/n323 ), .C(n1636), 
        .Y(\i_MIPS/ALU_Control/n15 ) );
  MX2X1 U3981 ( .A(n8007), .B(n8006), .S0(n5587), .Y(n8008) );
  BUFX20 U3982 ( .A(n5365), .Y(n5361) );
  AOI32X2 U3983 ( .A0(n10347), .A1(n10346), .A2(n10352), .B0(n10345), .B1(
        n10348), .Y(n10351) );
  INVX12 U3984 ( .A(n4147), .Y(mem_addr_I[28]) );
  AO22X2 U3985 ( .A0(net113445), .A1(n11468), .B0(net102346), .B1(n11499), .Y(
        n7734) );
  INVXL U3986 ( .A(net107042), .Y(n3830) );
  OAI221X2 U3987 ( .A0(n6376), .A1(n6375), .B0(n6374), .B1(n6373), .C0(n6372), 
        .Y(net98994) );
  NAND2XL U3988 ( .A(n10639), .B(n10638), .Y(n11540) );
  NAND2BX4 U3989 ( .AN(n7455), .B(n3796), .Y(n7547) );
  NAND2XL U3990 ( .A(n3777), .B(n10630), .Y(n11541) );
  OR4X8 U3991 ( .A(n4447), .B(n4448), .C(n4446), .D(n4449), .Y(n11368) );
  OAI22X2 U3992 ( .A0(n5249), .A1(n3201), .B0(n5204), .B1(n324), .Y(n4448) );
  OAI2BB2X2 U3993 ( .B0(\i_MIPS/n178 ), .B1(net110227), .A0N(n4444), .A1N(n173), .Y(\i_MIPS/N119 ) );
  OAI2BB2X4 U3994 ( .B0(\i_MIPS/n305 ), .B1(n5594), .A0N(n5593), .A1N(
        \i_MIPS/ID_EX[75] ), .Y(n6235) );
  AOI2BB1X4 U3995 ( .A0N(n8090), .A1N(n8546), .B0(n8089), .Y(n8091) );
  NAND3BX4 U3996 ( .AN(n10507), .B(n10506), .C(n10505), .Y(n11543) );
  NAND2X4 U3997 ( .A(net110255), .B(n4543), .Y(n10506) );
  CLKAND2X8 U3998 ( .A(n4822), .B(n6947), .Y(n4615) );
  INVX8 U3999 ( .A(n6571), .Y(n6573) );
  NAND2X6 U4000 ( .A(n8151), .B(n7847), .Y(n7798) );
  AOI2BB1X4 U4001 ( .A0N(\i_MIPS/n346 ), .A1N(n4818), .B0(n4671), .Y(n7019) );
  AOI211XL U4002 ( .A0(n6665), .A1(n177), .B0(n4671), .C0(n4668), .Y(n6668) );
  INVXL U4003 ( .A(n8152), .Y(n8159) );
  NAND3BX4 U4004 ( .AN(n8451), .B(n8450), .C(n9258), .Y(n8452) );
  CLKINVX20 U4005 ( .A(n11013), .Y(n3833) );
  NAND4X4 U4006 ( .A(n6498), .B(n6497), .C(n6496), .D(n6495), .Y(net98971) );
  AO22X4 U4007 ( .A0(n7358), .A1(n9259), .B0(n9258), .B1(n7357), .Y(n7361) );
  NAND2X1 U4008 ( .A(n7272), .B(n8718), .Y(n7357) );
  XOR3X1 U4009 ( .A(net111405), .B(n10965), .C(n10964), .Y(n10967) );
  INVX8 U4010 ( .A(n7959), .Y(n6627) );
  NAND2BX4 U4011 ( .AN(n8072), .B(n8521), .Y(n7959) );
  BUFX20 U4012 ( .A(net112701), .Y(net112691) );
  AOI222X2 U4013 ( .A0(n5475), .A1(n11502), .B0(mem_rdata_D[116]), .B1(n116), 
        .C0(n12977), .C1(n5473), .Y(n10521) );
  NAND4X2 U4014 ( .A(n8597), .B(n8596), .C(n8595), .D(n8594), .Y(n11502) );
  NAND4X6 U4015 ( .A(n8453), .B(n8454), .C(n8455), .D(n8452), .Y(net99605) );
  MX2X1 U4016 ( .A(n9280), .B(n9279), .S0(n8441), .Y(n8442) );
  NOR4BX2 U4017 ( .AN(n4501), .B(n4633), .C(n4634), .D(n4635), .Y(n9288) );
  NAND2BX4 U4018 ( .AN(n6595), .B(n8346), .Y(n6596) );
  NAND2XL U4019 ( .A(n10621), .B(n10620), .Y(n11529) );
  INVX3 U4020 ( .A(net98472), .Y(net105004) );
  NOR2BX4 U4021 ( .AN(n4820), .B(\i_MIPS/n367 ), .Y(n4672) );
  NOR4X4 U4022 ( .A(n10492), .B(n10491), .C(n10490), .D(n10489), .Y(n10496) );
  AO22X4 U4023 ( .A0(n4552), .A1(n9259), .B0(n9258), .B1(n8716), .Y(n8720) );
  NAND2X2 U4024 ( .A(n10352), .B(n10349), .Y(n10334) );
  NAND2X4 U4025 ( .A(n6247), .B(n7099), .Y(n6348) );
  CLKINVX3 U4026 ( .A(net102088), .Y(net113083) );
  NAND2X4 U4027 ( .A(n10348), .B(n10362), .Y(n10353) );
  NOR3X2 U4028 ( .A(n4701), .B(n4702), .C(n4703), .Y(n6202) );
  XNOR2X1 U4029 ( .A(n10132), .B(\i_MIPS/IR_ID[18] ), .Y(n4701) );
  AND2XL U4030 ( .A(n3315), .B(net99316), .Y(n4540) );
  NAND2X4 U4031 ( .A(n9271), .B(n5589), .Y(n8546) );
  AOI222X4 U4032 ( .A0(n8667), .A1(n9271), .B0(n9139), .B1(n8666), .C0(n4547), 
        .C1(n9267), .Y(n8668) );
  INVX12 U4033 ( .A(n9004), .Y(n9271) );
  CLKINVX3 U4034 ( .A(n5266), .Y(n5242) );
  NAND2XL U4035 ( .A(n7042), .B(n7709), .Y(n7034) );
  NAND2X6 U4036 ( .A(n4587), .B(n7698), .Y(n7561) );
  NAND2XL U4037 ( .A(n3736), .B(n10668), .Y(n11535) );
  INVXL U4038 ( .A(n7181), .Y(n3837) );
  INVX3 U4039 ( .A(n3837), .Y(n3838) );
  BUFX16 U4040 ( .A(net100105), .Y(net112705) );
  AO22XL U4041 ( .A0(ICACHE_addr[17]), .A1(mem_read_I), .B0(n4796), .B1(n11376), .Y(n12833) );
  INVX20 U4042 ( .A(n4807), .Y(n4805) );
  BUFX20 U4043 ( .A(n4631), .Y(n4807) );
  AND2X8 U4044 ( .A(n9272), .B(n3525), .Y(n4631) );
  NAND2X8 U4045 ( .A(n8095), .B(n7971), .Y(n8332) );
  AND3X8 U4046 ( .A(n6767), .B(n8717), .C(n8823), .Y(n4007) );
  NAND2X4 U4047 ( .A(\i_MIPS/ALUin1[12] ), .B(n3527), .Y(n6638) );
  OAI221X2 U4048 ( .A0(net112697), .A1(n1885), .B0(net112583), .B1(n318), .C0(
        n6059), .Y(n6060) );
  INVX16 U4049 ( .A(n4428), .Y(n4722) );
  AO22X4 U4050 ( .A0(n7549), .A1(n4925), .B0(n9258), .B1(n7548), .Y(n7552) );
  BUFX20 U4051 ( .A(net111967), .Y(net111917) );
  INVX4 U4052 ( .A(n8142), .Y(n8540) );
  AOI2BB2X4 U4053 ( .B0(net113041), .B1(net99313), .A0N(net102087), .A1N(n3840), .Y(net134133) );
  AO21X4 U4054 ( .A0(net99359), .A1(net99360), .B0(net112731), .Y(net102565)
         );
  AO22X4 U4055 ( .A0(net113447), .A1(n11475), .B0(net102346), .B1(n11506), .Y(
        n8973) );
  NAND2X6 U4056 ( .A(net99386), .B(net99387), .Y(n4123) );
  AOI2BB1X4 U4057 ( .A0N(n8146), .A1N(n4520), .B0(n7798), .Y(n7799) );
  CLKBUFX20 U4058 ( .A(n9264), .Y(n4798) );
  CLKINVX20 U4059 ( .A(n4798), .Y(n9258) );
  OR2X8 U4060 ( .A(net112561), .B(n1880), .Y(n4163) );
  INVX3 U4061 ( .A(n7625), .Y(n7627) );
  BUFX20 U4062 ( .A(net110259), .Y(net110253) );
  OAI21X1 U4063 ( .A0(n4488), .A1(net112609), .B0(n11389), .Y(n10138) );
  NAND2X6 U4064 ( .A(n3553), .B(net99541), .Y(n4124) );
  INVX1 U4065 ( .A(n6673), .Y(n6366) );
  INVX3 U4066 ( .A(n6674), .Y(n6363) );
  CLKMX2X3 U4067 ( .A(n9141), .B(n4799), .S0(n7848), .Y(n7694) );
  BUFX20 U4068 ( .A(n4452), .Y(n4799) );
  OR2X8 U4069 ( .A(net112569), .B(n1881), .Y(n4205) );
  OAI221X2 U4070 ( .A0(n9264), .A1(n286), .B0(n7621), .B1(n3746), .C0(n8805), 
        .Y(n7625) );
  NAND3X6 U4071 ( .A(n4219), .B(n4220), .C(n6121), .Y(n6122) );
  INVX8 U4072 ( .A(n6122), .Y(n10678) );
  MX2XL U4073 ( .A(\i_MIPS/ID_EX[75] ), .B(\i_MIPS/Sign_Extend_ID[2] ), .S0(
        n5508), .Y(\i_MIPS/n510 ) );
  OAI2BB1X4 U4074 ( .A0N(n11048), .A1N(n11192), .B0(n11047), .Y(n11049) );
  AO22X4 U4075 ( .A0(n11046), .A1(n11045), .B0(n11044), .B1(n11043), .Y(n11192) );
  OAI2BB2XL U4076 ( .B0(\i_MIPS/n239 ), .B1(net110219), .A0N(n175), .A1N(
        n11051), .Y(\i_MIPS/N93 ) );
  NAND3BX4 U4077 ( .AN(n11006), .B(n11005), .C(n11004), .Y(\i_MIPS/PC/n37 ) );
  XNOR3X1 U4078 ( .A(net111409), .B(net99765), .C(net99753), .Y(n3847) );
  XOR2X4 U4079 ( .A(net99962), .B(ICACHE_addr[22]), .Y(net99753) );
  OR2X2 U4080 ( .A(net98430), .B(n3502), .Y(n4193) );
  NOR2BX1 U4081 ( .AN(net110227), .B(\i_MIPS/Control_ID/n12 ), .Y(n4588) );
  NAND3BX4 U4082 ( .AN(n10881), .B(n10880), .C(n10879), .Y(\i_MIPS/PC/n42 ) );
  AOI2BB1X2 U4083 ( .A0N(n10272), .A1N(n10267), .B0(n10305), .Y(n10213) );
  BUFX20 U4084 ( .A(n4513), .Y(n5478) );
  MXI2X1 U4085 ( .A(n11173), .B(n11172), .S0(n5491), .Y(n11174) );
  BUFX20 U4086 ( .A(n5485), .Y(n5486) );
  BUFX20 U4087 ( .A(n11205), .Y(n5479) );
  MXI2X6 U4088 ( .A(n10796), .B(n10795), .S0(n5490), .Y(n10797) );
  AOI222X4 U4089 ( .A0(net109795), .A1(n11401), .B0(mem_rdata_D[12]), .B1(n116), .C0(n12985), .C1(net109805), .Y(n10796) );
  MX2X1 U4090 ( .A(\D_cache/cache[0][108] ), .B(n10797), .S0(net112643), .Y(
        \D_cache/n932 ) );
  OAI211X2 U4091 ( .A0(n10353), .A1(n10352), .B0(n10351), .C0(n10350), .Y(
        n10355) );
  AOI222X4 U4092 ( .A0(n5480), .A1(n11469), .B0(mem_rdata_D[82]), .B1(n116), 
        .C0(n12979), .C1(n5477), .Y(n10612) );
  MXI2X4 U4093 ( .A(n10612), .B(n10611), .S0(n5492), .Y(n10613) );
  XNOR2X2 U4094 ( .A(n4688), .B(ICACHE_addr[18]), .Y(n11020) );
  AOI2BB1X4 U4095 ( .A0N(n10325), .A1N(n10327), .B0(n10489), .Y(n10326) );
  CLKINVX1 U4096 ( .A(n10490), .Y(n10325) );
  AND4X8 U4097 ( .A(n9587), .B(n9590), .C(n9588), .D(n9589), .Y(n3848) );
  AO22X1 U4098 ( .A0(n174), .A1(n10222), .B0(net113592), .B1(
        \i_MIPS/IR_ID[31] ), .Y(\i_MIPS/N86 ) );
  AO22X1 U4099 ( .A0(n173), .A1(n10243), .B0(net113592), .B1(
        \i_MIPS/IR_ID[30] ), .Y(\i_MIPS/N85 ) );
  CLKAND2X12 U4100 ( .A(n6660), .B(n6447), .Y(n4171) );
  OR2X8 U4101 ( .A(n11087), .B(net110247), .Y(n4191) );
  CLKAND2X8 U4102 ( .A(n4192), .B(n4193), .Y(n10815) );
  OAI222X2 U4103 ( .A0(n4524), .A1(net110241), .B0(n10732), .B1(n10698), .C0(
        \i_MIPS/PC/n31 ), .C1(net110213), .Y(n10507) );
  AOI222X4 U4104 ( .A0(n5474), .A1(n11507), .B0(mem_rdata_D[121]), .B1(n116), 
        .C0(n12972), .C1(n5472), .Y(n10424) );
  MXI2X4 U4105 ( .A(n10424), .B(n10423), .S0(n5496), .Y(n10425) );
  AOI2BB2X1 U4106 ( .B0(n10943), .B1(net110205), .A0N(net98430), .A1N(n10944), 
        .Y(n10946) );
  OAI2BB2X2 U4107 ( .B0(net110241), .B1(n3849), .A0N(ICACHE_addr[0]), .A1N(
        net113592), .Y(net98447) );
  AOI2BB2X1 U4108 ( .B0(n11019), .B1(net110205), .A0N(net98430), .A1N(n11020), 
        .Y(n11022) );
  NAND3BX4 U4109 ( .AN(n9428), .B(n4423), .C(n4503), .Y(n11140) );
  BUFX6 U4110 ( .A(n5318), .Y(n5315) );
  AOI222X4 U4111 ( .A0(n5474), .A1(n11497), .B0(mem_rdata_D[111]), .B1(n116), 
        .C0(n12982), .C1(n5472), .Y(n10187) );
  AOI222X4 U4112 ( .A0(n5488), .A1(n11421), .B0(mem_rdata_D[32]), .B1(n117), 
        .C0(n12997), .C1(n5484), .Y(n10861) );
  MXI2X4 U4113 ( .A(n10861), .B(n10860), .S0(n5499), .Y(n10862) );
  INVXL U4114 ( .A(n9211), .Y(n3851) );
  AOI2BB2X4 U4115 ( .B0(net113039), .B1(net99430), .A0N(net102087), .A1N(n3853), .Y(n3872) );
  XOR2X4 U4116 ( .A(n3854), .B(n4385), .Y(n6166) );
  CLKAND2X8 U4117 ( .A(n10658), .B(n3774), .Y(n3854) );
  OAI211X2 U4118 ( .A0(n8779), .A1(n8778), .B0(net113437), .C0(net112607), .Y(
        net100104) );
  CLKMX2X2 U4119 ( .A(DCACHE_addr[29]), .B(n3851), .S0(n5509), .Y(
        \i_MIPS/n438 ) );
  OAI211X2 U4120 ( .A0(n8119), .A1(n8118), .B0(net113439), .C0(net112609), .Y(
        net99429) );
  OAI211X2 U4121 ( .A0(n8974), .A1(n8973), .B0(net102344), .C0(net112607), .Y(
        net99360) );
  NOR4X8 U4122 ( .A(n4107), .B(n4108), .C(n4110), .D(n4109), .Y(net102398) );
  OAI221XL U4123 ( .A0(net104351), .A1(net112709), .B0(n3520), .B1(net112721), 
        .C0(net104353), .Y(net99284) );
  NAND3BX2 U4124 ( .AN(n7887), .B(n4926), .C(n7886), .Y(n7888) );
  NAND4X2 U4125 ( .A(n4928), .B(n7712), .C(n7857), .D(n7707), .Y(n7716) );
  OA22XL U4126 ( .A0(\i_MIPS/Control_ID/n15 ), .A1(net113592), .B0(n5511), 
        .B1(n4434), .Y(n9810) );
  AO22XL U4127 ( .A0(n4973), .A1(n189), .B0(n4966), .B1(n734), .Y(n7686) );
  OA22XL U4128 ( .A0(n6657), .A1(n9014), .B0(n9160), .B1(n6656), .Y(n6684) );
  NAND2X1 U4129 ( .A(n9258), .B(n6669), .Y(n6657) );
  BUFX8 U4130 ( .A(n3750), .Y(net111947) );
  OA22X4 U4131 ( .A0(\i_MIPS/n353 ), .A1(n4812), .B0(\i_MIPS/n354 ), .B1(n4805), .Y(n6353) );
  NAND2X8 U4132 ( .A(n4553), .B(n8150), .Y(n8515) );
  OAI222X2 U4133 ( .A0(n8350), .A1(n8886), .B0(n9281), .B1(n9275), .C0(n8349), 
        .C1(n8660), .Y(n8356) );
  OAI2BB2XL U4134 ( .B0(\i_MIPS/n215 ), .B1(net110221), .A0N(n173), .A1N(
        n11053), .Y(\i_MIPS/N58 ) );
  CLKAND2X12 U4135 ( .A(\i_MIPS/IR_ID[19] ), .B(\i_MIPS/n316 ), .Y(n4657) );
  MX2XL U4136 ( .A(DCACHE_addr[20]), .B(n3694), .S0(n5507), .Y(\i_MIPS/n447 )
         );
  NAND3XL U4137 ( .A(n4166), .B(n3702), .C(n9210), .Y(net99254) );
  AOI2BB1X1 U4138 ( .A0N(\i_MIPS/n368 ), .A1N(n4826), .B0(n4672), .Y(n6945) );
  NAND2X4 U4139 ( .A(net134107), .B(net100042), .Y(n4083) );
  NAND3BX4 U4140 ( .AN(n9578), .B(n4663), .C(n4695), .Y(n9585) );
  MX2XL U4141 ( .A(\i_MIPS/ID_EX[72] ), .B(net99254), .S0(n5509), .Y(
        \i_MIPS/n375 ) );
  OA22X1 U4142 ( .A0(net112077), .A1(n1237), .B0(net111953), .B1(n2842), .Y(
        n8855) );
  BUFX12 U4143 ( .A(n12837), .Y(mem_addr_I[8]) );
  OA22X4 U4144 ( .A0(net112663), .A1(n2352), .B0(net112561), .B1(n850), .Y(
        n5948) );
  INVX1 U4145 ( .A(mem_read_I), .Y(n4324) );
  NAND4BX4 U4146 ( .AN(n6576), .B(n8517), .C(n8516), .D(n6575), .Y(n6579) );
  OAI211X2 U4147 ( .A0(n8927), .A1(n8926), .B0(n8924), .C0(n8925), .Y(n3866)
         );
  INVX2 U4148 ( .A(n6848), .Y(n6770) );
  INVXL U4149 ( .A(n11053), .Y(n11058) );
  NAND3BX4 U4150 ( .AN(n7483), .B(n7482), .C(n7481), .Y(net99110) );
  NAND4X4 U4151 ( .A(n8198), .B(n8197), .C(n8196), .D(n8195), .Y(n11405) );
  CLKMX2X3 U4152 ( .A(n8619), .B(n8618), .S0(net108963), .Y(net103218) );
  OA22X2 U4153 ( .A0(net112449), .A1(n2439), .B0(net112325), .B1(n463), .Y(
        n6124) );
  AOI33X2 U4154 ( .A0(n8523), .A1(n8553), .A2(n9258), .B0(n8522), .B1(n8530), 
        .B2(n9258), .Y(n8560) );
  NAND4X4 U4155 ( .A(n7725), .B(n7724), .C(n7723), .D(n7722), .Y(n11406) );
  NAND4X2 U4156 ( .A(n9496), .B(n9495), .C(n9494), .D(n9493), .Y(n11326) );
  NAND2X6 U4157 ( .A(n6577), .B(\i_MIPS/n352 ), .Y(n7781) );
  NAND2X8 U4158 ( .A(n6569), .B(\i_MIPS/n352 ), .Y(n8071) );
  OAI221X2 U4159 ( .A0(\i_MIPS/n351 ), .A1(n4825), .B0(\i_MIPS/n352 ), .B1(
        n4818), .C0(n6353), .Y(n6852) );
  NAND4X2 U4160 ( .A(n9501), .B(n9500), .C(n9499), .D(n9498), .Y(n11294) );
  XOR2X4 U4161 ( .A(n3251), .B(n6090), .Y(n6097) );
  OAI221X4 U4162 ( .A0(n4798), .A1(n3831), .B0(n8527), .B1(n9262), .C0(n8805), 
        .Y(n6942) );
  NOR4X2 U4163 ( .A(n6820), .B(n6819), .C(n6818), .D(n6817), .Y(n6821) );
  NAND4X8 U4164 ( .A(n9834), .B(n9833), .C(n9832), .D(n9831), .Y(n10884) );
  NAND2BX4 U4165 ( .AN(n5457), .B(n11237), .Y(n9831) );
  NAND4X2 U4166 ( .A(n8589), .B(n8588), .C(n8587), .D(n8586), .Y(n11409) );
  MX2XL U4167 ( .A(n3506), .B(n181), .S0(n5511), .Y(\i_MIPS/n433 ) );
  BUFX12 U4168 ( .A(n12834), .Y(mem_addr_I[18]) );
  BUFX12 U4169 ( .A(n12833), .Y(mem_addr_I[19]) );
  BUFX12 U4170 ( .A(n12832), .Y(mem_addr_I[20]) );
  AO22X1 U4171 ( .A0(ICACHE_addr[18]), .A1(mem_read_I), .B0(n4794), .B1(n11377), .Y(n12832) );
  AOI222X4 U4172 ( .A0(n5487), .A1(n11437), .B0(mem_rdata_D[49]), .B1(n117), 
        .C0(n12980), .C1(n5483), .Y(n10605) );
  MXI2X4 U4173 ( .A(n10605), .B(n10604), .S0(n5492), .Y(n10606) );
  OAI222X2 U4174 ( .A0(\i_MIPS/PC/n26 ), .A1(net110215), .B0(net130420), .B1(
        net110241), .C0(net99760), .C1(n3602), .Y(n4136) );
  XOR3X2 U4175 ( .A(net111409), .B(net99765), .C(net99753), .Y(net99760) );
  OA22X2 U4176 ( .A0(n4139), .A1(net140281), .B0(net98430), .B1(net99753), .Y(
        n4137) );
  BUFX12 U4177 ( .A(n12831), .Y(mem_addr_I[21]) );
  AO22X1 U4178 ( .A0(ICACHE_addr[19]), .A1(mem_read_I), .B0(n4796), .B1(n11378), .Y(n12831) );
  BUFX12 U4179 ( .A(n12830), .Y(mem_addr_I[22]) );
  AO22X1 U4180 ( .A0(ICACHE_addr[20]), .A1(mem_read_I), .B0(n4796), .B1(n11379), .Y(n12830) );
  BUFX12 U4181 ( .A(n12829), .Y(mem_addr_I[23]) );
  BUFX12 U4182 ( .A(n12828), .Y(mem_addr_I[24]) );
  BUFX12 U4183 ( .A(n12827), .Y(mem_addr_I[25]) );
  NAND3X8 U4184 ( .A(n11045), .B(n9611), .C(n11048), .Y(n10306) );
  INVXL U4185 ( .A(n3317), .Y(n3881) );
  MXI2X1 U4186 ( .A(n10602), .B(n10601), .S0(n5492), .Y(n10603) );
  NAND2X4 U4187 ( .A(n6655), .B(\i_MIPS/n343 ), .Y(n9014) );
  NAND2X4 U4188 ( .A(\i_MIPS/ALUin1[28] ), .B(n6655), .Y(n9160) );
  BUFX12 U4189 ( .A(n12826), .Y(mem_addr_I[26]) );
  AO22X1 U4190 ( .A0(ICACHE_addr[24]), .A1(mem_read_I), .B0(n4796), .B1(n3589), 
        .Y(n12826) );
  AO22X2 U4191 ( .A0(n9312), .A1(n433), .B0(n4985), .B1(n1996), .Y(n8038) );
  AO22X2 U4192 ( .A0(n9312), .A1(n434), .B0(n4985), .B1(n1997), .Y(n8029) );
  AO22X2 U4193 ( .A0(n9312), .A1(n437), .B0(n4985), .B1(n2000), .Y(n7941) );
  AO22X2 U4194 ( .A0(n9312), .A1(n435), .B0(n4985), .B1(n1998), .Y(n7932) );
  AO22XL U4195 ( .A0(n9312), .A1(n487), .B0(n4985), .B1(n2231), .Y(n7684) );
  AO22XL U4196 ( .A0(n9312), .A1(n488), .B0(n4985), .B1(n2232), .Y(n7675) );
  CLKBUFX8 U4197 ( .A(n4982), .Y(n4985) );
  CLKAND2X4 U4198 ( .A(n4707), .B(n7698), .Y(n4578) );
  NAND2X8 U4199 ( .A(n4578), .B(n8148), .Y(n8736) );
  INVX1 U4200 ( .A(n6850), .Y(n6461) );
  MX2XL U4201 ( .A(n3500), .B(net99284), .S0(n5509), .Y(\i_MIPS/n401 ) );
  AOI222X1 U4202 ( .A0(net109795), .A1(n11391), .B0(mem_rdata_D[1]), .B1(n117), 
        .C0(n12996), .C1(net109805), .Y(n10845) );
  AOI222X1 U4203 ( .A0(net109795), .A1(n11402), .B0(mem_rdata_D[13]), .B1(n117), .C0(n12984), .C1(net109805), .Y(n10808) );
  AND2X1 U4204 ( .A(n12997), .B(net109805), .Y(n4180) );
  AOI222X1 U4205 ( .A0(net109795), .A1(n11397), .B0(mem_rdata_D[8]), .B1(n116), 
        .C0(n12989), .C1(net109805), .Y(n10824) );
  CLKBUFX6 U4206 ( .A(net130594), .Y(net109805) );
  NAND4X2 U4207 ( .A(n8016), .B(n8015), .C(n8014), .D(n8013), .Y(n11411) );
  NAND2BX4 U4208 ( .AN(n5452), .B(n11333), .Y(n9832) );
  INVX3 U4209 ( .A(n10363), .Y(n10364) );
  NAND4X2 U4210 ( .A(n9506), .B(n9505), .C(n9504), .D(n9503), .Y(n11230) );
  NAND4X6 U4211 ( .A(n9838), .B(n9837), .C(n9836), .D(n9835), .Y(n10873) );
  CLKINVX1 U4212 ( .A(mem_read_I), .Y(n4349) );
  AO21X4 U4213 ( .A0(n4809), .A1(\i_MIPS/ALUin1[29] ), .B0(n4682), .Y(n6356)
         );
  INVX3 U4214 ( .A(n6666), .Y(n9164) );
  NAND2X1 U4215 ( .A(n6658), .B(\i_MIPS/n342 ), .Y(n6666) );
  MX2XL U4216 ( .A(n3633), .B(n3881), .S0(n5510), .Y(\i_MIPS/n415 ) );
  MX2XL U4217 ( .A(n12953), .B(net99313), .S0(n5510), .Y(\i_MIPS/n452 ) );
  BUFX12 U4218 ( .A(n12938), .Y(mem_wdata_I[1]) );
  AND2XL U4219 ( .A(n4796), .B(n11231), .Y(n12938) );
  BUFX12 U4220 ( .A(n12937), .Y(mem_wdata_I[2]) );
  AND2XL U4221 ( .A(n4796), .B(n11232), .Y(n12937) );
  BUFX12 U4222 ( .A(n12936), .Y(mem_wdata_I[3]) );
  AND2XL U4223 ( .A(n11547), .B(n11233), .Y(n12936) );
  AOI2BB1X4 U4224 ( .A0N(n8073), .A1N(n7959), .B0(n7958), .Y(n7960) );
  OAI221X4 U4225 ( .A0(\i_MIPS/Register/register[18][18] ), .A1(n4922), .B0(
        \i_MIPS/Register/register[26][18] ), .B1(n4915), .C0(n7905), .Y(n7908)
         );
  BUFX16 U4226 ( .A(n4919), .Y(n4922) );
  NAND4X2 U4227 ( .A(n7904), .B(n7903), .C(n7902), .D(n7901), .Y(n7909) );
  OAI32X2 U4228 ( .A0(n3838), .A1(n3817), .A2(n7182), .B0(n3817), .B1(n7179), 
        .Y(n7092) );
  AOI2BB2X2 U4229 ( .B0(\i_MIPS/IF_ID[79] ), .B1(n149), .A0N(net110189), .A1N(
        \i_MIPS/n194 ), .Y(n10286) );
  AO22XL U4230 ( .A0(n4898), .A1(n489), .B0(n4893), .B1(n2233), .Y(n8370) );
  AO22X4 U4231 ( .A0(n4898), .A1(n327), .B0(n4893), .B1(n1904), .Y(n8244) );
  AO22X4 U4232 ( .A0(n4898), .A1(n328), .B0(n4893), .B1(n1905), .Y(n8235) );
  AO22X4 U4233 ( .A0(n4898), .A1(n329), .B0(n4893), .B1(n1906), .Y(n8177) );
  AO22X4 U4234 ( .A0(n4898), .A1(n330), .B0(n4893), .B1(n1907), .Y(n8186) );
  AO22X4 U4235 ( .A0(n4898), .A1(n331), .B0(n4893), .B1(n1908), .Y(n8379) );
  AO22X4 U4236 ( .A0(n4898), .A1(n429), .B0(n4893), .B1(n1992), .Y(n8462) );
  AO22X4 U4237 ( .A0(n4898), .A1(n346), .B0(n4893), .B1(n1928), .Y(n8471) );
  AO21X4 U4238 ( .A0(net100103), .A1(net100104), .B0(net112729), .Y(net102901)
         );
  OA22X2 U4239 ( .A0(n5162), .A1(n455), .B0(n5119), .B1(n3240), .Y(n5994) );
  BUFX12 U4240 ( .A(n4889), .Y(n4892) );
  CLKBUFX2 U4241 ( .A(n9115), .Y(n4889) );
  NAND4X2 U4242 ( .A(n7376), .B(n7375), .C(n7374), .D(n7373), .Y(n7381) );
  NAND2X1 U4243 ( .A(n8263), .B(n7693), .Y(n6857) );
  OAI211X2 U4244 ( .A0(n8350), .A1(n141), .B0(n7202), .C0(n7201), .Y(n7203) );
  BUFX12 U4245 ( .A(n12935), .Y(mem_wdata_I[8]) );
  AND2XL U4246 ( .A(n4794), .B(n11238), .Y(n12935) );
  BUFX12 U4247 ( .A(n12896), .Y(mem_wdata_I[54]) );
  AND2XL U4248 ( .A(n4795), .B(n11284), .Y(n12896) );
  BUFX12 U4249 ( .A(n12934), .Y(mem_wdata_I[9]) );
  AND2XL U4250 ( .A(n4796), .B(n11239), .Y(n12934) );
  BUFX12 U4251 ( .A(n12893), .Y(mem_wdata_I[57]) );
  AND2XL U4252 ( .A(n4795), .B(n11287), .Y(n12893) );
  BUFX12 U4253 ( .A(n12890), .Y(mem_wdata_I[60]) );
  AND2XL U4254 ( .A(n4795), .B(n11290), .Y(n12890) );
  AND3X4 U4255 ( .A(n4661), .B(n9570), .C(n4640), .Y(n9589) );
  AO21X4 U4256 ( .A0(n10935), .A1(n11105), .B0(n10330), .Y(n11011) );
  BUFX12 U4257 ( .A(n12933), .Y(mem_wdata_I[10]) );
  AND2XL U4258 ( .A(n4796), .B(n11240), .Y(n12933) );
  OA22X4 U4259 ( .A0(net112237), .A1(n2367), .B0(net112163), .B1(n864), .Y(
        n6386) );
  BUFX12 U4260 ( .A(n12932), .Y(mem_wdata_I[11]) );
  AND2XL U4261 ( .A(n4794), .B(n11241), .Y(n12932) );
  OA22X1 U4262 ( .A0(n5164), .A1(n1238), .B0(n5121), .B1(n2843), .Y(n9350) );
  BUFX12 U4263 ( .A(n12931), .Y(mem_wdata_I[12]) );
  AND2XL U4264 ( .A(n4796), .B(n11242), .Y(n12931) );
  OA22X2 U4265 ( .A0(n9007), .A1(n9006), .B0(n9005), .B1(n9004), .Y(n9008) );
  BUFX12 U4266 ( .A(n12930), .Y(mem_wdata_I[13]) );
  AND2XL U4267 ( .A(n4796), .B(n11243), .Y(n12930) );
  AOI32X2 U4268 ( .A0(n8156), .A1(n8157), .A2(n8159), .B0(n8155), .B1(n8154), 
        .Y(n8161) );
  OAI221X2 U4269 ( .A0(net103869), .A1(net112707), .B0(n3547), .B1(net112721), 
        .C0(net103871), .Y(net99555) );
  AOI222X1 U4270 ( .A0(n5475), .A1(n11504), .B0(mem_rdata_D[118]), .B1(n117), 
        .C0(n12975), .C1(n5473), .Y(n10545) );
  NAND4X2 U4271 ( .A(n8024), .B(n8023), .C(n8022), .D(n8021), .Y(n11504) );
  BUFX12 U4272 ( .A(n12929), .Y(mem_wdata_I[14]) );
  AND2XL U4273 ( .A(n4794), .B(n11244), .Y(n12929) );
  OA22X2 U4274 ( .A0(n11196), .A1(net140280), .B0(net98430), .B1(n3516), .Y(
        n11198) );
  BUFX12 U4275 ( .A(n12928), .Y(mem_wdata_I[15]) );
  AND2XL U4276 ( .A(n4794), .B(n11245), .Y(n12928) );
  BUFX12 U4277 ( .A(n12887), .Y(mem_wdata_I[63]) );
  AND2XL U4278 ( .A(n4795), .B(n11293), .Y(n12887) );
  BUFX12 U4279 ( .A(n12927), .Y(mem_wdata_I[16]) );
  AND2XL U4280 ( .A(n4796), .B(n11246), .Y(n12927) );
  BUFX12 U4281 ( .A(n12899), .Y(mem_wdata_I[49]) );
  AND2XL U4282 ( .A(n4796), .B(n11279), .Y(n12899) );
  BUFX12 U4283 ( .A(n12884), .Y(mem_wdata_I[66]) );
  AND2XL U4284 ( .A(n4795), .B(n11296), .Y(n12884) );
  BUFX12 U4285 ( .A(n12926), .Y(mem_wdata_I[17]) );
  AND2XL U4286 ( .A(n4794), .B(n11247), .Y(n12926) );
  BUFX12 U4287 ( .A(n12925), .Y(mem_wdata_I[18]) );
  AND2XL U4288 ( .A(n4794), .B(n11248), .Y(n12925) );
  BUFX12 U4289 ( .A(n12924), .Y(mem_wdata_I[19]) );
  AND2XL U4290 ( .A(n4796), .B(n11249), .Y(n12924) );
  BUFX12 U4291 ( .A(n12923), .Y(mem_wdata_I[20]) );
  AND2XL U4292 ( .A(n4796), .B(n11250), .Y(n12923) );
  BUFX12 U4293 ( .A(n12922), .Y(mem_wdata_I[21]) );
  AND2XL U4294 ( .A(n11547), .B(n11251), .Y(n12922) );
  BUFX12 U4295 ( .A(n12898), .Y(mem_wdata_I[52]) );
  AND2XL U4296 ( .A(n4796), .B(n11282), .Y(n12898) );
  BUFX12 U4297 ( .A(n12881), .Y(mem_wdata_I[69]) );
  AND2XL U4298 ( .A(n4795), .B(n11299), .Y(n12881) );
  BUFX12 U4299 ( .A(n12921), .Y(mem_wdata_I[22]) );
  AND2XL U4300 ( .A(n4794), .B(n11252), .Y(n12921) );
  OA22XL U4301 ( .A0(net112065), .A1(n1456), .B0(net111941), .B1(n3069), .Y(
        n8013) );
  BUFX12 U4302 ( .A(n12897), .Y(mem_wdata_I[53]) );
  AND2XL U4303 ( .A(n4794), .B(n11283), .Y(n12897) );
  BUFX12 U4304 ( .A(n12895), .Y(mem_wdata_I[55]) );
  AND2XL U4305 ( .A(n4796), .B(n11285), .Y(n12895) );
  BUFX12 U4306 ( .A(n12920), .Y(mem_wdata_I[23]) );
  AND2XL U4307 ( .A(n4796), .B(n11253), .Y(n12920) );
  BUFX12 U4308 ( .A(n12878), .Y(mem_wdata_I[72]) );
  AND2XL U4309 ( .A(n4795), .B(n11302), .Y(n12878) );
  BUFX12 U4310 ( .A(n12894), .Y(mem_wdata_I[56]) );
  AND2XL U4311 ( .A(n4794), .B(n11286), .Y(n12894) );
  BUFX12 U4312 ( .A(n12892), .Y(mem_wdata_I[58]) );
  AND2XL U4313 ( .A(n4796), .B(n11288), .Y(n12892) );
  BUFX12 U4314 ( .A(n12919), .Y(mem_wdata_I[24]) );
  AND2XL U4315 ( .A(n4796), .B(n11254), .Y(n12919) );
  BUFX12 U4316 ( .A(n12875), .Y(mem_wdata_I[75]) );
  AND2XL U4317 ( .A(n4795), .B(n11305), .Y(n12875) );
  BUFX12 U4318 ( .A(n12891), .Y(mem_wdata_I[59]) );
  AND2XL U4319 ( .A(n4794), .B(n11289), .Y(n12891) );
  BUFX12 U4320 ( .A(n12889), .Y(mem_wdata_I[61]) );
  AND2XL U4321 ( .A(n4796), .B(n11291), .Y(n12889) );
  BUFX12 U4322 ( .A(n12918), .Y(mem_wdata_I[25]) );
  AND2XL U4323 ( .A(n4794), .B(n11255), .Y(n12918) );
  BUFX12 U4324 ( .A(n12872), .Y(mem_wdata_I[78]) );
  AND2XL U4325 ( .A(n4795), .B(n11308), .Y(n12872) );
  BUFX12 U4326 ( .A(n12888), .Y(mem_wdata_I[62]) );
  AND2XL U4327 ( .A(n4794), .B(n11292), .Y(n12888) );
  BUFX12 U4328 ( .A(n12886), .Y(mem_wdata_I[64]) );
  AND2XL U4329 ( .A(n4796), .B(n11294), .Y(n12886) );
  BUFX12 U4330 ( .A(n12917), .Y(mem_wdata_I[26]) );
  AND2XL U4331 ( .A(n4796), .B(n11256), .Y(n12917) );
  BUFX12 U4332 ( .A(n12869), .Y(mem_wdata_I[81]) );
  AND2XL U4333 ( .A(n4795), .B(n11311), .Y(n12869) );
  BUFX12 U4334 ( .A(n12885), .Y(mem_wdata_I[65]) );
  AND2XL U4335 ( .A(n4794), .B(n11295), .Y(n12885) );
  BUFX12 U4336 ( .A(n12883), .Y(mem_wdata_I[67]) );
  AND2XL U4337 ( .A(n4796), .B(n11297), .Y(n12883) );
  BUFX12 U4338 ( .A(n12916), .Y(mem_wdata_I[27]) );
  AND2XL U4339 ( .A(n4794), .B(n11257), .Y(n12916) );
  BUFX12 U4340 ( .A(n12866), .Y(mem_wdata_I[84]) );
  AND2XL U4341 ( .A(n4795), .B(n11314), .Y(n12866) );
  BUFX12 U4342 ( .A(n12882), .Y(mem_wdata_I[68]) );
  AND2XL U4343 ( .A(n4794), .B(n11298), .Y(n12882) );
  BUFX12 U4344 ( .A(n12880), .Y(mem_wdata_I[70]) );
  AND2XL U4345 ( .A(n4796), .B(n11300), .Y(n12880) );
  BUFX12 U4346 ( .A(n12825), .Y(mem_addr_I[27]) );
  BUFX12 U4347 ( .A(n12915), .Y(mem_wdata_I[28]) );
  AND2XL U4348 ( .A(n4794), .B(n11258), .Y(n12915) );
  BUFX12 U4349 ( .A(n12863), .Y(mem_wdata_I[87]) );
  AND2XL U4350 ( .A(n4795), .B(n11317), .Y(n12863) );
  BUFX12 U4351 ( .A(n12879), .Y(mem_wdata_I[71]) );
  AND2XL U4352 ( .A(n4794), .B(n11301), .Y(n12879) );
  BUFX12 U4353 ( .A(n12877), .Y(mem_wdata_I[73]) );
  AND2XL U4354 ( .A(n4796), .B(n11303), .Y(n12877) );
  BUFX12 U4355 ( .A(n12914), .Y(mem_wdata_I[29]) );
  AND2XL U4356 ( .A(n4796), .B(n11259), .Y(n12914) );
  BUFX12 U4357 ( .A(n12860), .Y(mem_wdata_I[90]) );
  AND2XL U4358 ( .A(n4795), .B(n11320), .Y(n12860) );
  BUFX12 U4359 ( .A(n12876), .Y(mem_wdata_I[74]) );
  AND2XL U4360 ( .A(n4794), .B(n11304), .Y(n12876) );
  BUFX12 U4361 ( .A(n12874), .Y(mem_wdata_I[76]) );
  AND2XL U4362 ( .A(n4796), .B(n11306), .Y(n12874) );
  BUFX12 U4363 ( .A(n12913), .Y(mem_wdata_I[30]) );
  AND2XL U4364 ( .A(n4796), .B(n11260), .Y(n12913) );
  BUFX12 U4365 ( .A(n12857), .Y(mem_wdata_I[93]) );
  AND2XL U4366 ( .A(n4795), .B(n11323), .Y(n12857) );
  BUFX12 U4367 ( .A(n12873), .Y(mem_wdata_I[77]) );
  AND2XL U4368 ( .A(n4794), .B(n11307), .Y(n12873) );
  BUFX12 U4369 ( .A(n12871), .Y(mem_wdata_I[79]) );
  AND2XL U4370 ( .A(n4796), .B(n11309), .Y(n12871) );
  BUFX12 U4371 ( .A(n12912), .Y(mem_wdata_I[31]) );
  AND2XL U4372 ( .A(n4796), .B(n11261), .Y(n12912) );
  BUFX12 U4373 ( .A(n12854), .Y(mem_wdata_I[96]) );
  AND2XL U4374 ( .A(n4795), .B(n11326), .Y(n12854) );
  BUFX12 U4375 ( .A(n12870), .Y(mem_wdata_I[80]) );
  AND2XL U4376 ( .A(n4794), .B(n11310), .Y(n12870) );
  BUFX12 U4377 ( .A(n12868), .Y(mem_wdata_I[82]) );
  AND2XL U4378 ( .A(n4796), .B(n11312), .Y(n12868) );
  BUFX12 U4379 ( .A(n12911), .Y(mem_wdata_I[32]) );
  AND2XL U4380 ( .A(n4794), .B(n11262), .Y(n12911) );
  BUFX12 U4381 ( .A(n12851), .Y(mem_wdata_I[99]) );
  AND2XL U4382 ( .A(n4795), .B(n11329), .Y(n12851) );
  BUFX12 U4383 ( .A(n12867), .Y(mem_wdata_I[83]) );
  AND2XL U4384 ( .A(n4794), .B(n11313), .Y(n12867) );
  BUFX12 U4385 ( .A(n12910), .Y(mem_wdata_I[33]) );
  AND2XL U4386 ( .A(n4796), .B(n11263), .Y(n12910) );
  BUFX12 U4387 ( .A(n12865), .Y(mem_wdata_I[85]) );
  AND2XL U4388 ( .A(n4796), .B(n11315), .Y(n12865) );
  INVXL U4389 ( .A(net106271), .Y(n3961) );
  BUFX12 U4390 ( .A(n12849), .Y(mem_wdata_I[102]) );
  AND2XL U4391 ( .A(n4795), .B(n11332), .Y(n12849) );
  BUFX12 U4392 ( .A(n12864), .Y(mem_wdata_I[86]) );
  AND2XL U4393 ( .A(n4794), .B(n11316), .Y(n12864) );
  XNOR2X4 U4394 ( .A(n11373), .B(ICACHE_addr[14]), .Y(n3964) );
  BUFX12 U4395 ( .A(n12909), .Y(mem_wdata_I[34]) );
  AND2XL U4396 ( .A(n11547), .B(n11264), .Y(n12909) );
  BUFX12 U4397 ( .A(n12862), .Y(mem_wdata_I[88]) );
  AND2XL U4398 ( .A(n4796), .B(n11318), .Y(n12862) );
  BUFX12 U4399 ( .A(n12846), .Y(mem_wdata_I[105]) );
  AND2XL U4400 ( .A(n4795), .B(n11335), .Y(n12846) );
  BUFX12 U4401 ( .A(n12861), .Y(mem_wdata_I[89]) );
  AND2XL U4402 ( .A(n4794), .B(n11319), .Y(n12861) );
  BUFX12 U4403 ( .A(n12908), .Y(mem_wdata_I[35]) );
  AND2XL U4404 ( .A(n4796), .B(n11265), .Y(n12908) );
  BUFX12 U4405 ( .A(n12859), .Y(mem_wdata_I[91]) );
  AND2XL U4406 ( .A(n4796), .B(n11321), .Y(n12859) );
  BUFX12 U4407 ( .A(n12843), .Y(mem_wdata_I[108]) );
  AND2XL U4408 ( .A(n4795), .B(n11338), .Y(n12843) );
  BUFX12 U4409 ( .A(n12858), .Y(mem_wdata_I[92]) );
  AND2XL U4410 ( .A(n4794), .B(n11322), .Y(n12858) );
  BUFX12 U4411 ( .A(n12907), .Y(mem_wdata_I[37]) );
  AND2XL U4412 ( .A(n4794), .B(n11267), .Y(n12907) );
  BUFX12 U4413 ( .A(n12856), .Y(mem_wdata_I[94]) );
  AND2XL U4414 ( .A(n4796), .B(n11324), .Y(n12856) );
  NAND4X8 U4415 ( .A(n5972), .B(n5971), .C(n5970), .D(n5969), .Y(n11384) );
  BUFX12 U4416 ( .A(n12841), .Y(mem_wdata_I[111]) );
  AND2XL U4417 ( .A(n4795), .B(n11341), .Y(n12841) );
  BUFX12 U4418 ( .A(n12906), .Y(mem_wdata_I[39]) );
  AND2XL U4419 ( .A(n4794), .B(n11269), .Y(n12906) );
  BUFX12 U4420 ( .A(n12855), .Y(mem_wdata_I[95]) );
  AND2XL U4421 ( .A(n4794), .B(n11325), .Y(n12855) );
  BUFX12 U4422 ( .A(n12853), .Y(mem_wdata_I[97]) );
  AND2XL U4423 ( .A(n4796), .B(n11327), .Y(n12853) );
  BUFX12 U4424 ( .A(n12839), .Y(mem_wdata_I[114]) );
  AND2XL U4425 ( .A(n4795), .B(n11344), .Y(n12839) );
  BUFX12 U4426 ( .A(n12905), .Y(mem_wdata_I[41]) );
  AND2XL U4427 ( .A(n4796), .B(n11271), .Y(n12905) );
  BUFX12 U4428 ( .A(n12852), .Y(mem_wdata_I[98]) );
  AND2XL U4429 ( .A(n4794), .B(n11328), .Y(n12852) );
  BUFX12 U4430 ( .A(n12850), .Y(mem_wdata_I[100]) );
  AND2XL U4431 ( .A(n4796), .B(n11330), .Y(n12850) );
  BUFX12 U4432 ( .A(n12904), .Y(mem_wdata_I[43]) );
  AND2XL U4433 ( .A(n4796), .B(n11273), .Y(n12904) );
  BUFX12 U4434 ( .A(n12838), .Y(mem_wdata_I[117]) );
  AND2XL U4435 ( .A(n4795), .B(n11347), .Y(n12838) );
  BUFX12 U4436 ( .A(n12847), .Y(mem_wdata_I[104]) );
  AND2XL U4437 ( .A(n4794), .B(n11334), .Y(n12847) );
  BUFX12 U4438 ( .A(n12848), .Y(mem_wdata_I[103]) );
  AND2XL U4439 ( .A(n4796), .B(n11333), .Y(n12848) );
  MX2XL U4440 ( .A(DCACHE_addr[18]), .B(net99639), .S0(n5509), .Y(
        \i_MIPS/n449 ) );
  MX2XL U4441 ( .A(DCACHE_addr[7]), .B(n3961), .S0(n5510), .Y(\i_MIPS/n460 )
         );
  NAND4X2 U4442 ( .A(n10496), .B(n10495), .C(n10497), .D(n10494), .Y(n10504)
         );
  OA22X4 U4443 ( .A0(net112245), .A1(n2389), .B0(net112163), .B1(n884), .Y(
        n7064) );
  OA22X4 U4444 ( .A0(net112245), .A1(n2393), .B0(net112163), .B1(n888), .Y(
        n7052) );
  OA22X4 U4445 ( .A0(net112245), .A1(n2395), .B0(net112161), .B1(n890), .Y(
        n7056) );
  OA22X4 U4446 ( .A0(net112245), .A1(n2398), .B0(net112163), .B1(n893), .Y(
        n6973) );
  NOR2BX4 U4447 ( .AN(\i_MIPS/IR_ID[18] ), .B(\i_MIPS/n318 ), .Y(n4652) );
  NAND2X4 U4448 ( .A(n4660), .B(n4652), .Y(n4480) );
  BUFX12 U4449 ( .A(n4975), .Y(n4971) );
  AO22X4 U4450 ( .A0(net113039), .A1(n10407), .B0(net102300), .B1(n8384), .Y(
        net103630) );
  MX2X1 U4451 ( .A(n8383), .B(n8382), .S0(n5587), .Y(n8384) );
  OA22X2 U4452 ( .A0(n5162), .A1(n456), .B0(n5119), .B1(n3241), .Y(n5990) );
  BUFX6 U4453 ( .A(n5187), .Y(n5162) );
  OAI221X4 U4454 ( .A0(n7867), .A1(n8088), .B0(n7285), .B1(n7693), .C0(n6362), 
        .Y(n6674) );
  OAI32X2 U4455 ( .A0(\i_MIPS/ID_EX[56] ), .A1(\i_MIPS/ID_EX[55] ), .A2(n6947), 
        .B0(n6620), .B1(\i_MIPS/n356 ), .Y(n6623) );
  NAND4X2 U4456 ( .A(n6204), .B(n6203), .C(n6298), .D(n6202), .Y(net101981) );
  INVX8 U4457 ( .A(net99538), .Y(net103060) );
  AOI211X2 U4458 ( .A0(n8822), .A1(n6436), .B0(n6435), .C0(n6434), .Y(n6437)
         );
  BUFX4 U4459 ( .A(n5405), .Y(n5379) );
  NAND3BX4 U4460 ( .AN(net113540), .B(net108204), .C(n3671), .Y(net100084) );
  NAND3BX4 U4461 ( .AN(n3672), .B(n3752), .C(net108204), .Y(net100105) );
  AOI222X1 U4462 ( .A0(net109791), .A1(net98185), .B0(mem_rdata_D[6]), .B1(
        n117), .C0(n12991), .C1(net109801), .Y(net100025) );
  NAND4X2 U4463 ( .A(net105032), .B(net105033), .C(net105034), .D(net105035), 
        .Y(net98185) );
  AO21X4 U4464 ( .A0(net100019), .A1(net100020), .B0(net113077), .Y(net100013)
         );
  OAI211X4 U4465 ( .A0(net105006), .A1(n4077), .B0(net113439), .C0(net112607), 
        .Y(net100020) );
  OA22X2 U4466 ( .A0(n11089), .A1(net140281), .B0(net98430), .B1(n11088), .Y(
        n11091) );
  MX2XL U4467 ( .A(n10461), .B(n3584), .S0(n5509), .Y(\i_MIPS/n383 ) );
  AOI32X2 U4468 ( .A0(n8149), .A1(\i_MIPS/ID_EX[83] ), .A2(n8148), .B0(n6429), 
        .B1(n6428), .Y(n6438) );
  NAND3BX2 U4469 ( .AN(n9259), .B(n4798), .C(n8805), .Y(n6428) );
  CLKINVX20 U4470 ( .A(n4723), .Y(n5595) );
  AOI21X2 U4471 ( .A0(n7356), .A1(n3801), .B0(n7273), .Y(n4551) );
  OA22X4 U4472 ( .A0(n5164), .A1(n1951), .B0(n5119), .B1(n375), .Y(n6031) );
  AOI211X2 U4473 ( .A0(n8263), .A1(n8098), .B0(n8097), .C0(n8096), .Y(n8099)
         );
  BUFX12 U4474 ( .A(n12903), .Y(mem_wdata_I[44]) );
  AND2XL U4475 ( .A(n4794), .B(n11274), .Y(n12903) );
  BUFX12 U4476 ( .A(n12844), .Y(mem_wdata_I[107]) );
  AND2XL U4477 ( .A(n4794), .B(n11337), .Y(n12844) );
  BUFX12 U4478 ( .A(n12845), .Y(mem_wdata_I[106]) );
  AND2XL U4479 ( .A(n4796), .B(n11336), .Y(n12845) );
  BUFX12 U4480 ( .A(n12902), .Y(mem_wdata_I[45]) );
  AND2XL U4481 ( .A(n4796), .B(n11275), .Y(n12902) );
  BUFX12 U4482 ( .A(n12842), .Y(mem_wdata_I[110]) );
  AND2XL U4483 ( .A(n4794), .B(n11340), .Y(n12842) );
  BUFX12 U4484 ( .A(n12901), .Y(mem_wdata_I[46]) );
  AND2XL U4485 ( .A(n4794), .B(n11276), .Y(n12901) );
  BUFX12 U4486 ( .A(n12840), .Y(mem_wdata_I[113]) );
  AND2XL U4487 ( .A(n4794), .B(n11343), .Y(n12840) );
  BUFX12 U4488 ( .A(n12900), .Y(mem_wdata_I[47]) );
  AND2XL U4489 ( .A(n4794), .B(n11277), .Y(n12900) );
  AOI2BB1X4 U4490 ( .A0N(n7708), .A1N(n6572), .B0(n8146), .Y(n6576) );
  NAND2X4 U4491 ( .A(n3643), .B(\i_MIPS/n359 ), .Y(n6602) );
  OAI221X2 U4492 ( .A0(\i_MIPS/n360 ), .A1(n4825), .B0(\i_MIPS/n359 ), .B1(
        n4817), .C0(n6948), .Y(n7872) );
  OAI2BB1X4 U4493 ( .A0N(n6348), .A1N(n6633), .B0(n6638), .Y(n6349) );
  NAND3BX2 U4494 ( .AN(ICACHE_addr[1]), .B(\i_MIPS/PC/n4 ), .C(n9572), .Y(
        n9575) );
  INVXL U4495 ( .A(n8995), .Y(n3995) );
  OAI221X4 U4496 ( .A0(\i_MIPS/Register/register[18][26] ), .A1(n4923), .B0(
        \i_MIPS/Register/register[26][26] ), .B1(n4917), .C0(n8377), .Y(n8380)
         );
  BUFX16 U4497 ( .A(n4919), .Y(n4923) );
  NAND2BX4 U4498 ( .AN(n4348), .B(n11339), .Y(n3998) );
  OR2X2 U4499 ( .A(n4348), .B(n4000), .Y(n3999) );
  OAI21X4 U4500 ( .A0(n4714), .A1(n6207), .B0(n3530), .Y(n4496) );
  NAND2BX2 U4501 ( .AN(n4348), .B(n11353), .Y(n4001) );
  CLKAND2X12 U4502 ( .A(\i_MIPS/IR_ID[17] ), .B(\i_MIPS/n312 ), .Y(n4660) );
  BUFX16 U4503 ( .A(n4931), .Y(n4932) );
  AO22X4 U4504 ( .A0(n5000), .A1(n347), .B0(n4996), .B1(n1929), .Y(n7940) );
  AO22X4 U4505 ( .A0(n5000), .A1(n333), .B0(n4996), .B1(n1910), .Y(n7931) );
  AO22X4 U4506 ( .A0(n5000), .A1(n334), .B0(n4996), .B1(n1911), .Y(n8037) );
  AO22X4 U4507 ( .A0(n5000), .A1(n335), .B0(n4996), .B1(n1912), .Y(n8028) );
  AO22X4 U4508 ( .A0(n5000), .A1(n348), .B0(n4996), .B1(n1930), .Y(n7683) );
  OA22X2 U4509 ( .A0(n5162), .A1(n457), .B0(n5119), .B1(n2011), .Y(n5998) );
  INVXL U4510 ( .A(net103060), .Y(n4002) );
  NAND2BX4 U4511 ( .AN(n5453), .B(n11328), .Y(n9606) );
  MX2XL U4512 ( .A(DCACHE_addr[25]), .B(n4002), .S0(n5508), .Y(\i_MIPS/n442 )
         );
  MX2XL U4513 ( .A(DCACHE_addr[4]), .B(net98472), .S0(n5507), .Y(\i_MIPS/n463 ) );
  NAND4X4 U4514 ( .A(n8295), .B(n8294), .C(n8293), .D(n8292), .Y(n11412) );
  AO22X4 U4515 ( .A0(n4991), .A1(n350), .B0(n4984), .B1(n1932), .Y(n6185) );
  NAND2X4 U4516 ( .A(\i_MIPS/ALUin1[4] ), .B(n3720), .Y(n7359) );
  OA22X4 U4517 ( .A0(n5164), .A1(n1952), .B0(n5120), .B1(n376), .Y(n6027) );
  NAND4X2 U4518 ( .A(n8964), .B(n8963), .C(n8962), .D(n8961), .Y(n11413) );
  OA22X4 U4519 ( .A0(net112063), .A1(n2400), .B0(net111939), .B1(n895), .Y(
        n7912) );
  BUFX12 U4520 ( .A(net111957), .Y(net111939) );
  OAI211X2 U4521 ( .A0(n7824), .A1(n7823), .B0(net113439), .C0(net112609), .Y(
        n10184) );
  OAI32X2 U4522 ( .A0(\i_MIPS/ID_EX[88] ), .A1(\i_MIPS/ID_EX[87] ), .A2(n6947), 
        .B0(n6621), .B1(\i_MIPS/n356 ), .Y(n6622) );
  AOI222X2 U4523 ( .A0(n5475), .A1(n11483), .B0(mem_rdata_D[96]), .B1(n116), 
        .C0(n12997), .C1(n5473), .Y(n10852) );
  NAND4X2 U4524 ( .A(n6542), .B(n6541), .C(n6540), .D(n6539), .Y(n11483) );
  AO21X4 U4525 ( .A0(net98967), .A1(net98968), .B0(net113079), .Y(net98964) );
  AO21X4 U4526 ( .A0(net98967), .A1(net98968), .B0(net112727), .Y(net98899) );
  OAI211X4 U4527 ( .A0(n6544), .A1(n6543), .B0(net113437), .C0(n3709), .Y(
        net98968) );
  OR2X2 U4528 ( .A(net112229), .B(n2024), .Y(n4221) );
  NAND2BX2 U4529 ( .AN(n4348), .B(n11342), .Y(n4008) );
  OA22X4 U4530 ( .A0(n5250), .A1(n1953), .B0(n5228), .B1(n377), .Y(n6030) );
  NAND2BX2 U4531 ( .AN(n4334), .B(n11349), .Y(n4009) );
  CLKINVX20 U4532 ( .A(n4009), .Y(mem_wdata_I[119]) );
  AOI222XL U4533 ( .A0(n5487), .A1(n11427), .B0(mem_rdata_D[39]), .B1(n117), 
        .C0(n12990), .C1(n5483), .Y(n10748) );
  NAND4X2 U4534 ( .A(n7487), .B(n7486), .C(n7485), .D(n7484), .Y(n11427) );
  AO22X4 U4535 ( .A0(net113445), .A1(n11474), .B0(net102346), .B1(n11505), .Y(
        n8304) );
  AOI222X1 U4536 ( .A0(n5475), .A1(n11505), .B0(mem_rdata_D[119]), .B1(n116), 
        .C0(n12974), .C1(n5473), .Y(n10557) );
  NAND2BX2 U4537 ( .AN(n4323), .B(n11345), .Y(n4013) );
  CLKINVX20 U4538 ( .A(n4013), .Y(mem_wdata_I[115]) );
  NAND4X2 U4539 ( .A(n7499), .B(n7498), .C(n7497), .D(n7496), .Y(n11489) );
  NAND2BX2 U4540 ( .AN(n4323), .B(n11352), .Y(n4014) );
  CLKINVX20 U4541 ( .A(n4014), .Y(mem_wdata_I[122]) );
  AOI222X1 U4542 ( .A0(net109791), .A1(n11404), .B0(mem_rdata_D[15]), .B1(n117), .C0(n12982), .C1(net109801), .Y(n10193) );
  OAI211X4 U4543 ( .A0(n7068), .A1(n7067), .B0(net113437), .C0(n3709), .Y(
        net99978) );
  AO22X4 U4544 ( .A0(n4972), .A1(n230), .B0(n4967), .B1(n1916), .Y(n7424) );
  AO22X4 U4545 ( .A0(n4972), .A1(n339), .B0(n4967), .B1(n1917), .Y(n7415) );
  AO22X4 U4546 ( .A0(n4972), .A1(n187), .B0(n4967), .B1(n1919), .Y(n7262) );
  AO22X4 U4547 ( .A0(n4972), .A1(n288), .B0(n4965), .B1(n1920), .Y(n7253) );
  BUFX12 U4548 ( .A(n4975), .Y(n4972) );
  NAND4X2 U4549 ( .A(n9248), .B(n9247), .C(n9246), .D(n9245), .Y(n11419) );
  INVX2 U4550 ( .A(n11419), .Y(n10689) );
  INVX3 U4551 ( .A(n8437), .Y(n8916) );
  NAND4X2 U4552 ( .A(n9090), .B(n9089), .C(n9088), .D(n9087), .Y(n11420) );
  NAND3BX4 U4553 ( .AN(n7027), .B(n7026), .C(n4928), .Y(n7049) );
  NOR4X4 U4554 ( .A(n6811), .B(n6810), .C(n6809), .D(n6808), .Y(n6822) );
  AO22XL U4555 ( .A0(n4895), .A1(n473), .B0(n4891), .B1(n2039), .Y(n6809) );
  OR2X8 U4556 ( .A(n11018), .B(net110247), .Y(n4422) );
  CLKMX2X4 U4557 ( .A(n7353), .B(n6431), .S0(n5590), .Y(n6779) );
  NAND4X4 U4558 ( .A(n7636), .B(n7635), .C(n7634), .D(n7633), .Y(n11422) );
  XOR2X4 U4559 ( .A(n11364), .B(\i_MIPS/PC/n9 ), .Y(n4018) );
  AOI2BB1X2 U4560 ( .A0N(n8737), .A1N(n3591), .B0(n8735), .Y(n8738) );
  NAND2BX2 U4561 ( .AN(n4334), .B(n11348), .Y(n4019) );
  CLKINVX20 U4562 ( .A(n4019), .Y(mem_wdata_I[118]) );
  OAI221X2 U4563 ( .A0(\i_MIPS/n370 ), .A1(n4826), .B0(\i_MIPS/n369 ), .B1(
        n4818), .C0(n6257), .Y(n6776) );
  XOR2XL U4564 ( .A(n9607), .B(n4005), .Y(n11195) );
  NAND4X2 U4565 ( .A(n8850), .B(n8849), .C(n8848), .D(n8847), .Y(n11423) );
  AO22X4 U4566 ( .A0(net113447), .A1(n11455), .B0(net102346), .B1(n11486), .Y(
        n8778) );
  NAND4X4 U4567 ( .A(n8777), .B(n8776), .C(n8775), .D(n8774), .Y(n11486) );
  NAND2BX2 U4568 ( .AN(n4348), .B(n11351), .Y(n4022) );
  AOI222X2 U4569 ( .A0(n5475), .A1(n11499), .B0(mem_rdata_D[113]), .B1(n116), 
        .C0(n12980), .C1(n5473), .Y(n10596) );
  AO21X4 U4570 ( .A0(net99311), .A1(net99312), .B0(net113077), .Y(net99293) );
  AO21X4 U4571 ( .A0(net99311), .A1(net99312), .B0(net112729), .Y(net104706)
         );
  OAI211X4 U4572 ( .A0(n7735), .A1(n7734), .B0(net113439), .C0(net112609), .Y(
        net99312) );
  NAND4X4 U4573 ( .A(n8094), .B(n8091), .C(n8092), .D(n8093), .Y(n8097) );
  OAI222X4 U4574 ( .A0(n8814), .A1(n8816), .B0(n7561), .B1(n7963), .C0(n8726), 
        .C1(n7969), .Y(n7564) );
  NAND2X2 U4575 ( .A(n7558), .B(n4707), .Y(n7963) );
  AOI211X2 U4576 ( .A0(n7565), .A1(n8822), .B0(n7564), .C0(n7563), .Y(n7566)
         );
  OAI221X2 U4577 ( .A0(net106270), .A1(net112709), .B0(net106271), .B1(
        net112723), .C0(net106272), .Y(net99056) );
  OAI222X4 U4578 ( .A0(n8659), .A1(n8346), .B0(n8345), .B1(n8437), .C0(n8360), 
        .C1(n8805), .Y(n8357) );
  OAI211X2 U4579 ( .A0(n7158), .A1(n7157), .B0(net113437), .C0(n3709), .Y(
        net99038) );
  CLKBUFX2 U4580 ( .A(net112095), .Y(net112043) );
  BUFX16 U4581 ( .A(net112095), .Y(net112037) );
  INVX4 U4582 ( .A(n6201), .Y(n6298) );
  OA22X1 U4583 ( .A0(net112071), .A1(n1239), .B0(net111947), .B1(n2844), .Y(
        n8397) );
  OA21X4 U4584 ( .A0(\i_MIPS/n362 ), .A1(n4819), .B0(n7280), .Y(n7037) );
  OA22X2 U4585 ( .A0(n5248), .A1(n1611), .B0(n5203), .B1(n3242), .Y(n5989) );
  NAND4X2 U4586 ( .A(n6971), .B(n6970), .C(n6969), .D(n6968), .Y(n11465) );
  OA22XL U4587 ( .A0(net112461), .A1(n1457), .B0(net112337), .B1(n3070), .Y(
        n6970) );
  AOI222X2 U4588 ( .A0(n8812), .A1(n3636), .B0(n8811), .B1(n8810), .C0(n8809), 
        .C1(n8808), .Y(n8813) );
  XOR2X4 U4589 ( .A(n3565), .B(\i_MIPS/PC/n33 ), .Y(n4024) );
  OAI33X2 U4590 ( .A0(n8078), .A1(n8076), .A2(n3600), .B0(n3699), .B1(n8076), 
        .B2(n9262), .Y(n8101) );
  AOI2BB2X2 U4591 ( .B0(\i_MIPS/IF_ID[84] ), .B1(n148), .A0N(net110191), .A1N(
        \i_MIPS/n199 ), .Y(n11153) );
  AO22X4 U4592 ( .A0(n115), .A1(ICACHE_addr[18]), .B0(n5463), .B1(n11377), .Y(
        n10997) );
  OR2X1 U4593 ( .A(n4559), .B(net110243), .Y(n4213) );
  OR2X1 U4594 ( .A(n4532), .B(net110243), .Y(n4416) );
  XOR3X2 U4595 ( .A(n10897), .B(n10896), .C(n10895), .Y(n10899) );
  XOR2X4 U4596 ( .A(n2), .B(n4560), .Y(n4121) );
  AOI222X1 U4597 ( .A0(net109791), .A1(n11399), .B0(mem_rdata_D[10]), .B1(n116), .C0(n12987), .C1(net109801), .Y(n10590) );
  MXI2X4 U4598 ( .A(n8088), .B(n7283), .S0(n5589), .Y(n4519) );
  OAI222X4 U4599 ( .A0(n9284), .A1(n6674), .B0(n8087), .B1(n9286), .C0(n8659), 
        .C1(n9170), .Y(n6679) );
  NAND2X4 U4600 ( .A(n9143), .B(\i_MIPS/n340 ), .Y(n11220) );
  INVX2 U4601 ( .A(n9142), .Y(n9143) );
  AO22X4 U4602 ( .A0(net99407), .A1(net113039), .B0(net102300), .B1(n8008), 
        .Y(net104271) );
  AOI2BB1X2 U4603 ( .A0N(n9007), .A1N(n7695), .B0(n8089), .Y(n7702) );
  BUFX6 U4604 ( .A(n4620), .Y(n4871) );
  AO22X4 U4605 ( .A0(net113447), .A1(n11463), .B0(net102346), .B1(n11494), .Y(
        n6285) );
  AOI222X1 U4606 ( .A0(n5481), .A1(n11463), .B0(mem_rdata_D[76]), .B1(n117), 
        .C0(n12985), .C1(n5478), .Y(n10793) );
  NAND4X2 U4607 ( .A(n6280), .B(n6279), .C(n6278), .D(n6277), .Y(n11463) );
  OAI221X2 U4608 ( .A0(net103707), .A1(net112707), .B0(net103708), .B1(
        net112721), .C0(net103709), .Y(n4025) );
  OAI221XL U4609 ( .A0(net103707), .A1(net112707), .B0(net103708), .B1(
        net112721), .C0(net103709), .Y(net99378) );
  AOI222X1 U4610 ( .A0(net109791), .A1(n11417), .B0(mem_rdata_D[28]), .B1(n117), .C0(n12969), .C1(net109801), .Y(n10402) );
  OAI221X1 U4611 ( .A0(\i_MIPS/Register/register[2][18] ), .A1(n4946), .B0(
        \i_MIPS/Register/register[10][18] ), .B1(n4484), .C0(n7930), .Y(n7938)
         );
  AO22X4 U4612 ( .A0(n4990), .A1(n340), .B0(n4981), .B1(n1921), .Y(n7422) );
  AO22X4 U4613 ( .A0(n9312), .A1(n343), .B0(n4981), .B1(n1924), .Y(n7260) );
  AO22X4 U4614 ( .A0(n4989), .A1(n344), .B0(n4981), .B1(n1925), .Y(n7251) );
  XOR2X4 U4615 ( .A(n3732), .B(n4533), .Y(n4102) );
  NAND4X2 U4616 ( .A(n6384), .B(n6383), .C(n6382), .D(n6381), .Y(n11402) );
  AND4X8 U4617 ( .A(n6129), .B(n6128), .C(n6127), .D(n6130), .Y(n4026) );
  INVX12 U4618 ( .A(net98881), .Y(net101969) );
  NAND4X4 U4619 ( .A(n7495), .B(n7494), .C(n7493), .D(n7492), .Y(n11458) );
  OA22X1 U4620 ( .A0(net112679), .A1(n1240), .B0(net112573), .B1(n2845), .Y(
        n7495) );
  OR2X6 U4621 ( .A(\i_MIPS/n345 ), .B(n4810), .Y(n4196) );
  OAI222X2 U4622 ( .A0(\i_MIPS/PC/n28 ), .A1(net110215), .B0(n4531), .B1(
        net110241), .C0(n3602), .C1(n10355), .Y(n10360) );
  OA22X4 U4623 ( .A0(net112511), .A1(n1954), .B0(net112379), .B1(n378), .Y(
        n6051) );
  OR2X2 U4624 ( .A(net100082), .B(n2025), .Y(n4219) );
  OAI2BB1X4 U4625 ( .A0N(n10207), .A1N(n10212), .B0(n10206), .Y(n10208) );
  OAI211X4 U4626 ( .A0(n7287), .A1(n3529), .B0(n7550), .C0(n7459), .Y(n4028)
         );
  MX2X1 U4627 ( .A(n9324), .B(n9323), .S0(net108959), .Y(n9326) );
  NAND2X6 U4628 ( .A(n3303), .B(n1609), .Y(n6118) );
  OAI221X2 U4629 ( .A0(n6628), .A1(n6494), .B0(n6493), .B1(n6492), .C0(n8891), 
        .Y(n6495) );
  XOR2X4 U4630 ( .A(n10697), .B(ICACHE_addr[27]), .Y(n10698) );
  NAND3BX1 U4631 ( .AN(n8154), .B(n8147), .C(n9258), .Y(n8166) );
  NAND3BX4 U4632 ( .AN(n9552), .B(n4661), .C(n4640), .Y(n5984) );
  INVX2 U4633 ( .A(n8804), .Y(n8807) );
  CLKAND2X12 U4634 ( .A(net113607), .B(n11440), .Y(mem_wdata_D[52]) );
  AOI222X1 U4635 ( .A0(n5487), .A1(n11440), .B0(mem_rdata_D[52]), .B1(n117), 
        .C0(n12977), .C1(n5483), .Y(n10530) );
  NAND3BX1 U4636 ( .AN(n8077), .B(n4928), .C(n3699), .Y(n8100) );
  NAND2BX4 U4637 ( .AN(n5453), .B(n11330), .Y(n9619) );
  NAND2BX4 U4638 ( .AN(n6224), .B(n7181), .Y(n6599) );
  XOR2X4 U4639 ( .A(n3199), .B(n6086), .Y(n6098) );
  NAND2X2 U4640 ( .A(n7198), .B(n4707), .Y(n8345) );
  INVXL U4641 ( .A(n3314), .Y(n4030) );
  AOI222X1 U4642 ( .A0(n5486), .A1(n11425), .B0(mem_rdata_D[36]), .B1(n117), 
        .C0(n12993), .C1(n5482), .Y(n10163) );
  CLKINVX1 U4643 ( .A(n11425), .Y(n10162) );
  NAND4X2 U4644 ( .A(n7396), .B(n7395), .C(n7394), .D(n7393), .Y(n11425) );
  AND2XL U4645 ( .A(net100048), .B(net100049), .Y(n4545) );
  AOI32X2 U4646 ( .A0(n8163), .A1(n8162), .A2(n9258), .B0(n8161), .B1(n8160), 
        .Y(n8164) );
  CLKINVX1 U4647 ( .A(n11421), .Y(n10860) );
  NAND4X2 U4648 ( .A(n6530), .B(n6529), .C(n6528), .D(n6527), .Y(n11421) );
  NAND3BX4 U4649 ( .AN(n8556), .B(n8555), .C(n4924), .Y(n8557) );
  OA22X2 U4650 ( .A0(n11152), .A1(net140280), .B0(net98430), .B1(n11151), .Y(
        n11154) );
  AO22X1 U4651 ( .A0(n5001), .A1(n648), .B0(n4997), .B1(n2169), .Y(n8601) );
  AO22X1 U4652 ( .A0(n4979), .A1(n553), .B0(n4976), .B1(n2056), .Y(n8603) );
  OA22X4 U4653 ( .A0(net112499), .A1(n2401), .B0(net112325), .B1(n379), .Y(
        n6149) );
  OAI2BB2X1 U4654 ( .B0(\i_MIPS/n171 ), .B1(net110225), .A0N(n173), .A1N(n3847), .Y(\i_MIPS/N112 ) );
  OAI211X2 U4655 ( .A0(n7869), .A1(n7791), .B0(n7790), .C0(n7789), .Y(n8725)
         );
  NAND4BX4 U4656 ( .AN(n7632), .B(n7631), .C(n7630), .D(n7629), .Y(net98929)
         );
  CLKINVX8 U4657 ( .A(n10382), .Y(n10499) );
  NAND4X4 U4658 ( .A(n6871), .B(n6870), .C(n6869), .D(n6868), .Y(n11429) );
  OA22X2 U4659 ( .A0(net112235), .A1(n921), .B0(net112165), .B1(n2458), .Y(
        n6869) );
  NAND4X2 U4660 ( .A(n6717), .B(n6716), .C(n6715), .D(n6714), .Y(n11480) );
  OA22XL U4661 ( .A0(net112233), .A1(n1458), .B0(net112165), .B1(n3071), .Y(
        n6715) );
  NAND2BX4 U4662 ( .AN(n6597), .B(n9168), .Y(n8643) );
  CLKAND2X12 U4663 ( .A(net113607), .B(n11479), .Y(mem_wdata_D[92]) );
  AOI222X1 U4664 ( .A0(n5479), .A1(n11479), .B0(mem_rdata_D[92]), .B1(n117), 
        .C0(n12969), .C1(n5476), .Y(n10399) );
  NAND4X2 U4665 ( .A(n6792), .B(n6791), .C(n6790), .D(n6789), .Y(n11397) );
  NAND3BX4 U4666 ( .AN(n4521), .B(n10216), .C(n11074), .Y(n10217) );
  OA22X4 U4667 ( .A0(net112453), .A1(n2402), .B0(net112329), .B1(n896), .Y(
        n6160) );
  BUFX16 U4668 ( .A(n4919), .Y(n4920) );
  OAI221X1 U4669 ( .A0(\i_MIPS/Register/register[18][13] ), .A1(n4920), .B0(
        \i_MIPS/Register/register[26][13] ), .B1(n4915), .C0(n6408), .Y(n6411)
         );
  OAI221X1 U4670 ( .A0(\i_MIPS/Register/register[2][13] ), .A1(n4920), .B0(
        \i_MIPS/Register/register[10][13] ), .B1(n4915), .C0(n6399), .Y(n6402)
         );
  NAND2X2 U4671 ( .A(n6234), .B(\i_MIPS/ALUin1[1] ), .Y(n8714) );
  OA22X1 U4672 ( .A0(net112681), .A1(n1241), .B0(net112565), .B1(n2846), .Y(
        n6392) );
  NAND4X2 U4673 ( .A(n6276), .B(n6275), .C(n6274), .D(n6273), .Y(n11401) );
  AO21X4 U4674 ( .A0(net99014), .A1(net99015), .B0(net112727), .Y(net107238)
         );
  NAND3BX4 U4675 ( .AN(n6604), .B(n6603), .C(n6602), .Y(n6610) );
  AOI2BB1X4 U4676 ( .A0N(n3704), .A1N(n3773), .B0(n6601), .Y(n6604) );
  NAND2X1 U4677 ( .A(net99737), .B(net113551), .Y(n10349) );
  INVX6 U4678 ( .A(n4887), .Y(n4882) );
  OA22X2 U4679 ( .A0(net112245), .A1(n2419), .B0(net112161), .B1(n465), .Y(
        n7146) );
  NAND4BX4 U4680 ( .AN(n10253), .B(n10254), .C(net110213), .D(net99855), .Y(
        n10252) );
  AOI2BB1X4 U4681 ( .A0N(n4798), .A1N(n8649), .B0(n4800), .Y(n8650) );
  CLKAND2X12 U4682 ( .A(net113606), .B(n11449), .Y(mem_wdata_D[61]) );
  AOI222X1 U4683 ( .A0(n5486), .A1(n11449), .B0(mem_rdata_D[61]), .B1(n116), 
        .C0(n12968), .C1(n5482), .Y(n10484) );
  CLKINVX1 U4684 ( .A(n11449), .Y(n10483) );
  NAND4X2 U4685 ( .A(n6709), .B(n6708), .C(n6707), .D(n6706), .Y(n11449) );
  NAND2X2 U4686 ( .A(\i_MIPS/ALUin1[27] ), .B(n6565), .Y(n8648) );
  OA22X4 U4687 ( .A0(\i_MIPS/n343 ), .A1(n4811), .B0(\i_MIPS/n344 ), .B1(n4804), .Y(n7020) );
  CLKAND2X12 U4688 ( .A(n4822), .B(\i_MIPS/ALUin1[27] ), .Y(n4668) );
  NAND2X2 U4689 ( .A(n6615), .B(\i_MIPS/n344 ), .Y(n8647) );
  XNOR3X2 U4690 ( .A(n10874), .B(n4586), .C(n10873), .Y(n10876) );
  INVX2 U4691 ( .A(n10873), .Y(n10878) );
  NOR2BX4 U4692 ( .AN(\i_MIPS/IR_ID[23] ), .B(\i_MIPS/n231 ), .Y(n4654) );
  NAND4BX4 U4693 ( .AN(n7764), .B(n7763), .C(n7762), .D(n7761), .Y(n7775) );
  NAND3X2 U4694 ( .A(n9018), .B(n9258), .C(n9015), .Y(n9022) );
  OAI211X2 U4695 ( .A0(n7182), .A1(n3838), .B0(n7180), .C0(n7179), .Y(n7184)
         );
  NAND3BX4 U4696 ( .AN(n10288), .B(n10287), .C(n10286), .Y(\i_MIPS/PC/n48 ) );
  NAND4X4 U4697 ( .A(n7318), .B(n7317), .C(n7316), .D(n7315), .Y(n11426) );
  AOI222X4 U4698 ( .A0(n5479), .A1(n11467), .B0(mem_rdata_D[80]), .B1(n117), 
        .C0(n12981), .C1(n5476), .Y(n10453) );
  NAND4X2 U4699 ( .A(net105044), .B(net105045), .C(net105046), .D(net105047), 
        .Y(net98153) );
  NAND3BX4 U4700 ( .AN(n10904), .B(n10903), .C(n10902), .Y(\i_MIPS/PC/n44 ) );
  NAND4X2 U4701 ( .A(n9086), .B(n9085), .C(n9084), .D(n9083), .Y(n11451) );
  OAI222X1 U4702 ( .A0(n3693), .A1(net110213), .B0(n4529), .B1(net110243), 
        .C0(n11052), .C1(net110247), .Y(n11056) );
  NAND4X2 U4703 ( .A(n8291), .B(n8290), .C(n8289), .D(n8288), .Y(n11443) );
  NAND4X4 U4704 ( .A(n6538), .B(n6537), .C(n6536), .D(n6535), .Y(n11452) );
  INVX20 U4705 ( .A(net130576), .Y(net110189) );
  NAND2BX1 U4706 ( .AN(net113725), .B(n11429), .Y(n4041) );
  XOR2X4 U4707 ( .A(n11369), .B(\i_MIPS/PC/n14 ), .Y(n4042) );
  NAND4X2 U4708 ( .A(n8960), .B(n8959), .C(n8958), .D(n8957), .Y(n11444) );
  NAND4X2 U4709 ( .A(n7242), .B(n7241), .C(n7240), .D(n7239), .Y(n11461) );
  NAND4X4 U4710 ( .A(n7644), .B(n7643), .C(n7642), .D(n7641), .Y(n11453) );
  NAND4X2 U4711 ( .A(n7234), .B(n7233), .C(n7232), .D(n7231), .Y(n11430) );
  OAI221X4 U4712 ( .A0(\i_MIPS/n361 ), .A1(n4825), .B0(\i_MIPS/n360 ), .B1(
        n4818), .C0(n6361), .Y(n8098) );
  AOI222X1 U4713 ( .A0(n5481), .A1(n11482), .B0(mem_rdata_D[95]), .B1(n116), 
        .C0(n5478), .C1(n12966), .Y(n11207) );
  NAND4X2 U4714 ( .A(n9094), .B(n9093), .C(n9092), .D(n9091), .Y(n11482) );
  NAND2X2 U4715 ( .A(n9932), .B(n9931), .Y(n11217) );
  OAI211X4 U4716 ( .A0(n9100), .A1(n9099), .B0(net102344), .C0(n3709), .Y(
        n9931) );
  NAND2BX4 U4717 ( .AN(n5452), .B(n11335), .Y(n9652) );
  AOI222X1 U4718 ( .A0(net109791), .A1(n11403), .B0(mem_rdata_D[14]), .B1(n117), .C0(n12983), .C1(net109801), .Y(n10442) );
  OAI211X4 U4719 ( .A0(n6977), .A1(n6976), .B0(net113437), .C0(net112607), .Y(
        net99582) );
  XOR2X4 U4720 ( .A(n10863), .B(\i_MIPS/n233 ), .Y(n4664) );
  NOR4X8 U4721 ( .A(n6169), .B(n6168), .C(n6167), .D(n6166), .Y(n6170) );
  NAND4X2 U4722 ( .A(n8479), .B(n8478), .C(n8477), .D(n8476), .Y(n11445) );
  NAND4X4 U4723 ( .A(n7152), .B(n7151), .C(n7150), .D(n7149), .Y(n11462) );
  NAND2BX4 U4724 ( .AN(n10213), .B(n10265), .Y(n10215) );
  NAND2X2 U4725 ( .A(n4488), .B(n11389), .Y(n11514) );
  NAND2X2 U4726 ( .A(n4604), .B(n10159), .Y(net98396) );
  NAND4X2 U4727 ( .A(n7144), .B(n7143), .C(n7142), .D(n7141), .Y(n11431) );
  NAND4X2 U4728 ( .A(n9047), .B(n9046), .C(n9045), .D(n9044), .Y(n11448) );
  NAND4X4 U4729 ( .A(n6796), .B(n6795), .C(n6794), .D(n6793), .Y(n11459) );
  NAND4X2 U4730 ( .A(n8396), .B(n8395), .C(n8394), .D(n8393), .Y(n11477) );
  NAND4X2 U4731 ( .A(n8202), .B(n8201), .C(n8200), .D(n8199), .Y(n11467) );
  AO22X1 U4732 ( .A0(ICACHE_addr[15]), .A1(mem_read_I), .B0(n4795), .B1(n11374), .Y(n12835) );
  OAI222X2 U4733 ( .A0(n4525), .A1(net110241), .B0(n10732), .B1(n10736), .C0(
        \i_MIPS/PC/n33 ), .C1(net110213), .Y(n10735) );
  MXI2X1 U4734 ( .A(n10450), .B(n10449), .S0(n5495), .Y(n10451) );
  NAND4X4 U4735 ( .A(n9059), .B(n9058), .C(n9057), .D(n9056), .Y(n11510) );
  AND3X8 U4736 ( .A(n7780), .B(n7800), .C(n4926), .Y(n7797) );
  MXI2X4 U4737 ( .A(\i_MIPS/ID_EX[112] ), .B(\i_MIPS/ID_EX[85] ), .S0(
        \i_MIPS/ID_EX_5 ), .Y(n6293) );
  MX2XL U4738 ( .A(DCACHE_addr[0]), .B(net99087), .S0(n5511), .Y(\i_MIPS/n467 ) );
  NAND2XL U4739 ( .A(n12965), .B(net113087), .Y(n10751) );
  AO21X1 U4740 ( .A0(n10153), .A1(n10152), .B0(n10151), .Y(n10159) );
  AOI222X1 U4741 ( .A0(n5480), .A1(n11475), .B0(mem_rdata_D[88]), .B1(n117), 
        .C0(n12973), .C1(n5477), .Y(n10573) );
  NAND4X2 U4742 ( .A(n8968), .B(n8967), .C(n8966), .D(n8965), .Y(n11475) );
  INVXL U4743 ( .A(net104525), .Y(n4066) );
  AOI2BB1X4 U4744 ( .A0N(n11106), .A1N(n11105), .B0(n11104), .Y(n11108) );
  INVX4 U4745 ( .A(n4724), .Y(n11106) );
  NAND3BX4 U4746 ( .AN(n6224), .B(n4522), .C(n6768), .Y(n6605) );
  OAI211X2 U4747 ( .A0(n3892), .A1(n6769), .B0(n4028), .C0(n4522), .Y(n7090)
         );
  NOR2BX4 U4748 ( .AN(\i_MIPS/IR_ID[16] ), .B(\i_MIPS/n314 ), .Y(n4686) );
  AO22X1 U4749 ( .A0(n4980), .A1(n554), .B0(n4976), .B1(n2057), .Y(n6338) );
  AO22X1 U4750 ( .A0(n4978), .A1(n555), .B0(n4976), .B1(n2058), .Y(n6329) );
  AO22X1 U4751 ( .A0(n4978), .A1(n556), .B0(n9309), .B1(n2059), .Y(n6836) );
  NOR2BX4 U4752 ( .AN(n4827), .B(\i_MIPS/n366 ), .Y(n4667) );
  BUFX12 U4753 ( .A(n5485), .Y(n5488) );
  OA22X4 U4754 ( .A0(net112431), .A1(n1955), .B0(net112381), .B1(n380), .Y(
        n6055) );
  OA22X4 U4755 ( .A0(n8659), .A1(n7847), .B0(n7699), .B1(n8437), .Y(n7700) );
  NAND2X8 U4756 ( .A(\i_MIPS/ALUin1[22] ), .B(n6585), .Y(n8250) );
  NAND2BX4 U4757 ( .AN(n5457), .B(n11239), .Y(n9651) );
  AOI21X2 U4758 ( .A0(n7108), .A1(n7785), .B0(n1891), .Y(n4547) );
  INVX8 U4759 ( .A(n4815), .Y(n4810) );
  OA21X4 U4760 ( .A0(\i_MIPS/ALUin1[18] ), .A1(n4819), .B0(n8531), .Y(n8532)
         );
  OAI211X2 U4761 ( .A0(n10366), .A1(n10365), .B0(n10377), .C0(n10497), .Y(
        n10367) );
  AOI211XL U4762 ( .A0(n8998), .A1(n177), .B0(n4670), .C0(n4666), .Y(n9000) );
  AOI21X4 U4763 ( .A0(n7875), .A1(n7874), .B0(n7873), .Y(n4568) );
  AOI2BB1X4 U4764 ( .A0N(\i_MIPS/n343 ), .A1N(n4826), .B0(n4668), .Y(n6355) );
  OAI211X4 U4765 ( .A0(n8430), .A1(n163), .B0(n8429), .C0(n4924), .Y(n8454) );
  AO22X4 U4766 ( .A0(net113457), .A1(n11439), .B0(net113463), .B1(n11408), .Y(
        n7824) );
  AOI222X1 U4767 ( .A0(net109791), .A1(n11408), .B0(mem_rdata_D[19]), .B1(n116), .C0(n12978), .C1(net109801), .Y(n10179) );
  CLKAND2X12 U4768 ( .A(net109181), .B(n11408), .Y(mem_wdata_D[19]) );
  NAND4X2 U4769 ( .A(n7814), .B(n7813), .C(n7812), .D(n7811), .Y(n11408) );
  NAND3BX4 U4770 ( .AN(n9577), .B(n4665), .C(n4662), .Y(n9586) );
  NAND4X8 U4771 ( .A(n9652), .B(n9651), .C(n9654), .D(n9653), .Y(n11073) );
  OA22X4 U4772 ( .A0(n5334), .A1(n3278), .B0(n5290), .B1(n1622), .Y(n6025) );
  OA22X4 U4773 ( .A0(n5334), .A1(n3279), .B0(n5318), .B1(n1623), .Y(n6029) );
  OAI211X2 U4774 ( .A0(n9262), .A1(n7806), .B0(n7805), .C0(n7804), .Y(net99267) );
  OAI211X2 U4775 ( .A0(n6222), .A1(n6221), .B0(n6219), .C0(n6220), .Y(n6445)
         );
  AO22X4 U4776 ( .A0(net113447), .A1(n11471), .B0(net102346), .B1(n11502), .Y(
        n8598) );
  OAI222X2 U4777 ( .A0(n7557), .A1(n7869), .B0(n8819), .B1(n7285), .C0(n4802), 
        .C1(n7970), .Y(n9285) );
  CLKMX2X4 U4778 ( .A(n7872), .B(n7194), .S0(n5590), .Y(n7970) );
  MX2X2 U4779 ( .A(n8444), .B(n7697), .S0(n5589), .Y(n8086) );
  OAI221X4 U4780 ( .A0(\i_MIPS/ALUin1[20] ), .A1(n4810), .B0(
        \i_MIPS/ALUin1[21] ), .B1(n4803), .C0(n6670), .Y(n8444) );
  MX2XL U4781 ( .A(n3492), .B(n3732), .S0(n5507), .Y(\i_MIPS/n395 ) );
  NAND2X6 U4782 ( .A(n3583), .B(net99693), .Y(n4126) );
  NAND2BX4 U4783 ( .AN(n5452), .B(n11339), .Y(n10055) );
  CLKAND2X12 U4784 ( .A(net113916), .B(n11438), .Y(mem_wdata_D[50]) );
  OA22X2 U4785 ( .A0(\i_MIPS/IF_ID[64] ), .A1(net99849), .B0(
        \i_MIPS/IF_ID[64] ), .B1(net98881), .Y(n10256) );
  NAND3BX2 U4786 ( .AN(n8428), .B(n8449), .C(n9258), .Y(n8455) );
  AO21X4 U4787 ( .A0(n4516), .A1(n8427), .B0(n8914), .Y(n8449) );
  AOI222X1 U4788 ( .A0(n5487), .A1(n11438), .B0(mem_rdata_D[50]), .B1(n117), 
        .C0(n12979), .C1(n5483), .Y(n10618) );
  AO21X4 U4789 ( .A0(net99288), .A1(net99289), .B0(net112729), .Y(net104353)
         );
  CLKMX2X2 U4790 ( .A(\i_MIPS/Reg_W[3] ), .B(n10130), .S0(n5511), .Y(
        \i_MIPS/n474 ) );
  INVX3 U4791 ( .A(n6291), .Y(n10130) );
  OAI2BB1X4 U4792 ( .A0N(n6449), .A1N(n8712), .B0(n8711), .Y(n6453) );
  AOI31X2 U4793 ( .A0(n6486), .A1(n6485), .A2(n6484), .B0(n8251), .Y(n6494) );
  NOR4X4 U4794 ( .A(n6631), .B(n6482), .C(n6481), .D(n6480), .Y(n6486) );
  NAND4X2 U4795 ( .A(n8487), .B(n8486), .C(n8485), .D(n8484), .Y(n11476) );
  INVX20 U4796 ( .A(net130576), .Y(net110191) );
  AO21X4 U4797 ( .A0(n10901), .A1(n10900), .B0(n4618), .Y(n10305) );
  CLKAND2X12 U4798 ( .A(net109181), .B(n11396), .Y(mem_wdata_D[7]) );
  NAND4X2 U4799 ( .A(n7491), .B(n7490), .C(n7489), .D(n7488), .Y(n11396) );
  XOR2X4 U4800 ( .A(n178), .B(n4078), .Y(n4073) );
  AO22X2 U4801 ( .A0(net113447), .A1(n11457), .B0(net102346), .B1(n11488), .Y(
        n7331) );
  MX2XL U4802 ( .A(DCACHE_addr[9]), .B(net99039), .S0(n5510), .Y(\i_MIPS/n458 ) );
  AOI222X1 U4803 ( .A0(net109791), .A1(n11395), .B0(mem_rdata_D[5]), .B1(n116), 
        .C0(n12992), .C1(net109801), .Y(n10759) );
  CLKAND2X12 U4804 ( .A(net109181), .B(n11395), .Y(mem_wdata_D[5]) );
  AOI32X2 U4805 ( .A0(n6217), .A1(n6216), .A2(n6215), .B0(n6218), .B1(
        \i_MIPS/ID_EX[75] ), .Y(n6222) );
  MXI2X2 U4806 ( .A(n9280), .B(n9279), .S0(n9278), .Y(n4633) );
  INVX20 U4807 ( .A(n4632), .Y(n9280) );
  OA22XL U4808 ( .A0(net112679), .A1(n1459), .B0(net112573), .B1(n3072), .Y(
        net105032) );
  OA22X1 U4809 ( .A0(net112471), .A1(n1242), .B0(net112347), .B1(n2847), .Y(
        net105033) );
  OA22X1 U4810 ( .A0(net112245), .A1(n1243), .B0(net112163), .B1(n2848), .Y(
        net105034) );
  OA22X1 U4811 ( .A0(net112059), .A1(n1244), .B0(net111935), .B1(n2849), .Y(
        net105035) );
  CLKBUFX3 U4812 ( .A(net112091), .Y(net112059) );
  CLKBUFX3 U4813 ( .A(net111967), .Y(net111935) );
  INVXL U4814 ( .A(net98185), .Y(net100026) );
  XOR2X4 U4815 ( .A(n4086), .B(net99064), .Y(n4081) );
  XOR2X4 U4816 ( .A(n4085), .B(n3317), .Y(n4079) );
  AO21X4 U4817 ( .A0(net99334), .A1(net99335), .B0(net113077), .Y(net99316) );
  XOR2X4 U4818 ( .A(n4083), .B(n4084), .Y(n4082) );
  AOI22X2 U4819 ( .A0(net113041), .A1(net99447), .B0(net102300), .B1(net105373), .Y(net134107) );
  OAI221X2 U4820 ( .A0(net104868), .A1(net112709), .B0(net104831), .B1(
        net112723), .C0(net104869), .Y(net98915) );
  XOR2X4 U4821 ( .A(net100015), .B(n4076), .Y(n4074) );
  OAI221X2 U4822 ( .A0(net105003), .A1(net112709), .B0(net105004), .B1(
        net112723), .C0(net105005), .Y(net100015) );
  CLKINVX3 U4823 ( .A(net105120), .Y(net99089) );
  NAND4X8 U4824 ( .A(net102400), .B(n4071), .C(net102397), .D(net102398), .Y(
        net99850) );
  NAND2XL U4825 ( .A(net113533), .B(net113089), .Y(net100019) );
  AND2XL U4826 ( .A(n3198), .B(net100013), .Y(net130474) );
  AO22X1 U4827 ( .A0(net113445), .A1(net98121), .B0(net102346), .B1(net98089), 
        .Y(n4077) );
  BUFX20 U4828 ( .A(net102345), .Y(net113445) );
  AO21X4 U4829 ( .A0(net100019), .A1(net100020), .B0(net112729), .Y(net105005)
         );
  AND2XL U4830 ( .A(n4140), .B(n4141), .Y(net130420) );
  INVX1 U4831 ( .A(net99759), .Y(n4139) );
  NAND4X1 U4832 ( .A(net100748), .B(net100749), .C(net100750), .D(net100751), 
        .Y(net99759) );
  CLKINVX1 U4833 ( .A(net99933), .Y(n4142) );
  AOI32X2 U4834 ( .A0(net98880), .A1(net131142), .A2(net126164), .B0(net99850), 
        .B1(n4145), .Y(n4144) );
  AND2X2 U4835 ( .A(\i_MIPS/IF_ID[97] ), .B(\i_MIPS/n233 ), .Y(net126164) );
  CLKINVX1 U4836 ( .A(net99664), .Y(n4145) );
  NOR2X8 U4837 ( .A(n3812), .B(n4031), .Y(net102400) );
  XNOR2X4 U4838 ( .A(n4123), .B(net99401), .Y(n4101) );
  OAI2BB1X2 U4839 ( .A0N(net99405), .A1N(net114113), .B0(net113083), .Y(
        net99387) );
  XNOR2X4 U4840 ( .A(net99555), .B(n4124), .Y(n4103) );
  OR2X8 U4841 ( .A(net140551), .B(net113075), .Y(net99541) );
  XNOR2X4 U4842 ( .A(n4122), .B(n4025), .Y(n4104) );
  XOR2X4 U4843 ( .A(n4532), .B(n4135), .Y(n4096) );
  INVX12 U4844 ( .A(net130301), .Y(net112707) );
  AO21X4 U4845 ( .A0(net99603), .A1(net99604), .B0(net112729), .Y(net103392)
         );
  XNOR2X4 U4846 ( .A(n4126), .B(net99531), .Y(n4098) );
  XOR2X4 U4847 ( .A(n182), .B(n4134), .Y(n4091) );
  AO21X4 U4848 ( .A0(net100103), .A1(net100104), .B0(net113075), .Y(net99450)
         );
  XNOR2X4 U4849 ( .A(net99354), .B(n4125), .Y(n4093) );
  AO21X4 U4850 ( .A0(net99359), .A1(net99360), .B0(net113075), .Y(n4141) );
  XOR2X4 U4851 ( .A(net99654), .B(n4527), .Y(n4094) );
  AOI22X4 U4852 ( .A0(net113039), .A1(net99971), .B0(net102300), .B1(net102500), .Y(net134093) );
  AO21X4 U4853 ( .A0(net99969), .A1(net99970), .B0(net113075), .Y(net99671) );
  XOR2X4 U4854 ( .A(net98946), .B(n4114), .Y(n4107) );
  XOR2X4 U4855 ( .A(net99056), .B(n4113), .Y(n4108) );
  AO21X2 U4856 ( .A0(net99060), .A1(net99061), .B0(net113077), .Y(net99042) );
  XOR2X4 U4857 ( .A(net99576), .B(n4112), .Y(n4109) );
  XOR2X4 U4858 ( .A(n4029), .B(n4111), .Y(n4110) );
  OAI221X2 U4859 ( .A0(net105929), .A1(net112709), .B0(net105930), .B1(
        net112723), .C0(net105931), .Y(net99607) );
  XOR2X4 U4860 ( .A(net99009), .B(n4120), .Y(n4115) );
  AO21X2 U4861 ( .A0(net99014), .A1(net99015), .B0(net113075), .Y(net99936) );
  XOR2X4 U4862 ( .A(net98988), .B(n4119), .Y(n4116) );
  AO21X2 U4863 ( .A0(net98992), .A1(net98993), .B0(net113079), .Y(net98974) );
  XOR2X4 U4864 ( .A(n4127), .B(n4128), .Y(n4117) );
  AO21X4 U4865 ( .A0(net98970), .A1(net98971), .B0(net112723), .Y(net98898) );
  NAND2X1 U4866 ( .A(net112713), .B(net106881), .Y(net98900) );
  NAND2X1 U4867 ( .A(net102300), .B(net106535), .Y(net99476) );
  NAND3BX4 U4868 ( .AN(n11155), .B(n11154), .C(n11153), .Y(\i_MIPS/PC/n53 ) );
  NAND2X2 U4869 ( .A(net112607), .B(n11389), .Y(n10151) );
  OA22X4 U4870 ( .A0(net112041), .A1(n2404), .B0(net111917), .B1(n898), .Y(
        n6162) );
  AO22X4 U4871 ( .A0(net113455), .A1(n11447), .B0(net113461), .B1(n11416), .Y(
        n8690) );
  AO22X2 U4872 ( .A0(net113455), .A1(n11444), .B0(net113461), .B1(n11413), .Y(
        n8974) );
  NAND2X4 U4873 ( .A(n6659), .B(\i_MIPS/n342 ), .Y(n9150) );
  NAND2X2 U4874 ( .A(n11226), .B(n9150), .Y(n6669) );
  NAND2X2 U4875 ( .A(\i_MIPS/ALUin1[29] ), .B(n6658), .Y(n11226) );
  NAND2X8 U4876 ( .A(n6170), .B(n6171), .Y(net100095) );
  NAND3BX4 U4877 ( .AN(n9581), .B(n9580), .C(n9579), .Y(n9584) );
  INVX8 U4878 ( .A(n6577), .Y(n6569) );
  BUFX20 U4879 ( .A(n4981), .Y(n4984) );
  OAI211X4 U4880 ( .A0(n8724), .A1(n7880), .B0(n7782), .C0(n4501), .Y(n7796)
         );
  OAI221X4 U4881 ( .A0(net112663), .A1(n1631), .B0(net112561), .B1(n3296), 
        .C0(n6160), .Y(n6161) );
  NAND2X6 U4882 ( .A(n3736), .B(n10668), .Y(n6155) );
  NAND4X2 U4883 ( .A(n8012), .B(n8011), .C(n8010), .D(n8009), .Y(n11442) );
  OAI221X4 U4884 ( .A0(n6442), .A1(n3638), .B0(n7367), .B1(n8817), .C0(n6441), 
        .Y(net106977) );
  OA22X4 U4885 ( .A0(net112089), .A1(n1956), .B0(net111915), .B1(n381), .Y(
        n6132) );
  BUFX20 U4886 ( .A(net112187), .Y(net112143) );
  BUFX4 U4887 ( .A(net112377), .Y(net112355) );
  OAI32X2 U4888 ( .A0(n8651), .A1(n4798), .A2(n4594), .B0(n8650), .B1(n1987), 
        .Y(n8653) );
  BUFX4 U4889 ( .A(net112339), .Y(net112363) );
  BUFX4 U4890 ( .A(net112339), .Y(net112359) );
  BUFX4 U4891 ( .A(net112333), .Y(net112357) );
  CLKAND2X12 U4892 ( .A(net113607), .B(n11475), .Y(mem_wdata_D[88]) );
  NAND4X2 U4893 ( .A(n8105), .B(n8104), .C(n8103), .D(n8102), .Y(n11441) );
  AND3X2 U4894 ( .A(n4665), .B(n9548), .C(n4662), .Y(n9564) );
  OA22XL U4895 ( .A0(net112667), .A1(n1460), .B0(net112565), .B1(n3073), .Y(
        n7810) );
  NAND4X4 U4896 ( .A(n7810), .B(n7809), .C(n7808), .D(n7807), .Y(n11439) );
  NAND4X2 U4897 ( .A(n8483), .B(n8482), .C(n8481), .D(n8480), .Y(n11414) );
  OA22XL U4898 ( .A0(net112667), .A1(n1461), .B0(net112565), .B1(n3074), .Y(
        n8483) );
  AO21X4 U4899 ( .A0(n7612), .A1(n7875), .B0(n7613), .Y(n7695) );
  INVX16 U4900 ( .A(n4502), .Y(n4503) );
  INVX1 U4901 ( .A(n10952), .Y(n10953) );
  AOI222X1 U4902 ( .A0(n5475), .A1(n11492), .B0(mem_rdata_D[106]), .B1(n116), 
        .C0(n12987), .C1(n5473), .Y(n10584) );
  OAI211X2 U4903 ( .A0(n11225), .A1(n9160), .B0(n9158), .C0(n9159), .Y(n9261)
         );
  AO22X4 U4904 ( .A0(net113455), .A1(n11440), .B0(net113461), .B1(n11409), .Y(
        n8599) );
  BUFX20 U4905 ( .A(net112165), .Y(net112155) );
  NAND4X2 U4906 ( .A(n8765), .B(n8764), .C(n8763), .D(n8762), .Y(n11424) );
  NAND4X2 U4907 ( .A(n6860), .B(n6859), .C(n6858), .D(n6857), .Y(n6862) );
  BUFX12 U4908 ( .A(net111965), .Y(net111937) );
  NAND4X2 U4909 ( .A(n7729), .B(n7728), .C(n7727), .D(n7726), .Y(n11468) );
  NAND4BX2 U4910 ( .AN(n7167), .B(n7166), .C(n7165), .D(n7164), .Y(n7178) );
  OA22XL U4911 ( .A0(\i_MIPS/Register/register[4][11] ), .A1(n4952), .B0(
        \i_MIPS/Register/register[12][11] ), .B1(n4949), .Y(n7166) );
  NAND3BX4 U4912 ( .AN(n9571), .B(n4651), .C(n4685), .Y(n9560) );
  MXI2X1 U4913 ( .A(n10545), .B(n10544), .S0(n5493), .Y(n10546) );
  NAND2X6 U4914 ( .A(n10630), .B(n3311), .Y(n6054) );
  OAI211X2 U4915 ( .A0(n7410), .A1(n7409), .B0(net113437), .C0(n3709), .Y(
        net100049) );
  CLKAND2X12 U4916 ( .A(net109181), .B(n11394), .Y(mem_wdata_D[4]) );
  AOI222X4 U4917 ( .A0(n5474), .A1(n11511), .B0(mem_rdata_D[125]), .B1(n116), 
        .C0(n12968), .C1(n5472), .Y(n10475) );
  NAND4X4 U4918 ( .A(n6875), .B(n6874), .C(n6873), .D(n6872), .Y(n11398) );
  OA22X1 U4919 ( .A0(net112679), .A1(n1245), .B0(net112577), .B1(n2850), .Y(
        n6875) );
  OA22X2 U4920 ( .A0(net112235), .A1(n938), .B0(net112165), .B1(n2463), .Y(
        n6873) );
  OAI211X4 U4921 ( .A0(n6885), .A1(n6884), .B0(net113437), .C0(net112607), .Y(
        net99061) );
  AO21X4 U4922 ( .A0(net99334), .A1(net99335), .B0(net112727), .Y(net105579)
         );
  OA22X2 U4923 ( .A0(net112465), .A1(n939), .B0(net112341), .B1(n2464), .Y(
        n7245) );
  AO22X2 U4924 ( .A0(net113457), .A1(n11443), .B0(net113463), .B1(n11412), .Y(
        n8305) );
  AO22X2 U4925 ( .A0(net113457), .A1(n11438), .B0(net113463), .B1(n11407), .Y(
        n7929) );
  AO22X1 U4926 ( .A0(net113447), .A1(n11482), .B0(net102346), .B1(n11513), .Y(
        n9099) );
  OAI211X4 U4927 ( .A0(n6286), .A1(n6285), .B0(net113437), .C0(net112607), .Y(
        net99015) );
  INVX3 U4928 ( .A(n10717), .Y(n10721) );
  INVX3 U4929 ( .A(n10322), .Y(n10329) );
  OA22X2 U4930 ( .A0(n5332), .A1(n458), .B0(n5289), .B1(n2012), .Y(n5996) );
  AO22X1 U4931 ( .A0(net113445), .A1(n11473), .B0(net102346), .B1(n11504), .Y(
        n8025) );
  AO22X4 U4932 ( .A0(n10568), .A1(net113039), .B0(net102300), .B1(n8956), .Y(
        net102651) );
  NAND4X4 U4933 ( .A(n7818), .B(n7817), .C(n7816), .D(n7815), .Y(n11470) );
  NOR3BX4 U4934 ( .AN(n4724), .B(n10936), .C(n11105), .Y(n10939) );
  AO21X4 U4935 ( .A0(n9010), .A1(n7785), .B0(n1891), .Y(n9006) );
  OAI221X4 U4936 ( .A0(\i_MIPS/n340 ), .A1(n4824), .B0(\i_MIPS/n341 ), .B1(
        n4816), .C0(n6223), .Y(n7365) );
  CLKAND2X3 U4937 ( .A(n10448), .B(n10447), .Y(net140551) );
  AO21X4 U4938 ( .A0(n10447), .A1(n10448), .B0(net112729), .Y(net103871) );
  OAI211X2 U4939 ( .A0(n8402), .A1(n8401), .B0(net113439), .C0(net112607), .Y(
        n10408) );
  XOR2X4 U4940 ( .A(n10736), .B(net111405), .Y(n10725) );
  XOR2X4 U4941 ( .A(n10716), .B(ICACHE_addr[29]), .Y(n10736) );
  NAND2X2 U4942 ( .A(n10715), .B(ICACHE_addr[28]), .Y(n10716) );
  AO21X4 U4943 ( .A0(net99429), .A1(net99428), .B0(net112729), .Y(net104025)
         );
  BUFX8 U4944 ( .A(net112519), .Y(net112499) );
  NAND4X4 U4945 ( .A(n8769), .B(n8768), .C(n8767), .D(n8766), .Y(n11393) );
  OA22X2 U4946 ( .A0(net112487), .A1(n2441), .B0(net112363), .B1(n466), .Y(
        n8768) );
  BUFX16 U4947 ( .A(net111979), .Y(net111967) );
  OA22X2 U4948 ( .A0(\i_MIPS/n367 ), .A1(n4812), .B0(\i_MIPS/n366 ), .B1(n4805), .Y(n6358) );
  AOI21X4 U4949 ( .A0(net111405), .A1(net99753), .B0(n4610), .Y(n4599) );
  CLKMX2X6 U4950 ( .A(n7194), .B(n7557), .S0(n5589), .Y(n7876) );
  NAND2X4 U4951 ( .A(n10307), .B(n10209), .Y(n10911) );
  OAI22X4 U4952 ( .A0(n10689), .A1(net102094), .B0(n10692), .B1(net102095), 
        .Y(n4603) );
  INVX3 U4953 ( .A(n11450), .Y(n10692) );
  BUFX20 U4954 ( .A(n3722), .Y(net112153) );
  BUFX20 U4955 ( .A(n3722), .Y(net112151) );
  NAND2X8 U4956 ( .A(n6228), .B(\i_MIPS/n363 ), .Y(n6847) );
  OAI221X2 U4957 ( .A0(net100082), .A1(n1886), .B0(net112139), .B1(n319), .C0(
        n6061), .Y(n6062) );
  OAI222X4 U4958 ( .A0(n8438), .A1(n8437), .B0(n8436), .B1(n8660), .C0(n8659), 
        .C1(n8435), .Y(n8447) );
  OAI222X4 U4959 ( .A0(n9007), .A1(n8434), .B0(n8451), .B1(n8805), .C0(n9004), 
        .C1(n8433), .Y(n8448) );
  CLKINVX20 U4960 ( .A(n4790), .Y(mem_addr_D[29]) );
  INVX4 U4961 ( .A(n4770), .Y(n4790) );
  AOI211X2 U4962 ( .A0(n8822), .A1(n7610), .B0(n6862), .C0(n6861), .Y(n6863)
         );
  AO21X4 U4963 ( .A0(n3666), .A1(n4802), .B0(n7788), .Y(n8727) );
  OA22X2 U4964 ( .A0(n5248), .A1(n448), .B0(n5203), .B1(n3243), .Y(n5993) );
  BUFX20 U4965 ( .A(n5361), .Y(n5333) );
  OA22XL U4966 ( .A0(net112667), .A1(n1462), .B0(net112565), .B1(n3075), .Y(
        n8299) );
  OA22XL U4967 ( .A0(net112667), .A1(n1463), .B0(net112565), .B1(n3076), .Y(
        n8388) );
  OA22XL U4968 ( .A0(net112667), .A1(n1464), .B0(net112565), .B1(n3077), .Y(
        n8303) );
  OA22XL U4969 ( .A0(net112667), .A1(n1465), .B0(net112565), .B1(n3078), .Y(
        n8585) );
  BUFX20 U4970 ( .A(n5361), .Y(n5332) );
  AO22X1 U4971 ( .A0(net113447), .A1(n11452), .B0(net102346), .B1(n11483), .Y(
        n6543) );
  AO22X1 U4972 ( .A0(net113447), .A1(n11480), .B0(net102346), .B1(n11511), .Y(
        n6722) );
  AO22X1 U4973 ( .A0(net113447), .A1(n11459), .B0(net102346), .B1(n11490), .Y(
        n6801) );
  AO22X1 U4974 ( .A0(net113447), .A1(n11460), .B0(net102346), .B1(n11491), .Y(
        n6884) );
  OA22X1 U4975 ( .A0(\i_MIPS/ALUin1[23] ), .A1(n4811), .B0(\i_MIPS/ALUin1[24] ), .B1(n4804), .Y(n8885) );
  OAI221X4 U4976 ( .A0(\i_MIPS/n371 ), .A1(n4818), .B0(\i_MIPS/n369 ), .B1(
        n4804), .C0(n6946), .Y(n8819) );
  OAI221X4 U4977 ( .A0(\i_MIPS/n347 ), .A1(n4810), .B0(\i_MIPS/n348 ), .B1(
        n4804), .C0(n7019), .Y(n7783) );
  OAI221X4 U4978 ( .A0(\i_MIPS/n361 ), .A1(n4810), .B0(\i_MIPS/n360 ), .B1(
        n4804), .C0(n7037), .Y(n8265) );
  AOI32X2 U4979 ( .A0(n6664), .A1(n9014), .A2(n6663), .B0(n9019), .B1(n6662), 
        .Y(n6683) );
  AO21X4 U4980 ( .A0(n8087), .A1(n7875), .B0(n7613), .Y(n7699) );
  OA22X2 U4981 ( .A0(\i_MIPS/n350 ), .A1(n4812), .B0(\i_MIPS/n351 ), .B1(n4805), .Y(n6258) );
  OAI221X4 U4982 ( .A0(\i_MIPS/n348 ), .A1(n4826), .B0(\i_MIPS/n349 ), .B1(
        n4818), .C0(n6258), .Y(n6764) );
  OA22X2 U4983 ( .A0(n5332), .A1(n1630), .B0(n5289), .B1(n3293), .Y(n5982) );
  OA22X2 U4984 ( .A0(n11079), .A1(net140280), .B0(net98430), .B1(n11078), .Y(
        n11081) );
  XOR2X4 U4985 ( .A(n3245), .B(n6118), .Y(n6129) );
  CLKAND2X12 U4986 ( .A(net113608), .B(n11485), .Y(mem_wdata_D[98]) );
  OAI211X4 U4987 ( .A0(n7501), .A1(n7500), .B0(net113439), .C0(n3709), .Y(
        net99109) );
  MX2X2 U4988 ( .A(n7196), .B(n6954), .S0(n5590), .Y(n7555) );
  OAI211X4 U4989 ( .A0(\i_MIPS/ALUin1[16] ), .A1(n4818), .B0(n8531), .C0(n6952), .Y(n7196) );
  NAND2XL U4990 ( .A(n10651), .B(n10650), .Y(n11527) );
  OA22X4 U4991 ( .A0(net112093), .A1(n1957), .B0(net111969), .B1(n385), .Y(
        n6057) );
  NAND4X2 U4992 ( .A(n6713), .B(n6712), .C(n6711), .D(n6710), .Y(n11418) );
  AO22X1 U4993 ( .A0(net113455), .A1(n11449), .B0(net113461), .B1(n11418), .Y(
        n6723) );
  CLKAND2X12 U4994 ( .A(net109181), .B(n11418), .Y(mem_wdata_D[29]) );
  OAI211X4 U4995 ( .A0(n6723), .A1(n6722), .B0(net113437), .C0(n3709), .Y(
        net99503) );
  NAND4X4 U4996 ( .A(n8020), .B(n8019), .C(n8018), .D(n8017), .Y(n11473) );
  NAND4X4 U4997 ( .A(n10104), .B(n10103), .C(n10102), .D(n10101), .Y(n10295)
         );
  AOI2BB1X4 U4998 ( .A0N(\i_MIPS/n344 ), .A1N(n4826), .B0(n4670), .Y(n6259) );
  CLKAND2X3 U4999 ( .A(n4820), .B(\i_MIPS/ALUin1[26] ), .Y(n4670) );
  NAND2BX4 U5000 ( .AN(n5456), .B(n11235), .Y(n9626) );
  XOR2X4 U5001 ( .A(n4748), .B(n6148), .Y(n6158) );
  OAI33X4 U5002 ( .A0(n3657), .A1(n3600), .A2(n9185), .B0(n9183), .B1(n9185), 
        .B2(n9262), .Y(n9186) );
  NAND2X4 U5003 ( .A(n4660), .B(n4656), .Y(n4487) );
  AO21X4 U5004 ( .A0(net99537), .A1(net99536), .B0(net112729), .Y(net103061)
         );
  AOI222X2 U5005 ( .A0(n4554), .A1(n7279), .B0(n7278), .B1(n7277), .C0(n7276), 
        .C1(n7275), .Y(n7292) );
  NAND2X8 U5006 ( .A(\i_MIPS/ALUin1[5] ), .B(n3788), .Y(n7459) );
  OA22XL U5007 ( .A0(net112491), .A1(n1466), .B0(net112355), .B1(n3079), .Y(
        n8112) );
  OA22XL U5008 ( .A0(net112233), .A1(n2851), .B0(net112151), .B1(n845), .Y(
        n8111) );
  CLKMX2X4 U5009 ( .A(n8542), .B(n6776), .S0(n5590), .Y(n8145) );
  INVX3 U5010 ( .A(n8145), .Y(n8887) );
  XOR3X2 U5011 ( .A(n11075), .B(n11074), .C(n11073), .Y(n11077) );
  OAI211X4 U5012 ( .A0(n6394), .A1(n6393), .B0(net113437), .C0(n3709), .Y(
        net98993) );
  NAND2X4 U5013 ( .A(n10274), .B(n10273), .Y(n10302) );
  NAND4X4 U5014 ( .A(n9677), .B(n9676), .C(n9675), .D(n9674), .Y(n10273) );
  XOR2X4 U5015 ( .A(n6123), .B(n3244), .Y(n6128) );
  BUFX20 U5016 ( .A(n11205), .Y(n5481) );
  AO22X2 U5017 ( .A0(net113445), .A1(n11477), .B0(net102346), .B1(n11508), .Y(
        n8401) );
  OA22X4 U5018 ( .A0(net112237), .A1(n2414), .B0(net112155), .B1(n905), .Y(
        n8682) );
  OA22X2 U5019 ( .A0(net112237), .A1(n2442), .B0(net112155), .B1(n467), .Y(
        n8767) );
  OA22X2 U5020 ( .A0(net112237), .A1(n942), .B0(net112155), .B1(n2467), .Y(
        n8763) );
  OA22XL U5021 ( .A0(net112237), .A1(n1467), .B0(net112155), .B1(n3080), .Y(
        n8587) );
  OA22XL U5022 ( .A0(net112237), .A1(n1468), .B0(net112155), .B1(n3081), .Y(
        n8674) );
  OAI2BB1X4 U5023 ( .A0N(n7190), .A1N(n7187), .B0(n7186), .Y(n7098) );
  OAI221X4 U5024 ( .A0(\i_MIPS/n341 ), .A1(n4824), .B0(\i_MIPS/n342 ), .B1(
        n4816), .C0(n7020), .Y(n7791) );
  AO22X1 U5025 ( .A0(n5000), .A1(n218), .B0(n4996), .B1(n2170), .Y(n6917) );
  CLKAND2X12 U5026 ( .A(net113607), .B(n11447), .Y(mem_wdata_D[59]) );
  CLKINVX1 U5027 ( .A(n11447), .Y(n10471) );
  NAND4X2 U5028 ( .A(n8676), .B(n8675), .C(n8674), .D(n8673), .Y(n11447) );
  NAND2X2 U5029 ( .A(n7284), .B(n4707), .Y(n8085) );
  NAND4X2 U5030 ( .A(n8773), .B(n8772), .C(n8771), .D(n8770), .Y(n11455) );
  OA22XL U5031 ( .A0(net112237), .A1(n2852), .B0(net112155), .B1(n846), .Y(
        n8775) );
  INVX3 U5032 ( .A(n6165), .Y(n10658) );
  OA22X2 U5033 ( .A0(net112235), .A1(n944), .B0(net112153), .B1(n2469), .Y(
        n7808) );
  NAND3BX4 U5034 ( .AN(n4425), .B(n4503), .C(n4424), .Y(n11136) );
  INVXL U5035 ( .A(n4794), .Y(n4334) );
  INVXL U5036 ( .A(n4794), .Y(n4323) );
  XOR2X4 U5037 ( .A(n3252), .B(n6115), .Y(n6130) );
  MXI2X4 U5038 ( .A(n10593), .B(n10592), .S0(n5492), .Y(n10594) );
  AOI222X4 U5039 ( .A0(n5487), .A1(n11430), .B0(mem_rdata_D[42]), .B1(n117), 
        .C0(n12987), .C1(n5483), .Y(n10593) );
  BUFX20 U5040 ( .A(n5485), .Y(n5487) );
  NAND3BX2 U5041 ( .AN(n8655), .B(n4550), .C(n9156), .Y(n8656) );
  NAND4BX4 U5042 ( .AN(n8101), .B(n8100), .C(n8099), .D(n3247), .Y(net99430)
         );
  AOI2BB1X1 U5043 ( .A0N(\i_MIPS/ALUin1[17] ), .A1N(n4806), .B0(n4597), .Y(
        n6671) );
  OAI221X2 U5044 ( .A0(net112263), .A1(n711), .B0(net112137), .B1(n221), .C0(
        n6045), .Y(n6046) );
  CLKAND2X12 U5045 ( .A(net113607), .B(n11478), .Y(mem_wdata_D[91]) );
  NAND4X4 U5046 ( .A(n8680), .B(n8679), .C(n8678), .D(n8677), .Y(n11416) );
  OA22X2 U5047 ( .A0(net112665), .A1(n945), .B0(net112555), .B1(n2470), .Y(
        n8680) );
  OAI222X1 U5048 ( .A0(n4424), .A1(net110213), .B0(net130474), .B1(net110243), 
        .C0(n11067), .C1(net110247), .Y(n11072) );
  NOR4X8 U5049 ( .A(n6069), .B(n6071), .C(n6070), .D(n6072), .Y(n6073) );
  OA22XL U5050 ( .A0(net112665), .A1(n1469), .B0(net112565), .B1(n3082), .Y(
        n8850) );
  OA22XL U5051 ( .A0(net112237), .A1(n1470), .B0(net112155), .B1(n3083), .Y(
        n8848) );
  NAND4BX2 U5052 ( .AN(n6703), .B(n6702), .C(n6701), .D(n6700), .Y(n6704) );
  AO22X1 U5053 ( .A0(n5000), .A1(n219), .B0(n4996), .B1(n2171), .Y(n6908) );
  XOR2X4 U5054 ( .A(n6104), .B(n12942), .Y(n6110) );
  NAND2X6 U5055 ( .A(n10645), .B(n10644), .Y(n6104) );
  AOI222X1 U5056 ( .A0(net109791), .A1(n11396), .B0(mem_rdata_D[7]), .B1(n116), 
        .C0(n12990), .C1(net109801), .Y(n10745) );
  CLKAND2X12 U5057 ( .A(n8818), .B(n8348), .Y(n4554) );
  NAND3BX4 U5058 ( .AN(n7372), .B(n7371), .C(n7370), .Y(net99447) );
  NAND4X4 U5059 ( .A(n8862), .B(n8861), .C(n8860), .D(n8859), .Y(n11485) );
  OA22XL U5060 ( .A0(net112665), .A1(n1471), .B0(net112565), .B1(n3084), .Y(
        n8858) );
  OA22XL U5061 ( .A0(net112237), .A1(n1472), .B0(net112155), .B1(n3085), .Y(
        n8856) );
  INVX8 U5062 ( .A(n9137), .Y(n9283) );
  NAND3BX4 U5063 ( .AN(n4425), .B(n4005), .C(n4424), .Y(n11135) );
  NAND2BX4 U5064 ( .AN(n10328), .B(n10322), .Y(n10948) );
  AO21X4 U5065 ( .A0(net111409), .A1(n11020), .B0(n4609), .Y(n10328) );
  AND2X8 U5066 ( .A(n4599), .B(n10498), .Y(n4564) );
  NAND4X2 U5067 ( .A(n4696), .B(n9582), .C(n4697), .D(n4694), .Y(n9551) );
  AOI2BB2X2 U5068 ( .B0(\i_MIPS/IF_ID[96] ), .B1(n147), .A0N(net110189), .A1N(
        \i_MIPS/n211 ), .Y(n10733) );
  INVXL U5069 ( .A(n8665), .Y(n8667) );
  CLKAND2X12 U5070 ( .A(n4796), .B(n11357), .Y(mem_wdata_I[127]) );
  CLKAND2X12 U5071 ( .A(net109181), .B(n11392), .Y(mem_wdata_D[2]) );
  AO22XL U5072 ( .A0(net113457), .A1(n11422), .B0(net113463), .B1(n11391), .Y(
        n7650) );
  OAI221X4 U5073 ( .A0(\i_MIPS/n371 ), .A1(n4824), .B0(\i_MIPS/n370 ), .B1(
        n4816), .C0(n7038), .Y(n7473) );
  NAND3BX4 U5074 ( .AN(n6444), .B(n4567), .C(n6263), .Y(n7968) );
  MX2X1 U5075 ( .A(n9141), .B(n4799), .S0(n7036), .Y(n7045) );
  OA22X2 U5076 ( .A0(n11003), .A1(net140280), .B0(n11002), .B1(net98430), .Y(
        n11005) );
  OAI222X2 U5077 ( .A0(n9610), .A1(n5454), .B0(n9609), .B1(n5452), .C0(n9608), 
        .C1(n5456), .Y(n11181) );
  CLKAND2X12 U5078 ( .A(net113606), .B(n11486), .Y(mem_wdata_D[99]) );
  AO22X4 U5079 ( .A0(n7858), .A1(n6627), .B0(n6627), .B1(n7776), .Y(n6648) );
  INVX20 U5080 ( .A(n4722), .Y(n4723) );
  NAND4X4 U5081 ( .A(n10001), .B(n10000), .C(n9999), .D(n9998), .Y(n10906) );
  NAND3BX4 U5082 ( .AN(n6784), .B(n6782), .C(n6783), .Y(net98952) );
  BUFX20 U5083 ( .A(net112687), .Y(net112673) );
  NAND2X2 U5084 ( .A(n4601), .B(net112607), .Y(n10695) );
  XOR2X4 U5085 ( .A(n3253), .B(n6095), .Y(n6096) );
  XOR2X4 U5086 ( .A(n10376), .B(ICACHE_addr[26]), .Y(n10390) );
  NAND2X2 U5087 ( .A(n10486), .B(ICACHE_addr[25]), .Y(n10376) );
  INVX12 U5088 ( .A(n10390), .Y(n10500) );
  AOI211X2 U5089 ( .A0(n8908), .A1(n9283), .B0(n8907), .C0(n8906), .Y(n8934)
         );
  OAI33X2 U5090 ( .A0(n4020), .A1(n8904), .A2(n9262), .B0(n9262), .B1(n8903), 
        .B2(n3548), .Y(n8907) );
  NAND2X4 U5091 ( .A(n4809), .B(\i_MIPS/ALUin1[30] ), .Y(n9274) );
  BUFX20 U5092 ( .A(n4513), .Y(n5476) );
  CLKAND2X12 U5093 ( .A(n10161), .B(n10147), .Y(n4513) );
  NOR2X2 U5094 ( .A(n135), .B(n186), .Y(net114092) );
  XOR2X4 U5095 ( .A(n3254), .B(n6042), .Y(n6076) );
  INVX4 U5096 ( .A(n6039), .Y(n10635) );
  OAI222X4 U5097 ( .A0(n3709), .A1(n4669), .B0(net113919), .B1(net100096), 
        .C0(mem_ready_D), .C1(n11389), .Y(n10158) );
  OAI221X2 U5098 ( .A0(net112657), .A1(n712), .B0(net112563), .B1(n3249), .C0(
        n6082), .Y(n6083) );
  AOI2BB1X4 U5099 ( .A0N(n11012), .A1N(n11011), .B0(n11010), .Y(n11014) );
  OA22X4 U5100 ( .A0(n9615), .A1(n5452), .B0(n9612), .B1(n5457), .Y(n9613) );
  NAND2BX4 U5101 ( .AN(n7097), .B(n3747), .Y(n7190) );
  OA22X2 U5102 ( .A0(n3611), .A1(n1612), .B0(n5383), .B1(n3294), .Y(n5987) );
  NAND3BX4 U5103 ( .AN(n10211), .B(n10307), .C(n3598), .Y(n10910) );
  NAND2BX4 U5104 ( .AN(n5458), .B(n11232), .Y(n9605) );
  AOI221X2 U5105 ( .A0(n7470), .A1(n7469), .B0(n7468), .B1(n7467), .C0(n7466), 
        .Y(n7482) );
  OA21X2 U5106 ( .A0(\i_MIPS/n365 ), .A1(n4826), .B0(n7281), .Y(n6357) );
  AO21X4 U5107 ( .A0(n8645), .A1(n4801), .B0(n8643), .Y(n8649) );
  NAND2X4 U5108 ( .A(n7785), .B(n9130), .Y(n7880) );
  NAND2X2 U5109 ( .A(n10344), .B(n10349), .Y(n10378) );
  XOR2X4 U5110 ( .A(n3246), .B(n6047), .Y(n6075) );
  OA22X4 U5111 ( .A0(net112429), .A1(n1959), .B0(net112301), .B1(n387), .Y(
        n6043) );
  AO21X4 U5112 ( .A0(net99383), .A1(net99382), .B0(net112729), .Y(net103709)
         );
  CLKAND2X12 U5113 ( .A(net113608), .B(n11492), .Y(mem_wdata_D[106]) );
  XOR2X4 U5114 ( .A(n3255), .B(n6050), .Y(n6074) );
  OA22X4 U5115 ( .A0(net112431), .A1(n1960), .B0(net112301), .B1(n388), .Y(
        n6048) );
  BUFX20 U5116 ( .A(n4575), .Y(n5482) );
  AOI222X1 U5117 ( .A0(n5486), .A1(n11447), .B0(mem_rdata_D[59]), .B1(n116), 
        .C0(n12970), .C1(n5482), .Y(n10472) );
  AOI222X4 U5118 ( .A0(n8822), .A1(n4593), .B0(n4568), .B1(n3599), .C0(n8820), 
        .C1(n8819), .Y(n8825) );
  OA22X4 U5119 ( .A0(net112089), .A1(n1961), .B0(net111915), .B1(n389), .Y(
        n6153) );
  NAND2X6 U5120 ( .A(n4198), .B(net112607), .Y(net99335) );
  NAND3BX4 U5121 ( .AN(n11360), .B(n11359), .C(n11358), .Y(n11363) );
  INVX8 U5122 ( .A(n9328), .Y(n11360) );
  AOI22X1 U5123 ( .A0(ICACHE_addr[26]), .A1(mem_read_I), .B0(n4796), .B1(
        n11385), .Y(n4147) );
  XOR2X4 U5124 ( .A(n3256), .B(n6134), .Y(n6141) );
  OA22X1 U5125 ( .A0(net112665), .A1(n1246), .B0(net112563), .B1(n2853), .Y(
        n8117) );
  BUFX8 U5126 ( .A(net112269), .Y(net112259) );
  AO21X4 U5127 ( .A0(n7612), .A1(n7785), .B0(n1891), .Y(n6673) );
  AOI211X2 U5128 ( .A0(n7200), .A1(n7290), .B0(n6371), .C0(n6370), .Y(n6372)
         );
  OAI221X2 U5129 ( .A0(net112265), .A1(n2045), .B0(net112139), .B1(n705), .C0(
        n6079), .Y(n6080) );
  NAND2X4 U5130 ( .A(n4778), .B(\i_MIPS/n334 ), .Y(n10139) );
  OAI221X2 U5131 ( .A0(net112265), .A1(n713), .B0(net112143), .B1(n3250), .C0(
        n6084), .Y(n6085) );
  AOI222X1 U5132 ( .A0(net109795), .A1(n11400), .B0(mem_rdata_D[11]), .B1(n116), .C0(n12986), .C1(net109805), .Y(n10784) );
  AOI2BB1X4 U5133 ( .A0N(n4602), .A1N(n4603), .B0(net100096), .Y(n4601) );
  NAND4X8 U5134 ( .A(n4459), .B(n4460), .C(n5978), .D(n5977), .Y(n11373) );
  OAI2BB1X4 U5135 ( .A0N(n10319), .A1N(n10318), .B0(n10323), .Y(n10964) );
  AOI211X2 U5136 ( .A0(n8654), .A1(n9283), .B0(n8653), .C0(n8652), .Y(n8670)
         );
  NAND4BX4 U5137 ( .AN(n8671), .B(n8670), .C(n8669), .D(n8668), .Y(net99538)
         );
  OAI221X2 U5138 ( .A0(net112657), .A1(n2046), .B0(net112563), .B1(n706), .C0(
        n6091), .Y(n6092) );
  CLKAND2X12 U5139 ( .A(net113606), .B(n11487), .Y(mem_wdata_D[100]) );
  AOI2BB1X2 U5140 ( .A0N(\i_MIPS/n355 ), .A1N(n4806), .B0(n4690), .Y(n6262) );
  OR4X8 U5141 ( .A(n9189), .B(n9186), .C(n9187), .D(n9188), .Y(n10629) );
  BUFX20 U5142 ( .A(n5274), .Y(n5250) );
  NAND2X2 U5143 ( .A(n4444), .B(net110253), .Y(n10734) );
  BUFX20 U5144 ( .A(net112517), .Y(net112507) );
  BUFX4 U5145 ( .A(n11212), .Y(n5485) );
  INVX4 U5146 ( .A(n6147), .Y(n10664) );
  OAI221X2 U5147 ( .A0(net112231), .A1(n2048), .B0(net112139), .B1(n320), .C0(
        n6146), .Y(n6147) );
  OA22X4 U5148 ( .A0(net112041), .A1(n1963), .B0(net111915), .B1(n391), .Y(
        n6146) );
  NAND4X8 U5149 ( .A(n9619), .B(n9618), .C(n9617), .D(n9616), .Y(n11063) );
  NAND2BX4 U5150 ( .AN(n5456), .B(n11234), .Y(n9618) );
  NAND2BX2 U5151 ( .AN(n10275), .B(n10302), .Y(n10277) );
  BUFX20 U5152 ( .A(n5274), .Y(n5249) );
  OAI221X2 U5153 ( .A0(net112659), .A1(n2049), .B0(net112575), .B1(n708), .C0(
        n6105), .Y(n6106) );
  OA22X4 U5154 ( .A0(net112449), .A1(n1964), .B0(net112325), .B1(n392), .Y(
        n6105) );
  OAI221X2 U5155 ( .A0(net112229), .A1(n2051), .B0(net112145), .B1(n710), .C0(
        n6107), .Y(n6108) );
  OA22X4 U5156 ( .A0(net112037), .A1(n1965), .B0(net111905), .B1(n393), .Y(
        n6107) );
  OAI221X2 U5157 ( .A0(net112241), .A1(n3258), .B0(net112143), .B1(n1615), 
        .C0(n6102), .Y(n6103) );
  INVX4 U5158 ( .A(n6103), .Y(n10644) );
  CLKXOR2X8 U5159 ( .A(n3314), .B(n4445), .Y(net98881) );
  BUFX20 U5160 ( .A(n5316), .Y(n5289) );
  CLKINVX4 U5161 ( .A(n6474), .Y(n6464) );
  XOR3X4 U5162 ( .A(net111409), .B(n10699), .C(n4544), .Y(n4543) );
  OA22X4 U5163 ( .A0(n5333), .A1(n1966), .B0(n5290), .B1(n394), .Y(n6012) );
  BUFX20 U5164 ( .A(n5316), .Y(n5290) );
  XOR2X4 U5165 ( .A(n11536), .B(n12944), .Y(n6109) );
  NAND2X4 U5166 ( .A(n10296), .B(n10295), .Y(n10917) );
  OAI221X4 U5167 ( .A0(\i_MIPS/n364 ), .A1(n4825), .B0(\i_MIPS/n363 ), .B1(
        n4817), .C0(n6949), .Y(n7194) );
  OAI221X4 U5168 ( .A0(\i_MIPS/n366 ), .A1(n4810), .B0(\i_MIPS/n365 ), .B1(
        n4803), .C0(n6945), .Y(n7557) );
  OAI221X2 U5169 ( .A0(net112697), .A1(n1887), .B0(net112583), .B1(n321), .C0(
        n6055), .Y(n6056) );
  BUFX20 U5170 ( .A(n4925), .Y(n4928) );
  OA22X2 U5171 ( .A0(n10357), .A1(net140281), .B0(net98430), .B1(n10363), .Y(
        n10359) );
  AOI33X4 U5172 ( .A0(n9258), .A1(n3698), .A2(n7884), .B0(n9258), .B1(n7862), 
        .B2(n7854), .Y(n7891) );
  OAI221X2 U5173 ( .A0(n8265), .A1(n7867), .B0(n7285), .B1(n7473), .C0(n7041), 
        .Y(n9129) );
  AOI2BB1X4 U5174 ( .A0N(n10954), .A1N(n4608), .B0(n10953), .Y(n10955) );
  AOI222X2 U5175 ( .A0(n6844), .A1(n3636), .B0(n6775), .B1(n6774), .C0(n6773), 
        .C1(n6772), .Y(n6783) );
  AO22X4 U5176 ( .A0(n6770), .A1(n4924), .B0(n9258), .B1(n6845), .Y(n6773) );
  OAI221X4 U5177 ( .A0(n4798), .A1(n6845), .B0(n6770), .B1(n9262), .C0(n8805), 
        .Y(n6774) );
  INVX1 U5178 ( .A(n6106), .Y(n10642) );
  MXI2X1 U5179 ( .A(n10514), .B(n10513), .S0(n5494), .Y(n10515) );
  AOI221X2 U5180 ( .A0(net140278), .A1(n11189), .B0(n3546), .B1(n11187), .C0(
        net98447), .Y(n11190) );
  OAI31X2 U5181 ( .A0(n6626), .A1(n6625), .A2(n6624), .B0(n7852), .Y(n7776) );
  AO21X4 U5182 ( .A0(n6633), .A1(n6632), .B0(n6472), .Y(n6473) );
  NAND3X4 U5183 ( .A(ICACHE_addr[12]), .B(ICACHE_addr[11]), .C(n10261), .Y(
        n10294) );
  NAND2X2 U5184 ( .A(net98880), .B(net131142), .Y(n11185) );
  OAI221X4 U5185 ( .A0(n9284), .A1(n8275), .B0(n9007), .B1(n8274), .C0(n4501), 
        .Y(n8276) );
  NAND2X4 U5186 ( .A(\i_MIPS/ALUin1[8] ), .B(n6228), .Y(n6771) );
  NAND2BX2 U5187 ( .AN(n5457), .B(n11241), .Y(n9971) );
  AO22X1 U5188 ( .A0(net113457), .A1(n11437), .B0(net113463), .B1(n11406), .Y(
        n7735) );
  OR2X1 U5189 ( .A(net112693), .B(n2350), .Y(n4148) );
  OR2X1 U5190 ( .A(n7560), .B(n7869), .Y(n4150) );
  INVX1 U5191 ( .A(n7874), .Y(n7560) );
  OR2X2 U5192 ( .A(n5383), .B(n2026), .Y(n4153) );
  NAND2BX4 U5193 ( .AN(n7799), .B(n4515), .Y(n8514) );
  OR2X8 U5194 ( .A(n4611), .B(n10870), .Y(n4156) );
  NAND2X6 U5195 ( .A(n4155), .B(n4156), .Y(n4586) );
  CLKAND2X8 U5196 ( .A(n10872), .B(n10871), .Y(n4611) );
  INVX3 U5197 ( .A(n9625), .Y(n10870) );
  NAND2X6 U5198 ( .A(n6589), .B(\i_MIPS/n347 ), .Y(n8905) );
  MX2XL U5199 ( .A(n9209), .B(n9208), .S0(net108959), .Y(n9212) );
  CLKAND2X12 U5200 ( .A(n6263), .B(n6447), .Y(n4585) );
  AND2X2 U5201 ( .A(n6447), .B(n8648), .Y(n6497) );
  NAND2X4 U5202 ( .A(\i_MIPS/ALUin1[10] ), .B(n6244), .Y(n7193) );
  NAND2X8 U5203 ( .A(n4587), .B(n4578), .Y(n8536) );
  NAND2X8 U5204 ( .A(n4577), .B(n4587), .Y(n9004) );
  OR2X1 U5205 ( .A(\i_MIPS/PC/n17 ), .B(net110213), .Y(n4172) );
  OR2X1 U5206 ( .A(\i_MIPS/PC/n16 ), .B(net110215), .Y(n4175) );
  OAI211X2 U5207 ( .A0(n10283), .A1(n10282), .B0(n10281), .C0(n10280), .Y(
        n10285) );
  AND2X2 U5208 ( .A(mem_rdata_D[0]), .B(n117), .Y(n4179) );
  BUFX12 U5209 ( .A(net98396), .Y(net109795) );
  NAND4X4 U5210 ( .A(n6534), .B(n6533), .C(n6532), .D(n6531), .Y(n11390) );
  INVXL U5211 ( .A(net113075), .Y(net140445) );
  XNOR3X2 U5212 ( .A(n11196), .B(n11192), .C(n3516), .Y(n11194) );
  OA22X4 U5213 ( .A0(net112033), .A1(n1967), .B0(net111931), .B1(n395), .Y(
        n6089) );
  AO21X4 U5214 ( .A0(n8664), .A1(n3816), .B0(n8663), .Y(n4188) );
  OR2X1 U5215 ( .A(\i_MIPS/PC/n15 ), .B(net110213), .Y(n4189) );
  XOR3X2 U5216 ( .A(n11085), .B(n11084), .C(n11083), .Y(n11087) );
  OAI211X2 U5217 ( .A0(n3610), .A1(n3502), .B0(n10815), .C0(n10816), .Y(
        \i_MIPS/PC/n34 ) );
  OAI221X4 U5218 ( .A0(n7867), .A1(n7286), .B0(n4797), .B1(n7611), .C0(n7476), 
        .Y(n8434) );
  OA21X4 U5219 ( .A0(n7248), .A1(n7247), .B0(net113437), .Y(n4198) );
  NOR2X2 U5220 ( .A(net112037), .B(n1894), .Y(n4206) );
  NAND2X2 U5221 ( .A(n4613), .B(n9579), .Y(n9337) );
  OR2X1 U5222 ( .A(n6934), .B(n6930), .Y(n4208) );
  NAND2BX4 U5223 ( .AN(n7094), .B(n6639), .Y(n6927) );
  BUFX16 U5224 ( .A(net112693), .Y(net112659) );
  OR2X1 U5225 ( .A(\i_MIPS/PC/n20 ), .B(net110215), .Y(n4212) );
  XOR2XL U5226 ( .A(n11093), .B(n11095), .Y(n4215) );
  XOR2X4 U5227 ( .A(n11094), .B(n4215), .Y(n11097) );
  OA21X4 U5228 ( .A0(n7332), .A1(n7331), .B0(net113437), .Y(n4216) );
  NAND2X6 U5229 ( .A(n4216), .B(net112607), .Y(net100039) );
  NAND2X2 U5230 ( .A(net100038), .B(net100039), .Y(n10764) );
  AO21X2 U5231 ( .A0(net100038), .A1(net100039), .B0(net112727), .Y(net105427)
         );
  OAI211X2 U5232 ( .A0(n6649), .A1(n6648), .B0(n6646), .C0(n6647), .Y(n9154)
         );
  INVXL U5233 ( .A(n4488), .Y(n4751) );
  CLKAND2X12 U5234 ( .A(net113608), .B(n11495), .Y(mem_wdata_D[109]) );
  BUFX8 U5235 ( .A(n11204), .Y(n4231) );
  BUFX8 U5236 ( .A(n10803), .Y(n4232) );
  BUFX8 U5237 ( .A(n10791), .Y(n4233) );
  BUFX8 U5238 ( .A(n10779), .Y(n4234) );
  BUFX8 U5239 ( .A(n11171), .Y(n4235) );
  BUFX8 U5240 ( .A(n10166), .Y(n4247) );
  BUFX8 U5241 ( .A(n10144), .Y(n4248) );
  BUFX8 U5242 ( .A(n10168), .Y(n4249) );
  BUFX8 U5243 ( .A(n10150), .Y(n4250) );
  BUFX8 U5244 ( .A(n10156), .Y(n4252) );
  XOR3X1 U5245 ( .A(net111405), .B(n11118), .C(n11117), .Y(n11146) );
  BUFX8 U5246 ( .A(n10476), .Y(n4254) );
  BUFX8 U5247 ( .A(n10397), .Y(n4255) );
  BUFX8 U5248 ( .A(n10413), .Y(n4257) );
  BUFX8 U5249 ( .A(n10558), .Y(n4259) );
  BUFX8 U5250 ( .A(n10174), .Y(n4261) );
  BUFX8 U5251 ( .A(n10585), .Y(n4264) );
  BUFX8 U5252 ( .A(n10688), .Y(n4266) );
  BUFX8 U5253 ( .A(n10416), .Y(n4269) );
  BUFX8 U5254 ( .A(n10428), .Y(n4270) );
  BUFX8 U5255 ( .A(n10561), .Y(n4271) );
  BUFX8 U5256 ( .A(n10525), .Y(n4273) );
  BUFX8 U5257 ( .A(n10177), .Y(n4274) );
  BUFX8 U5258 ( .A(n10454), .Y(n4275) );
  BUFX8 U5259 ( .A(n10191), .Y(n4276) );
  BUFX8 U5260 ( .A(n10440), .Y(n4277) );
  BUFX8 U5261 ( .A(n10770), .Y(n4278) );
  BUFX8 U5262 ( .A(n10743), .Y(n4279) );
  BUFX8 U5263 ( .A(n10757), .Y(n4280) );
  BUFX8 U5264 ( .A(n10512), .Y(n4281) );
  BUFX8 U5265 ( .A(n10691), .Y(n4303) );
  BUFX8 U5266 ( .A(n10419), .Y(n4306) );
  BUFX8 U5267 ( .A(n10431), .Y(n4307) );
  BUFX8 U5268 ( .A(n10540), .Y(n4311) );
  BUFX8 U5269 ( .A(n10528), .Y(n4312) );
  BUFX8 U5270 ( .A(n10616), .Y(n4313) );
  AO22X1 U5271 ( .A0(net113455), .A1(n11431), .B0(net113461), .B1(n11400), .Y(
        n7158) );
  XOR2X4 U5272 ( .A(n10270), .B(n10271), .Y(n10214) );
  AO21X4 U5273 ( .A0(net100048), .A1(net100049), .B0(net112727), .Y(net105286)
         );
  XOR3X2 U5274 ( .A(net111409), .B(n10381), .C(n10367), .Y(n10369) );
  NAND2X2 U5275 ( .A(n11107), .B(n10937), .Y(n10330) );
  CLKINVX6 U5276 ( .A(n11107), .Y(n10936) );
  NAND2X4 U5277 ( .A(n3515), .B(n9678), .Y(n11047) );
  AOI33X2 U5278 ( .A0(n3866), .A1(n9258), .A2(n8931), .B0(n8928), .B1(n8929), 
        .B2(n9258), .Y(n8932) );
  OAI211X2 U5279 ( .A0(n8927), .A1(n8926), .B0(n8924), .C0(n8925), .Y(n8930)
         );
  CLKMX2X2 U5280 ( .A(\i_MIPS/ALUin1[2] ), .B(net98449), .S0(n5505), .Y(
        \i_MIPS/n560 ) );
  OAI31X2 U5281 ( .A0(n10383), .A1(n4595), .A2(n10382), .B0(n10488), .Y(n10384) );
  NAND3BX4 U5282 ( .AN(n8341), .B(n4924), .C(n8340), .Y(n8363) );
  NAND3BX2 U5283 ( .AN(n7983), .B(n4924), .C(n7982), .Y(n7984) );
  MX2X2 U5284 ( .A(n4799), .B(n9141), .S0(n8095), .Y(n8096) );
  OAI211X4 U5285 ( .A0(n8329), .A1(n6590), .B0(n6614), .C0(n4516), .Y(n9167)
         );
  XOR2X4 U5286 ( .A(n11372), .B(ICACHE_addr[13]), .Y(n9566) );
  AOI21X4 U5287 ( .A0(n7710), .A1(n7709), .B0(n7708), .Y(n4520) );
  AOI33X4 U5288 ( .A0(n9015), .A1(n9171), .A2(n6654), .B0(n6653), .B1(n3562), 
        .B2(n11224), .Y(n6685) );
  OAI221X2 U5289 ( .A0(n8527), .A1(n7859), .B0(n7858), .B1(n7857), .C0(n7856), 
        .Y(n7885) );
  OAI211X4 U5290 ( .A0(net114031), .A1(net99664), .B0(n10389), .C0(n10388), 
        .Y(n10732) );
  OA21X1 U5291 ( .A0(\i_MIPS/ALUin1[13] ), .A1(n4819), .B0(n7104), .Y(n7105)
         );
  CLKAND2X12 U5292 ( .A(net113916), .B(n11473), .Y(mem_wdata_D[86]) );
  CLKAND2X12 U5293 ( .A(net113916), .B(n11470), .Y(mem_wdata_D[83]) );
  CLKAND2X12 U5294 ( .A(net113916), .B(n11468), .Y(mem_wdata_D[81]) );
  CLKAND2X12 U5295 ( .A(net113916), .B(n11441), .Y(mem_wdata_D[53]) );
  CLKAND2X12 U5296 ( .A(net113916), .B(n11439), .Y(mem_wdata_D[51]) );
  CLKAND2X12 U5297 ( .A(net113608), .B(n11442), .Y(mem_wdata_D[54]) );
  CLKAND2X12 U5298 ( .A(net113608), .B(n11510), .Y(mem_wdata_D[124]) );
  CLKAND2X12 U5299 ( .A(net113916), .B(n11474), .Y(mem_wdata_D[87]) );
  INVX20 U5300 ( .A(n4321), .Y(mem_addr_I[16]) );
  NOR2X2 U5301 ( .A(n4322), .B(n4323), .Y(n4325) );
  NOR2X2 U5302 ( .A(n4324), .B(\i_MIPS/PC/n18 ), .Y(n4326) );
  NOR2X8 U5303 ( .A(n4325), .B(n4326), .Y(n4321) );
  INVXL U5304 ( .A(n11371), .Y(n4328) );
  CLKINVX1 U5305 ( .A(mem_read_I), .Y(n4329) );
  INVX20 U5306 ( .A(n4332), .Y(mem_addr_I[13]) );
  CLKINVX1 U5307 ( .A(n11370), .Y(n4333) );
  CLKINVX1 U5308 ( .A(mem_read_I), .Y(n4335) );
  NOR2X2 U5309 ( .A(n4333), .B(n4334), .Y(n4336) );
  NOR2X2 U5310 ( .A(n4335), .B(\i_MIPS/PC/n15 ), .Y(n4337) );
  NOR2X8 U5311 ( .A(n4336), .B(n4337), .Y(n4332) );
  INVX20 U5312 ( .A(n4338), .Y(mem_addr_I[11]) );
  INVXL U5313 ( .A(n11368), .Y(n4339) );
  NOR2X2 U5314 ( .A(n4339), .B(n11361), .Y(n4340) );
  NOR2X2 U5315 ( .A(n4335), .B(\i_MIPS/PC/n13 ), .Y(n4341) );
  NOR2X8 U5316 ( .A(n4340), .B(n4341), .Y(n4338) );
  INVX20 U5317 ( .A(n4342), .Y(mem_addr_I[7]) );
  NOR2X2 U5318 ( .A(n4343), .B(n11361), .Y(n4344) );
  NOR2X8 U5319 ( .A(n4344), .B(n4345), .Y(n4342) );
  INVX20 U5320 ( .A(n4346), .Y(mem_addr_I[15]) );
  INVXL U5321 ( .A(n11372), .Y(n4347) );
  NOR2X2 U5322 ( .A(n4347), .B(n4348), .Y(n4350) );
  NOR2X2 U5323 ( .A(n4349), .B(\i_MIPS/PC/n17 ), .Y(n4351) );
  NOR2X6 U5324 ( .A(n4350), .B(n4351), .Y(n4346) );
  CLKAND2X12 U5325 ( .A(net109185), .B(n11437), .Y(mem_wdata_D[49]) );
  CLKAND2X12 U5326 ( .A(net113608), .B(n11450), .Y(mem_wdata_D[62]) );
  CLKAND2X12 U5327 ( .A(net113916), .B(n11466), .Y(mem_wdata_D[79]) );
  CLKAND2X12 U5328 ( .A(n4796), .B(n11272), .Y(mem_wdata_I[42]) );
  CLKAND2X12 U5329 ( .A(n4796), .B(n11270), .Y(mem_wdata_I[40]) );
  CLKAND2X12 U5330 ( .A(n4796), .B(n11268), .Y(mem_wdata_I[38]) );
  CLKAND2X12 U5331 ( .A(n4794), .B(n11266), .Y(mem_wdata_I[36]) );
  INVX12 U5332 ( .A(\i_MIPS/n310 ), .Y(DCACHE_wen) );
  INVX12 U5333 ( .A(\i_MIPS/n248 ), .Y(DCACHE_wdata[30]) );
  INVX12 U5334 ( .A(\i_MIPS/n278 ), .Y(DCACHE_wdata[15]) );
  INVX12 U5335 ( .A(\i_MIPS/n280 ), .Y(DCACHE_wdata[14]) );
  INVX12 U5336 ( .A(\i_MIPS/n250 ), .Y(DCACHE_wdata[29]) );
  INVX12 U5337 ( .A(\i_MIPS/n254 ), .Y(DCACHE_wdata[27]) );
  INVX12 U5338 ( .A(\i_MIPS/n256 ), .Y(DCACHE_wdata[26]) );
  INVX12 U5339 ( .A(\i_MIPS/n260 ), .Y(DCACHE_wdata[24]) );
  INVX12 U5340 ( .A(\i_MIPS/n268 ), .Y(DCACHE_wdata[20]) );
  INVX12 U5341 ( .A(\i_MIPS/n272 ), .Y(DCACHE_wdata[18]) );
  INVX12 U5342 ( .A(\i_MIPS/n274 ), .Y(DCACHE_wdata[17]) );
  INVX12 U5343 ( .A(\i_MIPS/n276 ), .Y(DCACHE_wdata[16]) );
  INVX12 U5344 ( .A(\i_MIPS/n282 ), .Y(DCACHE_wdata[13]) );
  INVX12 U5345 ( .A(\i_MIPS/n284 ), .Y(DCACHE_wdata[12]) );
  INVX12 U5346 ( .A(\i_MIPS/n286 ), .Y(DCACHE_wdata[11]) );
  INVX12 U5347 ( .A(\i_MIPS/n290 ), .Y(DCACHE_wdata[9]) );
  INVX12 U5348 ( .A(\i_MIPS/n292 ), .Y(DCACHE_wdata[8]) );
  INVX12 U5349 ( .A(\i_MIPS/n252 ), .Y(DCACHE_wdata[28]) );
  INVX12 U5350 ( .A(\i_MIPS/n258 ), .Y(DCACHE_wdata[25]) );
  INVX12 U5351 ( .A(\i_MIPS/n262 ), .Y(DCACHE_wdata[23]) );
  INVX12 U5352 ( .A(\i_MIPS/n264 ), .Y(DCACHE_wdata[22]) );
  INVX12 U5353 ( .A(\i_MIPS/n266 ), .Y(DCACHE_wdata[21]) );
  INVX12 U5354 ( .A(\i_MIPS/n270 ), .Y(DCACHE_wdata[19]) );
  INVX12 U5355 ( .A(\i_MIPS/n288 ), .Y(DCACHE_wdata[10]) );
  INVX12 U5356 ( .A(\i_MIPS/n294 ), .Y(DCACHE_wdata[7]) );
  INVX12 U5357 ( .A(\i_MIPS/n296 ), .Y(net139803) );
  INVX12 U5358 ( .A(\i_MIPS/n298 ), .Y(DCACHE_wdata[5]) );
  INVX12 U5359 ( .A(\i_MIPS/n300 ), .Y(DCACHE_wdata[4]) );
  INVX12 U5360 ( .A(\i_MIPS/n302 ), .Y(DCACHE_wdata[3]) );
  INVX12 U5361 ( .A(\i_MIPS/n304 ), .Y(DCACHE_wdata[2]) );
  INVX12 U5362 ( .A(\i_MIPS/n306 ), .Y(DCACHE_wdata[1]) );
  INVX12 U5363 ( .A(\i_MIPS/n308 ), .Y(DCACHE_wdata[0]) );
  INVX12 U5364 ( .A(\i_MIPS/n246 ), .Y(DCACHE_wdata[31]) );
  AO22XL U5365 ( .A0(n12941), .A1(mem_read_D), .B0(net113608), .B1(n11539), 
        .Y(n4770) );
  INVX12 U5366 ( .A(n4385), .Y(DCACHE_addr[22]) );
  INVX16 U5367 ( .A(n2315), .Y(DCACHE_addr[20]) );
  INVX16 U5368 ( .A(n3252), .Y(DCACHE_addr[7]) );
  INVX16 U5369 ( .A(n3199), .Y(DCACHE_addr[14]) );
  INVX16 U5370 ( .A(n3256), .Y(DCACHE_addr[18]) );
  INVX16 U5371 ( .A(n3251), .Y(DCACHE_addr[25]) );
  INVX16 U5372 ( .A(n3253), .Y(DCACHE_addr[9]) );
  INVX12 U5373 ( .A(n4393), .Y(DCACHE_addr[24]) );
  INVX12 U5374 ( .A(n4395), .Y(DCACHE_addr[26]) );
  AO22XL U5375 ( .A0(n12942), .A1(mem_read_D), .B0(net109183), .B1(n11538), 
        .Y(n4769) );
  INVX16 U5376 ( .A(n3255), .Y(DCACHE_addr[5]) );
  NAND2XL U5377 ( .A(n12963), .B(net113089), .Y(net99108) );
  INVX16 U5378 ( .A(n285), .Y(DCACHE_addr[11]) );
  NAND2XL U5379 ( .A(n12957), .B(net113087), .Y(net98992) );
  INVX16 U5380 ( .A(n3254), .Y(DCACHE_addr[13]) );
  NAND2XL U5381 ( .A(n12955), .B(net113087), .Y(net99977) );
  INVX16 U5382 ( .A(n283), .Y(DCACHE_addr[12]) );
  INVX16 U5383 ( .A(n3246), .Y(DCACHE_addr[28]) );
  AO22XL U5384 ( .A0(DCACHE_addr[28]), .A1(mem_read_D), .B0(net113608), .B1(
        n11540), .Y(n4771) );
  NAND2X1 U5385 ( .A(n12940), .B(\i_MIPS/n336 ), .Y(n10696) );
  INVX16 U5386 ( .A(n3245), .Y(DCACHE_addr[8]) );
  INVX16 U5387 ( .A(n3244), .Y(DCACHE_addr[6]) );
  OR2X1 U5388 ( .A(\i_MIPS/PC/n14 ), .B(net110215), .Y(n4404) );
  OR2X6 U5389 ( .A(n10916), .B(n10915), .Y(n4407) );
  NAND3X4 U5390 ( .A(n4407), .B(n4408), .C(n4590), .Y(n11103) );
  AOI211X2 U5391 ( .A0(n9013), .A1(n9283), .B0(n9011), .C0(n9012), .Y(n9023)
         );
  OR2X1 U5392 ( .A(\i_MIPS/PC/n27 ), .B(net110215), .Y(n4415) );
  OR2X1 U5393 ( .A(\i_MIPS/PC/n22 ), .B(net110213), .Y(n4420) );
  NAND3X6 U5394 ( .A(n4420), .B(n4421), .C(n4422), .Y(n11023) );
  NOR2XL U5395 ( .A(\i_MIPS/PC/n5 ), .B(net110215), .Y(n4429) );
  INVXL U5396 ( .A(n11000), .Y(n11001) );
  BUFX12 U5397 ( .A(net112507), .Y(net112449) );
  INVX3 U5398 ( .A(n5008), .Y(n5007) );
  BUFX2 U5399 ( .A(net112503), .Y(net112467) );
  BUFX2 U5400 ( .A(n5450), .Y(n5423) );
  CLKBUFX4 U5401 ( .A(n4910), .Y(n4913) );
  OR2XL U5402 ( .A(net113725), .B(n10462), .Y(n4775) );
  CLKBUFX2 U5403 ( .A(n5402), .Y(n5390) );
  CLKBUFX2 U5404 ( .A(n5141), .Y(n5126) );
  INVX8 U5405 ( .A(n4871), .Y(n4865) );
  CLKBUFX2 U5406 ( .A(n5141), .Y(n5127) );
  INVX1 U5407 ( .A(n8931), .Y(n8904) );
  NAND3X1 U5408 ( .A(n10157), .B(n10160), .C(n10159), .Y(n11212) );
  INVX1 U5409 ( .A(n4693), .Y(n5462) );
  BUFX4 U5410 ( .A(n4630), .Y(n4955) );
  AOI21X2 U5411 ( .A0(n6347), .A1(n6602), .B0(n6346), .Y(n4636) );
  AO22XL U5412 ( .A0(n4977), .A1(n514), .B0(n4976), .B1(n2267), .Y(n7345) );
  OA22X2 U5413 ( .A0(n5264), .A1(n947), .B0(n5219), .B1(n2472), .Y(n9943) );
  OA22X2 U5414 ( .A0(n5178), .A1(n949), .B0(n5134), .B1(n2474), .Y(n9944) );
  BUFX20 U5415 ( .A(net101983), .Y(net112727) );
  OA22XL U5416 ( .A0(n5430), .A1(n1054), .B0(n5386), .B1(n2626), .Y(n9378) );
  OA22XL U5417 ( .A0(n5165), .A1(n1055), .B0(n5121), .B1(n2627), .Y(n9381) );
  OA22XL U5418 ( .A0(n5251), .A1(n1056), .B0(n5205), .B1(n2628), .Y(n9380) );
  OA22XL U5419 ( .A0(n5441), .A1(n2854), .B0(n5395), .B1(n847), .Y(n9937) );
  AO22XL U5420 ( .A0(n5000), .A1(n246), .B0(n4996), .B1(n1874), .Y(n7600) );
  AO22XL U5421 ( .A0(n5000), .A1(n247), .B0(n4996), .B1(n1875), .Y(n7591) );
  OA22XL U5422 ( .A0(n5445), .A1(n1057), .B0(n5399), .B1(n2629), .Y(n10223) );
  OA22X1 U5423 ( .A0(n5342), .A1(n2506), .B0(n5298), .B1(n744), .Y(n9671) );
  OA22X2 U5424 ( .A0(n5349), .A1(n2444), .B0(n5305), .B1(n469), .Y(n9942) );
  OA22X1 U5425 ( .A0(n5339), .A1(n736), .B0(n5295), .B1(n2317), .Y(n9514) );
  OA22X1 U5426 ( .A0(n5341), .A1(n2507), .B0(n5297), .B1(n745), .Y(n9647) );
  OA22XL U5427 ( .A0(\i_MIPS/Register/register[4][14] ), .A1(n4953), .B0(
        \i_MIPS/Register/register[12][14] ), .B1(n4948), .Y(n6914) );
  OA22XL U5428 ( .A0(\i_MIPS/Register/register[0][14] ), .A1(n4961), .B0(
        \i_MIPS/Register/register[8][14] ), .B1(n4957), .Y(n6913) );
  NAND3X1 U5429 ( .A(n3647), .B(ICACHE_addr[5]), .C(n9451), .Y(n9431) );
  OA22XL U5430 ( .A0(n5340), .A1(n2526), .B0(n5296), .B1(n774), .Y(n9539) );
  OA22XL U5431 ( .A0(n5349), .A1(n1474), .B0(n5305), .B1(n3087), .Y(n9938) );
  OA22XL U5432 ( .A0(n5335), .A1(n1058), .B0(n5291), .B1(n2630), .Y(n9379) );
  OA22XL U5433 ( .A0(n5342), .A1(n1059), .B0(n5298), .B1(n2631), .Y(n9666) );
  AO22XL U5434 ( .A0(n5000), .A1(n515), .B0(n4996), .B1(n2268), .Y(n7533) );
  AO22XL U5435 ( .A0(n5000), .A1(n516), .B0(n4996), .B1(n2269), .Y(n7524) );
  OA22XL U5436 ( .A0(n5339), .A1(n746), .B0(n5295), .B1(n2325), .Y(n9509) );
  OA22XL U5437 ( .A0(net112051), .A1(n1475), .B0(net111927), .B1(n3088), .Y(
        n7141) );
  OA22XL U5438 ( .A0(net112057), .A1(n1476), .B0(net111933), .B1(n3089), .Y(
        n7401) );
  OA22XL U5439 ( .A0(net112081), .A1(n1477), .B0(net111957), .B1(n3090), .Y(
        n9052) );
  OA22XL U5440 ( .A0(n5343), .A1(n2527), .B0(n5299), .B1(n775), .Y(n9703) );
  AO22XL U5441 ( .A0(n9312), .A1(n255), .B0(n4986), .B1(n2234), .Y(n8611) );
  AO22X1 U5442 ( .A0(n4979), .A1(n557), .B0(n4976), .B1(n2060), .Y(n8612) );
  MX2X2 U5443 ( .A(n8955), .B(n8954), .S0(n5587), .Y(n8956) );
  AOI21X4 U5444 ( .A0(n4778), .A1(n352), .B0(n10158), .Y(n4604) );
  OA22XL U5445 ( .A0(n5257), .A1(n1060), .B0(n5211), .B1(n2632), .Y(n9643) );
  OA22XL U5446 ( .A0(n5171), .A1(n1061), .B0(n5128), .B1(n2633), .Y(n9644) );
  OA22XL U5447 ( .A0(net112071), .A1(n1478), .B0(net111947), .B1(n3091), .Y(
        n8480) );
  CLKBUFX2 U5448 ( .A(n3611), .Y(n5432) );
  INVX3 U5449 ( .A(n8646), .Y(n9166) );
  CLKBUFX2 U5450 ( .A(net101983), .Y(net112731) );
  AO22X1 U5451 ( .A0(n5000), .A1(n558), .B0(n4996), .B1(n2061), .Y(n7674) );
  CLKBUFX2 U5452 ( .A(net112499), .Y(net112485) );
  CLKBUFX3 U5453 ( .A(n5402), .Y(n5389) );
  AO22XL U5454 ( .A0(n4628), .A1(n297), .B0(n4566), .B1(n1870), .Y(n6504) );
  AO22XL U5455 ( .A0(n4628), .A1(n296), .B0(n4566), .B1(n1869), .Y(n6521) );
  OA22XL U5456 ( .A0(\i_MIPS/Register/register[16][14] ), .A1(n4961), .B0(
        \i_MIPS/Register/register[24][14] ), .B1(n4957), .Y(n6922) );
  OA22XL U5457 ( .A0(\i_MIPS/Register/register[17][2] ), .A1(n4834), .B0(
        \i_MIPS/Register/register[25][2] ), .B1(n4830), .Y(n8839) );
  OA22XL U5458 ( .A0(\i_MIPS/Register/register[21][27] ), .A1(n4850), .B0(
        \i_MIPS/Register/register[29][27] ), .B1(n4843), .Y(n8631) );
  OA22XL U5459 ( .A0(\i_MIPS/Register/register[22][2] ), .A1(n4914), .B0(
        \i_MIPS/Register/register[30][2] ), .B1(n4908), .Y(n8840) );
  OA22XL U5460 ( .A0(n5345), .A1(n1062), .B0(n5301), .B1(n2634), .Y(n9795) );
  OA22XL U5461 ( .A0(n5354), .A1(n1063), .B0(n5310), .B1(n2635), .Y(n10224) );
  MX2XL U5462 ( .A(\i_MIPS/ID_EX[69] ), .B(net99654), .S0(n5509), .Y(
        \i_MIPS/n381 ) );
  INVX3 U5463 ( .A(n10251), .Y(n11039) );
  CLKBUFX4 U5464 ( .A(n4943), .Y(n4945) );
  CLKINVX6 U5465 ( .A(n4869), .Y(n4868) );
  AO22X1 U5466 ( .A0(net113457), .A1(n11445), .B0(net113463), .B1(n11414), .Y(
        n8493) );
  INVXL U5467 ( .A(n8067), .Y(n7961) );
  NAND2XL U5468 ( .A(n8712), .B(n8711), .Y(n8722) );
  CLKINVX4 U5469 ( .A(n11517), .Y(n11545) );
  OA22X1 U5470 ( .A0(n5268), .A1(n980), .B0(n5223), .B1(n2528), .Y(n10225) );
  OA22X1 U5471 ( .A0(n5260), .A1(n981), .B0(n5214), .B1(n2529), .Y(n9762) );
  OA22X1 U5472 ( .A0(n5437), .A1(n982), .B0(n5392), .B1(n2530), .Y(n9760) );
  OA22XL U5473 ( .A0(\i_MIPS/Register/register[20][14] ), .A1(n4954), .B0(
        \i_MIPS/Register/register[28][14] ), .B1(n4948), .Y(n6923) );
  OA22X1 U5474 ( .A0(n5336), .A1(n983), .B0(n5292), .B1(n2531), .Y(n9399) );
  OA22XL U5475 ( .A0(\i_MIPS/Register/register[1][5] ), .A1(n4833), .B0(
        \i_MIPS/Register/register[9][5] ), .B1(n4830), .Y(n7297) );
  OA22XL U5476 ( .A0(\i_MIPS/Register/register[5][5] ), .A1(n4849), .B0(
        \i_MIPS/Register/register[13][5] ), .B1(n4841), .Y(n7296) );
  CLKBUFX2 U5477 ( .A(net112499), .Y(net112481) );
  CLKBUFX2 U5478 ( .A(n5421), .Y(n5433) );
  CLKBUFX2 U5479 ( .A(n5142), .Y(n5124) );
  INVX8 U5480 ( .A(n4847), .Y(n4841) );
  INVX6 U5481 ( .A(n4879), .Y(n4874) );
  CLKBUFX3 U5482 ( .A(n3611), .Y(n5435) );
  CLKBUFX2 U5483 ( .A(n5142), .Y(n5122) );
  CLKBUFX2 U5484 ( .A(n3611), .Y(n5431) );
  CLKMX2X2 U5485 ( .A(n4799), .B(n9141), .S0(n8905), .Y(n8906) );
  XOR3X2 U5486 ( .A(net111409), .B(n10343), .C(n10334), .Y(n10336) );
  CLKINVX3 U5487 ( .A(n9138), .Y(n8261) );
  AO22XL U5488 ( .A0(n4977), .A1(n490), .B0(n4976), .B1(n2235), .Y(n7171) );
  OA22XL U5489 ( .A0(n5253), .A1(n1064), .B0(n5207), .B1(n2636), .Y(n9434) );
  OA22XL U5490 ( .A0(n5432), .A1(n1065), .B0(n5388), .B1(n2637), .Y(n9432) );
  OA22XL U5491 ( .A0(n5167), .A1(n1066), .B0(n5123), .B1(n2638), .Y(n9435) );
  INVX1 U5492 ( .A(n7966), .Y(n7967) );
  NAND3BX2 U5493 ( .AN(n11515), .B(n11548), .C(n11514), .Y(n11517) );
  OA22XL U5494 ( .A0(n5442), .A1(n1067), .B0(n5396), .B1(n2639), .Y(n9641) );
  OA22XL U5495 ( .A0(n5254), .A1(n1068), .B0(n5208), .B1(n2640), .Y(n9480) );
  OA22XL U5496 ( .A0(n5433), .A1(n1069), .B0(n5399), .B1(n2641), .Y(n9478) );
  OA22XL U5497 ( .A0(n5168), .A1(n1070), .B0(n5124), .B1(n2642), .Y(n9481) );
  OA22XL U5498 ( .A0(n5256), .A1(n1071), .B0(n5210), .B1(n2643), .Y(n9593) );
  OA22XL U5499 ( .A0(n5431), .A1(n2532), .B0(n5389), .B1(n776), .Y(n9591) );
  OA22XL U5500 ( .A0(n5170), .A1(n1072), .B0(n5126), .B1(n2644), .Y(n9594) );
  OA22X1 U5501 ( .A0(n5265), .A1(n984), .B0(n5220), .B1(n2533), .Y(n9962) );
  OA22X1 U5502 ( .A0(n5442), .A1(n985), .B0(n5396), .B1(n2534), .Y(n9960) );
  OA22X1 U5503 ( .A0(n5179), .A1(n986), .B0(n5135), .B1(n2535), .Y(n9963) );
  INVX6 U5504 ( .A(n312), .Y(n5454) );
  OA22XL U5505 ( .A0(n5183), .A1(n1073), .B0(n5139), .B1(n2645), .Y(n10226) );
  OA22XL U5506 ( .A0(n5174), .A1(n1074), .B0(n5129), .B1(n2646), .Y(n9763) );
  OA22X4 U5507 ( .A0(net112101), .A1(n421), .B0(net111969), .B1(n3261), .Y(
        n6040) );
  OA22XL U5508 ( .A0(n5337), .A1(n2536), .B0(n5293), .B1(n777), .Y(n9433) );
  NAND2X2 U5509 ( .A(n9429), .B(n3645), .Y(n9430) );
  INVX3 U5510 ( .A(n9431), .Y(n9429) );
  AO22XL U5511 ( .A0(n5002), .A1(n491), .B0(n4997), .B1(n2236), .Y(n7259) );
  AO22XL U5512 ( .A0(n5002), .A1(n492), .B0(n4997), .B1(n2237), .Y(n7250) );
  AO22XL U5513 ( .A0(n5002), .A1(n517), .B0(n4997), .B1(n2270), .Y(n7009) );
  AO22XL U5514 ( .A0(n5002), .A1(n518), .B0(n4997), .B1(n2271), .Y(n7000) );
  AO22XL U5515 ( .A0(n5001), .A1(n519), .B0(n4997), .B1(n2272), .Y(n7169) );
  AO22XL U5516 ( .A0(n5002), .A1(n520), .B0(n4997), .B1(n2273), .Y(n7441) );
  AO22XL U5517 ( .A0(n5002), .A1(n521), .B0(n4997), .B1(n2274), .Y(n7160) );
  AO22XL U5518 ( .A0(n5000), .A1(n522), .B0(n4997), .B1(n2275), .Y(n7432) );
  OA22XL U5519 ( .A0(net112679), .A1(n1479), .B0(net112577), .B1(n3092), .Y(
        n6967) );
  OA22XL U5520 ( .A0(net112069), .A1(n1480), .B0(net111945), .B1(n3093), .Y(
        n8199) );
  OA22XL U5521 ( .A0(net112073), .A1(n1481), .B0(net111949), .B1(n3094), .Y(
        n8484) );
  OA22XL U5522 ( .A0(net112079), .A1(n1482), .B0(net111955), .B1(n3095), .Y(
        n9044) );
  OA22XL U5523 ( .A0(net112055), .A1(n1483), .B0(net111931), .B1(n3096), .Y(
        n7327) );
  OA22X4 U5524 ( .A0(net112087), .A1(n423), .B0(net111955), .B1(n3263), .Y(
        n6084) );
  OA22X4 U5525 ( .A0(net112097), .A1(n424), .B0(net111905), .B1(n3264), .Y(
        n6079) );
  OA22XL U5526 ( .A0(\i_MIPS/Register/register[6][11] ), .A1(n4911), .B0(
        \i_MIPS/Register/register[14][11] ), .B1(n4903), .Y(n7125) );
  OA22X1 U5527 ( .A0(n5340), .A1(n737), .B0(n5296), .B1(n2318), .Y(n9543) );
  OA22X1 U5528 ( .A0(net112053), .A1(n1247), .B0(net111929), .B1(n2855), .Y(
        n7149) );
  OA22X1 U5529 ( .A0(net112043), .A1(n1248), .B0(net111919), .B1(n2856), .Y(
        n6531) );
  OA22XL U5530 ( .A0(\i_MIPS/Register/register[1][2] ), .A1(n4834), .B0(
        \i_MIPS/Register/register[9][2] ), .B1(n4829), .Y(n8830) );
  OA22XL U5531 ( .A0(n5341), .A1(n747), .B0(n5297), .B1(n2326), .Y(n9642) );
  OA22XL U5532 ( .A0(n5338), .A1(n2537), .B0(n5294), .B1(n778), .Y(n9479) );
  OA22XL U5533 ( .A0(\i_MIPS/Register/register[17][11] ), .A1(n4833), .B0(
        \i_MIPS/Register/register[25][11] ), .B1(n4830), .Y(n7133) );
  OA22XL U5534 ( .A0(net112043), .A1(n1484), .B0(net111919), .B1(n3097), .Y(
        n6527) );
  OA22XL U5535 ( .A0(net112043), .A1(n1485), .B0(net111919), .B1(n3098), .Y(
        n6381) );
  OA22XL U5536 ( .A0(net112043), .A1(n1486), .B0(net111919), .B1(n3099), .Y(
        n6385) );
  OA22XL U5537 ( .A0(net112053), .A1(n1487), .B0(net111929), .B1(n3100), .Y(
        n7243) );
  OA22XL U5538 ( .A0(\i_MIPS/Register/register[22][11] ), .A1(n4911), .B0(
        \i_MIPS/Register/register[30][11] ), .B1(n4903), .Y(n7134) );
  OA22XL U5539 ( .A0(\i_MIPS/Register/register[22][20] ), .A1(n4913), .B0(
        \i_MIPS/Register/register[30][20] ), .B1(n4907), .Y(n8574) );
  OA22XL U5540 ( .A0(\i_MIPS/Register/register[22][11] ), .A1(n4936), .B0(
        \i_MIPS/Register/register[30][11] ), .B1(n4930), .Y(n7168) );
  OA22XL U5541 ( .A0(n5340), .A1(n2538), .B0(n5296), .B1(n779), .Y(n9592) );
  CLKBUFX3 U5542 ( .A(net111983), .Y(net111963) );
  INVX3 U5543 ( .A(n4880), .Y(n4877) );
  BUFX4 U5544 ( .A(n4970), .Y(n4969) );
  INVX1 U5545 ( .A(n11218), .Y(n11152) );
  INVX1 U5546 ( .A(n10958), .Y(n10960) );
  INVX1 U5547 ( .A(n10370), .Y(n10371) );
  INVX1 U5548 ( .A(n10337), .Y(n10338) );
  INVX1 U5549 ( .A(n10968), .Y(n10970) );
  AO22X1 U5550 ( .A0(net113447), .A1(n11461), .B0(net102346), .B1(n11492), .Y(
        n7247) );
  NAND2BX2 U5551 ( .AN(n5454), .B(n11301), .Y(n9834) );
  NAND2BX2 U5552 ( .AN(n5461), .B(n11269), .Y(n9833) );
  INVXL U5553 ( .A(n7852), .Y(n7778) );
  AOI21X2 U5554 ( .A0(n8661), .A1(n8647), .B0(n6652), .Y(n4563) );
  CLKINVX1 U5555 ( .A(n8440), .Y(n8451) );
  CLKINVX1 U5556 ( .A(n8553), .Y(n8556) );
  BUFX4 U5557 ( .A(net98432), .Y(net110239) );
  AND2X8 U5558 ( .A(net112727), .B(net112723), .Y(net130301) );
  NAND2X2 U5559 ( .A(n4693), .B(n11265), .Y(n9614) );
  INVX1 U5560 ( .A(n7034), .Y(n7027) );
  CLKINVX1 U5561 ( .A(n9277), .Y(n9278) );
  CLKINVX1 U5562 ( .A(n8429), .Y(n8428) );
  CLKBUFX2 U5563 ( .A(n4619), .Y(n4860) );
  NAND4X6 U5564 ( .A(n6010), .B(n6009), .C(n6008), .D(n6007), .Y(n11386) );
  AO21X4 U5565 ( .A0(net111409), .A1(n10959), .B0(n4608), .Y(n10327) );
  CLKINVX3 U5566 ( .A(n7856), .Y(n6625) );
  INVX3 U5567 ( .A(n10389), .Y(n10865) );
  AO22XL U5568 ( .A0(n9312), .A1(n263), .B0(n4986), .B1(n2276), .Y(n8131) );
  AO22XL U5569 ( .A0(n9312), .A1(n264), .B0(n4986), .B1(n2277), .Y(n8122) );
  AO22XL U5570 ( .A0(n9312), .A1(n256), .B0(n4986), .B1(n2238), .Y(n8505) );
  AO22XL U5571 ( .A0(n9312), .A1(n257), .B0(n4986), .B1(n2239), .Y(n8496) );
  AO22XL U5572 ( .A0(n9312), .A1(n258), .B0(n4986), .B1(n2240), .Y(n8317) );
  AO22XL U5573 ( .A0(n9312), .A1(n259), .B0(n4986), .B1(n2241), .Y(n8308) );
  AO22XL U5574 ( .A0(n9312), .A1(n260), .B0(n4986), .B1(n2242), .Y(n8602) );
  AO22XL U5575 ( .A0(n9312), .A1(n261), .B0(n4986), .B1(n2243), .Y(n8220) );
  AO22XL U5576 ( .A0(n9312), .A1(n262), .B0(n4986), .B1(n2244), .Y(n8211) );
  AOI22X4 U5577 ( .A0(net113083), .A1(n9126), .B0(net113167), .B1(n9125), .Y(
        n4605) );
  OA22XL U5578 ( .A0(n5441), .A1(n2857), .B0(n5395), .B1(n848), .Y(n9933) );
  OA22XL U5579 ( .A0(n5178), .A1(n1488), .B0(n5134), .B1(n3101), .Y(n9936) );
  OA22XL U5580 ( .A0(n5264), .A1(n1489), .B0(n5219), .B1(n3102), .Y(n9935) );
  INVX3 U5581 ( .A(n11029), .Y(n11025) );
  INVX3 U5582 ( .A(n11020), .Y(n10292) );
  AOI2BB1XL U5583 ( .A0N(n8800), .A1N(n177), .B0(n6416), .Y(n6442) );
  CLKMX2X2 U5584 ( .A(n6905), .B(n6904), .S0(n5588), .Y(n6906) );
  NOR4X1 U5585 ( .A(n6894), .B(n6893), .C(n6892), .D(n6891), .Y(n6905) );
  CLKMX2X2 U5586 ( .A(n6997), .B(n6996), .S0(n5588), .Y(n6998) );
  CLKMX2X2 U5587 ( .A(n7588), .B(n7587), .S0(n5588), .Y(n7589) );
  NOR4X1 U5588 ( .A(n7577), .B(n7576), .C(n7575), .D(n7574), .Y(n7588) );
  CLKMX2X2 U5589 ( .A(n7521), .B(n7520), .S0(n5588), .Y(n7522) );
  OA22X1 U5590 ( .A0(n5261), .A1(n987), .B0(n5215), .B1(n2539), .Y(n9796) );
  OA22X1 U5591 ( .A0(n5437), .A1(n988), .B0(n5392), .B1(n2540), .Y(n9748) );
  OA22X1 U5592 ( .A0(n5260), .A1(n989), .B0(n5214), .B1(n2541), .Y(n9750) );
  OA22X1 U5593 ( .A0(n5169), .A1(n738), .B0(n5125), .B1(n2319), .Y(n9516) );
  OA22X1 U5594 ( .A0(n5255), .A1(n739), .B0(n5209), .B1(n2320), .Y(n9515) );
  AO22X1 U5595 ( .A0(n4978), .A1(n649), .B0(n9309), .B1(n2172), .Y(n6919) );
  AO22XL U5596 ( .A0(n9312), .A1(n523), .B0(n4981), .B1(n2278), .Y(n7442) );
  AO22XL U5597 ( .A0(n9312), .A1(n493), .B0(n4981), .B1(n2245), .Y(n7433) );
  AO22XL U5598 ( .A0(n9312), .A1(n524), .B0(n4981), .B1(n2279), .Y(n7010) );
  AO22XL U5599 ( .A0(n9312), .A1(n525), .B0(n4981), .B1(n2280), .Y(n7001) );
  AO22XL U5600 ( .A0(n9312), .A1(n526), .B0(n4981), .B1(n2281), .Y(n7335) );
  OA22X1 U5601 ( .A0(n5435), .A1(n990), .B0(n5390), .B1(n2542), .Y(n9665) );
  OA22X1 U5602 ( .A0(n5172), .A1(n991), .B0(n5127), .B1(n2543), .Y(n9668) );
  OA22X1 U5603 ( .A0(n5258), .A1(n992), .B0(n5212), .B1(n2544), .Y(n9667) );
  OA22X1 U5604 ( .A0(n5432), .A1(n993), .B0(n5398), .B1(n2545), .Y(n9821) );
  OA22X1 U5605 ( .A0(n5176), .A1(n994), .B0(n5131), .B1(n2546), .Y(n9824) );
  OA22X1 U5606 ( .A0(n5262), .A1(n995), .B0(n5216), .B1(n2547), .Y(n9823) );
  OA22XL U5607 ( .A0(n5257), .A1(n1075), .B0(n5211), .B1(n2647), .Y(n9648) );
  OA22XL U5608 ( .A0(n5171), .A1(n1076), .B0(n5128), .B1(n2648), .Y(n9649) );
  OA22XL U5609 ( .A0(n5436), .A1(n1077), .B0(n5388), .B1(n2649), .Y(n9826) );
  OA22XL U5610 ( .A0(n5176), .A1(n1078), .B0(n5131), .B1(n2650), .Y(n9829) );
  OA22XL U5611 ( .A0(n5262), .A1(n1079), .B0(n5216), .B1(n2651), .Y(n9828) );
  OA22XL U5612 ( .A0(n5442), .A1(n1080), .B0(n5396), .B1(n2652), .Y(n9965) );
  OA22XL U5613 ( .A0(n5179), .A1(n1081), .B0(n5135), .B1(n2653), .Y(n9968) );
  OA22XL U5614 ( .A0(n5265), .A1(n1082), .B0(n5220), .B1(n2654), .Y(n9967) );
  OAI22X1 U5615 ( .A0(n5172), .A1(n907), .B0(n5127), .B1(n2418), .Y(n4476) );
  OAI22XL U5616 ( .A0(n5166), .A1(n924), .B0(n5122), .B1(n2438), .Y(n4478) );
  OAI22XL U5617 ( .A0(n5168), .A1(n714), .B0(n5124), .B1(n2314), .Y(n4477) );
  INVX1 U5618 ( .A(n10714), .Y(n10715) );
  OA22X1 U5619 ( .A0(net112075), .A1(n2807), .B0(net111951), .B1(n805), .Y(
        n8766) );
  AND2X8 U5620 ( .A(net110227), .B(\i_MIPS/IF_ID[97] ), .Y(n4494) );
  OA22X1 U5621 ( .A0(n5346), .A1(n996), .B0(n5302), .B1(n2548), .Y(n9822) );
  OA22X1 U5622 ( .A0(n5350), .A1(n997), .B0(n5306), .B1(n2549), .Y(n9961) );
  OA22X1 U5623 ( .A0(\i_MIPS/Register/register[21][5] ), .A1(n4849), .B0(
        \i_MIPS/Register/register[29][5] ), .B1(n4841), .Y(n7305) );
  AO22X1 U5624 ( .A0(n5002), .A1(n650), .B0(n4998), .B1(n2173), .Y(n9200) );
  AO22X1 U5625 ( .A0(n5002), .A1(n651), .B0(n4998), .B1(n2174), .Y(n9191) );
  AO22X1 U5626 ( .A0(n5002), .A1(n485), .B0(n4998), .B1(n2052), .Y(n9072) );
  AO22X1 U5627 ( .A0(n5002), .A1(n559), .B0(n4998), .B1(n2062), .Y(n9063) );
  AO22X1 U5628 ( .A0(n5002), .A1(n560), .B0(n4998), .B1(n2063), .Y(n8985) );
  AO22X1 U5629 ( .A0(n5002), .A1(n652), .B0(n4998), .B1(n2175), .Y(n8701) );
  AO22X1 U5630 ( .A0(n5002), .A1(n653), .B0(n4998), .B1(n2176), .Y(n8790) );
  AO22X1 U5631 ( .A0(n5002), .A1(n561), .B0(n4998), .B1(n2064), .Y(n8976) );
  AO22X1 U5632 ( .A0(n5002), .A1(n654), .B0(n4998), .B1(n2177), .Y(n8692) );
  AO22X1 U5633 ( .A0(n5002), .A1(n562), .B0(n4998), .B1(n2065), .Y(n8781) );
  AO22X1 U5634 ( .A0(n5002), .A1(n655), .B0(n4997), .B1(n2178), .Y(n7343) );
  AO22X1 U5635 ( .A0(n5002), .A1(n656), .B0(n4997), .B1(n2179), .Y(n7334) );
  OA22X1 U5636 ( .A0(n5344), .A1(n998), .B0(n5300), .B1(n2550), .Y(n9749) );
  OA22X1 U5637 ( .A0(n5345), .A1(n2508), .B0(n5301), .B1(n748), .Y(n9771) );
  OA22X1 U5638 ( .A0(net112045), .A1(n2808), .B0(net111921), .B1(n806), .Y(
        n6710) );
  AO21XL U5639 ( .A0(\i_MIPS/ID_EX[95] ), .A1(n5517), .B0(n4499), .Y(
        \i_MIPS/n490 ) );
  AO21XL U5640 ( .A0(\i_MIPS/ID_EX[100] ), .A1(n5517), .B0(n4499), .Y(
        \i_MIPS/n485 ) );
  AO21XL U5641 ( .A0(\i_MIPS/ID_EX[101] ), .A1(n5518), .B0(n4499), .Y(
        \i_MIPS/n484 ) );
  AO21XL U5642 ( .A0(\i_MIPS/ID_EX[104] ), .A1(n5513), .B0(n4499), .Y(
        \i_MIPS/n481 ) );
  OA22XL U5643 ( .A0(net112053), .A1(n1490), .B0(net111929), .B1(n3103), .Y(
        n7153) );
  OA22XL U5644 ( .A0(net112045), .A1(n1491), .B0(net111921), .B1(n3104), .Y(
        n6718) );
  OA22XL U5645 ( .A0(n5338), .A1(n2551), .B0(n5294), .B1(n780), .Y(n9470) );
  OA22XL U5646 ( .A0(n5340), .A1(n1083), .B0(n5296), .B1(n2655), .Y(n9524) );
  OA22XL U5647 ( .A0(n5335), .A1(n1084), .B0(n5291), .B1(n2656), .Y(n9384) );
  OA22XL U5648 ( .A0(n5336), .A1(n1085), .B0(n5292), .B1(n2657), .Y(n9423) );
  OA22XL U5649 ( .A0(n5350), .A1(n1086), .B0(n5306), .B1(n2658), .Y(n9966) );
  OA22XL U5650 ( .A0(net112079), .A1(n1492), .B0(net111955), .B1(n3105), .Y(
        n9048) );
  OA22XL U5651 ( .A0(net112079), .A1(n1493), .B0(net111955), .B1(n3106), .Y(
        n8969) );
  OA22XL U5652 ( .A0(net112045), .A1(n2858), .B0(net111921), .B1(n849), .Y(
        n6539) );
  OA22XL U5653 ( .A0(net112055), .A1(n1494), .B0(net111931), .B1(n3107), .Y(
        n7397) );
  MX2XL U5654 ( .A(n3791), .B(net100015), .S0(n5510), .Y(\i_MIPS/n425 ) );
  MX2XL U5655 ( .A(\i_MIPS/ID_EX[50] ), .B(net99056), .S0(n5510), .Y(
        \i_MIPS/n419 ) );
  CLKINVX3 U5656 ( .A(n5304), .Y(n5279) );
  CLKINVX3 U5657 ( .A(n5307), .Y(n5281) );
  CLKINVX3 U5658 ( .A(n5348), .Y(n5324) );
  CLKINVX3 U5659 ( .A(n5382), .Y(n5366) );
  CLKINVX3 U5660 ( .A(n5287), .Y(n5282) );
  CLKINVX3 U5661 ( .A(n5328), .Y(n5327) );
  CLKINVX3 U5662 ( .A(n5377), .Y(n5373) );
  CLKINVX3 U5663 ( .A(n5304), .Y(n5283) );
  CLKINVX3 U5664 ( .A(n5304), .Y(n5284) );
  CLKINVX3 U5665 ( .A(n5288), .Y(n5280) );
  CLKINVX3 U5666 ( .A(n5426), .Y(n5410) );
  CLKINVX3 U5667 ( .A(n5304), .Y(n5278) );
  CLKINVX3 U5668 ( .A(n5307), .Y(n5277) );
  CLKINVX3 U5669 ( .A(n5286), .Y(n5285) );
  CLKINVX2 U5670 ( .A(net112555), .Y(net112527) );
  CLKINVX2 U5671 ( .A(net112147), .Y(net112115) );
  CLKINVX2 U5672 ( .A(net112657), .Y(net112637) );
  CLKINVX2 U5673 ( .A(net112555), .Y(net112535) );
  CLKINVX2 U5674 ( .A(net112151), .Y(net112125) );
  CLKINVX2 U5675 ( .A(net112555), .Y(net112537) );
  CLKINVX2 U5676 ( .A(net112655), .Y(net112639) );
  CLKINVX2 U5677 ( .A(net112681), .Y(net112629) );
  CLKINVX2 U5678 ( .A(net112341), .Y(net112285) );
  CLKINVX2 U5679 ( .A(net112473), .Y(net112409) );
  CLKINVX2 U5680 ( .A(net112555), .Y(net112533) );
  CLKINVX2 U5681 ( .A(net112657), .Y(net112635) );
  CLKINVX2 U5682 ( .A(net112145), .Y(net112119) );
  CLKINVX2 U5683 ( .A(net112555), .Y(net112531) );
  CLKINVX2 U5684 ( .A(net112659), .Y(net112633) );
  CLKINVX2 U5685 ( .A(net112147), .Y(net112113) );
  CLKINVX2 U5686 ( .A(net112555), .Y(net112525) );
  CLKINVX2 U5687 ( .A(net112673), .Y(net112627) );
  CLKINVX2 U5688 ( .A(net112155), .Y(net112127) );
  CLKINVX2 U5689 ( .A(net112575), .Y(net112539) );
  CLKINVX2 U5690 ( .A(net112655), .Y(net112641) );
  CLKINVX2 U5691 ( .A(net112573), .Y(net112545) );
  CLKINVX2 U5692 ( .A(net112651), .Y(net112647) );
  CLKINVX2 U5693 ( .A(net112145), .Y(net112117) );
  CLKINVX2 U5694 ( .A(net112555), .Y(net112529) );
  CLKINVX2 U5695 ( .A(net112659), .Y(net112631) );
  CLKINVX2 U5696 ( .A(net112139), .Y(net112129) );
  CLKINVX2 U5697 ( .A(net112139), .Y(net112131) );
  CLKINVX2 U5698 ( .A(net112569), .Y(net112543) );
  CLKINVX2 U5699 ( .A(net112671), .Y(net112645) );
  CLKINVX2 U5700 ( .A(net112061), .Y(net112011) );
  CLKINVX2 U5701 ( .A(net112425), .Y(net112423) );
  CLKINVX2 U5702 ( .A(net112583), .Y(net112547) );
  CLKINVX2 U5703 ( .A(net112651), .Y(net112649) );
  BUFX2 U5704 ( .A(n5449), .Y(n5427) );
  CLKBUFX2 U5705 ( .A(n5143), .Y(n5118) );
  CLKBUFX2 U5706 ( .A(n5143), .Y(n5117) );
  BUFX8 U5707 ( .A(n4969), .Y(n4974) );
  BUFX8 U5708 ( .A(n4983), .Y(n4987) );
  INVXL U5709 ( .A(n10378), .Y(n10347) );
  CLKBUFX2 U5710 ( .A(n154), .Y(n5518) );
  CLKBUFX2 U5711 ( .A(n5143), .Y(n5121) );
  CLKBUFX2 U5712 ( .A(n5429), .Y(n5430) );
  CLKBUFX2 U5713 ( .A(n5403), .Y(n5386) );
  CLKBUFX2 U5714 ( .A(net112507), .Y(net112455) );
  CLKBUFX2 U5715 ( .A(n3611), .Y(n5434) );
  CLKBUFX2 U5716 ( .A(n4983), .Y(n4988) );
  CLKBUFX2 U5717 ( .A(n3611), .Y(n5436) );
  CLKBUFX2 U5718 ( .A(n5141), .Y(n5128) );
  CLKBUFX2 U5719 ( .A(n5402), .Y(n5391) );
  INVX3 U5720 ( .A(n7544), .Y(n7111) );
  INVX3 U5721 ( .A(n10918), .Y(n10921) );
  CLKBUFX2 U5722 ( .A(n5143), .Y(n5140) );
  CLKBUFX2 U5723 ( .A(n5409), .Y(n5401) );
  CLKBUFX2 U5724 ( .A(n5365), .Y(n5360) );
  CLKBUFX2 U5725 ( .A(n5144), .Y(n5186) );
  CLKBUFX2 U5726 ( .A(n5275), .Y(n5273) );
  CLKBUFX2 U5727 ( .A(n5188), .Y(n5185) );
  CLKBUFX2 U5728 ( .A(n5365), .Y(n5359) );
  CLKBUFX2 U5729 ( .A(n5318), .Y(n5314) );
  CLKBUFX2 U5730 ( .A(n5163), .Y(n5184) );
  CLKBUFX2 U5731 ( .A(n5363), .Y(n5358) );
  CLKBUFX2 U5732 ( .A(n5229), .Y(n5226) );
  CLKBUFX2 U5733 ( .A(n5275), .Y(n5271) );
  OR2XL U5734 ( .A(net113725), .B(n10777), .Y(n4773) );
  OR2XL U5735 ( .A(net113725), .B(n10608), .Y(n4776) );
  OR2XL U5736 ( .A(net113725), .B(n10569), .Y(n4780) );
  OR2XL U5737 ( .A(net113667), .B(n10411), .Y(n4782) );
  NAND2BXL U5738 ( .AN(n3819), .B(n11182), .Y(n11189) );
  CLKBUFX2 U5739 ( .A(n3611), .Y(n5447) );
  CLKBUFX2 U5740 ( .A(n5143), .Y(n5139) );
  CLKBUFX2 U5741 ( .A(n5290), .Y(n5312) );
  CLKBUFX2 U5742 ( .A(n5228), .Y(n5224) );
  CLKBUFX2 U5743 ( .A(n5330), .Y(n5356) );
  CLKBUFX2 U5744 ( .A(n5274), .Y(n5270) );
  INVX1 U5745 ( .A(n10356), .Y(n10357) );
  AOI2BB1XL U5746 ( .A0N(n10500), .A1N(n168), .B0(n4595), .Y(n10501) );
  AO22XL U5747 ( .A0(net113455), .A1(n11421), .B0(net113461), .B1(n11390), .Y(
        n6544) );
  AO22XL U5748 ( .A0(net113445), .A1(n11469), .B0(net102346), .B1(n11500), .Y(
        n7928) );
  INVX1 U5749 ( .A(n8082), .Y(n8076) );
  NAND2X2 U5750 ( .A(n8426), .B(n8351), .Y(n6593) );
  AND2X2 U5751 ( .A(n7111), .B(n8666), .Y(n7113) );
  AO22X4 U5752 ( .A0(n8807), .A1(n9259), .B0(n9258), .B1(n8806), .Y(n8809) );
  OAI211X2 U5753 ( .A0(n6469), .A1(n6477), .B0(n6468), .C0(n6467), .Y(n6478)
         );
  INVXL U5754 ( .A(n8088), .Y(n8090) );
  NAND2X2 U5755 ( .A(n4778), .B(n4589), .Y(n10157) );
  NAND2XL U5756 ( .A(n11224), .B(n9150), .Y(n9152) );
  NAND2XL U5757 ( .A(n9141), .B(n9143), .Y(n9147) );
  INVX3 U5758 ( .A(n10214), .Y(n10216) );
  NAND2X2 U5759 ( .A(n5590), .B(n4707), .Y(n7867) );
  INVX1 U5760 ( .A(n8344), .Y(n8360) );
  INVX1 U5761 ( .A(n8282), .Y(n8273) );
  INVX1 U5762 ( .A(n8162), .Y(n8157) );
  AO22XL U5763 ( .A0(n4800), .A1(n8530), .B0(n8529), .B1(n3636), .Y(n8552) );
  AO22XL U5764 ( .A0(n4800), .A1(n7964), .B0(n8254), .B1(n3636), .Y(n7978) );
  INVXL U5765 ( .A(n6477), .Y(n6479) );
  INVXL U5766 ( .A(n8338), .Y(n8341) );
  OA22X4 U5767 ( .A0(n9946), .A1(n5454), .B0(n9945), .B1(n5461), .Y(n9947) );
  INVX3 U5768 ( .A(n6512), .Y(n9310) );
  CLKMX2X4 U5769 ( .A(n8265), .B(n7474), .S0(n5590), .Y(n7787) );
  INVXL U5770 ( .A(n7951), .Y(n7953) );
  INVXL U5771 ( .A(n8542), .Y(n8547) );
  NAND2BXL U5772 ( .AN(n5461), .B(n11280), .Y(n10047) );
  NAND2BXL U5773 ( .AN(n5461), .B(n11279), .Y(n11147) );
  NAND2BXL U5774 ( .AN(n5456), .B(n11247), .Y(n11148) );
  NAND2BXL U5775 ( .AN(n5461), .B(n11282), .Y(n10023) );
  NAND2BXL U5776 ( .AN(n5461), .B(n11278), .Y(n10076) );
  NAND2BXL U5777 ( .AN(n5461), .B(n11281), .Y(n9994) );
  NAND2BXL U5778 ( .AN(n5461), .B(n11286), .Y(n9903) );
  NAND2BXL U5779 ( .AN(n5456), .B(n11254), .Y(n9904) );
  NAND2BXL U5780 ( .AN(n5461), .B(n11287), .Y(n10125) );
  NAND2BXL U5781 ( .AN(n5461), .B(n11283), .Y(n9879) );
  NAND2BXL U5782 ( .AN(n5456), .B(n11251), .Y(n9880) );
  NAND2BXL U5783 ( .AN(n5461), .B(n11285), .Y(n9927) );
  NAND2BXL U5784 ( .AN(n5461), .B(n11284), .Y(net100751) );
  NAND2BXL U5785 ( .AN(n5456), .B(n11252), .Y(net100750) );
  INVX3 U5786 ( .A(n11068), .Y(n11065) );
  XOR3XL U5787 ( .A(n11043), .B(n11003), .C(n11042), .Y(n11000) );
  NAND2BXL U5788 ( .AN(n5456), .B(n11257), .Y(n9737) );
  INVXL U5789 ( .A(n6764), .Y(n6766) );
  NAND2BXL U5790 ( .AN(n5456), .B(n11261), .Y(n9757) );
  NAND2BXL U5791 ( .AN(n5456), .B(n11260), .Y(n9805) );
  NAND2BXL U5792 ( .AN(n5456), .B(n11258), .Y(n9781) );
  INVXL U5793 ( .A(n7622), .Y(n7620) );
  INVX1 U5794 ( .A(n11326), .Y(n9609) );
  INVX1 U5795 ( .A(n7980), .Y(n7983) );
  INVX1 U5796 ( .A(n7884), .Y(n7887) );
  INVX1 U5797 ( .A(n8079), .Y(n8077) );
  AND2XL U5798 ( .A(n3218), .B(net100035), .Y(n4529) );
  AND3XL U5799 ( .A(net99476), .B(net99475), .C(net99477), .Y(n4524) );
  AND2XL U5800 ( .A(net99386), .B(net99387), .Y(n4528) );
  AND2XL U5801 ( .A(net99363), .B(net99364), .Y(n4557) );
  AND3XL U5802 ( .A(net98966), .B(net98964), .C(net98965), .Y(n4546) );
  AND2XL U5803 ( .A(net99711), .B(net99712), .Y(n4531) );
  AND2XL U5804 ( .A(n3312), .B(net99634), .Y(n4534) );
  CLKBUFX2 U5805 ( .A(n4619), .Y(n4861) );
  CLKBUFX2 U5806 ( .A(n4619), .Y(n4862) );
  CLKBUFX2 U5807 ( .A(n4619), .Y(n4863) );
  INVX1 U5808 ( .A(n7555), .Y(n7565) );
  CLKBUFX2 U5809 ( .A(n4623), .Y(n4853) );
  CLKBUFX2 U5810 ( .A(n4622), .Y(n4839) );
  CLKBUFX2 U5811 ( .A(n4623), .Y(n4854) );
  CLKBUFX2 U5812 ( .A(n4622), .Y(n4840) );
  INVXL U5813 ( .A(n9269), .Y(n9270) );
  BUFX4 U5814 ( .A(n4619), .Y(n4859) );
  NAND2XL U5815 ( .A(n4693), .B(n11262), .Y(n11182) );
  INVXL U5816 ( .A(n11435), .Y(n10195) );
  INVXL U5817 ( .A(n11434), .Y(n10444) );
  INVXL U5818 ( .A(n11433), .Y(n10810) );
  INVXL U5819 ( .A(n11499), .Y(n10595) );
  INVXL U5820 ( .A(n11509), .Y(n10462) );
  INVXL U5821 ( .A(n11508), .Y(n10411) );
  INVXL U5822 ( .A(n11506), .Y(n10569) );
  INVXL U5823 ( .A(n11502), .Y(n10520) );
  INVXL U5824 ( .A(n11498), .Y(n10449) );
  INVXL U5825 ( .A(n11497), .Y(n10186) );
  INVXL U5826 ( .A(n11496), .Y(n10435) );
  INVXL U5827 ( .A(n11491), .Y(n10765) );
  INVXL U5828 ( .A(n11490), .Y(n10817) );
  AO21X4 U5829 ( .A0(n10271), .A1(n10270), .B0(n10269), .Y(n10303) );
  OA22X4 U5830 ( .A0(n5425), .A1(n1601), .B0(n5381), .B1(n3265), .Y(n5973) );
  OA22X4 U5831 ( .A0(n5160), .A1(n3226), .B0(n5118), .B1(n1587), .Y(n5976) );
  OA22X4 U5832 ( .A0(n5243), .A1(n3227), .B0(n5229), .B1(n1588), .Y(n5975) );
  OA22X4 U5833 ( .A0(n5424), .A1(n425), .B0(n5380), .B1(n3266), .Y(n5969) );
  OA22X4 U5834 ( .A0(n5160), .A1(n1968), .B0(n5117), .B1(n396), .Y(n5972) );
  OA22X4 U5835 ( .A0(n5243), .A1(n1969), .B0(n5204), .B1(n397), .Y(n5971) );
  OA22X4 U5836 ( .A0(n5250), .A1(n3229), .B0(n5230), .B1(n400), .Y(n5963) );
  AOI211XL U5837 ( .A0(n8801), .A1(n177), .B0(n4672), .C0(n4667), .Y(n8815) );
  OA22X4 U5838 ( .A0(n5422), .A1(n1602), .B0(n5383), .B1(n3267), .Y(n5957) );
  OA22X4 U5839 ( .A0(n5156), .A1(n3230), .B0(n5115), .B1(n1589), .Y(n5960) );
  OA22X4 U5840 ( .A0(n5246), .A1(n3231), .B0(n5230), .B1(n1590), .Y(n5959) );
  OAI211X2 U5841 ( .A0(n7287), .A1(n3529), .B0(n7550), .C0(n7459), .Y(n6768)
         );
  NAND2X2 U5842 ( .A(n6242), .B(\i_MIPS/n364 ), .Y(n7477) );
  NAND2X4 U5843 ( .A(n6587), .B(\i_MIPS/n345 ), .Y(n8351) );
  INVXL U5844 ( .A(n8718), .Y(n8723) );
  AO21X4 U5845 ( .A0(n10878), .A1(n10877), .B0(n4611), .Y(n10314) );
  NAND2X2 U5846 ( .A(n8922), .B(n8925), .Y(n6590) );
  NAND2X2 U5847 ( .A(n11089), .B(n11088), .Y(n10264) );
  OA22X4 U5848 ( .A0(n5155), .A1(n3281), .B0(n5112), .B1(n1591), .Y(n4453) );
  OA22X4 U5849 ( .A0(n5244), .A1(n3282), .B0(n5203), .B1(n1592), .Y(n4454) );
  OA22X4 U5850 ( .A0(n5161), .A1(n3283), .B0(n5142), .B1(n1593), .Y(n4455) );
  OA22X4 U5851 ( .A0(n5248), .A1(n3284), .B0(n5202), .B1(n1594), .Y(n4456) );
  OA22X4 U5852 ( .A0(n5159), .A1(n3232), .B0(n5116), .B1(n1595), .Y(n4457) );
  OA22X4 U5853 ( .A0(n5245), .A1(n3233), .B0(n5200), .B1(n1596), .Y(n4458) );
  OA22X4 U5854 ( .A0(n5161), .A1(n1971), .B0(n5141), .B1(n401), .Y(n4459) );
  OA22X4 U5855 ( .A0(n5243), .A1(n426), .B0(n5228), .B1(n3268), .Y(n4460) );
  OA22X4 U5856 ( .A0(n5155), .A1(n1972), .B0(n5114), .B1(n402), .Y(n4461) );
  OA22X4 U5857 ( .A0(n5245), .A1(n1973), .B0(n5204), .B1(n403), .Y(n4462) );
  OA22X4 U5858 ( .A0(n5164), .A1(n3234), .B0(n5113), .B1(n404), .Y(n4463) );
  OA22X4 U5859 ( .A0(n5244), .A1(n3307), .B0(n5201), .B1(n405), .Y(n4464) );
  OA22X4 U5860 ( .A0(n5158), .A1(n1603), .B0(n5116), .B1(n3305), .Y(n4468) );
  OA22X4 U5861 ( .A0(n5247), .A1(n1604), .B0(n5228), .B1(n3306), .Y(n4469) );
  AO21X4 U5862 ( .A0(n10930), .A1(n10929), .B0(n10919), .Y(n11104) );
  AO22X4 U5863 ( .A0(net99583), .A1(net113041), .B0(net102300), .B1(n6998), 
        .Y(net106078) );
  AO22X4 U5864 ( .A0(net113041), .A1(net99110), .B0(net102300), .B1(n7522), 
        .Y(net105120) );
  OA22X4 U5865 ( .A0(n5186), .A1(n3298), .B0(n5115), .B1(n1633), .Y(n4472) );
  OA22X4 U5866 ( .A0(n5243), .A1(n3299), .B0(n5200), .B1(n1634), .Y(n4473) );
  OA22X4 U5867 ( .A0(n5429), .A1(n3300), .B0(n5384), .B1(n1635), .Y(n4474) );
  AND2XL U5868 ( .A(n9260), .B(n9277), .Y(n9294) );
  NAND4X2 U5869 ( .A(n9516), .B(n9515), .C(n9514), .D(n9513), .Y(n11233) );
  NAND2X2 U5870 ( .A(n10151), .B(n11168), .Y(n11515) );
  NAND4X2 U5871 ( .A(n9649), .B(n9648), .C(n9647), .D(n9646), .Y(n11239) );
  NAND4X2 U5872 ( .A(n9639), .B(n9638), .C(n9637), .D(n9636), .Y(n11271) );
  OA22XL U5873 ( .A0(n5435), .A1(n1087), .B0(n5402), .B1(n2659), .Y(n9636) );
  OA22XL U5874 ( .A0(n5171), .A1(n1088), .B0(n5134), .B1(n2660), .Y(n9639) );
  OA22XL U5875 ( .A0(n5257), .A1(n1089), .B0(n5211), .B1(n2661), .Y(n9638) );
  NAND4X2 U5876 ( .A(n9634), .B(n9633), .C(n9632), .D(n9631), .Y(n11303) );
  OA22XL U5877 ( .A0(n5435), .A1(n2803), .B0(n5396), .B1(n1223), .Y(n9631) );
  OA22XL U5878 ( .A0(n5171), .A1(n1090), .B0(n5123), .B1(n2662), .Y(n9634) );
  OA22XL U5879 ( .A0(n5257), .A1(n1091), .B0(n5211), .B1(n2663), .Y(n9633) );
  NAND4X2 U5880 ( .A(n9386), .B(n9385), .C(n9384), .D(n9383), .Y(n11275) );
  OA22XL U5881 ( .A0(n5430), .A1(n1092), .B0(n5386), .B1(n2664), .Y(n9383) );
  NAND4X2 U5882 ( .A(n9376), .B(n9375), .C(n9374), .D(n9373), .Y(n11307) );
  OA22XL U5883 ( .A0(n5165), .A1(n1093), .B0(n5121), .B1(n2665), .Y(n9376) );
  OA22XL U5884 ( .A0(n5251), .A1(n1094), .B0(n5205), .B1(n2666), .Y(n9375) );
  OA22XL U5885 ( .A0(n5430), .A1(n1095), .B0(n5386), .B1(n2667), .Y(n9373) );
  NAND4X2 U5886 ( .A(n9819), .B(n9818), .C(n9817), .D(n9816), .Y(n11269) );
  OA22XL U5887 ( .A0(n5436), .A1(n1096), .B0(n5388), .B1(n2668), .Y(n9816) );
  OA22XL U5888 ( .A0(n5176), .A1(n1097), .B0(n5131), .B1(n2669), .Y(n9819) );
  NAND4BX2 U5889 ( .AN(n4475), .B(n9449), .C(n9448), .D(n9447), .Y(n11268) );
  NAND4X2 U5890 ( .A(n9644), .B(n9643), .C(n9642), .D(n9641), .Y(n11335) );
  OA22XL U5891 ( .A0(n5432), .A1(n1098), .B0(n5388), .B1(n2670), .Y(n9442) );
  OA22XL U5892 ( .A0(n5167), .A1(n1099), .B0(n5123), .B1(n2671), .Y(n9445) );
  OA22XL U5893 ( .A0(n5253), .A1(n1100), .B0(n5207), .B1(n2672), .Y(n9444) );
  NAND4BX2 U5894 ( .AN(n4476), .B(n9672), .C(n9671), .D(n9670), .Y(n11272) );
  NAND4X2 U5895 ( .A(n9668), .B(n9667), .C(n9666), .D(n9665), .Y(n11240) );
  NAND4BX2 U5896 ( .AN(n4477), .B(n9471), .C(n9470), .D(n9469), .Y(n11266) );
  NAND4X2 U5897 ( .A(n9467), .B(n9466), .C(n9465), .D(n9464), .Y(n11298) );
  OA22XL U5898 ( .A0(n5433), .A1(n2552), .B0(n5396), .B1(n781), .Y(n9464) );
  OA22XL U5899 ( .A0(n5168), .A1(n1101), .B0(n5124), .B1(n2673), .Y(n9467) );
  OA22XL U5900 ( .A0(n5254), .A1(n2553), .B0(n5208), .B1(n782), .Y(n9466) );
  OA22XL U5901 ( .A0(n5432), .A1(n1102), .B0(n5388), .B1(n2674), .Y(n9437) );
  OA22XL U5902 ( .A0(n5167), .A1(n1103), .B0(n5123), .B1(n2675), .Y(n9440) );
  OA22XL U5903 ( .A0(n5253), .A1(n1104), .B0(n5207), .B1(n2676), .Y(n9439) );
  NAND4BX2 U5904 ( .AN(n4478), .B(n9415), .C(n9414), .D(n9413), .Y(n11270) );
  NAND4X2 U5905 ( .A(n9824), .B(n9823), .C(n9822), .D(n9821), .Y(n11333) );
  OA22XL U5906 ( .A0(n5432), .A1(n2554), .B0(n5388), .B1(n783), .Y(n9454) );
  OA22XL U5907 ( .A0(n5167), .A1(n1105), .B0(n5123), .B1(n2677), .Y(n9457) );
  OA22XL U5908 ( .A0(n5253), .A1(n1106), .B0(n5207), .B1(n2678), .Y(n9456) );
  OA22XL U5909 ( .A0(n5166), .A1(n1107), .B0(n5122), .B1(n2679), .Y(n9420) );
  OA22XL U5910 ( .A0(n5252), .A1(n1108), .B0(n5206), .B1(n2680), .Y(n9419) );
  OA22XL U5911 ( .A0(n5431), .A1(n1109), .B0(n5387), .B1(n2681), .Y(n9417) );
  OA22XL U5912 ( .A0(n5166), .A1(n1110), .B0(n5122), .B1(n2682), .Y(n9411) );
  OA22XL U5913 ( .A0(n5252), .A1(n1111), .B0(n5206), .B1(n2683), .Y(n9410) );
  OA22XL U5914 ( .A0(n5431), .A1(n1112), .B0(n5387), .B1(n2684), .Y(n9408) );
  OA22XL U5915 ( .A0(n5166), .A1(n1113), .B0(n5122), .B1(n2685), .Y(n9425) );
  OA22XL U5916 ( .A0(n5252), .A1(n1114), .B0(n5206), .B1(n2686), .Y(n9424) );
  OA22XL U5917 ( .A0(n5431), .A1(n2555), .B0(n5387), .B1(n784), .Y(n9422) );
  OA22XL U5918 ( .A0(n5432), .A1(n2556), .B0(n5388), .B1(n785), .Y(n9459) );
  OA22XL U5919 ( .A0(n5167), .A1(n1115), .B0(n5123), .B1(n2687), .Y(n9462) );
  OA22XL U5920 ( .A0(n5253), .A1(n1116), .B0(n5207), .B1(n2688), .Y(n9461) );
  NAND4X2 U5921 ( .A(n9936), .B(n9935), .C(n9934), .D(n9933), .Y(n11245) );
  NAND4X2 U5922 ( .A(n9350), .B(n9349), .C(n9348), .D(n9347), .Y(n11341) );
  OA22XL U5923 ( .A0(n5429), .A1(n1495), .B0(n5385), .B1(n3108), .Y(n9347) );
  OA22XL U5924 ( .A0(n5250), .A1(n1496), .B0(n5205), .B1(n3109), .Y(n9349) );
  NAND4X2 U5925 ( .A(n9944), .B(n9943), .C(n9942), .D(n9941), .Y(n11277) );
  NAND4X2 U5926 ( .A(n9940), .B(n9939), .C(n9938), .D(n9937), .Y(n11309) );
  OA22XL U5927 ( .A0(net112241), .A1(n807), .B0(net112159), .B1(n2340), .Y(
        n9250) );
  OA22XL U5928 ( .A0(net112083), .A1(n808), .B0(net111959), .B1(n2341), .Y(
        n9245) );
  OA22XL U5929 ( .A0(net112493), .A1(n809), .B0(net112353), .B1(n2342), .Y(
        n9247) );
  OA22XL U5930 ( .A0(net112241), .A1(n810), .B0(net112159), .B1(n2343), .Y(
        n9246) );
  OA22XL U5931 ( .A0(net112083), .A1(n811), .B0(net111959), .B1(n2344), .Y(
        n9237) );
  OA22XL U5932 ( .A0(net112459), .A1(n812), .B0(net112353), .B1(n2345), .Y(
        n9239) );
  OA22XL U5933 ( .A0(net112239), .A1(n813), .B0(net112161), .B1(n2346), .Y(
        n9238) );
  OA22XL U5934 ( .A0(net112465), .A1(n1497), .B0(net112341), .B1(n3110), .Y(
        n7155) );
  INVX1 U5935 ( .A(n9162), .Y(n9145) );
  INVX1 U5936 ( .A(n9161), .Y(n9144) );
  INVXL U5937 ( .A(n7107), .Y(n7109) );
  NAND2XL U5938 ( .A(n8897), .B(n8250), .Y(n6492) );
  NAND4XL U5939 ( .A(n6661), .B(n6660), .C(n3727), .D(n9160), .Y(n6676) );
  AO22XL U5940 ( .A0(n4978), .A1(n248), .B0(n4976), .B1(n307), .Y(n7602) );
  AO22XL U5941 ( .A0(n4978), .A1(n293), .B0(n4976), .B1(n1873), .Y(n7593) );
  AO22XL U5942 ( .A0(n4978), .A1(n527), .B0(n4976), .B1(n2282), .Y(n7535) );
  AO22XL U5943 ( .A0(n4978), .A1(n528), .B0(n4976), .B1(n2283), .Y(n7526) );
  AO22XL U5944 ( .A0(n4979), .A1(n529), .B0(n4976), .B1(n2284), .Y(n8132) );
  AO22XL U5945 ( .A0(n4979), .A1(n530), .B0(n9309), .B1(n2285), .Y(n8123) );
  AO22XL U5946 ( .A0(n4977), .A1(n531), .B0(n4976), .B1(n2286), .Y(n7443) );
  AO22XL U5947 ( .A0(n4977), .A1(n532), .B0(n4976), .B1(n2287), .Y(n7434) );
  AO22XL U5948 ( .A0(n4978), .A1(n533), .B0(n9309), .B1(n2288), .Y(n7942) );
  AO22XL U5949 ( .A0(n4978), .A1(n534), .B0(n9309), .B1(n2289), .Y(n7933) );
  AO22XL U5950 ( .A0(n4978), .A1(n494), .B0(n4976), .B1(n2246), .Y(n7685) );
  AO22XL U5951 ( .A0(n4978), .A1(n495), .B0(n9309), .B1(n2247), .Y(n7676) );
  AO22XL U5952 ( .A0(n4978), .A1(n535), .B0(n9309), .B1(n2290), .Y(n6186) );
  AO22XL U5953 ( .A0(n4978), .A1(n536), .B0(n9309), .B1(n2291), .Y(n6177) );
  AO22XL U5954 ( .A0(n4978), .A1(n496), .B0(n9309), .B1(n2248), .Y(n6827) );
  AO22XL U5955 ( .A0(n4978), .A1(n498), .B0(n9309), .B1(n2250), .Y(n6910) );
  AO22XL U5956 ( .A0(n4978), .A1(n499), .B0(n4976), .B1(n2251), .Y(n6756) );
  AO22XL U5957 ( .A0(n4977), .A1(n500), .B0(n4976), .B1(n2252), .Y(n6747) );
  AO22XL U5958 ( .A0(n4977), .A1(n537), .B0(n4976), .B1(n2292), .Y(n7011) );
  AO22XL U5959 ( .A0(n4977), .A1(n538), .B0(n4976), .B1(n2293), .Y(n7002) );
  AO22XL U5960 ( .A0(n4979), .A1(n501), .B0(n9309), .B1(n2253), .Y(n8318) );
  AO22XL U5961 ( .A0(n4979), .A1(n502), .B0(n9309), .B1(n2254), .Y(n8309) );
  AO22XL U5962 ( .A0(n4980), .A1(n539), .B0(n9309), .B1(n2294), .Y(n8987) );
  AO22XL U5963 ( .A0(n9310), .A1(n540), .B0(n9309), .B1(n2295), .Y(n8978) );
  AO22XL U5964 ( .A0(n4980), .A1(n503), .B0(n9309), .B1(n2255), .Y(n8792) );
  AO22XL U5965 ( .A0(n4977), .A1(n504), .B0(n9309), .B1(n2256), .Y(n8783) );
  AO22XL U5966 ( .A0(n4979), .A1(n505), .B0(n9309), .B1(n2257), .Y(n8221) );
  AO22XL U5967 ( .A0(n4977), .A1(n506), .B0(n9309), .B1(n2258), .Y(n7261) );
  AO22XL U5968 ( .A0(n4977), .A1(n507), .B0(n9309), .B1(n2259), .Y(n7252) );
  AO22XL U5969 ( .A0(n4979), .A1(n508), .B0(n9309), .B1(n2260), .Y(n8212) );
  AO22XL U5970 ( .A0(n4978), .A1(n295), .B0(n4976), .B1(n1867), .Y(n7838) );
  AO22XL U5971 ( .A0(n4977), .A1(n509), .B0(n4976), .B1(n2261), .Y(n7162) );
  AO22XL U5972 ( .A0(n4977), .A1(n542), .B0(n9309), .B1(n2297), .Y(n7336) );
  INVX3 U5973 ( .A(n10969), .Y(n10965) );
  INVXL U5974 ( .A(n3796), .Y(n6459) );
  NAND2XL U5975 ( .A(n8144), .B(n7704), .Y(n7706) );
  NAND2X1 U5976 ( .A(n4500), .B(n4581), .Y(n4481) );
  INVXL U5977 ( .A(n8888), .Y(n8908) );
  INVXL U5978 ( .A(n8642), .Y(n8654) );
  MX2XL U5979 ( .A(n9280), .B(n9279), .S0(n7620), .Y(n7631) );
  INVXL U5980 ( .A(n7099), .Y(n6466) );
  INVX3 U5981 ( .A(net99753), .Y(net99737) );
  CLKBUFX20 U5982 ( .A(n11545), .Y(mem_read_D) );
  OA21XL U5983 ( .A0(n9164), .A1(n9163), .B0(n9170), .Y(n9178) );
  NAND4X2 U5984 ( .A(n7927), .B(n7926), .C(n7925), .D(n7924), .Y(n11500) );
  OA22XL U5985 ( .A0(net112233), .A1(n1498), .B0(net112151), .B1(n3111), .Y(
        n7925) );
  NAND4X2 U5986 ( .A(n9814), .B(n9813), .C(n9812), .D(n9811), .Y(n11301) );
  OA22XL U5987 ( .A0(n5436), .A1(n1117), .B0(n5398), .B1(n2689), .Y(n9811) );
  OA22XL U5988 ( .A0(n5176), .A1(n1118), .B0(n5131), .B1(n2690), .Y(n9814) );
  OA22XL U5989 ( .A0(n5262), .A1(n1119), .B0(n5216), .B1(n2691), .Y(n9813) );
  OAI2BB1X4 U5990 ( .A0N(n9277), .A1N(n9179), .B0(n9260), .Y(n9184) );
  NAND4X2 U5991 ( .A(n9491), .B(n9490), .C(n9489), .D(n9488), .Y(n11264) );
  OA22XL U5992 ( .A0(n5433), .A1(n1120), .B0(n5387), .B1(n2692), .Y(n9488) );
  OA22XL U5993 ( .A0(n5168), .A1(n1121), .B0(n5124), .B1(n2693), .Y(n9491) );
  OA22XL U5994 ( .A0(n5254), .A1(n1122), .B0(n5208), .B1(n2694), .Y(n9490) );
  NAND4X2 U5995 ( .A(n9486), .B(n9485), .C(n9484), .D(n9483), .Y(n11296) );
  OA22XL U5996 ( .A0(n5433), .A1(n1123), .B0(n5387), .B1(n2695), .Y(n9483) );
  OA22XL U5997 ( .A0(n5168), .A1(n1124), .B0(n5124), .B1(n2696), .Y(n9486) );
  OA22XL U5998 ( .A0(n5254), .A1(n1125), .B0(n5208), .B1(n2697), .Y(n9485) );
  NAND4X2 U5999 ( .A(n9476), .B(n9475), .C(n9474), .D(n9473), .Y(n11328) );
  OA22XL U6000 ( .A0(n5433), .A1(n1126), .B0(n5391), .B1(n2698), .Y(n9473) );
  OA22XL U6001 ( .A0(n5168), .A1(n1127), .B0(n5124), .B1(n2699), .Y(n9476) );
  OA22XL U6002 ( .A0(n5254), .A1(n1128), .B0(n5208), .B1(n2700), .Y(n9475) );
  NAND4BX2 U6003 ( .AN(n4486), .B(n9540), .C(n9539), .D(n9538), .Y(n11331) );
  NAND4X2 U6004 ( .A(n9663), .B(n9662), .C(n9661), .D(n9660), .Y(n11304) );
  OA22XL U6005 ( .A0(n5435), .A1(n1129), .B0(n5390), .B1(n2701), .Y(n9660) );
  OA22XL U6006 ( .A0(n5172), .A1(n1130), .B0(n5127), .B1(n2702), .Y(n9663) );
  OA22XL U6007 ( .A0(n5258), .A1(n1131), .B0(n5212), .B1(n2703), .Y(n9662) );
  NAND4X2 U6008 ( .A(n9536), .B(n9535), .C(n9534), .D(n9533), .Y(n11267) );
  OA22XL U6009 ( .A0(n5435), .A1(n1132), .B0(n5389), .B1(n2704), .Y(n9533) );
  OA22XL U6010 ( .A0(n5170), .A1(n1133), .B0(n5126), .B1(n2705), .Y(n9536) );
  OA22XL U6011 ( .A0(n5256), .A1(n1134), .B0(n5210), .B1(n2706), .Y(n9535) );
  OA22XL U6012 ( .A0(n5435), .A1(n1135), .B0(n5389), .B1(n2707), .Y(n9528) );
  OA22XL U6013 ( .A0(n5170), .A1(n1136), .B0(n5126), .B1(n2708), .Y(n9531) );
  OA22XL U6014 ( .A0(n5256), .A1(n1137), .B0(n5210), .B1(n2709), .Y(n9530) );
  NAND4X2 U6015 ( .A(n9598), .B(n9597), .C(n9596), .D(n9595), .Y(n11263) );
  OA22XL U6016 ( .A0(n5442), .A1(n2557), .B0(n5398), .B1(n786), .Y(n9595) );
  OA22XL U6017 ( .A0(n5171), .A1(n1138), .B0(n5134), .B1(n2710), .Y(n9598) );
  OA22XL U6018 ( .A0(n5257), .A1(n1139), .B0(n5211), .B1(n2711), .Y(n9597) );
  NAND4X2 U6019 ( .A(n9594), .B(n9593), .C(n9592), .D(n9591), .Y(n11295) );
  OA22XL U6020 ( .A0(n5429), .A1(n1140), .B0(n5385), .B1(n2712), .Y(n9357) );
  OA22XL U6021 ( .A0(n5164), .A1(n1141), .B0(n5121), .B1(n2713), .Y(n9360) );
  OA22XL U6022 ( .A0(n5250), .A1(n1142), .B0(n5213), .B1(n2714), .Y(n9359) );
  NAND4X2 U6023 ( .A(n9481), .B(n9480), .C(n9479), .D(n9478), .Y(n11232) );
  NAND4X2 U6024 ( .A(n9545), .B(n9544), .C(n9543), .D(n9542), .Y(n11235) );
  OA22XL U6025 ( .A0(n5446), .A1(n1143), .B0(n5389), .B1(n2715), .Y(n9542) );
  OA22XL U6026 ( .A0(n5170), .A1(n1144), .B0(n5126), .B1(n2716), .Y(n9545) );
  OA22XL U6027 ( .A0(n5256), .A1(n1145), .B0(n5210), .B1(n2717), .Y(n9544) );
  OA22XL U6028 ( .A0(n5429), .A1(n1146), .B0(n5385), .B1(n2718), .Y(n9352) );
  OA22XL U6029 ( .A0(n5164), .A1(n1147), .B0(n5123), .B1(n2719), .Y(n9355) );
  OA22XL U6030 ( .A0(n5250), .A1(n1148), .B0(n5213), .B1(n2720), .Y(n9354) );
  OA22XL U6031 ( .A0(n5431), .A1(n1149), .B0(n5389), .B1(n2721), .Y(n9523) );
  OA22XL U6032 ( .A0(n5170), .A1(n1150), .B0(n5126), .B1(n2722), .Y(n9526) );
  OA22XL U6033 ( .A0(n5256), .A1(n1151), .B0(n5210), .B1(n2723), .Y(n9525) );
  OA22XL U6034 ( .A0(net112453), .A1(n1499), .B0(net112329), .B1(n3112), .Y(
        n6283) );
  OA22XL U6035 ( .A0(net112041), .A1(n1500), .B0(net111917), .B1(n3113), .Y(
        n6281) );
  NAND2XL U6036 ( .A(n7956), .B(n8250), .Y(n7964) );
  NAND2XL U6037 ( .A(n8521), .B(n8520), .Y(n8530) );
  NAND2XL U6038 ( .A(n7853), .B(n7852), .Y(n7862) );
  INVX3 U6039 ( .A(n11078), .Y(n11075) );
  NOR4XL U6040 ( .A(n6624), .B(n6483), .C(n6625), .D(n6487), .Y(n6484) );
  INVXL U6041 ( .A(n7853), .Y(n6483) );
  AO22XL U6042 ( .A0(n4977), .A1(n543), .B0(n9309), .B1(n2298), .Y(n9202) );
  AO22XL U6043 ( .A0(n9310), .A1(n544), .B0(n9309), .B1(n2299), .Y(n9193) );
  AO22XL U6044 ( .A0(n4859), .A1(n293), .B0(n4869), .B1(n1873), .Y(n7654) );
  AO22XL U6045 ( .A0(n4845), .A1(n294), .B0(n4852), .B1(n1866), .Y(n7653) );
  NAND2XL U6046 ( .A(n11221), .B(n11220), .Y(n9181) );
  INVX3 U6047 ( .A(n10929), .Y(n10905) );
  INVX3 U6048 ( .A(n11088), .Y(n11085) );
  INVXL U6049 ( .A(n8524), .Y(n6487) );
  INVXL U6050 ( .A(n7693), .Y(n8436) );
  AOI2BB1XL U6051 ( .A0N(n9127), .A1N(n9272), .B0(n4682), .Y(n9135) );
  INVXL U6052 ( .A(n6946), .Y(n6416) );
  AND2XL U6053 ( .A(n10448), .B(n10447), .Y(n4572) );
  AND2XL U6054 ( .A(net99536), .B(net99537), .Y(n4574) );
  AO22XL U6055 ( .A0(n4951), .A1(n299), .B0(n4956), .B1(n1872), .Y(n6505) );
  AO22XL U6056 ( .A0(n4951), .A1(n298), .B0(n4956), .B1(n1871), .Y(n6522) );
  AO22XL U6057 ( .A0(n432), .A1(n234), .B0(n4839), .B1(n1832), .Y(n7766) );
  AO22XL U6058 ( .A0(n432), .A1(n235), .B0(n4838), .B1(n1833), .Y(n7757) );
  AO22XL U6059 ( .A0(n432), .A1(n246), .B0(n4837), .B1(n1874), .Y(n7661) );
  AO22XL U6060 ( .A0(n432), .A1(n247), .B0(n4836), .B1(n1875), .Y(n7652) );
  AO22XL U6061 ( .A0(n432), .A1(n249), .B0(n4840), .B1(n1868), .Y(n9214) );
  NAND2XL U6062 ( .A(n3766), .B(n7193), .Y(n7205) );
  AND2XL U6063 ( .A(n9162), .B(n9161), .Y(n4592) );
  INVXL U6064 ( .A(n7193), .Y(n7204) );
  CLKBUFX2 U6065 ( .A(n312), .Y(n5455) );
  NAND4X2 U6066 ( .A(n6721), .B(n6720), .C(n6719), .D(n6718), .Y(n11511) );
  OA22XL U6067 ( .A0(net112457), .A1(n1501), .B0(net112333), .B1(n3114), .Y(
        n6720) );
  OA22XL U6068 ( .A0(net112233), .A1(n1502), .B0(net112165), .B1(n3115), .Y(
        n6719) );
  OA22XL U6069 ( .A0(net112679), .A1(n1503), .B0(net112577), .B1(n3116), .Y(
        n6721) );
  NAND4X2 U6070 ( .A(n6788), .B(n6787), .C(n6786), .D(n6785), .Y(n11428) );
  OA22XL U6071 ( .A0(net112459), .A1(n1504), .B0(net112335), .B1(n3117), .Y(
        n6787) );
  OA22XL U6072 ( .A0(net112235), .A1(n1505), .B0(net112165), .B1(n3118), .Y(
        n6786) );
  OA22XL U6073 ( .A0(net112679), .A1(n1506), .B0(net112577), .B1(n3119), .Y(
        n6788) );
  NAND4X2 U6074 ( .A(n7062), .B(n7061), .C(n7060), .D(n7059), .Y(n11466) );
  NAND4X2 U6075 ( .A(n9968), .B(n9967), .C(n9966), .D(n9965), .Y(n11273) );
  OA22XL U6076 ( .A0(n5442), .A1(n1152), .B0(n5396), .B1(n2724), .Y(n9955) );
  OA22XL U6077 ( .A0(n5179), .A1(n1153), .B0(n5135), .B1(n2725), .Y(n9958) );
  OA22XL U6078 ( .A0(n5265), .A1(n1154), .B0(n5220), .B1(n2726), .Y(n9957) );
  OA22XL U6079 ( .A0(net112083), .A1(n1155), .B0(net111959), .B1(n2727), .Y(
        n4490) );
  AND2XL U6080 ( .A(n6432), .B(\i_MIPS/n371 ), .Y(n6433) );
  NOR3X1 U6081 ( .A(n229), .B(n287), .C(n4705), .Y(\i_MIPS/Register/n105 ) );
  OA22XL U6082 ( .A0(n5183), .A1(n1156), .B0(n5137), .B1(n2728), .Y(n10230) );
  OA22XL U6083 ( .A0(n5268), .A1(n1157), .B0(n5223), .B1(n2729), .Y(n10229) );
  OA22XL U6084 ( .A0(n5445), .A1(n1158), .B0(n5399), .B1(n2730), .Y(n10227) );
  OA22XL U6085 ( .A0(n5175), .A1(n2558), .B0(n5130), .B1(n787), .Y(n9778) );
  OA22XL U6086 ( .A0(n5261), .A1(n2559), .B0(n5215), .B1(n788), .Y(n9777) );
  OA22XL U6087 ( .A0(n5438), .A1(n2560), .B0(n5387), .B1(n789), .Y(n9775) );
  OA22XL U6088 ( .A0(n5174), .A1(n2561), .B0(n5129), .B1(n790), .Y(n9768) );
  OA22XL U6089 ( .A0(n5260), .A1(n2562), .B0(n5214), .B1(n791), .Y(n9767) );
  OA22XL U6090 ( .A0(n5437), .A1(n2563), .B0(n5392), .B1(n792), .Y(n9765) );
  OA22XL U6091 ( .A0(n5173), .A1(n1159), .B0(n5128), .B1(n2731), .Y(n9734) );
  OA22XL U6092 ( .A0(n5259), .A1(n1160), .B0(n5213), .B1(n2732), .Y(n9733) );
  OA22XL U6093 ( .A0(n5436), .A1(n1161), .B0(n5391), .B1(n2733), .Y(n9731) );
  OA22XL U6094 ( .A0(n5173), .A1(n1162), .B0(n5128), .B1(n2734), .Y(n9724) );
  OA22XL U6095 ( .A0(n5259), .A1(n1163), .B0(n5213), .B1(n2735), .Y(n9723) );
  OA22XL U6096 ( .A0(n5436), .A1(n1164), .B0(n5391), .B1(n2736), .Y(n9721) );
  OA22XL U6097 ( .A0(n5173), .A1(n1165), .B0(n5128), .B1(n2737), .Y(n9729) );
  OA22XL U6098 ( .A0(n5259), .A1(n1166), .B0(n5213), .B1(n2738), .Y(n9728) );
  OA22XL U6099 ( .A0(n5436), .A1(n1167), .B0(n5391), .B1(n2739), .Y(n9726) );
  OA22XL U6100 ( .A0(n5183), .A1(n1734), .B0(n5136), .B1(n3418), .Y(n10123) );
  OA22XL U6101 ( .A0(n5268), .A1(n1735), .B0(n5223), .B1(n3419), .Y(n10122) );
  OA22XL U6102 ( .A0(n5445), .A1(n1736), .B0(n5399), .B1(n3420), .Y(n10120) );
  OA22XL U6103 ( .A0(n5183), .A1(n1737), .B0(n5136), .B1(n3421), .Y(n10113) );
  OA22XL U6104 ( .A0(n5268), .A1(n1738), .B0(n5223), .B1(n3422), .Y(n10112) );
  OA22XL U6105 ( .A0(n5445), .A1(n1739), .B0(n5399), .B1(n3423), .Y(n10110) );
  OA22XL U6106 ( .A0(n5178), .A1(n1740), .B0(n5134), .B1(n3424), .Y(n9925) );
  OA22XL U6107 ( .A0(n5264), .A1(n1741), .B0(n5219), .B1(n3425), .Y(n9924) );
  OA22XL U6108 ( .A0(n5441), .A1(n1742), .B0(n5395), .B1(n3426), .Y(n9922) );
  OA22XL U6109 ( .A0(n5176), .A1(n1743), .B0(n5131), .B1(n3427), .Y(n9847) );
  OA22XL U6110 ( .A0(n5262), .A1(n1744), .B0(n5216), .B1(n3428), .Y(n9846) );
  OA22XL U6111 ( .A0(n5439), .A1(n1745), .B0(n5393), .B1(n3429), .Y(n9844) );
  OA22XL U6112 ( .A0(n5179), .A1(n1746), .B0(n5135), .B1(n3430), .Y(n9982) );
  OA22XL U6113 ( .A0(n5265), .A1(n1747), .B0(n5220), .B1(n3431), .Y(n9981) );
  OA22XL U6114 ( .A0(n5442), .A1(n1748), .B0(n5396), .B1(n3432), .Y(n9979) );
  OA22XL U6115 ( .A0(n5177), .A1(n1749), .B0(n5138), .B1(n3433), .Y(n11133) );
  OA22XL U6116 ( .A0(n5269), .A1(n1750), .B0(n5221), .B1(n3434), .Y(n11132) );
  OA22XL U6117 ( .A0(n5446), .A1(n1751), .B0(n5400), .B1(n3435), .Y(n11130) );
  OA22XL U6118 ( .A0(n5177), .A1(n1752), .B0(n5138), .B1(n3436), .Y(n11144) );
  OA22XL U6119 ( .A0(n5269), .A1(n1753), .B0(n5221), .B1(n3437), .Y(n11143) );
  OA22XL U6120 ( .A0(n5446), .A1(n1754), .B0(n5400), .B1(n3438), .Y(n11141) );
  OA22XL U6121 ( .A0(n5177), .A1(n1755), .B0(n5138), .B1(n3439), .Y(n11128) );
  OA22XL U6122 ( .A0(n5269), .A1(n1756), .B0(n5217), .B1(n3440), .Y(n11127) );
  OA22XL U6123 ( .A0(n5446), .A1(n1757), .B0(n5400), .B1(n3441), .Y(n11125) );
  OA22XL U6124 ( .A0(n5182), .A1(n1758), .B0(n5137), .B1(n3442), .Y(n10074) );
  OA22XL U6125 ( .A0(n5267), .A1(n1759), .B0(n5222), .B1(n3443), .Y(n10073) );
  OA22XL U6126 ( .A0(n5444), .A1(n1760), .B0(n5398), .B1(n3444), .Y(n10071) );
  OA22XL U6127 ( .A0(n5172), .A1(n1761), .B0(n5127), .B1(n3445), .Y(n9682) );
  OA22XL U6128 ( .A0(n5258), .A1(n1762), .B0(n5212), .B1(n3446), .Y(n9681) );
  OA22XL U6129 ( .A0(n5435), .A1(n1763), .B0(n5390), .B1(n3447), .Y(n9679) );
  OA22XL U6130 ( .A0(n5182), .A1(n1764), .B0(n5137), .B1(n3448), .Y(n10108) );
  OA22XL U6131 ( .A0(n5267), .A1(n1765), .B0(n5222), .B1(n3449), .Y(n10107) );
  OA22XL U6132 ( .A0(n5444), .A1(n1766), .B0(n5398), .B1(n3450), .Y(n10105) );
  OA22XL U6133 ( .A0(n5183), .A1(n1767), .B0(n5136), .B1(n3451), .Y(n10118) );
  OA22XL U6134 ( .A0(n5268), .A1(n1768), .B0(n5223), .B1(n3452), .Y(n10117) );
  OA22XL U6135 ( .A0(n5445), .A1(n1769), .B0(n5399), .B1(n3453), .Y(n10115) );
  OA22XL U6136 ( .A0(n5178), .A1(n1770), .B0(n5134), .B1(n3454), .Y(n9920) );
  OA22XL U6137 ( .A0(n5264), .A1(n1771), .B0(n5219), .B1(n3455), .Y(n9919) );
  OA22XL U6138 ( .A0(n5441), .A1(n1772), .B0(n5395), .B1(n3456), .Y(n9917) );
  OA22XL U6139 ( .A0(n5176), .A1(n1773), .B0(n5131), .B1(n3457), .Y(n9842) );
  OA22XL U6140 ( .A0(n5262), .A1(n1774), .B0(n5216), .B1(n3458), .Y(n9841) );
  OA22XL U6141 ( .A0(n5439), .A1(n1775), .B0(n5393), .B1(n3459), .Y(n9839) );
  OA22XL U6142 ( .A0(n5179), .A1(n1776), .B0(n5135), .B1(n3460), .Y(n9977) );
  OA22XL U6143 ( .A0(n5265), .A1(n1777), .B0(n5220), .B1(n3461), .Y(n9976) );
  OA22XL U6144 ( .A0(n5442), .A1(n1778), .B0(n5396), .B1(n3462), .Y(n9974) );
  OA22XL U6145 ( .A0(n5179), .A1(n1779), .B0(n5135), .B1(n3463), .Y(n9987) );
  OA22XL U6146 ( .A0(n5265), .A1(n1780), .B0(n5220), .B1(n3464), .Y(n9986) );
  OA22XL U6147 ( .A0(n5442), .A1(n1781), .B0(n5396), .B1(n3465), .Y(n9984) );
  OA22XL U6148 ( .A0(n5177), .A1(n1782), .B0(n5138), .B1(n3466), .Y(n11123) );
  OA22XL U6149 ( .A0(n5269), .A1(n1783), .B0(n5217), .B1(n3467), .Y(n11122) );
  OA22XL U6150 ( .A0(n5446), .A1(n1784), .B0(n5400), .B1(n3468), .Y(n11120) );
  NAND2XL U6151 ( .A(DCACHE_addr[2]), .B(net113087), .Y(net100048) );
  NAND2XL U6152 ( .A(DCACHE_addr[16]), .B(net113089), .Y(net99288) );
  NAND2XL U6153 ( .A(DCACHE_addr[21]), .B(net113089), .Y(net99382) );
  NAND2XL U6154 ( .A(n10671), .B(n10670), .Y(n11532) );
  NAND2XL U6155 ( .A(n1632), .B(n3297), .Y(n11531) );
  NAND2XL U6156 ( .A(n3734), .B(n10664), .Y(n11523) );
  NAND2XL U6157 ( .A(n3202), .B(n10666), .Y(n11528) );
  NAND2XL U6158 ( .A(n10656), .B(n10655), .Y(n11522) );
  NAND2XL U6159 ( .A(n10648), .B(n10647), .Y(n11525) );
  NAND2XL U6160 ( .A(n10635), .B(n10634), .Y(n11526) );
  NAND2XL U6161 ( .A(n2437), .B(n10673), .Y(n11530) );
  NAND2XL U6162 ( .A(n10632), .B(n3745), .Y(n11518) );
  AOI2BB1XL U6163 ( .A0N(n9273), .A1N(n177), .B0(n4673), .Y(n9276) );
  NAND2X1 U6164 ( .A(\i_MIPS/Register/n117 ), .B(\i_MIPS/Register/n104 ), .Y(
        \i_MIPS/Register/n116 ) );
  NAND2X1 U6165 ( .A(\i_MIPS/Register/n115 ), .B(\i_MIPS/Register/n104 ), .Y(
        \i_MIPS/Register/n114 ) );
  NAND2X1 U6166 ( .A(\i_MIPS/Register/n113 ), .B(\i_MIPS/Register/n104 ), .Y(
        \i_MIPS/Register/n112 ) );
  NAND2X1 U6167 ( .A(\i_MIPS/Register/n111 ), .B(\i_MIPS/Register/n104 ), .Y(
        \i_MIPS/Register/n110 ) );
  NAND2X1 U6168 ( .A(\i_MIPS/Register/n109 ), .B(\i_MIPS/Register/n104 ), .Y(
        \i_MIPS/Register/n108 ) );
  NAND2X1 U6169 ( .A(\i_MIPS/Register/n107 ), .B(\i_MIPS/Register/n104 ), .Y(
        \i_MIPS/Register/n106 ) );
  NAND2X1 U6170 ( .A(\i_MIPS/Register/n119 ), .B(\i_MIPS/Register/n104 ), .Y(
        \i_MIPS/Register/n118 ) );
  NAND2X1 U6171 ( .A(\i_MIPS/Register/n131 ), .B(\i_MIPS/Register/n119 ), .Y(
        \i_MIPS/Register/n138 ) );
  NAND2X1 U6172 ( .A(\i_MIPS/Register/n131 ), .B(\i_MIPS/Register/n117 ), .Y(
        \i_MIPS/Register/n137 ) );
  NAND2X1 U6173 ( .A(\i_MIPS/Register/n131 ), .B(\i_MIPS/Register/n115 ), .Y(
        \i_MIPS/Register/n136 ) );
  NAND2X1 U6174 ( .A(\i_MIPS/Register/n131 ), .B(\i_MIPS/Register/n113 ), .Y(
        \i_MIPS/Register/n135 ) );
  NAND2X1 U6175 ( .A(\i_MIPS/Register/n131 ), .B(\i_MIPS/Register/n111 ), .Y(
        \i_MIPS/Register/n134 ) );
  NAND2X1 U6176 ( .A(\i_MIPS/Register/n131 ), .B(\i_MIPS/Register/n109 ), .Y(
        \i_MIPS/Register/n133 ) );
  NAND2X1 U6177 ( .A(\i_MIPS/Register/n131 ), .B(\i_MIPS/Register/n107 ), .Y(
        \i_MIPS/Register/n132 ) );
  NAND2X1 U6178 ( .A(\i_MIPS/Register/n131 ), .B(\i_MIPS/Register/n105 ), .Y(
        \i_MIPS/Register/n130 ) );
  NAND2X1 U6179 ( .A(\i_MIPS/Register/n122 ), .B(\i_MIPS/Register/n119 ), .Y(
        \i_MIPS/Register/n129 ) );
  NAND2X1 U6180 ( .A(\i_MIPS/Register/n122 ), .B(\i_MIPS/Register/n117 ), .Y(
        \i_MIPS/Register/n128 ) );
  NAND2X1 U6181 ( .A(\i_MIPS/Register/n122 ), .B(\i_MIPS/Register/n115 ), .Y(
        \i_MIPS/Register/n127 ) );
  NAND2X1 U6182 ( .A(\i_MIPS/Register/n122 ), .B(\i_MIPS/Register/n113 ), .Y(
        \i_MIPS/Register/n126 ) );
  NAND2X1 U6183 ( .A(\i_MIPS/Register/n122 ), .B(\i_MIPS/Register/n111 ), .Y(
        \i_MIPS/Register/n125 ) );
  NAND2X1 U6184 ( .A(\i_MIPS/Register/n122 ), .B(\i_MIPS/Register/n109 ), .Y(
        \i_MIPS/Register/n124 ) );
  NAND2X1 U6185 ( .A(\i_MIPS/Register/n122 ), .B(\i_MIPS/Register/n107 ), .Y(
        \i_MIPS/Register/n123 ) );
  NAND2X1 U6186 ( .A(\i_MIPS/Register/n122 ), .B(\i_MIPS/Register/n105 ), .Y(
        \i_MIPS/Register/n121 ) );
  AO21X1 U6187 ( .A0(\i_MIPS/Register/n104 ), .A1(\i_MIPS/Register/n105 ), 
        .B0(n4638), .Y(n10836) );
  NAND4X2 U6188 ( .A(n4491), .B(n9331), .C(n9330), .D(n9329), .Y(n9345) );
  OA22XL U6189 ( .A0(n5173), .A1(n1168), .B0(n5128), .B1(n2740), .Y(n9719) );
  OA22XL U6190 ( .A0(n5259), .A1(n1169), .B0(n5213), .B1(n2741), .Y(n9718) );
  OA22XL U6191 ( .A0(n5436), .A1(n1170), .B0(n5391), .B1(n2742), .Y(n9716) );
  OA22XL U6192 ( .A0(n5175), .A1(n1171), .B0(n5130), .B1(n2743), .Y(n9802) );
  OA22XL U6193 ( .A0(n5261), .A1(n1172), .B0(n5215), .B1(n2744), .Y(n9801) );
  OA22XL U6194 ( .A0(n5438), .A1(n1173), .B0(n5393), .B1(n2745), .Y(n9799) );
  OA22XL U6195 ( .A0(n5174), .A1(n1174), .B0(n5129), .B1(n2746), .Y(n9755) );
  OA22XL U6196 ( .A0(n5260), .A1(n1175), .B0(n5214), .B1(n2747), .Y(n9754) );
  OA22XL U6197 ( .A0(n5437), .A1(n1176), .B0(n5392), .B1(n2748), .Y(n9752) );
  OA22XL U6198 ( .A0(n5175), .A1(n1177), .B0(n5130), .B1(n2749), .Y(n9797) );
  OA22XL U6199 ( .A0(n5438), .A1(n1178), .B0(n5399), .B1(n2750), .Y(n9794) );
  OA22XL U6200 ( .A0(n5174), .A1(n1179), .B0(n5129), .B1(n2751), .Y(n9751) );
  OA22XL U6201 ( .A0(n5175), .A1(n1180), .B0(n5130), .B1(n2752), .Y(n9792) );
  OA22XL U6202 ( .A0(n5261), .A1(n1181), .B0(n5215), .B1(n2753), .Y(n9791) );
  OA22XL U6203 ( .A0(n5438), .A1(n1182), .B0(n5384), .B1(n2754), .Y(n9789) );
  OA22XL U6204 ( .A0(n5174), .A1(n1183), .B0(n5129), .B1(n2755), .Y(n9747) );
  OA22XL U6205 ( .A0(n5260), .A1(n1184), .B0(n5214), .B1(n2756), .Y(n9746) );
  OA22XL U6206 ( .A0(n5437), .A1(n1185), .B0(n5392), .B1(n2757), .Y(n9744) );
  OA22XL U6207 ( .A0(n5175), .A1(n1186), .B0(n5130), .B1(n2758), .Y(n9773) );
  OA22XL U6208 ( .A0(n5261), .A1(n1187), .B0(n5215), .B1(n2759), .Y(n9772) );
  OA22XL U6209 ( .A0(n5438), .A1(n2564), .B0(n5401), .B1(n793), .Y(n9770) );
  NAND2X1 U6210 ( .A(\i_MIPS/Register/n140 ), .B(\i_MIPS/Register/n119 ), .Y(
        \i_MIPS/Register/n147 ) );
  NAND2X1 U6211 ( .A(\i_MIPS/Register/n140 ), .B(\i_MIPS/Register/n111 ), .Y(
        \i_MIPS/Register/n143 ) );
  NAND2X1 U6212 ( .A(\i_MIPS/Register/n140 ), .B(\i_MIPS/Register/n109 ), .Y(
        \i_MIPS/Register/n142 ) );
  NAND2X1 U6213 ( .A(\i_MIPS/Register/n140 ), .B(\i_MIPS/Register/n107 ), .Y(
        \i_MIPS/Register/n141 ) );
  NAND2X1 U6214 ( .A(\i_MIPS/Register/n140 ), .B(\i_MIPS/Register/n117 ), .Y(
        \i_MIPS/Register/n146 ) );
  NAND2X1 U6215 ( .A(\i_MIPS/Register/n140 ), .B(\i_MIPS/Register/n115 ), .Y(
        \i_MIPS/Register/n145 ) );
  NAND2X1 U6216 ( .A(\i_MIPS/Register/n140 ), .B(\i_MIPS/Register/n113 ), .Y(
        \i_MIPS/Register/n144 ) );
  NAND2X1 U6217 ( .A(\i_MIPS/Register/n140 ), .B(\i_MIPS/Register/n105 ), .Y(
        \i_MIPS/Register/n139 ) );
  NAND2XL U6218 ( .A(\i_MIPS/IF_ID_28 ), .B(net130576), .Y(n10393) );
  OAI221X2 U6219 ( .A0(net112257), .A1(n1617), .B0(net112137), .B1(n224), .C0(
        n6052), .Y(n6053) );
  AO22XL U6220 ( .A0(n176), .A1(n11028), .B0(net113592), .B1(
        \i_MIPS/IR_ID[19] ), .Y(\i_MIPS/N74 ) );
  AO22XL U6221 ( .A0(n175), .A1(n10943), .B0(net113592), .B1(n10080), .Y(
        \i_MIPS/N71 ) );
  OA22X4 U6222 ( .A0(net112087), .A1(n1974), .B0(net111955), .B1(n406), .Y(
        n6093) );
  OA22X4 U6223 ( .A0(net112087), .A1(n1975), .B0(net111915), .B1(n407), .Y(
        n6066) );
  BUFX20 U6224 ( .A(\i_MIPS/ID_EX[82] ), .Y(n4802) );
  OA22XL U6225 ( .A0(n9276), .A1(n9275), .B0(n9275), .B1(n9274), .Y(n9289) );
  INVXL U6226 ( .A(n11466), .Y(n10189) );
  INVXL U6227 ( .A(n11437), .Y(n10604) );
  INVXL U6228 ( .A(n11406), .Y(n10601) );
  INVXL U6229 ( .A(n11468), .Y(n10598) );
  INVXL U6230 ( .A(n11459), .Y(n10820) );
  INVXL U6231 ( .A(n11428), .Y(n10826) );
  AOI2BB1XL U6232 ( .A0N(n3827), .A1N(n3592), .B0(n4600), .Y(n6952) );
  INVXL U6233 ( .A(n9128), .Y(n9132) );
  OA22XL U6234 ( .A0(\i_MIPS/Register/register[6][20] ), .A1(n4913), .B0(
        \i_MIPS/Register/register[14][20] ), .B1(n4907), .Y(n8565) );
  OA22XL U6235 ( .A0(\i_MIPS/Register/register[6][16] ), .A1(n4913), .B0(
        \i_MIPS/Register/register[14][16] ), .B1(n4907), .Y(n8175) );
  OA22XL U6236 ( .A0(\i_MIPS/Register/register[6][21] ), .A1(n4912), .B0(
        \i_MIPS/Register/register[14][21] ), .B1(n4906), .Y(n8051) );
  OA22XL U6237 ( .A0(\i_MIPS/Register/register[6][23] ), .A1(n4913), .B0(
        \i_MIPS/Register/register[14][23] ), .B1(n4907), .Y(n8233) );
  OA22XL U6238 ( .A0(\i_MIPS/Register/register[6][27] ), .A1(n4913), .B0(
        \i_MIPS/Register/register[14][27] ), .B1(n4907), .Y(n8624) );
  OA22XL U6239 ( .A0(\i_MIPS/Register/register[6][4] ), .A1(n4911), .B0(
        \i_MIPS/Register/register[14][4] ), .B1(n4903), .Y(n7377) );
  MXI2X1 U6240 ( .A(\i_MIPS/n370 ), .B(net98901), .S0(n5502), .Y(\i_MIPS/n561 ) );
  OA22XL U6241 ( .A0(\i_MIPS/Register/register[6][19] ), .A1(n4912), .B0(
        \i_MIPS/Register/register[14][19] ), .B1(n4906), .Y(n7756) );
  MXI2XL U6242 ( .A(n4704), .B(\i_MIPS/n222 ), .S0(n5507), .Y(\i_MIPS/n502 )
         );
  MXI2XL U6243 ( .A(\i_MIPS/n258 ), .B(\i_MIPS/n259 ), .S0(n5506), .Y(
        \i_MIPS/n386 ) );
  MXI2XL U6244 ( .A(n4709), .B(\i_MIPS/n225 ), .S0(n5507), .Y(\i_MIPS/n499 )
         );
  MXI2XL U6245 ( .A(\i_MIPS/n298 ), .B(\i_MIPS/n299 ), .S0(n5505), .Y(
        \i_MIPS/n426 ) );
  MXI2XL U6246 ( .A(\i_MIPS/n276 ), .B(\i_MIPS/n277 ), .S0(n5505), .Y(
        \i_MIPS/n404 ) );
  MXI2XL U6247 ( .A(\i_MIPS/n270 ), .B(\i_MIPS/n271 ), .S0(n5505), .Y(
        \i_MIPS/n398 ) );
  MXI2XL U6248 ( .A(\i_MIPS/n268 ), .B(\i_MIPS/n269 ), .S0(n5505), .Y(
        \i_MIPS/n396 ) );
  MXI2XL U6249 ( .A(\i_MIPS/n286 ), .B(\i_MIPS/n287 ), .S0(n5503), .Y(
        \i_MIPS/n414 ) );
  MXI2XL U6250 ( .A(\i_MIPS/n284 ), .B(\i_MIPS/n285 ), .S0(n5503), .Y(
        \i_MIPS/n412 ) );
  MXI2XL U6251 ( .A(\i_MIPS/n282 ), .B(\i_MIPS/n283 ), .S0(n5503), .Y(
        \i_MIPS/n410 ) );
  MXI2XL U6252 ( .A(\i_MIPS/n266 ), .B(\i_MIPS/n267 ), .S0(n5503), .Y(
        \i_MIPS/n394 ) );
  MXI2XL U6253 ( .A(\i_MIPS/n264 ), .B(\i_MIPS/n265 ), .S0(n5503), .Y(
        \i_MIPS/n392 ) );
  MXI2XL U6254 ( .A(\i_MIPS/n260 ), .B(\i_MIPS/n261 ), .S0(n5503), .Y(
        \i_MIPS/n388 ) );
  MXI2XL U6255 ( .A(n4712), .B(\i_MIPS/n223 ), .S0(n5508), .Y(\i_MIPS/n501 )
         );
  MXI2XL U6256 ( .A(n4713), .B(\i_MIPS/n226 ), .S0(n5508), .Y(\i_MIPS/n498 )
         );
  MXI2XL U6257 ( .A(\i_MIPS/n288 ), .B(\i_MIPS/n289 ), .S0(n5502), .Y(
        \i_MIPS/n416 ) );
  MXI2XL U6258 ( .A(\i_MIPS/n274 ), .B(\i_MIPS/n275 ), .S0(n5502), .Y(
        \i_MIPS/n402 ) );
  MXI2XL U6259 ( .A(\i_MIPS/n272 ), .B(\i_MIPS/n273 ), .S0(n5502), .Y(
        \i_MIPS/n400 ) );
  MXI2XL U6260 ( .A(\i_MIPS/n300 ), .B(\i_MIPS/n301 ), .S0(n5505), .Y(
        \i_MIPS/n428 ) );
  MXI2XL U6261 ( .A(\i_MIPS/n338 ), .B(\i_MIPS/n339 ), .S0(n5506), .Y(
        \i_MIPS/n529 ) );
  MXI2XL U6262 ( .A(\i_MIPS/n321 ), .B(\i_MIPS/n320 ), .S0(n5506), .Y(
        \i_MIPS/n517 ) );
  MXI2XL U6263 ( .A(\i_MIPS/n319 ), .B(\i_MIPS/n318 ), .S0(n5506), .Y(
        \i_MIPS/n516 ) );
  MXI2XL U6264 ( .A(\i_MIPS/n371 ), .B(n4546), .S0(n5503), .Y(\i_MIPS/n562 )
         );
  MXI2XL U6265 ( .A(\i_MIPS/n368 ), .B(n4556), .S0(n5503), .Y(\i_MIPS/n559 )
         );
  MXI2XL U6266 ( .A(\i_MIPS/n358 ), .B(n4538), .S0(n5503), .Y(\i_MIPS/n549 )
         );
  MXI2XL U6267 ( .A(\i_MIPS/n344 ), .B(n4530), .S0(n5503), .Y(\i_MIPS/n535 )
         );
  MXI2XL U6268 ( .A(\i_MIPS/n342 ), .B(n4524), .S0(n5503), .Y(\i_MIPS/n533 )
         );
  MXI2XL U6269 ( .A(\i_MIPS/n333 ), .B(\i_MIPS/n332 ), .S0(n5504), .Y(
        \i_MIPS/n523 ) );
  MXI2XL U6270 ( .A(\i_MIPS/n331 ), .B(\i_MIPS/n330 ), .S0(n5503), .Y(
        \i_MIPS/n522 ) );
  MXI2XL U6271 ( .A(\i_MIPS/n327 ), .B(\i_MIPS/n326 ), .S0(n5504), .Y(
        \i_MIPS/n520 ) );
  MXI2XL U6272 ( .A(\i_MIPS/n325 ), .B(\i_MIPS/n324 ), .S0(n5504), .Y(
        \i_MIPS/n519 ) );
  MXI2XL U6273 ( .A(\i_MIPS/n323 ), .B(\i_MIPS/n322 ), .S0(n5504), .Y(
        \i_MIPS/n518 ) );
  MXI2XL U6274 ( .A(\i_MIPS/n315 ), .B(\i_MIPS/n314 ), .S0(n5504), .Y(
        \i_MIPS/n514 ) );
  MXI2XL U6275 ( .A(\i_MIPS/n353 ), .B(n4559), .S0(n5502), .Y(\i_MIPS/n544 )
         );
  MXI2XL U6276 ( .A(\i_MIPS/n373 ), .B(\i_MIPS/n372 ), .S0(n5505), .Y(
        \i_MIPS/n563 ) );
  MXI2XL U6277 ( .A(\i_MIPS/n343 ), .B(n3552), .S0(n5505), .Y(\i_MIPS/n534 )
         );
  MXI2XL U6278 ( .A(\i_MIPS/n317 ), .B(\i_MIPS/n316 ), .S0(n5505), .Y(
        \i_MIPS/n515 ) );
  MXI2XL U6279 ( .A(\i_MIPS/n313 ), .B(\i_MIPS/n312 ), .S0(n5505), .Y(
        \i_MIPS/n513 ) );
  AOI2BB1XL U6280 ( .A0N(n8731), .A1N(n177), .B0(n4674), .Y(n7618) );
  OA22X1 U6281 ( .A0(net112673), .A1(n2809), .B0(net112571), .B1(n814), .Y(
        n7725) );
  INVX3 U6282 ( .A(n4771), .Y(n4791) );
  INVX16 U6283 ( .A(n4791), .Y(mem_addr_D[30]) );
  AO21X1 U6284 ( .A0(\i_MIPS/ID_EX[89] ), .A1(n5516), .B0(n4499), .Y(
        \i_MIPS/n496 ) );
  AO21X1 U6285 ( .A0(\i_MIPS/ID_EX[90] ), .A1(n5513), .B0(n4499), .Y(
        \i_MIPS/n495 ) );
  AO21X1 U6286 ( .A0(\i_MIPS/ID_EX[91] ), .A1(n5516), .B0(n4499), .Y(
        \i_MIPS/n494 ) );
  AO21X1 U6287 ( .A0(\i_MIPS/ID_EX[92] ), .A1(n5516), .B0(n4499), .Y(
        \i_MIPS/n493 ) );
  AO21X1 U6288 ( .A0(\i_MIPS/ID_EX[93] ), .A1(n5515), .B0(n4499), .Y(
        \i_MIPS/n492 ) );
  AO21X1 U6289 ( .A0(\i_MIPS/ID_EX[94] ), .A1(n5517), .B0(n4499), .Y(
        \i_MIPS/n491 ) );
  AO21X1 U6290 ( .A0(\i_MIPS/ID_EX[96] ), .A1(n5517), .B0(n4499), .Y(
        \i_MIPS/n489 ) );
  AO21X1 U6291 ( .A0(\i_MIPS/ID_EX[97] ), .A1(n5516), .B0(n4499), .Y(
        \i_MIPS/n488 ) );
  AO21X1 U6292 ( .A0(\i_MIPS/ID_EX[98] ), .A1(n5517), .B0(n4499), .Y(
        \i_MIPS/n487 ) );
  OA22XL U6293 ( .A0(\i_MIPS/Register/register[4][6] ), .A1(n4952), .B0(
        \i_MIPS/Register/register[12][6] ), .B1(n4949), .Y(n7530) );
  OA22XL U6294 ( .A0(\i_MIPS/Register/register[0][6] ), .A1(n4962), .B0(
        \i_MIPS/Register/register[8][6] ), .B1(n4958), .Y(n7529) );
  OA22XL U6295 ( .A0(\i_MIPS/Register/register[4][7] ), .A1(n4952), .B0(
        \i_MIPS/Register/register[12][7] ), .B1(n4949), .Y(n7438) );
  OA22XL U6296 ( .A0(\i_MIPS/Register/register[0][7] ), .A1(n4962), .B0(
        \i_MIPS/Register/register[8][7] ), .B1(n4958), .Y(n7437) );
  OA22XL U6297 ( .A0(\i_MIPS/Register/register[4][18] ), .A1(n4953), .B0(
        \i_MIPS/Register/register[12][18] ), .B1(n4949), .Y(n7937) );
  OA22XL U6298 ( .A0(\i_MIPS/Register/register[0][18] ), .A1(n4963), .B0(
        \i_MIPS/Register/register[8][18] ), .B1(n4959), .Y(n7936) );
  OA22XL U6299 ( .A0(\i_MIPS/Register/register[4][17] ), .A1(n4953), .B0(
        \i_MIPS/Register/register[12][17] ), .B1(n4949), .Y(n7680) );
  OA22XL U6300 ( .A0(\i_MIPS/Register/register[0][17] ), .A1(n4963), .B0(
        \i_MIPS/Register/register[8][17] ), .B1(n4959), .Y(n7679) );
  OA22XL U6301 ( .A0(\i_MIPS/Register/register[4][12] ), .A1(n4954), .B0(
        \i_MIPS/Register/register[12][12] ), .B1(n4948), .Y(n6181) );
  OA22XL U6302 ( .A0(\i_MIPS/Register/register[0][12] ), .A1(n4961), .B0(
        \i_MIPS/Register/register[8][12] ), .B1(n4957), .Y(n6180) );
  OA22XL U6303 ( .A0(\i_MIPS/Register/register[4][9] ), .A1(n4952), .B0(
        \i_MIPS/Register/register[12][9] ), .B1(n4948), .Y(n6831) );
  OA22XL U6304 ( .A0(\i_MIPS/Register/register[0][9] ), .A1(n4961), .B0(
        \i_MIPS/Register/register[8][9] ), .B1(n4957), .Y(n6830) );
  OA22XL U6305 ( .A0(\i_MIPS/Register/register[4][8] ), .A1(n4953), .B0(
        \i_MIPS/Register/register[12][8] ), .B1(n4948), .Y(n6751) );
  OA22XL U6306 ( .A0(\i_MIPS/Register/register[0][8] ), .A1(n4961), .B0(
        \i_MIPS/Register/register[8][8] ), .B1(n4957), .Y(n6750) );
  OA22XL U6307 ( .A0(\i_MIPS/Register/register[4][10] ), .A1(n4952), .B0(
        \i_MIPS/Register/register[12][10] ), .B1(n4949), .Y(n7256) );
  OA22XL U6308 ( .A0(\i_MIPS/Register/register[0][10] ), .A1(n4962), .B0(
        \i_MIPS/Register/register[8][10] ), .B1(n4958), .Y(n7255) );
  OA22XL U6309 ( .A0(\i_MIPS/Register/register[4][5] ), .A1(n4952), .B0(
        \i_MIPS/Register/register[12][5] ), .B1(n4949), .Y(n7340) );
  OA22XL U6310 ( .A0(\i_MIPS/Register/register[0][5] ), .A1(n4962), .B0(
        \i_MIPS/Register/register[8][5] ), .B1(n4958), .Y(n7339) );
  OA22XL U6311 ( .A0(\i_MIPS/Register/register[20][1] ), .A1(n4953), .B0(
        \i_MIPS/Register/register[28][1] ), .B1(n4949), .Y(n7606) );
  OA22XL U6312 ( .A0(\i_MIPS/Register/register[16][1] ), .A1(n4963), .B0(
        \i_MIPS/Register/register[24][1] ), .B1(n4959), .Y(n7605) );
  OA22XL U6313 ( .A0(\i_MIPS/Register/register[20][6] ), .A1(n4952), .B0(
        \i_MIPS/Register/register[28][6] ), .B1(n4948), .Y(n7539) );
  OA22XL U6314 ( .A0(\i_MIPS/Register/register[16][6] ), .A1(n4962), .B0(
        \i_MIPS/Register/register[24][6] ), .B1(n4958), .Y(n7538) );
  OA22XL U6315 ( .A0(\i_MIPS/Register/register[20][7] ), .A1(n4952), .B0(
        \i_MIPS/Register/register[28][7] ), .B1(n4949), .Y(n7447) );
  OA22XL U6316 ( .A0(\i_MIPS/Register/register[16][7] ), .A1(n4962), .B0(
        \i_MIPS/Register/register[24][7] ), .B1(n4958), .Y(n7446) );
  OA22XL U6317 ( .A0(\i_MIPS/Register/register[20][18] ), .A1(n4953), .B0(
        \i_MIPS/Register/register[28][18] ), .B1(n4949), .Y(n7946) );
  OA22XL U6318 ( .A0(\i_MIPS/Register/register[16][18] ), .A1(n4963), .B0(
        \i_MIPS/Register/register[24][18] ), .B1(n4959), .Y(n7945) );
  OA22XL U6319 ( .A0(\i_MIPS/Register/register[20][17] ), .A1(n4953), .B0(
        \i_MIPS/Register/register[28][17] ), .B1(n4949), .Y(n7689) );
  OA22XL U6320 ( .A0(\i_MIPS/Register/register[16][17] ), .A1(n4963), .B0(
        \i_MIPS/Register/register[24][17] ), .B1(n4959), .Y(n7688) );
  OA22XL U6321 ( .A0(\i_MIPS/Register/register[20][12] ), .A1(n4952), .B0(
        \i_MIPS/Register/register[28][12] ), .B1(n4948), .Y(n6190) );
  OA22XL U6322 ( .A0(\i_MIPS/Register/register[16][12] ), .A1(n4961), .B0(
        \i_MIPS/Register/register[24][12] ), .B1(n4957), .Y(n6189) );
  OA22XL U6323 ( .A0(\i_MIPS/Register/register[20][9] ), .A1(n4953), .B0(
        \i_MIPS/Register/register[28][9] ), .B1(n4948), .Y(n6840) );
  OA22XL U6324 ( .A0(\i_MIPS/Register/register[16][9] ), .A1(n4961), .B0(
        \i_MIPS/Register/register[24][9] ), .B1(n4957), .Y(n6839) );
  OA22XL U6325 ( .A0(\i_MIPS/Register/register[20][8] ), .A1(n4954), .B0(
        \i_MIPS/Register/register[28][8] ), .B1(n4948), .Y(n6760) );
  OA22XL U6326 ( .A0(\i_MIPS/Register/register[16][8] ), .A1(n4961), .B0(
        \i_MIPS/Register/register[24][8] ), .B1(n4957), .Y(n6759) );
  OA22XL U6327 ( .A0(\i_MIPS/Register/register[20][15] ), .A1(n4952), .B0(
        \i_MIPS/Register/register[28][15] ), .B1(n4949), .Y(n7015) );
  OA22XL U6328 ( .A0(\i_MIPS/Register/register[16][15] ), .A1(n4962), .B0(
        \i_MIPS/Register/register[24][15] ), .B1(n4958), .Y(n7014) );
  OA22XL U6329 ( .A0(\i_MIPS/Register/register[20][10] ), .A1(n4952), .B0(
        \i_MIPS/Register/register[28][10] ), .B1(n4949), .Y(n7265) );
  OA22XL U6330 ( .A0(\i_MIPS/Register/register[16][10] ), .A1(n4962), .B0(
        \i_MIPS/Register/register[24][10] ), .B1(n4958), .Y(n7264) );
  OA22XL U6331 ( .A0(\i_MIPS/Register/register[20][19] ), .A1(n4953), .B0(
        \i_MIPS/Register/register[28][19] ), .B1(n4949), .Y(n7842) );
  OA22XL U6332 ( .A0(\i_MIPS/Register/register[16][19] ), .A1(n4963), .B0(
        \i_MIPS/Register/register[24][19] ), .B1(n4959), .Y(n7841) );
  OA22XL U6333 ( .A0(\i_MIPS/Register/register[20][5] ), .A1(n4952), .B0(
        \i_MIPS/Register/register[28][5] ), .B1(n4949), .Y(n7349) );
  OA22XL U6334 ( .A0(\i_MIPS/Register/register[16][5] ), .A1(n4962), .B0(
        \i_MIPS/Register/register[24][5] ), .B1(n4958), .Y(n7348) );
  AO22XL U6335 ( .A0(n5001), .A1(n545), .B0(n4997), .B1(n2300), .Y(n8130) );
  AO22XL U6336 ( .A0(n5001), .A1(n546), .B0(n4997), .B1(n2301), .Y(n8121) );
  AO22XL U6337 ( .A0(n5001), .A1(n549), .B0(n4997), .B1(n2304), .Y(n8316) );
  AO22XL U6338 ( .A0(n5001), .A1(n510), .B0(n4997), .B1(n2262), .Y(n8307) );
  AO22XL U6339 ( .A0(n5001), .A1(n550), .B0(n4997), .B1(n2305), .Y(n8610) );
  AO22XL U6340 ( .A0(n5001), .A1(n511), .B0(n4997), .B1(n2263), .Y(n8219) );
  AO22XL U6341 ( .A0(n5001), .A1(n512), .B0(n4997), .B1(n2264), .Y(n8210) );
  AO22XL U6342 ( .A0(n5000), .A1(n206), .B0(n4996), .B1(n2306), .Y(n6336) );
  AO22XL U6343 ( .A0(n5001), .A1(n207), .B0(n4996), .B1(n2307), .Y(n6327) );
  AO22XL U6344 ( .A0(n5000), .A1(n208), .B0(n4996), .B1(n2308), .Y(n6184) );
  AO22XL U6345 ( .A0(n5000), .A1(n209), .B0(n4996), .B1(n2309), .Y(n6175) );
  AO22XL U6346 ( .A0(n5000), .A1(n210), .B0(n4996), .B1(n2310), .Y(n6834) );
  AO22XL U6347 ( .A0(n5000), .A1(n211), .B0(n4996), .B1(n2311), .Y(n6825) );
  AO22XL U6348 ( .A0(n5001), .A1(n212), .B0(n4996), .B1(n2312), .Y(n6754) );
  AO22XL U6349 ( .A0(n5000), .A1(n213), .B0(n4996), .B1(n2313), .Y(n6745) );
  OA22XL U6350 ( .A0(net112665), .A1(n1507), .B0(net112563), .B1(n3120), .Y(
        n8109) );
  OA22XL U6351 ( .A0(net112673), .A1(n815), .B0(net112571), .B1(n2347), .Y(
        n9248) );
  OA22XL U6352 ( .A0(net112671), .A1(n816), .B0(net112569), .B1(n2348), .Y(
        n9240) );
  OA22XL U6353 ( .A0(\i_MIPS/Register/register[1][20] ), .A1(n4834), .B0(
        \i_MIPS/Register/register[9][20] ), .B1(n4829), .Y(n8564) );
  OA22XL U6354 ( .A0(\i_MIPS/Register/register[23][27] ), .A1(n4884), .B0(
        \i_MIPS/Register/register[31][27] ), .B1(n4876), .Y(n8629) );
  OA22XL U6355 ( .A0(n5346), .A1(n2565), .B0(n5302), .B1(n794), .Y(n9817) );
  OA22XL U6356 ( .A0(n5346), .A1(n1189), .B0(n5302), .B1(n2761), .Y(n9812) );
  OA22XL U6357 ( .A0(n5337), .A1(n1190), .B0(n5293), .B1(n2762), .Y(n9438) );
  OA22XL U6358 ( .A0(n5341), .A1(n749), .B0(n5297), .B1(n2327), .Y(n9637) );
  OA22XL U6359 ( .A0(n5341), .A1(n750), .B0(n5297), .B1(n2328), .Y(n9632) );
  OA22XL U6360 ( .A0(n5336), .A1(n1191), .B0(n5292), .B1(n2763), .Y(n9418) );
  OA22XL U6361 ( .A0(n5336), .A1(n1192), .B0(n5292), .B1(n2764), .Y(n9414) );
  OA22XL U6362 ( .A0(n5336), .A1(n1193), .B0(n5292), .B1(n2765), .Y(n9409) );
  OA22XL U6363 ( .A0(n5338), .A1(n751), .B0(n5294), .B1(n2329), .Y(n9465) );
  OA22XL U6364 ( .A0(n5337), .A1(n752), .B0(n5293), .B1(n2330), .Y(n9460) );
  OA22XL U6365 ( .A0(n5337), .A1(n753), .B0(n5293), .B1(n2331), .Y(n9455) );
  OA22XL U6366 ( .A0(n5335), .A1(n754), .B0(n5291), .B1(n2332), .Y(n9374) );
  OA22XL U6367 ( .A0(n5349), .A1(n817), .B0(n5305), .B1(n2349), .Y(n9934) );
  OA22XL U6368 ( .A0(net112069), .A1(n1508), .B0(net111945), .B1(n3121), .Y(
        n8203) );
  OA22XL U6369 ( .A0(net112073), .A1(n1509), .B0(net111949), .B1(n3122), .Y(
        n8594) );
  OA22XL U6370 ( .A0(net112069), .A1(n1510), .B0(net111945), .B1(n3123), .Y(
        n8300) );
  OA22XL U6371 ( .A0(net112069), .A1(n1511), .B0(net111945), .B1(n3124), .Y(
        n8296) );
  OA22XL U6372 ( .A0(net112079), .A1(n1513), .B0(net111955), .B1(n3126), .Y(
        n8961) );
  OA22XL U6373 ( .A0(net112077), .A1(n1514), .B0(net111953), .B1(n3127), .Y(
        n8847) );
  OA22XL U6374 ( .A0(net112079), .A1(n1515), .B0(net111955), .B1(n3128), .Y(
        n8965) );
  OA22XL U6375 ( .A0(net112079), .A1(n1516), .B0(net111955), .B1(n3129), .Y(
        n8957) );
  OA22XL U6376 ( .A0(net112077), .A1(n1517), .B0(net111953), .B1(n3130), .Y(
        n8770) );
  OA22XL U6377 ( .A0(net112075), .A1(n1518), .B0(net111951), .B1(n3131), .Y(
        n8762) );
  OA22XL U6378 ( .A0(net112069), .A1(n1519), .B0(net111945), .B1(n3132), .Y(
        n8288) );
  OA22XL U6379 ( .A0(net112067), .A1(n1520), .B0(net111943), .B1(n3133), .Y(
        n8191) );
  OA22XL U6380 ( .A0(net112071), .A1(n1521), .B0(net111947), .B1(n3134), .Y(
        n8393) );
  OA22XL U6381 ( .A0(net112071), .A1(n1522), .B0(net111947), .B1(n3135), .Y(
        n8385) );
  OA22XL U6382 ( .A0(net112073), .A1(n1523), .B0(net111949), .B1(n3136), .Y(
        n8586) );
  OA22XL U6383 ( .A0(net112067), .A1(n2859), .B0(net111943), .B1(n1230), .Y(
        n8110) );
  OA22XL U6384 ( .A0(net112067), .A1(n1524), .B0(net111943), .B1(n3137), .Y(
        n8102) );
  OA22XL U6385 ( .A0(net112073), .A1(n1525), .B0(net111949), .B1(n3138), .Y(
        n8590) );
  OA22XL U6386 ( .A0(net112063), .A1(n1526), .B0(net111939), .B1(n3139), .Y(
        n7815) );
  OA22XL U6387 ( .A0(net112063), .A1(n1527), .B0(net111939), .B1(n3140), .Y(
        n7807) );
  OA22XL U6388 ( .A0(net112071), .A1(n1528), .B0(net111947), .B1(n3141), .Y(
        n8476) );
  OA22XL U6389 ( .A0(net112065), .A1(n1529), .B0(net111941), .B1(n3142), .Y(
        n8017) );
  OA22XL U6390 ( .A0(net112065), .A1(n1530), .B0(net111941), .B1(n3143), .Y(
        n8009) );
  OA22XL U6391 ( .A0(\i_MIPS/Register/register[22][18] ), .A1(n4912), .B0(
        \i_MIPS/Register/register[30][18] ), .B1(n4906), .Y(n7905) );
  OA22XL U6392 ( .A0(\i_MIPS/Register/register[22][26] ), .A1(n4913), .B0(
        \i_MIPS/Register/register[30][26] ), .B1(n4907), .Y(n8377) );
  OA22XL U6393 ( .A0(\i_MIPS/Register/register[6][26] ), .A1(n4913), .B0(
        \i_MIPS/Register/register[14][26] ), .B1(n4907), .Y(n8368) );
  OA22XL U6394 ( .A0(\i_MIPS/Register/register[22][17] ), .A1(n4912), .B0(
        \i_MIPS/Register/register[30][17] ), .B1(n4906), .Y(n7749) );
  OA22XL U6395 ( .A0(\i_MIPS/Register/register[6][17] ), .A1(n4912), .B0(
        \i_MIPS/Register/register[14][17] ), .B1(n4906), .Y(n7740) );
  OA22XL U6396 ( .A0(\i_MIPS/Register/register[22][21] ), .A1(n4913), .B0(
        \i_MIPS/Register/register[30][21] ), .B1(n4907), .Y(n8060) );
  OA22XL U6397 ( .A0(\i_MIPS/Register/register[22][23] ), .A1(n4913), .B0(
        \i_MIPS/Register/register[30][23] ), .B1(n4907), .Y(n8242) );
  OA22XL U6398 ( .A0(\i_MIPS/Register/register[22][27] ), .A1(n4913), .B0(
        \i_MIPS/Register/register[30][27] ), .B1(n4907), .Y(n8633) );
  OA22XL U6399 ( .A0(\i_MIPS/Register/register[22][4] ), .A1(n4911), .B0(
        \i_MIPS/Register/register[30][4] ), .B1(n4903), .Y(n7386) );
  OA22XL U6400 ( .A0(\i_MIPS/Register/register[22][19] ), .A1(n4912), .B0(
        \i_MIPS/Register/register[30][19] ), .B1(n4906), .Y(n7765) );
  OA22XL U6401 ( .A0(\i_MIPS/Register/register[6][23] ), .A1(n4938), .B0(
        \i_MIPS/Register/register[14][23] ), .B1(n4931), .Y(n8306) );
  OA22XL U6402 ( .A0(\i_MIPS/Register/register[22][23] ), .A1(n4938), .B0(
        \i_MIPS/Register/register[30][23] ), .B1(n4931), .Y(n8315) );
  OA22XL U6403 ( .A0(\i_MIPS/Register/register[22][3] ), .A1(n4914), .B0(
        \i_MIPS/Register/register[30][3] ), .B1(n4908), .Y(n8755) );
  AO21XL U6404 ( .A0(\i_MIPS/ID_EX[102] ), .A1(n5515), .B0(n4499), .Y(
        \i_MIPS/n483 ) );
  OA22XL U6405 ( .A0(\i_MIPS/Register/register[4][25] ), .A1(n4954), .B0(
        \i_MIPS/Register/register[12][25] ), .B1(n4950), .Y(n8501) );
  MX2XL U6406 ( .A(\D_cache/cache[7][142] ), .B(n10682), .S0(net111885), .Y(
        \D_cache/n653 ) );
  XNOR2X4 U6407 ( .A(n5587), .B(\i_MIPS/Reg_W[4] ), .Y(n6301) );
  NOR2XL U6408 ( .A(\i_MIPS/Reg_W[4] ), .B(\i_MIPS/Reg_W[3] ), .Y(
        \i_MIPS/forward_unit/n25 ) );
  NAND2X8 U6409 ( .A(n8821), .B(\i_MIPS/ALU/N303 ), .Y(n4501) );
  MX2XL U6410 ( .A(n3524), .B(\i_MIPS/Sign_Extend_ID[6] ), .S0(n5507), .Y(
        \i_MIPS/n506 ) );
  MX2XL U6411 ( .A(\D_cache/cache[7][29] ), .B(n4254), .S0(net111867), .Y(
        \D_cache/n1557 ) );
  MX2XL U6412 ( .A(\D_cache/cache[7][28] ), .B(n4255), .S0(net111871), .Y(
        \D_cache/n1565 ) );
  MX2XL U6413 ( .A(\D_cache/cache[7][27] ), .B(n4256), .S0(net111865), .Y(
        \D_cache/n1573 ) );
  MX2XL U6414 ( .A(\D_cache/cache[7][26] ), .B(n4257), .S0(net111871), .Y(
        \D_cache/n1581 ) );
  MX2XL U6415 ( .A(\D_cache/cache[7][25] ), .B(n10425), .S0(net111883), .Y(
        \D_cache/n1589 ) );
  MX2XL U6416 ( .A(\D_cache/cache[7][19] ), .B(n4261), .S0(net111883), .Y(
        \D_cache/n1637 ) );
  MX2XL U6417 ( .A(\D_cache/cache[7][16] ), .B(n4263), .S0(net111865), .Y(
        \D_cache/n1661 ) );
  MX2XL U6418 ( .A(\D_cache/cache[7][15] ), .B(n10188), .S0(net111871), .Y(
        \D_cache/n1669 ) );
  MX2XL U6419 ( .A(\D_cache/cache[7][14] ), .B(n10437), .S0(net111865), .Y(
        \D_cache/n1677 ) );
  MX2XL U6420 ( .A(\D_cache/cache[7][61] ), .B(n4267), .S0(net111867), .Y(
        \D_cache/n1301 ) );
  MX2XL U6421 ( .A(\D_cache/cache[7][60] ), .B(n10400), .S0(net111871), .Y(
        \D_cache/n1309 ) );
  MX2XL U6422 ( .A(\D_cache/cache[7][59] ), .B(n4268), .S0(net111871), .Y(
        \D_cache/n1317 ) );
  MX2XL U6423 ( .A(\D_cache/cache[7][58] ), .B(n4269), .S0(net111871), .Y(
        \D_cache/n1325 ) );
  MX2XL U6424 ( .A(\D_cache/cache[7][57] ), .B(n4270), .S0(net111865), .Y(
        \D_cache/n1333 ) );
  MX2XL U6425 ( .A(\D_cache/cache[7][51] ), .B(n4274), .S0(net111877), .Y(
        \D_cache/n1381 ) );
  MX2XL U6426 ( .A(\D_cache/cache[7][48] ), .B(n4275), .S0(net111865), .Y(
        \D_cache/n1405 ) );
  MX2XL U6427 ( .A(\D_cache/cache[7][47] ), .B(n4276), .S0(net111871), .Y(
        \D_cache/n1413 ) );
  MX2XL U6428 ( .A(\D_cache/cache[7][46] ), .B(n4277), .S0(net111865), .Y(
        \D_cache/n1421 ) );
  MX2XL U6429 ( .A(\D_cache/cache[7][35] ), .B(n4281), .S0(net111867), .Y(
        \D_cache/n1509 ) );
  MX2XL U6430 ( .A(\D_cache/cache[7][94] ), .B(n4283), .S0(net111885), .Y(
        \D_cache/n1037 ) );
  MX2XL U6431 ( .A(\D_cache/cache[7][93] ), .B(n4284), .S0(net111867), .Y(
        \D_cache/n1045 ) );
  MX2XL U6432 ( .A(\D_cache/cache[7][92] ), .B(n4285), .S0(net111871), .Y(
        \D_cache/n1053 ) );
  MX2XL U6433 ( .A(\D_cache/cache[7][91] ), .B(n4286), .S0(net111867), .Y(
        \D_cache/n1061 ) );
  MX2XL U6434 ( .A(\D_cache/cache[7][90] ), .B(n4287), .S0(net111883), .Y(
        \D_cache/n1069 ) );
  MX2XL U6435 ( .A(\D_cache/cache[7][89] ), .B(n4288), .S0(net111865), .Y(
        \D_cache/n1077 ) );
  MX2XL U6436 ( .A(\D_cache/cache[7][88] ), .B(n4289), .S0(net111879), .Y(
        \D_cache/n1085 ) );
  MX2XL U6437 ( .A(\D_cache/cache[7][87] ), .B(n4290), .S0(net111879), .Y(
        \D_cache/n1093 ) );
  MX2XL U6438 ( .A(\D_cache/cache[7][86] ), .B(n4291), .S0(net111877), .Y(
        \D_cache/n1101 ) );
  MX2XL U6439 ( .A(\D_cache/cache[7][85] ), .B(n4292), .S0(net111877), .Y(
        \D_cache/n1109 ) );
  MX2XL U6440 ( .A(\D_cache/cache[7][84] ), .B(n4293), .S0(net111877), .Y(
        \D_cache/n1117 ) );
  MX2XL U6441 ( .A(\D_cache/cache[7][83] ), .B(n4294), .S0(net111877), .Y(
        \D_cache/n1125 ) );
  MX2XL U6442 ( .A(\D_cache/cache[7][82] ), .B(n4295), .S0(net111873), .Y(
        \D_cache/n1133 ) );
  MX2XL U6443 ( .A(\D_cache/cache[7][81] ), .B(n10606), .S0(net111877), .Y(
        \D_cache/n1141 ) );
  MX2XL U6444 ( .A(\D_cache/cache[7][80] ), .B(n4296), .S0(net111865), .Y(
        \D_cache/n1149 ) );
  MX2XL U6445 ( .A(\D_cache/cache[7][79] ), .B(n4297), .S0(net111871), .Y(
        \D_cache/n1157 ) );
  MX2XL U6446 ( .A(\D_cache/cache[7][78] ), .B(n4298), .S0(net111865), .Y(
        \D_cache/n1165 ) );
  MX2XL U6447 ( .A(\D_cache/cache[7][74] ), .B(n10594), .S0(net111879), .Y(
        \D_cache/n1197 ) );
  MX2XL U6448 ( .A(\D_cache/cache[7][73] ), .B(n4299), .S0(net111867), .Y(
        \D_cache/n1205 ) );
  MX2XL U6449 ( .A(\D_cache/cache[7][71] ), .B(n4300), .S0(net111885), .Y(
        \D_cache/n1221 ) );
  MX2XL U6450 ( .A(\D_cache/cache[7][70] ), .B(n4282), .S0(net111883), .Y(
        \D_cache/n1229 ) );
  MX2XL U6451 ( .A(\D_cache/cache[7][69] ), .B(n4301), .S0(net111865), .Y(
        \D_cache/n1237 ) );
  MX2XL U6452 ( .A(\D_cache/cache[7][67] ), .B(n4302), .S0(net111867), .Y(
        \D_cache/n1253 ) );
  MX2XL U6453 ( .A(\D_cache/cache[7][126] ), .B(n4303), .S0(net111885), .Y(
        \D_cache/n781 ) );
  MX2XL U6454 ( .A(\D_cache/cache[7][125] ), .B(n4304), .S0(net111867), .Y(
        \D_cache/n789 ) );
  MX2XL U6455 ( .A(\D_cache/cache[7][124] ), .B(n10403), .S0(net111871), .Y(
        \D_cache/n797 ) );
  MX2XL U6456 ( .A(\D_cache/cache[7][123] ), .B(n4305), .S0(net111867), .Y(
        \D_cache/n805 ) );
  MX2XL U6457 ( .A(\D_cache/cache[7][122] ), .B(n4306), .S0(net111871), .Y(
        \D_cache/n813 ) );
  MX2XL U6458 ( .A(\D_cache/cache[7][121] ), .B(n4307), .S0(net111865), .Y(
        \D_cache/n821 ) );
  MX2XL U6459 ( .A(\D_cache/cache[7][120] ), .B(n4308), .S0(net111879), .Y(
        \D_cache/n829 ) );
  MX2XL U6460 ( .A(\D_cache/cache[7][119] ), .B(n4309), .S0(net111871), .Y(
        \D_cache/n837 ) );
  MX2XL U6461 ( .A(\D_cache/cache[7][118] ), .B(n4310), .S0(net111877), .Y(
        \D_cache/n845 ) );
  MX2XL U6462 ( .A(\D_cache/cache[7][117] ), .B(n4311), .S0(net111877), .Y(
        \D_cache/n853 ) );
  MX2XL U6463 ( .A(\D_cache/cache[7][116] ), .B(n4312), .S0(net111877), .Y(
        \D_cache/n861 ) );
  MX2XL U6464 ( .A(\D_cache/cache[7][115] ), .B(n10180), .S0(net111877), .Y(
        \D_cache/n869 ) );
  MX2XL U6465 ( .A(\D_cache/cache[7][114] ), .B(n4313), .S0(net111873), .Y(
        \D_cache/n877 ) );
  MX2XL U6466 ( .A(\D_cache/cache[7][113] ), .B(n4314), .S0(net111879), .Y(
        \D_cache/n885 ) );
  MX2XL U6467 ( .A(\D_cache/cache[7][112] ), .B(n4315), .S0(net111865), .Y(
        \D_cache/n893 ) );
  MX2XL U6468 ( .A(\D_cache/cache[7][111] ), .B(n10194), .S0(net111871), .Y(
        \D_cache/n901 ) );
  MX2XL U6469 ( .A(\D_cache/cache[7][110] ), .B(n10443), .S0(net111865), .Y(
        \D_cache/n909 ) );
  MX2XL U6470 ( .A(\D_cache/cache[7][106] ), .B(n10591), .S0(net111879), .Y(
        \D_cache/n941 ) );
  MX2XL U6471 ( .A(\D_cache/cache[7][105] ), .B(n4316), .S0(net111885), .Y(
        \D_cache/n949 ) );
  MX2XL U6472 ( .A(\D_cache/cache[7][103] ), .B(n10746), .S0(net111885), .Y(
        \D_cache/n965 ) );
  MX2XL U6473 ( .A(\D_cache/cache[7][101] ), .B(n10760), .S0(net111879), .Y(
        \D_cache/n981 ) );
  MX2XL U6474 ( .A(\D_cache/cache[7][99] ), .B(n4317), .S0(net111867), .Y(
        \D_cache/n997 ) );
  MX2XL U6475 ( .A(\D_cache/cache[7][30] ), .B(n4253), .S0(net111885), .Y(
        \D_cache/n1549 ) );
  MX2XL U6476 ( .A(\D_cache/cache[7][24] ), .B(n4258), .S0(net111879), .Y(
        \D_cache/n1597 ) );
  MX2XL U6477 ( .A(\D_cache/cache[7][23] ), .B(n4259), .S0(net111877), .Y(
        \D_cache/n1605 ) );
  MX2XL U6478 ( .A(\D_cache/cache[7][22] ), .B(n4260), .S0(net111877), .Y(
        \D_cache/n1613 ) );
  MX2XL U6479 ( .A(\D_cache/cache[7][21] ), .B(n10534), .S0(net111877), .Y(
        \D_cache/n1621 ) );
  MX2XL U6480 ( .A(\D_cache/cache[7][20] ), .B(n10522), .S0(net111867), .Y(
        \D_cache/n1629 ) );
  MX2XL U6481 ( .A(\D_cache/cache[7][18] ), .B(n4262), .S0(net111873), .Y(
        \D_cache/n1645 ) );
  MX2XL U6482 ( .A(\D_cache/cache[7][17] ), .B(n10597), .S0(net111879), .Y(
        \D_cache/n1653 ) );
  MX2XL U6483 ( .A(\D_cache/cache[7][10] ), .B(n4264), .S0(net111879), .Y(
        \D_cache/n1709 ) );
  MX2XL U6484 ( .A(\D_cache/cache[7][9] ), .B(n10767), .S0(net111879), .Y(
        \D_cache/n1717 ) );
  MX2XL U6485 ( .A(\D_cache/cache[7][7] ), .B(n4265), .S0(net111885), .Y(
        \D_cache/n1733 ) );
  MX2XL U6486 ( .A(\D_cache/cache[7][62] ), .B(n4266), .S0(net111885), .Y(
        \D_cache/n1293 ) );
  MX2XL U6487 ( .A(\D_cache/cache[7][56] ), .B(n10574), .S0(net111879), .Y(
        \D_cache/n1341 ) );
  MX2XL U6488 ( .A(\D_cache/cache[7][55] ), .B(n4271), .S0(net111877), .Y(
        \D_cache/n1349 ) );
  MX2XL U6489 ( .A(\D_cache/cache[7][54] ), .B(n10549), .S0(net111877), .Y(
        \D_cache/n1357 ) );
  MX2XL U6490 ( .A(\D_cache/cache[7][52] ), .B(n4273), .S0(net111867), .Y(
        \D_cache/n1373 ) );
  MX2XL U6491 ( .A(\D_cache/cache[7][50] ), .B(n10613), .S0(net111873), .Y(
        \D_cache/n1389 ) );
  MX2XL U6492 ( .A(\D_cache/cache[7][49] ), .B(n10600), .S0(net111879), .Y(
        \D_cache/n1397 ) );
  MX2XL U6493 ( .A(\D_cache/cache[7][42] ), .B(n10588), .S0(net111879), .Y(
        \D_cache/n1453 ) );
  MX2XL U6494 ( .A(\D_cache/cache[7][41] ), .B(n4278), .S0(net111881), .Y(
        \D_cache/n1461 ) );
  MX2XL U6495 ( .A(\D_cache/cache[7][39] ), .B(n4279), .S0(net111885), .Y(
        \D_cache/n1477 ) );
  MX2XL U6496 ( .A(\D_cache/cache[7][37] ), .B(n4280), .S0(net111865), .Y(
        \D_cache/n1493 ) );
  MX2XL U6497 ( .A(\D_cache/cache[7][13] ), .B(n4232), .S0(net111881), .Y(
        \D_cache/n1685 ) );
  MX2XL U6498 ( .A(\D_cache/cache[7][12] ), .B(n4233), .S0(net111867), .Y(
        \D_cache/n1693 ) );
  MX2XL U6499 ( .A(\D_cache/cache[7][11] ), .B(n4234), .S0(net111865), .Y(
        \D_cache/n1701 ) );
  MX2XL U6500 ( .A(\D_cache/cache[7][8] ), .B(n10819), .S0(net111881), .Y(
        \D_cache/n1725 ) );
  MX2XL U6501 ( .A(\D_cache/cache[7][2] ), .B(n4235), .S0(net111883), .Y(
        \D_cache/n1773 ) );
  MX2XL U6502 ( .A(\D_cache/cache[7][1] ), .B(n10840), .S0(net111881), .Y(
        \D_cache/n1781 ) );
  MX2XL U6503 ( .A(\D_cache/cache[7][0] ), .B(n10853), .S0(net111883), .Y(
        \D_cache/n1796 ) );
  MX2XL U6504 ( .A(\D_cache/cache[7][45] ), .B(n4236), .S0(net111881), .Y(
        \D_cache/n1429 ) );
  MX2XL U6505 ( .A(\D_cache/cache[7][44] ), .B(n10794), .S0(net111885), .Y(
        \D_cache/n1437 ) );
  MX2XL U6506 ( .A(\D_cache/cache[7][43] ), .B(n4239), .S0(net111885), .Y(
        \D_cache/n1445 ) );
  MX2XL U6507 ( .A(\D_cache/cache[7][40] ), .B(n4237), .S0(net111881), .Y(
        \D_cache/n1469 ) );
  MX2XL U6508 ( .A(\D_cache/cache[7][34] ), .B(n4240), .S0(net111883), .Y(
        \D_cache/n1517 ) );
  MX2XL U6509 ( .A(\D_cache/cache[7][33] ), .B(n4238), .S0(net111881), .Y(
        \D_cache/n1525 ) );
  MX2XL U6510 ( .A(\D_cache/cache[7][32] ), .B(n10856), .S0(net111883), .Y(
        \D_cache/n1533 ) );
  MX2XL U6511 ( .A(\D_cache/cache[7][95] ), .B(n4245), .S0(net111873), .Y(
        \D_cache/n1029 ) );
  MX2XL U6512 ( .A(\D_cache/cache[7][77] ), .B(n4241), .S0(net111881), .Y(
        \D_cache/n1173 ) );
  MX2XL U6513 ( .A(\D_cache/cache[7][76] ), .B(n10800), .S0(net111881), .Y(
        \D_cache/n1181 ) );
  MX2XL U6514 ( .A(\D_cache/cache[7][75] ), .B(n4244), .S0(net111879), .Y(
        \D_cache/n1189 ) );
  MX2XL U6515 ( .A(\D_cache/cache[7][72] ), .B(n4242), .S0(net111881), .Y(
        \D_cache/n1213 ) );
  MX2XL U6516 ( .A(\D_cache/cache[7][66] ), .B(n4246), .S0(net111883), .Y(
        \D_cache/n1261 ) );
  MX2XL U6517 ( .A(\D_cache/cache[7][65] ), .B(n4243), .S0(net111883), .Y(
        \D_cache/n1269 ) );
  MX2XL U6518 ( .A(\D_cache/cache[7][64] ), .B(n10862), .S0(net111883), .Y(
        \D_cache/n1277 ) );
  MX2XL U6519 ( .A(\D_cache/cache[7][63] ), .B(n11208), .S0(net111883), .Y(
        \D_cache/n1285 ) );
  MX2XL U6520 ( .A(\D_cache/cache[7][31] ), .B(n4231), .S0(net111883), .Y(
        \D_cache/n1541 ) );
  MX2XL U6521 ( .A(\D_cache/cache[7][109] ), .B(n10809), .S0(net111881), .Y(
        \D_cache/n917 ) );
  MX2XL U6522 ( .A(\D_cache/cache[7][108] ), .B(n10797), .S0(net111881), .Y(
        \D_cache/n925 ) );
  MX2XL U6523 ( .A(\D_cache/cache[7][107] ), .B(n10785), .S0(net111881), .Y(
        \D_cache/n933 ) );
  MX2XL U6524 ( .A(\D_cache/cache[7][104] ), .B(n10825), .S0(net111881), .Y(
        \D_cache/n957 ) );
  MX2XL U6525 ( .A(\D_cache/cache[7][98] ), .B(n11177), .S0(net111883), .Y(
        \D_cache/n1005 ) );
  MX2XL U6526 ( .A(\D_cache/cache[7][97] ), .B(n10846), .S0(net111879), .Y(
        \D_cache/n1013 ) );
  MX2XL U6527 ( .A(\D_cache/cache[7][96] ), .B(n10859), .S0(net111883), .Y(
        \D_cache/n1021 ) );
  MX2XL U6528 ( .A(\D_cache/cache[7][127] ), .B(n11211), .S0(net111883), .Y(
        \D_cache/n773 ) );
  MX2XL U6529 ( .A(\D_cache/cache[7][6] ), .B(n4247), .S0(net111883), .Y(
        \D_cache/n1741 ) );
  MX2XL U6530 ( .A(\D_cache/cache[7][4] ), .B(n4248), .S0(net111881), .Y(
        \D_cache/n1757 ) );
  MX2XL U6531 ( .A(\D_cache/cache[7][3] ), .B(n10509), .S0(net111867), .Y(
        \D_cache/n1765 ) );
  MX2XL U6532 ( .A(\D_cache/cache[7][38] ), .B(n4249), .S0(net111871), .Y(
        \D_cache/n1485 ) );
  MX2XL U6533 ( .A(\D_cache/cache[7][36] ), .B(n4250), .S0(net111879), .Y(
        \D_cache/n1501 ) );
  MX2XL U6534 ( .A(\D_cache/cache[7][68] ), .B(n4251), .S0(net111877), .Y(
        \D_cache/n1245 ) );
  MX2XL U6535 ( .A(\D_cache/cache[7][102] ), .B(n10169), .S0(net111883), .Y(
        \D_cache/n973 ) );
  MX2XL U6536 ( .A(\D_cache/cache[7][100] ), .B(n4252), .S0(net111867), .Y(
        \D_cache/n989 ) );
  MX2XL U6537 ( .A(n3505), .B(n4638), .S0(n5508), .Y(\i_MIPS/n530 ) );
  MX2XL U6538 ( .A(\D_cache/cache[7][145] ), .B(n121), .S0(net111877), .Y(
        \D_cache/n629 ) );
  MX2XL U6539 ( .A(\D_cache/cache[7][150] ), .B(n119), .S0(net111871), .Y(
        \D_cache/n589 ) );
  MX2XL U6540 ( .A(\D_cache/cache[7][134] ), .B(n127), .S0(net111865), .Y(
        \D_cache/n717 ) );
  MX2XL U6541 ( .A(\D_cache/cache[7][132] ), .B(n145), .S0(net111877), .Y(
        \D_cache/n733 ) );
  MX2XL U6542 ( .A(\D_cache/cache[7][149] ), .B(n120), .S0(net111871), .Y(
        \D_cache/n597 ) );
  MX2XL U6543 ( .A(\D_cache/cache[7][147] ), .B(n122), .S0(net111871), .Y(
        \D_cache/n613 ) );
  MX2XL U6544 ( .A(\D_cache/cache[7][151] ), .B(n132), .S0(net111871), .Y(
        \D_cache/n581 ) );
  MX2XL U6545 ( .A(\D_cache/cache[7][135] ), .B(n130), .S0(net111865), .Y(
        \D_cache/n709 ) );
  MX2XL U6546 ( .A(\D_cache/cache[7][137] ), .B(n136), .S0(net111871), .Y(
        \D_cache/n693 ) );
  MX2XL U6547 ( .A(\D_cache/cache[7][148] ), .B(n144), .S0(net111885), .Y(
        \D_cache/n605 ) );
  MX2XL U6548 ( .A(\D_cache/cache[7][138] ), .B(n129), .S0(net111865), .Y(
        \D_cache/n685 ) );
  MX2XL U6549 ( .A(\D_cache/cache[7][133] ), .B(n123), .S0(net111885), .Y(
        \D_cache/n725 ) );
  MX2XL U6550 ( .A(\D_cache/cache[7][129] ), .B(n137), .S0(net111885), .Y(
        \D_cache/n757 ) );
  MX2XL U6551 ( .A(\D_cache/cache[7][152] ), .B(n126), .S0(net111873), .Y(
        \D_cache/n573 ) );
  MX2XL U6552 ( .A(\D_cache/cache[7][143] ), .B(n143), .S0(net111873), .Y(
        \D_cache/n645 ) );
  MX2XL U6553 ( .A(\D_cache/cache[7][141] ), .B(n125), .S0(net111873), .Y(
        \D_cache/n661 ) );
  MX2XL U6554 ( .A(\D_cache/cache[7][128] ), .B(n118), .S0(net111873), .Y(
        \D_cache/n765 ) );
  MX2XL U6555 ( .A(\D_cache/cache[7][136] ), .B(n142), .S0(net111873), .Y(
        \D_cache/n701 ) );
  NAND2XL U6556 ( .A(n12950), .B(\i_MIPS/n336 ), .Y(net99637) );
  NAND2XL U6557 ( .A(n12959), .B(net113087), .Y(net99037) );
  NAND2XL U6558 ( .A(n12946), .B(\i_MIPS/n336 ), .Y(net99359) );
  NAND2XL U6559 ( .A(n12943), .B(\i_MIPS/n336 ), .Y(net99536) );
  NAND2XL U6560 ( .A(n12944), .B(net113089), .Y(n10409) );
  NAND2XL U6561 ( .A(n12948), .B(net113089), .Y(net99405) );
  NAND2XL U6562 ( .A(n9366), .B(ICACHE_addr[13]), .Y(n9367) );
  OA22XL U6563 ( .A0(\i_MIPS/Register/register[6][5] ), .A1(n4911), .B0(
        \i_MIPS/Register/register[14][5] ), .B1(n4903), .Y(n7298) );
  OA22XL U6564 ( .A0(\i_MIPS/Register/register[6][7] ), .A1(n4911), .B0(
        \i_MIPS/Register/register[14][7] ), .B1(n4903), .Y(n7506) );
  OA22XL U6565 ( .A0(\i_MIPS/Register/register[6][8] ), .A1(n4909), .B0(
        \i_MIPS/Register/register[14][8] ), .B1(n4906), .Y(n6807) );
  OA22XL U6566 ( .A0(\i_MIPS/Register/register[6][29] ), .A1(n4911), .B0(
        \i_MIPS/Register/register[14][29] ), .B1(n4906), .Y(n6728) );
  OA22XL U6567 ( .A0(\i_MIPS/Register/register[6][15] ), .A1(n4911), .B0(
        \i_MIPS/Register/register[14][15] ), .B1(n4903), .Y(n7073) );
  OA22XL U6568 ( .A0(\i_MIPS/Register/register[6][19] ), .A1(n4937), .B0(
        \i_MIPS/Register/register[14][19] ), .B1(n4930), .Y(n7826) );
  OAI221XL U6569 ( .A0(\i_MIPS/ALUin1[21] ), .A1(n4825), .B0(
        \i_MIPS/ALUin1[22] ), .B1(n4816), .C0(n8885), .Y(n8997) );
  OAI221XL U6570 ( .A0(\i_MIPS/ALUin1[24] ), .A1(n4824), .B0(
        \i_MIPS/ALUin1[25] ), .B1(n4816), .C0(n8640), .Y(n9136) );
  OAI221XL U6571 ( .A0(\i_MIPS/ALUin1[7] ), .A1(n4825), .B0(\i_MIPS/ALUin1[6] ), .B1(n4817), .C0(n6417), .Y(n7367) );
  OAI221XL U6572 ( .A0(\i_MIPS/ALUin1[9] ), .A1(n4824), .B0(\i_MIPS/ALUin1[8] ), .B1(n4816), .C0(n7556), .Y(n8816) );
  CLKBUFX3 U6573 ( .A(\i_MIPS/IR_ID[25] ), .Y(n5587) );
  OA22XL U6574 ( .A0(\i_MIPS/Register/register[4][31] ), .A1(n4953), .B0(
        \i_MIPS/Register/register[12][31] ), .B1(n4950), .Y(n9197) );
  OA22XL U6575 ( .A0(\i_MIPS/Register/register[0][31] ), .A1(n4963), .B0(
        \i_MIPS/Register/register[8][31] ), .B1(n4957), .Y(n9196) );
  OA22XL U6576 ( .A0(\i_MIPS/Register/register[4][30] ), .A1(n4952), .B0(
        \i_MIPS/Register/register[12][30] ), .B1(n4950), .Y(n9304) );
  OA22XL U6577 ( .A0(\i_MIPS/Register/register[0][30] ), .A1(n4963), .B0(
        \i_MIPS/Register/register[8][30] ), .B1(n4957), .Y(n9303) );
  OA22XL U6578 ( .A0(\i_MIPS/Register/register[5][6] ), .A1(n4851), .B0(
        \i_MIPS/Register/register[13][6] ), .B1(n4842), .Y(n7571) );
  OA22XL U6579 ( .A0(\i_MIPS/Register/register[7][6] ), .A1(n4883), .B0(
        \i_MIPS/Register/register[15][6] ), .B1(n4875), .Y(n7569) );
  OA22XL U6580 ( .A0(\i_MIPS/Register/register[1][6] ), .A1(n4834), .B0(
        \i_MIPS/Register/register[9][6] ), .B1(n4831), .Y(n7572) );
  OA22XL U6581 ( .A0(\i_MIPS/Register/register[1][14] ), .A1(n4832), .B0(
        \i_MIPS/Register/register[9][14] ), .B1(n4829), .Y(n6981) );
  OA22XL U6582 ( .A0(\i_MIPS/Register/register[1][9] ), .A1(n4832), .B0(
        \i_MIPS/Register/register[9][9] ), .B1(n4829), .Y(n6889) );
  OA22XL U6583 ( .A0(\i_MIPS/Register/register[7][7] ), .A1(n4882), .B0(
        \i_MIPS/Register/register[15][7] ), .B1(n4874), .Y(n7502) );
  OA22XL U6584 ( .A0(\i_MIPS/Register/register[1][7] ), .A1(n4833), .B0(
        \i_MIPS/Register/register[9][7] ), .B1(n4830), .Y(n7505) );
  OA22XL U6585 ( .A0(\i_MIPS/Register/register[1][13] ), .A1(n4832), .B0(
        \i_MIPS/Register/register[9][13] ), .B1(n4829), .Y(n6398) );
  OA22XL U6586 ( .A0(\i_MIPS/Register/register[5][21] ), .A1(n4850), .B0(
        \i_MIPS/Register/register[13][21] ), .B1(n4842), .Y(n8049) );
  OA22XL U6587 ( .A0(\i_MIPS/Register/register[7][21] ), .A1(n4883), .B0(
        \i_MIPS/Register/register[15][21] ), .B1(n4875), .Y(n8047) );
  OA22XL U6588 ( .A0(\i_MIPS/Register/register[1][21] ), .A1(n4835), .B0(
        \i_MIPS/Register/register[9][21] ), .B1(n4831), .Y(n8050) );
  OA22XL U6589 ( .A0(\i_MIPS/Register/register[1][4] ), .A1(n4833), .B0(
        \i_MIPS/Register/register[9][4] ), .B1(n4830), .Y(n7376) );
  OA22XL U6590 ( .A0(\i_MIPS/Register/register[1][11] ), .A1(n4833), .B0(
        \i_MIPS/Register/register[9][11] ), .B1(n4830), .Y(n7124) );
  OA22XL U6591 ( .A0(\i_MIPS/Register/register[7][5] ), .A1(n4882), .B0(
        \i_MIPS/Register/register[15][5] ), .B1(n4874), .Y(n7294) );
  OA22XL U6592 ( .A0(\i_MIPS/Register/register[1][8] ), .A1(n4832), .B0(
        \i_MIPS/Register/register[9][8] ), .B1(n4829), .Y(n6806) );
  OA22XL U6593 ( .A0(\i_MIPS/Register/register[1][29] ), .A1(n4832), .B0(
        \i_MIPS/Register/register[9][29] ), .B1(n4829), .Y(n6727) );
  OA22XL U6594 ( .A0(\i_MIPS/Register/register[5][15] ), .A1(n4849), .B0(
        \i_MIPS/Register/register[13][15] ), .B1(n4841), .Y(n7071) );
  OA22XL U6595 ( .A0(\i_MIPS/Register/register[7][15] ), .A1(n4882), .B0(
        \i_MIPS/Register/register[15][15] ), .B1(n4874), .Y(n7069) );
  OA22XL U6596 ( .A0(\i_MIPS/Register/register[1][15] ), .A1(n4833), .B0(
        \i_MIPS/Register/register[9][15] ), .B1(n4830), .Y(n7072) );
  OA22XL U6597 ( .A0(\i_MIPS/Register/register[5][12] ), .A1(n4848), .B0(
        \i_MIPS/Register/register[13][12] ), .B1(n4843), .Y(n6307) );
  OA22XL U6598 ( .A0(\i_MIPS/Register/register[7][12] ), .A1(n4881), .B0(
        \i_MIPS/Register/register[15][12] ), .B1(n4873), .Y(n6305) );
  OA22XL U6599 ( .A0(\i_MIPS/Register/register[1][12] ), .A1(n4832), .B0(
        \i_MIPS/Register/register[9][12] ), .B1(n4829), .Y(n6308) );
  OA22XL U6600 ( .A0(\i_MIPS/Register/register[20][31] ), .A1(n4954), .B0(
        \i_MIPS/Register/register[28][31] ), .B1(n4950), .Y(n9206) );
  OA22XL U6601 ( .A0(\i_MIPS/Register/register[16][31] ), .A1(n4961), .B0(
        \i_MIPS/Register/register[24][31] ), .B1(n4957), .Y(n9205) );
  OA22XL U6602 ( .A0(\i_MIPS/Register/register[20][30] ), .A1(n4953), .B0(
        \i_MIPS/Register/register[28][30] ), .B1(n4950), .Y(n9321) );
  OA22XL U6603 ( .A0(\i_MIPS/Register/register[16][30] ), .A1(n4962), .B0(
        \i_MIPS/Register/register[24][30] ), .B1(n4957), .Y(n9320) );
  NAND2XL U6604 ( .A(n10261), .B(ICACHE_addr[11]), .Y(n10262) );
  OA22XL U6605 ( .A0(net112679), .A1(n1531), .B0(net112577), .B1(n3144), .Y(
        n6963) );
  OA22XL U6606 ( .A0(net112679), .A1(n1532), .B0(net112577), .B1(n3145), .Y(
        n6883) );
  OA22XL U6607 ( .A0(net112679), .A1(n1533), .B0(net112577), .B1(n3146), .Y(
        n6800) );
  OA22XL U6608 ( .A0(net112679), .A1(n1534), .B0(net112577), .B1(n3147), .Y(
        n6792) );
  OA22XL U6609 ( .A0(net112657), .A1(n1536), .B0(net112573), .B1(n3149), .Y(
        n7491) );
  OA22XL U6610 ( .A0(\i_MIPS/Register/register[17][31] ), .A1(n4835), .B0(
        \i_MIPS/Register/register[25][31] ), .B1(n4831), .Y(n9113) );
  OA22XL U6611 ( .A0(\i_MIPS/Register/register[1][31] ), .A1(n4835), .B0(
        \i_MIPS/Register/register[9][31] ), .B1(n4829), .Y(n9104) );
  OA22XL U6612 ( .A0(\i_MIPS/Register/register[17][3] ), .A1(n4834), .B0(
        \i_MIPS/Register/register[25][3] ), .B1(n4831), .Y(n8754) );
  OA22XL U6613 ( .A0(\i_MIPS/Register/register[17][20] ), .A1(n4834), .B0(
        \i_MIPS/Register/register[25][20] ), .B1(n4831), .Y(n8573) );
  OA22XL U6614 ( .A0(\i_MIPS/Register/register[17][21] ), .A1(n4835), .B0(
        \i_MIPS/Register/register[25][21] ), .B1(n4831), .Y(n8059) );
  OA22XL U6615 ( .A0(\i_MIPS/Register/register[17][23] ), .A1(n4834), .B0(
        \i_MIPS/Register/register[25][23] ), .B1(n4830), .Y(n8241) );
  OA22XL U6616 ( .A0(\i_MIPS/Register/register[17][18] ), .A1(n4832), .B0(
        \i_MIPS/Register/register[25][18] ), .B1(n4831), .Y(n7904) );
  OA22XL U6617 ( .A0(\i_MIPS/Register/register[17][17] ), .A1(n4835), .B0(
        \i_MIPS/Register/register[25][17] ), .B1(n4831), .Y(n7748) );
  OA22XL U6618 ( .A0(\i_MIPS/Register/register[17][27] ), .A1(n4834), .B0(
        \i_MIPS/Register/register[25][27] ), .B1(n4831), .Y(n8632) );
  OA22XL U6619 ( .A0(\i_MIPS/Register/register[17][13] ), .A1(n4832), .B0(
        \i_MIPS/Register/register[25][13] ), .B1(n4829), .Y(n6407) );
  OA22XL U6620 ( .A0(\i_MIPS/Register/register[17][14] ), .A1(n4833), .B0(
        \i_MIPS/Register/register[25][14] ), .B1(n4830), .Y(n6990) );
  OA22XL U6621 ( .A0(\i_MIPS/Register/register[17][7] ), .A1(n4833), .B0(
        \i_MIPS/Register/register[25][7] ), .B1(n4830), .Y(n7514) );
  OA22XL U6622 ( .A0(\i_MIPS/Register/register[17][4] ), .A1(n4833), .B0(
        \i_MIPS/Register/register[25][4] ), .B1(n4830), .Y(n7385) );
  OA22XL U6623 ( .A0(\i_MIPS/Register/register[17][5] ), .A1(n4833), .B0(
        \i_MIPS/Register/register[25][5] ), .B1(n4830), .Y(n7306) );
  OA22XL U6624 ( .A0(\i_MIPS/Register/register[17][6] ), .A1(n4832), .B0(
        \i_MIPS/Register/register[25][6] ), .B1(n4831), .Y(n7581) );
  OA22XL U6625 ( .A0(\i_MIPS/Register/register[17][9] ), .A1(n4832), .B0(
        \i_MIPS/Register/register[25][9] ), .B1(n4829), .Y(n6898) );
  OA22XL U6626 ( .A0(\i_MIPS/Register/register[17][8] ), .A1(n4832), .B0(
        \i_MIPS/Register/register[25][8] ), .B1(n4829), .Y(n6815) );
  OA22XL U6627 ( .A0(\i_MIPS/Register/register[17][15] ), .A1(n4833), .B0(
        \i_MIPS/Register/register[25][15] ), .B1(n4830), .Y(n7081) );
  OA22XL U6628 ( .A0(\i_MIPS/Register/register[17][12] ), .A1(n4832), .B0(
        \i_MIPS/Register/register[25][12] ), .B1(n4829), .Y(n6317) );
  OA22XL U6629 ( .A0(\i_MIPS/Register/register[19][31] ), .A1(n4868), .B0(
        \i_MIPS/Register/register[27][31] ), .B1(n4858), .Y(n9111) );
  OA22XL U6630 ( .A0(\i_MIPS/Register/register[3][31] ), .A1(n4868), .B0(
        \i_MIPS/Register/register[11][31] ), .B1(n4858), .Y(n9102) );
  OA22XL U6631 ( .A0(\i_MIPS/Register/register[21][31] ), .A1(n4851), .B0(
        \i_MIPS/Register/register[29][31] ), .B1(n4844), .Y(n9112) );
  OA22XL U6632 ( .A0(\i_MIPS/Register/register[5][31] ), .A1(n4851), .B0(
        \i_MIPS/Register/register[13][31] ), .B1(n4844), .Y(n9103) );
  OA22XL U6633 ( .A0(\i_MIPS/Register/register[3][21] ), .A1(n4866), .B0(
        \i_MIPS/Register/register[11][21] ), .B1(n4858), .Y(n8048) );
  OA22XL U6634 ( .A0(\i_MIPS/Register/register[19][21] ), .A1(n4866), .B0(
        \i_MIPS/Register/register[27][21] ), .B1(n4856), .Y(n8057) );
  OA22XL U6635 ( .A0(\i_MIPS/Register/register[3][27] ), .A1(n4867), .B0(
        \i_MIPS/Register/register[11][27] ), .B1(n4857), .Y(n8621) );
  OA22XL U6636 ( .A0(\i_MIPS/Register/register[19][27] ), .A1(n4867), .B0(
        \i_MIPS/Register/register[27][27] ), .B1(n4857), .Y(n8630) );
  OA22XL U6637 ( .A0(\i_MIPS/Register/register[3][18] ), .A1(n4866), .B0(
        \i_MIPS/Register/register[11][18] ), .B1(n4856), .Y(n7893) );
  OA22XL U6638 ( .A0(\i_MIPS/Register/register[19][18] ), .A1(n4866), .B0(
        \i_MIPS/Register/register[27][18] ), .B1(n4855), .Y(n7902) );
  OA22XL U6639 ( .A0(\i_MIPS/Register/register[3][6] ), .A1(n4866), .B0(
        \i_MIPS/Register/register[11][6] ), .B1(n4857), .Y(n7570) );
  OA22XL U6640 ( .A0(\i_MIPS/Register/register[19][6] ), .A1(n4866), .B0(
        \i_MIPS/Register/register[27][6] ), .B1(n4856), .Y(n7579) );
  OA22XL U6641 ( .A0(\i_MIPS/Register/register[19][14] ), .A1(n4865), .B0(
        \i_MIPS/Register/register[27][14] ), .B1(n4856), .Y(n6988) );
  OA22XL U6642 ( .A0(\i_MIPS/Register/register[3][7] ), .A1(n4865), .B0(
        \i_MIPS/Register/register[11][7] ), .B1(n4856), .Y(n7503) );
  OA22XL U6643 ( .A0(\i_MIPS/Register/register[19][7] ), .A1(n4865), .B0(
        \i_MIPS/Register/register[27][7] ), .B1(n4856), .Y(n7512) );
  OA22XL U6644 ( .A0(\i_MIPS/Register/register[3][5] ), .A1(n4865), .B0(
        \i_MIPS/Register/register[11][5] ), .B1(n4856), .Y(n7295) );
  OA22XL U6645 ( .A0(\i_MIPS/Register/register[19][5] ), .A1(n4865), .B0(
        \i_MIPS/Register/register[27][5] ), .B1(n4856), .Y(n7304) );
  OA22XL U6646 ( .A0(\i_MIPS/Register/register[19][29] ), .A1(n4864), .B0(
        \i_MIPS/Register/register[27][29] ), .B1(n4855), .Y(n6734) );
  OA22XL U6647 ( .A0(\i_MIPS/Register/register[3][15] ), .A1(n4865), .B0(
        \i_MIPS/Register/register[11][15] ), .B1(n4856), .Y(n7070) );
  OA22XL U6648 ( .A0(\i_MIPS/Register/register[19][15] ), .A1(n4865), .B0(
        \i_MIPS/Register/register[27][15] ), .B1(n4856), .Y(n7079) );
  OA22XL U6649 ( .A0(\i_MIPS/Register/register[3][12] ), .A1(n4864), .B0(
        \i_MIPS/Register/register[11][12] ), .B1(n4855), .Y(n6306) );
  OA22XL U6650 ( .A0(\i_MIPS/Register/register[19][12] ), .A1(n4864), .B0(
        \i_MIPS/Register/register[27][12] ), .B1(n4855), .Y(n6315) );
  OA22XL U6651 ( .A0(\i_MIPS/Register/register[21][18] ), .A1(n4851), .B0(
        \i_MIPS/Register/register[29][18] ), .B1(n4842), .Y(n7903) );
  OA22XL U6652 ( .A0(\i_MIPS/Register/register[21][21] ), .A1(n4850), .B0(
        \i_MIPS/Register/register[29][21] ), .B1(n4842), .Y(n8058) );
  OA22XL U6653 ( .A0(\i_MIPS/Register/register[21][6] ), .A1(n4851), .B0(
        \i_MIPS/Register/register[29][6] ), .B1(n4842), .Y(n7580) );
  OA22XL U6654 ( .A0(\i_MIPS/Register/register[21][14] ), .A1(n4849), .B0(
        \i_MIPS/Register/register[29][14] ), .B1(n4841), .Y(n6989) );
  OA22XL U6655 ( .A0(\i_MIPS/Register/register[21][7] ), .A1(n4849), .B0(
        \i_MIPS/Register/register[29][7] ), .B1(n4841), .Y(n7513) );
  OA22XL U6656 ( .A0(\i_MIPS/Register/register[21][15] ), .A1(n4849), .B0(
        \i_MIPS/Register/register[29][15] ), .B1(n4841), .Y(n7080) );
  OA22XL U6657 ( .A0(\i_MIPS/Register/register[21][12] ), .A1(n4848), .B0(
        \i_MIPS/Register/register[29][12] ), .B1(n4843), .Y(n6316) );
  OA22XL U6658 ( .A0(net112681), .A1(n1537), .B0(net112565), .B1(n3150), .Y(
        n6380) );
  OA22XL U6659 ( .A0(net112681), .A1(n1538), .B0(net112577), .B1(n3151), .Y(
        n6284) );
  OA22XL U6660 ( .A0(\i_MIPS/Register/register[4][19] ), .A1(n4953), .B0(
        \i_MIPS/Register/register[12][19] ), .B1(n4949), .Y(n7833) );
  OA22XL U6661 ( .A0(\i_MIPS/Register/register[20][25] ), .A1(n4954), .B0(
        \i_MIPS/Register/register[28][25] ), .B1(n4950), .Y(n8510) );
  OA22XL U6662 ( .A0(\i_MIPS/Register/register[4][1] ), .A1(n4953), .B0(
        \i_MIPS/Register/register[12][1] ), .B1(n4949), .Y(n7597) );
  OA22XL U6663 ( .A0(\i_MIPS/Register/register[23][31] ), .A1(n4885), .B0(
        \i_MIPS/Register/register[31][31] ), .B1(n4877), .Y(n9110) );
  OA22XL U6664 ( .A0(\i_MIPS/Register/register[7][31] ), .A1(n4885), .B0(
        \i_MIPS/Register/register[15][31] ), .B1(n4877), .Y(n9101) );
  OA22XL U6665 ( .A0(\i_MIPS/Register/register[23][21] ), .A1(n4883), .B0(
        \i_MIPS/Register/register[31][21] ), .B1(n4875), .Y(n8056) );
  OA22XL U6666 ( .A0(\i_MIPS/Register/register[23][18] ), .A1(n4883), .B0(
        \i_MIPS/Register/register[31][18] ), .B1(n4875), .Y(n7901) );
  OA22XL U6667 ( .A0(\i_MIPS/Register/register[23][14] ), .A1(n4882), .B0(
        \i_MIPS/Register/register[31][14] ), .B1(n4874), .Y(n6987) );
  OA22XL U6668 ( .A0(\i_MIPS/Register/register[23][7] ), .A1(n4882), .B0(
        \i_MIPS/Register/register[31][7] ), .B1(n4874), .Y(n7511) );
  OA22XL U6669 ( .A0(\i_MIPS/Register/register[23][5] ), .A1(n4882), .B0(
        \i_MIPS/Register/register[31][5] ), .B1(n4874), .Y(n7303) );
  OA22XL U6670 ( .A0(\i_MIPS/Register/register[23][6] ), .A1(n4883), .B0(
        \i_MIPS/Register/register[31][6] ), .B1(n4875), .Y(n7578) );
  OA22XL U6671 ( .A0(\i_MIPS/Register/register[23][15] ), .A1(n4882), .B0(
        \i_MIPS/Register/register[31][15] ), .B1(n4874), .Y(n7078) );
  OA22XL U6672 ( .A0(\i_MIPS/Register/register[23][12] ), .A1(n4881), .B0(
        \i_MIPS/Register/register[31][12] ), .B1(n4873), .Y(n6314) );
  OA22XL U6673 ( .A0(\i_MIPS/Register/register[0][19] ), .A1(n4963), .B0(
        \i_MIPS/Register/register[8][19] ), .B1(n4959), .Y(n7832) );
  OA22XL U6674 ( .A0(\i_MIPS/Register/register[16][25] ), .A1(n4962), .B0(
        \i_MIPS/Register/register[24][25] ), .B1(n4959), .Y(n8509) );
  OA22XL U6675 ( .A0(\i_MIPS/Register/register[0][25] ), .A1(n4963), .B0(
        \i_MIPS/Register/register[8][25] ), .B1(n4959), .Y(n8500) );
  OA22XL U6676 ( .A0(\i_MIPS/Register/register[0][1] ), .A1(n4963), .B0(
        \i_MIPS/Register/register[8][1] ), .B1(n4958), .Y(n7596) );
  OA22XL U6677 ( .A0(\i_MIPS/Register/register[23][0] ), .A1(n6515), .B0(
        \i_MIPS/Register/register[31][0] ), .B1(n6514), .Y(n6516) );
  OA22XL U6678 ( .A0(\i_MIPS/Register/register[7][0] ), .A1(n6515), .B0(
        \i_MIPS/Register/register[15][0] ), .B1(n6514), .Y(n6499) );
  OA22XL U6679 ( .A0(n5339), .A1(n1194), .B0(n5295), .B1(n2766), .Y(n9519) );
  OA22XL U6680 ( .A0(n5342), .A1(n1195), .B0(n5298), .B1(n2767), .Y(n9661) );
  OA22XL U6681 ( .A0(n5341), .A1(n1196), .B0(n5297), .B1(n2768), .Y(n9656) );
  OA22XL U6682 ( .A0(n5335), .A1(n755), .B0(n5291), .B1(n2333), .Y(n9369) );
  OA22XL U6683 ( .A0(n5338), .A1(n2566), .B0(n5294), .B1(n795), .Y(n9489) );
  OA22XL U6684 ( .A0(n5338), .A1(n2567), .B0(n5294), .B1(n796), .Y(n9484) );
  OA22XL U6685 ( .A0(n5338), .A1(n2568), .B0(n5294), .B1(n797), .Y(n9474) );
  OA22XL U6686 ( .A0(n5340), .A1(n756), .B0(n5296), .B1(n2334), .Y(n9534) );
  OA22XL U6687 ( .A0(n5350), .A1(n1197), .B0(n5306), .B1(n2769), .Y(n9956) );
  OA22XL U6688 ( .A0(n5340), .A1(n757), .B0(n5296), .B1(n2335), .Y(n9529) );
  OA22XL U6689 ( .A0(n5341), .A1(n2569), .B0(n5297), .B1(n798), .Y(n9596) );
  OA22XL U6690 ( .A0(n5339), .A1(n1198), .B0(n5295), .B1(n2770), .Y(n9504) );
  OA22XL U6691 ( .A0(n5339), .A1(n2570), .B0(n5295), .B1(n799), .Y(n9494) );
  OA22XL U6692 ( .A0(n5339), .A1(n1199), .B0(n5295), .B1(n2771), .Y(n9499) );
  OA22XL U6693 ( .A0(n5336), .A1(n1200), .B0(n5292), .B1(n2772), .Y(n9404) );
  OA22XL U6694 ( .A0(n5335), .A1(n1201), .B0(n5291), .B1(n2773), .Y(n9394) );
  OA22XL U6695 ( .A0(n5335), .A1(n1202), .B0(n5291), .B1(n2774), .Y(n9389) );
  OA22XL U6696 ( .A0(n5353), .A1(n1203), .B0(n5309), .B1(n2775), .Y(n10097) );
  OA22XL U6697 ( .A0(n5353), .A1(n1204), .B0(n5309), .B1(n2776), .Y(n10087) );
  OA22XL U6698 ( .A0(n5349), .A1(n1205), .B0(n5305), .B1(n2777), .Y(n9951) );
  OA22XL U6699 ( .A0(net112041), .A1(n1539), .B0(net111917), .B1(n3152), .Y(
        n6277) );
  OA22XL U6700 ( .A0(net112041), .A1(n1540), .B0(net111917), .B1(n3153), .Y(
        n6269) );
  OA22XL U6701 ( .A0(net112055), .A1(n1541), .B0(net111931), .B1(n3154), .Y(
        n7393) );
  OA22XL U6702 ( .A0(net112053), .A1(n1542), .B0(net111929), .B1(n3155), .Y(
        n7235) );
  OA22XL U6703 ( .A0(net112053), .A1(n1543), .B0(net111929), .B1(n3156), .Y(
        n7239) );
  OA22XL U6704 ( .A0(net112053), .A1(n1544), .B0(net111929), .B1(n3157), .Y(
        n7231) );
  OA22XL U6705 ( .A0(net112055), .A1(n1545), .B0(net111931), .B1(n3158), .Y(
        n7319) );
  OA22XL U6706 ( .A0(net112055), .A1(n1546), .B0(net111931), .B1(n3159), .Y(
        n7323) );
  OA22XL U6707 ( .A0(net112055), .A1(n1547), .B0(net111931), .B1(n3160), .Y(
        n7315) );
  OA22XL U6708 ( .A0(net112047), .A1(n1548), .B0(net111923), .B1(n3161), .Y(
        n6785) );
  OA22XL U6709 ( .A0(net112061), .A1(n1549), .B0(net111937), .B1(n3162), .Y(
        n7645) );
  OA22XL U6710 ( .A0(net112061), .A1(n1550), .B0(net111937), .B1(n3163), .Y(
        n7641) );
  OA22XL U6711 ( .A0(net112045), .A1(n1551), .B0(net111921), .B1(n3164), .Y(
        n6535) );
  OA22XL U6712 ( .A0(net112045), .A1(n1552), .B0(net111921), .B1(n3165), .Y(
        n6714) );
  OA22XL U6713 ( .A0(net112045), .A1(n1553), .B0(net111921), .B1(n3166), .Y(
        n6706) );
  OA22XL U6714 ( .A0(net112057), .A1(n1554), .B0(net111933), .B1(n3167), .Y(
        n7484) );
  OA22XL U6715 ( .A0(net112059), .A1(n1555), .B0(net111935), .B1(n3168), .Y(
        net105047) );
  OA22XL U6716 ( .A0(net112081), .A1(n1556), .B0(net111957), .B1(n3169), .Y(
        n9087) );
  OA22XL U6717 ( .A0(net112081), .A1(n1557), .B0(net111957), .B1(n3170), .Y(
        n9091) );
  OA22XL U6718 ( .A0(net112081), .A1(n1558), .B0(net111957), .B1(n3171), .Y(
        n9083) );
  OA22XL U6719 ( .A0(\i_MIPS/Register/register[6][16] ), .A1(n4938), .B0(
        \i_MIPS/Register/register[14][16] ), .B1(n4931), .Y(n8209) );
  OA22XL U6720 ( .A0(\i_MIPS/Register/register[6][27] ), .A1(n4938), .B0(
        \i_MIPS/Register/register[14][27] ), .B1(n4931), .Y(n8691) );
  OA22XL U6721 ( .A0(\i_MIPS/Register/register[22][16] ), .A1(n4938), .B0(
        \i_MIPS/Register/register[30][16] ), .B1(n4931), .Y(n8218) );
  OA22XL U6722 ( .A0(\i_MIPS/Register/register[22][27] ), .A1(n4934), .B0(
        \i_MIPS/Register/register[30][27] ), .B1(n4931), .Y(n8700) );
  OA22XL U6723 ( .A0(\i_MIPS/Register/register[6][21] ), .A1(n4937), .B0(
        \i_MIPS/Register/register[14][21] ), .B1(n4930), .Y(n8120) );
  OA22XL U6724 ( .A0(\i_MIPS/Register/register[22][21] ), .A1(n4937), .B0(
        \i_MIPS/Register/register[30][21] ), .B1(n4931), .Y(n8129) );
  OA22XL U6725 ( .A0(\i_MIPS/Register/register[22][19] ), .A1(n4937), .B0(
        \i_MIPS/Register/register[30][19] ), .B1(n4930), .Y(n7835) );
  OA22XL U6726 ( .A0(\i_MIPS/Register/register[6][18] ), .A1(n4937), .B0(
        \i_MIPS/Register/register[14][18] ), .B1(n4930), .Y(n7930) );
  OA22XL U6727 ( .A0(\i_MIPS/Register/register[22][18] ), .A1(n4937), .B0(
        \i_MIPS/Register/register[30][18] ), .B1(n4930), .Y(n7939) );
  OA22XL U6728 ( .A0(\i_MIPS/Register/register[22][17] ), .A1(n4937), .B0(
        \i_MIPS/Register/register[30][17] ), .B1(n4930), .Y(n7682) );
  OA22XL U6729 ( .A0(\i_MIPS/Register/register[22][5] ), .A1(n4911), .B0(
        \i_MIPS/Register/register[30][5] ), .B1(n4903), .Y(n7307) );
  OA22XL U6730 ( .A0(\i_MIPS/Register/register[22][6] ), .A1(n4912), .B0(
        \i_MIPS/Register/register[30][6] ), .B1(n4906), .Y(n7582) );
  OA22XL U6731 ( .A0(\i_MIPS/Register/register[6][6] ), .A1(n4912), .B0(
        \i_MIPS/Register/register[14][6] ), .B1(n4906), .Y(n7573) );
  OA22XL U6732 ( .A0(\i_MIPS/Register/register[22][13] ), .A1(n4909), .B0(
        \i_MIPS/Register/register[30][13] ), .B1(n4903), .Y(n6408) );
  OA22XL U6733 ( .A0(\i_MIPS/Register/register[22][14] ), .A1(n4911), .B0(
        \i_MIPS/Register/register[30][14] ), .B1(n4903), .Y(n6991) );
  OA22XL U6734 ( .A0(\i_MIPS/Register/register[6][11] ), .A1(n4936), .B0(
        \i_MIPS/Register/register[14][11] ), .B1(n4930), .Y(n7159) );
  OA22XL U6735 ( .A0(\i_MIPS/Register/register[22][9] ), .A1(n4909), .B0(
        \i_MIPS/Register/register[30][9] ), .B1(n4906), .Y(n6899) );
  OA22XL U6736 ( .A0(\i_MIPS/Register/register[6][9] ), .A1(n4909), .B0(
        \i_MIPS/Register/register[14][9] ), .B1(n4903), .Y(n6890) );
  OA22XL U6737 ( .A0(\i_MIPS/Register/register[22][7] ), .A1(n4911), .B0(
        \i_MIPS/Register/register[30][7] ), .B1(n4903), .Y(n7515) );
  OA22XL U6738 ( .A0(\i_MIPS/Register/register[22][8] ), .A1(n4909), .B0(
        \i_MIPS/Register/register[30][8] ), .B1(n4903), .Y(n6816) );
  OA22XL U6739 ( .A0(\i_MIPS/Register/register[22][29] ), .A1(n4911), .B0(
        \i_MIPS/Register/register[30][29] ), .B1(n4906), .Y(n6737) );
  OA22XL U6740 ( .A0(\i_MIPS/Register/register[22][10] ), .A1(n4936), .B0(
        \i_MIPS/Register/register[30][10] ), .B1(n4930), .Y(n7258) );
  OA22XL U6741 ( .A0(\i_MIPS/Register/register[6][5] ), .A1(n4936), .B0(
        \i_MIPS/Register/register[14][5] ), .B1(n4930), .Y(n7333) );
  OA22XL U6742 ( .A0(\i_MIPS/Register/register[22][5] ), .A1(n4936), .B0(
        \i_MIPS/Register/register[30][5] ), .B1(n4930), .Y(n7342) );
  OA22XL U6743 ( .A0(\i_MIPS/Register/register[22][15] ), .A1(n4911), .B0(
        \i_MIPS/Register/register[30][15] ), .B1(n4903), .Y(n7082) );
  OA22XL U6744 ( .A0(\i_MIPS/Register/register[22][1] ), .A1(n4912), .B0(
        \i_MIPS/Register/register[30][1] ), .B1(n4906), .Y(n7660) );
  OA22XL U6745 ( .A0(\i_MIPS/Register/register[6][1] ), .A1(n4912), .B0(
        \i_MIPS/Register/register[14][1] ), .B1(n4906), .Y(n7651) );
  OA22XL U6746 ( .A0(\i_MIPS/Register/register[6][12] ), .A1(n4909), .B0(
        \i_MIPS/Register/register[14][12] ), .B1(n4906), .Y(n6309) );
  OA22XL U6747 ( .A0(\i_MIPS/Register/register[6][29] ), .A1(n4935), .B0(
        \i_MIPS/Register/register[14][29] ), .B1(n4929), .Y(n6686) );
  OA22XL U6748 ( .A0(\i_MIPS/Register/register[22][29] ), .A1(n4935), .B0(
        \i_MIPS/Register/register[30][29] ), .B1(n4929), .Y(n6695) );
  OA22XL U6749 ( .A0(\i_MIPS/Register/register[6][7] ), .A1(n4936), .B0(
        \i_MIPS/Register/register[14][7] ), .B1(n4930), .Y(n7431) );
  OA22XL U6750 ( .A0(\i_MIPS/Register/register[22][7] ), .A1(n4936), .B0(
        \i_MIPS/Register/register[30][7] ), .B1(n4930), .Y(n7440) );
  OA22XL U6751 ( .A0(\i_MIPS/Register/register[6][6] ), .A1(n4937), .B0(
        \i_MIPS/Register/register[14][6] ), .B1(n4930), .Y(n7523) );
  OA22XL U6752 ( .A0(\i_MIPS/Register/register[22][6] ), .A1(n4937), .B0(
        \i_MIPS/Register/register[30][6] ), .B1(n4930), .Y(n7532) );
  OA22XL U6753 ( .A0(\i_MIPS/Register/register[6][13] ), .A1(n4935), .B0(
        \i_MIPS/Register/register[14][13] ), .B1(n4929), .Y(n6326) );
  OA22XL U6754 ( .A0(\i_MIPS/Register/register[6][15] ), .A1(n4936), .B0(
        \i_MIPS/Register/register[14][15] ), .B1(n4929), .Y(n6999) );
  OA22XL U6755 ( .A0(\i_MIPS/Register/register[22][13] ), .A1(n4935), .B0(
        \i_MIPS/Register/register[30][13] ), .B1(n4929), .Y(n6335) );
  OA22XL U6756 ( .A0(\i_MIPS/Register/register[22][15] ), .A1(n4936), .B0(
        \i_MIPS/Register/register[30][15] ), .B1(n4929), .Y(n7008) );
  OA22XL U6757 ( .A0(\i_MIPS/Register/register[6][14] ), .A1(n4935), .B0(
        \i_MIPS/Register/register[14][14] ), .B1(n4929), .Y(n6907) );
  OA22XL U6758 ( .A0(\i_MIPS/Register/register[22][14] ), .A1(n4936), .B0(
        \i_MIPS/Register/register[30][14] ), .B1(n4930), .Y(n6916) );
  OA22XL U6759 ( .A0(\i_MIPS/Register/register[6][12] ), .A1(n4935), .B0(
        \i_MIPS/Register/register[14][12] ), .B1(n4929), .Y(n6174) );
  OA22XL U6760 ( .A0(\i_MIPS/Register/register[22][1] ), .A1(n4937), .B0(
        \i_MIPS/Register/register[30][1] ), .B1(n4930), .Y(n7599) );
  OA22XL U6761 ( .A0(\i_MIPS/Register/register[22][12] ), .A1(n4935), .B0(
        \i_MIPS/Register/register[30][12] ), .B1(n4929), .Y(n6183) );
  OA22XL U6762 ( .A0(\i_MIPS/Register/register[6][9] ), .A1(n4935), .B0(
        \i_MIPS/Register/register[14][9] ), .B1(n4929), .Y(n6824) );
  OA22XL U6763 ( .A0(\i_MIPS/Register/register[22][9] ), .A1(n4935), .B0(
        \i_MIPS/Register/register[30][9] ), .B1(n4929), .Y(n6833) );
  OA22XL U6764 ( .A0(\i_MIPS/Register/register[6][8] ), .A1(n4935), .B0(
        \i_MIPS/Register/register[14][8] ), .B1(n4929), .Y(n6744) );
  OA22XL U6765 ( .A0(\i_MIPS/Register/register[22][8] ), .A1(n4935), .B0(
        \i_MIPS/Register/register[30][8] ), .B1(n4929), .Y(n6753) );
  OA22XL U6766 ( .A0(\i_MIPS/Register/register[6][3] ), .A1(n4938), .B0(
        \i_MIPS/Register/register[14][3] ), .B1(n4932), .Y(n8780) );
  OA22XL U6767 ( .A0(\i_MIPS/Register/register[22][3] ), .A1(n4938), .B0(
        \i_MIPS/Register/register[30][3] ), .B1(n4932), .Y(n8789) );
  OA22XL U6768 ( .A0(\i_MIPS/Register/register[22][30] ), .A1(n4914), .B0(
        \i_MIPS/Register/register[30][30] ), .B1(n4908), .Y(n9222) );
  OA22XL U6769 ( .A0(\i_MIPS/Register/register[6][30] ), .A1(n4914), .B0(
        \i_MIPS/Register/register[14][30] ), .B1(n4908), .Y(n9213) );
  OA22XL U6770 ( .A0(\i_MIPS/Register/register[22][31] ), .A1(n4914), .B0(
        \i_MIPS/Register/register[30][31] ), .B1(n4908), .Y(n9114) );
  OA22XL U6771 ( .A0(\i_MIPS/Register/register[6][31] ), .A1(n4914), .B0(
        \i_MIPS/Register/register[14][31] ), .B1(n4908), .Y(n9105) );
  OA22XL U6772 ( .A0(\i_MIPS/Register/register[22][30] ), .A1(n4938), .B0(
        \i_MIPS/Register/register[30][30] ), .B1(n4932), .Y(n9306) );
  MX2XL U6773 ( .A(\I_cache/cache[7][142] ), .B(n11034), .S0(n5368), .Y(n11680) );
  MX2XL U6774 ( .A(\I_cache/cache[6][151] ), .B(n3512), .S0(n5410), .Y(n11609)
         );
  MX2XL U6775 ( .A(\I_cache/cache[3][151] ), .B(n3512), .S0(n5190), .Y(n11612)
         );
  MX2XL U6776 ( .A(\I_cache/cache[1][151] ), .B(n3512), .S0(n5103), .Y(n11614)
         );
  MX2XL U6777 ( .A(\I_cache/cache[2][139] ), .B(n10976), .S0(n5233), .Y(n11709) );
  MX2XL U6778 ( .A(\I_cache/cache[4][15] ), .B(n9351), .S0(n5321), .Y(n12699)
         );
  MX2XL U6779 ( .A(\I_cache/cache[7][128] ), .B(n10978), .S0(n5366), .Y(n11792) );
  MX2XL U6780 ( .A(\I_cache/cache[7][131] ), .B(n10994), .S0(n5367), .Y(n11768) );
  MX2XL U6781 ( .A(\I_cache/cache[2][131] ), .B(n10994), .S0(n5233), .Y(n11773) );
  MX2XL U6782 ( .A(\I_cache/cache[0][131] ), .B(n10994), .S0(n5146), .Y(n11775) );
  MX2XL U6783 ( .A(\I_cache/cache[7][130] ), .B(n10993), .S0(n5367), .Y(n11776) );
  MX2XL U6784 ( .A(\I_cache/cache[2][130] ), .B(n10993), .S0(n5233), .Y(n11781) );
  MX2XL U6785 ( .A(\I_cache/cache[0][130] ), .B(n10993), .S0(n5146), .Y(n11783) );
  MX2XL U6786 ( .A(\I_cache/cache[7][144] ), .B(n3514), .S0(n5366), .Y(n11664)
         );
  MX2XL U6787 ( .A(\I_cache/cache[7][15] ), .B(n9351), .S0(n5366), .Y(n12696)
         );
  MX2XL U6788 ( .A(\I_cache/cache[6][15] ), .B(n9351), .S0(n5418), .Y(n12697)
         );
  MX2XL U6789 ( .A(\I_cache/cache[5][15] ), .B(n9351), .S0(n5284), .Y(n12698)
         );
  MX2XL U6790 ( .A(\I_cache/cache[3][15] ), .B(n9351), .S0(n5198), .Y(n12700)
         );
  MX2XL U6791 ( .A(\I_cache/cache[2][15] ), .B(n9351), .S0(n5240), .Y(n12701)
         );
  MX2XL U6792 ( .A(\I_cache/cache[1][15] ), .B(n9351), .S0(n5102), .Y(n12702)
         );
  MX2XL U6793 ( .A(\I_cache/cache[0][15] ), .B(n9351), .S0(n5153), .Y(n12703)
         );
  MX2XL U6794 ( .A(\I_cache/cache[7][151] ), .B(n3512), .S0(n5366), .Y(n11608)
         );
  MX2XL U6795 ( .A(\I_cache/cache[7][152] ), .B(n10977), .S0(n5366), .Y(n11600) );
  MX2XL U6796 ( .A(\I_cache/cache[7][139] ), .B(n10976), .S0(n5366), .Y(n11704) );
  MX2XL U6797 ( .A(\I_cache/cache[7][140] ), .B(n11157), .S0(n5367), .Y(n11696) );
  MX2XL U6798 ( .A(\I_cache/cache[2][140] ), .B(n11157), .S0(n5233), .Y(n11701) );
  MX2XL U6799 ( .A(\I_cache/cache[0][140] ), .B(n11157), .S0(n5146), .Y(n11703) );
  MX2XL U6800 ( .A(\I_cache/cache[7][136] ), .B(n10980), .S0(n5370), .Y(n11728) );
  MX2XL U6801 ( .A(\I_cache/cache[0][136] ), .B(n10980), .S0(n5149), .Y(n11735) );
  MX2XL U6802 ( .A(\I_cache/cache[6][128] ), .B(n10978), .S0(n5410), .Y(n11793) );
  MX2XL U6803 ( .A(\I_cache/cache[3][128] ), .B(n10978), .S0(n5190), .Y(n11796) );
  MX2XL U6804 ( .A(\I_cache/cache[1][128] ), .B(n10978), .S0(n5103), .Y(n11798) );
  MX2XL U6805 ( .A(\I_cache/cache[7][132] ), .B(n10986), .S0(n5370), .Y(n11760) );
  MX2XL U6806 ( .A(\I_cache/cache[7][148] ), .B(n10983), .S0(n5367), .Y(n11632) );
  MX2XL U6807 ( .A(\I_cache/cache[7][133] ), .B(n10988), .S0(n5370), .Y(n11752) );
  MX2XL U6808 ( .A(\I_cache/cache[6][131] ), .B(n10994), .S0(n5411), .Y(n11769) );
  MX2XL U6809 ( .A(\I_cache/cache[3][131] ), .B(n10994), .S0(n5191), .Y(n11772) );
  MX2XL U6810 ( .A(\I_cache/cache[1][131] ), .B(n10994), .S0(n5104), .Y(n11774) );
  MX2XL U6811 ( .A(\I_cache/cache[7][150] ), .B(n10991), .S0(n5368), .Y(n11616) );
  MX2XL U6812 ( .A(\I_cache/cache[7][145] ), .B(n10990), .S0(n5373), .Y(n11656) );
  MX2XL U6813 ( .A(\I_cache/cache[7][134] ), .B(n10987), .S0(n5374), .Y(n11744) );
  MX2XL U6814 ( .A(\I_cache/cache[6][130] ), .B(n10993), .S0(n5411), .Y(n11777) );
  MX2XL U6815 ( .A(\I_cache/cache[3][130] ), .B(n10993), .S0(n5191), .Y(n11780) );
  MX2XL U6816 ( .A(\I_cache/cache[1][130] ), .B(n10993), .S0(n5104), .Y(n11782) );
  MX2XL U6817 ( .A(\I_cache/cache[6][144] ), .B(n3514), .S0(n5410), .Y(n11665)
         );
  MX2XL U6818 ( .A(\I_cache/cache[3][144] ), .B(n3514), .S0(n5190), .Y(n11668)
         );
  MX2XL U6819 ( .A(\I_cache/cache[1][144] ), .B(n3514), .S0(n5103), .Y(n11670)
         );
  MX2XL U6820 ( .A(\I_cache/cache[7][137] ), .B(n3510), .S0(n5369), .Y(n11720)
         );
  MX2XL U6821 ( .A(\I_cache/cache[7][111] ), .B(n11007), .S0(n5368), .Y(n11928) );
  MX2XL U6822 ( .A(\I_cache/cache[0][111] ), .B(n11007), .S0(n5147), .Y(n11935) );
  MX2XL U6823 ( .A(\I_cache/cache[7][79] ), .B(n11009), .S0(n5368), .Y(n12184)
         );
  MX2XL U6824 ( .A(\I_cache/cache[0][79] ), .B(n11009), .S0(n5147), .Y(n12191)
         );
  MX2XL U6825 ( .A(\I_cache/cache[7][47] ), .B(n11008), .S0(n5368), .Y(n12440)
         );
  MX2XL U6826 ( .A(\I_cache/cache[0][47] ), .B(n11008), .S0(n5147), .Y(n12447)
         );
  MX2XL U6827 ( .A(\I_cache/cache[0][142] ), .B(n11034), .S0(n5147), .Y(n11687) );
  MX2XL U6828 ( .A(\I_cache/cache[7][135] ), .B(n10981), .S0(n5367), .Y(n11736) );
  MX2XL U6829 ( .A(\I_cache/cache[7][143] ), .B(n10996), .S0(n5368), .Y(n11672) );
  MX2XL U6830 ( .A(\I_cache/cache[0][143] ), .B(n10996), .S0(n5147), .Y(n11679) );
  MX2XL U6831 ( .A(\I_cache/cache[0][141] ), .B(n10997), .S0(n5147), .Y(n11695) );
  MX2XL U6832 ( .A(\I_cache/cache[7][149] ), .B(n10985), .S0(n5370), .Y(n11624) );
  MX2XL U6833 ( .A(\I_cache/cache[7][138] ), .B(n10989), .S0(n5366), .Y(n11712) );
  MX2XL U6834 ( .A(\I_cache/cache[7][146] ), .B(n10992), .S0(n5368), .Y(n11648) );
  MX2XL U6835 ( .A(\I_cache/cache[6][139] ), .B(n10976), .S0(n5410), .Y(n11705) );
  MX2XL U6836 ( .A(\I_cache/cache[3][139] ), .B(n10976), .S0(n5190), .Y(n11708) );
  MX2XL U6837 ( .A(\I_cache/cache[1][139] ), .B(n10976), .S0(n5103), .Y(n11710) );
  MX2XL U6838 ( .A(\I_cache/cache[7][129] ), .B(n10995), .S0(n5368), .Y(n11784) );
  MX2XL U6839 ( .A(\I_cache/cache[2][111] ), .B(n11007), .S0(n5234), .Y(n11933) );
  MX2XL U6840 ( .A(\I_cache/cache[2][79] ), .B(n11009), .S0(n5234), .Y(n12189)
         );
  MX2XL U6841 ( .A(\I_cache/cache[2][47] ), .B(n11008), .S0(n5234), .Y(n12445)
         );
  MX2XL U6842 ( .A(\I_cache/cache[2][141] ), .B(n10997), .S0(n5234), .Y(n11693) );
  MX2XL U6843 ( .A(\I_cache/cache[6][132] ), .B(n10986), .S0(n5412), .Y(n11761) );
  MX2XL U6844 ( .A(\I_cache/cache[3][132] ), .B(n10986), .S0(n5198), .Y(n11764) );
  MX2XL U6845 ( .A(\I_cache/cache[6][148] ), .B(n10983), .S0(n5410), .Y(n11633) );
  MX2XL U6846 ( .A(\I_cache/cache[3][148] ), .B(n10983), .S0(n5192), .Y(n11636) );
  MX2XL U6847 ( .A(\I_cache/cache[2][148] ), .B(n10983), .S0(n5238), .Y(n11637) );
  MX2XL U6848 ( .A(\I_cache/cache[6][133] ), .B(n10988), .S0(n5418), .Y(n11753) );
  MX2XL U6849 ( .A(\I_cache/cache[3][133] ), .B(n10988), .S0(n5194), .Y(n11756) );
  MX2XL U6850 ( .A(\I_cache/cache[2][133] ), .B(n10988), .S0(n5240), .Y(n11757) );
  MX2XL U6851 ( .A(\I_cache/cache[6][150] ), .B(n10991), .S0(n5412), .Y(n11617) );
  MX2XL U6852 ( .A(\I_cache/cache[3][150] ), .B(n10991), .S0(n5190), .Y(n11620) );
  MX2XL U6853 ( .A(\I_cache/cache[2][150] ), .B(n10991), .S0(n5242), .Y(n11621) );
  MX2XL U6854 ( .A(\I_cache/cache[6][145] ), .B(n10990), .S0(n5411), .Y(n11657) );
  MX2XL U6855 ( .A(\I_cache/cache[3][145] ), .B(n10990), .S0(n5198), .Y(n11660) );
  MX2XL U6856 ( .A(\I_cache/cache[2][145] ), .B(n10990), .S0(n5241), .Y(n11661) );
  MX2XL U6857 ( .A(\I_cache/cache[6][134] ), .B(n10987), .S0(n5415), .Y(n11745) );
  MX2XL U6858 ( .A(\I_cache/cache[3][134] ), .B(n10987), .S0(n5191), .Y(n11748) );
  MX2XL U6859 ( .A(\I_cache/cache[2][134] ), .B(n10987), .S0(n5239), .Y(n11749) );
  MX2XL U6860 ( .A(\I_cache/cache[2][144] ), .B(n3514), .S0(n5236), .Y(n11669)
         );
  MX2XL U6861 ( .A(\I_cache/cache[6][137] ), .B(n3510), .S0(n5410), .Y(n11721)
         );
  MX2XL U6862 ( .A(\I_cache/cache[3][137] ), .B(n3510), .S0(n5192), .Y(n11724)
         );
  MX2XL U6863 ( .A(\I_cache/cache[2][137] ), .B(n3510), .S0(n5236), .Y(n11725)
         );
  MX2XL U6864 ( .A(\I_cache/cache[6][111] ), .B(n11007), .S0(n5412), .Y(n11929) );
  MX2XL U6865 ( .A(\I_cache/cache[5][111] ), .B(n11007), .S0(n5284), .Y(n11930) );
  MX2XL U6866 ( .A(\I_cache/cache[6][79] ), .B(n11009), .S0(n5412), .Y(n12185)
         );
  MX2XL U6867 ( .A(\I_cache/cache[5][79] ), .B(n11009), .S0(n5277), .Y(n12186)
         );
  MX2XL U6868 ( .A(\I_cache/cache[6][47] ), .B(n11008), .S0(n5412), .Y(n12441)
         );
  MX2XL U6869 ( .A(\I_cache/cache[5][47] ), .B(n11008), .S0(n5284), .Y(n12442)
         );
  MX2XL U6870 ( .A(\I_cache/cache[6][142] ), .B(n11034), .S0(n5412), .Y(n11681) );
  MX2XL U6871 ( .A(\I_cache/cache[2][135] ), .B(n10981), .S0(n5234), .Y(n11741) );
  MX2XL U6872 ( .A(\I_cache/cache[6][138] ), .B(n10989), .S0(n5414), .Y(n11713) );
  MX2XL U6873 ( .A(\I_cache/cache[3][138] ), .B(n10989), .S0(n5196), .Y(n11716) );
  MX2XL U6874 ( .A(\I_cache/cache[2][138] ), .B(n10989), .S0(n5238), .Y(n11717) );
  MX2XL U6875 ( .A(\I_cache/cache[6][146] ), .B(n10992), .S0(n5418), .Y(n11649) );
  MX2XL U6876 ( .A(\I_cache/cache[3][146] ), .B(n10992), .S0(n5194), .Y(n11652) );
  MX2XL U6877 ( .A(\I_cache/cache[2][146] ), .B(n10992), .S0(n5240), .Y(n11653) );
  MX2XL U6878 ( .A(\I_cache/cache[5][129] ), .B(n10995), .S0(n5278), .Y(n11786) );
  MX2XL U6879 ( .A(\I_cache/cache[4][111] ), .B(n11007), .S0(n5321), .Y(n11931) );
  MX2XL U6880 ( .A(\I_cache/cache[4][79] ), .B(n11009), .S0(n5321), .Y(n12187)
         );
  MX2XL U6881 ( .A(\I_cache/cache[4][47] ), .B(n11008), .S0(n5321), .Y(n12443)
         );
  MX2XL U6882 ( .A(\I_cache/cache[1][132] ), .B(n10986), .S0(n5102), .Y(n11766) );
  MX2XL U6883 ( .A(\I_cache/cache[1][148] ), .B(n10983), .S0(n5102), .Y(n11638) );
  MX2XL U6884 ( .A(\I_cache/cache[0][148] ), .B(n10983), .S0(n5149), .Y(n11639) );
  MX2XL U6885 ( .A(\I_cache/cache[1][133] ), .B(n10988), .S0(n5102), .Y(n11758) );
  MX2XL U6886 ( .A(\I_cache/cache[0][133] ), .B(n10988), .S0(n5149), .Y(n11759) );
  MX2XL U6887 ( .A(\I_cache/cache[1][150] ), .B(n10991), .S0(n5102), .Y(n11622) );
  MX2XL U6888 ( .A(\I_cache/cache[0][150] ), .B(n10991), .S0(n5147), .Y(n11623) );
  MX2XL U6889 ( .A(\I_cache/cache[1][134] ), .B(n10987), .S0(n5102), .Y(n11750) );
  MX2XL U6890 ( .A(\I_cache/cache[0][134] ), .B(n10987), .S0(n5149), .Y(n11751) );
  MX2XL U6891 ( .A(\I_cache/cache[0][144] ), .B(n3514), .S0(n5145), .Y(n11671)
         );
  MX2XL U6892 ( .A(\I_cache/cache[1][137] ), .B(n3510), .S0(n5102), .Y(n11726)
         );
  MX2XL U6893 ( .A(\I_cache/cache[0][137] ), .B(n3510), .S0(n5145), .Y(n11727)
         );
  MX2XL U6894 ( .A(\I_cache/cache[3][111] ), .B(n11007), .S0(n5192), .Y(n11932) );
  MX2XL U6895 ( .A(\I_cache/cache[1][111] ), .B(n11007), .S0(n5105), .Y(n11934) );
  MX2XL U6896 ( .A(\I_cache/cache[3][79] ), .B(n11009), .S0(n5192), .Y(n12188)
         );
  MX2XL U6897 ( .A(\I_cache/cache[1][79] ), .B(n11009), .S0(n5105), .Y(n12190)
         );
  MX2XL U6898 ( .A(\I_cache/cache[3][47] ), .B(n11008), .S0(n5192), .Y(n12444)
         );
  MX2XL U6899 ( .A(\I_cache/cache[1][47] ), .B(n11008), .S0(n5105), .Y(n12446)
         );
  MX2XL U6900 ( .A(\I_cache/cache[0][135] ), .B(n10981), .S0(n5153), .Y(n11743) );
  MX2XL U6901 ( .A(\I_cache/cache[1][138] ), .B(n10989), .S0(n5102), .Y(n11718) );
  MX2XL U6902 ( .A(\I_cache/cache[0][138] ), .B(n10989), .S0(n5146), .Y(n11719) );
  MX2XL U6903 ( .A(\I_cache/cache[1][146] ), .B(n10992), .S0(n5102), .Y(n11654) );
  MX2XL U6904 ( .A(\I_cache/cache[0][146] ), .B(n10992), .S0(n5147), .Y(n11655) );
  MX2XL U6905 ( .A(\I_cache/cache[4][145] ), .B(n10990), .S0(n5321), .Y(n11659) );
  MX2XL U6906 ( .A(\I_cache/cache[5][145] ), .B(n10990), .S0(n5284), .Y(n11658) );
  NAND2XL U6907 ( .A(n12961), .B(net113087), .Y(net99060) );
  NAND2XL U6908 ( .A(\i_MIPS/EX_MEM[6] ), .B(net113089), .Y(n10830) );
  NAND2XL U6909 ( .A(\i_MIPS/EX_MEM[5] ), .B(net113087), .Y(net98967) );
  NAND2XL U6910 ( .A(n12953), .B(net113089), .Y(net99311) );
  NAND2XL U6911 ( .A(n12949), .B(net113089), .Y(net99428) );
  OA22XL U6912 ( .A0(n5344), .A1(n1206), .B0(n5300), .B1(n2778), .Y(n9753) );
  OA22XL U6913 ( .A0(n5354), .A1(n1207), .B0(n5310), .B1(n2779), .Y(n10228) );
  OA22XL U6914 ( .A0(n5345), .A1(n1208), .B0(n5301), .B1(n2780), .Y(n9800) );
  OA22XL U6915 ( .A0(n5344), .A1(n1209), .B0(n5300), .B1(n2781), .Y(n9745) );
  OA22XL U6916 ( .A0(n5344), .A1(n1210), .B0(n5300), .B1(n2782), .Y(n9761) );
  OA22XL U6917 ( .A0(n5342), .A1(n1211), .B0(n5298), .B1(n2783), .Y(n9693) );
  OA22XL U6918 ( .A0(n5345), .A1(n1212), .B0(n5301), .B1(n2784), .Y(n9790) );
  OA22XL U6919 ( .A0(n5345), .A1(n1213), .B0(n5301), .B1(n2785), .Y(n9776) );
  OA22XL U6920 ( .A0(n5344), .A1(n1214), .B0(n5300), .B1(n2786), .Y(n9766) );
  OA22XL U6921 ( .A0(n5342), .A1(n1215), .B0(n5298), .B1(n2787), .Y(n9698) );
  OA22XL U6922 ( .A0(n5343), .A1(n1216), .B0(n5299), .B1(n2788), .Y(n9717) );
  OA22XL U6923 ( .A0(n5343), .A1(n1217), .B0(n5299), .B1(n2789), .Y(n9732) );
  OA22XL U6924 ( .A0(n5343), .A1(n1218), .B0(n5299), .B1(n2790), .Y(n9727) );
  OA22XL U6925 ( .A0(n5343), .A1(n1219), .B0(n5299), .B1(n2791), .Y(n9722) );
  OA22XL U6926 ( .A0(n5353), .A1(n1785), .B0(n5309), .B1(n3469), .Y(n10106) );
  OA22XL U6927 ( .A0(n5354), .A1(n1786), .B0(n5310), .B1(n3470), .Y(n10116) );
  OA22XL U6928 ( .A0(n5354), .A1(n1787), .B0(n5310), .B1(n3471), .Y(n10121) );
  OA22XL U6929 ( .A0(n5354), .A1(n1788), .B0(n5310), .B1(n3472), .Y(n10111) );
  OA22XL U6930 ( .A0(n5346), .A1(n1789), .B0(n5302), .B1(n3473), .Y(n9840) );
  OA22XL U6931 ( .A0(n5346), .A1(n1790), .B0(n5302), .B1(n3474), .Y(n9845) );
  OA22XL U6932 ( .A0(n5350), .A1(n1791), .B0(n5306), .B1(n3475), .Y(n9975) );
  OA22XL U6933 ( .A0(n5350), .A1(n1792), .B0(n5306), .B1(n3476), .Y(n9985) );
  OA22XL U6934 ( .A0(n5350), .A1(n1793), .B0(n5306), .B1(n3477), .Y(n9980) );
  OA22XL U6935 ( .A0(n5353), .A1(n1794), .B0(n5309), .B1(n3478), .Y(n10072) );
  OA22XL U6936 ( .A0(n5342), .A1(n1795), .B0(n5298), .B1(n3479), .Y(n9680) );
  OA22XL U6937 ( .A0(n5355), .A1(n1796), .B0(n5311), .B1(n3480), .Y(n11121) );
  OA22XL U6938 ( .A0(n5355), .A1(n1797), .B0(n5311), .B1(n3481), .Y(n11131) );
  OA22XL U6939 ( .A0(n5355), .A1(n1798), .B0(n5311), .B1(n3482), .Y(n11142) );
  OA22XL U6940 ( .A0(n5355), .A1(n1799), .B0(n5311), .B1(n3483), .Y(n11126) );
  AO21XL U6941 ( .A0(n3321), .A1(net111881), .B0(\D_cache/cache[7][154] ), .Y(
        \D_cache/n557 ) );
  AO21XL U6942 ( .A0(n3321), .A1(net112011), .B0(\D_cache/cache[6][154] ), .Y(
        \D_cache/n558 ) );
  AO21XL U6943 ( .A0(n3321), .A1(net112121), .B0(\D_cache/cache[5][154] ), .Y(
        \D_cache/n559 ) );
  AO21XL U6944 ( .A0(n3321), .A1(net112211), .B0(\D_cache/cache[4][154] ), .Y(
        \D_cache/n560 ) );
  AO21XL U6945 ( .A0(n3321), .A1(net112283), .B0(\D_cache/cache[3][154] ), .Y(
        \D_cache/n561 ) );
  AO21XL U6946 ( .A0(n3321), .A1(net112423), .B0(\D_cache/cache[2][154] ), .Y(
        \D_cache/n562 ) );
  AO21XL U6947 ( .A0(n3321), .A1(net112547), .B0(\D_cache/cache[1][154] ), .Y(
        \D_cache/n563 ) );
  AO21XL U6948 ( .A0(n3321), .A1(net112649), .B0(\D_cache/cache[0][154] ), .Y(
        \D_cache/n564 ) );
  AO21XL U6949 ( .A0(n4793), .A1(n5325), .B0(\I_cache/cache[4][154] ), .Y(
        n11587) );
  AO21XL U6950 ( .A0(n4793), .A1(n5371), .B0(\I_cache/cache[7][154] ), .Y(
        n11584) );
  AO21XL U6951 ( .A0(n4793), .A1(n5416), .B0(\I_cache/cache[6][154] ), .Y(
        n11585) );
  AO21XL U6952 ( .A0(n4793), .A1(n5285), .B0(\I_cache/cache[5][154] ), .Y(
        n11586) );
  AO21XL U6953 ( .A0(n4793), .A1(n5195), .B0(\I_cache/cache[3][154] ), .Y(
        n11588) );
  AO21XL U6954 ( .A0(n4793), .A1(n5242), .B0(\I_cache/cache[2][154] ), .Y(
        n11589) );
  AO21XL U6955 ( .A0(n4793), .A1(n5111), .B0(\I_cache/cache[1][154] ), .Y(
        n11590) );
  AO21XL U6956 ( .A0(n4793), .A1(n5148), .B0(\I_cache/cache[0][154] ), .Y(
        n11591) );
  XOR2X4 U6957 ( .A(n11386), .B(ICACHE_addr[27]), .Y(n9549) );
  CLKBUFX3 U6958 ( .A(n154), .Y(n5514) );
  CLKBUFX3 U6959 ( .A(n154), .Y(n5515) );
  CLKBUFX3 U6960 ( .A(n154), .Y(n5513) );
  CLKBUFX3 U6961 ( .A(n154), .Y(n5512) );
  CLKBUFX3 U6962 ( .A(n5518), .Y(n5517) );
  CLKBUFX3 U6963 ( .A(n5518), .Y(n5516) );
  CLKBUFX3 U6964 ( .A(n10835), .Y(n5096) );
  CLKBUFX3 U6965 ( .A(n10835), .Y(n5095) );
  INVX3 U6966 ( .A(n5443), .Y(n5414) );
  INVX3 U6967 ( .A(n5351), .Y(n5323) );
  INVX3 U6968 ( .A(n5247), .Y(n5236) );
  INVX3 U6969 ( .A(n5158), .Y(n5149) );
  INVX3 U6970 ( .A(n5423), .Y(n5413) );
  INVX3 U6971 ( .A(n5328), .Y(n5322) );
  INVX3 U6972 ( .A(n5263), .Y(n5235) );
  INVX3 U6973 ( .A(n5159), .Y(n5148) );
  INVX3 U6974 ( .A(n5425), .Y(n5411) );
  INVX3 U6975 ( .A(n5348), .Y(n5320) );
  INVX3 U6976 ( .A(n5263), .Y(n5233) );
  INVX3 U6977 ( .A(n5160), .Y(n5146) );
  INVX3 U6978 ( .A(n5177), .Y(n5145) );
  INVX3 U6979 ( .A(n5422), .Y(n5416) );
  INVX3 U6980 ( .A(n5348), .Y(n5325) );
  INVX3 U6981 ( .A(n5246), .Y(n5238) );
  INVX3 U6982 ( .A(n5443), .Y(n5419) );
  INVX3 U6983 ( .A(n5243), .Y(n5241) );
  INVX3 U6984 ( .A(n5177), .Y(n5154) );
  INVX3 U6985 ( .A(n5329), .Y(n5321) );
  INVX3 U6986 ( .A(n5266), .Y(n5234) );
  INVX3 U6987 ( .A(n5177), .Y(n5147) );
  INVX3 U6988 ( .A(n5351), .Y(n5326) );
  INVX3 U6989 ( .A(n5245), .Y(n5239) );
  INVX3 U6990 ( .A(n5177), .Y(n5152) );
  INVX3 U6991 ( .A(n5244), .Y(n5240) );
  INVX3 U6992 ( .A(net112081), .Y(net111999) );
  INVX3 U6993 ( .A(net112047), .Y(net111995) );
  INVX3 U6994 ( .A(net112081), .Y(net111989) );
  INVX3 U6995 ( .A(net112443), .Y(net112401) );
  INVX3 U6996 ( .A(net112063), .Y(net112009) );
  INVX3 U6997 ( .A(net112443), .Y(net112405) );
  INVX3 U6998 ( .A(net112033), .Y(net111991) );
  INVX3 U6999 ( .A(net112431), .Y(net112417) );
  INVX3 U7000 ( .A(net112429), .Y(net112419) );
  INVX3 U7001 ( .A(n5132), .Y(n5102) );
  INVX3 U7002 ( .A(n5397), .Y(n5370) );
  INVX3 U7003 ( .A(n5217), .Y(n5194) );
  INVX3 U7004 ( .A(n5116), .Y(n5107) );
  INVX3 U7005 ( .A(n5379), .Y(n5369) );
  INVX3 U7006 ( .A(n5221), .Y(n5193) );
  INVX3 U7007 ( .A(n5132), .Y(n5106) );
  INVX3 U7008 ( .A(n5381), .Y(n5367) );
  INVX3 U7009 ( .A(n5218), .Y(n5191) );
  INVX3 U7010 ( .A(n5118), .Y(n5104) );
  INVX3 U7011 ( .A(n5378), .Y(n5371) );
  INVX3 U7012 ( .A(n5218), .Y(n5195) );
  INVX3 U7013 ( .A(n5221), .Y(n5190) );
  INVX3 U7014 ( .A(n5136), .Y(n5103) );
  INVX3 U7015 ( .A(n5394), .Y(n5372) );
  INVX3 U7016 ( .A(n5115), .Y(n5109) );
  INVX3 U7017 ( .A(n5397), .Y(n5374) );
  INVX3 U7018 ( .A(n5200), .Y(n5199) );
  INVX3 U7019 ( .A(n5136), .Y(n5110) );
  INVX3 U7020 ( .A(n5217), .Y(n5192) );
  INVX3 U7021 ( .A(n5117), .Y(n5105) );
  INVX3 U7022 ( .A(net112343), .Y(net112289) );
  INVX3 U7023 ( .A(net111941), .Y(net111865) );
  INVX3 U7024 ( .A(net112337), .Y(net112277) );
  INVX3 U7025 ( .A(net111929), .Y(net111879) );
  INVX3 U7026 ( .A(net112345), .Y(net112291) );
  INVX3 U7027 ( .A(net111929), .Y(net111885) );
  INVX3 U7028 ( .A(net111929), .Y(net111867) );
  INVX3 U7029 ( .A(n3688), .Y(net112279) );
  INVX3 U7030 ( .A(net111929), .Y(net111881) );
  INVX3 U7031 ( .A(net111941), .Y(net111883) );
  INVX3 U7032 ( .A(net112235), .Y(net112215) );
  CLKBUFX3 U7033 ( .A(net110231), .Y(net110219) );
  CLKBUFX3 U7034 ( .A(n5499), .Y(n5493) );
  CLKBUFX3 U7035 ( .A(n5498), .Y(n5494) );
  CLKBUFX3 U7036 ( .A(n5498), .Y(n5495) );
  CLKBUFX3 U7037 ( .A(n5498), .Y(n5497) );
  CLKBUFX3 U7038 ( .A(n5498), .Y(n5496) );
  CLKBUFX3 U7039 ( .A(n5499), .Y(n5492) );
  CLKBUFX3 U7040 ( .A(n5499), .Y(n5490) );
  CLKBUFX3 U7041 ( .A(n5499), .Y(n5491) );
  CLKBUFX3 U7042 ( .A(n5498), .Y(n5489) );
  CLKBUFX3 U7043 ( .A(net110233), .Y(net110221) );
  CLKBUFX3 U7044 ( .A(n5188), .Y(n5161) );
  CLKBUFX3 U7045 ( .A(n5449), .Y(n5426) );
  CLKBUFX3 U7046 ( .A(n5188), .Y(n5160) );
  CLKBUFX3 U7047 ( .A(net112097), .Y(net112033) );
  CLKBUFX3 U7048 ( .A(net112101), .Y(net112019) );
  CLKBUFX3 U7049 ( .A(n5231), .Y(n5200) );
  CLKBUFX3 U7050 ( .A(n5404), .Y(n5382) );
  CLKBUFX3 U7051 ( .A(n5316), .Y(n5287) );
  CLKBUFX3 U7052 ( .A(net111977), .Y(net111889) );
  CLKBUFX3 U7053 ( .A(net112385), .Y(net112319) );
  CLKBUFX3 U7054 ( .A(net112093), .Y(net112051) );
  CLKBUFX3 U7055 ( .A(n5272), .Y(n5256) );
  CLKBUFX3 U7056 ( .A(n5185), .Y(n5170) );
  CLKBUFX3 U7057 ( .A(net112499), .Y(net112477) );
  CLKBUFX3 U7058 ( .A(net112093), .Y(net112049) );
  CLKBUFX3 U7059 ( .A(net112093), .Y(net112047) );
  CLKBUFX3 U7060 ( .A(net112093), .Y(net112045) );
  CLKBUFX3 U7061 ( .A(n5360), .Y(n5336) );
  CLKBUFX3 U7062 ( .A(n5360), .Y(n5338) );
  CLKBUFX3 U7063 ( .A(n5359), .Y(n5340) );
  CLKBUFX3 U7064 ( .A(n5359), .Y(n5342) );
  CLKBUFX3 U7065 ( .A(net112503), .Y(net112469) );
  CLKBUFX3 U7066 ( .A(n5273), .Y(n5252) );
  CLKBUFX3 U7067 ( .A(n5186), .Y(n5166) );
  CLKBUFX3 U7068 ( .A(n5273), .Y(n5254) );
  CLKBUFX3 U7069 ( .A(n5186), .Y(n5168) );
  CLKBUFX3 U7070 ( .A(n5360), .Y(n5337) );
  CLKBUFX3 U7071 ( .A(n5273), .Y(n5253) );
  CLKBUFX3 U7072 ( .A(n5186), .Y(n5167) );
  CLKBUFX3 U7073 ( .A(n5358), .Y(n5346) );
  CLKBUFX3 U7074 ( .A(n5271), .Y(n5262) );
  CLKBUFX3 U7075 ( .A(n5184), .Y(n5176) );
  CLKBUFX3 U7076 ( .A(n5359), .Y(n5341) );
  CLKBUFX3 U7077 ( .A(n5272), .Y(n5257) );
  CLKBUFX3 U7078 ( .A(n5185), .Y(n5171) );
  CLKBUFX3 U7079 ( .A(n5357), .Y(n5350) );
  CLKBUFX3 U7080 ( .A(n5270), .Y(n5265) );
  CLKBUFX3 U7081 ( .A(n5158), .Y(n5179) );
  CLKBUFX3 U7082 ( .A(n5428), .Y(n5442) );
  CLKBUFX3 U7083 ( .A(n5361), .Y(n5335) );
  CLKBUFX3 U7084 ( .A(n5274), .Y(n5251) );
  CLKBUFX3 U7085 ( .A(n5187), .Y(n5165) );
  CLKBUFX3 U7086 ( .A(n5272), .Y(n5258) );
  CLKBUFX3 U7087 ( .A(n5185), .Y(n5172) );
  CLKBUFX3 U7088 ( .A(n3611), .Y(n5441) );
  CLKBUFX3 U7089 ( .A(n5272), .Y(n5264) );
  CLKBUFX3 U7090 ( .A(n5273), .Y(n5255) );
  CLKBUFX3 U7091 ( .A(n5159), .Y(n5178) );
  CLKBUFX3 U7092 ( .A(n5186), .Y(n5169) );
  CLKBUFX3 U7093 ( .A(n5360), .Y(n5339) );
  CLKBUFX3 U7094 ( .A(n5357), .Y(n5349) );
  CLKBUFX3 U7095 ( .A(net112087), .Y(net112069) );
  CLKBUFX3 U7096 ( .A(net112497), .Y(net112489) );
  CLKBUFX3 U7097 ( .A(net112087), .Y(net112073) );
  CLKBUFX3 U7098 ( .A(net112089), .Y(net112067) );
  CLKBUFX3 U7099 ( .A(net112091), .Y(net112053) );
  CLKBUFX3 U7100 ( .A(net112087), .Y(net112075) );
  CLKBUFX3 U7101 ( .A(net112085), .Y(net112079) );
  CLKBUFX3 U7102 ( .A(net112089), .Y(net112065) );
  CLKBUFX3 U7103 ( .A(net112091), .Y(net112057) );
  CLKBUFX3 U7104 ( .A(net112091), .Y(net112055) );
  CLKBUFX3 U7105 ( .A(n5356), .Y(n5354) );
  CLKBUFX3 U7106 ( .A(n5358), .Y(n5345) );
  CLKBUFX3 U7107 ( .A(n5441), .Y(n5438) );
  CLKBUFX3 U7108 ( .A(n5271), .Y(n5261) );
  CLKBUFX3 U7109 ( .A(n5184), .Y(n5175) );
  CLKBUFX3 U7110 ( .A(n5358), .Y(n5344) );
  CLKBUFX3 U7111 ( .A(n5441), .Y(n5437) );
  CLKBUFX3 U7112 ( .A(n5271), .Y(n5260) );
  CLKBUFX3 U7113 ( .A(n5184), .Y(n5174) );
  CLKBUFX3 U7114 ( .A(n5359), .Y(n5343) );
  CLKBUFX3 U7115 ( .A(n5272), .Y(n5259) );
  CLKBUFX3 U7116 ( .A(n5185), .Y(n5173) );
  CLKBUFX3 U7117 ( .A(n5447), .Y(n5445) );
  CLKBUFX3 U7118 ( .A(n5270), .Y(n5268) );
  CLKBUFX3 U7119 ( .A(n5165), .Y(n5183) );
  CLKBUFX3 U7120 ( .A(n5357), .Y(n5348) );
  CLKBUFX3 U7121 ( .A(n5439), .Y(n5440) );
  CLKBUFX3 U7122 ( .A(n5358), .Y(n5347) );
  CLKBUFX3 U7123 ( .A(n5271), .Y(n5263) );
  CLKBUFX3 U7124 ( .A(n5184), .Y(n5177) );
  CLKBUFX3 U7125 ( .A(n5357), .Y(n5351) );
  CLKBUFX3 U7126 ( .A(n5269), .Y(n5266) );
  CLKBUFX3 U7127 ( .A(n5181), .Y(n5180) );
  CLKBUFX3 U7128 ( .A(n5356), .Y(n5352) );
  CLKBUFX3 U7129 ( .A(n5447), .Y(n5443) );
  CLKBUFX3 U7130 ( .A(n5173), .Y(n5181) );
  CLKBUFX3 U7131 ( .A(n5356), .Y(n5353) );
  CLKBUFX3 U7132 ( .A(n5447), .Y(n5444) );
  CLKBUFX3 U7133 ( .A(n5270), .Y(n5267) );
  CLKBUFX3 U7134 ( .A(n5165), .Y(n5182) );
  CLKBUFX3 U7135 ( .A(n5227), .Y(n5210) );
  CLKBUFX3 U7136 ( .A(n5315), .Y(n5292) );
  CLKBUFX3 U7137 ( .A(n5315), .Y(n5294) );
  CLKBUFX3 U7138 ( .A(n5315), .Y(n5296) );
  CLKBUFX3 U7139 ( .A(n5313), .Y(n5298) );
  CLKBUFX3 U7140 ( .A(n5228), .Y(n5206) );
  CLKBUFX3 U7141 ( .A(n5228), .Y(n5208) );
  CLKBUFX3 U7142 ( .A(n5315), .Y(n5293) );
  CLKBUFX3 U7143 ( .A(n5228), .Y(n5207) );
  CLKBUFX3 U7144 ( .A(n5142), .Y(n5123) );
  CLKBUFX3 U7145 ( .A(n5140), .Y(n5131) );
  CLKBUFX3 U7146 ( .A(n5315), .Y(n5297) );
  CLKBUFX3 U7147 ( .A(n5227), .Y(n5211) );
  CLKBUFX3 U7148 ( .A(n5313), .Y(n5306) );
  CLKBUFX3 U7149 ( .A(n5225), .Y(n5220) );
  CLKBUFX3 U7150 ( .A(n5140), .Y(n5135) );
  CLKBUFX3 U7151 ( .A(n5409), .Y(n5396) );
  CLKBUFX3 U7152 ( .A(n5227), .Y(n5212) );
  CLKBUFX3 U7153 ( .A(n5315), .Y(n5295) );
  CLKBUFX3 U7154 ( .A(n5228), .Y(n5209) );
  CLKBUFX3 U7155 ( .A(n5225), .Y(n5219) );
  CLKBUFX3 U7156 ( .A(n5142), .Y(n5134) );
  CLKBUFX3 U7157 ( .A(net111961), .Y(net111951) );
  CLKBUFX3 U7158 ( .A(net111969), .Y(net111927) );
  CLKBUFX3 U7159 ( .A(net111967), .Y(net111933) );
  CLKBUFX3 U7160 ( .A(net111965), .Y(net111943) );
  CLKBUFX3 U7161 ( .A(net112319), .Y(net112369) );
  CLKBUFX3 U7162 ( .A(net111969), .Y(net111921) );
  CLKBUFX3 U7163 ( .A(net112301), .Y(net112367) );
  CLKBUFX3 U7164 ( .A(net111963), .Y(net111919) );
  CLKBUFX3 U7165 ( .A(net111969), .Y(net111925) );
  CLKBUFX3 U7166 ( .A(net111969), .Y(net111923) );
  CLKBUFX3 U7167 ( .A(n5312), .Y(n5310) );
  CLKBUFX3 U7168 ( .A(n5314), .Y(n5301) );
  CLKBUFX3 U7169 ( .A(n5226), .Y(n5215) );
  CLKBUFX3 U7170 ( .A(n5140), .Y(n5130) );
  CLKBUFX3 U7171 ( .A(n5314), .Y(n5300) );
  CLKBUFX3 U7172 ( .A(n5401), .Y(n5392) );
  CLKBUFX3 U7173 ( .A(n5226), .Y(n5214) );
  CLKBUFX3 U7174 ( .A(n5140), .Y(n5129) );
  CLKBUFX3 U7175 ( .A(n5287), .Y(n5299) );
  CLKBUFX3 U7176 ( .A(n5227), .Y(n5213) );
  CLKBUFX3 U7177 ( .A(n5224), .Y(n5223) );
  CLKBUFX3 U7178 ( .A(n5313), .Y(n5304) );
  CLKBUFX3 U7179 ( .A(n5393), .Y(n5394) );
  CLKBUFX3 U7180 ( .A(n5225), .Y(n5218) );
  CLKBUFX3 U7181 ( .A(n5132), .Y(n5133) );
  CLKBUFX3 U7182 ( .A(n5314), .Y(n5303) );
  CLKBUFX3 U7183 ( .A(n5401), .Y(n5393) );
  CLKBUFX3 U7184 ( .A(n5226), .Y(n5217) );
  CLKBUFX3 U7185 ( .A(n5140), .Y(n5132) );
  CLKBUFX3 U7186 ( .A(n5313), .Y(n5307) );
  CLKBUFX3 U7187 ( .A(n5393), .Y(n5397) );
  CLKBUFX3 U7188 ( .A(n5312), .Y(n5308) );
  CLKBUFX3 U7189 ( .A(n5224), .Y(n5221) );
  CLKBUFX3 U7190 ( .A(n5139), .Y(n5136) );
  CLKBUFX3 U7191 ( .A(n5312), .Y(n5309) );
  CLKBUFX3 U7192 ( .A(n5224), .Y(n5222) );
  CLKBUFX3 U7193 ( .A(n5139), .Y(n5137) );
  CLKBUFX3 U7194 ( .A(n5356), .Y(n5355) );
  CLKBUFX3 U7195 ( .A(n5447), .Y(n5446) );
  CLKBUFX3 U7196 ( .A(n5270), .Y(n5269) );
  CLKBUFX3 U7197 ( .A(n3750), .Y(net111959) );
  CLKBUFX3 U7198 ( .A(n5312), .Y(n5311) );
  CLKBUFX3 U7199 ( .A(n5139), .Y(n5138) );
  CLKBUFX3 U7200 ( .A(n9116), .Y(n4895) );
  INVX3 U7201 ( .A(n4566), .Y(n4963) );
  INVX3 U7202 ( .A(n4566), .Y(n4962) );
  INVX3 U7203 ( .A(n4566), .Y(n4961) );
  CLKINVX1 U7204 ( .A(n5076), .Y(n5075) );
  CLKBUFX3 U7205 ( .A(n5915), .Y(n5913) );
  CLKBUFX3 U7206 ( .A(n5915), .Y(n5912) );
  CLKBUFX3 U7207 ( .A(n5915), .Y(n5911) );
  CLKBUFX3 U7208 ( .A(n5915), .Y(n5910) );
  CLKBUFX3 U7209 ( .A(n5915), .Y(n5909) );
  CLKBUFX3 U7210 ( .A(n5915), .Y(n5908) );
  CLKBUFX3 U7211 ( .A(n5915), .Y(n5907) );
  CLKBUFX3 U7212 ( .A(n5915), .Y(n5906) );
  CLKBUFX3 U7213 ( .A(n5915), .Y(n5905) );
  CLKBUFX3 U7214 ( .A(n5915), .Y(n5904) );
  CLKBUFX3 U7215 ( .A(n5915), .Y(n5903) );
  CLKBUFX3 U7216 ( .A(n5916), .Y(n5902) );
  CLKBUFX3 U7217 ( .A(n5916), .Y(n5901) );
  CLKBUFX3 U7218 ( .A(n5916), .Y(n5900) );
  CLKBUFX3 U7219 ( .A(n5916), .Y(n5899) );
  CLKBUFX3 U7220 ( .A(n5916), .Y(n5898) );
  CLKBUFX3 U7221 ( .A(n5916), .Y(n5897) );
  CLKBUFX3 U7222 ( .A(n5916), .Y(n5896) );
  CLKBUFX3 U7223 ( .A(n5916), .Y(n5895) );
  CLKBUFX3 U7224 ( .A(n5916), .Y(n5894) );
  CLKBUFX3 U7225 ( .A(n5916), .Y(n5893) );
  CLKBUFX3 U7226 ( .A(n5916), .Y(n5892) );
  CLKBUFX3 U7227 ( .A(n5916), .Y(n5891) );
  CLKBUFX3 U7228 ( .A(n5917), .Y(n5890) );
  CLKBUFX3 U7229 ( .A(n5917), .Y(n5889) );
  CLKBUFX3 U7230 ( .A(n5917), .Y(n5888) );
  CLKBUFX3 U7231 ( .A(n5917), .Y(n5887) );
  CLKBUFX3 U7232 ( .A(n5917), .Y(n5886) );
  CLKBUFX3 U7233 ( .A(n5917), .Y(n5885) );
  CLKBUFX3 U7234 ( .A(n5917), .Y(n5884) );
  CLKBUFX3 U7235 ( .A(n5917), .Y(n5883) );
  CLKBUFX3 U7236 ( .A(n5917), .Y(n5882) );
  CLKBUFX3 U7237 ( .A(n5917), .Y(n5881) );
  CLKBUFX3 U7238 ( .A(n5917), .Y(n5880) );
  CLKBUFX3 U7239 ( .A(n5917), .Y(n5879) );
  CLKBUFX3 U7240 ( .A(n5918), .Y(n5878) );
  CLKBUFX3 U7241 ( .A(n5918), .Y(n5877) );
  CLKBUFX3 U7242 ( .A(n5918), .Y(n5876) );
  CLKBUFX3 U7243 ( .A(n5918), .Y(n5875) );
  CLKBUFX3 U7244 ( .A(n5918), .Y(n5874) );
  CLKBUFX3 U7245 ( .A(n5918), .Y(n5873) );
  CLKBUFX3 U7246 ( .A(n5918), .Y(n5872) );
  CLKBUFX3 U7247 ( .A(n5918), .Y(n5871) );
  CLKBUFX3 U7248 ( .A(n5918), .Y(n5870) );
  CLKBUFX3 U7249 ( .A(n5918), .Y(n5869) );
  CLKBUFX3 U7250 ( .A(n5918), .Y(n5868) );
  CLKBUFX3 U7251 ( .A(n5918), .Y(n5867) );
  CLKBUFX3 U7252 ( .A(n5919), .Y(n5866) );
  CLKBUFX3 U7253 ( .A(n5919), .Y(n5865) );
  CLKBUFX3 U7254 ( .A(n5919), .Y(n5864) );
  CLKBUFX3 U7255 ( .A(n5919), .Y(n5863) );
  CLKBUFX3 U7256 ( .A(n5919), .Y(n5862) );
  CLKBUFX3 U7257 ( .A(n5919), .Y(n5861) );
  CLKBUFX3 U7258 ( .A(n5919), .Y(n5860) );
  CLKBUFX3 U7259 ( .A(n5919), .Y(n5859) );
  CLKBUFX3 U7260 ( .A(n5919), .Y(n5858) );
  CLKBUFX3 U7261 ( .A(n5919), .Y(n5857) );
  CLKBUFX3 U7262 ( .A(n5919), .Y(n5856) );
  CLKBUFX3 U7263 ( .A(n5919), .Y(n5855) );
  CLKBUFX3 U7264 ( .A(n5920), .Y(n5854) );
  CLKBUFX3 U7265 ( .A(n5920), .Y(n5853) );
  CLKBUFX3 U7266 ( .A(n5920), .Y(n5852) );
  CLKBUFX3 U7267 ( .A(n5920), .Y(n5851) );
  CLKBUFX3 U7268 ( .A(n5920), .Y(n5850) );
  CLKBUFX3 U7269 ( .A(n5920), .Y(n5849) );
  CLKBUFX3 U7270 ( .A(n5920), .Y(n5848) );
  CLKBUFX3 U7271 ( .A(n5920), .Y(n5847) );
  CLKBUFX3 U7272 ( .A(n5920), .Y(n5846) );
  CLKBUFX3 U7273 ( .A(n5920), .Y(n5845) );
  CLKBUFX3 U7274 ( .A(n5920), .Y(n5844) );
  CLKBUFX3 U7275 ( .A(n5920), .Y(n5843) );
  CLKBUFX3 U7276 ( .A(n5921), .Y(n5842) );
  CLKBUFX3 U7277 ( .A(n5921), .Y(n5841) );
  CLKBUFX3 U7278 ( .A(n5921), .Y(n5840) );
  CLKBUFX3 U7279 ( .A(n5921), .Y(n5839) );
  CLKBUFX3 U7280 ( .A(n5921), .Y(n5838) );
  CLKBUFX3 U7281 ( .A(n5921), .Y(n5837) );
  CLKBUFX3 U7282 ( .A(n5921), .Y(n5836) );
  CLKBUFX3 U7283 ( .A(n5921), .Y(n5835) );
  CLKBUFX3 U7284 ( .A(n5921), .Y(n5834) );
  CLKBUFX3 U7285 ( .A(n5921), .Y(n5833) );
  CLKBUFX3 U7286 ( .A(n5921), .Y(n5832) );
  CLKBUFX3 U7287 ( .A(n5921), .Y(n5831) );
  CLKBUFX3 U7288 ( .A(n5922), .Y(n5830) );
  CLKBUFX3 U7289 ( .A(n5922), .Y(n5829) );
  CLKBUFX3 U7290 ( .A(n5922), .Y(n5828) );
  CLKBUFX3 U7291 ( .A(n5922), .Y(n5827) );
  CLKBUFX3 U7292 ( .A(n5922), .Y(n5826) );
  CLKBUFX3 U7293 ( .A(n5922), .Y(n5825) );
  CLKBUFX3 U7294 ( .A(n5922), .Y(n5824) );
  CLKBUFX3 U7295 ( .A(n5922), .Y(n5823) );
  CLKBUFX3 U7296 ( .A(n5922), .Y(n5822) );
  CLKBUFX3 U7297 ( .A(n5922), .Y(n5821) );
  CLKBUFX3 U7298 ( .A(n5922), .Y(n5820) );
  CLKBUFX3 U7299 ( .A(n5922), .Y(n5819) );
  CLKBUFX3 U7300 ( .A(n5923), .Y(n5818) );
  CLKBUFX3 U7301 ( .A(n5923), .Y(n5817) );
  CLKBUFX3 U7302 ( .A(n5923), .Y(n5816) );
  CLKBUFX3 U7303 ( .A(n5923), .Y(n5815) );
  CLKBUFX3 U7304 ( .A(n5923), .Y(n5814) );
  CLKBUFX3 U7305 ( .A(n5923), .Y(n5813) );
  CLKBUFX3 U7306 ( .A(n5923), .Y(n5812) );
  CLKBUFX3 U7307 ( .A(n5931), .Y(n5707) );
  CLKBUFX3 U7308 ( .A(n5931), .Y(n5706) );
  CLKBUFX3 U7309 ( .A(n5931), .Y(n5705) );
  CLKBUFX3 U7310 ( .A(n5931), .Y(n5704) );
  CLKBUFX3 U7311 ( .A(n5931), .Y(n5703) );
  CLKBUFX3 U7312 ( .A(n5931), .Y(n5702) );
  CLKBUFX3 U7313 ( .A(n5931), .Y(n5701) );
  CLKBUFX3 U7314 ( .A(n5931), .Y(n5700) );
  CLKBUFX3 U7315 ( .A(n5931), .Y(n5699) );
  CLKBUFX3 U7316 ( .A(n5932), .Y(n5698) );
  CLKBUFX3 U7317 ( .A(n5932), .Y(n5697) );
  CLKBUFX3 U7318 ( .A(n5932), .Y(n5696) );
  CLKBUFX3 U7319 ( .A(n5932), .Y(n5695) );
  CLKBUFX3 U7320 ( .A(n5932), .Y(n5694) );
  CLKBUFX3 U7321 ( .A(n5932), .Y(n5693) );
  CLKBUFX3 U7322 ( .A(n5932), .Y(n5692) );
  CLKBUFX3 U7323 ( .A(n5932), .Y(n5691) );
  CLKBUFX3 U7324 ( .A(n5932), .Y(n5690) );
  CLKBUFX3 U7325 ( .A(n5932), .Y(n5689) );
  CLKBUFX3 U7326 ( .A(n5932), .Y(n5688) );
  CLKBUFX3 U7327 ( .A(n5932), .Y(n5687) );
  CLKBUFX3 U7328 ( .A(n5933), .Y(n5686) );
  CLKBUFX3 U7329 ( .A(n5933), .Y(n5685) );
  CLKBUFX3 U7330 ( .A(n5933), .Y(n5684) );
  CLKBUFX3 U7331 ( .A(n5933), .Y(n5683) );
  CLKBUFX3 U7332 ( .A(n5933), .Y(n5682) );
  CLKBUFX3 U7333 ( .A(n5933), .Y(n5681) );
  CLKBUFX3 U7334 ( .A(n5933), .Y(n5680) );
  CLKBUFX3 U7335 ( .A(n5933), .Y(n5679) );
  CLKBUFX3 U7336 ( .A(n5933), .Y(n5678) );
  CLKBUFX3 U7337 ( .A(n5933), .Y(n5677) );
  CLKBUFX3 U7338 ( .A(n5933), .Y(n5676) );
  CLKBUFX3 U7339 ( .A(n5933), .Y(n5675) );
  CLKBUFX3 U7340 ( .A(n5934), .Y(n5674) );
  CLKBUFX3 U7341 ( .A(n5934), .Y(n5673) );
  CLKBUFX3 U7342 ( .A(n5934), .Y(n5672) );
  CLKBUFX3 U7343 ( .A(n5934), .Y(n5671) );
  CLKBUFX3 U7344 ( .A(n5934), .Y(n5670) );
  CLKBUFX3 U7345 ( .A(n5934), .Y(n5669) );
  CLKBUFX3 U7346 ( .A(n5934), .Y(n5668) );
  CLKBUFX3 U7347 ( .A(n5934), .Y(n5667) );
  CLKBUFX3 U7348 ( .A(n5934), .Y(n5666) );
  CLKBUFX3 U7349 ( .A(n5934), .Y(n5665) );
  CLKBUFX3 U7350 ( .A(n5934), .Y(n5664) );
  CLKBUFX3 U7351 ( .A(n5934), .Y(n5663) );
  CLKBUFX3 U7352 ( .A(n5935), .Y(n5662) );
  CLKBUFX3 U7353 ( .A(n5935), .Y(n5661) );
  CLKBUFX3 U7354 ( .A(n5935), .Y(n5660) );
  CLKBUFX3 U7355 ( .A(n5935), .Y(n5659) );
  CLKBUFX3 U7356 ( .A(n5935), .Y(n5658) );
  CLKBUFX3 U7357 ( .A(n5935), .Y(n5657) );
  CLKBUFX3 U7358 ( .A(n5935), .Y(n5656) );
  CLKBUFX3 U7359 ( .A(n5935), .Y(n5655) );
  CLKBUFX3 U7360 ( .A(n5935), .Y(n5654) );
  CLKBUFX3 U7361 ( .A(n5935), .Y(n5653) );
  CLKBUFX3 U7362 ( .A(n5935), .Y(n5652) );
  CLKBUFX3 U7363 ( .A(n5935), .Y(n5651) );
  CLKBUFX3 U7364 ( .A(n5939), .Y(n5650) );
  CLKBUFX3 U7365 ( .A(n5939), .Y(n5649) );
  CLKBUFX3 U7366 ( .A(n5915), .Y(n5648) );
  CLKBUFX3 U7367 ( .A(n5937), .Y(n5647) );
  CLKBUFX3 U7368 ( .A(n5914), .Y(n5646) );
  CLKBUFX3 U7369 ( .A(n5939), .Y(n5645) );
  CLKBUFX3 U7370 ( .A(n5930), .Y(n5644) );
  CLKBUFX3 U7371 ( .A(n5926), .Y(n5643) );
  CLKBUFX3 U7372 ( .A(n5922), .Y(n5642) );
  CLKBUFX3 U7373 ( .A(n5919), .Y(n5641) );
  CLKBUFX3 U7374 ( .A(n5924), .Y(n5640) );
  CLKBUFX3 U7375 ( .A(n5931), .Y(n5639) );
  CLKBUFX3 U7376 ( .A(n5936), .Y(n5638) );
  CLKBUFX3 U7377 ( .A(n5936), .Y(n5637) );
  CLKBUFX3 U7378 ( .A(n5936), .Y(n5636) );
  CLKBUFX3 U7379 ( .A(n5936), .Y(n5635) );
  CLKBUFX3 U7380 ( .A(n5936), .Y(n5634) );
  CLKBUFX3 U7381 ( .A(n5936), .Y(n5633) );
  CLKBUFX3 U7382 ( .A(n5936), .Y(n5632) );
  CLKBUFX3 U7383 ( .A(n5936), .Y(n5631) );
  CLKBUFX3 U7384 ( .A(n5936), .Y(n5630) );
  CLKBUFX3 U7385 ( .A(n5936), .Y(n5629) );
  CLKBUFX3 U7386 ( .A(n5936), .Y(n5628) );
  CLKBUFX3 U7387 ( .A(n5936), .Y(n5627) );
  CLKBUFX3 U7388 ( .A(n5923), .Y(n5811) );
  CLKBUFX3 U7389 ( .A(n5923), .Y(n5810) );
  CLKBUFX3 U7390 ( .A(n5923), .Y(n5809) );
  CLKBUFX3 U7391 ( .A(n5923), .Y(n5808) );
  CLKBUFX3 U7392 ( .A(n5923), .Y(n5807) );
  CLKBUFX3 U7393 ( .A(n5924), .Y(n5806) );
  CLKBUFX3 U7394 ( .A(n5924), .Y(n5805) );
  CLKBUFX3 U7395 ( .A(n5924), .Y(n5804) );
  CLKBUFX3 U7396 ( .A(n5924), .Y(n5803) );
  CLKBUFX3 U7397 ( .A(n5924), .Y(n5802) );
  CLKBUFX3 U7398 ( .A(n5924), .Y(n5801) );
  CLKBUFX3 U7399 ( .A(n5924), .Y(n5800) );
  CLKBUFX3 U7400 ( .A(n5924), .Y(n5799) );
  CLKBUFX3 U7401 ( .A(n5924), .Y(n5798) );
  CLKBUFX3 U7402 ( .A(n5924), .Y(n5797) );
  CLKBUFX3 U7403 ( .A(n5924), .Y(n5796) );
  CLKBUFX3 U7404 ( .A(n5924), .Y(n5795) );
  CLKBUFX3 U7405 ( .A(n5925), .Y(n5794) );
  CLKBUFX3 U7406 ( .A(n5925), .Y(n5793) );
  CLKBUFX3 U7407 ( .A(n5925), .Y(n5792) );
  CLKBUFX3 U7408 ( .A(n5925), .Y(n5791) );
  CLKBUFX3 U7409 ( .A(n5925), .Y(n5790) );
  CLKBUFX3 U7410 ( .A(n5925), .Y(n5789) );
  CLKBUFX3 U7411 ( .A(n5925), .Y(n5788) );
  CLKBUFX3 U7412 ( .A(n5925), .Y(n5787) );
  CLKBUFX3 U7413 ( .A(n5925), .Y(n5786) );
  CLKBUFX3 U7414 ( .A(n5925), .Y(n5785) );
  CLKBUFX3 U7415 ( .A(n5925), .Y(n5784) );
  CLKBUFX3 U7416 ( .A(n5925), .Y(n5783) );
  CLKBUFX3 U7417 ( .A(n5926), .Y(n5782) );
  CLKBUFX3 U7418 ( .A(n5926), .Y(n5781) );
  CLKBUFX3 U7419 ( .A(n5926), .Y(n5780) );
  CLKBUFX3 U7420 ( .A(n5926), .Y(n5779) );
  CLKBUFX3 U7421 ( .A(n5926), .Y(n5778) );
  CLKBUFX3 U7422 ( .A(n5926), .Y(n5777) );
  CLKBUFX3 U7423 ( .A(n5926), .Y(n5776) );
  CLKBUFX3 U7424 ( .A(n5926), .Y(n5775) );
  CLKBUFX3 U7425 ( .A(n5926), .Y(n5774) );
  CLKBUFX3 U7426 ( .A(n5926), .Y(n5773) );
  CLKBUFX3 U7427 ( .A(n5926), .Y(n5772) );
  CLKBUFX3 U7428 ( .A(n5926), .Y(n5771) );
  CLKBUFX3 U7429 ( .A(n5927), .Y(n5770) );
  CLKBUFX3 U7430 ( .A(n5927), .Y(n5769) );
  CLKBUFX3 U7431 ( .A(n5927), .Y(n5768) );
  CLKBUFX3 U7432 ( .A(n5927), .Y(n5767) );
  CLKBUFX3 U7433 ( .A(n5927), .Y(n5766) );
  CLKBUFX3 U7434 ( .A(n5927), .Y(n5765) );
  CLKBUFX3 U7435 ( .A(n5927), .Y(n5764) );
  CLKBUFX3 U7436 ( .A(n5927), .Y(n5763) );
  CLKBUFX3 U7437 ( .A(n5927), .Y(n5762) );
  CLKBUFX3 U7438 ( .A(n5927), .Y(n5761) );
  CLKBUFX3 U7439 ( .A(n5927), .Y(n5760) );
  CLKBUFX3 U7440 ( .A(n5927), .Y(n5759) );
  CLKBUFX3 U7441 ( .A(n5928), .Y(n5758) );
  CLKBUFX3 U7442 ( .A(n5928), .Y(n5757) );
  CLKBUFX3 U7443 ( .A(n5928), .Y(n5756) );
  CLKBUFX3 U7444 ( .A(n5928), .Y(n5755) );
  CLKBUFX3 U7445 ( .A(n5928), .Y(n5754) );
  CLKBUFX3 U7446 ( .A(n5928), .Y(n5753) );
  CLKBUFX3 U7447 ( .A(n5928), .Y(n5752) );
  CLKBUFX3 U7448 ( .A(n5928), .Y(n5751) );
  CLKBUFX3 U7449 ( .A(n5928), .Y(n5750) );
  CLKBUFX3 U7450 ( .A(n5928), .Y(n5749) );
  CLKBUFX3 U7451 ( .A(n5928), .Y(n5748) );
  CLKBUFX3 U7452 ( .A(n5928), .Y(n5747) );
  CLKBUFX3 U7453 ( .A(n5929), .Y(n5746) );
  CLKBUFX3 U7454 ( .A(n5929), .Y(n5745) );
  CLKBUFX3 U7455 ( .A(n5929), .Y(n5744) );
  CLKBUFX3 U7456 ( .A(n5929), .Y(n5743) );
  CLKBUFX3 U7457 ( .A(n5929), .Y(n5742) );
  CLKBUFX3 U7458 ( .A(n5929), .Y(n5741) );
  CLKBUFX3 U7459 ( .A(n5929), .Y(n5740) );
  CLKBUFX3 U7460 ( .A(n5929), .Y(n5739) );
  CLKBUFX3 U7461 ( .A(n5929), .Y(n5738) );
  CLKBUFX3 U7462 ( .A(n5929), .Y(n5737) );
  CLKBUFX3 U7463 ( .A(n5929), .Y(n5736) );
  CLKBUFX3 U7464 ( .A(n5929), .Y(n5735) );
  CLKBUFX3 U7465 ( .A(n5930), .Y(n5734) );
  CLKBUFX3 U7466 ( .A(n5930), .Y(n5733) );
  CLKBUFX3 U7467 ( .A(n5930), .Y(n5732) );
  CLKBUFX3 U7468 ( .A(n5930), .Y(n5731) );
  CLKBUFX3 U7469 ( .A(n5930), .Y(n5730) );
  CLKBUFX3 U7470 ( .A(n5930), .Y(n5729) );
  CLKBUFX3 U7471 ( .A(n5930), .Y(n5728) );
  CLKBUFX3 U7472 ( .A(n5930), .Y(n5727) );
  CLKBUFX3 U7473 ( .A(n5930), .Y(n5726) );
  CLKBUFX3 U7474 ( .A(n5930), .Y(n5725) );
  CLKBUFX3 U7475 ( .A(n5930), .Y(n5724) );
  CLKBUFX3 U7476 ( .A(n5930), .Y(n5723) );
  CLKBUFX3 U7477 ( .A(rst_n), .Y(n5722) );
  CLKBUFX3 U7478 ( .A(n5926), .Y(n5721) );
  CLKBUFX3 U7479 ( .A(n5919), .Y(n5720) );
  CLKBUFX3 U7480 ( .A(n5931), .Y(n5719) );
  CLKBUFX3 U7481 ( .A(n5940), .Y(n5718) );
  CLKBUFX3 U7482 ( .A(n5916), .Y(n5717) );
  CLKBUFX3 U7483 ( .A(n5920), .Y(n5716) );
  CLKBUFX3 U7484 ( .A(n5927), .Y(n5715) );
  CLKBUFX3 U7485 ( .A(n5929), .Y(n5714) );
  CLKBUFX3 U7486 ( .A(n5921), .Y(n5713) );
  CLKBUFX3 U7487 ( .A(n5936), .Y(n5712) );
  CLKBUFX3 U7488 ( .A(n5932), .Y(n5711) );
  CLKBUFX3 U7489 ( .A(n5931), .Y(n5710) );
  CLKBUFX3 U7490 ( .A(n5931), .Y(n5709) );
  CLKBUFX3 U7491 ( .A(n5931), .Y(n5708) );
  CLKBUFX3 U7492 ( .A(n5915), .Y(n5914) );
  CLKINVX1 U7493 ( .A(n11363), .Y(n11546) );
  INVX12 U7494 ( .A(n4762), .Y(mem_wdata_D[46]) );
  OR2X1 U7495 ( .A(net113725), .B(n10444), .Y(n4762) );
  INVX12 U7496 ( .A(n4763), .Y(mem_wdata_D[47]) );
  OR2X1 U7497 ( .A(net113725), .B(n10195), .Y(n4763) );
  INVX12 U7498 ( .A(n4760), .Y(mem_wdata_D[104]) );
  OR2X1 U7499 ( .A(net113725), .B(n10817), .Y(n4760) );
  INVX12 U7500 ( .A(n4765), .Y(mem_wdata_D[105]) );
  OR2X1 U7501 ( .A(net113725), .B(n10765), .Y(n4765) );
  INVX12 U7502 ( .A(n4761), .Y(mem_wdata_D[108]) );
  OR2X1 U7503 ( .A(net113725), .B(n10789), .Y(n4761) );
  INVX12 U7504 ( .A(n4759), .Y(mem_wdata_D[110]) );
  OR2X1 U7505 ( .A(net113725), .B(n10435), .Y(n4759) );
  INVX12 U7506 ( .A(n4764), .Y(mem_wdata_D[111]) );
  OR2X1 U7507 ( .A(net113725), .B(n10186), .Y(n4764) );
  INVX12 U7508 ( .A(n4766), .Y(mem_wdata_D[112]) );
  OR2X1 U7509 ( .A(net113667), .B(n10449), .Y(n4766) );
  INVX12 U7510 ( .A(n4768), .Y(mem_wdata_D[113]) );
  OR2X1 U7511 ( .A(net113725), .B(n10595), .Y(n4768) );
  INVX12 U7512 ( .A(n4758), .Y(mem_wdata_D[45]) );
  OR2X1 U7513 ( .A(net113725), .B(n10810), .Y(n4758) );
  INVX12 U7514 ( .A(n4773), .Y(mem_wdata_D[107]) );
  INVX12 U7515 ( .A(n4776), .Y(mem_wdata_D[114]) );
  INVX12 U7516 ( .A(n4774), .Y(mem_wdata_D[116]) );
  OR2X1 U7517 ( .A(net113725), .B(n10520), .Y(n4774) );
  INVX12 U7518 ( .A(n4780), .Y(mem_wdata_D[120]) );
  INVX12 U7519 ( .A(n4782), .Y(mem_wdata_D[122]) );
  INVX12 U7520 ( .A(n4775), .Y(mem_wdata_D[123]) );
  INVX12 U7521 ( .A(n4777), .Y(mem_wdata_D[125]) );
  OR2X1 U7522 ( .A(net113725), .B(n10474), .Y(n4777) );
  NAND3BX1 U7523 ( .AN(n10251), .B(n10250), .C(n10249), .Y(n10253) );
  CLKINVX1 U7524 ( .A(n10248), .Y(n10250) );
  OR3X2 U7525 ( .A(n10243), .B(n10222), .C(n11164), .Y(n10251) );
  CLKINVX1 U7526 ( .A(n10907), .Y(n10922) );
  CLKINVX1 U7527 ( .A(n10301), .Y(n10279) );
  CLKINVX1 U7528 ( .A(n6932), .Y(n6933) );
  AND2X2 U7529 ( .A(n10245), .B(n10248), .Y(n4511) );
  CLKINVX1 U7530 ( .A(n6677), .Y(n6663) );
  CLKINVX1 U7531 ( .A(n10344), .Y(n10345) );
  CLKINVX1 U7532 ( .A(n8661), .Y(n8658) );
  CLKINVX1 U7533 ( .A(n11028), .Y(n11030) );
  CLKBUFX3 U7534 ( .A(n4933), .Y(n4935) );
  CLKINVX1 U7535 ( .A(n6473), .Y(n6475) );
  CLKBUFX3 U7536 ( .A(n10681), .Y(n5060) );
  INVX3 U7537 ( .A(n5501), .Y(n5500) );
  INVX3 U7538 ( .A(net111845), .Y(net111835) );
  CLKBUFX3 U7539 ( .A(n1840), .Y(net111845) );
  INVX3 U7540 ( .A(net111845), .Y(net111837) );
  INVX3 U7541 ( .A(n5047), .Y(n5045) );
  CLKBUFX3 U7542 ( .A(n1835), .Y(n5047) );
  INVX3 U7543 ( .A(n5047), .Y(n5046) );
  INVX3 U7544 ( .A(n5059), .Y(n5057) );
  INVX3 U7545 ( .A(n5076), .Y(n5074) );
  INVX3 U7546 ( .A(n5059), .Y(n5058) );
  INVX3 U7547 ( .A(n432), .Y(n4831) );
  INVX3 U7548 ( .A(n432), .Y(n4830) );
  INVX3 U7549 ( .A(n432), .Y(n4829) );
  INVX3 U7550 ( .A(n4623), .Y(n4850) );
  INVX3 U7551 ( .A(n4854), .Y(n4848) );
  INVX3 U7552 ( .A(n4630), .Y(n4954) );
  INVX3 U7553 ( .A(n4955), .Y(n4953) );
  INVX3 U7554 ( .A(n4955), .Y(n4952) );
  INVX3 U7555 ( .A(n5008), .Y(n5006) );
  CLKBUFX3 U7556 ( .A(n4545), .Y(n5008) );
  CLKBUFX3 U7557 ( .A(n5143), .Y(n5141) );
  CLKBUFX3 U7558 ( .A(n5408), .Y(n5402) );
  CLKBUFX3 U7559 ( .A(n9307), .Y(n4964) );
  CLKBUFX3 U7560 ( .A(n9311), .Y(n4983) );
  CLKBUFX3 U7561 ( .A(net110239), .Y(net110229) );
  CLKBUFX3 U7562 ( .A(net110239), .Y(net110231) );
  CLKBUFX3 U7563 ( .A(n11213), .Y(n5498) );
  CLKBUFX3 U7564 ( .A(n5464), .Y(n5471) );
  CLKBUFX3 U7565 ( .A(n5498), .Y(n5499) );
  NAND2X1 U7566 ( .A(n5098), .B(n5524), .Y(n10835) );
  CLKINVX1 U7567 ( .A(n4638), .Y(n5524) );
  INVX3 U7568 ( .A(n4638), .Y(n5522) );
  INVX3 U7569 ( .A(n4638), .Y(n5523) );
  CLKBUFX3 U7570 ( .A(n5937), .Y(n5626) );
  CLKBUFX3 U7571 ( .A(n5937), .Y(n5625) );
  CLKBUFX3 U7572 ( .A(n5937), .Y(n5624) );
  CLKBUFX3 U7573 ( .A(n5937), .Y(n5623) );
  CLKBUFX3 U7574 ( .A(n5937), .Y(n5622) );
  CLKBUFX3 U7575 ( .A(n5937), .Y(n5621) );
  CLKBUFX3 U7576 ( .A(n5937), .Y(n5619) );
  CLKBUFX3 U7577 ( .A(n5937), .Y(n5618) );
  CLKBUFX3 U7578 ( .A(n5937), .Y(n5617) );
  CLKBUFX3 U7579 ( .A(n5937), .Y(n5616) );
  CLKBUFX3 U7580 ( .A(n5937), .Y(n5615) );
  CLKBUFX3 U7581 ( .A(n5938), .Y(n5614) );
  CLKBUFX3 U7582 ( .A(n5938), .Y(n5613) );
  CLKBUFX3 U7583 ( .A(n5938), .Y(n5612) );
  CLKBUFX3 U7584 ( .A(n5938), .Y(n5611) );
  CLKBUFX3 U7585 ( .A(n5938), .Y(n5610) );
  CLKBUFX3 U7586 ( .A(n5938), .Y(n5609) );
  CLKBUFX3 U7587 ( .A(n5938), .Y(n5605) );
  CLKBUFX3 U7588 ( .A(n5938), .Y(n5604) );
  CLKBUFX3 U7589 ( .A(n5938), .Y(n5603) );
  CLKBUFX3 U7590 ( .A(n5939), .Y(n5602) );
  CLKBUFX3 U7591 ( .A(n5939), .Y(n5601) );
  CLKBUFX3 U7592 ( .A(n5939), .Y(n5600) );
  CLKBUFX3 U7593 ( .A(n5940), .Y(n5599) );
  CLKBUFX3 U7594 ( .A(n5939), .Y(n5598) );
  CLKBUFX3 U7595 ( .A(n5940), .Y(n5597) );
  CLKBUFX3 U7596 ( .A(n5914), .Y(n5596) );
  CLKBUFX3 U7597 ( .A(n5937), .Y(n5620) );
  CLKBUFX3 U7598 ( .A(n5938), .Y(n5606) );
  CLKBUFX3 U7599 ( .A(n5938), .Y(n5608) );
  CLKBUFX3 U7600 ( .A(n5938), .Y(n5607) );
  CLKBUFX3 U7601 ( .A(n5940), .Y(n5915) );
  CLKBUFX3 U7602 ( .A(n5940), .Y(n5916) );
  CLKBUFX3 U7603 ( .A(n5939), .Y(n5917) );
  CLKBUFX3 U7604 ( .A(rst_n), .Y(n5918) );
  CLKBUFX3 U7605 ( .A(n5922), .Y(n5919) );
  CLKBUFX3 U7606 ( .A(n5940), .Y(n5920) );
  CLKBUFX3 U7607 ( .A(n5940), .Y(n5921) );
  CLKBUFX3 U7608 ( .A(rst_n), .Y(n5922) );
  CLKBUFX3 U7609 ( .A(n5940), .Y(n5932) );
  CLKBUFX3 U7610 ( .A(n5939), .Y(n5933) );
  CLKBUFX3 U7611 ( .A(n5939), .Y(n5934) );
  CLKBUFX3 U7612 ( .A(n5939), .Y(n5935) );
  CLKBUFX3 U7613 ( .A(n5940), .Y(n5936) );
  CLKBUFX3 U7614 ( .A(n5939), .Y(n5923) );
  CLKBUFX3 U7615 ( .A(rst_n), .Y(n5924) );
  CLKBUFX3 U7616 ( .A(n5939), .Y(n5925) );
  CLKBUFX3 U7617 ( .A(rst_n), .Y(n5926) );
  CLKBUFX3 U7618 ( .A(n5940), .Y(n5927) );
  CLKBUFX3 U7619 ( .A(n5939), .Y(n5928) );
  CLKBUFX3 U7620 ( .A(n5940), .Y(n5929) );
  CLKBUFX3 U7621 ( .A(rst_n), .Y(n5930) );
  CLKBUFX3 U7622 ( .A(n5924), .Y(n5931) );
  INVX1 U7623 ( .A(n11057), .Y(n11050) );
  INVX12 U7624 ( .A(n1804), .Y(mem_wdata_D[118]) );
  INVX12 U7625 ( .A(n1806), .Y(mem_wdata_D[126]) );
  INVX12 U7626 ( .A(n1807), .Y(mem_wdata_D[127]) );
  AO22X1 U7627 ( .A0(net113445), .A1(n11458), .B0(net102346), .B1(n11489), .Y(
        n7500) );
  AO22X1 U7628 ( .A0(net113455), .A1(n11429), .B0(net113461), .B1(n11398), .Y(
        n6885) );
  AO22X1 U7629 ( .A0(net113455), .A1(n11434), .B0(net113461), .B1(n11403), .Y(
        n6977) );
  AO22X1 U7630 ( .A0(net113455), .A1(n11432), .B0(net113461), .B1(n11401), .Y(
        n6286) );
  AO22X1 U7631 ( .A0(net113447), .A1(n11464), .B0(net102346), .B1(n11495), .Y(
        n6393) );
  AO22X1 U7632 ( .A0(net113447), .A1(n11466), .B0(net102346), .B1(n11497), .Y(
        n7067) );
  AO22X1 U7633 ( .A0(net113455), .A1(n11435), .B0(net113461), .B1(n11404), .Y(
        n7068) );
  XOR2X1 U7634 ( .A(n10295), .B(n10296), .Y(n10276) );
  XOR2X1 U7635 ( .A(n10906), .B(n10905), .Y(n10918) );
  NAND2XL U7636 ( .A(n7846), .B(n8150), .Y(n7851) );
  AND2X2 U7637 ( .A(n10974), .B(n9345), .Y(n4512) );
  OA22X1 U7638 ( .A0(n10353), .A1(n10349), .B0(n10348), .B1(n10362), .Y(n10350) );
  AOI2BB1X1 U7639 ( .A0N(n10276), .A1N(n10264), .B0(n10279), .Y(n10283) );
  AND2X2 U7640 ( .A(n10279), .B(n10278), .Y(n10282) );
  AND2X2 U7641 ( .A(n4521), .B(n10216), .Y(n10219) );
  AND2X2 U7642 ( .A(n10922), .B(n10921), .Y(n10925) );
  CLKINVX1 U7643 ( .A(n6669), .Y(n6672) );
  CLKINVX1 U7644 ( .A(n8541), .Y(n8548) );
  CLKMX2X2 U7645 ( .A(n9141), .B(n4799), .S0(n6369), .Y(n6370) );
  CLKINVX1 U7646 ( .A(n6603), .Y(n6369) );
  NAND2BX1 U7647 ( .AN(n5454), .B(n11303), .Y(n9654) );
  NAND2BX1 U7648 ( .AN(n5462), .B(n11271), .Y(n9653) );
  NAND2BX1 U7649 ( .AN(n5454), .B(n11302), .Y(n9687) );
  NAND2BX1 U7650 ( .AN(n5461), .B(n11270), .Y(n9686) );
  NAND2BX1 U7651 ( .AN(n5454), .B(n11307), .Y(n10054) );
  NAND2BX1 U7652 ( .AN(n5461), .B(n11275), .Y(n10052) );
  NAND2BX1 U7653 ( .AN(n5461), .B(n11273), .Y(n9970) );
  NAND2BX1 U7654 ( .AN(n5454), .B(n11300), .Y(n9836) );
  NAND2BX1 U7655 ( .AN(n5461), .B(n11268), .Y(n9835) );
  NAND2BX1 U7656 ( .AN(n5454), .B(n11308), .Y(n10000) );
  NAND2BX1 U7657 ( .AN(n5461), .B(n11276), .Y(n9998) );
  NAND2BX1 U7658 ( .AN(n5454), .B(n11306), .Y(n10103) );
  NAND2BX1 U7659 ( .AN(n5462), .B(n11267), .Y(n9628) );
  INVX1 U7660 ( .A(n10497), .Y(n10503) );
  CLKMX2X2 U7661 ( .A(n9280), .B(n9279), .S0(n8264), .Y(n8268) );
  NAND2BX1 U7662 ( .AN(n5454), .B(n11298), .Y(n9617) );
  NAND2BX1 U7663 ( .AN(n5462), .B(n11266), .Y(n9616) );
  NAND2BX1 U7664 ( .AN(n5454), .B(n11321), .Y(n9738) );
  NAND2BX1 U7665 ( .AN(n5461), .B(n11289), .Y(n9736) );
  NAND2BXL U7666 ( .AN(n5453), .B(n11353), .Y(n9739) );
  NAND4X1 U7667 ( .A(n9783), .B(n9782), .C(n9781), .D(n9780), .Y(n10248) );
  NAND2BX1 U7668 ( .AN(n5454), .B(n11322), .Y(n9782) );
  NAND2BX1 U7669 ( .AN(n5461), .B(n11290), .Y(n9780) );
  NAND2BXL U7670 ( .AN(n5452), .B(n11354), .Y(n9783) );
  NAND2X1 U7671 ( .A(n4569), .B(n8818), .Y(n8826) );
  INVX12 U7672 ( .A(n1805), .Y(mem_wdata_D[119]) );
  NAND2BX1 U7673 ( .AN(n5454), .B(n11296), .Y(n9604) );
  NAND2BX1 U7674 ( .AN(n5462), .B(n11264), .Y(n9603) );
  NAND2BX1 U7675 ( .AN(n5454), .B(n11304), .Y(n9676) );
  NAND2BX1 U7676 ( .AN(n5461), .B(n11272), .Y(n9674) );
  INVXL U7677 ( .A(n11059), .Y(n11060) );
  AND2XL U7678 ( .A(n11058), .B(n11057), .Y(n11061) );
  INVXL U7679 ( .A(n10893), .Y(n10894) );
  CLKINVX1 U7680 ( .A(n10348), .Y(n10346) );
  NAND2BX1 U7681 ( .AN(n5454), .B(n11295), .Y(n9600) );
  NAND2BX1 U7682 ( .AN(n5461), .B(n11263), .Y(n9599) );
  NAND4X1 U7683 ( .A(n10242), .B(n10241), .C(n10240), .D(n10239), .Y(n11164)
         );
  NAND2BX1 U7684 ( .AN(n5454), .B(n11323), .Y(n10241) );
  NAND2BX1 U7685 ( .AN(n5461), .B(n11291), .Y(n10239) );
  NAND2BXL U7686 ( .AN(n5452), .B(n11355), .Y(n10242) );
  NAND4X1 U7687 ( .A(n9759), .B(n9758), .C(n9757), .D(n9756), .Y(n10222) );
  NAND2BX1 U7688 ( .AN(n5454), .B(n11325), .Y(n9758) );
  NAND2BX1 U7689 ( .AN(n5461), .B(n11293), .Y(n9756) );
  NAND2BXL U7690 ( .AN(n5452), .B(n11357), .Y(n9759) );
  NAND4X1 U7691 ( .A(n9715), .B(n9714), .C(n9713), .D(n9712), .Y(n10244) );
  NAND2BX1 U7692 ( .AN(n5454), .B(n11320), .Y(n9714) );
  NAND2BX1 U7693 ( .AN(n5461), .B(n11288), .Y(n9712) );
  NAND4X1 U7694 ( .A(n10026), .B(n10025), .C(n10024), .D(n10023), .Y(n10958)
         );
  NAND2BX1 U7695 ( .AN(n5454), .B(n11314), .Y(n10025) );
  NAND2BXL U7696 ( .AN(n5456), .B(n11250), .Y(n10024) );
  NAND4X1 U7697 ( .A(n9997), .B(n9996), .C(n9995), .D(n9994), .Y(n11028) );
  NAND2BX1 U7698 ( .AN(n5454), .B(n11313), .Y(n9996) );
  NAND2BXL U7699 ( .AN(n5456), .B(n11249), .Y(n9995) );
  NAND4X1 U7700 ( .A(n10050), .B(n10049), .C(n10048), .D(n10047), .Y(n11019)
         );
  NAND2BX1 U7701 ( .AN(n5454), .B(n11312), .Y(n10049) );
  NAND2BXL U7702 ( .AN(n5456), .B(n11248), .Y(n10048) );
  NAND4X1 U7703 ( .A(n11150), .B(n11149), .C(n11148), .D(n11147), .Y(n11218)
         );
  NAND2BX1 U7704 ( .AN(n5454), .B(n11311), .Y(n11149) );
  NAND4X1 U7705 ( .A(n10079), .B(n10078), .C(n10077), .D(n10076), .Y(n10943)
         );
  NAND2BX1 U7706 ( .AN(n5454), .B(n11310), .Y(n10078) );
  NAND2BXL U7707 ( .AN(n5456), .B(n11246), .Y(n10077) );
  INVXL U7708 ( .A(n7846), .Y(n7848) );
  INVXL U7709 ( .A(n7561), .Y(n6364) );
  NAND4X1 U7710 ( .A(n10128), .B(n10127), .C(n10126), .D(n10125), .Y(n10370)
         );
  NAND2BX1 U7711 ( .AN(n5454), .B(n11319), .Y(n10127) );
  NAND2BXL U7712 ( .AN(n5456), .B(n11255), .Y(n10126) );
  NAND4X1 U7713 ( .A(n9906), .B(n9905), .C(n9904), .D(n9903), .Y(n10356) );
  NAND2BX1 U7714 ( .AN(n5454), .B(n11318), .Y(n9905) );
  NAND4X1 U7715 ( .A(n9930), .B(n9929), .C(n9928), .D(n9927), .Y(n10337) );
  NAND2BX1 U7716 ( .AN(n5454), .B(n11317), .Y(n9929) );
  NAND2BXL U7717 ( .AN(n5456), .B(n11253), .Y(n9928) );
  NAND2BX1 U7718 ( .AN(n5454), .B(n11316), .Y(net100749) );
  NAND4X1 U7719 ( .A(n9882), .B(n9881), .C(n9880), .D(n9879), .Y(n10968) );
  NAND2BX1 U7720 ( .AN(n5454), .B(n11315), .Y(n9881) );
  INVXL U7721 ( .A(n7781), .Y(n8519) );
  INVXL U7722 ( .A(n8426), .Y(n8441) );
  NAND4X1 U7723 ( .A(n9807), .B(n9806), .C(n9805), .D(n9804), .Y(n10243) );
  NAND2BX1 U7724 ( .AN(n5454), .B(n11324), .Y(n9806) );
  NAND2BX1 U7725 ( .AN(n5461), .B(n11292), .Y(n9804) );
  NAND2BXL U7726 ( .AN(n5452), .B(n11356), .Y(n9807) );
  CLKINVX1 U7727 ( .A(n9150), .Y(n11225) );
  INVXL U7728 ( .A(n8520), .Y(n6491) );
  NAND2X1 U7729 ( .A(n9345), .B(n9572), .Y(n11359) );
  CLKINVX1 U7730 ( .A(n8911), .Y(n8912) );
  AOI2BB1XL U7731 ( .A0N(n9140), .A1N(n9139), .B0(n9138), .Y(n9149) );
  AND2XL U7732 ( .A(n10582), .B(n10581), .Y(n4526) );
  AND2XL U7733 ( .A(n3583), .B(net99693), .Y(n4530) );
  AND2XL U7734 ( .A(n3203), .B(net98932), .Y(n4541) );
  AND2XL U7735 ( .A(net99089), .B(net99090), .Y(n4542) );
  NAND2BXL U7736 ( .AN(n5456), .B(n11259), .Y(n10240) );
  NAND2BXL U7737 ( .AN(n5452), .B(n11352), .Y(n9715) );
  NAND2BXL U7738 ( .AN(n5452), .B(n11351), .Y(n10128) );
  NAND2BXL U7739 ( .AN(n5452), .B(n11350), .Y(n9906) );
  NAND2BXL U7740 ( .AN(n5453), .B(n11349), .Y(n9930) );
  NAND2BXL U7741 ( .AN(n5453), .B(n11348), .Y(net100748) );
  NAND2BXL U7742 ( .AN(n5453), .B(n11347), .Y(n9882) );
  NAND2BXL U7743 ( .AN(n5452), .B(n11346), .Y(n10026) );
  NAND2BXL U7744 ( .AN(n5452), .B(n11345), .Y(n9997) );
  NAND2BXL U7745 ( .AN(n5452), .B(n11344), .Y(n10050) );
  NAND2BXL U7746 ( .AN(n5452), .B(n11343), .Y(n11150) );
  NAND2BXL U7747 ( .AN(n5452), .B(n11342), .Y(n10079) );
  CLKINVX1 U7748 ( .A(n7356), .Y(n7358) );
  AOI21XL U7749 ( .A0(n8914), .A1(n8426), .B0(n8326), .Y(n4548) );
  AND2X2 U7750 ( .A(n5455), .B(n11297), .Y(n4549) );
  INVXL U7751 ( .A(n8920), .Y(n8264) );
  INVXL U7752 ( .A(n7709), .Y(n7036) );
  CLKINVX1 U7753 ( .A(n11309), .Y(n9946) );
  CLKINVX1 U7754 ( .A(n11277), .Y(n9945) );
  AND2XL U7755 ( .A(n3204), .B(net99042), .Y(n4558) );
  CLKINVX1 U7756 ( .A(n8543), .Y(n8544) );
  CLKINVX1 U7757 ( .A(n11230), .Y(n9608) );
  CLKINVX1 U7758 ( .A(n11294), .Y(n9610) );
  CLKINVX1 U7759 ( .A(n6676), .Y(n6662) );
  INVX1 U7760 ( .A(n11042), .Y(n11046) );
  MX2XL U7761 ( .A(n9280), .B(n9279), .S0(n8146), .Y(n8167) );
  AO22X1 U7762 ( .A0(net113447), .A1(n11478), .B0(net102346), .B1(n11509), .Y(
        n8689) );
  CLKINVX1 U7763 ( .A(n8530), .Y(n8528) );
  CLKINVX1 U7764 ( .A(n7862), .Y(n7860) );
  CLKINVX1 U7765 ( .A(n7964), .Y(n7962) );
  CLKBUFX3 U7766 ( .A(n4624), .Y(n4847) );
  CLKBUFX3 U7767 ( .A(n4624), .Y(n4846) );
  CLKBUFX3 U7768 ( .A(n4624), .Y(n4845) );
  CLKBUFX3 U7769 ( .A(n4625), .Y(n4878) );
  CLKBUFX3 U7770 ( .A(n4625), .Y(n4879) );
  CLKBUFX3 U7771 ( .A(n4621), .Y(n4887) );
  CLKBUFX3 U7772 ( .A(n4621), .Y(n4888) );
  CLKBUFX3 U7773 ( .A(n4621), .Y(n4886) );
  CLKBUFX3 U7774 ( .A(n4623), .Y(n4852) );
  CLKBUFX3 U7775 ( .A(n4628), .Y(n4960) );
  AND2X2 U7776 ( .A(n4584), .B(n4582), .Y(n4566) );
  CLKINVX1 U7777 ( .A(n11217), .Y(n5501) );
  CLKINVX1 U7778 ( .A(n10607), .Y(n5059) );
  CLKINVX1 U7779 ( .A(n10764), .Y(n5076) );
  INVXL U7780 ( .A(n7971), .Y(n7972) );
  AOI2BB1X1 U7781 ( .A0N(n8436), .A1N(n7880), .B0(n7694), .Y(n7703) );
  OA22XL U7782 ( .A0(n9007), .A1(n8910), .B0(n9004), .B1(n8909), .Y(n8919) );
  CLKBUFX3 U7783 ( .A(n4479), .Y(n4905) );
  CLKBUFX3 U7784 ( .A(n4629), .Y(n4951) );
  INVX3 U7785 ( .A(n5011), .Y(n5009) );
  INVX3 U7786 ( .A(n5011), .Y(n5010) );
  CLKBUFX3 U7787 ( .A(n1837), .Y(n5011) );
  INVX3 U7788 ( .A(n5035), .Y(n5033) );
  CLKBUFX3 U7789 ( .A(n1858), .Y(n5035) );
  INVX3 U7790 ( .A(n5029), .Y(n5027) );
  CLKBUFX3 U7791 ( .A(n4572), .Y(n5029) );
  INVX3 U7792 ( .A(n5020), .Y(n5018) );
  CLKBUFX3 U7793 ( .A(n1853), .Y(n5020) );
  INVX3 U7794 ( .A(n5026), .Y(n5024) );
  CLKBUFX3 U7795 ( .A(n1856), .Y(n5026) );
  INVX3 U7796 ( .A(n5088), .Y(n5086) );
  CLKBUFX3 U7797 ( .A(n1849), .Y(n5088) );
  INVX3 U7798 ( .A(n5082), .Y(n5080) );
  CLKBUFX3 U7799 ( .A(n4573), .Y(n5082) );
  INVX3 U7800 ( .A(n5053), .Y(n5051) );
  CLKBUFX3 U7801 ( .A(n4571), .Y(n5053) );
  INVX3 U7802 ( .A(n5091), .Y(n5089) );
  CLKBUFX3 U7803 ( .A(n1838), .Y(n5091) );
  INVX3 U7804 ( .A(n5070), .Y(n5068) );
  CLKBUFX3 U7805 ( .A(n1839), .Y(n5070) );
  INVX3 U7806 ( .A(n5035), .Y(n5034) );
  INVX3 U7807 ( .A(n5029), .Y(n5028) );
  INVX3 U7808 ( .A(n5020), .Y(n5019) );
  INVX3 U7809 ( .A(n5026), .Y(n5025) );
  INVX3 U7810 ( .A(n5088), .Y(n5087) );
  INVX3 U7811 ( .A(n5082), .Y(n5081) );
  INVX3 U7812 ( .A(n5053), .Y(n5052) );
  INVX3 U7813 ( .A(n5091), .Y(n5090) );
  INVX3 U7814 ( .A(n5070), .Y(n5069) );
  INVX3 U7815 ( .A(n5023), .Y(n5021) );
  CLKBUFX3 U7816 ( .A(n1855), .Y(n5023) );
  INVX3 U7817 ( .A(n5050), .Y(n5048) );
  CLKBUFX3 U7818 ( .A(n1836), .Y(n5050) );
  INVX3 U7819 ( .A(n5056), .Y(n5054) );
  CLKBUFX3 U7820 ( .A(n1852), .Y(n5056) );
  INVX3 U7821 ( .A(n5085), .Y(n5083) );
  CLKBUFX3 U7822 ( .A(n1857), .Y(n5085) );
  INVX3 U7823 ( .A(n5079), .Y(n5077) );
  CLKBUFX3 U7824 ( .A(n1843), .Y(n5079) );
  INVX3 U7825 ( .A(n5005), .Y(n5003) );
  CLKBUFX3 U7826 ( .A(n1842), .Y(n5005) );
  INVX3 U7827 ( .A(n5101), .Y(n5099) );
  CLKBUFX3 U7828 ( .A(n1854), .Y(n5101) );
  INVX3 U7829 ( .A(n5023), .Y(n5022) );
  INVX3 U7830 ( .A(n5050), .Y(n5049) );
  INVX3 U7831 ( .A(n5056), .Y(n5055) );
  INVX3 U7832 ( .A(n5085), .Y(n5084) );
  INVX3 U7833 ( .A(n5079), .Y(n5078) );
  INVX3 U7834 ( .A(n5005), .Y(n5004) );
  INVX3 U7835 ( .A(n5101), .Y(n5100) );
  INVX3 U7836 ( .A(n5017), .Y(n5015) );
  INVX3 U7837 ( .A(n5017), .Y(n5016) );
  INVX3 U7838 ( .A(n5041), .Y(n5039) );
  CLKBUFX3 U7839 ( .A(n223), .Y(n5041) );
  INVX3 U7840 ( .A(n5094), .Y(n5092) );
  CLKBUFX3 U7841 ( .A(n1841), .Y(n5094) );
  INVX3 U7842 ( .A(n5041), .Y(n5040) );
  INVX3 U7843 ( .A(n5094), .Y(n5093) );
  NAND2X1 U7844 ( .A(n4707), .B(n3787), .Y(n7864) );
  INVX3 U7845 ( .A(n5038), .Y(n5036) );
  CLKBUFX3 U7846 ( .A(n1995), .Y(n5038) );
  INVX3 U7847 ( .A(n5038), .Y(n5037) );
  INVX3 U7848 ( .A(n5073), .Y(n5071) );
  CLKBUFX3 U7849 ( .A(n222), .Y(n5073) );
  INVX3 U7850 ( .A(n5073), .Y(n5072) );
  INVX3 U7851 ( .A(n5067), .Y(n5065) );
  CLKBUFX3 U7852 ( .A(n1834), .Y(n5067) );
  INVX3 U7853 ( .A(n5014), .Y(n5012) );
  CLKBUFX3 U7854 ( .A(n1850), .Y(n5014) );
  INVX3 U7855 ( .A(n5032), .Y(n5030) );
  INVX3 U7856 ( .A(n5044), .Y(n5042) );
  CLKBUFX3 U7857 ( .A(n1851), .Y(n5044) );
  INVX3 U7858 ( .A(n1834), .Y(n5066) );
  INVX3 U7859 ( .A(n5014), .Y(n5013) );
  INVX3 U7860 ( .A(n5032), .Y(n5031) );
  CLKBUFX3 U7861 ( .A(n4574), .Y(n5032) );
  INVX3 U7862 ( .A(n5044), .Y(n5043) );
  CLKINVX1 U7863 ( .A(n7777), .Y(n7858) );
  CLKINVX1 U7864 ( .A(n8929), .Y(n8903) );
  CLKBUFX3 U7865 ( .A(n11161), .Y(n5464) );
  CLKINVX1 U7866 ( .A(n9181), .Y(n9185) );
  CLKBUFX3 U7867 ( .A(n4481), .Y(n4919) );
  CLKBUFX3 U7868 ( .A(n4487), .Y(n4934) );
  CLKBUFX3 U7869 ( .A(n4485), .Y(n4918) );
  CLKBUFX3 U7870 ( .A(n4484), .Y(n4941) );
  CLKBUFX3 U7871 ( .A(n4484), .Y(n4940) );
  CLKBUFX3 U7872 ( .A(n4487), .Y(n4933) );
  CLKBUFX3 U7873 ( .A(n4480), .Y(n4929) );
  CLKBUFX3 U7874 ( .A(n4484), .Y(n4942) );
  CLKBUFX3 U7875 ( .A(n9308), .Y(n4970) );
  CLKBUFX3 U7876 ( .A(net102036), .Y(net113047) );
  CLKBUFX3 U7877 ( .A(n4625), .Y(n4880) );
  CLKINVX1 U7878 ( .A(net113081), .Y(net113079) );
  CLKINVX1 U7879 ( .A(net112729), .Y(net114085) );
  CLKINVX1 U7880 ( .A(n11511), .Y(n10474) );
  CLKINVX1 U7881 ( .A(n11500), .Y(n10608) );
  CLKINVX1 U7882 ( .A(n11493), .Y(n10777) );
  CLKINVX1 U7883 ( .A(n11494), .Y(n10789) );
  CLKINVX1 U7884 ( .A(n11165), .Y(n9688) );
  CLKBUFX3 U7885 ( .A(\i_MIPS/Register/n147 ), .Y(n5585) );
  CLKBUFX3 U7886 ( .A(\i_MIPS/Register/n147 ), .Y(n5586) );
  CLKBUFX3 U7887 ( .A(\i_MIPS/Register/n146 ), .Y(n5583) );
  CLKBUFX3 U7888 ( .A(\i_MIPS/Register/n146 ), .Y(n5584) );
  CLKBUFX3 U7889 ( .A(\i_MIPS/Register/n145 ), .Y(n5581) );
  CLKBUFX3 U7890 ( .A(\i_MIPS/Register/n145 ), .Y(n5582) );
  CLKBUFX3 U7891 ( .A(\i_MIPS/Register/n144 ), .Y(n5579) );
  CLKBUFX3 U7892 ( .A(\i_MIPS/Register/n144 ), .Y(n5580) );
  CLKBUFX3 U7893 ( .A(\i_MIPS/Register/n143 ), .Y(n5577) );
  CLKBUFX3 U7894 ( .A(\i_MIPS/Register/n143 ), .Y(n5578) );
  CLKBUFX3 U7895 ( .A(\i_MIPS/Register/n142 ), .Y(n5575) );
  CLKBUFX3 U7896 ( .A(\i_MIPS/Register/n142 ), .Y(n5576) );
  CLKBUFX3 U7897 ( .A(\i_MIPS/Register/n141 ), .Y(n5573) );
  CLKBUFX3 U7898 ( .A(\i_MIPS/Register/n141 ), .Y(n5574) );
  CLKBUFX3 U7899 ( .A(\i_MIPS/Register/n139 ), .Y(n5571) );
  CLKBUFX3 U7900 ( .A(\i_MIPS/Register/n139 ), .Y(n5572) );
  CLKBUFX3 U7901 ( .A(\i_MIPS/Register/n138 ), .Y(n5569) );
  CLKBUFX3 U7902 ( .A(\i_MIPS/Register/n138 ), .Y(n5570) );
  CLKBUFX3 U7903 ( .A(\i_MIPS/Register/n137 ), .Y(n5567) );
  CLKBUFX3 U7904 ( .A(\i_MIPS/Register/n137 ), .Y(n5568) );
  CLKBUFX3 U7905 ( .A(\i_MIPS/Register/n136 ), .Y(n5565) );
  CLKBUFX3 U7906 ( .A(\i_MIPS/Register/n136 ), .Y(n5566) );
  CLKBUFX3 U7907 ( .A(\i_MIPS/Register/n135 ), .Y(n5563) );
  CLKBUFX3 U7908 ( .A(\i_MIPS/Register/n135 ), .Y(n5564) );
  CLKBUFX3 U7909 ( .A(\i_MIPS/Register/n134 ), .Y(n5561) );
  CLKBUFX3 U7910 ( .A(\i_MIPS/Register/n134 ), .Y(n5562) );
  CLKBUFX3 U7911 ( .A(\i_MIPS/Register/n133 ), .Y(n5559) );
  CLKBUFX3 U7912 ( .A(\i_MIPS/Register/n133 ), .Y(n5560) );
  CLKBUFX3 U7913 ( .A(\i_MIPS/Register/n132 ), .Y(n5557) );
  CLKBUFX3 U7914 ( .A(\i_MIPS/Register/n132 ), .Y(n5558) );
  CLKBUFX3 U7915 ( .A(\i_MIPS/Register/n130 ), .Y(n5555) );
  CLKBUFX3 U7916 ( .A(\i_MIPS/Register/n130 ), .Y(n5556) );
  CLKBUFX3 U7917 ( .A(\i_MIPS/Register/n129 ), .Y(n5553) );
  CLKBUFX3 U7918 ( .A(\i_MIPS/Register/n129 ), .Y(n5554) );
  CLKBUFX3 U7919 ( .A(\i_MIPS/Register/n128 ), .Y(n5551) );
  CLKBUFX3 U7920 ( .A(\i_MIPS/Register/n128 ), .Y(n5552) );
  CLKBUFX3 U7921 ( .A(\i_MIPS/Register/n127 ), .Y(n5549) );
  CLKBUFX3 U7922 ( .A(\i_MIPS/Register/n127 ), .Y(n5550) );
  CLKBUFX3 U7923 ( .A(\i_MIPS/Register/n126 ), .Y(n5547) );
  CLKBUFX3 U7924 ( .A(\i_MIPS/Register/n126 ), .Y(n5548) );
  CLKBUFX3 U7925 ( .A(\i_MIPS/Register/n125 ), .Y(n5545) );
  CLKBUFX3 U7926 ( .A(\i_MIPS/Register/n125 ), .Y(n5546) );
  CLKBUFX3 U7927 ( .A(\i_MIPS/Register/n124 ), .Y(n5543) );
  CLKBUFX3 U7928 ( .A(\i_MIPS/Register/n124 ), .Y(n5544) );
  CLKBUFX3 U7929 ( .A(\i_MIPS/Register/n123 ), .Y(n5541) );
  CLKBUFX3 U7930 ( .A(\i_MIPS/Register/n123 ), .Y(n5542) );
  CLKBUFX3 U7931 ( .A(\i_MIPS/Register/n121 ), .Y(n5539) );
  CLKBUFX3 U7932 ( .A(\i_MIPS/Register/n121 ), .Y(n5540) );
  CLKBUFX3 U7933 ( .A(\i_MIPS/Register/n112 ), .Y(n5531) );
  CLKBUFX3 U7934 ( .A(\i_MIPS/Register/n112 ), .Y(n5532) );
  CLKBUFX3 U7935 ( .A(\i_MIPS/Register/n108 ), .Y(n5527) );
  CLKBUFX3 U7936 ( .A(\i_MIPS/Register/n108 ), .Y(n5528) );
  CLKBUFX3 U7937 ( .A(\i_MIPS/Register/n106 ), .Y(n5525) );
  CLKBUFX3 U7938 ( .A(\i_MIPS/Register/n106 ), .Y(n5526) );
  CLKBUFX3 U7939 ( .A(\i_MIPS/Register/n116 ), .Y(n5535) );
  CLKBUFX3 U7940 ( .A(\i_MIPS/Register/n116 ), .Y(n5536) );
  CLKBUFX3 U7941 ( .A(\i_MIPS/Register/n114 ), .Y(n5533) );
  CLKBUFX3 U7942 ( .A(\i_MIPS/Register/n114 ), .Y(n5534) );
  CLKBUFX3 U7943 ( .A(\i_MIPS/Register/n110 ), .Y(n5529) );
  CLKBUFX3 U7944 ( .A(\i_MIPS/Register/n110 ), .Y(n5530) );
  CLKBUFX3 U7945 ( .A(n10836), .Y(n5097) );
  CLKBUFX3 U7946 ( .A(n10836), .Y(n5098) );
  CLKBUFX3 U7947 ( .A(\i_MIPS/Register/n118 ), .Y(n5537) );
  CLKBUFX3 U7948 ( .A(\i_MIPS/Register/n118 ), .Y(n5538) );
  CLKBUFX3 U7949 ( .A(n5940), .Y(n5937) );
  CLKBUFX3 U7950 ( .A(n5940), .Y(n5938) );
  AND2XL U7951 ( .A(n6632), .B(n6936), .Y(n6373) );
  AND2XL U7952 ( .A(n7180), .B(n7183), .Y(n6867) );
  INVX12 U7953 ( .A(n1808), .Y(mem_addr_D[18]) );
  AOI21X2 U7954 ( .A0(n10137), .A1(n10139), .B0(n10136), .Y(n10519) );
  NOR2XL U7955 ( .A(n4488), .B(n11168), .Y(n10136) );
  OAI21XL U7956 ( .A0(n11548), .A1(n11515), .B0(n4488), .Y(n10137) );
  OA22X1 U7957 ( .A0(net112493), .A1(n2810), .B0(net112369), .B1(n818), .Y(
        n9058) );
  OA22X1 U7958 ( .A0(net112239), .A1(n2811), .B0(net112161), .B1(n819), .Y(
        n9057) );
  OA22X1 U7959 ( .A0(net112485), .A1(n1249), .B0(net112361), .B1(n2860), .Y(
        n8490) );
  OA22X1 U7960 ( .A0(net112073), .A1(n1250), .B0(net111949), .B1(n2861), .Y(
        n8488) );
  CLKMX2X2 U7961 ( .A(n7018), .B(n7017), .S0(net108963), .Y(net105929) );
  CLKMX2X2 U7962 ( .A(n7692), .B(n7691), .S0(net108963), .Y(net104704) );
  OA22XL U7963 ( .A0(net112241), .A1(n1559), .B0(net112159), .B1(n3172), .Y(
        n7719) );
  OA22XL U7964 ( .A0(net112673), .A1(n1560), .B0(net112571), .B1(n3173), .Y(
        n7721) );
  OA22XL U7965 ( .A0(net112241), .A1(n1561), .B0(net112159), .B1(n3174), .Y(
        n7727) );
  OA22XL U7966 ( .A0(net112673), .A1(n1562), .B0(net112571), .B1(n3175), .Y(
        n7729) );
  OA22X1 U7967 ( .A0(net112489), .A1(n1251), .B0(net112303), .B1(n2862), .Y(
        n8849) );
  OA22X1 U7968 ( .A0(net112671), .A1(n1252), .B0(net112569), .B1(n2863), .Y(
        n9047) );
  OA22X1 U7969 ( .A0(net112491), .A1(n1253), .B0(net112367), .B1(n2864), .Y(
        n9046) );
  OA22X1 U7970 ( .A0(net112239), .A1(n2812), .B0(net112153), .B1(n820), .Y(
        n9045) );
  OA22X1 U7971 ( .A0(net112671), .A1(n1254), .B0(net112569), .B1(n2865), .Y(
        n9055) );
  OA22X1 U7972 ( .A0(net112493), .A1(n1255), .B0(net112369), .B1(n2866), .Y(
        n9054) );
  OA22X1 U7973 ( .A0(net112239), .A1(n1256), .B0(net112161), .B1(n2867), .Y(
        n9053) );
  OA22X1 U7974 ( .A0(net112671), .A1(n1257), .B0(net112569), .B1(n2868), .Y(
        n8960) );
  OA22X1 U7975 ( .A0(net112491), .A1(n1258), .B0(net112367), .B1(n2869), .Y(
        n8959) );
  OA22X1 U7976 ( .A0(net112239), .A1(n2813), .B0(net112153), .B1(n821), .Y(
        n8958) );
  OA22X1 U7977 ( .A0(net112481), .A1(n1259), .B0(net112357), .B1(n2870), .Y(
        n8290) );
  OA22X1 U7978 ( .A0(net112235), .A1(n1260), .B0(net112153), .B1(n2871), .Y(
        n8289) );
  OA22X1 U7979 ( .A0(net112671), .A1(n1261), .B0(net112569), .B1(n2872), .Y(
        n9094) );
  OA22X1 U7980 ( .A0(net112239), .A1(n1263), .B0(net112153), .B1(n2874), .Y(
        n9092) );
  OA22X1 U7981 ( .A0(net112671), .A1(n1264), .B0(net112569), .B1(n2875), .Y(
        n9086) );
  OA22X1 U7982 ( .A0(net112239), .A1(n1266), .B0(net112159), .B1(n2877), .Y(
        n9084) );
  OA22X1 U7983 ( .A0(net112681), .A1(n1267), .B0(net112565), .B1(n2878), .Y(
        n8765) );
  OA22X1 U7984 ( .A0(net112487), .A1(n1268), .B0(net112363), .B1(n2879), .Y(
        n8764) );
  OA22X1 U7985 ( .A0(net112491), .A1(n1269), .B0(net112367), .B1(n2880), .Y(
        n8967) );
  OA22X1 U7986 ( .A0(net112671), .A1(n1270), .B0(net112569), .B1(n2881), .Y(
        n8968) );
  OA22X1 U7987 ( .A0(net112239), .A1(n1271), .B0(net112153), .B1(n2882), .Y(
        n8966) );
  OA22X1 U7988 ( .A0(net112667), .A1(n1272), .B0(net112573), .B1(n2883), .Y(
        n7318) );
  OA22X1 U7989 ( .A0(net112467), .A1(n1273), .B0(net112343), .B1(n2884), .Y(
        n7317) );
  OA22X1 U7990 ( .A0(net112245), .A1(n1228), .B0(net112163), .B1(n2885), .Y(
        n7316) );
  OA22X1 U7991 ( .A0(net112489), .A1(n1274), .B0(net112303), .B1(n2886), .Y(
        n8772) );
  OA22X1 U7992 ( .A0(net112665), .A1(n1275), .B0(net112565), .B1(n2887), .Y(
        n8773) );
  OA22X1 U7993 ( .A0(net112237), .A1(n1276), .B0(net112155), .B1(n2888), .Y(
        n8771) );
  OA22X1 U7994 ( .A0(net112679), .A1(n1277), .B0(net112573), .B1(n2889), .Y(
        n7326) );
  OA22X1 U7995 ( .A0(net112467), .A1(n1278), .B0(net112343), .B1(n2890), .Y(
        n7325) );
  OA22X1 U7996 ( .A0(net112681), .A1(n1279), .B0(net112575), .B1(n2891), .Y(
        n7234) );
  OA22X1 U7997 ( .A0(net112465), .A1(n1280), .B0(net112341), .B1(n2892), .Y(
        n7233) );
  OA22X1 U7998 ( .A0(net112245), .A1(n1281), .B0(net112163), .B1(n2893), .Y(
        n7232) );
  OA22X1 U7999 ( .A0(net112463), .A1(n1282), .B0(net112339), .B1(n2894), .Y(
        n7143) );
  OA22X1 U8000 ( .A0(net112465), .A1(n1283), .B0(net112341), .B1(n2895), .Y(
        n7241) );
  OA22X1 U8001 ( .A0(net112665), .A1(n1284), .B0(net112563), .B1(n2896), .Y(
        n8194) );
  OA22X1 U8002 ( .A0(net112483), .A1(n1285), .B0(net112355), .B1(n2897), .Y(
        n8193) );
  OA22X1 U8003 ( .A0(net112679), .A1(n1286), .B0(net112575), .B1(n2898), .Y(
        n7152) );
  OA22X1 U8004 ( .A0(net112465), .A1(n1287), .B0(net112341), .B1(n2899), .Y(
        n7151) );
  OA22X1 U8005 ( .A0(net112245), .A1(n1288), .B0(net112161), .B1(n2900), .Y(
        n7150) );
  OA22X1 U8006 ( .A0(net112679), .A1(n1289), .B0(net112573), .B1(n2901), .Y(
        n7404) );
  OA22X1 U8007 ( .A0(net112469), .A1(n1290), .B0(net112345), .B1(n2902), .Y(
        n7403) );
  OA22X1 U8008 ( .A0(net112481), .A1(n1291), .B0(net112357), .B1(n2903), .Y(
        n8201) );
  OA22X1 U8009 ( .A0(net112665), .A1(n1292), .B0(net112563), .B1(n2904), .Y(
        n8202) );
  OA22X1 U8010 ( .A0(net112233), .A1(n1293), .B0(net112151), .B1(n2905), .Y(
        n8200) );
  OA22X1 U8011 ( .A0(net112679), .A1(n1294), .B0(net112573), .B1(n2906), .Y(
        n7396) );
  OA22X1 U8012 ( .A0(net112467), .A1(n1295), .B0(net112343), .B1(n2907), .Y(
        n7395) );
  OA22X1 U8013 ( .A0(net112483), .A1(n1296), .B0(net112359), .B1(n2908), .Y(
        n8395) );
  OA22X1 U8014 ( .A0(net112235), .A1(n1297), .B0(net112153), .B1(n2909), .Y(
        n8394) );
  OA22X1 U8015 ( .A0(net112665), .A1(n1298), .B0(net112565), .B1(n2910), .Y(
        n8684) );
  OA22X1 U8016 ( .A0(net112483), .A1(n1299), .B0(net112359), .B1(n2911), .Y(
        n8387) );
  OA22X1 U8017 ( .A0(net112235), .A1(n1300), .B0(net112153), .B1(n2912), .Y(
        n8386) );
  OA22X1 U8018 ( .A0(net112487), .A1(n1301), .B0(net112363), .B1(n2913), .Y(
        n8675) );
  OA22X1 U8019 ( .A0(net112665), .A1(n1302), .B0(net112565), .B1(n2914), .Y(
        n8676) );
  OA22X1 U8020 ( .A0(net112469), .A1(n1303), .B0(net112351), .B1(n2915), .Y(
        n7809) );
  OA22XL U8021 ( .A0(net112673), .A1(n1563), .B0(net112571), .B1(n3176), .Y(
        n7644) );
  OA22X1 U8022 ( .A0(net112473), .A1(n1304), .B0(net112349), .B1(n2916), .Y(
        n7643) );
  OA22XL U8023 ( .A0(net112241), .A1(n1564), .B0(net112159), .B1(n3177), .Y(
        n7642) );
  OA22XL U8024 ( .A0(net112673), .A1(n1565), .B0(net112571), .B1(n3178), .Y(
        n7636) );
  OA22X1 U8025 ( .A0(net112471), .A1(n1305), .B0(net112347), .B1(n2917), .Y(
        n7635) );
  OA22XL U8026 ( .A0(net112241), .A1(n1566), .B0(net112159), .B1(n3179), .Y(
        n7634) );
  OA22X2 U8027 ( .A0(net112455), .A1(n952), .B0(net112351), .B1(n2477), .Y(
        n7817) );
  OA22XL U8028 ( .A0(net112231), .A1(n1567), .B0(net112159), .B1(n3180), .Y(
        n7816) );
  OA22X1 U8029 ( .A0(net112485), .A1(n1306), .B0(net112361), .B1(n2918), .Y(
        n8592) );
  OA22X1 U8030 ( .A0(net112665), .A1(n1307), .B0(net112565), .B1(n2919), .Y(
        n8593) );
  OA22X1 U8031 ( .A0(net112237), .A1(n1308), .B0(net112155), .B1(n2920), .Y(
        n8591) );
  OA22X1 U8032 ( .A0(net112457), .A1(n1309), .B0(net112333), .B1(n2921), .Y(
        n6716) );
  OA22X1 U8033 ( .A0(net112679), .A1(n1310), .B0(net112577), .B1(n2922), .Y(
        n6717) );
  OA22X1 U8034 ( .A0(net112457), .A1(n1311), .B0(net112333), .B1(n2923), .Y(
        n6708) );
  OA22X1 U8035 ( .A0(net112679), .A1(n1312), .B0(net112577), .B1(n2924), .Y(
        n6709) );
  OA22X1 U8036 ( .A0(net112233), .A1(n1313), .B0(net112165), .B1(n2925), .Y(
        n6707) );
  OA22X1 U8037 ( .A0(net112665), .A1(n1314), .B0(net112563), .B1(n2926), .Y(
        n8113) );
  OA22X1 U8038 ( .A0(net112235), .A1(n1315), .B0(net112153), .B1(n2927), .Y(
        n8583) );
  OA22X1 U8039 ( .A0(net112477), .A1(n1316), .B0(net112353), .B1(n2928), .Y(
        n8019) );
  OA22X1 U8040 ( .A0(net112233), .A1(n1317), .B0(net112151), .B1(n2929), .Y(
        n8018) );
  OA22X1 U8041 ( .A0(net112665), .A1(n1318), .B0(net112563), .B1(n2930), .Y(
        n8020) );
  OA22X1 U8042 ( .A0(net112483), .A1(n1319), .B0(net112355), .B1(n2931), .Y(
        n8104) );
  OA22X1 U8043 ( .A0(net112665), .A1(n1320), .B0(net112563), .B1(n2932), .Y(
        n8105) );
  OA22X1 U8044 ( .A0(net112477), .A1(n1321), .B0(net112353), .B1(n2933), .Y(
        n8011) );
  OA22X1 U8045 ( .A0(net112233), .A1(n1322), .B0(net112151), .B1(n2934), .Y(
        n8010) );
  OA22X1 U8046 ( .A0(net112665), .A1(n1323), .B0(net112563), .B1(n2935), .Y(
        n8012) );
  NAND4X1 U8047 ( .A(n7915), .B(n7914), .C(n7913), .D(n7912), .Y(n11438) );
  OA22X2 U8048 ( .A0(net112663), .A1(n954), .B0(net112561), .B1(n2479), .Y(
        n7915) );
  OA22X2 U8049 ( .A0(net112471), .A1(n955), .B0(net112351), .B1(n2480), .Y(
        n7914) );
  OA22XL U8050 ( .A0(net112231), .A1(n1568), .B0(net112145), .B1(n3181), .Y(
        n7913) );
  OA22X1 U8051 ( .A0(net112665), .A1(n1324), .B0(net112563), .B1(n2936), .Y(
        n7923) );
  OA22X1 U8052 ( .A0(net112477), .A1(n1325), .B0(net112353), .B1(n2937), .Y(
        n7922) );
  OA22X1 U8053 ( .A0(net112233), .A1(n2814), .B0(net112151), .B1(n822), .Y(
        n7921) );
  OA22X1 U8054 ( .A0(net112681), .A1(n1326), .B0(net112565), .B1(n2938), .Y(
        n6530) );
  OA22X1 U8055 ( .A0(net112455), .A1(n1327), .B0(net112331), .B1(n2939), .Y(
        n6529) );
  OA22X1 U8056 ( .A0(net112681), .A1(n1328), .B0(net112565), .B1(n2940), .Y(
        n6538) );
  OA22X1 U8057 ( .A0(net112457), .A1(n1329), .B0(net112333), .B1(n2941), .Y(
        n6537) );
  OA22X1 U8058 ( .A0(net112237), .A1(n1330), .B0(net112153), .B1(n2942), .Y(
        n6536) );
  OA22X1 U8059 ( .A0(net112485), .A1(n1331), .B0(net112361), .B1(n2943), .Y(
        n8486) );
  OA22X1 U8060 ( .A0(net112235), .A1(n1332), .B0(net112153), .B1(n2944), .Y(
        n8485) );
  OA22X1 U8061 ( .A0(net112667), .A1(n1333), .B0(net112565), .B1(n2945), .Y(
        n8487) );
  OA22X1 U8062 ( .A0(net112483), .A1(n1334), .B0(net112359), .B1(n2946), .Y(
        n8478) );
  OA22X1 U8063 ( .A0(net112235), .A1(n1335), .B0(net112153), .B1(n2947), .Y(
        n8477) );
  OA22X1 U8064 ( .A0(net112667), .A1(n1336), .B0(net112565), .B1(n2948), .Y(
        n8479) );
  OA22X1 U8065 ( .A0(net112469), .A1(n1337), .B0(net112345), .B1(n2949), .Y(
        n7494) );
  OA22X1 U8066 ( .A0(net112245), .A1(n1338), .B0(net112163), .B1(n2950), .Y(
        n7493) );
  OA22X1 U8067 ( .A0(net112057), .A1(n1339), .B0(net111933), .B1(n2951), .Y(
        n7492) );
  OA22X1 U8068 ( .A0(net112469), .A1(n1340), .B0(net112345), .B1(n2952), .Y(
        n7486) );
  OA22X1 U8069 ( .A0(net112679), .A1(n1341), .B0(net112573), .B1(n2953), .Y(
        n7487) );
  OA22X1 U8070 ( .A0(net112471), .A1(n1342), .B0(net112347), .B1(n2954), .Y(
        net105021) );
  OA22XL U8071 ( .A0(net112241), .A1(n1569), .B0(net112159), .B1(n3182), .Y(
        net105022) );
  OA22X1 U8072 ( .A0(net112059), .A1(n1343), .B0(net111935), .B1(n2955), .Y(
        net105023) );
  OA22X1 U8073 ( .A0(net112455), .A1(n1344), .B0(net112331), .B1(n2956), .Y(
        n6387) );
  OA22X1 U8074 ( .A0(net112681), .A1(n1345), .B0(net112565), .B1(n2957), .Y(
        n6388) );
  OA22X1 U8075 ( .A0(net112471), .A1(n1346), .B0(net112347), .B1(n2958), .Y(
        net105045) );
  OA22X1 U8076 ( .A0(net112245), .A1(n1347), .B0(net112161), .B1(n2959), .Y(
        net105046) );
  OA22X1 U8077 ( .A0(net112667), .A1(n1348), .B0(net112573), .B1(n2960), .Y(
        net105044) );
  OA22X1 U8078 ( .A0(net112461), .A1(n1349), .B0(net112337), .B1(n2961), .Y(
        n6878) );
  OA22X1 U8079 ( .A0(net112235), .A1(n1229), .B0(net112165), .B1(n2962), .Y(
        n6877) );
  OA22X1 U8080 ( .A0(net112679), .A1(n1350), .B0(net112577), .B1(n2963), .Y(
        n6879) );
  OA22X1 U8081 ( .A0(net112453), .A1(n1351), .B0(net112329), .B1(n2964), .Y(
        n6279) );
  OA22X1 U8082 ( .A0(net112681), .A1(n1352), .B0(net112577), .B1(n2965), .Y(
        n6280) );
  OA22X1 U8083 ( .A0(net112459), .A1(n1353), .B0(net112335), .B1(n2966), .Y(
        n6870) );
  OA22X1 U8084 ( .A0(net112679), .A1(n1354), .B0(net112577), .B1(n2967), .Y(
        n6871) );
  OA22X1 U8085 ( .A0(net112453), .A1(n1355), .B0(net112329), .B1(n2968), .Y(
        n6271) );
  OA22X1 U8086 ( .A0(net112681), .A1(n1356), .B0(net112577), .B1(n2969), .Y(
        n6272) );
  OA22X1 U8087 ( .A0(net112459), .A1(n1357), .B0(net112335), .B1(n2970), .Y(
        n6795) );
  OA22X1 U8088 ( .A0(net112679), .A1(n1358), .B0(net112577), .B1(n2971), .Y(
        n6796) );
  OA22X1 U8089 ( .A0(net112665), .A1(n1359), .B0(net112565), .B1(n2972), .Y(
        n8854) );
  OA22X1 U8090 ( .A0(net112489), .A1(n1360), .B0(net112303), .B1(n2973), .Y(
        n8853) );
  OA22X1 U8091 ( .A0(net112237), .A1(n2815), .B0(net112155), .B1(n823), .Y(
        n8852) );
  OA22X1 U8092 ( .A0(net112491), .A1(n2816), .B0(net112367), .B1(n824), .Y(
        n9050) );
  OA22X1 U8093 ( .A0(net112671), .A1(n2817), .B0(net112569), .B1(n825), .Y(
        n9051) );
  OA22X1 U8094 ( .A0(net112239), .A1(n2818), .B0(net112161), .B1(n826), .Y(
        n9049) );
  OA22X1 U8095 ( .A0(net112671), .A1(n1361), .B0(net112569), .B1(n2974), .Y(
        n9090) );
  OA22X1 U8096 ( .A0(net112239), .A1(n1363), .B0(net112163), .B1(n2976), .Y(
        n9088) );
  OA22X1 U8097 ( .A0(net112491), .A1(n2819), .B0(net112367), .B1(n827), .Y(
        n8963) );
  OA22X1 U8098 ( .A0(net112671), .A1(n2820), .B0(net112569), .B1(n828), .Y(
        n8964) );
  OA22X1 U8099 ( .A0(net112239), .A1(n2821), .B0(net112163), .B1(n829), .Y(
        n8962) );
  OA22X1 U8100 ( .A0(net112657), .A1(n1365), .B0(net112573), .B1(n2978), .Y(
        n7330) );
  OA22X1 U8101 ( .A0(net112481), .A1(n1366), .B0(net112357), .B1(n2979), .Y(
        n8294) );
  OA22X1 U8102 ( .A0(net112667), .A1(n1367), .B0(net112565), .B1(n2980), .Y(
        n8295) );
  OA22X1 U8103 ( .A0(net112235), .A1(n2822), .B0(net112153), .B1(n830), .Y(
        n8293) );
  OA22X1 U8104 ( .A0(net112665), .A1(n2823), .B0(net112565), .B1(n831), .Y(
        n8769) );
  OA22X1 U8105 ( .A0(net112657), .A1(n1368), .B0(net112573), .B1(n2981), .Y(
        n7322) );
  OA22X1 U8106 ( .A0(net112673), .A1(n1369), .B0(net112575), .B1(n2982), .Y(
        n7238) );
  OA22X1 U8107 ( .A0(net112469), .A1(n1372), .B0(net112345), .B1(n2985), .Y(
        n7407) );
  OA22X1 U8108 ( .A0(net112679), .A1(n1373), .B0(net112573), .B1(n2986), .Y(
        n7408) );
  OA22X1 U8109 ( .A0(net112463), .A1(n1374), .B0(net112339), .B1(n2987), .Y(
        n7147) );
  OA22X1 U8110 ( .A0(net112483), .A1(n1375), .B0(net112355), .B1(n2988), .Y(
        n8197) );
  OA22X1 U8111 ( .A0(net112665), .A1(n1376), .B0(net112563), .B1(n2989), .Y(
        n8198) );
  OA22X1 U8112 ( .A0(net112233), .A1(n1377), .B0(net112151), .B1(n2990), .Y(
        n8196) );
  OA22X1 U8113 ( .A0(net112657), .A1(n1378), .B0(net112573), .B1(n2991), .Y(
        n7400) );
  OA22X1 U8114 ( .A0(net112467), .A1(n1379), .B0(net112343), .B1(n2992), .Y(
        n7399) );
  OA22XL U8115 ( .A0(net112673), .A1(n1570), .B0(net112571), .B1(n3183), .Y(
        n7648) );
  OA22XL U8116 ( .A0(net112241), .A1(n1571), .B0(net112159), .B1(n3184), .Y(
        n7646) );
  OA22XL U8117 ( .A0(net112231), .A1(n1572), .B0(net112159), .B1(n3185), .Y(
        n7820) );
  OA22X1 U8118 ( .A0(net112487), .A1(n1380), .B0(net112363), .B1(n2993), .Y(
        n8679) );
  OA22XL U8119 ( .A0(net112231), .A1(n1573), .B0(net112153), .B1(n3186), .Y(
        n7812) );
  OA22X1 U8120 ( .A0(net112471), .A1(n1381), .B0(net112347), .B1(n2994), .Y(
        n7639) );
  OA22XL U8121 ( .A0(net112241), .A1(n1574), .B0(net112159), .B1(n3187), .Y(
        n7638) );
  OA22X1 U8122 ( .A0(net112487), .A1(n2824), .B0(net112355), .B1(n832), .Y(
        n8116) );
  OA22X1 U8123 ( .A0(net112233), .A1(n2825), .B0(net112151), .B1(n833), .Y(
        n8115) );
  OA22X1 U8124 ( .A0(net112067), .A1(n2826), .B0(net111943), .B1(n834), .Y(
        n8114) );
  OA22X1 U8125 ( .A0(net112485), .A1(n1382), .B0(net112361), .B1(n2995), .Y(
        n8588) );
  OA22X1 U8126 ( .A0(net112665), .A1(n1383), .B0(net112565), .B1(n2996), .Y(
        n8589) );
  OA22X1 U8127 ( .A0(net112489), .A1(n1384), .B0(net112331), .B1(n2997), .Y(
        n8776) );
  OA22X1 U8128 ( .A0(net112665), .A1(n1385), .B0(net112565), .B1(n2998), .Y(
        n8777) );
  OA22X1 U8129 ( .A0(net112457), .A1(n1386), .B0(net112333), .B1(n2999), .Y(
        n6712) );
  OA22X1 U8130 ( .A0(net112233), .A1(n2827), .B0(net112165), .B1(n835), .Y(
        n6711) );
  OA22X1 U8131 ( .A0(net112679), .A1(n1387), .B0(net112577), .B1(n3000), .Y(
        n6713) );
  OA22X1 U8132 ( .A0(net112487), .A1(n2828), .B0(net112355), .B1(n836), .Y(
        n8108) );
  OA22X1 U8133 ( .A0(net112067), .A1(n2829), .B0(net111943), .B1(n837), .Y(
        n8106) );
  OA22X1 U8134 ( .A0(net112477), .A1(n1388), .B0(net112353), .B1(n3001), .Y(
        n8015) );
  OA22X1 U8135 ( .A0(net112233), .A1(n2830), .B0(net112151), .B1(n838), .Y(
        n8014) );
  OA22X1 U8136 ( .A0(net112665), .A1(n1389), .B0(net112563), .B1(n3002), .Y(
        n8016) );
  OA22XL U8137 ( .A0(net112231), .A1(n1575), .B0(net112153), .B1(n3188), .Y(
        n7917) );
  OA22X1 U8138 ( .A0(net112681), .A1(n1390), .B0(net112577), .B1(n3003), .Y(
        n6542) );
  OA22X1 U8139 ( .A0(net112457), .A1(n1391), .B0(net112333), .B1(n3004), .Y(
        n6541) );
  OA22X1 U8140 ( .A0(net112681), .A1(n1392), .B0(net112577), .B1(n3005), .Y(
        n6534) );
  OA22X1 U8141 ( .A0(net112455), .A1(n1393), .B0(net112331), .B1(n3006), .Y(
        n6533) );
  OA22X1 U8142 ( .A0(net112469), .A1(n1394), .B0(net112345), .B1(n3007), .Y(
        n7498) );
  OA22X1 U8143 ( .A0(net112057), .A1(n1395), .B0(net111933), .B1(n3008), .Y(
        n7496) );
  OA22X1 U8144 ( .A0(net112483), .A1(n1396), .B0(net112359), .B1(n3009), .Y(
        n8482) );
  OA22X1 U8145 ( .A0(net112235), .A1(n1397), .B0(net112153), .B1(n3010), .Y(
        n8481) );
  OA22X1 U8146 ( .A0(net112469), .A1(n1398), .B0(net112345), .B1(n3011), .Y(
        n7490) );
  OA22X1 U8147 ( .A0(net112057), .A1(n1399), .B0(net111933), .B1(n3012), .Y(
        n7488) );
  OA22X1 U8148 ( .A0(net112471), .A1(n1400), .B0(net112347), .B1(n3013), .Y(
        net105009) );
  OA22XL U8149 ( .A0(net112241), .A1(n1576), .B0(net112159), .B1(n3189), .Y(
        net105010) );
  OA22X1 U8150 ( .A0(net112059), .A1(n1401), .B0(net111935), .B1(n3014), .Y(
        net105011) );
  OA22X1 U8151 ( .A0(net112455), .A1(n1402), .B0(net112331), .B1(n3015), .Y(
        n6391) );
  OA22X1 U8152 ( .A0(net112043), .A1(n1403), .B0(net111919), .B1(n3016), .Y(
        n6389) );
  OA22X1 U8153 ( .A0(net112461), .A1(n1404), .B0(net112337), .B1(n3017), .Y(
        n6966) );
  OA22X1 U8154 ( .A0(net112235), .A1(n1405), .B0(net112165), .B1(n3018), .Y(
        n6965) );
  OA22X1 U8155 ( .A0(net112049), .A1(n1406), .B0(net111925), .B1(n3019), .Y(
        n6964) );
  OA22X1 U8156 ( .A0(net112455), .A1(n1407), .B0(net112331), .B1(n3020), .Y(
        n6383) );
  OA22X1 U8157 ( .A0(net112681), .A1(n1408), .B0(net112565), .B1(n3021), .Y(
        n6384) );
  OA22X1 U8158 ( .A0(net112459), .A1(n1409), .B0(net112335), .B1(n3022), .Y(
        n6874) );
  OA22X1 U8159 ( .A0(net112047), .A1(n1410), .B0(net111923), .B1(n3023), .Y(
        n6872) );
  OA22X1 U8160 ( .A0(net112453), .A1(n1411), .B0(net112329), .B1(n3024), .Y(
        n6275) );
  OA22X1 U8161 ( .A0(net112459), .A1(n1412), .B0(net112335), .B1(n3025), .Y(
        n6791) );
  OA22X1 U8162 ( .A0(net112235), .A1(n1413), .B0(net112165), .B1(n3026), .Y(
        n6790) );
  OA22X1 U8163 ( .A0(net112047), .A1(n1414), .B0(net111923), .B1(n3027), .Y(
        n6789) );
  OA22X1 U8164 ( .A0(net112463), .A1(n1415), .B0(net112339), .B1(n3028), .Y(
        n7057) );
  OA22X1 U8165 ( .A0(net112051), .A1(n1416), .B0(net111927), .B1(n3029), .Y(
        n7055) );
  OA22X1 U8166 ( .A0(net112473), .A1(n2831), .B0(net112349), .B1(n839), .Y(
        n7724) );
  OA22XL U8167 ( .A0(net112241), .A1(n1577), .B0(net112159), .B1(n3190), .Y(
        n7723) );
  OA22X1 U8168 ( .A0(net112061), .A1(n2832), .B0(net111937), .B1(n840), .Y(
        n7722) );
  OA22X1 U8169 ( .A0(net112489), .A1(n1417), .B0(net112331), .B1(n3030), .Y(
        n8857) );
  OA22X1 U8170 ( .A0(net112481), .A1(n1418), .B0(net112357), .B1(n3031), .Y(
        n8298) );
  OA22X1 U8171 ( .A0(net112235), .A1(n1419), .B0(net112153), .B1(n3032), .Y(
        n8297) );
  OA22X1 U8172 ( .A0(net112671), .A1(n1420), .B0(net112569), .B1(n3033), .Y(
        n9098) );
  OA22X1 U8173 ( .A0(net112239), .A1(n1422), .B0(net112159), .B1(n3035), .Y(
        n9096) );
  OA22X1 U8174 ( .A0(net112477), .A1(n1423), .B0(net112353), .B1(n3036), .Y(
        n8023) );
  OA22X1 U8175 ( .A0(net112671), .A1(n1424), .B0(net112569), .B1(n3037), .Y(
        n8862) );
  OA22X1 U8176 ( .A0(net112489), .A1(n1425), .B0(net112303), .B1(n3038), .Y(
        n8861) );
  OA22X1 U8177 ( .A0(net112239), .A1(n1426), .B0(net112159), .B1(n3039), .Y(
        n8860) );
  NAND4BX1 U8178 ( .AN(n7598), .B(n7597), .C(n7596), .D(n7595), .Y(n7609) );
  NAND4BX1 U8179 ( .AN(n7834), .B(n7833), .C(n7832), .D(n7831), .Y(n7845) );
  CLKMX2X2 U8180 ( .A(n7542), .B(n7541), .S0(net108963), .Y(net105003) );
  CLKMX2X2 U8181 ( .A(n6843), .B(n6842), .S0(net108963), .Y(net106270) );
  CLKMX2X2 U8182 ( .A(n6345), .B(n6344), .S0(net108963), .Y(net107041) );
  OA22X1 U8183 ( .A0(net112481), .A1(n1427), .B0(net112357), .B1(n3040), .Y(
        n8302) );
  NAND2X1 U8184 ( .A(n4802), .B(\i_MIPS/n340 ), .Y(n7476) );
  NAND2X1 U8185 ( .A(n4684), .B(n3787), .Y(n8911) );
  NAND4X1 U8186 ( .A(n9371), .B(n9370), .C(n9369), .D(n9368), .Y(n11339) );
  OA22X2 U8187 ( .A0(n5165), .A1(n911), .B0(n5121), .B1(n2428), .Y(n9371) );
  OA22X2 U8188 ( .A0(n5251), .A1(n912), .B0(n5205), .B1(n2429), .Y(n9370) );
  OA22X2 U8189 ( .A0(n5442), .A1(n440), .B0(n5392), .B1(n2002), .Y(n9646) );
  NAND4X1 U8190 ( .A(n9953), .B(n9952), .C(n9951), .D(n9950), .Y(n11337) );
  OA22X1 U8191 ( .A0(n5441), .A1(n999), .B0(n5395), .B1(n2571), .Y(n9950) );
  OA22X1 U8192 ( .A0(n5178), .A1(n1000), .B0(n5134), .B1(n2572), .Y(n9953) );
  OA22X1 U8193 ( .A0(n5264), .A1(n1001), .B0(n5219), .B1(n2573), .Y(n9952) );
  OA22X2 U8194 ( .A0(n5445), .A1(n2420), .B0(n5389), .B1(n443), .Y(n9538) );
  OA22X2 U8195 ( .A0(n5435), .A1(n915), .B0(n5390), .B1(n2432), .Y(n9670) );
  OA22X2 U8196 ( .A0(n5258), .A1(n916), .B0(n5212), .B1(n2433), .Y(n9672) );
  OA22X2 U8197 ( .A0(n5433), .A1(n441), .B0(n5399), .B1(n2003), .Y(n9469) );
  NAND4X1 U8198 ( .A(n9658), .B(n9657), .C(n9656), .D(n9655), .Y(n11336) );
  OA22X1 U8199 ( .A0(n5442), .A1(n1002), .B0(n5402), .B1(n2574), .Y(n9655) );
  OA22X2 U8200 ( .A0(n5171), .A1(n918), .B0(n5138), .B1(n2435), .Y(n9658) );
  OA22X2 U8201 ( .A0(n5257), .A1(n919), .B0(n5211), .B1(n2436), .Y(n9657) );
  NAND4X1 U8202 ( .A(n10234), .B(n10233), .C(n10232), .D(n10231), .Y(n11259)
         );
  OA22X1 U8203 ( .A0(n5183), .A1(n1003), .B0(n5139), .B1(n2575), .Y(n10234) );
  OA22X1 U8204 ( .A0(n5268), .A1(n1004), .B0(n5223), .B1(n2576), .Y(n10233) );
  OA22X1 U8205 ( .A0(n5445), .A1(n1005), .B0(n5399), .B1(n2577), .Y(n10231) );
  NAND4X1 U8206 ( .A(n10226), .B(n10225), .C(n10224), .D(n10223), .Y(n11355)
         );
  NAND4X1 U8207 ( .A(n10238), .B(n10237), .C(n10236), .D(n10235), .Y(n11291)
         );
  OA22X1 U8208 ( .A0(n5165), .A1(n1006), .B0(n5138), .B1(n2578), .Y(n10238) );
  OA22X1 U8209 ( .A0(n5269), .A1(n1007), .B0(n5218), .B1(n2579), .Y(n10237) );
  OA22X1 U8210 ( .A0(n5446), .A1(n1008), .B0(n5400), .B1(n2580), .Y(n10235) );
  NAND4X1 U8211 ( .A(n10230), .B(n10229), .C(n10228), .D(n10227), .Y(n11323)
         );
  NAND4X1 U8212 ( .A(n9751), .B(n9750), .C(n9749), .D(n9748), .Y(n11261) );
  NAND4X1 U8213 ( .A(n9743), .B(n9742), .C(n9741), .D(n9740), .Y(n11357) );
  OA22X1 U8214 ( .A0(n5174), .A1(n1009), .B0(n5129), .B1(n2581), .Y(n9743) );
  OA22X1 U8215 ( .A0(n5260), .A1(n1010), .B0(n5214), .B1(n2582), .Y(n9742) );
  OA22X1 U8216 ( .A0(n5437), .A1(n1011), .B0(n5392), .B1(n2583), .Y(n9740) );
  NAND4X1 U8217 ( .A(n9755), .B(n9754), .C(n9753), .D(n9752), .Y(n11293) );
  NAND4X1 U8218 ( .A(n9747), .B(n9746), .C(n9745), .D(n9744), .Y(n11325) );
  NAND4X1 U8219 ( .A(n9695), .B(n9694), .C(n9693), .D(n9692), .Y(n11352) );
  OA22X1 U8220 ( .A0(n5172), .A1(n2509), .B0(n5127), .B1(n758), .Y(n9695) );
  OA22X1 U8221 ( .A0(n5258), .A1(n2510), .B0(n5212), .B1(n759), .Y(n9694) );
  OA22X1 U8222 ( .A0(n5435), .A1(n2511), .B0(n5390), .B1(n760), .Y(n9692) );
  NAND4X1 U8223 ( .A(n9705), .B(n9704), .C(n9703), .D(n9702), .Y(n11256) );
  OA22X1 U8224 ( .A0(n5173), .A1(n1012), .B0(n5128), .B1(n2584), .Y(n9705) );
  OA22X1 U8225 ( .A0(n5259), .A1(n1013), .B0(n5213), .B1(n2585), .Y(n9704) );
  OA22X1 U8226 ( .A0(n5436), .A1(n2512), .B0(n5391), .B1(n761), .Y(n9702) );
  NAND4X1 U8227 ( .A(n9710), .B(n9709), .C(n9708), .D(n9707), .Y(n11288) );
  OA22X1 U8228 ( .A0(n5173), .A1(n1014), .B0(n5128), .B1(n2586), .Y(n9710) );
  OA22X1 U8229 ( .A0(n5259), .A1(n2513), .B0(n5213), .B1(n762), .Y(n9709) );
  OA22X1 U8230 ( .A0(n5436), .A1(n2514), .B0(n5391), .B1(n763), .Y(n9707) );
  NAND4X1 U8231 ( .A(n9700), .B(n9699), .C(n9698), .D(n9697), .Y(n11320) );
  OA22X1 U8232 ( .A0(n5172), .A1(n1015), .B0(n5127), .B1(n2587), .Y(n9700) );
  OA22X1 U8233 ( .A0(n5258), .A1(n1016), .B0(n5212), .B1(n2588), .Y(n9699) );
  OA22X1 U8234 ( .A0(n5435), .A1(n2515), .B0(n5390), .B1(n764), .Y(n9697) );
  NAND4X1 U8235 ( .A(n9797), .B(n9796), .C(n9795), .D(n9794), .Y(n11260) );
  NAND4X1 U8236 ( .A(n9787), .B(n9786), .C(n9785), .D(n9784), .Y(n11356) );
  OA22X1 U8237 ( .A0(n5175), .A1(n1017), .B0(n5130), .B1(n2589), .Y(n9787) );
  OA22X1 U8238 ( .A0(n5261), .A1(n1018), .B0(n5215), .B1(n2590), .Y(n9786) );
  OA22X1 U8239 ( .A0(n5438), .A1(n1019), .B0(n5403), .B1(n2591), .Y(n9784) );
  NAND4X1 U8240 ( .A(n9802), .B(n9801), .C(n9800), .D(n9799), .Y(n11292) );
  NAND4X1 U8241 ( .A(n9792), .B(n9791), .C(n9790), .D(n9789), .Y(n11324) );
  NAND4X1 U8242 ( .A(n9773), .B(n9772), .C(n9771), .D(n9770), .Y(n11258) );
  NAND4X1 U8243 ( .A(n9763), .B(n9762), .C(n9761), .D(n9760), .Y(n11354) );
  NAND4X1 U8244 ( .A(n9778), .B(n9777), .C(n9776), .D(n9775), .Y(n11290) );
  NAND4X1 U8245 ( .A(n9768), .B(n9767), .C(n9766), .D(n9765), .Y(n11322) );
  NAND4X1 U8246 ( .A(n9729), .B(n9728), .C(n9727), .D(n9726), .Y(n11257) );
  NAND4X1 U8247 ( .A(n9719), .B(n9718), .C(n9717), .D(n9716), .Y(n11353) );
  NAND4X1 U8248 ( .A(n9734), .B(n9733), .C(n9732), .D(n9731), .Y(n11289) );
  NAND4X1 U8249 ( .A(n9724), .B(n9723), .C(n9722), .D(n9721), .Y(n11321) );
  NAND4X1 U8250 ( .A(n10108), .B(n10107), .C(n10106), .D(n10105), .Y(n11351)
         );
  NAND4X1 U8251 ( .A(n10118), .B(n10117), .C(n10116), .D(n10115), .Y(n11255)
         );
  NAND4X1 U8252 ( .A(n10123), .B(n10122), .C(n10121), .D(n10120), .Y(n11287)
         );
  NAND4X1 U8253 ( .A(n10113), .B(n10112), .C(n10111), .D(n10110), .Y(n11319)
         );
  NAND4X1 U8254 ( .A(n9886), .B(n9885), .C(n9884), .D(n9883), .Y(n11350) );
  OA22X1 U8255 ( .A0(n5180), .A1(n1638), .B0(n5133), .B1(n3322), .Y(n9886) );
  OA22X1 U8256 ( .A0(n5266), .A1(n1639), .B0(n5218), .B1(n3323), .Y(n9885) );
  OA22X1 U8257 ( .A0(n5440), .A1(n1640), .B0(n5394), .B1(n3324), .Y(n9883) );
  NAND4X1 U8258 ( .A(n9896), .B(n9895), .C(n9894), .D(n9893), .Y(n11254) );
  OA22X1 U8259 ( .A0(n5180), .A1(n1641), .B0(n5133), .B1(n3325), .Y(n9896) );
  OA22X1 U8260 ( .A0(n5266), .A1(n1642), .B0(n5218), .B1(n3326), .Y(n9895) );
  OA22X1 U8261 ( .A0(n5440), .A1(n1643), .B0(n5394), .B1(n3327), .Y(n9893) );
  NAND4X1 U8262 ( .A(n9901), .B(n9900), .C(n9899), .D(n9898), .Y(n11286) );
  OA22X1 U8263 ( .A0(n5180), .A1(n1644), .B0(n5133), .B1(n3328), .Y(n9901) );
  OA22X1 U8264 ( .A0(n5266), .A1(n1645), .B0(n5218), .B1(n3329), .Y(n9900) );
  OA22X1 U8265 ( .A0(n5440), .A1(n1646), .B0(n5394), .B1(n3330), .Y(n9898) );
  NAND4X1 U8266 ( .A(n9891), .B(n9890), .C(n9889), .D(n9888), .Y(n11318) );
  OA22X1 U8267 ( .A0(n5180), .A1(n1647), .B0(n5133), .B1(n3331), .Y(n9891) );
  OA22X1 U8268 ( .A0(n5266), .A1(n1648), .B0(n5218), .B1(n3332), .Y(n9890) );
  OA22X1 U8269 ( .A0(n5440), .A1(n1649), .B0(n5394), .B1(n3333), .Y(n9888) );
  NAND4X1 U8270 ( .A(n9910), .B(n9909), .C(n9908), .D(n9907), .Y(n11349) );
  OA22X1 U8271 ( .A0(n5180), .A1(n1650), .B0(n5133), .B1(n3334), .Y(n9910) );
  OA22X1 U8272 ( .A0(n5266), .A1(n1651), .B0(n5218), .B1(n3335), .Y(n9909) );
  OA22X1 U8273 ( .A0(n5440), .A1(n1652), .B0(n5394), .B1(n3336), .Y(n9907) );
  NAND4X1 U8274 ( .A(n9920), .B(n9919), .C(n9918), .D(n9917), .Y(n11253) );
  NAND4X1 U8275 ( .A(n9925), .B(n9924), .C(n9923), .D(n9922), .Y(n11285) );
  NAND4X1 U8276 ( .A(n9915), .B(n9914), .C(n9913), .D(n9912), .Y(n11317) );
  OA22X1 U8277 ( .A0(n5180), .A1(n1653), .B0(n5133), .B1(n3337), .Y(n9915) );
  OA22X1 U8278 ( .A0(n5266), .A1(n1654), .B0(n5218), .B1(n3338), .Y(n9914) );
  OA22X1 U8279 ( .A0(n5440), .A1(n1655), .B0(n5394), .B1(n3339), .Y(n9912) );
  NAND4X1 U8280 ( .A(n9842), .B(n9841), .C(n9840), .D(n9839), .Y(n11348) );
  NAND4X1 U8281 ( .A(n9852), .B(n9851), .C(n9850), .D(n9849), .Y(n11252) );
  OA22X1 U8282 ( .A0(n5177), .A1(n1656), .B0(n5132), .B1(n3340), .Y(n9852) );
  OA22X1 U8283 ( .A0(n5263), .A1(n1657), .B0(n5217), .B1(n3341), .Y(n9851) );
  OA22X1 U8284 ( .A0(n5439), .A1(n1658), .B0(n5393), .B1(n3342), .Y(n9849) );
  NAND4X1 U8285 ( .A(n9857), .B(n9856), .C(n9855), .D(n9854), .Y(n11284) );
  OA22X1 U8286 ( .A0(n5177), .A1(n1659), .B0(n5132), .B1(n3343), .Y(n9857) );
  OA22X1 U8287 ( .A0(n5263), .A1(n1660), .B0(n5217), .B1(n3344), .Y(n9856) );
  OA22X1 U8288 ( .A0(n5439), .A1(n1661), .B0(n5393), .B1(n3345), .Y(n9854) );
  NAND4X1 U8289 ( .A(n9847), .B(n9846), .C(n9845), .D(n9844), .Y(n11316) );
  NAND4X1 U8290 ( .A(n9862), .B(n9861), .C(n9860), .D(n9859), .Y(n11347) );
  OA22X1 U8291 ( .A0(n5177), .A1(n1662), .B0(n5132), .B1(n3346), .Y(n9862) );
  OA22X1 U8292 ( .A0(n5263), .A1(n1663), .B0(n5217), .B1(n3347), .Y(n9861) );
  OA22X1 U8293 ( .A0(n5439), .A1(n1664), .B0(n5393), .B1(n3348), .Y(n9859) );
  NAND4X1 U8294 ( .A(n9872), .B(n9871), .C(n9870), .D(n9869), .Y(n11251) );
  OA22X1 U8295 ( .A0(n5177), .A1(n1665), .B0(n5132), .B1(n3349), .Y(n9872) );
  OA22X1 U8296 ( .A0(n5263), .A1(n1666), .B0(n5217), .B1(n3350), .Y(n9871) );
  OA22X1 U8297 ( .A0(n5439), .A1(n1667), .B0(n5393), .B1(n3351), .Y(n9869) );
  NAND4X1 U8298 ( .A(n9877), .B(n9876), .C(n9875), .D(n9874), .Y(n11283) );
  OA22X1 U8299 ( .A0(n5177), .A1(n1668), .B0(n5132), .B1(n3352), .Y(n9877) );
  OA22X1 U8300 ( .A0(n5263), .A1(n1669), .B0(n5217), .B1(n3353), .Y(n9876) );
  OA22X1 U8301 ( .A0(n5439), .A1(n1670), .B0(n5393), .B1(n3354), .Y(n9874) );
  NAND4X1 U8302 ( .A(n9867), .B(n9866), .C(n9865), .D(n9864), .Y(n11315) );
  OA22X1 U8303 ( .A0(n5177), .A1(n1671), .B0(n5132), .B1(n3355), .Y(n9867) );
  OA22X1 U8304 ( .A0(n5263), .A1(n1672), .B0(n5217), .B1(n3356), .Y(n9866) );
  OA22X1 U8305 ( .A0(n5439), .A1(n1673), .B0(n5393), .B1(n3357), .Y(n9864) );
  NAND4X1 U8306 ( .A(n10006), .B(n10005), .C(n10004), .D(n10003), .Y(n11346)
         );
  OA22X1 U8307 ( .A0(n5180), .A1(n1674), .B0(n5133), .B1(n3358), .Y(n10006) );
  OA22X1 U8308 ( .A0(n5266), .A1(n1675), .B0(n5218), .B1(n3359), .Y(n10005) );
  OA22X1 U8309 ( .A0(n5440), .A1(n1676), .B0(n5397), .B1(n3360), .Y(n10003) );
  NAND4X1 U8310 ( .A(n10016), .B(n10015), .C(n10014), .D(n10013), .Y(n11250)
         );
  OA22X1 U8311 ( .A0(n5180), .A1(n1677), .B0(n5133), .B1(n3361), .Y(n10016) );
  OA22X1 U8312 ( .A0(n5266), .A1(n1678), .B0(n5218), .B1(n3362), .Y(n10015) );
  OA22X1 U8313 ( .A0(n5440), .A1(n1679), .B0(n5397), .B1(n3363), .Y(n10013) );
  NAND4X1 U8314 ( .A(n10021), .B(n10020), .C(n10019), .D(n10018), .Y(n11282)
         );
  OA22X1 U8315 ( .A0(n5180), .A1(n1680), .B0(n5133), .B1(n3364), .Y(n10021) );
  OA22X1 U8316 ( .A0(n5266), .A1(n1681), .B0(n5218), .B1(n3365), .Y(n10020) );
  OA22X1 U8317 ( .A0(n5440), .A1(n1682), .B0(n5397), .B1(n3366), .Y(n10018) );
  NAND4X1 U8318 ( .A(n10011), .B(n10010), .C(n10009), .D(n10008), .Y(n11314)
         );
  OA22X1 U8319 ( .A0(n5180), .A1(n1683), .B0(n5133), .B1(n3367), .Y(n10011) );
  OA22X1 U8320 ( .A0(n5266), .A1(n1684), .B0(n5218), .B1(n3368), .Y(n10010) );
  OA22X1 U8321 ( .A0(n5440), .A1(n1685), .B0(n5397), .B1(n3369), .Y(n10008) );
  NAND4X1 U8322 ( .A(n9977), .B(n9976), .C(n9975), .D(n9974), .Y(n11345) );
  NAND4X1 U8323 ( .A(n9987), .B(n9986), .C(n9985), .D(n9984), .Y(n11249) );
  NAND4X1 U8324 ( .A(n9992), .B(n9991), .C(n9990), .D(n9989), .Y(n11281) );
  OA22X1 U8325 ( .A0(n5180), .A1(n1686), .B0(n5133), .B1(n3370), .Y(n9992) );
  OA22X1 U8326 ( .A0(n5266), .A1(n1687), .B0(n5218), .B1(n3371), .Y(n9991) );
  OA22X1 U8327 ( .A0(n5440), .A1(n1688), .B0(n5397), .B1(n3372), .Y(n9989) );
  NAND4X1 U8328 ( .A(n9982), .B(n9981), .C(n9980), .D(n9979), .Y(n11313) );
  NAND4X1 U8329 ( .A(n10030), .B(n10029), .C(n10028), .D(n10027), .Y(n11344)
         );
  OA22X1 U8330 ( .A0(n5180), .A1(n1689), .B0(n5133), .B1(n3373), .Y(n10030) );
  OA22X1 U8331 ( .A0(n5266), .A1(n1690), .B0(n5218), .B1(n3374), .Y(n10029) );
  OA22X1 U8332 ( .A0(n5440), .A1(n1691), .B0(n5397), .B1(n3375), .Y(n10027) );
  NAND4X1 U8333 ( .A(n10040), .B(n10039), .C(n10038), .D(n10037), .Y(n11248)
         );
  OA22X1 U8334 ( .A0(n5181), .A1(n1692), .B0(n5136), .B1(n3376), .Y(n10040) );
  OA22X1 U8335 ( .A0(n5263), .A1(n1693), .B0(n5221), .B1(n3377), .Y(n10039) );
  OA22X1 U8336 ( .A0(n5443), .A1(n1694), .B0(n5394), .B1(n3378), .Y(n10037) );
  NAND4X1 U8337 ( .A(n10045), .B(n10044), .C(n10043), .D(n10042), .Y(n11280)
         );
  OA22X1 U8338 ( .A0(n5181), .A1(n1695), .B0(n5136), .B1(n3379), .Y(n10045) );
  OA22X1 U8339 ( .A0(n5263), .A1(n1696), .B0(n5221), .B1(n3380), .Y(n10044) );
  OA22X1 U8340 ( .A0(n5443), .A1(n1697), .B0(n5394), .B1(n3381), .Y(n10042) );
  NAND4X1 U8341 ( .A(n10035), .B(n10034), .C(n10033), .D(n10032), .Y(n11312)
         );
  OA22X1 U8342 ( .A0(n5181), .A1(n1698), .B0(n5136), .B1(n3382), .Y(n10035) );
  OA22X1 U8343 ( .A0(n5263), .A1(n1699), .B0(n5221), .B1(n3383), .Y(n10034) );
  OA22X1 U8344 ( .A0(n5443), .A1(n1700), .B0(n5394), .B1(n3384), .Y(n10032) );
  NAND4X1 U8345 ( .A(n11123), .B(n11122), .C(n11121), .D(n11120), .Y(n11343)
         );
  NAND4X1 U8346 ( .A(n11133), .B(n11132), .C(n11131), .D(n11130), .Y(n11247)
         );
  NAND4X1 U8347 ( .A(n11144), .B(n11143), .C(n11142), .D(n11141), .Y(n11279)
         );
  NAND4X1 U8348 ( .A(n11128), .B(n11127), .C(n11126), .D(n11125), .Y(n11311)
         );
  NAND4X1 U8349 ( .A(n10059), .B(n10058), .C(n10057), .D(n10056), .Y(n11342)
         );
  OA22X1 U8350 ( .A0(n5181), .A1(n1701), .B0(n5136), .B1(n3385), .Y(n10059) );
  OA22X1 U8351 ( .A0(n5263), .A1(n1702), .B0(n5221), .B1(n3386), .Y(n10058) );
  OA22X1 U8352 ( .A0(n5443), .A1(n1703), .B0(n5397), .B1(n3387), .Y(n10056) );
  NAND4X1 U8353 ( .A(n10069), .B(n10068), .C(n10067), .D(n10066), .Y(n11246)
         );
  OA22X1 U8354 ( .A0(n5181), .A1(n1704), .B0(n5136), .B1(n3388), .Y(n10069) );
  OA22X1 U8355 ( .A0(n5263), .A1(n1705), .B0(n5221), .B1(n3389), .Y(n10068) );
  OA22X1 U8356 ( .A0(n5443), .A1(n1706), .B0(n5397), .B1(n3390), .Y(n10066) );
  NAND4X1 U8357 ( .A(n10074), .B(n10073), .C(n10072), .D(n10071), .Y(n11278)
         );
  NAND4X1 U8358 ( .A(n10064), .B(n10063), .C(n10062), .D(n10061), .Y(n11310)
         );
  OA22X1 U8359 ( .A0(n5181), .A1(n1707), .B0(n5136), .B1(n3391), .Y(n10064) );
  OA22X1 U8360 ( .A0(n5263), .A1(n1708), .B0(n5221), .B1(n3392), .Y(n10063) );
  OA22X1 U8361 ( .A0(n5443), .A1(n1709), .B0(n5394), .B1(n3393), .Y(n10061) );
  NAND4X1 U8362 ( .A(n9401), .B(n9400), .C(n9399), .D(n9398), .Y(n11244) );
  OA22X1 U8363 ( .A0(n5166), .A1(n1020), .B0(n5122), .B1(n2592), .Y(n9401) );
  OA22X1 U8364 ( .A0(n5252), .A1(n1021), .B0(n5206), .B1(n2593), .Y(n9400) );
  OA22X1 U8365 ( .A0(n5431), .A1(n1022), .B0(n5387), .B1(n2594), .Y(n9398) );
  NAND4X1 U8366 ( .A(n9391), .B(n9390), .C(n9389), .D(n9388), .Y(n11340) );
  OA22X1 U8367 ( .A0(n5165), .A1(n1023), .B0(n5121), .B1(n2595), .Y(n9391) );
  OA22X1 U8368 ( .A0(n5251), .A1(n1024), .B0(n5205), .B1(n2596), .Y(n9390) );
  OA22X1 U8369 ( .A0(n5430), .A1(n1025), .B0(n5386), .B1(n2597), .Y(n9388) );
  NAND4X1 U8370 ( .A(n9406), .B(n9405), .C(n9404), .D(n9403), .Y(n11276) );
  OA22X1 U8371 ( .A0(n5166), .A1(n1026), .B0(n5122), .B1(n2598), .Y(n9406) );
  OA22X1 U8372 ( .A0(n5252), .A1(n1027), .B0(n5206), .B1(n2599), .Y(n9405) );
  OA22X1 U8373 ( .A0(n5431), .A1(n1028), .B0(n5387), .B1(n2600), .Y(n9403) );
  NAND4X1 U8374 ( .A(n9396), .B(n9395), .C(n9394), .D(n9393), .Y(n11308) );
  OA22X1 U8375 ( .A0(n5165), .A1(n1029), .B0(n5121), .B1(n2601), .Y(n9396) );
  OA22X1 U8376 ( .A0(n5251), .A1(n1030), .B0(n5205), .B1(n2602), .Y(n9395) );
  OA22X1 U8377 ( .A0(n5430), .A1(n1031), .B0(n5386), .B1(n2603), .Y(n9393) );
  NAND4X1 U8378 ( .A(n10094), .B(n10093), .C(n10092), .D(n10091), .Y(n11242)
         );
  OA22X1 U8379 ( .A0(n5182), .A1(n1032), .B0(n5137), .B1(n2604), .Y(n10094) );
  OA22X1 U8380 ( .A0(n5267), .A1(n1033), .B0(n5222), .B1(n2605), .Y(n10093) );
  NAND4X1 U8381 ( .A(n10084), .B(n10083), .C(n10082), .D(n10081), .Y(n11338)
         );
  OA22X1 U8382 ( .A0(n5182), .A1(n1034), .B0(n5137), .B1(n2606), .Y(n10084) );
  OA22X1 U8383 ( .A0(n5267), .A1(n1035), .B0(n5222), .B1(n2607), .Y(n10083) );
  OA22X1 U8384 ( .A0(n5444), .A1(n1036), .B0(n5398), .B1(n2608), .Y(n10081) );
  OA22X1 U8385 ( .A0(n5182), .A1(n1037), .B0(n5137), .B1(n2609), .Y(n10099) );
  OA22X1 U8386 ( .A0(n5267), .A1(n1038), .B0(n5222), .B1(n2610), .Y(n10098) );
  OA22X1 U8387 ( .A0(n5182), .A1(n1039), .B0(n5137), .B1(n2611), .Y(n10089) );
  OA22X1 U8388 ( .A0(n5267), .A1(n1040), .B0(n5222), .B1(n2612), .Y(n10088) );
  OA22X1 U8389 ( .A0(n5444), .A1(n1041), .B0(n5398), .B1(n2613), .Y(n10086) );
  OAI222XL U8390 ( .A0(n5097), .A1(n188), .B0(n5032), .B1(n5096), .C0(n5523), 
        .C1(\i_MIPS/n207 ), .Y(n11553) );
  OAI222XL U8391 ( .A0(n5097), .A1(n292), .B0(n5017), .B1(n5095), .C0(n5523), 
        .C1(\i_MIPS/n206 ), .Y(n11554) );
  OAI222XL U8392 ( .A0(n5097), .A1(n193), .B0(n1851), .B1(n5096), .C0(n5523), 
        .C1(\i_MIPS/n202 ), .Y(n11558) );
  OAI222XL U8393 ( .A0(n5097), .A1(n291), .B0(n5041), .B1(n5096), .C0(n5523), 
        .C1(\i_MIPS/n201 ), .Y(n11559) );
  OAI222XL U8394 ( .A0(n5098), .A1(n244), .B0(n1995), .B1(n5095), .C0(n5523), 
        .C1(\i_MIPS/n200 ), .Y(n11560) );
  OAI222XL U8395 ( .A0(n5098), .A1(n230), .B0(n5008), .B1(n5095), .C0(n5524), 
        .C1(\i_MIPS/n184 ), .Y(n11576) );
  OAI222XL U8396 ( .A0(n5097), .A1(n190), .B0(n5501), .B1(n5096), .C0(n5522), 
        .C1(\i_MIPS/n211 ), .Y(n11549) );
  OAI222XL U8397 ( .A0(n5097), .A1(n228), .B0(n1834), .B1(n5096), .C0(n5522), 
        .C1(\i_MIPS/n210 ), .Y(n11550) );
  OAI222XL U8398 ( .A0(n5097), .A1(n231), .B0(n1858), .B1(n5096), .C0(n5523), 
        .C1(\i_MIPS/n209 ), .Y(n11551) );
  OAI222XL U8399 ( .A0(n5097), .A1(n240), .B0(n1855), .B1(n5095), .C0(n5523), 
        .C1(\i_MIPS/n205 ), .Y(n11555) );
  OAI222XL U8400 ( .A0(n5097), .A1(n242), .B0(n1836), .B1(n5096), .C0(n5523), 
        .C1(\i_MIPS/n204 ), .Y(n11556) );
  OAI222XL U8401 ( .A0(n5097), .A1(n241), .B0(n1835), .B1(n5096), .C0(n5523), 
        .C1(\i_MIPS/n203 ), .Y(n11557) );
  OAI222XL U8402 ( .A0(n5098), .A1(n184), .B0(n1837), .B1(n5095), .C0(n5523), 
        .C1(\i_MIPS/n199 ), .Y(n11561) );
  OAI222XL U8403 ( .A0(n5097), .A1(n192), .B0(n5059), .B1(n5096), .C0(n5522), 
        .C1(\i_MIPS/n198 ), .Y(n11562) );
  OAI222XL U8404 ( .A0(n5098), .A1(n189), .B0(n1852), .B1(n5096), .C0(n5522), 
        .C1(\i_MIPS/n197 ), .Y(n11563) );
  OAI222XL U8405 ( .A0(n5098), .A1(n194), .B0(n5029), .B1(n5095), .C0(n5523), 
        .C1(\i_MIPS/n196 ), .Y(n11564) );
  OAI222XL U8406 ( .A0(n5098), .A1(n239), .B0(n1853), .B1(n5095), .C0(n5523), 
        .C1(\i_MIPS/n195 ), .Y(n11565) );
  OAI222XL U8407 ( .A0(n5098), .A1(n232), .B0(n1856), .B1(n5095), .C0(n5523), 
        .C1(\i_MIPS/n194 ), .Y(n11566) );
  OAI222XL U8408 ( .A0(n5097), .A1(n227), .B0(n1849), .B1(n5096), .C0(n5522), 
        .C1(\i_MIPS/n193 ), .Y(n11567) );
  OAI222XL U8409 ( .A0(n5097), .A1(n237), .B0(n1857), .B1(n5095), .C0(n5522), 
        .C1(\i_MIPS/n192 ), .Y(n11568) );
  OAI222XL U8410 ( .A0(n5097), .A1(n233), .B0(n4573), .B1(n5096), .C0(n5522), 
        .C1(\i_MIPS/n191 ), .Y(n11569) );
  OAI222XL U8411 ( .A0(n10836), .A1(n187), .B0(n5053), .B1(n5096), .C0(n5522), 
        .C1(\i_MIPS/n190 ), .Y(n11570) );
  OAI222XL U8412 ( .A0(n5097), .A1(n225), .B0(n1843), .B1(n5095), .C0(n5522), 
        .C1(\i_MIPS/n189 ), .Y(n11571) );
  OAI222XL U8413 ( .A0(n5097), .A1(n226), .B0(n1838), .B1(n10835), .C0(n5522), 
        .C1(\i_MIPS/n188 ), .Y(n11572) );
  OAI222XL U8414 ( .A0(n5097), .A1(n238), .B0(n1839), .B1(n5096), .C0(n5522), 
        .C1(\i_MIPS/n187 ), .Y(n11573) );
  OAI222XL U8415 ( .A0(n5098), .A1(n191), .B0(n1840), .B1(n5095), .C0(n5523), 
        .C1(\i_MIPS/n186 ), .Y(n11574) );
  OAI222XL U8416 ( .A0(n5098), .A1(n195), .B0(n5076), .B1(n5095), .C0(n5524), 
        .C1(\i_MIPS/n185 ), .Y(n11575) );
  OAI222XL U8417 ( .A0(n5098), .A1(n243), .B0(n1842), .B1(n5095), .C0(n5524), 
        .C1(\i_MIPS/n183 ), .Y(n11577) );
  NOR4XL U8418 ( .A(n6650), .B(n3686), .C(n6629), .D(n6651), .Y(n6496) );
  OA22XL U8419 ( .A0(n8726), .A1(n9265), .B0(n7974), .B1(n8729), .Y(n6957) );
  OA22XL U8420 ( .A0(n8659), .A1(n6598), .B0(n9001), .B1(n7561), .Y(n6267) );
  AOI2BB1X1 U8421 ( .A0N(n8736), .A1N(n7366), .B0(n6264), .Y(n6265) );
  NAND4X1 U8422 ( .A(n9521), .B(n9520), .C(n9519), .D(n9518), .Y(n11297) );
  OA22X1 U8423 ( .A0(n5434), .A1(n2516), .B0(n5395), .B1(n765), .Y(n9518) );
  OA22X1 U8424 ( .A0(n5169), .A1(n2517), .B0(n5125), .B1(n766), .Y(n9521) );
  OA22X1 U8425 ( .A0(n5255), .A1(n2518), .B0(n5209), .B1(n767), .Y(n9520) );
  NAND4X1 U8426 ( .A(n9682), .B(n9681), .C(n9680), .D(n9679), .Y(n11262) );
  OA22X1 U8427 ( .A0(n5434), .A1(n2519), .B0(n5387), .B1(n768), .Y(n9503) );
  OA22X1 U8428 ( .A0(n5169), .A1(n1042), .B0(n5125), .B1(n2614), .Y(n9506) );
  OA22X1 U8429 ( .A0(n5255), .A1(n1043), .B0(n5209), .B1(n2615), .Y(n9505) );
  OA22X1 U8430 ( .A0(n5434), .A1(n740), .B0(n5387), .B1(n2321), .Y(n9508) );
  OA22X1 U8431 ( .A0(n5169), .A1(n741), .B0(n5125), .B1(n2322), .Y(n9511) );
  OA22X1 U8432 ( .A0(n5255), .A1(n742), .B0(n5209), .B1(n2323), .Y(n9510) );
  OA22X1 U8433 ( .A0(n5434), .A1(n743), .B0(n5387), .B1(n2324), .Y(n9493) );
  OA22X1 U8434 ( .A0(n5169), .A1(n2520), .B0(n5125), .B1(n769), .Y(n9496) );
  OA22X1 U8435 ( .A0(n5255), .A1(n2521), .B0(n5209), .B1(n770), .Y(n9495) );
  OA22X1 U8436 ( .A0(n5434), .A1(n2522), .B0(n5387), .B1(n771), .Y(n9498) );
  OA22X1 U8437 ( .A0(n5169), .A1(n2523), .B0(n5125), .B1(n772), .Y(n9501) );
  OA22X1 U8438 ( .A0(n5255), .A1(n2524), .B0(n5209), .B1(n773), .Y(n9500) );
  NAND2XL U8439 ( .A(n6633), .B(n6638), .Y(n6254) );
  CLKINVX1 U8440 ( .A(n6609), .Y(n6365) );
  NOR4X1 U8441 ( .A(n9203), .B(n9202), .C(n9201), .D(n9200), .Y(n9204) );
  AO22X1 U8442 ( .A0(n4974), .A1(n190), .B0(n4967), .B1(n2180), .Y(n9203) );
  AO22X1 U8443 ( .A0(n9312), .A1(n657), .B0(n4987), .B1(n2181), .Y(n9201) );
  NOR4X1 U8444 ( .A(n9194), .B(n9193), .C(n9192), .D(n9191), .Y(n9195) );
  AO22X1 U8445 ( .A0(n4974), .A1(n658), .B0(n4967), .B1(n2182), .Y(n9194) );
  AO22X1 U8446 ( .A0(n9312), .A1(n659), .B0(n4987), .B1(n2183), .Y(n9192) );
  NOR4X1 U8447 ( .A(n9318), .B(n9317), .C(n9316), .D(n9315), .Y(n9319) );
  AO22X1 U8448 ( .A0(n4975), .A1(n228), .B0(n4968), .B1(n302), .Y(n9318) );
  AO22X1 U8449 ( .A0(n4980), .A1(n185), .B0(n4976), .B1(n201), .Y(n9317) );
  AO22X1 U8450 ( .A0(n9312), .A1(n197), .B0(n4988), .B1(n303), .Y(n9316) );
  NOR4X1 U8451 ( .A(n9301), .B(n9300), .C(n9299), .D(n9298), .Y(n9302) );
  AO22X1 U8452 ( .A0(n4975), .A1(n300), .B0(n4968), .B1(n1863), .Y(n9301) );
  AO22X1 U8453 ( .A0(n4980), .A1(n301), .B0(n4976), .B1(n1864), .Y(n9300) );
  AO22X1 U8454 ( .A0(n9312), .A1(n250), .B0(n4988), .B1(n1865), .Y(n9299) );
  NOR4X1 U8455 ( .A(n9217), .B(n9216), .C(n9215), .D(n9214), .Y(n9218) );
  AO22X1 U8456 ( .A0(n4879), .A1(n300), .B0(n4888), .B1(n1863), .Y(n9217) );
  AO22X1 U8457 ( .A0(n4863), .A1(n301), .B0(n4872), .B1(n1864), .Y(n9216) );
  AO22X1 U8458 ( .A0(n4845), .A1(n250), .B0(n4854), .B1(n1865), .Y(n9215) );
  NOR4X1 U8459 ( .A(n9230), .B(n9229), .C(n9228), .D(n9227), .Y(n9231) );
  AO22X1 U8460 ( .A0(n4880), .A1(n228), .B0(n4886), .B1(n302), .Y(n9230) );
  AO22X1 U8461 ( .A0(n4862), .A1(n185), .B0(n4870), .B1(n201), .Y(n9229) );
  AO22X1 U8462 ( .A0(n4845), .A1(n197), .B0(n4853), .B1(n303), .Y(n9228) );
  NOR4X1 U8463 ( .A(n7603), .B(n7602), .C(n7601), .D(n7600), .Y(n7604) );
  AO22X1 U8464 ( .A0(n4969), .A1(n183), .B0(n4966), .B1(n202), .Y(n7603) );
  AO22X1 U8465 ( .A0(n9312), .A1(n251), .B0(n4985), .B1(n304), .Y(n7601) );
  NOR4X1 U8466 ( .A(n7594), .B(n7593), .C(n7592), .D(n7591), .Y(n7595) );
  AO22X1 U8467 ( .A0(n4969), .A1(n198), .B0(n4966), .B1(n305), .Y(n7594) );
  AO22X1 U8468 ( .A0(n9312), .A1(n294), .B0(n4985), .B1(n1866), .Y(n7592) );
  NOR4X1 U8469 ( .A(n7536), .B(n7535), .C(n7534), .D(n7533), .Y(n7537) );
  AO22X1 U8470 ( .A0(n4969), .A1(n191), .B0(n4965), .B1(n724), .Y(n7536) );
  AO22X1 U8471 ( .A0(n9312), .A1(n660), .B0(n4985), .B1(n2184), .Y(n7534) );
  NOR4X1 U8472 ( .A(n7527), .B(n7526), .C(n7525), .D(n7524), .Y(n7528) );
  AO22X1 U8473 ( .A0(n4975), .A1(n220), .B0(n4966), .B1(n725), .Y(n7527) );
  AO22X1 U8474 ( .A0(n9312), .A1(n661), .B0(n4985), .B1(n2185), .Y(n7525) );
  NOR4X1 U8475 ( .A(n6837), .B(n6836), .C(n6835), .D(n6834), .Y(n6838) );
  AO22X1 U8476 ( .A0(n4971), .A1(n225), .B0(n4965), .B1(n2066), .Y(n6837) );
  AO22X1 U8477 ( .A0(n9312), .A1(n563), .B0(n4984), .B1(n2067), .Y(n6835) );
  NOR4X1 U8478 ( .A(n6828), .B(n6827), .C(n6826), .D(n6825), .Y(n6829) );
  AO22X1 U8479 ( .A0(n4971), .A1(n309), .B0(n4965), .B1(n2068), .Y(n6828) );
  AO22X1 U8480 ( .A0(n9312), .A1(n564), .B0(n4984), .B1(n2069), .Y(n6826) );
  NOR4X1 U8481 ( .A(n6187), .B(n6186), .C(n6185), .D(n6184), .Y(n6188) );
  AO22X1 U8482 ( .A0(n4971), .A1(n237), .B0(n4965), .B1(n2186), .Y(n6187) );
  NOR4X1 U8483 ( .A(n6178), .B(n6177), .C(n6176), .D(n6175), .Y(n6179) );
  AO22X1 U8484 ( .A0(n4971), .A1(n662), .B0(n4965), .B1(n2187), .Y(n6178) );
  AO22X1 U8485 ( .A0(n4992), .A1(n663), .B0(n4984), .B1(n2188), .Y(n6176) );
  NOR4X1 U8486 ( .A(n7444), .B(n7443), .C(n7442), .D(n7441), .Y(n7445) );
  AO22X1 U8487 ( .A0(n4972), .A1(n238), .B0(n4967), .B1(n2189), .Y(n7444) );
  NOR4X1 U8488 ( .A(n7435), .B(n7434), .C(n7433), .D(n7432), .Y(n7436) );
  AO22X1 U8489 ( .A0(n4972), .A1(n664), .B0(n4967), .B1(n2190), .Y(n7435) );
  NOR4X1 U8490 ( .A(n6757), .B(n6756), .C(n6755), .D(n6754), .Y(n6758) );
  AO22X1 U8491 ( .A0(n4971), .A1(n226), .B0(n4965), .B1(n2070), .Y(n6757) );
  AO22X1 U8492 ( .A0(n4989), .A1(n565), .B0(n4984), .B1(n2071), .Y(n6755) );
  NOR4X1 U8493 ( .A(n6748), .B(n6747), .C(n6746), .D(n6745), .Y(n6749) );
  AO22X1 U8494 ( .A0(n4971), .A1(n310), .B0(n4965), .B1(n2072), .Y(n6748) );
  AO22X1 U8495 ( .A0(n4989), .A1(n566), .B0(n4984), .B1(n2073), .Y(n6746) );
  NOR4X1 U8496 ( .A(n6920), .B(n6919), .C(n6918), .D(n6917), .Y(n6921) );
  NOR4X1 U8497 ( .A(n6911), .B(n6910), .C(n6909), .D(n6908), .Y(n6912) );
  NOR4X1 U8498 ( .A(n7012), .B(n7011), .C(n7010), .D(n7009), .Y(n7013) );
  AO22X1 U8499 ( .A0(n4972), .A1(n239), .B0(n4967), .B1(n2191), .Y(n7012) );
  NOR4X1 U8500 ( .A(n7003), .B(n7002), .C(n7001), .D(n7000), .Y(n7004) );
  AO22X1 U8501 ( .A0(n4972), .A1(n665), .B0(n4967), .B1(n2192), .Y(n7003) );
  NOR4X1 U8502 ( .A(n6339), .B(n6338), .C(n6337), .D(n6336), .Y(n6340) );
  AO22X1 U8503 ( .A0(n4971), .A1(n227), .B0(n4965), .B1(n2074), .Y(n6339) );
  AO22X1 U8504 ( .A0(n9312), .A1(n567), .B0(n4984), .B1(n2075), .Y(n6337) );
  NOR4X1 U8505 ( .A(n6330), .B(n6329), .C(n6328), .D(n6327), .Y(n6331) );
  AO22X1 U8506 ( .A0(n4971), .A1(n311), .B0(n4965), .B1(n2076), .Y(n6330) );
  AO22X1 U8507 ( .A0(n4992), .A1(n568), .B0(n4984), .B1(n2077), .Y(n6328) );
  NOR4X1 U8508 ( .A(n8133), .B(n8132), .C(n8131), .D(n8130), .Y(n8134) );
  AO22X1 U8509 ( .A0(n4973), .A1(n291), .B0(n4966), .B1(n2193), .Y(n8133) );
  NOR4X1 U8510 ( .A(n8124), .B(n8123), .C(n8122), .D(n8121), .Y(n8125) );
  AO22X1 U8511 ( .A0(n4973), .A1(n666), .B0(n4966), .B1(n2194), .Y(n8124) );
  NOR4X1 U8512 ( .A(n7943), .B(n7942), .C(n7941), .D(n7940), .Y(n7944) );
  AO22X1 U8513 ( .A0(n4973), .A1(n192), .B0(n4966), .B1(n726), .Y(n7943) );
  NOR4X1 U8514 ( .A(n7934), .B(n7933), .C(n7932), .D(n7931), .Y(n7935) );
  AO22X1 U8515 ( .A0(n4973), .A1(n214), .B0(n4966), .B1(n715), .Y(n7934) );
  NOR4X1 U8516 ( .A(n7262), .B(n7261), .C(n7260), .D(n7259), .Y(n7263) );
  NOR4X1 U8517 ( .A(n7253), .B(n7252), .C(n7251), .D(n7250), .Y(n7254) );
  NOR4X1 U8518 ( .A(n7769), .B(n7768), .C(n7767), .D(n7766), .Y(n7770) );
  AO22X1 U8519 ( .A0(n4880), .A1(n184), .B0(n4886), .B1(n203), .Y(n7769) );
  AO22X1 U8520 ( .A0(n4862), .A1(n295), .B0(n4871), .B1(n1867), .Y(n7768) );
  AO22X1 U8521 ( .A0(n4845), .A1(n289), .B0(n4853), .B1(n1859), .Y(n7767) );
  NOR4X1 U8522 ( .A(n7760), .B(n7759), .C(n7758), .D(n7757), .Y(n7761) );
  AO22X1 U8523 ( .A0(n4878), .A1(n199), .B0(n4887), .B1(n306), .Y(n7760) );
  AO22X1 U8524 ( .A0(n4861), .A1(n290), .B0(n4870), .B1(n1860), .Y(n7759) );
  AO22X1 U8525 ( .A0(n4847), .A1(n236), .B0(n4852), .B1(n1861), .Y(n7758) );
  NOR4X1 U8526 ( .A(n7677), .B(n7676), .C(n7675), .D(n7674), .Y(n7678) );
  NOR4X1 U8527 ( .A(n7664), .B(n7663), .C(n7662), .D(n7661), .Y(n7665) );
  AO22X1 U8528 ( .A0(n4880), .A1(n183), .B0(n4888), .B1(n202), .Y(n7664) );
  AO22X1 U8529 ( .A0(n4860), .A1(n248), .B0(n4872), .B1(n307), .Y(n7663) );
  AO22X1 U8530 ( .A0(n4846), .A1(n251), .B0(n4852), .B1(n304), .Y(n7662) );
  NOR4X1 U8531 ( .A(n7655), .B(n7654), .C(n7653), .D(n7652), .Y(n7656) );
  AO22X1 U8532 ( .A0(n4880), .A1(n198), .B0(n4886), .B1(n305), .Y(n7655) );
  AO22X1 U8533 ( .A0(n4974), .A1(n196), .B0(n4967), .B1(n2080), .Y(n8878) );
  AO22X1 U8534 ( .A0(n9310), .A1(n570), .B0(n4976), .B1(n2081), .Y(n8877) );
  AO22X1 U8535 ( .A0(n9312), .A1(n571), .B0(n4987), .B1(n2082), .Y(n8876) );
  NOR4X1 U8536 ( .A(n8869), .B(n8868), .C(n8867), .D(n8866), .Y(n8870) );
  AO22X1 U8537 ( .A0(n4974), .A1(n572), .B0(n4967), .B1(n2083), .Y(n8869) );
  AO22X1 U8538 ( .A0(n4980), .A1(n573), .B0(n9309), .B1(n2084), .Y(n8868) );
  AO22X1 U8539 ( .A0(n9312), .A1(n574), .B0(n4987), .B1(n2085), .Y(n8867) );
  NOR4X1 U8540 ( .A(n8319), .B(n8318), .C(n8317), .D(n8316), .Y(n8320) );
  AO22X1 U8541 ( .A0(n4973), .A1(n241), .B0(n4966), .B1(n2086), .Y(n8319) );
  NOR4X1 U8542 ( .A(n8310), .B(n8309), .C(n8308), .D(n8307), .Y(n8311) );
  AO22X1 U8543 ( .A0(n4973), .A1(n575), .B0(n4966), .B1(n2087), .Y(n8310) );
  AO22X1 U8544 ( .A0(n9312), .A1(n667), .B0(n4987), .B1(n2195), .Y(n8702) );
  AO22X1 U8545 ( .A0(n9312), .A1(n577), .B0(n4987), .B1(n2089), .Y(n8693) );
  AO22X1 U8546 ( .A0(n9312), .A1(n578), .B0(n4987), .B1(n2091), .Y(n8986) );
  NOR4X1 U8547 ( .A(n9075), .B(n9074), .C(n9073), .D(n9072), .Y(n9076) );
  AO22X1 U8548 ( .A0(n4974), .A1(n245), .B0(n4967), .B1(n2092), .Y(n9075) );
  AO22X1 U8549 ( .A0(n4977), .A1(n486), .B0(n9309), .B1(n2053), .Y(n9074) );
  AO22X1 U8550 ( .A0(n9312), .A1(n579), .B0(n4987), .B1(n2093), .Y(n9073) );
  NOR4X1 U8551 ( .A(n8793), .B(n8792), .C(n8791), .D(n8790), .Y(n8794) );
  AO22X1 U8552 ( .A0(n4974), .A1(n243), .B0(n4967), .B1(n2094), .Y(n8793) );
  AO22X1 U8553 ( .A0(n9312), .A1(n580), .B0(n4987), .B1(n2095), .Y(n8791) );
  AO22X1 U8554 ( .A0(n9312), .A1(n582), .B0(n4987), .B1(n2097), .Y(n8977) );
  AO22X1 U8555 ( .A0(n4969), .A1(n199), .B0(n4965), .B1(n306), .Y(n7830) );
  NOR4X1 U8556 ( .A(n9066), .B(n9065), .C(n9064), .D(n9063), .Y(n9067) );
  AO22X1 U8557 ( .A0(n4974), .A1(n583), .B0(n4967), .B1(n2098), .Y(n9066) );
  AO22X1 U8558 ( .A0(n4979), .A1(n668), .B0(n9309), .B1(n2196), .Y(n9065) );
  AO22X1 U8559 ( .A0(n9312), .A1(n584), .B0(n4987), .B1(n2099), .Y(n9064) );
  NOR4X1 U8560 ( .A(n8784), .B(n8783), .C(n8782), .D(n8781), .Y(n8785) );
  AO22X1 U8561 ( .A0(n4974), .A1(n585), .B0(n4967), .B1(n2100), .Y(n8784) );
  AO22X1 U8562 ( .A0(n9312), .A1(n586), .B0(n4987), .B1(n2101), .Y(n8782) );
  NOR4X1 U8563 ( .A(n8040), .B(n8039), .C(n8038), .D(n8037), .Y(n8041) );
  AO22X1 U8564 ( .A0(n4969), .A1(n193), .B0(n4965), .B1(n717), .Y(n8040) );
  AO22X1 U8565 ( .A0(n4978), .A1(n587), .B0(n4976), .B1(n2102), .Y(n8039) );
  NOR4X1 U8566 ( .A(n7424), .B(n7423), .C(n7422), .D(n7421), .Y(n7425) );
  AO22X1 U8567 ( .A0(n4977), .A1(n588), .B0(n9309), .B1(n2103), .Y(n7423) );
  NOR4X1 U8568 ( .A(n6699), .B(n6698), .C(n6697), .D(n6696), .Y(n6700) );
  NOR4X1 U8569 ( .A(n8031), .B(n8030), .C(n8029), .D(n8028), .Y(n8032) );
  AO22X1 U8570 ( .A0(n4969), .A1(n216), .B0(n4966), .B1(n718), .Y(n8031) );
  AO22X1 U8571 ( .A0(n4978), .A1(n589), .B0(n4976), .B1(n2104), .Y(n8030) );
  NOR4X1 U8572 ( .A(n8613), .B(n8612), .C(n8611), .D(n8610), .Y(n8614) );
  AO22X1 U8573 ( .A0(n4973), .A1(n244), .B0(n4966), .B1(n2105), .Y(n8613) );
  NOR4X1 U8574 ( .A(n8222), .B(n8221), .C(n8220), .D(n8219), .Y(n8223) );
  AO22X1 U8575 ( .A0(n4973), .A1(n194), .B0(n4966), .B1(n2106), .Y(n8222) );
  NOR4X1 U8576 ( .A(n8416), .B(n8415), .C(n8414), .D(n8413), .Y(n8417) );
  AO22X1 U8577 ( .A0(n4973), .A1(n292), .B0(n4966), .B1(n2107), .Y(n8416) );
  AO22X1 U8578 ( .A0(n4979), .A1(n590), .B0(n9309), .B1(n2108), .Y(n8415) );
  AO22X1 U8579 ( .A0(n9312), .A1(n265), .B0(n4986), .B1(n2109), .Y(n8414) );
  AO22X1 U8580 ( .A0(n4977), .A1(n591), .B0(n4976), .B1(n2110), .Y(n7414) );
  NOR4X1 U8581 ( .A(n8604), .B(n8603), .C(n8602), .D(n8601), .Y(n8605) );
  AO22X1 U8582 ( .A0(n4973), .A1(n592), .B0(n4966), .B1(n2111), .Y(n8604) );
  NOR4X1 U8583 ( .A(n8213), .B(n8212), .C(n8211), .D(n8210), .Y(n8214) );
  AO22X1 U8584 ( .A0(n4973), .A1(n593), .B0(n4966), .B1(n2112), .Y(n8213) );
  NOR4X1 U8585 ( .A(n6690), .B(n6689), .C(n6688), .D(n6687), .Y(n6691) );
  AO22X1 U8586 ( .A0(n4972), .A1(n195), .B0(n4967), .B1(n2197), .Y(n7346) );
  AO22X1 U8587 ( .A0(n4973), .A1(n594), .B0(n4966), .B1(n2113), .Y(n8407) );
  AO22X1 U8588 ( .A0(n4979), .A1(n595), .B0(n4976), .B1(n2114), .Y(n8406) );
  AO22X1 U8589 ( .A0(n9312), .A1(n266), .B0(n4986), .B1(n2115), .Y(n8405) );
  NOR4X1 U8590 ( .A(n7172), .B(n7171), .C(n7170), .D(n7169), .Y(n7173) );
  AO22X1 U8591 ( .A0(n4972), .A1(n669), .B0(n4967), .B1(n2198), .Y(n7337) );
  NOR4X1 U8592 ( .A(n7163), .B(n7162), .C(n7161), .D(n7160), .Y(n7164) );
  AO22X1 U8593 ( .A0(n4972), .A1(n596), .B0(n4967), .B1(n2116), .Y(n7163) );
  AO22X1 U8594 ( .A0(n4992), .A1(n597), .B0(n4981), .B1(n2117), .Y(n7161) );
  NAND2XL U8595 ( .A(n8718), .B(n8717), .Y(n8719) );
  NAND2XL U8596 ( .A(n7028), .B(n7029), .Y(n6940) );
  AO22X1 U8597 ( .A0(DCACHE_addr[29]), .A1(mem_read_D), .B0(net113608), .B1(
        n11541), .Y(n4772) );
  NAND4BBX4 U8598 ( .AN(n4579), .BN(n4580), .C(n6037), .D(n6036), .Y(n9328) );
  NAND3XL U8599 ( .A(n9556), .B(n9572), .C(n4614), .Y(n4579) );
  NAND3XL U8600 ( .A(n4651), .B(n4018), .C(n9554), .Y(n4580) );
  INVXL U8601 ( .A(n8351), .Y(n8352) );
  INVXL U8602 ( .A(n159), .Y(n7878) );
  AOI2BB1X1 U8603 ( .A0N(n8159), .A1N(n8158), .B0(n9262), .Y(n8160) );
  AOI2BB1X1 U8604 ( .A0N(n8715), .A1N(n6454), .B0(n6453), .Y(n6458) );
  CLKINVX1 U8605 ( .A(n9273), .Y(n8998) );
  CLKMX2X2 U8606 ( .A(n9280), .B(n9279), .S0(n9164), .Y(n6667) );
  CLKINVX1 U8607 ( .A(n9127), .Y(n6665) );
  AOI211X1 U8608 ( .A0(n6489), .A1(n6488), .B0(n6631), .C0(n6618), .Y(n6490)
         );
  NAND4XL U8609 ( .A(n7853), .B(n7856), .C(n8524), .D(n6634), .Y(n6488) );
  AOI2BB1XL U8610 ( .A0N(n6487), .A1N(n7852), .B0(n8525), .Y(n6489) );
  NAND2XL U8611 ( .A(n9014), .B(n9171), .Y(n9016) );
  NAND2XL U8612 ( .A(n9142), .B(\i_MIPS/n340 ), .Y(n9162) );
  CLKINVX1 U8613 ( .A(n4441), .Y(n7621) );
  NAND2XL U8614 ( .A(n8516), .B(n159), .Y(n7884) );
  OA22X2 U8615 ( .A0(net112455), .A1(n961), .B0(net112331), .B1(n2486), .Y(
        n6379) );
  OA22X2 U8616 ( .A0(net112239), .A1(n962), .B0(net112163), .B1(n2487), .Y(
        n6378) );
  OA22X1 U8617 ( .A0(net112043), .A1(n1428), .B0(net111919), .B1(n3041), .Y(
        n6377) );
  NAND4X1 U8618 ( .A(n7054), .B(n7053), .C(n7052), .D(n7051), .Y(n11435) );
  OA22X1 U8619 ( .A0(net112463), .A1(n1429), .B0(net112339), .B1(n3042), .Y(
        n7053) );
  OA22X1 U8620 ( .A0(net112051), .A1(n1430), .B0(net111927), .B1(n3043), .Y(
        n7051) );
  NAND2XL U8621 ( .A(n8151), .B(n8150), .Y(n8162) );
  OA22X1 U8622 ( .A0(net112473), .A1(n2833), .B0(net112349), .B1(n841), .Y(
        n7732) );
  OA22XL U8623 ( .A0(net112241), .A1(n1578), .B0(net112159), .B1(n3191), .Y(
        n7731) );
  OA22X1 U8624 ( .A0(net112061), .A1(n2834), .B0(net111937), .B1(n842), .Y(
        n7730) );
  OAI221XL U8625 ( .A0(n9275), .A1(n9136), .B0(n8641), .B1(n8886), .C0(n4501), 
        .Y(n8671) );
  NAND2XL U8626 ( .A(n7847), .B(n7846), .Y(n7712) );
  NAND2XL U8627 ( .A(n8068), .B(n8067), .Y(n8082) );
  NAND2XL U8628 ( .A(n8922), .B(n7971), .Y(n7980) );
  NAND2XL U8629 ( .A(n7781), .B(n8517), .Y(n7800) );
  NAND2XL U8630 ( .A(n7186), .B(n7099), .Y(n6477) );
  NAND2XL U8631 ( .A(n8901), .B(n8905), .Y(n8931) );
  NAND2XL U8632 ( .A(n8512), .B(n8543), .Y(n8553) );
  NAND2XL U8633 ( .A(n8426), .B(n8435), .Y(n8429) );
  NAND2XL U8634 ( .A(n8346), .B(n8351), .Y(n8338) );
  NAND2XL U8635 ( .A(n8095), .B(n8080), .Y(n8079) );
  NAND2X1 U8636 ( .A(n4683), .B(n5591), .Y(n9138) );
  NAND2XL U8637 ( .A(n8920), .B(n8925), .Y(n8258) );
  NAND2X1 U8638 ( .A(n9268), .B(\i_MIPS/n341 ), .Y(n9257) );
  CLKMX2X2 U8639 ( .A(n6743), .B(n6742), .S0(n5588), .Y(net106535) );
  NOR4X1 U8640 ( .A(n6732), .B(n6731), .C(n6730), .D(n6729), .Y(n6743) );
  NOR4X1 U8641 ( .A(n6741), .B(n6740), .C(n6739), .D(n6738), .Y(n6742) );
  NOR4X1 U8642 ( .A(n6553), .B(n6552), .C(n6551), .D(n6550), .Y(n6564) );
  NOR4X1 U8643 ( .A(n6562), .B(n6561), .C(n6560), .D(n6559), .Y(n6563) );
  CLKMX2X2 U8644 ( .A(n6526), .B(n6525), .S0(net108963), .Y(net106881) );
  NOR4X1 U8645 ( .A(n6507), .B(n6506), .C(n6505), .D(n6504), .Y(n6526) );
  NOR4X1 U8646 ( .A(n6524), .B(n6523), .C(n6522), .D(n6521), .Y(n6525) );
  NAND2XL U8647 ( .A(n3675), .B(\i_MIPS/n370 ), .Y(n7622) );
  NAND2XL U8648 ( .A(n8432), .B(n8431), .Y(n8440) );
  INVXL U8649 ( .A(n8922), .Y(n8254) );
  NAND4X1 U8650 ( .A(n6963), .B(n6962), .C(n6961), .D(n6960), .Y(n11434) );
  OA22X2 U8651 ( .A0(net112461), .A1(n963), .B0(net112337), .B1(n2488), .Y(
        n6962) );
  OA22X2 U8652 ( .A0(net112235), .A1(n964), .B0(net112165), .B1(n2489), .Y(
        n6961) );
  OA22X1 U8653 ( .A0(net112049), .A1(n1431), .B0(net111925), .B1(n3044), .Y(
        n6960) );
  OA22X1 U8654 ( .A0(net112237), .A1(n1432), .B0(net112155), .B1(n3045), .Y(
        n8595) );
  NAND4X1 U8655 ( .A(n6883), .B(n6882), .C(n6881), .D(n6880), .Y(n11491) );
  OA22X2 U8656 ( .A0(net112461), .A1(n967), .B0(net112337), .B1(n2492), .Y(
        n6882) );
  OA22X2 U8657 ( .A0(net112235), .A1(n922), .B0(net112165), .B1(n2493), .Y(
        n6881) );
  OA22X1 U8658 ( .A0(net112049), .A1(n1433), .B0(net111925), .B1(n3046), .Y(
        n6880) );
  NAND4X1 U8659 ( .A(n8972), .B(n8971), .C(n8970), .D(n8969), .Y(n11506) );
  OA22X2 U8660 ( .A0(net112491), .A1(n968), .B0(net112367), .B1(n2494), .Y(
        n8971) );
  OA22X1 U8661 ( .A0(net112239), .A1(n2835), .B0(net112153), .B1(n843), .Y(
        n8970) );
  OA22X2 U8662 ( .A0(net112671), .A1(n969), .B0(net112569), .B1(n2495), .Y(
        n8972) );
  OA22X2 U8663 ( .A0(net112487), .A1(n970), .B0(net112363), .B1(n2496), .Y(
        n8687) );
  OA22X1 U8664 ( .A0(net112237), .A1(n1434), .B0(net112155), .B1(n3047), .Y(
        n8686) );
  OA22X2 U8665 ( .A0(net112665), .A1(n971), .B0(net112565), .B1(n2497), .Y(
        n8688) );
  OA22X2 U8666 ( .A0(net112483), .A1(n920), .B0(net112359), .B1(n2498), .Y(
        n8399) );
  OA22X1 U8667 ( .A0(net112235), .A1(n2836), .B0(net112153), .B1(n844), .Y(
        n8398) );
  OA22X1 U8668 ( .A0(net112481), .A1(n1435), .B0(net112357), .B1(n3048), .Y(
        n8205) );
  OA22X2 U8669 ( .A0(net112233), .A1(n972), .B0(net112151), .B1(n2499), .Y(
        n8204) );
  OA22X2 U8670 ( .A0(net112665), .A1(n973), .B0(net112563), .B1(n2500), .Y(
        n8206) );
  NAND4X1 U8671 ( .A(n7066), .B(n7065), .C(n7064), .D(n7063), .Y(n11497) );
  OA22X1 U8672 ( .A0(net112463), .A1(n1436), .B0(net112339), .B1(n3049), .Y(
        n7065) );
  OA22X1 U8673 ( .A0(net112051), .A1(n1437), .B0(net111927), .B1(n3050), .Y(
        n7063) );
  NAND4X1 U8674 ( .A(n6975), .B(n6974), .C(n6973), .D(n6972), .Y(n11496) );
  OA22X2 U8675 ( .A0(net112461), .A1(n974), .B0(net112337), .B1(n2501), .Y(
        n6974) );
  OA22X1 U8676 ( .A0(net112049), .A1(n1438), .B0(net111925), .B1(n3051), .Y(
        n6972) );
  OA22X2 U8677 ( .A0(net112459), .A1(n975), .B0(net112335), .B1(n2502), .Y(
        n6799) );
  OA22X2 U8678 ( .A0(net112235), .A1(n976), .B0(net112165), .B1(n2503), .Y(
        n6798) );
  OA22X1 U8679 ( .A0(net112047), .A1(n1439), .B0(net111923), .B1(n3052), .Y(
        n6797) );
  CLKMX2X2 U8680 ( .A(n9236), .B(n9235), .S0(n5587), .Y(n9254) );
  NAND2XL U8681 ( .A(n6771), .B(n7179), .Y(n6772) );
  CLKINVX1 U8682 ( .A(n6587), .Y(n6594) );
  CLKINVX1 U8683 ( .A(n6771), .Y(n6844) );
  NAND2XL U8684 ( .A(n6847), .B(n6846), .Y(n6775) );
  NAND2XL U8685 ( .A(n3741), .B(n8823), .Y(n8808) );
  CLKINVX1 U8686 ( .A(n7354), .Y(n7273) );
  NAND2XL U8687 ( .A(n7359), .B(n7457), .Y(n7360) );
  CLKMX2X2 U8688 ( .A(n8639), .B(n8638), .S0(n5587), .Y(n8672) );
  NOR4X1 U8689 ( .A(n8628), .B(n8627), .C(n8626), .D(n8625), .Y(n8639) );
  NAND2XL U8690 ( .A(n7546), .B(n3670), .Y(n7554) );
  CLKINVX1 U8691 ( .A(n8997), .Y(n9013) );
  NAND2XL U8692 ( .A(n3634), .B(n7461), .Y(n7469) );
  CLKINVX1 U8693 ( .A(n11226), .Y(n9151) );
  NAND2XL U8694 ( .A(n7463), .B(n3632), .Y(n7468) );
  NAND2XL U8695 ( .A(n8803), .B(n8802), .Y(n8811) );
  CLKINVX1 U8696 ( .A(n8648), .Y(n6652) );
  AND2XL U8697 ( .A(net111409), .B(n10380), .Y(n4595) );
  CLKMX2X2 U8698 ( .A(n7313), .B(n7312), .S0(n5588), .Y(n7314) );
  CLKMX2X2 U8699 ( .A(n8580), .B(n8579), .S0(n5588), .Y(n8581) );
  NOR4X1 U8700 ( .A(n8569), .B(n8568), .C(n8567), .D(n8566), .Y(n8580) );
  NOR4X1 U8701 ( .A(n7996), .B(n7995), .C(n7994), .D(n7993), .Y(n8007) );
  NOR4X1 U8702 ( .A(n8237), .B(n8236), .C(n8235), .D(n8234), .Y(n8248) );
  CLKMX2X2 U8703 ( .A(n8475), .B(n8474), .S0(n5587), .Y(net103479) );
  NOR4X1 U8704 ( .A(n8464), .B(n8463), .C(n8462), .D(n8461), .Y(n8475) );
  NAND2XL U8705 ( .A(n7459), .B(n7458), .Y(n7275) );
  NAND2XL U8706 ( .A(n7562), .B(n7550), .Y(n7551) );
  NAND2XL U8707 ( .A(n7355), .B(n7354), .Y(n7363) );
  AO21X1 U8708 ( .A0(n11227), .A1(n11226), .B0(n11225), .Y(n11581) );
  INVXL U8709 ( .A(n11224), .Y(n11227) );
  MX2XL U8710 ( .A(\i_MIPS/n366 ), .B(\i_MIPS/n365 ), .S0(n3524), .Y(n8732) );
  CLKMX2X2 U8711 ( .A(n8642), .B(n8272), .S0(n5589), .Y(n9128) );
  CLKMX2X2 U8712 ( .A(n6414), .B(n6413), .S0(\i_MIPS/IR_ID[25] ), .Y(n6415) );
  NOR4X1 U8713 ( .A(n6403), .B(n6402), .C(n6401), .D(n6400), .Y(n6414) );
  NOR4X1 U8714 ( .A(n7129), .B(n7128), .C(n7127), .D(n7126), .Y(n7140) );
  CLKMX2X2 U8715 ( .A(n7088), .B(n7087), .S0(n5588), .Y(n7089) );
  NOR4X1 U8716 ( .A(n7077), .B(n7076), .C(n7075), .D(n7074), .Y(n7088) );
  CLKMX2X2 U8717 ( .A(n6324), .B(n6323), .S0(\i_MIPS/IR_ID[25] ), .Y(n6325) );
  NOR4X1 U8718 ( .A(n6313), .B(n6312), .C(n6311), .D(n6310), .Y(n6324) );
  CLKMX2X2 U8719 ( .A(n6822), .B(n6821), .S0(\i_MIPS/IR_ID[25] ), .Y(n6823) );
  NOR4X1 U8720 ( .A(n8835), .B(n8834), .C(n8833), .D(n8832), .Y(n8846) );
  CLKMX2X2 U8721 ( .A(n7392), .B(n7391), .S0(n5588), .Y(net105373) );
  CLKMX2X2 U8722 ( .A(n7230), .B(n7229), .S0(n5588), .Y(net105666) );
  NOR4X1 U8723 ( .A(n7219), .B(n7218), .C(n7217), .D(n7216), .Y(n7230) );
  CLKMX2X2 U8724 ( .A(n7911), .B(n7910), .S0(n5588), .Y(net104440) );
  NOR4X1 U8725 ( .A(n7900), .B(n7899), .C(n7898), .D(n7897), .Y(n7911) );
  CLKMX2X2 U8726 ( .A(n7697), .B(n7696), .S0(n5589), .Y(n8433) );
  INVXL U8727 ( .A(n8925), .Y(n8259) );
  INVXL U8728 ( .A(n8712), .Y(n6454) );
  MX2XL U8729 ( .A(\i_MIPS/n342 ), .B(\i_MIPS/n343 ), .S0(n3524), .Y(n9127) );
  MX2XL U8730 ( .A(\i_MIPS/n369 ), .B(\i_MIPS/n368 ), .S0(n3524), .Y(n8800) );
  MX2XL U8731 ( .A(\i_MIPS/n343 ), .B(\i_MIPS/n344 ), .S0(n3524), .Y(n9273) );
  MX2XL U8732 ( .A(\i_MIPS/n368 ), .B(\i_MIPS/n367 ), .S0(n3524), .Y(n8731) );
  INVXL U8733 ( .A(n7865), .Y(n6954) );
  NAND2XL U8734 ( .A(n286), .B(n3636), .Y(n6439) );
  CLKINVX1 U8735 ( .A(n8080), .Y(n8081) );
  CLKMX2X2 U8736 ( .A(n7352), .B(n7351), .S0(net108963), .Y(net105425) );
  CLKMX2X2 U8737 ( .A(n8228), .B(n8227), .S0(net108959), .Y(net103869) );
  AND2X2 U8738 ( .A(n4656), .B(n4584), .Y(n4630) );
  CLKINVX1 U8739 ( .A(n10410), .Y(n5017) );
  NAND2XL U8740 ( .A(n10409), .B(n10408), .Y(n10410) );
  CLKBUFX3 U8741 ( .A(\i_MIPS/n336 ), .Y(net113089) );
  CLKMX2X2 U8742 ( .A(n7670), .B(n7669), .S0(n5588), .Y(n7672) );
  CLKBUFX3 U8743 ( .A(\i_MIPS/n336 ), .Y(net113087) );
  INVX1 U8744 ( .A(n6657), .Y(n6654) );
  AND2XL U8745 ( .A(n8521), .B(n8250), .Y(n6485) );
  AO22X1 U8746 ( .A0(n5000), .A1(n200), .B0(n4998), .B1(n252), .Y(n9315) );
  AO22X1 U8747 ( .A0(n5001), .A1(n249), .B0(n4998), .B1(n1868), .Y(n9298) );
  AO22X1 U8748 ( .A0(n9118), .A1(n296), .B0(n4901), .B1(n1869), .Y(n6559) );
  AO22X1 U8749 ( .A0(n9118), .A1(n297), .B0(n4901), .B1(n1870), .Y(n6550) );
  AO22X1 U8750 ( .A0(n432), .A1(n200), .B0(n4836), .B1(n252), .Y(n9227) );
  CLKMX2X2 U8751 ( .A(n8139), .B(n8138), .S0(net108959), .Y(net104023) );
  AO22X1 U8752 ( .A0(n4895), .A1(n298), .B0(n4891), .B1(n1871), .Y(n6560) );
  AO22X1 U8753 ( .A0(n4895), .A1(n299), .B0(n4891), .B1(n1872), .Y(n6551) );
  INVXL U8754 ( .A(n8516), .Y(n7861) );
  AND3XL U8755 ( .A(n8261), .B(n4802), .C(n8818), .Y(n7466) );
  CLKMX2X2 U8756 ( .A(n7178), .B(n7177), .S0(net108963), .Y(net105735) );
  NOR4X1 U8757 ( .A(n8055), .B(n8054), .C(n8053), .D(n8052), .Y(n8066) );
  INVXL U8758 ( .A(n11389), .Y(n4750) );
  NOR4X1 U8759 ( .A(n9032), .B(n9031), .C(n9030), .D(n9029), .Y(n9043) );
  NAND3BXL U8760 ( .AN(n11360), .B(n11228), .C(n4793), .Y(n11161) );
  NAND3BX1 U8761 ( .AN(n9808), .B(n9688), .C(\i_MIPS/n324 ), .Y(
        \i_MIPS/Control_ID/n10 ) );
  NAND2X1 U8762 ( .A(\i_MIPS/n322 ), .B(\i_MIPS/n332 ), .Y(n11165) );
  CLKINVX1 U8763 ( .A(n4793), .Y(n11358) );
  NAND2X1 U8764 ( .A(n3303), .B(n1609), .Y(n11521) );
  NAND2X1 U8765 ( .A(n1608), .B(n3295), .Y(n11524) );
  NAND2X1 U8766 ( .A(n10679), .B(n10678), .Y(n11519) );
  NOR2BX1 U8767 ( .AN(n4717), .B(n9808), .Y(n4637) );
  AND2X2 U8768 ( .A(n4637), .B(\i_MIPS/n332 ), .Y(n4638) );
  NAND2X1 U8769 ( .A(\i_MIPS/Control_ID/n15 ), .B(\i_MIPS/Control_ID/n10 ), 
        .Y(\i_MIPS/control_out[7] ) );
  CLKBUFX3 U8770 ( .A(n5918), .Y(n5940) );
  CLKBUFX3 U8771 ( .A(n5930), .Y(n5939) );
  INVX12 U8772 ( .A(n1813), .Y(mem_addr_D[27]) );
  CLKINVX1 U8773 ( .A(net113667), .Y(net113983) );
  INVX12 U8774 ( .A(n1811), .Y(mem_addr_D[25]) );
  MXI2X2 U8775 ( .A(n10690), .B(n10689), .S0(n5491), .Y(n10691) );
  AOI222XL U8776 ( .A0(net109791), .A1(n11419), .B0(mem_rdata_D[30]), .B1(n116), .C0(n12967), .C1(net109801), .Y(n10690) );
  INVXL U8777 ( .A(n11418), .Y(n10480) );
  MXI2X2 U8778 ( .A(n10402), .B(n10401), .S0(n5497), .Y(n10403) );
  INVXL U8779 ( .A(n11417), .Y(n10401) );
  INVXL U8780 ( .A(n11416), .Y(n10468) );
  MXI2X2 U8781 ( .A(n10418), .B(n10417), .S0(n5496), .Y(n10419) );
  INVXL U8782 ( .A(n11415), .Y(n10417) );
  AOI222XL U8783 ( .A0(net109791), .A1(n11415), .B0(mem_rdata_D[26]), .B1(n117), .C0(n12971), .C1(net109801), .Y(n10418) );
  MXI2X2 U8784 ( .A(n10430), .B(n10429), .S0(n5496), .Y(n10431) );
  INVXL U8785 ( .A(n11414), .Y(n10429) );
  AOI222XL U8786 ( .A0(net109791), .A1(n11414), .B0(mem_rdata_D[25]), .B1(n117), .C0(n12972), .C1(net109801), .Y(n10430) );
  INVXL U8787 ( .A(n11413), .Y(n10575) );
  AOI222XL U8788 ( .A0(net109791), .A1(n11413), .B0(mem_rdata_D[24]), .B1(n117), .C0(n12973), .C1(net109801), .Y(n10576) );
  INVXL U8789 ( .A(n11412), .Y(n10562) );
  AOI222XL U8790 ( .A0(net109791), .A1(n11412), .B0(mem_rdata_D[23]), .B1(n117), .C0(n12974), .C1(net109801), .Y(n10563) );
  INVXL U8791 ( .A(n11411), .Y(n10550) );
  AOI222XL U8792 ( .A0(net109791), .A1(n11411), .B0(mem_rdata_D[22]), .B1(n116), .C0(n12975), .C1(net109801), .Y(n10551) );
  MXI2X2 U8793 ( .A(n10539), .B(n10538), .S0(n5494), .Y(n10540) );
  INVXL U8794 ( .A(n11410), .Y(n10538) );
  AOI222XL U8795 ( .A0(net109791), .A1(n11410), .B0(mem_rdata_D[21]), .B1(n116), .C0(n12976), .C1(net109801), .Y(n10539) );
  MXI2X2 U8796 ( .A(n10527), .B(n10526), .S0(n5494), .Y(n10528) );
  INVXL U8797 ( .A(n11409), .Y(n10526) );
  AOI222XL U8798 ( .A0(net109791), .A1(n11409), .B0(mem_rdata_D[20]), .B1(n117), .C0(n12977), .C1(net109801), .Y(n10527) );
  MXI2X2 U8799 ( .A(n10179), .B(n10178), .S0(n5497), .Y(n10180) );
  INVXL U8800 ( .A(n11408), .Y(n10178) );
  MXI2X2 U8801 ( .A(n10615), .B(n10614), .S0(n5492), .Y(n10616) );
  INVXL U8802 ( .A(n11407), .Y(n10614) );
  AOI222XL U8803 ( .A0(net109791), .A1(n11407), .B0(mem_rdata_D[18]), .B1(n116), .C0(n12979), .C1(net109801), .Y(n10615) );
  AOI222XL U8804 ( .A0(net109791), .A1(n11406), .B0(mem_rdata_D[17]), .B1(n117), .C0(n12980), .C1(net109801), .Y(n10602) );
  INVXL U8805 ( .A(n11405), .Y(n10455) );
  MXI2X2 U8806 ( .A(n10193), .B(n10192), .S0(n5497), .Y(n10194) );
  MXI2X2 U8807 ( .A(n10442), .B(n10441), .S0(n5496), .Y(n10443) );
  MXI2X2 U8808 ( .A(n10590), .B(n10589), .S0(n5492), .Y(n10591) );
  INVXL U8809 ( .A(n11399), .Y(n10589) );
  INVXL U8810 ( .A(n11398), .Y(n10771) );
  MXI2X2 U8811 ( .A(n10745), .B(n10744), .S0(n5491), .Y(n10746) );
  INVXL U8812 ( .A(n11396), .Y(n10744) );
  MXI2X2 U8813 ( .A(net100025), .B(net100026), .S0(n5497), .Y(n10169) );
  MXI2X2 U8814 ( .A(n10759), .B(n10758), .S0(n5491), .Y(n10760) );
  INVXL U8815 ( .A(n11395), .Y(n10758) );
  MXI2X2 U8816 ( .A(n10155), .B(n10154), .S0(n5497), .Y(n10156) );
  INVXL U8817 ( .A(n11394), .Y(n10154) );
  AOI222XL U8818 ( .A0(net109791), .A1(n11394), .B0(mem_rdata_D[4]), .B1(n116), 
        .C0(n12993), .C1(net109801), .Y(n10155) );
  INVXL U8819 ( .A(n11393), .Y(n10513) );
  MXI2X2 U8820 ( .A(n10808), .B(n10807), .S0(n5489), .Y(n10809) );
  INVXL U8821 ( .A(n11402), .Y(n10807) );
  INVXL U8822 ( .A(n11401), .Y(n10795) );
  MXI2X2 U8823 ( .A(n10784), .B(n10783), .S0(n5490), .Y(n10785) );
  INVXL U8824 ( .A(n11400), .Y(n10783) );
  MXI2X2 U8825 ( .A(n10824), .B(n10823), .S0(n5489), .Y(n10825) );
  INVXL U8826 ( .A(n11397), .Y(n10823) );
  MXI2X2 U8827 ( .A(n11176), .B(n11175), .S0(n5495), .Y(n11177) );
  INVXL U8828 ( .A(n11392), .Y(n11175) );
  MXI2X2 U8829 ( .A(n10845), .B(n10844), .S0(n5489), .Y(n10846) );
  INVXL U8830 ( .A(n11391), .Y(n10844) );
  NAND2XL U8831 ( .A(n12962), .B(net113087), .Y(net98950) );
  MXI2X2 U8832 ( .A(n11215), .B(n11214), .S0(n5496), .Y(n11216) );
  INVXL U8833 ( .A(n11451), .Y(n11214) );
  AOI222XL U8834 ( .A0(n5488), .A1(n11451), .B0(mem_rdata_D[63]), .B1(n117), 
        .C0(n12966), .C1(n5484), .Y(n11215) );
  MXI2X2 U8835 ( .A(n10687), .B(n10686), .S0(n5491), .Y(n10688) );
  AOI222XL U8836 ( .A0(n5480), .A1(n11481), .B0(mem_rdata_D[94]), .B1(n117), 
        .C0(n12967), .C1(n5477), .Y(n10687) );
  INVXL U8837 ( .A(n11480), .Y(n10477) );
  MXI2X2 U8838 ( .A(n10399), .B(n10398), .S0(n5497), .Y(n10400) );
  INVXL U8839 ( .A(n11479), .Y(n10398) );
  INVXL U8840 ( .A(n11478), .Y(n10465) );
  INVXL U8841 ( .A(n11477), .Y(n10414) );
  MXI2X2 U8842 ( .A(n10427), .B(n10426), .S0(n5496), .Y(n10428) );
  INVXL U8843 ( .A(n11476), .Y(n10426) );
  AOI222XL U8844 ( .A0(n5479), .A1(n11476), .B0(mem_rdata_D[89]), .B1(n116), 
        .C0(n12972), .C1(n5476), .Y(n10427) );
  MXI2X2 U8845 ( .A(n10573), .B(n10572), .S0(n5493), .Y(n10574) );
  INVXL U8846 ( .A(n11475), .Y(n10572) );
  INVXL U8847 ( .A(n11474), .Y(n10559) );
  INVXL U8848 ( .A(n11473), .Y(n10547) );
  INVXL U8849 ( .A(n11472), .Y(n10535) );
  MXI2X2 U8850 ( .A(n10524), .B(n10523), .S0(n5494), .Y(n10525) );
  INVXL U8851 ( .A(n11471), .Y(n10523) );
  INVXL U8852 ( .A(n11470), .Y(n10175) );
  AOI222XL U8853 ( .A0(n5479), .A1(n11470), .B0(mem_rdata_D[83]), .B1(n116), 
        .C0(n12978), .C1(n5476), .Y(n10176) );
  INVXL U8854 ( .A(n11469), .Y(n10611) );
  INVXL U8855 ( .A(n11467), .Y(n10452) );
  MXI2X2 U8856 ( .A(n10439), .B(n10438), .S0(n5496), .Y(n10440) );
  INVXL U8857 ( .A(n11465), .Y(n10438) );
  AOI222XL U8858 ( .A0(n5479), .A1(n11465), .B0(mem_rdata_D[78]), .B1(n116), 
        .C0(n12983), .C1(n5476), .Y(n10439) );
  INVXL U8859 ( .A(n11461), .Y(n10586) );
  INVXL U8860 ( .A(n11460), .Y(n10768) );
  MXI2X2 U8861 ( .A(n10742), .B(n10741), .S0(n5491), .Y(n10743) );
  INVXL U8862 ( .A(n11458), .Y(n10741) );
  AOI222XL U8863 ( .A0(n5480), .A1(n11458), .B0(mem_rdata_D[71]), .B1(n117), 
        .C0(n12990), .C1(n5477), .Y(n10742) );
  MXI2X2 U8864 ( .A(n10167), .B(net100029), .S0(n5489), .Y(n10168) );
  INVXL U8865 ( .A(net98121), .Y(net100029) );
  AOI222XL U8866 ( .A0(n5479), .A1(net98121), .B0(mem_rdata_D[70]), .B1(n116), 
        .C0(n12991), .C1(n5476), .Y(n10167) );
  MXI2X2 U8867 ( .A(n10756), .B(n10755), .S0(n5491), .Y(n10757) );
  INVXL U8868 ( .A(n11457), .Y(n10755) );
  AOI222XL U8869 ( .A0(n5480), .A1(n11457), .B0(mem_rdata_D[69]), .B1(n116), 
        .C0(n12992), .C1(n5477), .Y(n10756) );
  MXI2X2 U8870 ( .A(n10149), .B(n10148), .S0(n5489), .Y(n10150) );
  INVXL U8871 ( .A(n11456), .Y(n10148) );
  AOI222XL U8872 ( .A0(n5479), .A1(n11456), .B0(mem_rdata_D[68]), .B1(n116), 
        .C0(n12993), .C1(n5476), .Y(n10149) );
  MXI2X2 U8873 ( .A(n10511), .B(n10510), .S0(n5494), .Y(n10512) );
  INVXL U8874 ( .A(n11455), .Y(n10510) );
  AOI222XL U8875 ( .A0(n5479), .A1(n11455), .B0(mem_rdata_D[67]), .B1(n117), 
        .C0(n12994), .C1(n5476), .Y(n10511) );
  INVXL U8876 ( .A(n11510), .Y(n10395) );
  AOI222XL U8877 ( .A0(n5474), .A1(n11508), .B0(mem_rdata_D[122]), .B1(n116), 
        .C0(n12971), .C1(n5472), .Y(n10412) );
  INVXL U8878 ( .A(n11507), .Y(n10423) );
  MXI2X2 U8879 ( .A(n10557), .B(n10556), .S0(n5493), .Y(n10558) );
  INVXL U8880 ( .A(n11505), .Y(n10556) );
  INVXL U8881 ( .A(n11504), .Y(n10544) );
  INVXL U8882 ( .A(n11503), .Y(n10532) );
  MXI2X2 U8883 ( .A(n10521), .B(n10520), .S0(n5494), .Y(n10522) );
  MXI2X2 U8884 ( .A(n10173), .B(n10172), .S0(n5497), .Y(n10174) );
  INVXL U8885 ( .A(n11501), .Y(n10172) );
  AOI222XL U8886 ( .A0(n5474), .A1(n11501), .B0(mem_rdata_D[115]), .B1(n117), 
        .C0(n12978), .C1(n5472), .Y(n10173) );
  MXI2X2 U8887 ( .A(n10596), .B(n10595), .S0(n5492), .Y(n10597) );
  MXI2X2 U8888 ( .A(n10436), .B(n10435), .S0(n5496), .Y(n10437) );
  MXI2X2 U8889 ( .A(n10584), .B(n10583), .S0(n5492), .Y(n10585) );
  INVXL U8890 ( .A(n11492), .Y(n10583) );
  INVXL U8891 ( .A(n11489), .Y(n10738) );
  MXI2X2 U8892 ( .A(n10165), .B(net100032), .S0(n5495), .Y(n10166) );
  INVXL U8893 ( .A(net98089), .Y(net100032) );
  AOI222XL U8894 ( .A0(n5474), .A1(net98089), .B0(mem_rdata_D[102]), .B1(n116), 
        .C0(n12991), .C1(n5472), .Y(n10165) );
  MXI2X2 U8895 ( .A(n10753), .B(n10752), .S0(n5491), .Y(n10754) );
  INVXL U8896 ( .A(n11488), .Y(n10752) );
  MXI2X2 U8897 ( .A(n10143), .B(n10142), .S0(n5493), .Y(n10144) );
  INVXL U8898 ( .A(n11487), .Y(n10142) );
  AOI222XL U8899 ( .A0(n5474), .A1(n11487), .B0(mem_rdata_D[100]), .B1(n117), 
        .C0(n12993), .C1(n5472), .Y(n10143) );
  MXI2X2 U8900 ( .A(n10141), .B(n10140), .S0(n5497), .Y(n10509) );
  INVXL U8901 ( .A(n11486), .Y(n10140) );
  MXI2X2 U8902 ( .A(n10693), .B(n10692), .S0(n5491), .Y(n10694) );
  AOI222XL U8903 ( .A0(n5487), .A1(n11450), .B0(mem_rdata_D[62]), .B1(n117), 
        .C0(n12967), .C1(n5483), .Y(n10693) );
  MXI2X2 U8904 ( .A(n10484), .B(n10483), .S0(n5494), .Y(n10485) );
  MXI2X2 U8905 ( .A(n10405), .B(n10404), .S0(n5496), .Y(n10406) );
  INVXL U8906 ( .A(n11448), .Y(n10404) );
  MXI2X2 U8907 ( .A(n10421), .B(n10420), .S0(n5496), .Y(n10422) );
  INVXL U8908 ( .A(n11446), .Y(n10420) );
  AOI222XL U8909 ( .A0(n5486), .A1(n11446), .B0(mem_rdata_D[58]), .B1(n116), 
        .C0(n12971), .C1(n5482), .Y(n10421) );
  MXI2X2 U8910 ( .A(n10433), .B(n10432), .S0(n5496), .Y(n10434) );
  INVXL U8911 ( .A(n11445), .Y(n10432) );
  AOI222XL U8912 ( .A0(n5486), .A1(n11445), .B0(mem_rdata_D[57]), .B1(n116), 
        .C0(n12972), .C1(n5482), .Y(n10433) );
  MXI2X2 U8913 ( .A(n10579), .B(n10578), .S0(n5493), .Y(n10580) );
  INVXL U8914 ( .A(n11444), .Y(n10578) );
  AOI222XL U8915 ( .A0(n5487), .A1(n11444), .B0(mem_rdata_D[56]), .B1(n116), 
        .C0(n12973), .C1(n5483), .Y(n10579) );
  MXI2X2 U8916 ( .A(n10566), .B(n10565), .S0(n5493), .Y(n10567) );
  INVXL U8917 ( .A(n11443), .Y(n10565) );
  AOI222XL U8918 ( .A0(n5487), .A1(n11443), .B0(mem_rdata_D[55]), .B1(n116), 
        .C0(n12974), .C1(n5483), .Y(n10566) );
  MXI2X2 U8919 ( .A(n10554), .B(n10553), .S0(n5493), .Y(n10555) );
  INVXL U8920 ( .A(n11442), .Y(n10553) );
  AOI222XL U8921 ( .A0(n5487), .A1(n11442), .B0(mem_rdata_D[54]), .B1(n117), 
        .C0(n12975), .C1(n5483), .Y(n10554) );
  MXI2X2 U8922 ( .A(n10542), .B(n10541), .S0(n5494), .Y(n10543) );
  INVXL U8923 ( .A(n11441), .Y(n10541) );
  MXI2X2 U8924 ( .A(n10530), .B(n10529), .S0(n5494), .Y(n10531) );
  INVXL U8925 ( .A(n11440), .Y(n10529) );
  MXI2X2 U8926 ( .A(n10182), .B(n10181), .S0(n5497), .Y(n10183) );
  INVXL U8927 ( .A(n11439), .Y(n10181) );
  AOI222XL U8928 ( .A0(n5486), .A1(n11439), .B0(mem_rdata_D[51]), .B1(n116), 
        .C0(n12978), .C1(n5482), .Y(n10182) );
  MXI2X2 U8929 ( .A(n10618), .B(n10617), .S0(n5492), .Y(n10619) );
  INVXL U8930 ( .A(n11438), .Y(n10617) );
  INVXL U8931 ( .A(n11436), .Y(n10458) );
  MXI2X2 U8932 ( .A(n10196), .B(n10195), .S0(n5497), .Y(n10197) );
  AOI222XL U8933 ( .A0(n5486), .A1(n11435), .B0(mem_rdata_D[47]), .B1(n117), 
        .C0(n12982), .C1(n5482), .Y(n10196) );
  INVXL U8934 ( .A(n11430), .Y(n10592) );
  MXI2X2 U8935 ( .A(n10775), .B(n10774), .S0(n5490), .Y(n10776) );
  INVXL U8936 ( .A(n11429), .Y(n10774) );
  MXI2X2 U8937 ( .A(n10748), .B(n10747), .S0(n5491), .Y(n10749) );
  INVXL U8938 ( .A(n11427), .Y(n10747) );
  INVXL U8939 ( .A(net98153), .Y(net100023) );
  MXI2X2 U8940 ( .A(n10762), .B(n10761), .S0(n5491), .Y(n10763) );
  INVXL U8941 ( .A(n11426), .Y(n10761) );
  AOI222XL U8942 ( .A0(n5487), .A1(n11426), .B0(mem_rdata_D[37]), .B1(n117), 
        .C0(n12992), .C1(n5483), .Y(n10762) );
  MXI2X2 U8943 ( .A(n10163), .B(n10162), .S0(n5495), .Y(n10164) );
  MXI2X2 U8944 ( .A(n10517), .B(n10516), .S0(n5494), .Y(n10518) );
  INVXL U8945 ( .A(n11424), .Y(n10516) );
  AOI222XL U8946 ( .A0(n5486), .A1(n11424), .B0(mem_rdata_D[35]), .B1(n116), 
        .C0(n12994), .C1(n5482), .Y(n10517) );
  INVXL U8947 ( .A(n11464), .Y(n10804) );
  AOI222XL U8948 ( .A0(n5481), .A1(n11464), .B0(mem_rdata_D[77]), .B1(n116), 
        .C0(n12984), .C1(n5478), .Y(n10805) );
  MXI2X2 U8949 ( .A(n10793), .B(n10792), .S0(n5490), .Y(n10794) );
  INVXL U8950 ( .A(n11463), .Y(n10792) );
  INVXL U8951 ( .A(n11462), .Y(n10780) );
  AOI222XL U8952 ( .A0(n5481), .A1(n11462), .B0(mem_rdata_D[75]), .B1(n116), 
        .C0(n12986), .C1(n5478), .Y(n10781) );
  AOI222XL U8953 ( .A0(n5481), .A1(n11459), .B0(mem_rdata_D[72]), .B1(n116), 
        .C0(n12989), .C1(n5478), .Y(n10821) );
  INVXL U8954 ( .A(n11454), .Y(n11172) );
  INVXL U8955 ( .A(n11453), .Y(n10841) );
  AOI222XL U8956 ( .A0(n5481), .A1(n11453), .B0(mem_rdata_D[65]), .B1(n117), 
        .C0(n12996), .C1(n5478), .Y(n10842) );
  INVXL U8957 ( .A(n11452), .Y(n10854) );
  MXI2X2 U8958 ( .A(n10802), .B(n10801), .S0(n5489), .Y(n10803) );
  INVXL U8959 ( .A(n11495), .Y(n10801) );
  AOI222XL U8960 ( .A0(n5474), .A1(n11495), .B0(mem_rdata_D[109]), .B1(n117), 
        .C0(n12984), .C1(n5473), .Y(n10802) );
  MXI2X2 U8961 ( .A(n10790), .B(n10789), .S0(n5490), .Y(n10791) );
  AOI222XL U8962 ( .A0(n5474), .A1(n11494), .B0(mem_rdata_D[108]), .B1(n117), 
        .C0(n12985), .C1(n5473), .Y(n10790) );
  MXI2X2 U8963 ( .A(n10778), .B(n10777), .S0(n5490), .Y(n10779) );
  MXI2X2 U8964 ( .A(n10818), .B(n10817), .S0(n5489), .Y(n10819) );
  INVXL U8965 ( .A(n11485), .Y(n11169) );
  AOI222XL U8966 ( .A0(n5474), .A1(n11485), .B0(mem_rdata_D[98]), .B1(n117), 
        .C0(n12995), .C1(n5473), .Y(n11170) );
  MXI2X2 U8967 ( .A(n10839), .B(n10838), .S0(n5489), .Y(n10840) );
  INVXL U8968 ( .A(n11484), .Y(n10838) );
  INVXL U8969 ( .A(n11483), .Y(n10851) );
  MXI2X2 U8970 ( .A(n10811), .B(n10810), .S0(n5489), .Y(n10812) );
  INVXL U8971 ( .A(n11432), .Y(n10798) );
  MXI2X2 U8972 ( .A(n10787), .B(n10786), .S0(n5490), .Y(n10788) );
  INVXL U8973 ( .A(n11431), .Y(n10786) );
  AOI222XL U8974 ( .A0(n5488), .A1(n11431), .B0(mem_rdata_D[43]), .B1(n116), 
        .C0(n12986), .C1(n5484), .Y(n10787) );
  MXI2X2 U8975 ( .A(n10827), .B(n10826), .S0(n5489), .Y(n10828) );
  AOI222XL U8976 ( .A0(n5488), .A1(n11428), .B0(mem_rdata_D[40]), .B1(n117), 
        .C0(n12989), .C1(n5484), .Y(n10827) );
  MXI2X2 U8977 ( .A(n11179), .B(n11178), .S0(n5491), .Y(n11180) );
  INVXL U8978 ( .A(n11423), .Y(n11178) );
  AOI222XL U8979 ( .A0(n5488), .A1(n11423), .B0(mem_rdata_D[34]), .B1(n117), 
        .C0(n12995), .C1(n5484), .Y(n11179) );
  MXI2X2 U8980 ( .A(n10848), .B(n10847), .S0(n5489), .Y(n10849) );
  INVXL U8981 ( .A(n11422), .Y(n10847) );
  AOI222XL U8982 ( .A0(n5488), .A1(n11422), .B0(mem_rdata_D[33]), .B1(n116), 
        .C0(n12996), .C1(n5484), .Y(n10848) );
  NAND2X1 U8983 ( .A(n10201), .B(ICACHE_addr[21]), .Y(net99962) );
  MXI2X2 U8984 ( .A(n11210), .B(n11209), .S0(n5494), .Y(n11211) );
  INVXL U8985 ( .A(n11420), .Y(n11209) );
  MXI2X2 U8986 ( .A(n11203), .B(n11202), .S0(n5493), .Y(n11204) );
  INVXL U8987 ( .A(n11513), .Y(n11202) );
  AOI222XL U8988 ( .A0(n5474), .A1(n11513), .B0(mem_rdata_D[127]), .B1(n116), 
        .C0(n5473), .C1(n12966), .Y(n11203) );
  XOR2X1 U8989 ( .A(n10203), .B(ICACHE_addr[10]), .Y(n10270) );
  NAND2X1 U8990 ( .A(n10202), .B(ICACHE_addr[9]), .Y(n10203) );
  XOR2X1 U8991 ( .A(n10290), .B(ICACHE_addr[15]), .Y(n11113) );
  XOR2X1 U8992 ( .A(n10294), .B(ICACHE_addr[13]), .Y(n11098) );
  MXI2X2 U8993 ( .A(n11207), .B(n11206), .S0(n5495), .Y(n11208) );
  INVXL U8994 ( .A(n11482), .Y(n11206) );
  XOR2X1 U8995 ( .A(n10291), .B(ICACHE_addr[19]), .Y(n11029) );
  XOR2X1 U8996 ( .A(n10263), .B(ICACHE_addr[11]), .Y(n11088) );
  XOR2X1 U8997 ( .A(n10204), .B(ICACHE_addr[9]), .Y(n11078) );
  XOR2X1 U8998 ( .A(\i_MIPS/PC/n4 ), .B(ICACHE_addr[1]), .Y(n11002) );
  XOR2X1 U8999 ( .A(n9367), .B(ICACHE_addr[14]), .Y(n10929) );
  XOR2X1 U9000 ( .A(n10262), .B(ICACHE_addr[12]), .Y(n10299) );
  OA22XL U9001 ( .A0(\i_MIPS/ALUin1[24] ), .A1(n4812), .B0(\i_MIPS/ALUin1[25] ), .B1(n3592), .Y(n6675) );
  OA22XL U9002 ( .A0(\i_MIPS/ALUin1[5] ), .A1(n4812), .B0(\i_MIPS/ALUin1[4] ), 
        .B1(n4805), .Y(n6417) );
  OAI221XL U9003 ( .A0(\i_MIPS/ALUin1[10] ), .A1(n4824), .B0(
        \i_MIPS/ALUin1[9] ), .B1(n4816), .C0(n7472), .Y(n8733) );
  OAI221X1 U9004 ( .A0(\i_MIPS/ALUin1[12] ), .A1(n4810), .B0(
        \i_MIPS/ALUin1[11] ), .B1(n4803), .C0(n7105), .Y(n7451) );
  OA22XL U9005 ( .A0(\i_MIPS/ALUin1[10] ), .A1(n4812), .B0(\i_MIPS/ALUin1[9] ), 
        .B1(n4805), .Y(n6854) );
  OA22XL U9006 ( .A0(\i_MIPS/ALUin1[9] ), .A1(n4812), .B0(\i_MIPS/ALUin1[8] ), 
        .B1(n4805), .Y(n6430) );
  NAND2X1 U9007 ( .A(\i_MIPS/ALUin1[29] ), .B(n6659), .Y(n9170) );
  OAI222XL U9008 ( .A0(n5097), .A1(n196), .B0(n5073), .B1(n10835), .C0(n5522), 
        .C1(\i_MIPS/n182 ), .Y(n11578) );
  OAI222XL U9009 ( .A0(n5098), .A1(n245), .B0(n1850), .B1(n5095), .C0(n5523), 
        .C1(\i_MIPS/n208 ), .Y(n11552) );
  OAI222XL U9010 ( .A0(n5097), .A1(n183), .B0(n1841), .B1(n10835), .C0(n5522), 
        .C1(\i_MIPS/n181 ), .Y(n11579) );
  OAI222XL U9011 ( .A0(n5097), .A1(n1802), .B0(n5101), .B1(n10835), .C0(n5522), 
        .C1(\i_MIPS/n180 ), .Y(n11580) );
  XOR2X4 U9012 ( .A(n11385), .B(\i_MIPS/PC/n30 ), .Y(n4640) );
  AO22X2 U9013 ( .A0(n5063), .A1(DCACHE_addr[8]), .B0(n5061), .B1(n11521), .Y(
        n10677) );
  NAND2X1 U9014 ( .A(n6198), .B(n6197), .Y(n6205) );
  NAND4X1 U9015 ( .A(n6196), .B(n6195), .C(n6194), .D(n6302), .Y(n6206) );
  XNOR2XL U9016 ( .A(\i_MIPS/Reg_W[3] ), .B(\i_MIPS/IR_ID[19] ), .Y(n6197) );
  AO22X2 U9017 ( .A0(mem_rdata_I[3]), .A1(n114), .B0(n5465), .B1(n11233), .Y(
        n9517) );
  AO22X2 U9018 ( .A0(mem_rdata_I[31]), .A1(n115), .B0(n5465), .B1(n11261), .Y(
        n11037) );
  AO22X2 U9019 ( .A0(mem_rdata_I[29]), .A1(n114), .B0(n5470), .B1(n11259), .Y(
        n11160) );
  AO22X2 U9020 ( .A0(mem_rdata_I[26]), .A1(n115), .B0(n5467), .B1(n11256), .Y(
        n9706) );
  AO22X2 U9021 ( .A0(mem_rdata_I[25]), .A1(n114), .B0(n5469), .B1(n11255), .Y(
        n10119) );
  AO22X2 U9022 ( .A0(mem_rdata_I[24]), .A1(n115), .B0(n5467), .B1(n11254), .Y(
        n9897) );
  AO22X2 U9023 ( .A0(mem_rdata_I[23]), .A1(n115), .B0(n5467), .B1(n11253), .Y(
        n9921) );
  AO22X2 U9024 ( .A0(mem_rdata_I[21]), .A1(n115), .B0(n5467), .B1(n11251), .Y(
        n9873) );
  AO22X2 U9025 ( .A0(mem_rdata_I[20]), .A1(n115), .B0(n5468), .B1(n11250), .Y(
        n10017) );
  AO22X2 U9026 ( .A0(mem_rdata_I[19]), .A1(n114), .B0(n5468), .B1(n11249), .Y(
        n9988) );
  AO22X2 U9027 ( .A0(mem_rdata_I[18]), .A1(n115), .B0(n5469), .B1(n11248), .Y(
        n10041) );
  AO22X2 U9028 ( .A0(mem_rdata_I[17]), .A1(n113), .B0(n5470), .B1(n11247), .Y(
        n11134) );
  AO22X2 U9029 ( .A0(mem_rdata_I[16]), .A1(n115), .B0(n5469), .B1(n11246), .Y(
        n10070) );
  AO22X2 U9030 ( .A0(mem_rdata_I[14]), .A1(n115), .B0(n5465), .B1(n11244), .Y(
        n9402) );
  AO22X2 U9031 ( .A0(mem_rdata_I[13]), .A1(n115), .B0(n5465), .B1(n11243), .Y(
        n9382) );
  AO22X2 U9032 ( .A0(mem_rdata_I[12]), .A1(n115), .B0(n5469), .B1(n11242), .Y(
        n10095) );
  AO22X2 U9033 ( .A0(mem_rdata_I[11]), .A1(n114), .B0(n5468), .B1(n11241), .Y(
        n9964) );
  AO22X2 U9034 ( .A0(mem_rdata_I[9]), .A1(n115), .B0(n5469), .B1(n11239), .Y(
        n9650) );
  AO22X2 U9035 ( .A0(mem_rdata_I[8]), .A1(n115), .B0(n5468), .B1(n11238), .Y(
        n9426) );
  AO22X2 U9036 ( .A0(mem_rdata_I[6]), .A1(n113), .B0(n5468), .B1(n11236), .Y(
        n9441) );
  AO22X2 U9037 ( .A0(mem_rdata_I[5]), .A1(n115), .B0(n5465), .B1(n11235), .Y(
        n9546) );
  AO22X2 U9038 ( .A0(mem_rdata_I[4]), .A1(n115), .B0(n5468), .B1(n11234), .Y(
        n9463) );
  AO22X2 U9039 ( .A0(mem_rdata_I[2]), .A1(n114), .B0(n5465), .B1(n11232), .Y(
        n9482) );
  AO22X2 U9040 ( .A0(mem_rdata_I[1]), .A1(n113), .B0(n5469), .B1(n11231), .Y(
        n9361) );
  AO22X2 U9041 ( .A0(mem_rdata_I[63]), .A1(n113), .B0(n5471), .B1(n11293), .Y(
        n11038) );
  AO22X2 U9042 ( .A0(mem_rdata_I[61]), .A1(n115), .B0(n5470), .B1(n11291), .Y(
        n11163) );
  AO22X2 U9043 ( .A0(mem_rdata_I[58]), .A1(n113), .B0(n5469), .B1(n11288), .Y(
        n9711) );
  AO22X2 U9044 ( .A0(mem_rdata_I[57]), .A1(n113), .B0(n5466), .B1(n11287), .Y(
        n10124) );
  AO22X2 U9045 ( .A0(mem_rdata_I[56]), .A1(n113), .B0(n5467), .B1(n11286), .Y(
        n9902) );
  AO22X2 U9046 ( .A0(mem_rdata_I[55]), .A1(n113), .B0(n5467), .B1(n11285), .Y(
        n9926) );
  AO22X2 U9047 ( .A0(mem_rdata_I[53]), .A1(n113), .B0(n5467), .B1(n11283), .Y(
        n9878) );
  AO22X2 U9048 ( .A0(mem_rdata_I[52]), .A1(n113), .B0(n5468), .B1(n11282), .Y(
        n10022) );
  AO22X2 U9049 ( .A0(mem_rdata_I[51]), .A1(n113), .B0(n5468), .B1(n11281), .Y(
        n9993) );
  AO22X2 U9050 ( .A0(mem_rdata_I[50]), .A1(n113), .B0(n5469), .B1(n11280), .Y(
        n10046) );
  AO22X2 U9051 ( .A0(mem_rdata_I[49]), .A1(n113), .B0(n5470), .B1(n11279), .Y(
        n11145) );
  AO22X2 U9052 ( .A0(mem_rdata_I[48]), .A1(n115), .B0(n5469), .B1(n11278), .Y(
        n10075) );
  AO22X2 U9053 ( .A0(mem_rdata_I[46]), .A1(n114), .B0(n5465), .B1(n11276), .Y(
        n9407) );
  AO22X2 U9054 ( .A0(mem_rdata_I[45]), .A1(n114), .B0(n5465), .B1(n11275), .Y(
        n9387) );
  AO22X2 U9055 ( .A0(mem_rdata_I[44]), .A1(n113), .B0(n5469), .B1(n11274), .Y(
        n10100) );
  AO22X2 U9056 ( .A0(mem_rdata_I[43]), .A1(n115), .B0(n5468), .B1(n11273), .Y(
        n9969) );
  AO22X2 U9057 ( .A0(mem_rdata_I[42]), .A1(n113), .B0(n5469), .B1(n11272), .Y(
        n9673) );
  AO22X2 U9058 ( .A0(mem_rdata_I[41]), .A1(n113), .B0(n5469), .B1(n11271), .Y(
        n9640) );
  AO22X2 U9059 ( .A0(mem_rdata_I[40]), .A1(n115), .B0(n5468), .B1(n11270), .Y(
        n9416) );
  AO22X2 U9060 ( .A0(mem_rdata_I[39]), .A1(n114), .B0(n5466), .B1(n11269), .Y(
        n9820) );
  AO22X2 U9061 ( .A0(mem_rdata_I[38]), .A1(n113), .B0(n5468), .B1(n11268), .Y(
        n9450) );
  AO22X2 U9062 ( .A0(mem_rdata_I[36]), .A1(n113), .B0(n5468), .B1(n11266), .Y(
        n9472) );
  AO22X2 U9063 ( .A0(mem_rdata_I[34]), .A1(n115), .B0(n5465), .B1(n11264), .Y(
        n9492) );
  AO22X2 U9064 ( .A0(mem_rdata_I[33]), .A1(n114), .B0(n5470), .B1(n11263), .Y(
        n10999) );
  AO22X2 U9065 ( .A0(mem_rdata_I[95]), .A1(n113), .B0(n5468), .B1(n11325), .Y(
        n11036) );
  AO22X2 U9066 ( .A0(mem_rdata_I[93]), .A1(n115), .B0(n5470), .B1(n11323), .Y(
        n11159) );
  AO22X2 U9067 ( .A0(mem_rdata_I[92]), .A1(n114), .B0(n5467), .B1(n11322), .Y(
        n9769) );
  AO22X2 U9068 ( .A0(mem_rdata_I[91]), .A1(n113), .B0(n5467), .B1(n11321), .Y(
        n9725) );
  AO22X2 U9069 ( .A0(mem_rdata_I[90]), .A1(n114), .B0(n5465), .B1(n11320), .Y(
        n9701) );
  AO22X2 U9070 ( .A0(mem_rdata_I[89]), .A1(n115), .B0(n5470), .B1(n11319), .Y(
        n10114) );
  AO22X2 U9071 ( .A0(mem_rdata_I[88]), .A1(n113), .B0(n5467), .B1(n11318), .Y(
        n9892) );
  AO22X2 U9072 ( .A0(mem_rdata_I[87]), .A1(n115), .B0(n5467), .B1(n11317), .Y(
        n9916) );
  AO22X2 U9073 ( .A0(mem_rdata_I[85]), .A1(n114), .B0(n5467), .B1(n11315), .Y(
        n9868) );
  AO22X2 U9074 ( .A0(mem_rdata_I[84]), .A1(n114), .B0(n5468), .B1(n11314), .Y(
        n10012) );
  AO22X2 U9075 ( .A0(mem_rdata_I[83]), .A1(n114), .B0(n5468), .B1(n11313), .Y(
        n9983) );
  AO22X2 U9076 ( .A0(mem_rdata_I[82]), .A1(n114), .B0(n5469), .B1(n11312), .Y(
        n10036) );
  AO22X2 U9077 ( .A0(mem_rdata_I[81]), .A1(n114), .B0(n5470), .B1(n11311), .Y(
        n11129) );
  AO22X2 U9078 ( .A0(mem_rdata_I[80]), .A1(n114), .B0(n5469), .B1(n11310), .Y(
        n10065) );
  AO22X2 U9079 ( .A0(mem_rdata_I[78]), .A1(n114), .B0(n5468), .B1(n11308), .Y(
        n9397) );
  AO22X2 U9080 ( .A0(mem_rdata_I[77]), .A1(n115), .B0(n5468), .B1(n11307), .Y(
        n9377) );
  AO22X2 U9081 ( .A0(mem_rdata_I[76]), .A1(n113), .B0(n5469), .B1(n11306), .Y(
        n10090) );
  AO22X2 U9082 ( .A0(mem_rdata_I[74]), .A1(n114), .B0(n5466), .B1(n11304), .Y(
        n9664) );
  AO22X2 U9083 ( .A0(mem_rdata_I[72]), .A1(n114), .B0(n5465), .B1(n11302), .Y(
        n9412) );
  AO22X2 U9084 ( .A0(mem_rdata_I[70]), .A1(n113), .B0(n5468), .B1(n11300), .Y(
        n9446) );
  AO22X2 U9085 ( .A0(mem_rdata_I[68]), .A1(n115), .B0(n5468), .B1(n11298), .Y(
        n9468) );
  AO22X2 U9086 ( .A0(mem_rdata_I[66]), .A1(n114), .B0(n5465), .B1(n11296), .Y(
        n9487) );
  AO22X2 U9087 ( .A0(mem_rdata_I[65]), .A1(n115), .B0(n5466), .B1(n11295), .Y(
        n10998) );
  AO22X2 U9088 ( .A0(mem_rdata_I[127]), .A1(n115), .B0(n5469), .B1(n11357), 
        .Y(n11035) );
  AO22X2 U9089 ( .A0(mem_rdata_I[125]), .A1(n114), .B0(n5470), .B1(n11355), 
        .Y(n11158) );
  AO22X2 U9090 ( .A0(mem_rdata_I[124]), .A1(n113), .B0(n5467), .B1(n11354), 
        .Y(n9764) );
  AO22X2 U9091 ( .A0(mem_rdata_I[123]), .A1(n115), .B0(n5467), .B1(n11353), 
        .Y(n9720) );
  AO22X2 U9092 ( .A0(mem_rdata_I[121]), .A1(n114), .B0(n5469), .B1(n11351), 
        .Y(n10109) );
  AO22X2 U9093 ( .A0(mem_rdata_I[120]), .A1(n114), .B0(n5467), .B1(n11350), 
        .Y(n9887) );
  AO22X2 U9094 ( .A0(mem_rdata_I[119]), .A1(n114), .B0(n5467), .B1(n11349), 
        .Y(n9911) );
  AO22X2 U9095 ( .A0(mem_rdata_I[115]), .A1(n114), .B0(n5468), .B1(n11345), 
        .Y(n9978) );
  AO22X2 U9096 ( .A0(mem_rdata_I[114]), .A1(n113), .B0(n5468), .B1(n11344), 
        .Y(n10031) );
  AO22X2 U9097 ( .A0(mem_rdata_I[113]), .A1(n114), .B0(n5470), .B1(n11343), 
        .Y(n11124) );
  AO22X2 U9098 ( .A0(mem_rdata_I[110]), .A1(n113), .B0(n5466), .B1(n11340), 
        .Y(n9392) );
  AO22X2 U9099 ( .A0(mem_rdata_I[109]), .A1(n115), .B0(n5468), .B1(n11339), 
        .Y(n9372) );
  AO22X2 U9100 ( .A0(mem_rdata_I[108]), .A1(n114), .B0(n5469), .B1(n11338), 
        .Y(n10085) );
  AO22X2 U9101 ( .A0(mem_rdata_I[107]), .A1(n114), .B0(n5467), .B1(n11337), 
        .Y(n9954) );
  AO22X2 U9102 ( .A0(mem_rdata_I[106]), .A1(n113), .B0(n5469), .B1(n11336), 
        .Y(n9659) );
  AO22X2 U9103 ( .A0(mem_rdata_I[105]), .A1(n115), .B0(n5469), .B1(n11335), 
        .Y(n9645) );
  AO22X2 U9104 ( .A0(mem_rdata_I[104]), .A1(n114), .B0(n5468), .B1(n11334), 
        .Y(n9421) );
  AO22X2 U9105 ( .A0(mem_rdata_I[103]), .A1(n115), .B0(n5466), .B1(n11333), 
        .Y(n9825) );
  AO22X2 U9106 ( .A0(mem_rdata_I[102]), .A1(n113), .B0(n5468), .B1(n11332), 
        .Y(n9436) );
  AO22X2 U9107 ( .A0(mem_rdata_I[101]), .A1(n113), .B0(n5469), .B1(n11331), 
        .Y(n9541) );
  AO22X2 U9108 ( .A0(mem_rdata_I[100]), .A1(n114), .B0(n5468), .B1(n11330), 
        .Y(n9458) );
  AO22X2 U9109 ( .A0(mem_rdata_I[98]), .A1(n115), .B0(n5468), .B1(n11328), .Y(
        n9477) );
  AO22X2 U9110 ( .A0(mem_rdata_I[97]), .A1(n115), .B0(n5467), .B1(n11327), .Y(
        n9356) );
  AO22X2 U9111 ( .A0(n113), .A1(ICACHE_addr[24]), .B0(n5463), .B1(n3589), .Y(
        n10984) );
  AO22X2 U9112 ( .A0(n114), .A1(n3645), .B0(n5463), .B1(n11366), .Y(n10993) );
  AO22X2 U9113 ( .A0(n114), .A1(ICACHE_addr[26]), .B0(n5463), .B1(n11385), .Y(
        n10985) );
  AO22X2 U9114 ( .A0(n113), .A1(ICACHE_addr[20]), .B0(n5463), .B1(n11379), .Y(
        n10996) );
  AO22X2 U9115 ( .A0(mem_rdata_I[35]), .A1(n113), .B0(n5465), .B1(n11265), .Y(
        n9527) );
  AO22X2 U9116 ( .A0(mem_rdata_I[67]), .A1(n113), .B0(n5465), .B1(n11297), .Y(
        n9522) );
  AO22X2 U9117 ( .A0(mem_rdata_I[15]), .A1(n115), .B0(n5466), .B1(n11245), .Y(
        n11007) );
  AO22X2 U9118 ( .A0(mem_rdata_I[47]), .A1(n114), .B0(n5466), .B1(n11277), .Y(
        n11009) );
  AO22X2 U9119 ( .A0(mem_rdata_I[79]), .A1(n113), .B0(n5471), .B1(n11309), .Y(
        n11008) );
  AO22X2 U9120 ( .A0(mem_rdata_I[99]), .A1(n115), .B0(n5465), .B1(n11329), .Y(
        n9512) );
  AO22X2 U9121 ( .A0(n5064), .A1(n12949), .B0(n5061), .B1(n11531), .Y(n10682)
         );
  CLKBUFX2 U9122 ( .A(n4576), .Y(n5064) );
  AO22X2 U9123 ( .A0(n113), .A1(ICACHE_addr[29]), .B0(n5463), .B1(n3565), .Y(
        n10977) );
  AO22X2 U9124 ( .A0(n114), .A1(ICACHE_addr[11]), .B0(n5463), .B1(n11370), .Y(
        n10987) );
  AO22X2 U9125 ( .A0(n115), .A1(ICACHE_addr[10]), .B0(n5463), .B1(n11369), .Y(
        n10988) );
  OAI221XL U9126 ( .A0(\i_MIPS/Register/register[2][27] ), .A1(n4923), .B0(
        \i_MIPS/Register/register[10][27] ), .B1(n4917), .C0(n8624), .Y(n8627)
         );
  OAI221XL U9127 ( .A0(\i_MIPS/Register/register[2][20] ), .A1(n4923), .B0(
        \i_MIPS/Register/register[10][20] ), .B1(n4917), .C0(n8565), .Y(n8568)
         );
  OAI221XL U9128 ( .A0(\i_MIPS/Register/register[2][25] ), .A1(n4923), .B0(
        \i_MIPS/Register/register[10][25] ), .B1(n4915), .C0(n8460), .Y(n8463)
         );
  OA22X1 U9129 ( .A0(\i_MIPS/Register/register[6][25] ), .A1(n4913), .B0(
        \i_MIPS/Register/register[14][25] ), .B1(n4907), .Y(n8460) );
  OAI221XL U9130 ( .A0(\i_MIPS/Register/register[2][21] ), .A1(n4922), .B0(
        \i_MIPS/Register/register[10][21] ), .B1(n4915), .C0(n8051), .Y(n8054)
         );
  OAI221XL U9131 ( .A0(\i_MIPS/Register/register[2][23] ), .A1(n4923), .B0(
        \i_MIPS/Register/register[10][23] ), .B1(n4917), .C0(n8233), .Y(n8236)
         );
  OAI221XL U9132 ( .A0(\i_MIPS/Register/register[2][22] ), .A1(n4922), .B0(
        \i_MIPS/Register/register[10][22] ), .B1(n4917), .C0(n7992), .Y(n7995)
         );
  OA22X1 U9133 ( .A0(\i_MIPS/Register/register[6][22] ), .A1(n4912), .B0(
        \i_MIPS/Register/register[14][22] ), .B1(n4906), .Y(n7992) );
  OAI221XL U9134 ( .A0(\i_MIPS/Register/register[2][16] ), .A1(n4923), .B0(
        \i_MIPS/Register/register[10][16] ), .B1(n4917), .C0(n8175), .Y(n8178)
         );
  OAI221XL U9135 ( .A0(\i_MIPS/Register/register[2][28] ), .A1(n4921), .B0(
        \i_MIPS/Register/register[10][28] ), .B1(n4917), .C0(n9028), .Y(n9031)
         );
  OAI221XL U9136 ( .A0(\i_MIPS/Register/register[2][24] ), .A1(n4921), .B0(
        \i_MIPS/Register/register[10][24] ), .B1(n4917), .C0(n8940), .Y(n8943)
         );
  OAI221XL U9137 ( .A0(\i_MIPS/Register/register[2][2] ), .A1(n4921), .B0(
        \i_MIPS/Register/register[10][2] ), .B1(n4917), .C0(n8831), .Y(n8834)
         );
  OA22X1 U9138 ( .A0(\i_MIPS/Register/register[6][2] ), .A1(n4914), .B0(
        \i_MIPS/Register/register[14][2] ), .B1(n4908), .Y(n8831) );
  OAI221XL U9139 ( .A0(\i_MIPS/Register/register[2][18] ), .A1(n4922), .B0(
        \i_MIPS/Register/register[10][18] ), .B1(n4916), .C0(n7896), .Y(n7899)
         );
  OA22X1 U9140 ( .A0(\i_MIPS/Register/register[6][18] ), .A1(n4912), .B0(
        \i_MIPS/Register/register[14][18] ), .B1(n4906), .Y(n7896) );
  OAI221XL U9141 ( .A0(\i_MIPS/Register/register[2][17] ), .A1(n4922), .B0(
        \i_MIPS/Register/register[10][17] ), .B1(n4916), .C0(n7740), .Y(n7743)
         );
  OAI221XL U9142 ( .A0(\i_MIPS/Register/register[2][10] ), .A1(n4921), .B0(
        \i_MIPS/Register/register[10][10] ), .B1(n4916), .C0(n7215), .Y(n7218)
         );
  OA22X1 U9143 ( .A0(\i_MIPS/Register/register[6][10] ), .A1(n4911), .B0(
        \i_MIPS/Register/register[14][10] ), .B1(n4903), .Y(n7215) );
  OAI221XL U9144 ( .A0(\i_MIPS/Register/register[2][11] ), .A1(n4921), .B0(
        \i_MIPS/Register/register[10][11] ), .B1(n4916), .C0(n7125), .Y(n7128)
         );
  OAI221XL U9145 ( .A0(\i_MIPS/Register/register[2][4] ), .A1(n4921), .B0(
        \i_MIPS/Register/register[10][4] ), .B1(n4916), .C0(n7377), .Y(n7380)
         );
  OAI221XL U9146 ( .A0(\i_MIPS/Register/register[2][5] ), .A1(n4921), .B0(
        \i_MIPS/Register/register[10][5] ), .B1(n4916), .C0(n7298), .Y(n7301)
         );
  OAI221XL U9147 ( .A0(\i_MIPS/Register/register[2][7] ), .A1(n4921), .B0(
        \i_MIPS/Register/register[10][7] ), .B1(n4916), .C0(n7506), .Y(n7509)
         );
  OAI221XL U9148 ( .A0(\i_MIPS/Register/register[2][6] ), .A1(n4922), .B0(
        \i_MIPS/Register/register[10][6] ), .B1(n4916), .C0(n7573), .Y(n7576)
         );
  OA22X1 U9149 ( .A0(\i_MIPS/Register/register[6][13] ), .A1(n4909), .B0(
        \i_MIPS/Register/register[14][13] ), .B1(n4906), .Y(n6399) );
  OAI221XL U9150 ( .A0(\i_MIPS/Register/register[2][12] ), .A1(n4920), .B0(
        \i_MIPS/Register/register[10][12] ), .B1(n4915), .C0(n6309), .Y(n6312)
         );
  OAI221XL U9151 ( .A0(\i_MIPS/Register/register[2][15] ), .A1(n4921), .B0(
        \i_MIPS/Register/register[10][15] ), .B1(n4916), .C0(n7073), .Y(n7076)
         );
  OA22X1 U9152 ( .A0(\i_MIPS/Register/register[6][14] ), .A1(n4909), .B0(
        \i_MIPS/Register/register[14][14] ), .B1(n4906), .Y(n6982) );
  OAI221XL U9153 ( .A0(\i_MIPS/Register/register[18][0] ), .A1(n4920), .B0(
        \i_MIPS/Register/register[26][0] ), .B1(n4915), .C0(n6558), .Y(n6561)
         );
  OA22X1 U9154 ( .A0(\i_MIPS/Register/register[22][0] ), .A1(n4909), .B0(
        \i_MIPS/Register/register[30][0] ), .B1(n4906), .Y(n6558) );
  OAI221XL U9155 ( .A0(\i_MIPS/Register/register[2][0] ), .A1(n4920), .B0(
        \i_MIPS/Register/register[10][0] ), .B1(n4915), .C0(n6549), .Y(n6552)
         );
  OA22X1 U9156 ( .A0(\i_MIPS/Register/register[6][0] ), .A1(n4909), .B0(
        \i_MIPS/Register/register[14][0] ), .B1(n4903), .Y(n6549) );
  OA22X1 U9157 ( .A0(\i_MIPS/Register/register[6][0] ), .A1(n4935), .B0(
        \i_MIPS/Register/register[14][0] ), .B1(n4929), .Y(n6503) );
  INVX1 U9158 ( .A(n9129), .Y(n9131) );
  CLKINVX1 U9159 ( .A(\i_MIPS/n251 ), .Y(n10508) );
  INVX12 U9160 ( .A(n1812), .Y(mem_addr_D[26]) );
  INVX12 U9161 ( .A(n4789), .Y(mem_addr_D[28]) );
  CLKINVX1 U9162 ( .A(n4769), .Y(n4789) );
  INVX12 U9163 ( .A(n1810), .Y(mem_addr_D[24]) );
  INVX12 U9164 ( .A(n4787), .Y(mem_addr_D[22]) );
  INVX1 U9165 ( .A(n4767), .Y(n4787) );
  OAI2BB2XL U9166 ( .B0(net113725), .B1(n4788), .A0N(DCACHE_addr[20]), .A1N(
        mem_read_D), .Y(n4767) );
  CLKINVX1 U9167 ( .A(n11532), .Y(n4788) );
  NAND2X1 U9168 ( .A(n12945), .B(net113089), .Y(net99603) );
  NAND2XL U9169 ( .A(n3768), .B(\i_MIPS/ID_EX[78] ), .Y(n6221) );
  NOR4X1 U9170 ( .A(n9109), .B(n9108), .C(n9107), .D(n9106), .Y(n9124) );
  OAI221XL U9171 ( .A0(\i_MIPS/Register/register[2][31] ), .A1(n4921), .B0(
        \i_MIPS/Register/register[10][31] ), .B1(n4915), .C0(n9105), .Y(n9108)
         );
  NAND4X1 U9172 ( .A(n9104), .B(n9103), .C(n9102), .D(n9101), .Y(n9109) );
  NOR4X1 U9173 ( .A(n9122), .B(n9121), .C(n9120), .D(n9119), .Y(n9123) );
  OAI221XL U9174 ( .A0(\i_MIPS/Register/register[18][31] ), .A1(n4921), .B0(
        \i_MIPS/Register/register[26][31] ), .B1(n4915), .C0(n9114), .Y(n9121)
         );
  NAND4X1 U9175 ( .A(n9113), .B(n9112), .C(n9111), .D(n9110), .Y(n9122) );
  NOR4X1 U9176 ( .A(n7311), .B(n7310), .C(n7309), .D(n7308), .Y(n7312) );
  OAI221XL U9177 ( .A0(\i_MIPS/Register/register[18][5] ), .A1(n4921), .B0(
        \i_MIPS/Register/register[26][5] ), .B1(n4916), .C0(n7307), .Y(n7310)
         );
  NAND4X1 U9178 ( .A(n7306), .B(n7305), .C(n7304), .D(n7303), .Y(n7311) );
  AO22X1 U9179 ( .A0(n4896), .A1(n670), .B0(n4892), .B1(n2199), .Y(n7309) );
  NOR4X1 U9180 ( .A(n7519), .B(n7518), .C(n7517), .D(n7516), .Y(n7520) );
  OAI221XL U9181 ( .A0(\i_MIPS/Register/register[18][7] ), .A1(n4921), .B0(
        \i_MIPS/Register/register[26][7] ), .B1(n4916), .C0(n7515), .Y(n7518)
         );
  NAND4X1 U9182 ( .A(n7514), .B(n7513), .C(n7512), .D(n7511), .Y(n7519) );
  AO22X1 U9183 ( .A0(n4897), .A1(n671), .B0(n4894), .B1(n2200), .Y(n7517) );
  NOR4X1 U9184 ( .A(n7086), .B(n7085), .C(n7084), .D(n7083), .Y(n7087) );
  OAI221XL U9185 ( .A0(\i_MIPS/Register/register[18][15] ), .A1(n4921), .B0(
        \i_MIPS/Register/register[26][15] ), .B1(n4916), .C0(n7082), .Y(n7085)
         );
  NAND4X1 U9186 ( .A(n7081), .B(n7080), .C(n7079), .D(n7078), .Y(n7086) );
  AO22X1 U9187 ( .A0(n4896), .A1(n672), .B0(n4892), .B1(n2201), .Y(n7084) );
  NOR4X1 U9188 ( .A(n6995), .B(n6994), .C(n6993), .D(n6992), .Y(n6996) );
  OAI221XL U9189 ( .A0(\i_MIPS/Register/register[18][14] ), .A1(n4921), .B0(
        \i_MIPS/Register/register[26][14] ), .B1(n4916), .C0(n6991), .Y(n6994)
         );
  NAND4X1 U9190 ( .A(n6990), .B(n6989), .C(n6988), .D(n6987), .Y(n6995) );
  AO22X1 U9191 ( .A0(n4896), .A1(n673), .B0(n4892), .B1(n2202), .Y(n6993) );
  NOR4X1 U9192 ( .A(n7586), .B(n7585), .C(n7584), .D(n7583), .Y(n7587) );
  OAI221XL U9193 ( .A0(\i_MIPS/Register/register[18][6] ), .A1(n4922), .B0(
        \i_MIPS/Register/register[26][6] ), .B1(n4915), .C0(n7582), .Y(n7585)
         );
  NAND4X1 U9194 ( .A(n7581), .B(n7580), .C(n7579), .D(n7578), .Y(n7586) );
  AO22X1 U9195 ( .A0(n4897), .A1(n674), .B0(n4891), .B1(n2203), .Y(n7584) );
  NOR4X1 U9196 ( .A(n6412), .B(n6411), .C(n6410), .D(n6409), .Y(n6413) );
  NAND4X1 U9197 ( .A(n6407), .B(n6406), .C(n6405), .D(n6404), .Y(n6412) );
  AO22X1 U9198 ( .A0(n4895), .A1(n598), .B0(n4891), .B1(n2118), .Y(n6410) );
  NOR4X1 U9199 ( .A(n6903), .B(n6902), .C(n6901), .D(n6900), .Y(n6904) );
  NAND4X1 U9200 ( .A(n6898), .B(n6897), .C(n6896), .D(n6895), .Y(n6903) );
  AO22X1 U9201 ( .A0(n4895), .A1(n675), .B0(n4891), .B1(n2204), .Y(n6901) );
  NAND4X1 U9202 ( .A(n6815), .B(n6814), .C(n6813), .D(n6812), .Y(n6820) );
  AO22X1 U9203 ( .A0(n4895), .A1(n676), .B0(n4891), .B1(n2205), .Y(n6818) );
  NOR4X1 U9204 ( .A(n6322), .B(n6321), .C(n6320), .D(n6319), .Y(n6323) );
  OAI221XL U9205 ( .A0(\i_MIPS/Register/register[18][12] ), .A1(n4920), .B0(
        \i_MIPS/Register/register[26][12] ), .B1(n4915), .C0(n6318), .Y(n6321)
         );
  NAND4X1 U9206 ( .A(n6317), .B(n6316), .C(n6315), .D(n6314), .Y(n6322) );
  AO22X1 U9207 ( .A0(n4895), .A1(n677), .B0(n4891), .B1(n2206), .Y(n6320) );
  OAI221XL U9208 ( .A0(\i_MIPS/Register/register[18][24] ), .A1(n4921), .B0(
        \i_MIPS/Register/register[26][24] ), .B1(n4917), .C0(n8949), .Y(n8952)
         );
  AO22X1 U9209 ( .A0(n4898), .A1(n599), .B0(n4894), .B1(n2119), .Y(n8951) );
  NOR4X1 U9210 ( .A(n8188), .B(n8187), .C(n8186), .D(n8185), .Y(n8189) );
  OAI221XL U9211 ( .A0(\i_MIPS/Register/register[18][16] ), .A1(n4923), .B0(
        \i_MIPS/Register/register[26][16] ), .B1(n4915), .C0(n8184), .Y(n8187)
         );
  NAND4X1 U9212 ( .A(n8183), .B(n8182), .C(n8181), .D(n8180), .Y(n8188) );
  OAI221XL U9213 ( .A0(\i_MIPS/Register/register[18][23] ), .A1(n4923), .B0(
        \i_MIPS/Register/register[26][23] ), .B1(n4917), .C0(n8242), .Y(n8245)
         );
  NAND4X1 U9214 ( .A(n8241), .B(n8240), .C(n8239), .D(n8238), .Y(n8246) );
  NOR4X1 U9215 ( .A(n8005), .B(n8004), .C(n8003), .D(n8002), .Y(n8006) );
  OAI221XL U9216 ( .A0(\i_MIPS/Register/register[18][22] ), .A1(n4922), .B0(
        \i_MIPS/Register/register[26][22] ), .B1(n4917), .C0(n8001), .Y(n8004)
         );
  NAND4X1 U9217 ( .A(n8000), .B(n7999), .C(n7998), .D(n7997), .Y(n8005) );
  AO22X1 U9218 ( .A0(n4897), .A1(n600), .B0(n4894), .B1(n2120), .Y(n8003) );
  NOR4X1 U9219 ( .A(n8759), .B(n8758), .C(n8757), .D(n8756), .Y(n8760) );
  NAND4X1 U9220 ( .A(n8754), .B(n8753), .C(n8752), .D(n8751), .Y(n8759) );
  AO22X1 U9221 ( .A0(n4898), .A1(n601), .B0(n4894), .B1(n2121), .Y(n8757) );
  NOR4X1 U9222 ( .A(n8578), .B(n8577), .C(n8576), .D(n8575), .Y(n8579) );
  OAI221XL U9223 ( .A0(\i_MIPS/Register/register[18][20] ), .A1(n4923), .B0(
        \i_MIPS/Register/register[26][20] ), .B1(n4917), .C0(n8574), .Y(n8577)
         );
  NAND4X1 U9224 ( .A(n8573), .B(n8572), .C(n8571), .D(n8570), .Y(n8578) );
  AO22X1 U9225 ( .A0(n4898), .A1(n602), .B0(n4893), .B1(n2122), .Y(n8576) );
  NOR4X1 U9226 ( .A(n8064), .B(n8063), .C(n8062), .D(n8061), .Y(n8065) );
  OAI221XL U9227 ( .A0(\i_MIPS/Register/register[18][21] ), .A1(n4923), .B0(
        \i_MIPS/Register/register[26][21] ), .B1(n4917), .C0(n8060), .Y(n8063)
         );
  NAND4X1 U9228 ( .A(n8059), .B(n8058), .C(n8057), .D(n8056), .Y(n8064) );
  AO22X1 U9229 ( .A0(n4897), .A1(n603), .B0(n4894), .B1(n2123), .Y(n8062) );
  NOR4X1 U9230 ( .A(n8844), .B(n8843), .C(n8842), .D(n8841), .Y(n8845) );
  OAI221XL U9231 ( .A0(\i_MIPS/Register/register[18][2] ), .A1(n4921), .B0(
        \i_MIPS/Register/register[26][2] ), .B1(n4917), .C0(n8840), .Y(n8843)
         );
  NAND4X1 U9232 ( .A(n8839), .B(n8838), .C(n8837), .D(n8836), .Y(n8844) );
  AO22X1 U9233 ( .A0(n4898), .A1(n604), .B0(n4894), .B1(n2124), .Y(n8842) );
  NOR4X1 U9234 ( .A(n7390), .B(n7389), .C(n7388), .D(n7387), .Y(n7391) );
  OAI221XL U9235 ( .A0(\i_MIPS/Register/register[18][4] ), .A1(n4921), .B0(
        \i_MIPS/Register/register[26][4] ), .B1(n4916), .C0(n7386), .Y(n7389)
         );
  NAND4X1 U9236 ( .A(n7385), .B(n7384), .C(n7383), .D(n7382), .Y(n7390) );
  AO22X1 U9237 ( .A0(n4896), .A1(n605), .B0(n4892), .B1(n2125), .Y(n7388) );
  NOR4X1 U9238 ( .A(n7228), .B(n7227), .C(n7226), .D(n7225), .Y(n7229) );
  OAI221XL U9239 ( .A0(\i_MIPS/Register/register[18][10] ), .A1(n4921), .B0(
        \i_MIPS/Register/register[26][10] ), .B1(n4916), .C0(n7224), .Y(n7227)
         );
  NAND4X1 U9240 ( .A(n7223), .B(n7222), .C(n7221), .D(n7220), .Y(n7228) );
  AO22X1 U9241 ( .A0(n4896), .A1(n678), .B0(n4892), .B1(n2207), .Y(n7226) );
  NOR4X1 U9242 ( .A(n9041), .B(n9040), .C(n9039), .D(n9038), .Y(n9042) );
  NAND4X1 U9243 ( .A(n9036), .B(n9035), .C(n9034), .D(n9033), .Y(n9041) );
  AO22X1 U9244 ( .A0(n4896), .A1(n606), .B0(n4894), .B1(n2126), .Y(n9039) );
  NOR4X1 U9245 ( .A(n8473), .B(n8472), .C(n8471), .D(n8470), .Y(n8474) );
  OAI221XL U9246 ( .A0(\i_MIPS/Register/register[18][25] ), .A1(n4923), .B0(
        \i_MIPS/Register/register[26][25] ), .B1(n4917), .C0(n8469), .Y(n8472)
         );
  NAND4X1 U9247 ( .A(n8468), .B(n8467), .C(n8466), .D(n8465), .Y(n8473) );
  NOR4X1 U9248 ( .A(n7138), .B(n7137), .C(n7136), .D(n7135), .Y(n7139) );
  OAI221XL U9249 ( .A0(\i_MIPS/Register/register[18][11] ), .A1(n4921), .B0(
        \i_MIPS/Register/register[26][11] ), .B1(n4916), .C0(n7134), .Y(n7137)
         );
  NAND4X1 U9250 ( .A(n7133), .B(n7132), .C(n7131), .D(n7130), .Y(n7138) );
  AO22X1 U9251 ( .A0(n4896), .A1(n607), .B0(n4892), .B1(n2127), .Y(n7136) );
  NOR4X1 U9252 ( .A(n8637), .B(n8636), .C(n8635), .D(n8634), .Y(n8638) );
  OAI221XL U9253 ( .A0(\i_MIPS/Register/register[18][27] ), .A1(n4923), .B0(
        \i_MIPS/Register/register[26][27] ), .B1(n4917), .C0(n8633), .Y(n8636)
         );
  NAND4X1 U9254 ( .A(n8632), .B(n8631), .C(n8630), .D(n8629), .Y(n8637) );
  AO22X1 U9255 ( .A0(n4898), .A1(n608), .B0(n4893), .B1(n2128), .Y(n8635) );
  NOR4X1 U9256 ( .A(n7753), .B(n7752), .C(n7751), .D(n7750), .Y(n7754) );
  OAI221XL U9257 ( .A0(\i_MIPS/Register/register[18][17] ), .A1(n4922), .B0(
        \i_MIPS/Register/register[26][17] ), .B1(n4915), .C0(n7749), .Y(n7752)
         );
  NAND4X1 U9258 ( .A(n7748), .B(n7747), .C(n7746), .D(n7745), .Y(n7753) );
  AO22X1 U9259 ( .A0(n4897), .A1(n679), .B0(n4894), .B1(n2208), .Y(n7751) );
  AO22X1 U9260 ( .A0(n4897), .A1(n680), .B0(n4891), .B1(n2209), .Y(n7907) );
  CLKINVX1 U9261 ( .A(n11184), .Y(n11191) );
  OAI221XL U9262 ( .A0(\i_MIPS/Register/register[18][25] ), .A1(n4947), .B0(
        \i_MIPS/Register/register[26][25] ), .B1(n4939), .C0(n8503), .Y(n8511)
         );
  OAI221XL U9263 ( .A0(\i_MIPS/Register/register[2][25] ), .A1(n4947), .B0(
        \i_MIPS/Register/register[10][25] ), .B1(n4939), .C0(n8494), .Y(n8502)
         );
  OAI221XL U9264 ( .A0(\i_MIPS/Register/register[2][1] ), .A1(n4946), .B0(
        \i_MIPS/Register/register[10][1] ), .B1(n4940), .C0(n7590), .Y(n7598)
         );
  OA22X1 U9265 ( .A0(\i_MIPS/Register/register[6][1] ), .A1(n4937), .B0(
        \i_MIPS/Register/register[14][1] ), .B1(n4930), .Y(n7590) );
  NAND4X1 U9266 ( .A(\i_MIPS/IR_ID[29] ), .B(\i_MIPS/IR_ID[31] ), .C(n4717), 
        .D(n9809), .Y(n11200) );
  AND3XL U9267 ( .A(net110227), .B(\i_MIPS/n326 ), .C(\i_MIPS/n330 ), .Y(n9809) );
  XNOR2XL U9268 ( .A(\i_MIPS/IR_ID[16] ), .B(\i_MIPS/Reg_W[0] ), .Y(n6194) );
  XNOR2XL U9269 ( .A(\i_MIPS/IR_ID[17] ), .B(\i_MIPS/Reg_W[1] ), .Y(n6195) );
  XNOR2XL U9270 ( .A(\i_MIPS/IR_ID[18] ), .B(\i_MIPS/Reg_W[2] ), .Y(n6196) );
  XOR2X4 U9271 ( .A(n11388), .B(\i_MIPS/PC/n33 ), .Y(n4651) );
  XOR2X4 U9272 ( .A(n11384), .B(\i_MIPS/PC/n29 ), .Y(n4661) );
  XNOR2XL U9273 ( .A(\i_MIPS/Reg_W[3] ), .B(\i_MIPS/IR_ID[24] ), .Y(n6289) );
  AOI2BB1XL U9274 ( .A0N(\i_MIPS/ALUin1[15] ), .A1N(n3592), .B0(n4597), .Y(
        n7021) );
  XNOR2XL U9275 ( .A(\i_MIPS/Reg_W[1] ), .B(\i_MIPS/IR_ID[22] ), .Y(n6290) );
  XNOR2XL U9276 ( .A(\i_MIPS/Reg_W[2] ), .B(\i_MIPS/IR_ID[23] ), .Y(n6287) );
  XNOR2XL U9277 ( .A(\i_MIPS/Reg_W[0] ), .B(\i_MIPS/IR_ID[21] ), .Y(n6288) );
  XOR2X4 U9278 ( .A(n11378), .B(\i_MIPS/PC/n23 ), .Y(n4662) );
  XNOR2X1 U9279 ( .A(\i_MIPS/Reg_W[4] ), .B(net108959), .Y(n6198) );
  NAND2XL U9280 ( .A(\i_MIPS/ALU/N303 ), .B(n9143), .Y(n9161) );
  XOR2X4 U9281 ( .A(n11367), .B(n3650), .Y(n4663) );
  NAND2XL U9282 ( .A(\i_MIPS/ALU/N303 ), .B(n9142), .Y(n11221) );
  OAI2BB2XL U9283 ( .B0(\i_MIPS/n227 ), .B1(net110225), .A0N(n176), .A1N(n168), 
        .Y(\i_MIPS/N70 ) );
  OAI2BB2XL U9284 ( .B0(\i_MIPS/n226 ), .B1(net110227), .A0N(n173), .A1N(
        n10906), .Y(\i_MIPS/N69 ) );
  OAI2BB2XL U9285 ( .B0(\i_MIPS/n224 ), .B1(net110225), .A0N(n174), .A1N(
        n10295), .Y(\i_MIPS/N67 ) );
  OAI2BB2XL U9286 ( .B0(\i_MIPS/n212 ), .B1(net110221), .A0N(n176), .A1N(
        n11189), .Y(\i_MIPS/N55 ) );
  OAI2BB2XL U9287 ( .B0(\i_MIPS/n232 ), .B1(net110225), .A0N(n173), .A1N(
        n10370), .Y(\i_MIPS/N80 ) );
  OAI2BB2XL U9288 ( .B0(\i_MIPS/n231 ), .B1(net110225), .A0N(n176), .A1N(
        n10356), .Y(\i_MIPS/N79 ) );
  OAI2BB2XL U9289 ( .B0(\i_MIPS/n230 ), .B1(net110225), .A0N(n175), .A1N(
        n10337), .Y(\i_MIPS/N78 ) );
  OAI2BB2XL U9290 ( .B0(\i_MIPS/n229 ), .B1(net110225), .A0N(n174), .A1N(
        net99759), .Y(\i_MIPS/N77 ) );
  OAI2BB2XL U9291 ( .B0(\i_MIPS/n225 ), .B1(net110225), .A0N(n173), .A1N(
        n11093), .Y(\i_MIPS/N68 ) );
  OAI2BB2XL U9292 ( .B0(\i_MIPS/n221 ), .B1(net110221), .A0N(n174), .A1N(
        n11073), .Y(\i_MIPS/N64 ) );
  OAI2BB2XL U9293 ( .B0(\i_MIPS/n219 ), .B1(net110221), .A0N(n175), .A1N(
        n10884), .Y(\i_MIPS/N62 ) );
  OAI2BB2XL U9294 ( .B0(\i_MIPS/n217 ), .B1(net110221), .A0N(n175), .A1N(
        n10212), .Y(\i_MIPS/N60 ) );
  OAI2BB2XL U9295 ( .B0(\i_MIPS/n216 ), .B1(net110227), .A0N(n173), .A1N(
        n11063), .Y(\i_MIPS/N59 ) );
  OAI2BB2XL U9296 ( .B0(\i_MIPS/n214 ), .B1(net110221), .A0N(n175), .A1N(n9678), .Y(\i_MIPS/N57 ) );
  OAI2BB2XL U9297 ( .B0(\i_MIPS/n213 ), .B1(net110221), .A0N(n173), .A1N(
        n11044), .Y(\i_MIPS/N56 ) );
  OAI2BB2XL U9298 ( .B0(\i_MIPS/n182 ), .B1(net110227), .A0N(n174), .A1N(
        \i_MIPS/PC/n4 ), .Y(\i_MIPS/N25 ) );
  INVXL U9299 ( .A(n11052), .Y(n11051) );
  OAI2BB2XL U9300 ( .B0(\i_MIPS/n242 ), .B1(net110221), .A0N(n176), .A1N(
        n10875), .Y(\i_MIPS/N96 ) );
  CLKINVX1 U9301 ( .A(n10876), .Y(n10875) );
  OAI2BB2XL U9302 ( .B0(\i_MIPS/n243 ), .B1(net110221), .A0N(n176), .A1N(
        n10886), .Y(\i_MIPS/N97 ) );
  OAI2BB2XL U9303 ( .B0(\i_MIPS/n245 ), .B1(net110217), .A0N(n175), .A1N(
        n11076), .Y(\i_MIPS/N99 ) );
  OAI2BB2XL U9304 ( .B0(\i_MIPS/n172 ), .B1(net110225), .A0N(n173), .A1N(
        n10335), .Y(\i_MIPS/N113 ) );
  CLKINVX1 U9305 ( .A(n10336), .Y(n10335) );
  OAI2BB2XL U9306 ( .B0(\i_MIPS/n222 ), .B1(net110221), .A0N(n173), .A1N(
        n10273), .Y(\i_MIPS/N65 ) );
  OAI2BB2XL U9307 ( .B0(\i_MIPS/n183 ), .B1(net110217), .A0N(n175), .A1N(
        n11043), .Y(\i_MIPS/N26 ) );
  OAI2BB2XL U9308 ( .B0(\i_MIPS/n236 ), .B1(net110217), .A0N(n174), .A1N(
        n11184), .Y(\i_MIPS/N90 ) );
  OAI2BB2XL U9309 ( .B0(\i_MIPS/n237 ), .B1(net110219), .A0N(n173), .A1N(
        n11000), .Y(\i_MIPS/N91 ) );
  OAI2BB2XL U9310 ( .B0(\i_MIPS/n238 ), .B1(net110215), .A0N(n175), .A1N(
        n11193), .Y(\i_MIPS/N92 ) );
  CLKINVX1 U9311 ( .A(n11194), .Y(n11193) );
  CLKINVX1 U9312 ( .A(n11067), .Y(n11066) );
  OAI2BB2XL U9313 ( .B0(\i_MIPS/n162 ), .B1(net110217), .A0N(n176), .A1N(
        n11096), .Y(\i_MIPS/N103 ) );
  OAI2BB2XL U9314 ( .B0(\i_MIPS/n166 ), .B1(net110217), .A0N(n176), .A1N(
        n11119), .Y(\i_MIPS/N107 ) );
  OAI2BB2XL U9315 ( .B0(\i_MIPS/n199 ), .B1(net110217), .A0N(n11118), .A1N(
        n174), .Y(\i_MIPS/N42 ) );
  OAI2BB2XL U9316 ( .B0(\i_MIPS/n186 ), .B1(net110219), .A0N(n11065), .A1N(
        n173), .Y(\i_MIPS/N29 ) );
  OAI2BB2XL U9317 ( .B0(\i_MIPS/n208 ), .B1(net110227), .A0N(n10500), .A1N(
        n176), .Y(\i_MIPS/N51 ) );
  OAI2BB2XL U9318 ( .B0(\i_MIPS/n209 ), .B1(net110227), .A0N(n10699), .A1N(
        n176), .Y(\i_MIPS/N52 ) );
  OAI2BB2XL U9319 ( .B0(\i_MIPS/n197 ), .B1(net110217), .A0N(n11110), .A1N(
        n173), .Y(\i_MIPS/N40 ) );
  OAI2BB2XL U9320 ( .B0(\i_MIPS/n201 ), .B1(net110219), .A0N(n11025), .A1N(
        n174), .Y(\i_MIPS/N44 ) );
  OAI2BB2XL U9321 ( .B0(\i_MIPS/n194 ), .B1(net110225), .A0N(n10296), .A1N(
        n175), .Y(\i_MIPS/N37 ) );
  OAI2BB2XL U9322 ( .B0(\i_MIPS/n195 ), .B1(net110217), .A0N(n11095), .A1N(
        n173), .Y(\i_MIPS/N38 ) );
  OAI2BB2XL U9323 ( .B0(\i_MIPS/n204 ), .B1(net110225), .A0N(net99737), .A1N(
        n174), .Y(\i_MIPS/N47 ) );
  OAI2BB2XL U9324 ( .B0(\i_MIPS/n210 ), .B1(net110227), .A0N(n10713), .A1N(
        n176), .Y(\i_MIPS/N53 ) );
  OAI2BB2XL U9325 ( .B0(\i_MIPS/n192 ), .B1(net110225), .A0N(n10274), .A1N(
        n175), .Y(\i_MIPS/N35 ) );
  OAI2BB2XL U9326 ( .B0(\i_MIPS/n233 ), .B1(net110221), .A0N(n10865), .A1N(
        n175), .Y(\i_MIPS/N87 ) );
  OAI2BB2XL U9327 ( .B0(\i_MIPS/n211 ), .B1(net110227), .A0N(n10737), .A1N(
        n173), .Y(\i_MIPS/N54 ) );
  INVXL U9328 ( .A(n10736), .Y(n10737) );
  OAI2BB2XL U9329 ( .B0(\i_MIPS/n161 ), .B1(net110225), .A0N(n10284), .A1N(
        n174), .Y(\i_MIPS/N102 ) );
  CLKINVX1 U9330 ( .A(n10285), .Y(n10284) );
  OAI2BB2XL U9331 ( .B0(\i_MIPS/n180 ), .B1(net110221), .A0N(
        \i_MIPS/BranchAddr[0] ), .A1N(n175), .Y(\i_MIPS/N23 ) );
  OAI2BB2XL U9332 ( .B0(\i_MIPS/n181 ), .B1(net110221), .A0N(\i_MIPS/PC_o[1] ), 
        .A1N(n173), .Y(\i_MIPS/N24 ) );
  OAI2BB2XL U9333 ( .B0(\i_MIPS/n207 ), .B1(net110221), .A0N(n10381), .A1N(
        n174), .Y(\i_MIPS/N50 ) );
  OAI2BB2XL U9334 ( .B0(\i_MIPS/n234 ), .B1(net110227), .A0N(
        \i_MIPS/BranchAddr[0] ), .A1N(n176), .Y(\i_MIPS/N88 ) );
  OAI2BB2XL U9335 ( .B0(\i_MIPS/n235 ), .B1(net110221), .A0N(\i_MIPS/PC_o[1] ), 
        .A1N(n176), .Y(\i_MIPS/N89 ) );
  OAI2BB2XL U9336 ( .B0(\i_MIPS/n179 ), .B1(net110219), .A0N(n11041), .A1N(
        n174), .Y(\i_MIPS/N120 ) );
  AND3XL U9337 ( .A(n11040), .B(n11039), .C(n4511), .Y(n11041) );
  OAI2BB2XL U9338 ( .B0(\i_MIPS/n187 ), .B1(net110219), .A0N(n10207), .A1N(
        n174), .Y(\i_MIPS/N30 ) );
  OAI2BB2XL U9339 ( .B0(\i_MIPS/n198 ), .B1(net110219), .A0N(n10940), .A1N(
        n175), .Y(\i_MIPS/N41 ) );
  OAI2BB2XL U9340 ( .B0(\i_MIPS/n203 ), .B1(net110219), .A0N(n10965), .A1N(
        n175), .Y(\i_MIPS/N46 ) );
  OAI2BB2XL U9341 ( .B0(\i_MIPS/n189 ), .B1(net110219), .A0N(n10885), .A1N(
        n176), .Y(\i_MIPS/N32 ) );
  OAI2BB2XL U9342 ( .B0(\i_MIPS/n196 ), .B1(net110221), .A0N(n10905), .A1N(
        n173), .Y(\i_MIPS/N39 ) );
  OAI2BB2XL U9343 ( .B0(\i_MIPS/n188 ), .B1(net110219), .A0N(n10874), .A1N(
        n176), .Y(\i_MIPS/N31 ) );
  OAI2BB2XL U9344 ( .B0(\i_MIPS/n190 ), .B1(net110219), .A0N(n10897), .A1N(
        n176), .Y(\i_MIPS/N33 ) );
  OAI2BB2XL U9345 ( .B0(\i_MIPS/n200 ), .B1(net110217), .A0N(n10292), .A1N(
        n176), .Y(\i_MIPS/N43 ) );
  OAI2BB2XL U9346 ( .B0(\i_MIPS/n206 ), .B1(net110225), .A0N(n10364), .A1N(
        n175), .Y(\i_MIPS/N49 ) );
  NAND2XL U9347 ( .A(\i_MIPS/ALUin1[30] ), .B(n9268), .Y(n9260) );
  NAND2X1 U9348 ( .A(n11183), .B(n11182), .Y(n11184) );
  NAND4X1 U9349 ( .A(n6981), .B(n6980), .C(n6979), .D(n6978), .Y(n6986) );
  OA22X1 U9350 ( .A0(\i_MIPS/Register/register[5][14] ), .A1(n4848), .B0(
        \i_MIPS/Register/register[13][14] ), .B1(n4844), .Y(n6980) );
  OA22X1 U9351 ( .A0(\i_MIPS/Register/register[7][14] ), .A1(n4881), .B0(
        \i_MIPS/Register/register[15][14] ), .B1(n4873), .Y(n6978) );
  NAND4X1 U9352 ( .A(n7572), .B(n7571), .C(n7570), .D(n7569), .Y(n7577) );
  NAND4X1 U9353 ( .A(n7505), .B(n7504), .C(n7503), .D(n7502), .Y(n7510) );
  NAND4X1 U9354 ( .A(n6889), .B(n6888), .C(n6887), .D(n6886), .Y(n6894) );
  OA22X1 U9355 ( .A0(\i_MIPS/Register/register[5][9] ), .A1(n4848), .B0(
        \i_MIPS/Register/register[13][9] ), .B1(n4843), .Y(n6888) );
  OA22X1 U9356 ( .A0(\i_MIPS/Register/register[7][9] ), .A1(n4881), .B0(
        \i_MIPS/Register/register[15][9] ), .B1(n4873), .Y(n6886) );
  NAND4X1 U9357 ( .A(n6398), .B(n6397), .C(n6396), .D(n6395), .Y(n6403) );
  OA22X1 U9358 ( .A0(\i_MIPS/Register/register[5][13] ), .A1(n4848), .B0(
        \i_MIPS/Register/register[13][13] ), .B1(n4843), .Y(n6397) );
  OA22X1 U9359 ( .A0(\i_MIPS/Register/register[7][13] ), .A1(n4881), .B0(
        \i_MIPS/Register/register[15][13] ), .B1(n4873), .Y(n6395) );
  NAND4X1 U9360 ( .A(n8564), .B(n8563), .C(n8562), .D(n8561), .Y(n8569) );
  OA22X1 U9361 ( .A0(\i_MIPS/Register/register[5][20] ), .A1(n4850), .B0(
        \i_MIPS/Register/register[13][20] ), .B1(n4843), .Y(n8563) );
  OA22X1 U9362 ( .A0(\i_MIPS/Register/register[7][20] ), .A1(n4884), .B0(
        \i_MIPS/Register/register[15][20] ), .B1(n4876), .Y(n8561) );
  OA22X1 U9363 ( .A0(\i_MIPS/Register/register[5][26] ), .A1(n4850), .B0(
        \i_MIPS/Register/register[13][26] ), .B1(n4843), .Y(n8366) );
  OA22X1 U9364 ( .A0(\i_MIPS/Register/register[7][26] ), .A1(n4884), .B0(
        \i_MIPS/Register/register[15][26] ), .B1(n4876), .Y(n8364) );
  NAND4X1 U9365 ( .A(n8050), .B(n8049), .C(n8048), .D(n8047), .Y(n8055) );
  NAND4X1 U9366 ( .A(n8232), .B(n8231), .C(n8230), .D(n8229), .Y(n8237) );
  OA22X1 U9367 ( .A0(\i_MIPS/Register/register[5][23] ), .A1(n4850), .B0(
        \i_MIPS/Register/register[13][23] ), .B1(n4842), .Y(n8231) );
  OA22X1 U9368 ( .A0(\i_MIPS/Register/register[7][23] ), .A1(n4883), .B0(
        \i_MIPS/Register/register[15][23] ), .B1(n4875), .Y(n8229) );
  OA22X1 U9369 ( .A0(\i_MIPS/Register/register[1][23] ), .A1(n4832), .B0(
        \i_MIPS/Register/register[9][23] ), .B1(n4831), .Y(n8232) );
  NAND4X1 U9370 ( .A(n7991), .B(n7990), .C(n7989), .D(n7988), .Y(n7996) );
  OA22X1 U9371 ( .A0(\i_MIPS/Register/register[5][22] ), .A1(n4851), .B0(
        \i_MIPS/Register/register[13][22] ), .B1(n4842), .Y(n7990) );
  OA22X1 U9372 ( .A0(\i_MIPS/Register/register[7][22] ), .A1(n4883), .B0(
        \i_MIPS/Register/register[15][22] ), .B1(n4875), .Y(n7988) );
  OA22X1 U9373 ( .A0(\i_MIPS/Register/register[1][22] ), .A1(n4832), .B0(
        \i_MIPS/Register/register[9][22] ), .B1(n4831), .Y(n7991) );
  OA22X1 U9374 ( .A0(\i_MIPS/Register/register[5][16] ), .A1(n4850), .B0(
        \i_MIPS/Register/register[13][16] ), .B1(n4842), .Y(n8173) );
  OA22X1 U9375 ( .A0(\i_MIPS/Register/register[7][16] ), .A1(n4883), .B0(
        \i_MIPS/Register/register[15][16] ), .B1(n4875), .Y(n8171) );
  OA22X1 U9376 ( .A0(\i_MIPS/Register/register[1][16] ), .A1(n4835), .B0(
        \i_MIPS/Register/register[9][16] ), .B1(n4831), .Y(n8174) );
  OA22X1 U9377 ( .A0(\i_MIPS/Register/register[5][24] ), .A1(n4851), .B0(
        \i_MIPS/Register/register[13][24] ), .B1(n4844), .Y(n8938) );
  OA22X1 U9378 ( .A0(\i_MIPS/Register/register[7][24] ), .A1(n4885), .B0(
        \i_MIPS/Register/register[15][24] ), .B1(n4877), .Y(n8936) );
  NAND4X1 U9379 ( .A(n8830), .B(n8829), .C(n8828), .D(n8827), .Y(n8835) );
  OA22X1 U9380 ( .A0(\i_MIPS/Register/register[5][2] ), .A1(n4850), .B0(
        \i_MIPS/Register/register[13][2] ), .B1(n4843), .Y(n8829) );
  OA22X1 U9381 ( .A0(\i_MIPS/Register/register[7][2] ), .A1(n4884), .B0(
        \i_MIPS/Register/register[15][2] ), .B1(n4876), .Y(n8827) );
  NAND4X1 U9382 ( .A(n8745), .B(n8744), .C(n8743), .D(n8742), .Y(n8750) );
  OA22X1 U9383 ( .A0(\i_MIPS/Register/register[5][3] ), .A1(n4850), .B0(
        \i_MIPS/Register/register[13][3] ), .B1(n4843), .Y(n8744) );
  OA22X1 U9384 ( .A0(\i_MIPS/Register/register[7][3] ), .A1(n4884), .B0(
        \i_MIPS/Register/register[15][3] ), .B1(n4876), .Y(n8742) );
  OA22X1 U9385 ( .A0(\i_MIPS/Register/register[1][3] ), .A1(n4834), .B0(
        \i_MIPS/Register/register[9][3] ), .B1(n4829), .Y(n8745) );
  NAND4X1 U9386 ( .A(n7214), .B(n7213), .C(n7212), .D(n7211), .Y(n7219) );
  OA22X1 U9387 ( .A0(\i_MIPS/Register/register[5][10] ), .A1(n4849), .B0(
        \i_MIPS/Register/register[13][10] ), .B1(n4841), .Y(n7213) );
  OA22X1 U9388 ( .A0(\i_MIPS/Register/register[7][10] ), .A1(n4882), .B0(
        \i_MIPS/Register/register[15][10] ), .B1(n4874), .Y(n7211) );
  OA22X1 U9389 ( .A0(\i_MIPS/Register/register[1][10] ), .A1(n4833), .B0(
        \i_MIPS/Register/register[9][10] ), .B1(n4830), .Y(n7214) );
  OA22X1 U9390 ( .A0(\i_MIPS/Register/register[5][4] ), .A1(n4849), .B0(
        \i_MIPS/Register/register[13][4] ), .B1(n4841), .Y(n7375) );
  OA22X1 U9391 ( .A0(\i_MIPS/Register/register[7][4] ), .A1(n4882), .B0(
        \i_MIPS/Register/register[15][4] ), .B1(n4874), .Y(n7373) );
  NAND4X1 U9392 ( .A(n8623), .B(n8622), .C(n8621), .D(n8620), .Y(n8628) );
  OA22X1 U9393 ( .A0(\i_MIPS/Register/register[5][27] ), .A1(n4850), .B0(
        \i_MIPS/Register/register[13][27] ), .B1(n4843), .Y(n8622) );
  OA22X1 U9394 ( .A0(\i_MIPS/Register/register[7][27] ), .A1(n4884), .B0(
        \i_MIPS/Register/register[15][27] ), .B1(n4876), .Y(n8620) );
  NAND4X1 U9395 ( .A(n8459), .B(n8458), .C(n8457), .D(n8456), .Y(n8464) );
  OA22X1 U9396 ( .A0(\i_MIPS/Register/register[5][25] ), .A1(n4850), .B0(
        \i_MIPS/Register/register[13][25] ), .B1(n4843), .Y(n8458) );
  OA22X1 U9397 ( .A0(\i_MIPS/Register/register[7][25] ), .A1(n4884), .B0(
        \i_MIPS/Register/register[15][25] ), .B1(n4876), .Y(n8456) );
  OA22X1 U9398 ( .A0(\i_MIPS/Register/register[5][28] ), .A1(n4851), .B0(
        \i_MIPS/Register/register[13][28] ), .B1(n4844), .Y(n9026) );
  OA22X1 U9399 ( .A0(\i_MIPS/Register/register[7][28] ), .A1(n4885), .B0(
        \i_MIPS/Register/register[15][28] ), .B1(n4877), .Y(n9024) );
  OA22X1 U9400 ( .A0(\i_MIPS/Register/register[1][28] ), .A1(n4835), .B0(
        \i_MIPS/Register/register[9][28] ), .B1(n4831), .Y(n9027) );
  NAND4X1 U9401 ( .A(n7895), .B(n7894), .C(n7893), .D(n7892), .Y(n7900) );
  OA22X1 U9402 ( .A0(\i_MIPS/Register/register[5][18] ), .A1(n4851), .B0(
        \i_MIPS/Register/register[13][18] ), .B1(n4842), .Y(n7894) );
  OA22X1 U9403 ( .A0(\i_MIPS/Register/register[7][18] ), .A1(n4883), .B0(
        \i_MIPS/Register/register[15][18] ), .B1(n4875), .Y(n7892) );
  OA22X1 U9404 ( .A0(\i_MIPS/Register/register[1][18] ), .A1(n4833), .B0(
        \i_MIPS/Register/register[9][18] ), .B1(n4831), .Y(n7895) );
  NAND4X1 U9405 ( .A(n7739), .B(n7738), .C(n7737), .D(n7736), .Y(n7744) );
  OA22X1 U9406 ( .A0(\i_MIPS/Register/register[5][17] ), .A1(n4851), .B0(
        \i_MIPS/Register/register[13][17] ), .B1(n4842), .Y(n7738) );
  OA22X1 U9407 ( .A0(\i_MIPS/Register/register[7][17] ), .A1(n4883), .B0(
        \i_MIPS/Register/register[15][17] ), .B1(n4875), .Y(n7736) );
  OA22X1 U9408 ( .A0(\i_MIPS/Register/register[1][17] ), .A1(n4835), .B0(
        \i_MIPS/Register/register[9][17] ), .B1(n4831), .Y(n7739) );
  NAND4X1 U9409 ( .A(n7124), .B(n7123), .C(n7122), .D(n7121), .Y(n7129) );
  OA22X1 U9410 ( .A0(\i_MIPS/Register/register[5][11] ), .A1(n4849), .B0(
        \i_MIPS/Register/register[13][11] ), .B1(n4841), .Y(n7123) );
  OA22X1 U9411 ( .A0(\i_MIPS/Register/register[7][11] ), .A1(n4882), .B0(
        \i_MIPS/Register/register[15][11] ), .B1(n4874), .Y(n7121) );
  NAND4X1 U9412 ( .A(n6308), .B(n6307), .C(n6306), .D(n6305), .Y(n6313) );
  NAND4X1 U9413 ( .A(n7072), .B(n7071), .C(n7070), .D(n7069), .Y(n7077) );
  NAND4X1 U9414 ( .A(n6806), .B(n6805), .C(n6804), .D(n6803), .Y(n6811) );
  OA22X1 U9415 ( .A0(\i_MIPS/Register/register[5][8] ), .A1(n4848), .B0(
        \i_MIPS/Register/register[13][8] ), .B1(n4844), .Y(n6805) );
  OA22X1 U9416 ( .A0(\i_MIPS/Register/register[7][8] ), .A1(n4881), .B0(
        \i_MIPS/Register/register[15][8] ), .B1(n4873), .Y(n6803) );
  NAND4X1 U9417 ( .A(n6736), .B(n6735), .C(n6734), .D(n6733), .Y(n6741) );
  OA22X1 U9418 ( .A0(\i_MIPS/Register/register[21][29] ), .A1(n4848), .B0(
        \i_MIPS/Register/register[29][29] ), .B1(n4843), .Y(n6735) );
  OA22X1 U9419 ( .A0(\i_MIPS/Register/register[23][29] ), .A1(n4881), .B0(
        \i_MIPS/Register/register[31][29] ), .B1(n4873), .Y(n6733) );
  OA22X1 U9420 ( .A0(\i_MIPS/Register/register[17][29] ), .A1(n4832), .B0(
        \i_MIPS/Register/register[25][29] ), .B1(n4829), .Y(n6736) );
  NAND4X1 U9421 ( .A(n6727), .B(n6726), .C(n6725), .D(n6724), .Y(n6732) );
  OA22X1 U9422 ( .A0(\i_MIPS/Register/register[5][29] ), .A1(n4848), .B0(
        \i_MIPS/Register/register[13][29] ), .B1(n4843), .Y(n6726) );
  OA22X1 U9423 ( .A0(\i_MIPS/Register/register[7][29] ), .A1(n4881), .B0(
        \i_MIPS/Register/register[15][29] ), .B1(n4873), .Y(n6724) );
  NAND4X1 U9424 ( .A(n6557), .B(n6556), .C(n6555), .D(n6554), .Y(n6562) );
  OA22X1 U9425 ( .A0(\i_MIPS/Register/register[21][0] ), .A1(n4848), .B0(
        \i_MIPS/Register/register[29][0] ), .B1(n4844), .Y(n6556) );
  OA22X1 U9426 ( .A0(\i_MIPS/Register/register[23][0] ), .A1(n4881), .B0(
        \i_MIPS/Register/register[31][0] ), .B1(n4873), .Y(n6554) );
  OA22X1 U9427 ( .A0(\i_MIPS/Register/register[17][0] ), .A1(n4832), .B0(
        \i_MIPS/Register/register[25][0] ), .B1(n4829), .Y(n6557) );
  NAND4X1 U9428 ( .A(n6548), .B(n6547), .C(n6546), .D(n6545), .Y(n6553) );
  OA22X1 U9429 ( .A0(\i_MIPS/Register/register[5][0] ), .A1(n4848), .B0(
        \i_MIPS/Register/register[13][0] ), .B1(n4843), .Y(n6547) );
  OA22X1 U9430 ( .A0(\i_MIPS/Register/register[7][0] ), .A1(n4881), .B0(
        \i_MIPS/Register/register[15][0] ), .B1(n4873), .Y(n6545) );
  OA22X1 U9431 ( .A0(\i_MIPS/Register/register[1][0] ), .A1(n4832), .B0(
        \i_MIPS/Register/register[9][0] ), .B1(n4829), .Y(n6548) );
  NAND4X1 U9432 ( .A(n6519), .B(n6518), .C(n6517), .D(n6516), .Y(n6524) );
  OA22XL U9433 ( .A0(\i_MIPS/Register/register[17][0] ), .A1(n6509), .B0(
        \i_MIPS/Register/register[25][0] ), .B1(n6508), .Y(n6519) );
  OA22XL U9434 ( .A0(\i_MIPS/Register/register[21][0] ), .A1(n6511), .B0(
        \i_MIPS/Register/register[29][0] ), .B1(n6510), .Y(n6518) );
  OA22XL U9435 ( .A0(\i_MIPS/Register/register[19][0] ), .A1(n179), .B0(
        \i_MIPS/Register/register[27][0] ), .B1(n6512), .Y(n6517) );
  NAND4X1 U9436 ( .A(n6502), .B(n6501), .C(n6500), .D(n6499), .Y(n6507) );
  OA22XL U9437 ( .A0(\i_MIPS/Register/register[1][0] ), .A1(n6509), .B0(
        \i_MIPS/Register/register[9][0] ), .B1(n6508), .Y(n6502) );
  OA22XL U9438 ( .A0(\i_MIPS/Register/register[5][0] ), .A1(n6511), .B0(
        \i_MIPS/Register/register[13][0] ), .B1(n6510), .Y(n6501) );
  OA22XL U9439 ( .A0(\i_MIPS/Register/register[3][0] ), .A1(n180), .B0(
        \i_MIPS/Register/register[11][0] ), .B1(n6512), .Y(n6500) );
  NAND4BX1 U9440 ( .AN(n9198), .B(n9197), .C(n9196), .D(n9195), .Y(n9209) );
  OAI221XL U9441 ( .A0(\i_MIPS/Register/register[2][31] ), .A1(n4947), .B0(
        \i_MIPS/Register/register[10][31] ), .B1(n4940), .C0(n9190), .Y(n9198)
         );
  NAND4BX1 U9442 ( .AN(n9305), .B(n9304), .C(n9303), .D(n9302), .Y(n9324) );
  OAI221XL U9443 ( .A0(\i_MIPS/Register/register[2][30] ), .A1(n4947), .B0(
        \i_MIPS/Register/register[10][30] ), .B1(n4940), .C0(n9297), .Y(n9305)
         );
  NAND4BX1 U9444 ( .AN(n9221), .B(n9220), .C(n9219), .D(n9218), .Y(n9236) );
  OA22XL U9445 ( .A0(\i_MIPS/Register/register[4][30] ), .A1(n9224), .B0(
        \i_MIPS/Register/register[12][30] ), .B1(n9223), .Y(n9220) );
  OA22XL U9446 ( .A0(\i_MIPS/Register/register[0][30] ), .A1(n9226), .B0(
        \i_MIPS/Register/register[8][30] ), .B1(n9225), .Y(n9219) );
  OAI221XL U9447 ( .A0(\i_MIPS/Register/register[2][30] ), .A1(n4921), .B0(
        \i_MIPS/Register/register[10][30] ), .B1(n4917), .C0(n9213), .Y(n9221)
         );
  NAND4BX1 U9448 ( .AN(n7659), .B(n7658), .C(n7657), .D(n7656), .Y(n7670) );
  OA22XL U9449 ( .A0(\i_MIPS/Register/register[4][1] ), .A1(n9224), .B0(
        \i_MIPS/Register/register[12][1] ), .B1(n9223), .Y(n7658) );
  OA22XL U9450 ( .A0(\i_MIPS/Register/register[0][1] ), .A1(n9226), .B0(
        \i_MIPS/Register/register[8][1] ), .B1(n9225), .Y(n7657) );
  OAI221XL U9451 ( .A0(\i_MIPS/Register/register[2][1] ), .A1(n4922), .B0(
        \i_MIPS/Register/register[10][1] ), .B1(n4916), .C0(n7651), .Y(n7659)
         );
  NAND4BX1 U9452 ( .AN(n7531), .B(n7530), .C(n7529), .D(n7528), .Y(n7542) );
  OAI221XL U9453 ( .A0(\i_MIPS/Register/register[2][6] ), .A1(n4946), .B0(
        \i_MIPS/Register/register[10][6] ), .B1(n4940), .C0(n7523), .Y(n7531)
         );
  NAND4BX1 U9454 ( .AN(n6832), .B(n6831), .C(n6830), .D(n6829), .Y(n6843) );
  OAI221XL U9455 ( .A0(\i_MIPS/Register/register[2][9] ), .A1(n4944), .B0(
        \i_MIPS/Register/register[10][9] ), .B1(n4942), .C0(n6824), .Y(n6832)
         );
  NAND4BX1 U9456 ( .AN(n6182), .B(n6181), .C(n6180), .D(n6179), .Y(n6193) );
  OAI221XL U9457 ( .A0(\i_MIPS/Register/register[2][12] ), .A1(n4944), .B0(
        \i_MIPS/Register/register[10][12] ), .B1(n4942), .C0(n6174), .Y(n6182)
         );
  OAI221XL U9458 ( .A0(\i_MIPS/Register/register[2][7] ), .A1(n4945), .B0(
        \i_MIPS/Register/register[10][7] ), .B1(n4484), .C0(n7431), .Y(n7439)
         );
  NAND4BX1 U9459 ( .AN(n6752), .B(n6751), .C(n6750), .D(n6749), .Y(n6763) );
  OAI221XL U9460 ( .A0(\i_MIPS/Register/register[2][8] ), .A1(n4944), .B0(
        \i_MIPS/Register/register[10][8] ), .B1(n4942), .C0(n6744), .Y(n6752)
         );
  NAND4BX1 U9461 ( .AN(n6915), .B(n6914), .C(n6913), .D(n6912), .Y(n6926) );
  OAI221XL U9462 ( .A0(\i_MIPS/Register/register[2][14] ), .A1(n4944), .B0(
        \i_MIPS/Register/register[10][14] ), .B1(n4942), .C0(n6907), .Y(n6915)
         );
  NAND4BX1 U9463 ( .AN(n7007), .B(n7006), .C(n7005), .D(n7004), .Y(n7018) );
  OA22X1 U9464 ( .A0(\i_MIPS/Register/register[4][15] ), .A1(n4952), .B0(
        \i_MIPS/Register/register[12][15] ), .B1(n4948), .Y(n7006) );
  OA22X1 U9465 ( .A0(\i_MIPS/Register/register[0][15] ), .A1(n4961), .B0(
        \i_MIPS/Register/register[8][15] ), .B1(n4957), .Y(n7005) );
  OAI221XL U9466 ( .A0(\i_MIPS/Register/register[2][15] ), .A1(n4945), .B0(
        \i_MIPS/Register/register[10][15] ), .B1(n4940), .C0(n6999), .Y(n7007)
         );
  NAND4BX1 U9467 ( .AN(n6334), .B(n6333), .C(n6332), .D(n6331), .Y(n6345) );
  OA22X1 U9468 ( .A0(\i_MIPS/Register/register[4][13] ), .A1(n4953), .B0(
        \i_MIPS/Register/register[12][13] ), .B1(n4948), .Y(n6333) );
  OA22X1 U9469 ( .A0(\i_MIPS/Register/register[0][13] ), .A1(n4961), .B0(
        \i_MIPS/Register/register[8][13] ), .B1(n4957), .Y(n6332) );
  OAI221XL U9470 ( .A0(\i_MIPS/Register/register[2][13] ), .A1(n4944), .B0(
        \i_MIPS/Register/register[10][13] ), .B1(n4942), .C0(n6326), .Y(n6334)
         );
  OA22X1 U9471 ( .A0(\i_MIPS/Register/register[4][21] ), .A1(n4953), .B0(
        \i_MIPS/Register/register[12][21] ), .B1(n4949), .Y(n8127) );
  OA22X1 U9472 ( .A0(\i_MIPS/Register/register[0][21] ), .A1(n4963), .B0(
        \i_MIPS/Register/register[8][21] ), .B1(n4958), .Y(n8126) );
  NAND4BX1 U9473 ( .AN(n7938), .B(n7937), .C(n7936), .D(n7935), .Y(n7949) );
  NAND4BX1 U9474 ( .AN(n7257), .B(n7256), .C(n7255), .D(n7254), .Y(n7268) );
  OAI221XL U9475 ( .A0(\i_MIPS/Register/register[2][10] ), .A1(n4945), .B0(
        \i_MIPS/Register/register[10][10] ), .B1(n4940), .C0(n7249), .Y(n7257)
         );
  NAND4BX1 U9476 ( .AN(n7681), .B(n7680), .C(n7679), .D(n7678), .Y(n7692) );
  OA22X1 U9477 ( .A0(\i_MIPS/Register/register[4][2] ), .A1(n4954), .B0(
        \i_MIPS/Register/register[12][2] ), .B1(n4950), .Y(n8872) );
  OA22X1 U9478 ( .A0(\i_MIPS/Register/register[0][2] ), .A1(n4962), .B0(
        \i_MIPS/Register/register[8][2] ), .B1(n4957), .Y(n8871) );
  OAI221XL U9479 ( .A0(\i_MIPS/Register/register[2][2] ), .A1(n4944), .B0(
        \i_MIPS/Register/register[10][2] ), .B1(n4939), .C0(n8865), .Y(n8873)
         );
  NAND4BX1 U9480 ( .AN(n8314), .B(n8313), .C(n8312), .D(n8311), .Y(n8325) );
  OA22X1 U9481 ( .A0(\i_MIPS/Register/register[4][23] ), .A1(n4954), .B0(
        \i_MIPS/Register/register[12][23] ), .B1(n4949), .Y(n8313) );
  OA22X1 U9482 ( .A0(\i_MIPS/Register/register[0][23] ), .A1(n4962), .B0(
        \i_MIPS/Register/register[8][23] ), .B1(n4959), .Y(n8312) );
  OAI221XL U9483 ( .A0(\i_MIPS/Register/register[2][23] ), .A1(n4947), .B0(
        \i_MIPS/Register/register[10][23] ), .B1(n4939), .C0(n8306), .Y(n8314)
         );
  OA22X1 U9484 ( .A0(\i_MIPS/Register/register[4][27] ), .A1(n4954), .B0(
        \i_MIPS/Register/register[12][27] ), .B1(n4950), .Y(n8698) );
  OA22X1 U9485 ( .A0(\i_MIPS/Register/register[0][27] ), .A1(n4961), .B0(
        \i_MIPS/Register/register[8][27] ), .B1(n4959), .Y(n8697) );
  OAI221XL U9486 ( .A0(\i_MIPS/Register/register[2][27] ), .A1(n4947), .B0(
        \i_MIPS/Register/register[10][27] ), .B1(n4940), .C0(n8691), .Y(n8699)
         );
  OA22X1 U9487 ( .A0(\i_MIPS/Register/register[4][24] ), .A1(n4954), .B0(
        \i_MIPS/Register/register[12][24] ), .B1(n4950), .Y(n8982) );
  OA22X1 U9488 ( .A0(\i_MIPS/Register/register[0][24] ), .A1(n4963), .B0(
        \i_MIPS/Register/register[8][24] ), .B1(n4957), .Y(n8981) );
  NAND4BX1 U9489 ( .AN(n9070), .B(n9069), .C(n9068), .D(n9067), .Y(n9081) );
  OA22X1 U9490 ( .A0(\i_MIPS/Register/register[4][28] ), .A1(n4952), .B0(
        \i_MIPS/Register/register[12][28] ), .B1(n4950), .Y(n9069) );
  OA22X1 U9491 ( .A0(\i_MIPS/Register/register[0][28] ), .A1(n4963), .B0(
        \i_MIPS/Register/register[8][28] ), .B1(n4957), .Y(n9068) );
  OAI221XL U9492 ( .A0(\i_MIPS/Register/register[2][28] ), .A1(n4947), .B0(
        \i_MIPS/Register/register[10][28] ), .B1(n4939), .C0(n9062), .Y(n9070)
         );
  NAND4BX1 U9493 ( .AN(n8788), .B(n8787), .C(n8786), .D(n8785), .Y(n8799) );
  OA22X1 U9494 ( .A0(\i_MIPS/Register/register[4][3] ), .A1(n4954), .B0(
        \i_MIPS/Register/register[12][3] ), .B1(n4950), .Y(n8787) );
  OA22X1 U9495 ( .A0(\i_MIPS/Register/register[0][3] ), .A1(n4962), .B0(
        \i_MIPS/Register/register[8][3] ), .B1(n4959), .Y(n8786) );
  OAI221XL U9496 ( .A0(\i_MIPS/Register/register[2][3] ), .A1(n4947), .B0(
        \i_MIPS/Register/register[10][3] ), .B1(n4939), .C0(n8780), .Y(n8788)
         );
  NAND4BX1 U9497 ( .AN(n8035), .B(n8034), .C(n8033), .D(n8032), .Y(n8046) );
  OA22X1 U9498 ( .A0(\i_MIPS/Register/register[4][22] ), .A1(n4953), .B0(
        \i_MIPS/Register/register[12][22] ), .B1(n4949), .Y(n8034) );
  OA22X1 U9499 ( .A0(\i_MIPS/Register/register[0][22] ), .A1(n4963), .B0(
        \i_MIPS/Register/register[8][22] ), .B1(n4959), .Y(n8033) );
  OAI221XL U9500 ( .A0(\i_MIPS/Register/register[2][22] ), .A1(n4946), .B0(
        \i_MIPS/Register/register[10][22] ), .B1(n4939), .C0(n8027), .Y(n8035)
         );
  NAND4BX1 U9501 ( .AN(n7419), .B(n7418), .C(n7417), .D(n7416), .Y(n7430) );
  OA22X1 U9502 ( .A0(\i_MIPS/Register/register[4][4] ), .A1(n4952), .B0(
        \i_MIPS/Register/register[12][4] ), .B1(n4949), .Y(n7418) );
  OA22X1 U9503 ( .A0(\i_MIPS/Register/register[0][4] ), .A1(n4962), .B0(
        \i_MIPS/Register/register[8][4] ), .B1(n4958), .Y(n7417) );
  OAI221XL U9504 ( .A0(\i_MIPS/Register/register[2][4] ), .A1(n4945), .B0(
        \i_MIPS/Register/register[10][4] ), .B1(n4940), .C0(n7411), .Y(n7419)
         );
  NAND4BX1 U9505 ( .AN(n8608), .B(n8607), .C(n8606), .D(n8605), .Y(n8619) );
  OA22X1 U9506 ( .A0(\i_MIPS/Register/register[4][20] ), .A1(n4954), .B0(
        \i_MIPS/Register/register[12][20] ), .B1(n4950), .Y(n8607) );
  OA22X1 U9507 ( .A0(\i_MIPS/Register/register[0][20] ), .A1(n4963), .B0(
        \i_MIPS/Register/register[8][20] ), .B1(n4959), .Y(n8606) );
  OAI221XL U9508 ( .A0(\i_MIPS/Register/register[2][20] ), .A1(n4947), .B0(
        \i_MIPS/Register/register[10][20] ), .B1(n4939), .C0(n8600), .Y(n8608)
         );
  NAND4BX1 U9509 ( .AN(n8217), .B(n8216), .C(n8215), .D(n8214), .Y(n8228) );
  OA22X1 U9510 ( .A0(\i_MIPS/Register/register[4][16] ), .A1(n4953), .B0(
        \i_MIPS/Register/register[12][16] ), .B1(n4949), .Y(n8216) );
  OA22X1 U9511 ( .A0(\i_MIPS/Register/register[0][16] ), .A1(n4963), .B0(
        \i_MIPS/Register/register[8][16] ), .B1(n4958), .Y(n8215) );
  OAI221XL U9512 ( .A0(\i_MIPS/Register/register[2][16] ), .A1(n4947), .B0(
        \i_MIPS/Register/register[10][16] ), .B1(n4939), .C0(n8209), .Y(n8217)
         );
  NAND4BX1 U9513 ( .AN(n6694), .B(n6693), .C(n6692), .D(n6691), .Y(n6705) );
  OA22X1 U9514 ( .A0(\i_MIPS/Register/register[4][29] ), .A1(n4953), .B0(
        \i_MIPS/Register/register[12][29] ), .B1(n4948), .Y(n6693) );
  OA22X1 U9515 ( .A0(\i_MIPS/Register/register[0][29] ), .A1(n4961), .B0(
        \i_MIPS/Register/register[8][29] ), .B1(n4957), .Y(n6692) );
  OAI221XL U9516 ( .A0(\i_MIPS/Register/register[2][29] ), .A1(n4944), .B0(
        \i_MIPS/Register/register[10][29] ), .B1(n4942), .C0(n6686), .Y(n6694)
         );
  NAND4BX1 U9517 ( .AN(n8411), .B(n8410), .C(n8409), .D(n8408), .Y(n8422) );
  OA22X1 U9518 ( .A0(\i_MIPS/Register/register[4][26] ), .A1(n4954), .B0(
        \i_MIPS/Register/register[12][26] ), .B1(n4950), .Y(n8410) );
  OA22X1 U9519 ( .A0(\i_MIPS/Register/register[0][26] ), .A1(n4961), .B0(
        \i_MIPS/Register/register[8][26] ), .B1(n4959), .Y(n8409) );
  OAI221XL U9520 ( .A0(\i_MIPS/Register/register[2][26] ), .A1(n4947), .B0(
        \i_MIPS/Register/register[10][26] ), .B1(n4939), .C0(n8403), .Y(n8411)
         );
  OAI221XL U9521 ( .A0(\i_MIPS/Register/register[2][5] ), .A1(n4945), .B0(
        \i_MIPS/Register/register[10][5] ), .B1(n4940), .C0(n7333), .Y(n7341)
         );
  OA22X1 U9522 ( .A0(\i_MIPS/Register/register[0][11] ), .A1(n4962), .B0(
        \i_MIPS/Register/register[8][11] ), .B1(n4958), .Y(n7165) );
  OAI221XL U9523 ( .A0(\i_MIPS/Register/register[2][11] ), .A1(n4945), .B0(
        \i_MIPS/Register/register[10][11] ), .B1(n4940), .C0(n7159), .Y(n7167)
         );
  NAND4BX1 U9524 ( .AN(n9207), .B(n9206), .C(n9205), .D(n9204), .Y(n9208) );
  OAI221XL U9525 ( .A0(\i_MIPS/Register/register[18][31] ), .A1(n4944), .B0(
        \i_MIPS/Register/register[26][31] ), .B1(n4940), .C0(n9199), .Y(n9207)
         );
  NAND4BX1 U9526 ( .AN(n9322), .B(n9321), .C(n9320), .D(n9319), .Y(n9323) );
  OAI221XL U9527 ( .A0(\i_MIPS/Register/register[18][30] ), .A1(n4946), .B0(
        \i_MIPS/Register/register[26][30] ), .B1(n4940), .C0(n9306), .Y(n9322)
         );
  NAND4BX1 U9528 ( .AN(n9234), .B(n9233), .C(n9232), .D(n9231), .Y(n9235) );
  OA22XL U9529 ( .A0(\i_MIPS/Register/register[20][30] ), .A1(n9224), .B0(
        \i_MIPS/Register/register[28][30] ), .B1(n9223), .Y(n9233) );
  OA22XL U9530 ( .A0(\i_MIPS/Register/register[16][30] ), .A1(n9226), .B0(
        \i_MIPS/Register/register[24][30] ), .B1(n9225), .Y(n9232) );
  OAI221XL U9531 ( .A0(\i_MIPS/Register/register[18][30] ), .A1(n4921), .B0(
        \i_MIPS/Register/register[26][30] ), .B1(n4917), .C0(n9222), .Y(n9234)
         );
  NAND4BX1 U9532 ( .AN(n7607), .B(n7606), .C(n7605), .D(n7604), .Y(n7608) );
  OAI221XL U9533 ( .A0(\i_MIPS/Register/register[18][1] ), .A1(n4946), .B0(
        \i_MIPS/Register/register[26][1] ), .B1(n4941), .C0(n7599), .Y(n7607)
         );
  NAND4BX1 U9534 ( .AN(n7668), .B(n7667), .C(n7666), .D(n7665), .Y(n7669) );
  OA22XL U9535 ( .A0(\i_MIPS/Register/register[20][1] ), .A1(n9224), .B0(
        \i_MIPS/Register/register[28][1] ), .B1(n9223), .Y(n7667) );
  OA22XL U9536 ( .A0(\i_MIPS/Register/register[16][1] ), .A1(n9226), .B0(
        \i_MIPS/Register/register[24][1] ), .B1(n9225), .Y(n7666) );
  OAI221XL U9537 ( .A0(\i_MIPS/Register/register[18][1] ), .A1(n4922), .B0(
        \i_MIPS/Register/register[26][1] ), .B1(n4916), .C0(n7660), .Y(n7668)
         );
  NAND4BX1 U9538 ( .AN(n7540), .B(n7539), .C(n7538), .D(n7537), .Y(n7541) );
  OAI221XL U9539 ( .A0(\i_MIPS/Register/register[18][6] ), .A1(n4946), .B0(
        \i_MIPS/Register/register[26][6] ), .B1(n4941), .C0(n7532), .Y(n7540)
         );
  NAND4BX1 U9540 ( .AN(n6841), .B(n6840), .C(n6839), .D(n6838), .Y(n6842) );
  OAI221XL U9541 ( .A0(\i_MIPS/Register/register[18][9] ), .A1(n4944), .B0(
        \i_MIPS/Register/register[26][9] ), .B1(n4942), .C0(n6833), .Y(n6841)
         );
  NAND4BX1 U9542 ( .AN(n6191), .B(n6190), .C(n6189), .D(n6188), .Y(n6192) );
  OAI221XL U9543 ( .A0(\i_MIPS/Register/register[18][12] ), .A1(n4944), .B0(
        \i_MIPS/Register/register[26][12] ), .B1(n4942), .C0(n6183), .Y(n6191)
         );
  OAI221XL U9544 ( .A0(\i_MIPS/Register/register[18][7] ), .A1(n4945), .B0(
        \i_MIPS/Register/register[26][7] ), .B1(n4484), .C0(n7440), .Y(n7448)
         );
  NAND4BX1 U9545 ( .AN(n6761), .B(n6760), .C(n6759), .D(n6758), .Y(n6762) );
  OAI221XL U9546 ( .A0(\i_MIPS/Register/register[18][8] ), .A1(n4944), .B0(
        \i_MIPS/Register/register[26][8] ), .B1(n4942), .C0(n6753), .Y(n6761)
         );
  NAND4BX1 U9547 ( .AN(n6924), .B(n6923), .C(n6922), .D(n6921), .Y(n6925) );
  OAI221XL U9548 ( .A0(\i_MIPS/Register/register[18][14] ), .A1(n4945), .B0(
        \i_MIPS/Register/register[26][14] ), .B1(n4940), .C0(n6916), .Y(n6924)
         );
  NAND4BX1 U9549 ( .AN(n7016), .B(n7015), .C(n7014), .D(n7013), .Y(n7017) );
  OAI221XL U9550 ( .A0(\i_MIPS/Register/register[18][15] ), .A1(n4945), .B0(
        \i_MIPS/Register/register[26][15] ), .B1(n4942), .C0(n7008), .Y(n7016)
         );
  NAND4BX1 U9551 ( .AN(n6343), .B(n6342), .C(n6341), .D(n6340), .Y(n6344) );
  OA22X1 U9552 ( .A0(\i_MIPS/Register/register[20][13] ), .A1(n4952), .B0(
        \i_MIPS/Register/register[28][13] ), .B1(n4948), .Y(n6342) );
  OA22X1 U9553 ( .A0(\i_MIPS/Register/register[16][13] ), .A1(n4961), .B0(
        \i_MIPS/Register/register[24][13] ), .B1(n4957), .Y(n6341) );
  OAI221XL U9554 ( .A0(\i_MIPS/Register/register[18][13] ), .A1(n4944), .B0(
        \i_MIPS/Register/register[26][13] ), .B1(n4942), .C0(n6335), .Y(n6343)
         );
  NAND4BX1 U9555 ( .AN(n8137), .B(n8136), .C(n8135), .D(n8134), .Y(n8138) );
  OA22X1 U9556 ( .A0(\i_MIPS/Register/register[20][21] ), .A1(n4953), .B0(
        \i_MIPS/Register/register[28][21] ), .B1(n4949), .Y(n8136) );
  OA22X1 U9557 ( .A0(\i_MIPS/Register/register[16][21] ), .A1(n4963), .B0(
        \i_MIPS/Register/register[24][21] ), .B1(n4959), .Y(n8135) );
  OAI221XL U9558 ( .A0(\i_MIPS/Register/register[18][21] ), .A1(n4947), .B0(
        \i_MIPS/Register/register[26][21] ), .B1(n4939), .C0(n8129), .Y(n8137)
         );
  NAND4BX1 U9559 ( .AN(n7947), .B(n7946), .C(n7945), .D(n7944), .Y(n7948) );
  OAI221XL U9560 ( .A0(\i_MIPS/Register/register[18][18] ), .A1(n4946), .B0(
        \i_MIPS/Register/register[26][18] ), .B1(n4940), .C0(n7939), .Y(n7947)
         );
  NAND4BX1 U9561 ( .AN(n7266), .B(n7265), .C(n7264), .D(n7263), .Y(n7267) );
  OA22XL U9562 ( .A0(\i_MIPS/Register/register[20][19] ), .A1(n9224), .B0(
        \i_MIPS/Register/register[28][19] ), .B1(n9223), .Y(n7772) );
  OA22XL U9563 ( .A0(\i_MIPS/Register/register[16][19] ), .A1(n9226), .B0(
        \i_MIPS/Register/register[24][19] ), .B1(n9225), .Y(n7771) );
  NAND4BX1 U9564 ( .AN(n7690), .B(n7689), .C(n7688), .D(n7687), .Y(n7691) );
  OAI221XL U9565 ( .A0(\i_MIPS/Register/register[18][17] ), .A1(n4946), .B0(
        \i_MIPS/Register/register[26][17] ), .B1(n4941), .C0(n7682), .Y(n7690)
         );
  NAND4BX1 U9566 ( .AN(n8882), .B(n8881), .C(n8880), .D(n8879), .Y(n8883) );
  OA22X1 U9567 ( .A0(\i_MIPS/Register/register[20][2] ), .A1(n4954), .B0(
        \i_MIPS/Register/register[28][2] ), .B1(n4950), .Y(n8881) );
  OA22X1 U9568 ( .A0(\i_MIPS/Register/register[16][2] ), .A1(n4962), .B0(
        \i_MIPS/Register/register[24][2] ), .B1(n4957), .Y(n8880) );
  OAI221XL U9569 ( .A0(\i_MIPS/Register/register[18][2] ), .A1(n4947), .B0(
        \i_MIPS/Register/register[26][2] ), .B1(n4939), .C0(n8874), .Y(n8882)
         );
  NAND4BX1 U9570 ( .AN(n8323), .B(n8322), .C(n8321), .D(n8320), .Y(n8324) );
  OA22X1 U9571 ( .A0(\i_MIPS/Register/register[20][23] ), .A1(n4954), .B0(
        \i_MIPS/Register/register[28][23] ), .B1(n4950), .Y(n8322) );
  OA22X1 U9572 ( .A0(\i_MIPS/Register/register[16][23] ), .A1(n4963), .B0(
        \i_MIPS/Register/register[24][23] ), .B1(n4959), .Y(n8321) );
  OAI221XL U9573 ( .A0(\i_MIPS/Register/register[18][23] ), .A1(n4947), .B0(
        \i_MIPS/Register/register[26][23] ), .B1(n4939), .C0(n8315), .Y(n8323)
         );
  OA22X1 U9574 ( .A0(\i_MIPS/Register/register[20][27] ), .A1(n4954), .B0(
        \i_MIPS/Register/register[28][27] ), .B1(n4949), .Y(n8707) );
  OA22X1 U9575 ( .A0(\i_MIPS/Register/register[16][27] ), .A1(n4962), .B0(
        \i_MIPS/Register/register[24][27] ), .B1(n4959), .Y(n8706) );
  OAI221XL U9576 ( .A0(\i_MIPS/Register/register[18][27] ), .A1(n4947), .B0(
        \i_MIPS/Register/register[26][27] ), .B1(n4939), .C0(n8700), .Y(n8708)
         );
  OA22X1 U9577 ( .A0(\i_MIPS/Register/register[20][24] ), .A1(n4954), .B0(
        \i_MIPS/Register/register[28][24] ), .B1(n4950), .Y(n8991) );
  OA22X1 U9578 ( .A0(\i_MIPS/Register/register[16][24] ), .A1(n4961), .B0(
        \i_MIPS/Register/register[24][24] ), .B1(n4957), .Y(n8990) );
  NAND4BX1 U9579 ( .AN(n7843), .B(n7842), .C(n7841), .D(n7840), .Y(n7844) );
  OAI221XL U9580 ( .A0(\i_MIPS/Register/register[18][19] ), .A1(n4946), .B0(
        \i_MIPS/Register/register[26][19] ), .B1(n4940), .C0(n7835), .Y(n7843)
         );
  NAND4BX1 U9581 ( .AN(n9079), .B(n9078), .C(n9077), .D(n9076), .Y(n9080) );
  OA22X1 U9582 ( .A0(\i_MIPS/Register/register[20][28] ), .A1(n4953), .B0(
        \i_MIPS/Register/register[28][28] ), .B1(n4950), .Y(n9078) );
  OA22X1 U9583 ( .A0(\i_MIPS/Register/register[16][28] ), .A1(n4961), .B0(
        \i_MIPS/Register/register[24][28] ), .B1(n4957), .Y(n9077) );
  OAI221XL U9584 ( .A0(\i_MIPS/Register/register[18][28] ), .A1(n4947), .B0(
        \i_MIPS/Register/register[26][28] ), .B1(n4939), .C0(n9071), .Y(n9079)
         );
  NAND4BX1 U9585 ( .AN(n8797), .B(n8796), .C(n8795), .D(n8794), .Y(n8798) );
  OA22X1 U9586 ( .A0(\i_MIPS/Register/register[20][3] ), .A1(n4954), .B0(
        \i_MIPS/Register/register[28][3] ), .B1(n4949), .Y(n8796) );
  OA22X1 U9587 ( .A0(\i_MIPS/Register/register[16][3] ), .A1(n4963), .B0(
        \i_MIPS/Register/register[24][3] ), .B1(n4959), .Y(n8795) );
  OAI221XL U9588 ( .A0(\i_MIPS/Register/register[18][3] ), .A1(n4947), .B0(
        \i_MIPS/Register/register[26][3] ), .B1(n4939), .C0(n8789), .Y(n8797)
         );
  OA22X1 U9589 ( .A0(\i_MIPS/Register/register[20][22] ), .A1(n4953), .B0(
        \i_MIPS/Register/register[28][22] ), .B1(n4949), .Y(n8043) );
  OA22X1 U9590 ( .A0(\i_MIPS/Register/register[16][22] ), .A1(n4963), .B0(
        \i_MIPS/Register/register[24][22] ), .B1(n4958), .Y(n8042) );
  OAI221XL U9591 ( .A0(\i_MIPS/Register/register[18][22] ), .A1(n4946), .B0(
        \i_MIPS/Register/register[26][22] ), .B1(n4939), .C0(n8036), .Y(n8044)
         );
  OA22X1 U9592 ( .A0(\i_MIPS/Register/register[20][4] ), .A1(n4952), .B0(
        \i_MIPS/Register/register[28][4] ), .B1(n4948), .Y(n7427) );
  OA22X1 U9593 ( .A0(\i_MIPS/Register/register[16][4] ), .A1(n4962), .B0(
        \i_MIPS/Register/register[24][4] ), .B1(n4958), .Y(n7426) );
  OA22X1 U9594 ( .A0(\i_MIPS/Register/register[20][29] ), .A1(n4952), .B0(
        \i_MIPS/Register/register[28][29] ), .B1(n4948), .Y(n6702) );
  OA22X1 U9595 ( .A0(\i_MIPS/Register/register[16][29] ), .A1(n4961), .B0(
        \i_MIPS/Register/register[24][29] ), .B1(n4957), .Y(n6701) );
  OAI221XL U9596 ( .A0(\i_MIPS/Register/register[18][29] ), .A1(n4944), .B0(
        \i_MIPS/Register/register[26][29] ), .B1(n4942), .C0(n6695), .Y(n6703)
         );
  NAND4BX1 U9597 ( .AN(n8617), .B(n8616), .C(n8615), .D(n8614), .Y(n8618) );
  OA22X1 U9598 ( .A0(\i_MIPS/Register/register[20][20] ), .A1(n4954), .B0(
        \i_MIPS/Register/register[28][20] ), .B1(n4950), .Y(n8616) );
  OA22X1 U9599 ( .A0(\i_MIPS/Register/register[16][20] ), .A1(n4961), .B0(
        \i_MIPS/Register/register[24][20] ), .B1(n4959), .Y(n8615) );
  OAI221XL U9600 ( .A0(\i_MIPS/Register/register[18][20] ), .A1(n4947), .B0(
        \i_MIPS/Register/register[26][20] ), .B1(n4939), .C0(n8609), .Y(n8617)
         );
  NAND4BX1 U9601 ( .AN(n8226), .B(n8225), .C(n8224), .D(n8223), .Y(n8227) );
  OA22X1 U9602 ( .A0(\i_MIPS/Register/register[20][16] ), .A1(n4954), .B0(
        \i_MIPS/Register/register[28][16] ), .B1(n4949), .Y(n8225) );
  OA22X1 U9603 ( .A0(\i_MIPS/Register/register[16][16] ), .A1(n4961), .B0(
        \i_MIPS/Register/register[24][16] ), .B1(n4959), .Y(n8224) );
  OAI221XL U9604 ( .A0(\i_MIPS/Register/register[18][16] ), .A1(n4947), .B0(
        \i_MIPS/Register/register[26][16] ), .B1(n4939), .C0(n8218), .Y(n8226)
         );
  NAND4BX1 U9605 ( .AN(n8420), .B(n8419), .C(n8418), .D(n8417), .Y(n8421) );
  OA22X1 U9606 ( .A0(\i_MIPS/Register/register[20][26] ), .A1(n4954), .B0(
        \i_MIPS/Register/register[28][26] ), .B1(n4950), .Y(n8419) );
  OA22X1 U9607 ( .A0(\i_MIPS/Register/register[16][26] ), .A1(n4961), .B0(
        \i_MIPS/Register/register[24][26] ), .B1(n4959), .Y(n8418) );
  OAI221XL U9608 ( .A0(\i_MIPS/Register/register[18][26] ), .A1(n4947), .B0(
        \i_MIPS/Register/register[26][26] ), .B1(n4939), .C0(n8412), .Y(n8420)
         );
  OAI221XL U9609 ( .A0(\i_MIPS/Register/register[18][5] ), .A1(n4945), .B0(
        \i_MIPS/Register/register[26][5] ), .B1(n4942), .C0(n7342), .Y(n7350)
         );
  NAND4BX1 U9610 ( .AN(n7176), .B(n7175), .C(n7174), .D(n7173), .Y(n7177) );
  OA22X1 U9611 ( .A0(\i_MIPS/Register/register[20][11] ), .A1(n4952), .B0(
        \i_MIPS/Register/register[28][11] ), .B1(n4948), .Y(n7175) );
  OA22X1 U9612 ( .A0(\i_MIPS/Register/register[16][11] ), .A1(n4962), .B0(
        \i_MIPS/Register/register[24][11] ), .B1(n4958), .Y(n7174) );
  OAI221XL U9613 ( .A0(\i_MIPS/Register/register[18][11] ), .A1(n4945), .B0(
        \i_MIPS/Register/register[26][11] ), .B1(n4940), .C0(n7168), .Y(n7176)
         );
  AO21XL U9614 ( .A0(\i_MIPS/ALUin1[0] ), .A1(n6432), .B0(n7621), .Y(n6429) );
  MXI2X1 U9615 ( .A(\i_MIPS/n352 ), .B(net98501), .S0(n5505), .Y(\i_MIPS/n543 ) );
  OAI221X1 U9616 ( .A0(net112231), .A1(n1628), .B0(net112137), .B1(n3287), 
        .C0(n6162), .Y(n6163) );
  MXI2X1 U9617 ( .A(\i_MIPS/n341 ), .B(n4526), .S0(n5502), .Y(\i_MIPS/n532 )
         );
  MXI2X1 U9618 ( .A(\i_MIPS/n340 ), .B(n4525), .S0(n5502), .Y(\i_MIPS/n531 )
         );
  MXI2X1 U9619 ( .A(\i_MIPS/n367 ), .B(n4562), .S0(n5505), .Y(\i_MIPS/n558 )
         );
  MXI2X1 U9620 ( .A(\i_MIPS/n366 ), .B(n4529), .S0(n5505), .Y(\i_MIPS/n557 )
         );
  MXI2X1 U9621 ( .A(\i_MIPS/n365 ), .B(net130474), .S0(n5502), .Y(
        \i_MIPS/n556 ) );
  MXI2X1 U9622 ( .A(\i_MIPS/n364 ), .B(n4542), .S0(n5502), .Y(\i_MIPS/n555 )
         );
  MXI2X1 U9623 ( .A(\i_MIPS/n363 ), .B(n4541), .S0(n5503), .Y(\i_MIPS/n554 )
         );
  MXI2X1 U9624 ( .A(\i_MIPS/n362 ), .B(n4558), .S0(n5503), .Y(\i_MIPS/n553 )
         );
  MXI2X1 U9625 ( .A(\i_MIPS/n361 ), .B(n4540), .S0(n5502), .Y(\i_MIPS/n552 )
         );
  MXI2X1 U9626 ( .A(\i_MIPS/n360 ), .B(n4539), .S0(n5503), .Y(\i_MIPS/n551 )
         );
  MXI2X1 U9627 ( .A(\i_MIPS/n359 ), .B(n4561), .S0(n5503), .Y(\i_MIPS/n550 )
         );
  MXI2X1 U9628 ( .A(n6947), .B(n4537), .S0(n5505), .Y(\i_MIPS/n548 ) );
  MXI2X1 U9629 ( .A(\i_MIPS/n355 ), .B(n4535), .S0(n5502), .Y(\i_MIPS/n546 )
         );
  MXI2X1 U9630 ( .A(\i_MIPS/n354 ), .B(n4560), .S0(n5502), .Y(\i_MIPS/n545 )
         );
  MXI2X1 U9631 ( .A(\i_MIPS/n351 ), .B(n4534), .S0(n5505), .Y(\i_MIPS/n542 )
         );
  MXI2X1 U9632 ( .A(\i_MIPS/n350 ), .B(n4533), .S0(n5503), .Y(\i_MIPS/n541 )
         );
  MXI2X1 U9633 ( .A(\i_MIPS/n349 ), .B(n4528), .S0(n5504), .Y(\i_MIPS/n540 )
         );
  MXI2X1 U9634 ( .A(\i_MIPS/n348 ), .B(n4557), .S0(n5509), .Y(\i_MIPS/n539 )
         );
  MXI2X1 U9635 ( .A(\i_MIPS/n347 ), .B(net130420), .S0(n5506), .Y(
        \i_MIPS/n538 ) );
  MXI2X1 U9636 ( .A(\i_MIPS/n346 ), .B(n4532), .S0(n5506), .Y(\i_MIPS/n537 )
         );
  MXI2X1 U9637 ( .A(\i_MIPS/n345 ), .B(n4531), .S0(n5506), .Y(\i_MIPS/n536 )
         );
  CLKINVX1 U9638 ( .A(n7282), .Y(n7628) );
  MXI2X1 U9639 ( .A(\i_MIPS/n336 ), .B(\i_MIPS/n337 ), .S0(n5504), .Y(
        \i_MIPS/n526 ) );
  MXI2X1 U9640 ( .A(\i_MIPS/n334 ), .B(\i_MIPS/n335 ), .S0(n5504), .Y(
        \i_MIPS/n524 ) );
  MXI2X1 U9641 ( .A(\i_MIPS/n310 ), .B(\i_MIPS/n311 ), .S0(n5504), .Y(
        \i_MIPS/n479 ) );
  MXI2X1 U9642 ( .A(\i_MIPS/n308 ), .B(\i_MIPS/n309 ), .S0(n5504), .Y(
        \i_MIPS/n436 ) );
  MXI2X1 U9643 ( .A(\i_MIPS/n306 ), .B(\i_MIPS/n307 ), .S0(n5503), .Y(
        \i_MIPS/n434 ) );
  MXI2X1 U9644 ( .A(\i_MIPS/n296 ), .B(n3820), .S0(n5505), .Y(\i_MIPS/n424 )
         );
  MXI2X1 U9645 ( .A(\i_MIPS/n292 ), .B(\i_MIPS/n293 ), .S0(n5503), .Y(
        \i_MIPS/n420 ) );
  MXI2X1 U9646 ( .A(\i_MIPS/n290 ), .B(\i_MIPS/n291 ), .S0(n5503), .Y(
        \i_MIPS/n418 ) );
  MXI2X1 U9647 ( .A(\i_MIPS/n280 ), .B(\i_MIPS/n281 ), .S0(n5506), .Y(
        \i_MIPS/n408 ) );
  MXI2X1 U9648 ( .A(\i_MIPS/n278 ), .B(\i_MIPS/n279 ), .S0(n5505), .Y(
        \i_MIPS/n406 ) );
  MXI2X1 U9649 ( .A(\i_MIPS/n256 ), .B(\i_MIPS/n257 ), .S0(n5505), .Y(
        \i_MIPS/n384 ) );
  MXI2X1 U9650 ( .A(\i_MIPS/n254 ), .B(\i_MIPS/n255 ), .S0(n5510), .Y(
        \i_MIPS/n382 ) );
  MXI2X1 U9651 ( .A(\i_MIPS/n252 ), .B(\i_MIPS/n253 ), .S0(n5502), .Y(
        \i_MIPS/n380 ) );
  MXI2X1 U9652 ( .A(\i_MIPS/n250 ), .B(\i_MIPS/n251 ), .S0(n5504), .Y(
        \i_MIPS/n378 ) );
  MXI2X1 U9653 ( .A(\i_MIPS/n248 ), .B(\i_MIPS/n249 ), .S0(n5502), .Y(
        \i_MIPS/n376 ) );
  MXI2X1 U9654 ( .A(\i_MIPS/n246 ), .B(\i_MIPS/n247 ), .S0(n5504), .Y(
        \i_MIPS/n374 ) );
  NAND2XL U9655 ( .A(n9141), .B(\i_MIPS/ALU/N303 ), .Y(n9148) );
  XOR2X4 U9656 ( .A(n11379), .B(\i_MIPS/PC/n24 ), .Y(n4665) );
  NOR3X1 U9657 ( .A(\i_MIPS/Hazard_detection/n8 ), .B(
        \i_MIPS/Hazard_detection/n9 ), .C(\i_MIPS/Hazard_detection/n10 ), .Y(
        \i_MIPS/Hazard_detection/n7 ) );
  XOR2XL U9658 ( .A(\i_MIPS/ID_EX[114] ), .B(\i_MIPS/IR_ID[24] ), .Y(
        \i_MIPS/Hazard_detection/n8 ) );
  XOR2XL U9659 ( .A(\i_MIPS/ID_EX[112] ), .B(\i_MIPS/IR_ID[22] ), .Y(
        \i_MIPS/Hazard_detection/n9 ) );
  XOR2XL U9660 ( .A(n5588), .B(\i_MIPS/ID_EX[115] ), .Y(
        \i_MIPS/Hazard_detection/n10 ) );
  NOR3X1 U9661 ( .A(\i_MIPS/Hazard_detection/n11 ), .B(
        \i_MIPS/Hazard_detection/n12 ), .C(\i_MIPS/Hazard_detection/n13 ), .Y(
        \i_MIPS/Hazard_detection/n4 ) );
  XOR2XL U9662 ( .A(\i_MIPS/IR_ID[19] ), .B(\i_MIPS/ID_EX[114] ), .Y(
        \i_MIPS/Hazard_detection/n11 ) );
  XOR2XL U9663 ( .A(\i_MIPS/IR_ID[17] ), .B(\i_MIPS/ID_EX[112] ), .Y(
        \i_MIPS/Hazard_detection/n12 ) );
  XOR2XL U9664 ( .A(net108963), .B(\i_MIPS/ID_EX[115] ), .Y(
        \i_MIPS/Hazard_detection/n13 ) );
  NAND2XL U9665 ( .A(\i_MIPS/IF_ID_1 ), .B(net130576), .Y(n10832) );
  AOI2BB2X4 U9666 ( .B0(n4676), .B1(\I_cache/cache[4][135] ), .A0N(n5290), 
        .A1N(n3209), .Y(n5980) );
  AOI2BB2X4 U9667 ( .B0(n4677), .B1(\I_cache/cache[4][137] ), .A0N(n5317), 
        .A1N(n3210), .Y(n5978) );
  AOI2BB2X4 U9668 ( .B0(n4678), .B1(\I_cache/cache[4][148] ), .A0N(n5318), 
        .A1N(n3211), .Y(n5970) );
  AOI2BB2X4 U9669 ( .B0(n4679), .B1(\I_cache/cache[4][152] ), .A0N(n5287), 
        .A1N(n3212), .Y(n5958) );
  AOI2BB2X4 U9670 ( .B0(n4680), .B1(\I_cache/cache[4][151] ), .A0N(n5288), 
        .A1N(n3213), .Y(n5966) );
  AOI2BB2X4 U9671 ( .B0(n4681), .B1(\I_cache/cache[4][139] ), .A0N(n5288), 
        .A1N(n3215), .Y(n5953) );
  XOR2X4 U9672 ( .A(n11364), .B(\i_MIPS/PC/n9 ), .Y(n4685) );
  NAND2XL U9673 ( .A(n10198), .B(ICACHE_addr[19]), .Y(n9363) );
  AND2XL U9674 ( .A(n9362), .B(ICACHE_addr[17]), .Y(n4688) );
  MX2XL U9675 ( .A(DCACHE_addr[6]), .B(net98952), .S0(n5508), .Y(\i_MIPS/n461 ) );
  MX2XL U9676 ( .A(DCACHE_addr[8]), .B(net99336), .S0(n5510), .Y(\i_MIPS/n459 ) );
  MX2XL U9677 ( .A(DCACHE_addr[11]), .B(n3830), .S0(n5508), .Y(\i_MIPS/n456 )
         );
  MX2XL U9678 ( .A(DCACHE_addr[12]), .B(net99583), .S0(n5506), .Y(
        \i_MIPS/n455 ) );
  MX2XL U9679 ( .A(DCACHE_addr[14]), .B(n3667), .S0(n5506), .Y(\i_MIPS/n453 )
         );
  MX2XL U9680 ( .A(DCACHE_addr[28]), .B(n4727), .S0(n5509), .Y(\i_MIPS/n439 )
         );
  MX2XL U9681 ( .A(DCACHE_addr[5]), .B(net99110), .S0(n5510), .Y(\i_MIPS/n462 ) );
  CLKBUFX3 U9682 ( .A(\i_MIPS/IR_ID[20] ), .Y(net108959) );
  XOR2X4 U9683 ( .A(n11374), .B(\i_MIPS/PC/n19 ), .Y(n4694) );
  MX3XL U9684 ( .A(n8732), .B(n8731), .C(n8733), .S0(n177), .S1(n5590), .Y(
        n8737) );
  OA22XL U9685 ( .A0(net112673), .A1(n1579), .B0(net112571), .B1(n3192), .Y(
        n7733) );
  XOR2X4 U9686 ( .A(n11369), .B(\i_MIPS/PC/n14 ), .Y(n4697) );
  OA22XL U9687 ( .A0(\i_MIPS/Register/register[0][19] ), .A1(n9226), .B0(
        \i_MIPS/Register/register[8][19] ), .B1(n9225), .Y(n7762) );
  CLKMX2X2 U9688 ( .A(\I_cache/cache[7][153] ), .B(n4512), .S0(n5373), .Y(
        n11592) );
  CLKMX2X2 U9689 ( .A(\I_cache/cache[6][153] ), .B(n4512), .S0(n5417), .Y(
        n11593) );
  CLKMX2X2 U9690 ( .A(\I_cache/cache[5][153] ), .B(n4512), .S0(n5283), .Y(
        n11594) );
  CLKMX2X2 U9691 ( .A(\I_cache/cache[4][153] ), .B(n4512), .S0(n5326), .Y(
        n11595) );
  CLKMX2X2 U9692 ( .A(\I_cache/cache[3][153] ), .B(n4512), .S0(n5197), .Y(
        n11596) );
  CLKMX2X2 U9693 ( .A(\I_cache/cache[2][153] ), .B(n4512), .S0(n5239), .Y(
        n11597) );
  CLKMX2X2 U9694 ( .A(\I_cache/cache[1][153] ), .B(n4512), .S0(n5110), .Y(
        n11598) );
  CLKMX2X2 U9695 ( .A(\I_cache/cache[0][153] ), .B(n4512), .S0(n5152), .Y(
        n11599) );
  OA22X1 U9696 ( .A0(\i_MIPS/Register/register[23][24] ), .A1(n4885), .B0(
        \i_MIPS/Register/register[31][24] ), .B1(n4877), .Y(n8945) );
  OA22X1 U9697 ( .A0(\i_MIPS/Register/register[23][28] ), .A1(n4885), .B0(
        \i_MIPS/Register/register[31][28] ), .B1(n4877), .Y(n9033) );
  OA22X1 U9698 ( .A0(\i_MIPS/Register/register[23][20] ), .A1(n4884), .B0(
        \i_MIPS/Register/register[31][20] ), .B1(n4876), .Y(n8570) );
  OA22X1 U9699 ( .A0(\i_MIPS/Register/register[23][23] ), .A1(n4884), .B0(
        \i_MIPS/Register/register[31][23] ), .B1(n4876), .Y(n8238) );
  OA22X1 U9700 ( .A0(\i_MIPS/Register/register[23][22] ), .A1(n4883), .B0(
        \i_MIPS/Register/register[31][22] ), .B1(n4875), .Y(n7997) );
  OA22X1 U9701 ( .A0(\i_MIPS/Register/register[23][16] ), .A1(n4883), .B0(
        \i_MIPS/Register/register[31][16] ), .B1(n4875), .Y(n8180) );
  OA22X1 U9702 ( .A0(\i_MIPS/Register/register[23][2] ), .A1(n4884), .B0(
        \i_MIPS/Register/register[31][2] ), .B1(n4876), .Y(n8836) );
  OA22X1 U9703 ( .A0(\i_MIPS/Register/register[23][3] ), .A1(n4884), .B0(
        \i_MIPS/Register/register[31][3] ), .B1(n4876), .Y(n8751) );
  OA22X1 U9704 ( .A0(\i_MIPS/Register/register[23][13] ), .A1(n4881), .B0(
        \i_MIPS/Register/register[31][13] ), .B1(n4873), .Y(n6404) );
  OA22X1 U9705 ( .A0(\i_MIPS/Register/register[23][26] ), .A1(n4884), .B0(
        \i_MIPS/Register/register[31][26] ), .B1(n4876), .Y(n8373) );
  OA22X1 U9706 ( .A0(\i_MIPS/Register/register[23][25] ), .A1(n4884), .B0(
        \i_MIPS/Register/register[31][25] ), .B1(n4876), .Y(n8465) );
  OA22X1 U9707 ( .A0(\i_MIPS/Register/register[23][17] ), .A1(n4883), .B0(
        \i_MIPS/Register/register[31][17] ), .B1(n4875), .Y(n7745) );
  OA22X1 U9708 ( .A0(\i_MIPS/Register/register[23][10] ), .A1(n4882), .B0(
        \i_MIPS/Register/register[31][10] ), .B1(n4874), .Y(n7220) );
  OA22X1 U9709 ( .A0(\i_MIPS/Register/register[23][11] ), .A1(n4882), .B0(
        \i_MIPS/Register/register[31][11] ), .B1(n4874), .Y(n7130) );
  OA22X1 U9710 ( .A0(\i_MIPS/Register/register[23][4] ), .A1(n4882), .B0(
        \i_MIPS/Register/register[31][4] ), .B1(n4874), .Y(n7382) );
  OA22X1 U9711 ( .A0(\i_MIPS/Register/register[23][9] ), .A1(n4881), .B0(
        \i_MIPS/Register/register[31][9] ), .B1(n4873), .Y(n6895) );
  OA22X1 U9712 ( .A0(\i_MIPS/Register/register[23][8] ), .A1(n4881), .B0(
        \i_MIPS/Register/register[31][8] ), .B1(n4873), .Y(n6812) );
  OA22X1 U9713 ( .A0(net112051), .A1(n1440), .B0(net111927), .B1(n3053), .Y(
        n7059) );
  OA22X1 U9714 ( .A0(net112077), .A1(n1441), .B0(net111953), .B1(n3054), .Y(
        n8859) );
  OA22X1 U9715 ( .A0(net112077), .A1(n1442), .B0(net111953), .B1(n3055), .Y(
        n8851) );
  OA22X1 U9716 ( .A0(net112069), .A1(n1443), .B0(net111945), .B1(n3056), .Y(
        n8292) );
  OA22X1 U9717 ( .A0(net112067), .A1(n1444), .B0(net111943), .B1(n3057), .Y(
        n8195) );
  OA22X1 U9718 ( .A0(net112075), .A1(n1445), .B0(net111951), .B1(n3058), .Y(
        n8677) );
  OA22X1 U9719 ( .A0(net112063), .A1(n1446), .B0(net111939), .B1(n3059), .Y(
        n7811) );
  OA22X1 U9720 ( .A0(net112075), .A1(n1447), .B0(net111951), .B1(n3060), .Y(
        n8673) );
  OA22X1 U9721 ( .A0(net112065), .A1(n1448), .B0(net111941), .B1(n3061), .Y(
        n8021) );
  OA22X1 U9722 ( .A0(net112059), .A1(n1449), .B0(net111935), .B1(n3062), .Y(
        n7633) );
  OA22X1 U9723 ( .A0(net112063), .A1(n1450), .B0(net111939), .B1(n3063), .Y(
        n7916) );
  OA22X1 U9724 ( .A0(net112065), .A1(n1451), .B0(net111941), .B1(n3064), .Y(
        n7920) );
  OA22X1 U9725 ( .A0(net112049), .A1(n1452), .B0(net111925), .B1(n3065), .Y(
        n6968) );
  OA22X1 U9726 ( .A0(net112049), .A1(n1453), .B0(net111925), .B1(n3066), .Y(
        n6876) );
  OA22X1 U9727 ( .A0(net112047), .A1(n1454), .B0(net111923), .B1(n3067), .Y(
        n6868) );
  OA22X1 U9728 ( .A0(net112047), .A1(n1455), .B0(net111923), .B1(n3068), .Y(
        n6793) );
  OA22XL U9729 ( .A0(\i_MIPS/Register/register[4][19] ), .A1(n9224), .B0(
        \i_MIPS/Register/register[12][19] ), .B1(n9223), .Y(n7763) );
  MX2XL U9730 ( .A(\D_cache/cache[6][152] ), .B(n126), .S0(net111989), .Y(
        \D_cache/n574 ) );
  MX2XL U9731 ( .A(\D_cache/cache[5][152] ), .B(n126), .S0(net112123), .Y(
        \D_cache/n575 ) );
  MX2XL U9732 ( .A(\D_cache/cache[4][152] ), .B(n126), .S0(net112195), .Y(
        \D_cache/n576 ) );
  MX2XL U9733 ( .A(\D_cache/cache[3][152] ), .B(n126), .S0(net112285), .Y(
        \D_cache/n577 ) );
  MX2XL U9734 ( .A(\D_cache/cache[2][152] ), .B(n126), .S0(net112409), .Y(
        \D_cache/n578 ) );
  MX2XL U9735 ( .A(\D_cache/cache[1][152] ), .B(n126), .S0(net112533), .Y(
        \D_cache/n579 ) );
  MX2XL U9736 ( .A(\D_cache/cache[0][152] ), .B(n126), .S0(net112635), .Y(
        \D_cache/n580 ) );
  MX2XL U9737 ( .A(\I_cache/cache[5][132] ), .B(n10986), .S0(n5277), .Y(n11762) );
  MX2XL U9738 ( .A(\I_cache/cache[4][132] ), .B(n10986), .S0(n4680), .Y(n11763) );
  MX2XL U9739 ( .A(\I_cache/cache[2][132] ), .B(n10986), .S0(n5242), .Y(n11765) );
  MX2XL U9740 ( .A(\I_cache/cache[0][132] ), .B(n10986), .S0(n5149), .Y(n11767) );
  MX2XL U9741 ( .A(\I_cache/cache[5][128] ), .B(n10978), .S0(n5277), .Y(n11794) );
  MX2XL U9742 ( .A(\I_cache/cache[4][128] ), .B(n10978), .S0(n4680), .Y(n11795) );
  MX2XL U9743 ( .A(\I_cache/cache[2][128] ), .B(n10978), .S0(n5237), .Y(n11797) );
  MX2XL U9744 ( .A(\I_cache/cache[0][128] ), .B(n10978), .S0(n5145), .Y(n11799) );
  OA22X1 U9745 ( .A0(\i_MIPS/Register/register[19][20] ), .A1(n4867), .B0(
        \i_MIPS/Register/register[27][20] ), .B1(n4857), .Y(n8571) );
  OA22X1 U9746 ( .A0(\i_MIPS/Register/register[3][20] ), .A1(n4867), .B0(
        \i_MIPS/Register/register[11][20] ), .B1(n4857), .Y(n8562) );
  OA22X1 U9747 ( .A0(\i_MIPS/Register/register[19][26] ), .A1(n4867), .B0(
        \i_MIPS/Register/register[27][26] ), .B1(n4857), .Y(n8374) );
  OA22X1 U9748 ( .A0(\i_MIPS/Register/register[3][26] ), .A1(n4867), .B0(
        \i_MIPS/Register/register[11][26] ), .B1(n4857), .Y(n8365) );
  OA22X1 U9749 ( .A0(\i_MIPS/Register/register[19][23] ), .A1(n4867), .B0(
        \i_MIPS/Register/register[27][23] ), .B1(n4857), .Y(n8239) );
  OA22X1 U9750 ( .A0(\i_MIPS/Register/register[3][23] ), .A1(n4866), .B0(
        \i_MIPS/Register/register[11][23] ), .B1(n4855), .Y(n8230) );
  OA22X1 U9751 ( .A0(\i_MIPS/Register/register[19][22] ), .A1(n4866), .B0(
        \i_MIPS/Register/register[27][22] ), .B1(n4855), .Y(n7998) );
  OA22X1 U9752 ( .A0(\i_MIPS/Register/register[3][22] ), .A1(n4866), .B0(
        \i_MIPS/Register/register[11][22] ), .B1(n4857), .Y(n7989) );
  OA22X1 U9753 ( .A0(\i_MIPS/Register/register[19][16] ), .A1(n4866), .B0(
        \i_MIPS/Register/register[27][16] ), .B1(n4855), .Y(n8181) );
  OA22X1 U9754 ( .A0(\i_MIPS/Register/register[3][16] ), .A1(n4866), .B0(
        \i_MIPS/Register/register[11][16] ), .B1(n4857), .Y(n8172) );
  OA22X1 U9755 ( .A0(\i_MIPS/Register/register[19][2] ), .A1(n4867), .B0(
        \i_MIPS/Register/register[27][2] ), .B1(n4857), .Y(n8837) );
  OA22X1 U9756 ( .A0(\i_MIPS/Register/register[3][2] ), .A1(n4867), .B0(
        \i_MIPS/Register/register[11][2] ), .B1(n4857), .Y(n8828) );
  OA22X1 U9757 ( .A0(\i_MIPS/Register/register[19][3] ), .A1(n4867), .B0(
        \i_MIPS/Register/register[27][3] ), .B1(n4857), .Y(n8752) );
  OA22X1 U9758 ( .A0(\i_MIPS/Register/register[3][3] ), .A1(n4867), .B0(
        \i_MIPS/Register/register[11][3] ), .B1(n4857), .Y(n8743) );
  OA22X1 U9759 ( .A0(\i_MIPS/Register/register[19][10] ), .A1(n4865), .B0(
        \i_MIPS/Register/register[27][10] ), .B1(n4856), .Y(n7221) );
  OA22X1 U9760 ( .A0(\i_MIPS/Register/register[3][10] ), .A1(n4865), .B0(
        \i_MIPS/Register/register[11][10] ), .B1(n4856), .Y(n7212) );
  OA22X1 U9761 ( .A0(\i_MIPS/Register/register[19][4] ), .A1(n4865), .B0(
        \i_MIPS/Register/register[27][4] ), .B1(n4856), .Y(n7383) );
  OA22X1 U9762 ( .A0(\i_MIPS/Register/register[3][4] ), .A1(n4865), .B0(
        \i_MIPS/Register/register[11][4] ), .B1(n4856), .Y(n7374) );
  OA22X1 U9763 ( .A0(\i_MIPS/Register/register[19][13] ), .A1(n4864), .B0(
        \i_MIPS/Register/register[27][13] ), .B1(n4855), .Y(n6405) );
  OA22X1 U9764 ( .A0(\i_MIPS/Register/register[3][13] ), .A1(n4864), .B0(
        \i_MIPS/Register/register[11][13] ), .B1(n4855), .Y(n6396) );
  OA22X1 U9765 ( .A0(\i_MIPS/Register/register[3][14] ), .A1(n4864), .B0(
        \i_MIPS/Register/register[11][14] ), .B1(n4855), .Y(n6979) );
  OA22X1 U9766 ( .A0(\i_MIPS/Register/register[19][9] ), .A1(n4864), .B0(
        \i_MIPS/Register/register[27][9] ), .B1(n4855), .Y(n6896) );
  OA22X1 U9767 ( .A0(\i_MIPS/Register/register[3][9] ), .A1(n4864), .B0(
        \i_MIPS/Register/register[11][9] ), .B1(n4855), .Y(n6887) );
  OA22X1 U9768 ( .A0(\i_MIPS/Register/register[19][25] ), .A1(n4867), .B0(
        \i_MIPS/Register/register[27][25] ), .B1(n4857), .Y(n8466) );
  OA22X1 U9769 ( .A0(\i_MIPS/Register/register[3][25] ), .A1(n4867), .B0(
        \i_MIPS/Register/register[11][25] ), .B1(n4857), .Y(n8457) );
  OA22X1 U9770 ( .A0(\i_MIPS/Register/register[19][17] ), .A1(n4866), .B0(
        \i_MIPS/Register/register[27][17] ), .B1(n4857), .Y(n7746) );
  OA22X1 U9771 ( .A0(\i_MIPS/Register/register[3][17] ), .A1(n4866), .B0(
        \i_MIPS/Register/register[11][17] ), .B1(n4856), .Y(n7737) );
  OA22X1 U9772 ( .A0(\i_MIPS/Register/register[19][11] ), .A1(n4865), .B0(
        \i_MIPS/Register/register[27][11] ), .B1(n4856), .Y(n7131) );
  OA22X1 U9773 ( .A0(\i_MIPS/Register/register[3][11] ), .A1(n4865), .B0(
        \i_MIPS/Register/register[11][11] ), .B1(n4856), .Y(n7122) );
  OA22X1 U9774 ( .A0(\i_MIPS/Register/register[19][8] ), .A1(n4864), .B0(
        \i_MIPS/Register/register[27][8] ), .B1(n4855), .Y(n6813) );
  OA22X1 U9775 ( .A0(\i_MIPS/Register/register[3][8] ), .A1(n4864), .B0(
        \i_MIPS/Register/register[11][8] ), .B1(n4855), .Y(n6804) );
  OA22X1 U9776 ( .A0(\i_MIPS/Register/register[3][29] ), .A1(n4864), .B0(
        \i_MIPS/Register/register[11][29] ), .B1(n4855), .Y(n6725) );
  OA22X1 U9777 ( .A0(\i_MIPS/Register/register[19][0] ), .A1(n4864), .B0(
        \i_MIPS/Register/register[27][0] ), .B1(n4855), .Y(n6555) );
  OA22X1 U9778 ( .A0(\i_MIPS/Register/register[3][0] ), .A1(n4864), .B0(
        \i_MIPS/Register/register[11][0] ), .B1(n4855), .Y(n6546) );
  AO22X1 U9779 ( .A0(n9118), .A1(n474), .B0(n4900), .B1(n2027), .Y(n9119) );
  AO22X1 U9780 ( .A0(n9118), .A1(n475), .B0(n4901), .B1(n2028), .Y(n9106) );
  AO22X1 U9781 ( .A0(n9118), .A1(n609), .B0(n4901), .B1(n2129), .Y(n6738) );
  AO22X1 U9782 ( .A0(n9118), .A1(n610), .B0(n4901), .B1(n2130), .Y(n6729) );
  AO22X1 U9783 ( .A0(n9118), .A1(n272), .B0(n4899), .B1(n727), .Y(n7299) );
  AO22X1 U9784 ( .A0(n9118), .A1(n681), .B0(n4900), .B1(n2210), .Y(n7507) );
  AO22X1 U9785 ( .A0(n9118), .A1(n273), .B0(n4899), .B1(n728), .Y(n6983) );
  AO22X1 U9786 ( .A0(n9118), .A1(n267), .B0(n4899), .B1(n719), .Y(n7074) );
  AO22X1 U9787 ( .A0(n9118), .A1(n682), .B0(n4900), .B1(n2211), .Y(n7574) );
  AO22X1 U9788 ( .A0(n9118), .A1(n611), .B0(n4901), .B1(n2131), .Y(n6400) );
  AO22X1 U9789 ( .A0(n9118), .A1(n683), .B0(n4901), .B1(n2212), .Y(n6891) );
  AO22X1 U9790 ( .A0(n9118), .A1(n476), .B0(n4901), .B1(n2029), .Y(n6808) );
  AO22X1 U9791 ( .A0(n9118), .A1(n684), .B0(n4901), .B1(n2213), .Y(n6310) );
  AO22X1 U9792 ( .A0(n9118), .A1(n612), .B0(n4900), .B1(n2132), .Y(n8950) );
  AO22X1 U9793 ( .A0(n9118), .A1(n613), .B0(n4900), .B1(n2133), .Y(n8941) );
  AO22X1 U9794 ( .A0(n9118), .A1(n614), .B0(n4902), .B1(n2134), .Y(n8185) );
  AO22X1 U9795 ( .A0(n9118), .A1(n615), .B0(n4902), .B1(n2135), .Y(n8176) );
  AO22X1 U9796 ( .A0(n9118), .A1(n616), .B0(n4902), .B1(n2136), .Y(n8243) );
  AO22X1 U9797 ( .A0(n9118), .A1(n617), .B0(n4902), .B1(n2137), .Y(n8234) );
  AO22X1 U9798 ( .A0(n9118), .A1(n618), .B0(n4902), .B1(n2138), .Y(n8002) );
  AO22X1 U9799 ( .A0(n9118), .A1(n619), .B0(n4902), .B1(n2139), .Y(n7993) );
  AO22X1 U9800 ( .A0(n9118), .A1(n620), .B0(n4900), .B1(n2140), .Y(n8756) );
  AO22X1 U9801 ( .A0(n9118), .A1(n621), .B0(n4900), .B1(n2141), .Y(n8747) );
  AO22X1 U9802 ( .A0(n9118), .A1(n622), .B0(n4902), .B1(n2142), .Y(n8575) );
  AO22X1 U9803 ( .A0(n9118), .A1(n623), .B0(n4900), .B1(n2143), .Y(n8061) );
  AO22X1 U9804 ( .A0(n9118), .A1(n624), .B0(n4902), .B1(n2144), .Y(n8566) );
  AO22X1 U9805 ( .A0(n9118), .A1(n625), .B0(n4900), .B1(n2145), .Y(n8052) );
  AO22X1 U9806 ( .A0(n9118), .A1(n685), .B0(n4902), .B1(n2214), .Y(n7516) );
  AO22X1 U9807 ( .A0(n9118), .A1(n626), .B0(n4900), .B1(n2146), .Y(n8841) );
  AO22X1 U9808 ( .A0(n9118), .A1(n627), .B0(n4899), .B1(n2147), .Y(n8832) );
  AO22X1 U9809 ( .A0(n9118), .A1(n628), .B0(n4901), .B1(n2148), .Y(n6409) );
  AO22X1 U9810 ( .A0(n9118), .A1(n274), .B0(n4899), .B1(n729), .Y(n6992) );
  AO22X1 U9811 ( .A0(n9118), .A1(n686), .B0(n4900), .B1(n2215), .Y(n7583) );
  AO22X1 U9812 ( .A0(n9118), .A1(n275), .B0(n4899), .B1(n730), .Y(n7308) );
  AO22X1 U9813 ( .A0(n9118), .A1(n268), .B0(n4899), .B1(n720), .Y(n7387) );
  AO22X1 U9814 ( .A0(n9118), .A1(n269), .B0(n4899), .B1(n721), .Y(n7378) );
  AO22X1 U9815 ( .A0(n9118), .A1(n687), .B0(n4901), .B1(n2216), .Y(n6900) );
  AO22X1 U9816 ( .A0(n9118), .A1(n629), .B0(n4902), .B1(n2149), .Y(n8378) );
  AO22X1 U9817 ( .A0(n9118), .A1(n630), .B0(n4902), .B1(n2150), .Y(n8369) );
  AO22X1 U9818 ( .A0(n9118), .A1(n276), .B0(n4899), .B1(n731), .Y(n7225) );
  AO22X1 U9819 ( .A0(n9118), .A1(n277), .B0(n4899), .B1(n732), .Y(n7083) );
  AO22X1 U9820 ( .A0(n9118), .A1(n278), .B0(n4899), .B1(n733), .Y(n7216) );
  AO22X1 U9821 ( .A0(n9118), .A1(n631), .B0(n4900), .B1(n2151), .Y(n9038) );
  AO22X1 U9822 ( .A0(n9118), .A1(n477), .B0(n4902), .B1(n2030), .Y(n8470) );
  AO22X1 U9823 ( .A0(n9118), .A1(n632), .B0(n4900), .B1(n2152), .Y(n9029) );
  AO22X1 U9824 ( .A0(n9118), .A1(n478), .B0(n4902), .B1(n2031), .Y(n8461) );
  AO22X1 U9825 ( .A0(n9118), .A1(n479), .B0(n4901), .B1(n2032), .Y(n6817) );
  AO22X1 U9826 ( .A0(n9118), .A1(n270), .B0(n4899), .B1(n722), .Y(n7135) );
  AO22X1 U9827 ( .A0(n9118), .A1(n271), .B0(n4899), .B1(n723), .Y(n7126) );
  AO22X1 U9828 ( .A0(n9118), .A1(n633), .B0(n4902), .B1(n2153), .Y(n8634) );
  AO22X1 U9829 ( .A0(n9118), .A1(n688), .B0(n4902), .B1(n2217), .Y(n7750) );
  AO22X1 U9830 ( .A0(n9118), .A1(n634), .B0(n4902), .B1(n2154), .Y(n8625) );
  AO22X1 U9831 ( .A0(n9118), .A1(n689), .B0(n4900), .B1(n2218), .Y(n7741) );
  AO22X1 U9832 ( .A0(n5002), .A1(n480), .B0(n4998), .B1(n2033), .Y(n8875) );
  AO22X1 U9833 ( .A0(n5002), .A1(n481), .B0(n4998), .B1(n2034), .Y(n8866) );
  AO22X1 U9834 ( .A0(n9118), .A1(n690), .B0(n4900), .B1(n2219), .Y(n7906) );
  AO22X1 U9835 ( .A0(n9118), .A1(n691), .B0(n4900), .B1(n2220), .Y(n7897) );
  AO22X1 U9836 ( .A0(n5002), .A1(n482), .B0(n4997), .B1(n2035), .Y(n7421) );
  AO22X1 U9837 ( .A0(n5001), .A1(n483), .B0(n4997), .B1(n2036), .Y(n8413) );
  AO22X1 U9838 ( .A0(n5001), .A1(n217), .B0(n4998), .B1(n2155), .Y(n6696) );
  AO22X1 U9839 ( .A0(n5002), .A1(n484), .B0(n4997), .B1(n2037), .Y(n7412) );
  AO22X1 U9840 ( .A0(n5001), .A1(n692), .B0(n4997), .B1(n2221), .Y(n8404) );
  AO22X1 U9841 ( .A0(n5001), .A1(n205), .B0(n4996), .B1(n2038), .Y(n6687) );
  OA22XL U9842 ( .A0(n5334), .A1(n1220), .B0(n5291), .B1(n2792), .Y(n9330) );
  OA22XL U9843 ( .A0(n5334), .A1(n1221), .B0(n5299), .B1(n2793), .Y(n9353) );
  OA22XL U9844 ( .A0(n5334), .A1(n1222), .B0(n5299), .B1(n2794), .Y(n9358) );
  OA22X1 U9845 ( .A0(n5337), .A1(n1044), .B0(n5293), .B1(n2616), .Y(n9448) );
  OA22XL U9846 ( .A0(n5334), .A1(n1580), .B0(n5293), .B1(n3193), .Y(n9348) );
  OA22X1 U9847 ( .A0(n5354), .A1(n1045), .B0(n5310), .B1(n2617), .Y(n10232) );
  OA22X1 U9848 ( .A0(n5355), .A1(n1046), .B0(n5311), .B1(n2618), .Y(n10236) );
  OA22X1 U9849 ( .A0(n5344), .A1(n1047), .B0(n5300), .B1(n2619), .Y(n9741) );
  OA22X1 U9850 ( .A0(n5343), .A1(n1048), .B0(n5299), .B1(n2620), .Y(n9708) );
  OA22X1 U9851 ( .A0(n5345), .A1(n1049), .B0(n5301), .B1(n2621), .Y(n9785) );
  OA22X1 U9852 ( .A0(n5348), .A1(n1710), .B0(n5304), .B1(n3394), .Y(n9884) );
  OA22X1 U9853 ( .A0(n5348), .A1(n1711), .B0(n5304), .B1(n3395), .Y(n9894) );
  OA22X1 U9854 ( .A0(n5348), .A1(n1712), .B0(n5304), .B1(n3396), .Y(n9899) );
  OA22X1 U9855 ( .A0(n5348), .A1(n1713), .B0(n5304), .B1(n3397), .Y(n9889) );
  OA22X1 U9856 ( .A0(n5348), .A1(n1714), .B0(n5304), .B1(n3398), .Y(n9908) );
  OA22XL U9857 ( .A0(n5349), .A1(n1800), .B0(n5305), .B1(n3484), .Y(n9918) );
  OA22XL U9858 ( .A0(n5349), .A1(n1801), .B0(n5305), .B1(n3485), .Y(n9923) );
  OA22X1 U9859 ( .A0(n5348), .A1(n1715), .B0(n5304), .B1(n3399), .Y(n9913) );
  OA22X1 U9860 ( .A0(n5347), .A1(n1716), .B0(n5303), .B1(n3400), .Y(n9850) );
  OA22X1 U9861 ( .A0(n5347), .A1(n1717), .B0(n5303), .B1(n3401), .Y(n9855) );
  OA22X1 U9862 ( .A0(n5347), .A1(n1718), .B0(n5303), .B1(n3402), .Y(n9860) );
  OA22X1 U9863 ( .A0(n5347), .A1(n1719), .B0(n5303), .B1(n3403), .Y(n9870) );
  OA22X1 U9864 ( .A0(n5347), .A1(n1720), .B0(n5303), .B1(n3404), .Y(n9875) );
  OA22X1 U9865 ( .A0(n5347), .A1(n1721), .B0(n5303), .B1(n3405), .Y(n9865) );
  OA22X1 U9866 ( .A0(n5351), .A1(n1722), .B0(n5307), .B1(n3406), .Y(n10004) );
  OA22X1 U9867 ( .A0(n5351), .A1(n1723), .B0(n5307), .B1(n3407), .Y(n10014) );
  OA22X1 U9868 ( .A0(n5351), .A1(n1724), .B0(n5307), .B1(n3408), .Y(n10019) );
  OA22X1 U9869 ( .A0(n5351), .A1(n1725), .B0(n5307), .B1(n3409), .Y(n10009) );
  OA22X1 U9870 ( .A0(n5351), .A1(n1726), .B0(n5307), .B1(n3410), .Y(n9990) );
  OA22X1 U9871 ( .A0(n5351), .A1(n1727), .B0(n5307), .B1(n3411), .Y(n10028) );
  OA22X1 U9872 ( .A0(n5352), .A1(n1728), .B0(n5308), .B1(n3412), .Y(n10038) );
  OA22X1 U9873 ( .A0(n5352), .A1(n1729), .B0(n5308), .B1(n3413), .Y(n10043) );
  OA22X1 U9874 ( .A0(n5352), .A1(n1730), .B0(n5308), .B1(n3414), .Y(n10033) );
  OA22X1 U9875 ( .A0(n5352), .A1(n1731), .B0(n5308), .B1(n3415), .Y(n10057) );
  OA22X1 U9876 ( .A0(n5352), .A1(n1732), .B0(n5308), .B1(n3416), .Y(n10067) );
  OA22X1 U9877 ( .A0(n5352), .A1(n1733), .B0(n5308), .B1(n3417), .Y(n10062) );
  OA22X1 U9878 ( .A0(n5353), .A1(n1050), .B0(n5309), .B1(n2622), .Y(n10092) );
  OA22X1 U9879 ( .A0(n5353), .A1(n1051), .B0(n5309), .B1(n2623), .Y(n10082) );
  OA22X1 U9880 ( .A0(\i_MIPS/Register/register[22][25] ), .A1(n4913), .B0(
        \i_MIPS/Register/register[30][25] ), .B1(n4907), .Y(n8469) );
  OA22X1 U9881 ( .A0(\i_MIPS/Register/register[22][22] ), .A1(n4912), .B0(
        \i_MIPS/Register/register[30][22] ), .B1(n4906), .Y(n8001) );
  OA22X1 U9882 ( .A0(\i_MIPS/Register/register[22][10] ), .A1(n4911), .B0(
        \i_MIPS/Register/register[30][10] ), .B1(n4903), .Y(n7224) );
  OA22X1 U9883 ( .A0(\i_MIPS/Register/register[22][2] ), .A1(n4938), .B0(
        \i_MIPS/Register/register[30][2] ), .B1(n4932), .Y(n8874) );
  OA22X1 U9884 ( .A0(\i_MIPS/Register/register[6][2] ), .A1(n4938), .B0(
        \i_MIPS/Register/register[14][2] ), .B1(n4932), .Y(n8865) );
  OA22X1 U9885 ( .A0(\i_MIPS/Register/register[22][4] ), .A1(n4936), .B0(
        \i_MIPS/Register/register[30][4] ), .B1(n4929), .Y(n7420) );
  OA22X1 U9886 ( .A0(\i_MIPS/Register/register[22][22] ), .A1(n4937), .B0(
        \i_MIPS/Register/register[30][22] ), .B1(n4930), .Y(n8036) );
  OA22X1 U9887 ( .A0(\i_MIPS/Register/register[6][22] ), .A1(n4937), .B0(
        \i_MIPS/Register/register[14][22] ), .B1(n4930), .Y(n8027) );
  OA22X2 U9888 ( .A0(net112449), .A1(n977), .B0(net112325), .B1(n2504), .Y(
        n6100) );
  OA22X2 U9889 ( .A0(net112037), .A1(n978), .B0(net111965), .B1(n2505), .Y(
        n6102) );
  OA22X1 U9890 ( .A0(\i_MIPS/Register/register[21][23] ), .A1(n4850), .B0(
        \i_MIPS/Register/register[29][23] ), .B1(n4843), .Y(n8240) );
  OA22X1 U9891 ( .A0(\i_MIPS/Register/register[21][22] ), .A1(n4851), .B0(
        \i_MIPS/Register/register[29][22] ), .B1(n4842), .Y(n7999) );
  OA22X1 U9892 ( .A0(\i_MIPS/Register/register[21][16] ), .A1(n4851), .B0(
        \i_MIPS/Register/register[29][16] ), .B1(n4842), .Y(n8182) );
  OA22X1 U9893 ( .A0(\i_MIPS/Register/register[21][24] ), .A1(n4851), .B0(
        \i_MIPS/Register/register[29][24] ), .B1(n4844), .Y(n8947) );
  OA22X1 U9894 ( .A0(\i_MIPS/Register/register[21][2] ), .A1(n4850), .B0(
        \i_MIPS/Register/register[29][2] ), .B1(n4843), .Y(n8838) );
  OA22X1 U9895 ( .A0(\i_MIPS/Register/register[21][3] ), .A1(n4850), .B0(
        \i_MIPS/Register/register[29][3] ), .B1(n4843), .Y(n8753) );
  OA22X1 U9896 ( .A0(\i_MIPS/Register/register[21][20] ), .A1(n4850), .B0(
        \i_MIPS/Register/register[29][20] ), .B1(n4843), .Y(n8572) );
  OA22X1 U9897 ( .A0(\i_MIPS/Register/register[21][26] ), .A1(n4850), .B0(
        \i_MIPS/Register/register[29][26] ), .B1(n4843), .Y(n8375) );
  OA22X1 U9898 ( .A0(\i_MIPS/Register/register[21][25] ), .A1(n4850), .B0(
        \i_MIPS/Register/register[29][25] ), .B1(n4843), .Y(n8467) );
  OA22X1 U9899 ( .A0(\i_MIPS/Register/register[21][28] ), .A1(n4851), .B0(
        \i_MIPS/Register/register[29][28] ), .B1(n4844), .Y(n9035) );
  OA22X1 U9900 ( .A0(\i_MIPS/Register/register[21][17] ), .A1(n4850), .B0(
        \i_MIPS/Register/register[29][17] ), .B1(n4842), .Y(n7747) );
  OA22X1 U9901 ( .A0(\i_MIPS/Register/register[21][10] ), .A1(n4849), .B0(
        \i_MIPS/Register/register[29][10] ), .B1(n4841), .Y(n7222) );
  OA22X1 U9902 ( .A0(\i_MIPS/Register/register[21][11] ), .A1(n4849), .B0(
        \i_MIPS/Register/register[29][11] ), .B1(n4841), .Y(n7132) );
  OA22X1 U9903 ( .A0(\i_MIPS/Register/register[21][4] ), .A1(n4849), .B0(
        \i_MIPS/Register/register[29][4] ), .B1(n4841), .Y(n7384) );
  OA22X1 U9904 ( .A0(\i_MIPS/Register/register[21][13] ), .A1(n4848), .B0(
        \i_MIPS/Register/register[29][13] ), .B1(n4843), .Y(n6406) );
  OA22X1 U9905 ( .A0(\i_MIPS/Register/register[21][9] ), .A1(n4848), .B0(
        \i_MIPS/Register/register[29][9] ), .B1(n4843), .Y(n6897) );
  OA22X1 U9906 ( .A0(\i_MIPS/Register/register[21][8] ), .A1(n4848), .B0(
        \i_MIPS/Register/register[29][8] ), .B1(n4844), .Y(n6814) );
  AO22X1 U9907 ( .A0(n4895), .A1(n635), .B0(n4891), .B1(n2156), .Y(n6739) );
  AO22X1 U9908 ( .A0(n4895), .A1(n636), .B0(n4891), .B1(n2157), .Y(n6730) );
  AO22X1 U9909 ( .A0(n4896), .A1(n693), .B0(n4892), .B1(n2222), .Y(n7300) );
  AO22X1 U9910 ( .A0(n4897), .A1(n694), .B0(n4894), .B1(n2223), .Y(n7508) );
  AO22X1 U9911 ( .A0(n4897), .A1(n695), .B0(n4891), .B1(n2224), .Y(n7575) );
  AO22X1 U9912 ( .A0(n4896), .A1(n637), .B0(n4892), .B1(n2158), .Y(n7075) );
  AO22X1 U9913 ( .A0(n4895), .A1(n638), .B0(n4891), .B1(n2159), .Y(n6401) );
  AO22X1 U9914 ( .A0(n4895), .A1(n696), .B0(n4891), .B1(n2225), .Y(n6892) );
  AO22X1 U9915 ( .A0(n4898), .A1(n639), .B0(n4894), .B1(n2160), .Y(n8942) );
  AO22X1 U9916 ( .A0(n4895), .A1(n697), .B0(n4891), .B1(n2226), .Y(n6311) );
  AO22X1 U9917 ( .A0(n4897), .A1(n640), .B0(n4889), .B1(n2161), .Y(n7994) );
  AO22X1 U9918 ( .A0(n4896), .A1(n641), .B0(n4894), .B1(n2162), .Y(n8748) );
  AO22X1 U9919 ( .A0(n4897), .A1(n642), .B0(n4893), .B1(n2163), .Y(n8053) );
  AO22X1 U9920 ( .A0(n4898), .A1(n643), .B0(n4894), .B1(n2164), .Y(n8833) );
  AO22X1 U9921 ( .A0(n4896), .A1(n644), .B0(n4892), .B1(n2165), .Y(n7379) );
  AO22X1 U9922 ( .A0(n4896), .A1(n698), .B0(n4892), .B1(n2227), .Y(n7217) );
  AO22X1 U9923 ( .A0(n4898), .A1(n645), .B0(n4894), .B1(n2166), .Y(n9030) );
  AO22X1 U9924 ( .A0(n4896), .A1(n699), .B0(n4892), .B1(n2228), .Y(n7127) );
  AO22X1 U9925 ( .A0(n4898), .A1(n646), .B0(n4893), .B1(n2167), .Y(n8626) );
  AO22X1 U9926 ( .A0(n4897), .A1(n700), .B0(n4894), .B1(n2229), .Y(n7742) );
  AO22X1 U9927 ( .A0(n4897), .A1(n701), .B0(n4891), .B1(n2230), .Y(n7898) );
  MX2XL U9928 ( .A(\D_cache/cache[6][127] ), .B(n11211), .S0(net111991), .Y(
        \D_cache/n774 ) );
  MX2XL U9929 ( .A(\D_cache/cache[5][127] ), .B(n11211), .S0(net112131), .Y(
        \D_cache/n775 ) );
  MX2XL U9930 ( .A(\D_cache/cache[4][127] ), .B(n11211), .S0(net112211), .Y(
        \D_cache/n776 ) );
  MX2XL U9931 ( .A(\D_cache/cache[3][127] ), .B(n11211), .S0(net112295), .Y(
        \D_cache/n777 ) );
  MX2XL U9932 ( .A(\D_cache/cache[2][127] ), .B(n11211), .S0(net112419), .Y(
        \D_cache/n778 ) );
  MX2XL U9933 ( .A(\D_cache/cache[1][127] ), .B(n11211), .S0(net112543), .Y(
        \D_cache/n779 ) );
  MX2XL U9934 ( .A(\D_cache/cache[0][127] ), .B(n11211), .S0(net112645), .Y(
        \D_cache/n780 ) );
  MX2XL U9935 ( .A(\D_cache/cache[6][63] ), .B(n11208), .S0(net111991), .Y(
        \D_cache/n1286 ) );
  MX2XL U9936 ( .A(\D_cache/cache[5][63] ), .B(n11208), .S0(net112131), .Y(
        \D_cache/n1287 ) );
  MX2XL U9937 ( .A(\D_cache/cache[4][63] ), .B(n11208), .S0(net112211), .Y(
        \D_cache/n1288 ) );
  MX2XL U9938 ( .A(\D_cache/cache[3][63] ), .B(n11208), .S0(net112295), .Y(
        \D_cache/n1289 ) );
  MX2XL U9939 ( .A(\D_cache/cache[2][63] ), .B(n11208), .S0(net112419), .Y(
        \D_cache/n1290 ) );
  MX2XL U9940 ( .A(\D_cache/cache[1][63] ), .B(n11208), .S0(net112543), .Y(
        \D_cache/n1291 ) );
  MX2XL U9941 ( .A(\D_cache/cache[0][63] ), .B(n11208), .S0(net112645), .Y(
        \D_cache/n1292 ) );
  MX2XL U9942 ( .A(\D_cache/cache[6][31] ), .B(n4231), .S0(net111993), .Y(
        \D_cache/n1542 ) );
  MX2XL U9943 ( .A(\D_cache/cache[5][31] ), .B(n4231), .S0(net112131), .Y(
        \D_cache/n1543 ) );
  MX2XL U9944 ( .A(\D_cache/cache[4][31] ), .B(n4231), .S0(net112211), .Y(
        \D_cache/n1544 ) );
  MX2XL U9945 ( .A(\D_cache/cache[3][31] ), .B(n4231), .S0(net112295), .Y(
        \D_cache/n1545 ) );
  MX2XL U9946 ( .A(\D_cache/cache[2][31] ), .B(n4231), .S0(net112419), .Y(
        \D_cache/n1546 ) );
  MX2XL U9947 ( .A(\D_cache/cache[1][31] ), .B(n4231), .S0(net112543), .Y(
        \D_cache/n1547 ) );
  MX2XL U9948 ( .A(\D_cache/cache[0][31] ), .B(n4231), .S0(net112645), .Y(
        \D_cache/n1548 ) );
  MX2XL U9949 ( .A(\D_cache/cache[6][62] ), .B(n4266), .S0(net112009), .Y(
        \D_cache/n1294 ) );
  MX2XL U9950 ( .A(\D_cache/cache[5][62] ), .B(n4266), .S0(net112123), .Y(
        \D_cache/n1295 ) );
  MX2XL U9951 ( .A(\D_cache/cache[4][62] ), .B(n4266), .S0(net112215), .Y(
        \D_cache/n1296 ) );
  MX2XL U9952 ( .A(\D_cache/cache[3][62] ), .B(n4266), .S0(net112295), .Y(
        \D_cache/n1297 ) );
  MX2XL U9953 ( .A(\D_cache/cache[2][62] ), .B(n4266), .S0(net112419), .Y(
        \D_cache/n1298 ) );
  MX2XL U9954 ( .A(\D_cache/cache[1][62] ), .B(n4266), .S0(net112545), .Y(
        \D_cache/n1299 ) );
  MX2XL U9955 ( .A(\D_cache/cache[0][62] ), .B(n4266), .S0(net112647), .Y(
        \D_cache/n1300 ) );
  MX2XL U9956 ( .A(\D_cache/cache[6][61] ), .B(n4267), .S0(net111991), .Y(
        \D_cache/n1302 ) );
  MX2XL U9957 ( .A(\D_cache/cache[5][61] ), .B(n4267), .S0(net112115), .Y(
        \D_cache/n1303 ) );
  MX2XL U9958 ( .A(\D_cache/cache[4][61] ), .B(n4267), .S0(net112197), .Y(
        \D_cache/n1304 ) );
  MX2XL U9959 ( .A(\D_cache/cache[3][61] ), .B(n4267), .S0(net112279), .Y(
        \D_cache/n1305 ) );
  MX2XL U9960 ( .A(\D_cache/cache[2][61] ), .B(n4267), .S0(net112403), .Y(
        \D_cache/n1306 ) );
  MX2XL U9961 ( .A(\D_cache/cache[1][61] ), .B(n4267), .S0(net112527), .Y(
        \D_cache/n1307 ) );
  MX2XL U9962 ( .A(\D_cache/cache[0][61] ), .B(n4267), .S0(net112629), .Y(
        \D_cache/n1308 ) );
  MX2XL U9963 ( .A(\D_cache/cache[6][60] ), .B(n10400), .S0(net111995), .Y(
        \D_cache/n1310 ) );
  MX2XL U9964 ( .A(\D_cache/cache[5][60] ), .B(n10400), .S0(net112119), .Y(
        \D_cache/n1311 ) );
  MX2XL U9965 ( .A(\D_cache/cache[4][60] ), .B(n10400), .S0(net112201), .Y(
        \D_cache/n1312 ) );
  MX2XL U9966 ( .A(\D_cache/cache[3][60] ), .B(n10400), .S0(net112283), .Y(
        \D_cache/n1313 ) );
  MX2XL U9967 ( .A(\D_cache/cache[2][60] ), .B(n10400), .S0(net112403), .Y(
        \D_cache/n1314 ) );
  MX2XL U9968 ( .A(\D_cache/cache[1][60] ), .B(n10400), .S0(net112531), .Y(
        \D_cache/n1315 ) );
  MX2XL U9969 ( .A(\D_cache/cache[0][60] ), .B(n10400), .S0(net112633), .Y(
        \D_cache/n1316 ) );
  MX2XL U9970 ( .A(\D_cache/cache[6][59] ), .B(n4268), .S0(net111999), .Y(
        \D_cache/n1318 ) );
  MX2XL U9971 ( .A(\D_cache/cache[5][59] ), .B(n4268), .S0(net112121), .Y(
        \D_cache/n1319 ) );
  MX2XL U9972 ( .A(\D_cache/cache[4][59] ), .B(n4268), .S0(net112215), .Y(
        \D_cache/n1320 ) );
  MX2XL U9973 ( .A(\D_cache/cache[3][59] ), .B(n4268), .S0(net112281), .Y(
        \D_cache/n1321 ) );
  MX2XL U9974 ( .A(\D_cache/cache[2][59] ), .B(n4268), .S0(net112411), .Y(
        \D_cache/n1322 ) );
  MX2XL U9975 ( .A(\D_cache/cache[1][59] ), .B(n4268), .S0(net112527), .Y(
        \D_cache/n1323 ) );
  MX2XL U9976 ( .A(\D_cache/cache[0][59] ), .B(n4268), .S0(net112629), .Y(
        \D_cache/n1324 ) );
  MX2XL U9977 ( .A(\D_cache/cache[6][58] ), .B(n4269), .S0(net111995), .Y(
        \D_cache/n1326 ) );
  MX2XL U9978 ( .A(\D_cache/cache[5][58] ), .B(n4269), .S0(net112119), .Y(
        \D_cache/n1327 ) );
  MX2XL U9979 ( .A(\D_cache/cache[4][58] ), .B(n4269), .S0(net112201), .Y(
        \D_cache/n1328 ) );
  MX2XL U9980 ( .A(\D_cache/cache[3][58] ), .B(n4269), .S0(net112283), .Y(
        \D_cache/n1329 ) );
  MX2XL U9981 ( .A(\D_cache/cache[2][58] ), .B(n4269), .S0(net112411), .Y(
        \D_cache/n1330 ) );
  MX2XL U9982 ( .A(\D_cache/cache[1][58] ), .B(n4269), .S0(net112531), .Y(
        \D_cache/n1331 ) );
  MX2XL U9983 ( .A(\D_cache/cache[0][58] ), .B(n4269), .S0(net112631), .Y(
        \D_cache/n1332 ) );
  MX2XL U9984 ( .A(\D_cache/cache[6][57] ), .B(n4270), .S0(net111989), .Y(
        \D_cache/n1334 ) );
  MX2XL U9985 ( .A(\D_cache/cache[5][57] ), .B(n4270), .S0(net112113), .Y(
        \D_cache/n1335 ) );
  MX2XL U9986 ( .A(\D_cache/cache[4][57] ), .B(n4270), .S0(net112195), .Y(
        \D_cache/n1336 ) );
  MX2XL U9987 ( .A(\D_cache/cache[3][57] ), .B(n4270), .S0(net112277), .Y(
        \D_cache/n1337 ) );
  MX2XL U9988 ( .A(\D_cache/cache[2][57] ), .B(n4270), .S0(net112401), .Y(
        \D_cache/n1338 ) );
  MX2XL U9989 ( .A(\D_cache/cache[1][57] ), .B(n4270), .S0(net112525), .Y(
        \D_cache/n1339 ) );
  MX2XL U9990 ( .A(\D_cache/cache[0][57] ), .B(n4270), .S0(net112627), .Y(
        \D_cache/n1340 ) );
  MX2XL U9991 ( .A(\D_cache/cache[6][56] ), .B(n10574), .S0(net112003), .Y(
        \D_cache/n1342 ) );
  MX2XL U9992 ( .A(\D_cache/cache[5][56] ), .B(n10574), .S0(net112127), .Y(
        \D_cache/n1343 ) );
  MX2XL U9993 ( .A(\D_cache/cache[4][56] ), .B(n10574), .S0(net112211), .Y(
        \D_cache/n1344 ) );
  MX2XL U9994 ( .A(\D_cache/cache[3][56] ), .B(n10574), .S0(net112291), .Y(
        \D_cache/n1345 ) );
  MX2XL U9995 ( .A(\D_cache/cache[2][56] ), .B(n10574), .S0(net112415), .Y(
        \D_cache/n1346 ) );
  MX2XL U9996 ( .A(\D_cache/cache[1][56] ), .B(n10574), .S0(net112539), .Y(
        \D_cache/n1347 ) );
  MX2XL U9997 ( .A(\D_cache/cache[0][56] ), .B(n10574), .S0(net112641), .Y(
        \D_cache/n1348 ) );
  MX2XL U9998 ( .A(\D_cache/cache[6][55] ), .B(n4271), .S0(net112009), .Y(
        \D_cache/n1350 ) );
  MX2XL U9999 ( .A(\D_cache/cache[5][55] ), .B(n4271), .S0(net112125), .Y(
        \D_cache/n1351 ) );
  MX2XL U10000 ( .A(\D_cache/cache[4][55] ), .B(n4271), .S0(net112211), .Y(
        \D_cache/n1352 ) );
  MX2XL U10001 ( .A(\D_cache/cache[3][55] ), .B(n4271), .S0(net112289), .Y(
        \D_cache/n1353 ) );
  MX2XL U10002 ( .A(\D_cache/cache[2][55] ), .B(n4271), .S0(net112401), .Y(
        \D_cache/n1354 ) );
  MX2XL U10003 ( .A(\D_cache/cache[1][55] ), .B(n4271), .S0(net112537), .Y(
        \D_cache/n1355 ) );
  MX2XL U10004 ( .A(\D_cache/cache[0][55] ), .B(n4271), .S0(net112639), .Y(
        \D_cache/n1356 ) );
  MX2XL U10005 ( .A(\D_cache/cache[6][54] ), .B(n10549), .S0(net112005), .Y(
        \D_cache/n1358 ) );
  MX2XL U10006 ( .A(\D_cache/cache[5][54] ), .B(n10549), .S0(net112125), .Y(
        \D_cache/n1359 ) );
  MX2XL U10007 ( .A(\D_cache/cache[4][54] ), .B(n10549), .S0(net112211), .Y(
        \D_cache/n1360 ) );
  MX2XL U10008 ( .A(\D_cache/cache[3][54] ), .B(n10549), .S0(net112289), .Y(
        \D_cache/n1361 ) );
  MX2XL U10009 ( .A(\D_cache/cache[2][54] ), .B(n10549), .S0(net112415), .Y(
        \D_cache/n1362 ) );
  MX2XL U10010 ( .A(\D_cache/cache[1][54] ), .B(n10549), .S0(net112537), .Y(
        \D_cache/n1363 ) );
  MX2XL U10011 ( .A(\D_cache/cache[0][54] ), .B(n10549), .S0(net112639), .Y(
        \D_cache/n1364 ) );
  MX2XL U10012 ( .A(\D_cache/cache[6][53] ), .B(n4272), .S0(net111995), .Y(
        \D_cache/n1366 ) );
  MX2XL U10013 ( .A(\D_cache/cache[5][53] ), .B(n4272), .S0(net112125), .Y(
        \D_cache/n1367 ) );
  MX2XL U10014 ( .A(\D_cache/cache[4][53] ), .B(n4272), .S0(net112211), .Y(
        \D_cache/n1368 ) );
  MX2XL U10015 ( .A(\D_cache/cache[3][53] ), .B(n4272), .S0(net112289), .Y(
        \D_cache/n1369 ) );
  MX2XL U10016 ( .A(\D_cache/cache[2][53] ), .B(n4272), .S0(net112415), .Y(
        \D_cache/n1370 ) );
  MX2XL U10017 ( .A(\D_cache/cache[1][53] ), .B(n4272), .S0(net112537), .Y(
        \D_cache/n1371 ) );
  MX2XL U10018 ( .A(\D_cache/cache[0][53] ), .B(n4272), .S0(net112639), .Y(
        \D_cache/n1372 ) );
  MX2XL U10019 ( .A(\D_cache/cache[6][52] ), .B(n4273), .S0(net111991), .Y(
        \D_cache/n1374 ) );
  MX2XL U10020 ( .A(\D_cache/cache[5][52] ), .B(n4273), .S0(net112115), .Y(
        \D_cache/n1375 ) );
  MX2XL U10021 ( .A(\D_cache/cache[4][52] ), .B(n4273), .S0(net112197), .Y(
        \D_cache/n1376 ) );
  MX2XL U10022 ( .A(\D_cache/cache[3][52] ), .B(n4273), .S0(net112279), .Y(
        \D_cache/n1377 ) );
  MX2XL U10023 ( .A(\D_cache/cache[2][52] ), .B(n4273), .S0(net112403), .Y(
        \D_cache/n1378 ) );
  MX2XL U10024 ( .A(\D_cache/cache[1][52] ), .B(n4273), .S0(net112527), .Y(
        \D_cache/n1379 ) );
  MX2XL U10025 ( .A(\D_cache/cache[0][52] ), .B(n4273), .S0(net112629), .Y(
        \D_cache/n1380 ) );
  MX2XL U10026 ( .A(\D_cache/cache[6][51] ), .B(n4274), .S0(net111993), .Y(
        \D_cache/n1382 ) );
  MX2XL U10027 ( .A(\D_cache/cache[5][51] ), .B(n4274), .S0(net112117), .Y(
        \D_cache/n1383 ) );
  MX2XL U10028 ( .A(\D_cache/cache[4][51] ), .B(n4274), .S0(net112199), .Y(
        \D_cache/n1384 ) );
  MX2XL U10029 ( .A(\D_cache/cache[3][51] ), .B(n4274), .S0(net112281), .Y(
        \D_cache/n1385 ) );
  MX2XL U10030 ( .A(\D_cache/cache[2][51] ), .B(n4274), .S0(net112405), .Y(
        \D_cache/n1386 ) );
  MX2XL U10031 ( .A(\D_cache/cache[1][51] ), .B(n4274), .S0(net112529), .Y(
        \D_cache/n1387 ) );
  MX2XL U10032 ( .A(\D_cache/cache[0][51] ), .B(n4274), .S0(net112631), .Y(
        \D_cache/n1388 ) );
  MX2XL U10033 ( .A(\D_cache/cache[6][50] ), .B(n10613), .S0(net111999), .Y(
        \D_cache/n1390 ) );
  MX2XL U10034 ( .A(\D_cache/cache[5][50] ), .B(n10613), .S0(net112121), .Y(
        \D_cache/n1391 ) );
  MX2XL U10035 ( .A(\D_cache/cache[4][50] ), .B(n10613), .S0(net112197), .Y(
        \D_cache/n1392 ) );
  MX2XL U10036 ( .A(\D_cache/cache[3][50] ), .B(n10613), .S0(net112285), .Y(
        \D_cache/n1393 ) );
  MX2XL U10037 ( .A(\D_cache/cache[2][50] ), .B(n10613), .S0(net112409), .Y(
        \D_cache/n1394 ) );
  MX2XL U10038 ( .A(\D_cache/cache[1][50] ), .B(n10613), .S0(net112533), .Y(
        \D_cache/n1395 ) );
  MX2XL U10039 ( .A(\D_cache/cache[0][50] ), .B(n10613), .S0(net112635), .Y(
        \D_cache/n1396 ) );
  MX2XL U10040 ( .A(\D_cache/cache[6][49] ), .B(n10600), .S0(net112003), .Y(
        \D_cache/n1398 ) );
  MX2XL U10041 ( .A(\D_cache/cache[5][49] ), .B(n10600), .S0(net112127), .Y(
        \D_cache/n1399 ) );
  MX2XL U10042 ( .A(\D_cache/cache[4][49] ), .B(n10600), .S0(net112199), .Y(
        \D_cache/n1400 ) );
  MX2XL U10043 ( .A(\D_cache/cache[3][49] ), .B(n10600), .S0(net112291), .Y(
        \D_cache/n1401 ) );
  MX2XL U10044 ( .A(\D_cache/cache[2][49] ), .B(n10600), .S0(net112415), .Y(
        \D_cache/n1402 ) );
  MX2XL U10045 ( .A(\D_cache/cache[1][49] ), .B(n10600), .S0(net112539), .Y(
        \D_cache/n1403 ) );
  MX2XL U10046 ( .A(\D_cache/cache[0][49] ), .B(n10600), .S0(net112641), .Y(
        \D_cache/n1404 ) );
  MX2XL U10047 ( .A(\D_cache/cache[6][48] ), .B(n4275), .S0(net111989), .Y(
        \D_cache/n1406 ) );
  MX2XL U10048 ( .A(\D_cache/cache[5][48] ), .B(n4275), .S0(net112113), .Y(
        \D_cache/n1407 ) );
  MX2XL U10049 ( .A(\D_cache/cache[4][48] ), .B(n4275), .S0(net112195), .Y(
        \D_cache/n1408 ) );
  MX2XL U10050 ( .A(\D_cache/cache[3][48] ), .B(n4275), .S0(net112277), .Y(
        \D_cache/n1409 ) );
  MX2XL U10051 ( .A(\D_cache/cache[2][48] ), .B(n4275), .S0(net112405), .Y(
        \D_cache/n1410 ) );
  MX2XL U10052 ( .A(\D_cache/cache[1][48] ), .B(n4275), .S0(net112525), .Y(
        \D_cache/n1411 ) );
  MX2XL U10053 ( .A(\D_cache/cache[0][48] ), .B(n4275), .S0(net112627), .Y(
        \D_cache/n1412 ) );
  MX2XL U10054 ( .A(\D_cache/cache[6][47] ), .B(n4276), .S0(net111995), .Y(
        \D_cache/n1414 ) );
  MX2XL U10055 ( .A(\D_cache/cache[5][47] ), .B(n4276), .S0(net112119), .Y(
        \D_cache/n1415 ) );
  MX2XL U10056 ( .A(\D_cache/cache[4][47] ), .B(n4276), .S0(net112201), .Y(
        \D_cache/n1416 ) );
  MX2XL U10057 ( .A(\D_cache/cache[3][47] ), .B(n4276), .S0(net112283), .Y(
        \D_cache/n1417 ) );
  MX2XL U10058 ( .A(\D_cache/cache[2][47] ), .B(n4276), .S0(net112403), .Y(
        \D_cache/n1418 ) );
  MX2XL U10059 ( .A(\D_cache/cache[1][47] ), .B(n4276), .S0(net112531), .Y(
        \D_cache/n1419 ) );
  MX2XL U10060 ( .A(\D_cache/cache[0][47] ), .B(n4276), .S0(net112633), .Y(
        \D_cache/n1420 ) );
  MX2XL U10061 ( .A(\D_cache/cache[6][46] ), .B(n4277), .S0(net111989), .Y(
        \D_cache/n1422 ) );
  MX2XL U10062 ( .A(\D_cache/cache[5][46] ), .B(n4277), .S0(net112113), .Y(
        \D_cache/n1423 ) );
  MX2XL U10063 ( .A(\D_cache/cache[4][46] ), .B(n4277), .S0(net112195), .Y(
        \D_cache/n1424 ) );
  MX2XL U10064 ( .A(\D_cache/cache[3][46] ), .B(n4277), .S0(net112277), .Y(
        \D_cache/n1425 ) );
  MX2XL U10065 ( .A(\D_cache/cache[2][46] ), .B(n4277), .S0(net112401), .Y(
        \D_cache/n1426 ) );
  MX2XL U10066 ( .A(\D_cache/cache[1][46] ), .B(n4277), .S0(net112525), .Y(
        \D_cache/n1427 ) );
  MX2XL U10067 ( .A(\D_cache/cache[0][46] ), .B(n4277), .S0(net112627), .Y(
        \D_cache/n1428 ) );
  MX2XL U10068 ( .A(\D_cache/cache[6][42] ), .B(n10588), .S0(net112003), .Y(
        \D_cache/n1454 ) );
  MX2XL U10069 ( .A(\D_cache/cache[5][42] ), .B(n10588), .S0(net112127), .Y(
        \D_cache/n1455 ) );
  MX2XL U10070 ( .A(\D_cache/cache[4][42] ), .B(n10588), .S0(net112201), .Y(
        \D_cache/n1456 ) );
  MX2XL U10071 ( .A(\D_cache/cache[3][42] ), .B(n10588), .S0(net112291), .Y(
        \D_cache/n1457 ) );
  MX2XL U10072 ( .A(\D_cache/cache[2][42] ), .B(n10588), .S0(net112415), .Y(
        \D_cache/n1458 ) );
  MX2XL U10073 ( .A(\D_cache/cache[1][42] ), .B(n10588), .S0(net112539), .Y(
        \D_cache/n1459 ) );
  MX2XL U10074 ( .A(\D_cache/cache[0][42] ), .B(n10588), .S0(net112641), .Y(
        \D_cache/n1460 ) );
  MX2XL U10075 ( .A(\D_cache/cache[6][41] ), .B(n4278), .S0(net112011), .Y(
        \D_cache/n1462 ) );
  MX2XL U10076 ( .A(\D_cache/cache[5][41] ), .B(n4278), .S0(net112121), .Y(
        \D_cache/n1463 ) );
  MX2XL U10077 ( .A(\D_cache/cache[3][41] ), .B(n4278), .S0(net112291), .Y(
        \D_cache/n1465 ) );
  MX2XL U10078 ( .A(\D_cache/cache[2][41] ), .B(n4278), .S0(net112423), .Y(
        \D_cache/n1466 ) );
  MX2XL U10079 ( .A(\D_cache/cache[1][41] ), .B(n4278), .S0(net112547), .Y(
        \D_cache/n1467 ) );
  MX2XL U10080 ( .A(\D_cache/cache[0][41] ), .B(n4278), .S0(net112649), .Y(
        \D_cache/n1468 ) );
  MX2XL U10081 ( .A(\D_cache/cache[6][39] ), .B(n4279), .S0(net112009), .Y(
        \D_cache/n1478 ) );
  MX2XL U10082 ( .A(\D_cache/cache[5][39] ), .B(n4279), .S0(net112121), .Y(
        \D_cache/n1479 ) );
  MX2XL U10083 ( .A(\D_cache/cache[4][39] ), .B(n4279), .S0(net112215), .Y(
        \D_cache/n1480 ) );
  MX2XL U10084 ( .A(\D_cache/cache[3][39] ), .B(n4279), .S0(net112293), .Y(
        \D_cache/n1481 ) );
  MX2XL U10085 ( .A(\D_cache/cache[2][39] ), .B(n4279), .S0(net112417), .Y(
        \D_cache/n1482 ) );
  MX2XL U10086 ( .A(\D_cache/cache[1][39] ), .B(n4279), .S0(net112545), .Y(
        \D_cache/n1483 ) );
  MX2XL U10087 ( .A(\D_cache/cache[0][39] ), .B(n4279), .S0(net112647), .Y(
        \D_cache/n1484 ) );
  MX2XL U10088 ( .A(\D_cache/cache[6][38] ), .B(n4249), .S0(net111993), .Y(
        \D_cache/n1486 ) );
  MX2XL U10089 ( .A(\D_cache/cache[5][38] ), .B(n4249), .S0(net112117), .Y(
        \D_cache/n1487 ) );
  MX2XL U10090 ( .A(\D_cache/cache[4][38] ), .B(n4249), .S0(net112199), .Y(
        \D_cache/n1488 ) );
  MX2XL U10091 ( .A(\D_cache/cache[3][38] ), .B(n4249), .S0(net112281), .Y(
        \D_cache/n1489 ) );
  MX2XL U10092 ( .A(\D_cache/cache[2][38] ), .B(n4249), .S0(net112401), .Y(
        \D_cache/n1490 ) );
  MX2XL U10093 ( .A(\D_cache/cache[1][38] ), .B(n4249), .S0(net112529), .Y(
        \D_cache/n1491 ) );
  MX2XL U10094 ( .A(\D_cache/cache[0][38] ), .B(n4249), .S0(net112631), .Y(
        \D_cache/n1492 ) );
  MX2XL U10095 ( .A(\D_cache/cache[6][37] ), .B(n4280), .S0(net111989), .Y(
        \D_cache/n1494 ) );
  MX2XL U10096 ( .A(\D_cache/cache[5][37] ), .B(n4280), .S0(net112113), .Y(
        \D_cache/n1495 ) );
  MX2XL U10097 ( .A(\D_cache/cache[4][37] ), .B(n4280), .S0(net112195), .Y(
        \D_cache/n1496 ) );
  MX2XL U10098 ( .A(\D_cache/cache[3][37] ), .B(n4280), .S0(net112277), .Y(
        \D_cache/n1497 ) );
  MX2XL U10099 ( .A(\D_cache/cache[2][37] ), .B(n4280), .S0(net112401), .Y(
        \D_cache/n1498 ) );
  MX2XL U10100 ( .A(\D_cache/cache[1][37] ), .B(n4280), .S0(net112525), .Y(
        \D_cache/n1499 ) );
  MX2XL U10101 ( .A(\D_cache/cache[0][37] ), .B(n4280), .S0(net112627), .Y(
        \D_cache/n1500 ) );
  MX2XL U10102 ( .A(\D_cache/cache[6][36] ), .B(n4250), .S0(net111993), .Y(
        \D_cache/n1502 ) );
  MX2XL U10103 ( .A(\D_cache/cache[5][36] ), .B(n4250), .S0(net112117), .Y(
        \D_cache/n1503 ) );
  MX2XL U10104 ( .A(\D_cache/cache[4][36] ), .B(n4250), .S0(net112199), .Y(
        \D_cache/n1504 ) );
  MX2XL U10105 ( .A(\D_cache/cache[3][36] ), .B(n4250), .S0(net112281), .Y(
        \D_cache/n1505 ) );
  MX2XL U10106 ( .A(\D_cache/cache[2][36] ), .B(n4250), .S0(net112401), .Y(
        \D_cache/n1506 ) );
  MX2XL U10107 ( .A(\D_cache/cache[1][36] ), .B(n4250), .S0(net112529), .Y(
        \D_cache/n1507 ) );
  MX2XL U10108 ( .A(\D_cache/cache[0][36] ), .B(n4250), .S0(net112631), .Y(
        \D_cache/n1508 ) );
  MX2XL U10109 ( .A(\D_cache/cache[6][35] ), .B(n4281), .S0(net111991), .Y(
        \D_cache/n1510 ) );
  MX2XL U10110 ( .A(\D_cache/cache[5][35] ), .B(n4281), .S0(net112115), .Y(
        \D_cache/n1511 ) );
  MX2XL U10111 ( .A(\D_cache/cache[4][35] ), .B(n4281), .S0(net112197), .Y(
        \D_cache/n1512 ) );
  MX2XL U10112 ( .A(\D_cache/cache[3][35] ), .B(n4281), .S0(net112279), .Y(
        \D_cache/n1513 ) );
  MX2XL U10113 ( .A(\D_cache/cache[2][35] ), .B(n4281), .S0(net112403), .Y(
        \D_cache/n1514 ) );
  MX2XL U10114 ( .A(\D_cache/cache[1][35] ), .B(n4281), .S0(net112527), .Y(
        \D_cache/n1515 ) );
  MX2XL U10115 ( .A(\D_cache/cache[0][35] ), .B(n4281), .S0(net112629), .Y(
        \D_cache/n1516 ) );
  MX2XL U10116 ( .A(\D_cache/cache[6][30] ), .B(n4253), .S0(net112009), .Y(
        \D_cache/n1550 ) );
  MX2XL U10117 ( .A(\D_cache/cache[5][30] ), .B(n4253), .S0(net112123), .Y(
        \D_cache/n1551 ) );
  MX2XL U10118 ( .A(\D_cache/cache[4][30] ), .B(n4253), .S0(net112215), .Y(
        \D_cache/n1552 ) );
  MX2XL U10119 ( .A(\D_cache/cache[3][30] ), .B(n4253), .S0(net112277), .Y(
        \D_cache/n1553 ) );
  MX2XL U10120 ( .A(\D_cache/cache[2][30] ), .B(n4253), .S0(net112419), .Y(
        \D_cache/n1554 ) );
  MX2XL U10121 ( .A(\D_cache/cache[1][30] ), .B(n4253), .S0(net112545), .Y(
        \D_cache/n1555 ) );
  MX2XL U10122 ( .A(\D_cache/cache[0][30] ), .B(n4253), .S0(net112647), .Y(
        \D_cache/n1556 ) );
  MX2XL U10123 ( .A(\D_cache/cache[6][29] ), .B(n4254), .S0(net111991), .Y(
        \D_cache/n1558 ) );
  MX2XL U10124 ( .A(\D_cache/cache[5][29] ), .B(n4254), .S0(net112115), .Y(
        \D_cache/n1559 ) );
  MX2XL U10125 ( .A(\D_cache/cache[4][29] ), .B(n4254), .S0(net112197), .Y(
        \D_cache/n1560 ) );
  MX2XL U10126 ( .A(\D_cache/cache[3][29] ), .B(n4254), .S0(net112279), .Y(
        \D_cache/n1561 ) );
  MX2XL U10127 ( .A(\D_cache/cache[2][29] ), .B(n4254), .S0(net112403), .Y(
        \D_cache/n1562 ) );
  MX2XL U10128 ( .A(\D_cache/cache[1][29] ), .B(n4254), .S0(net112527), .Y(
        \D_cache/n1563 ) );
  MX2XL U10129 ( .A(\D_cache/cache[0][29] ), .B(n4254), .S0(net112629), .Y(
        \D_cache/n1564 ) );
  MX2XL U10130 ( .A(\D_cache/cache[6][28] ), .B(n4255), .S0(net111995), .Y(
        \D_cache/n1566 ) );
  MX2XL U10131 ( .A(\D_cache/cache[5][28] ), .B(n4255), .S0(net112119), .Y(
        \D_cache/n1567 ) );
  MX2XL U10132 ( .A(\D_cache/cache[4][28] ), .B(n4255), .S0(net112201), .Y(
        \D_cache/n1568 ) );
  MX2XL U10133 ( .A(\D_cache/cache[3][28] ), .B(n4255), .S0(net112283), .Y(
        \D_cache/n1569 ) );
  MX2XL U10134 ( .A(\D_cache/cache[2][28] ), .B(n4255), .S0(net112401), .Y(
        \D_cache/n1570 ) );
  MX2XL U10135 ( .A(\D_cache/cache[1][28] ), .B(n4255), .S0(net112531), .Y(
        \D_cache/n1571 ) );
  MX2XL U10136 ( .A(\D_cache/cache[0][28] ), .B(n4255), .S0(net112633), .Y(
        \D_cache/n1572 ) );
  MX2XL U10137 ( .A(\D_cache/cache[6][27] ), .B(n4256), .S0(net111989), .Y(
        \D_cache/n1574 ) );
  MX2XL U10138 ( .A(\D_cache/cache[5][27] ), .B(n4256), .S0(net112113), .Y(
        \D_cache/n1575 ) );
  MX2XL U10139 ( .A(\D_cache/cache[4][27] ), .B(n4256), .S0(net112195), .Y(
        \D_cache/n1576 ) );
  MX2XL U10140 ( .A(\D_cache/cache[3][27] ), .B(n4256), .S0(net112277), .Y(
        \D_cache/n1577 ) );
  MX2XL U10141 ( .A(\D_cache/cache[2][27] ), .B(n4256), .S0(net112405), .Y(
        \D_cache/n1578 ) );
  MX2XL U10142 ( .A(\D_cache/cache[1][27] ), .B(n4256), .S0(net112535), .Y(
        \D_cache/n1579 ) );
  MX2XL U10143 ( .A(\D_cache/cache[0][27] ), .B(n4256), .S0(net112629), .Y(
        \D_cache/n1580 ) );
  MX2XL U10144 ( .A(\D_cache/cache[6][26] ), .B(n4257), .S0(net111995), .Y(
        \D_cache/n1582 ) );
  MX2XL U10145 ( .A(\D_cache/cache[5][26] ), .B(n4257), .S0(net112119), .Y(
        \D_cache/n1583 ) );
  MX2XL U10146 ( .A(\D_cache/cache[4][26] ), .B(n4257), .S0(net112201), .Y(
        \D_cache/n1584 ) );
  MX2XL U10147 ( .A(\D_cache/cache[3][26] ), .B(n4257), .S0(net112283), .Y(
        \D_cache/n1585 ) );
  MX2XL U10148 ( .A(\D_cache/cache[1][26] ), .B(n4257), .S0(net112531), .Y(
        \D_cache/n1587 ) );
  MX2XL U10149 ( .A(\D_cache/cache[0][26] ), .B(n4257), .S0(net112633), .Y(
        \D_cache/n1588 ) );
  MX2XL U10150 ( .A(\D_cache/cache[6][25] ), .B(n10425), .S0(net111993), .Y(
        \D_cache/n1590 ) );
  MX2XL U10151 ( .A(\D_cache/cache[5][25] ), .B(n10425), .S0(net112117), .Y(
        \D_cache/n1591 ) );
  MX2XL U10152 ( .A(\D_cache/cache[4][25] ), .B(n10425), .S0(net112199), .Y(
        \D_cache/n1592 ) );
  MX2XL U10153 ( .A(\D_cache/cache[3][25] ), .B(n10425), .S0(net112281), .Y(
        \D_cache/n1593 ) );
  MX2XL U10154 ( .A(\D_cache/cache[2][25] ), .B(n10425), .S0(net112405), .Y(
        \D_cache/n1594 ) );
  MX2XL U10155 ( .A(\D_cache/cache[1][25] ), .B(n10425), .S0(net112525), .Y(
        \D_cache/n1595 ) );
  MX2XL U10156 ( .A(\D_cache/cache[0][25] ), .B(n10425), .S0(net112627), .Y(
        \D_cache/n1596 ) );
  MX2XL U10157 ( .A(\D_cache/cache[6][24] ), .B(n4258), .S0(net112003), .Y(
        \D_cache/n1598 ) );
  MX2XL U10158 ( .A(\D_cache/cache[5][24] ), .B(n4258), .S0(net112127), .Y(
        \D_cache/n1599 ) );
  MX2XL U10159 ( .A(\D_cache/cache[4][24] ), .B(n4258), .S0(net112211), .Y(
        \D_cache/n1600 ) );
  MX2XL U10160 ( .A(\D_cache/cache[3][24] ), .B(n4258), .S0(net112291), .Y(
        \D_cache/n1601 ) );
  MX2XL U10161 ( .A(\D_cache/cache[2][24] ), .B(n4258), .S0(net112415), .Y(
        \D_cache/n1602 ) );
  MX2XL U10162 ( .A(\D_cache/cache[1][24] ), .B(n4258), .S0(net112539), .Y(
        \D_cache/n1603 ) );
  MX2XL U10163 ( .A(\D_cache/cache[0][24] ), .B(n4258), .S0(net112641), .Y(
        \D_cache/n1604 ) );
  MX2XL U10164 ( .A(\D_cache/cache[6][23] ), .B(n4259), .S0(net112009), .Y(
        \D_cache/n1606 ) );
  MX2XL U10165 ( .A(\D_cache/cache[5][23] ), .B(n4259), .S0(net112125), .Y(
        \D_cache/n1607 ) );
  MX2XL U10166 ( .A(\D_cache/cache[4][23] ), .B(n4259), .S0(net112211), .Y(
        \D_cache/n1608 ) );
  MX2XL U10167 ( .A(\D_cache/cache[3][23] ), .B(n4259), .S0(net112289), .Y(
        \D_cache/n1609 ) );
  MX2XL U10168 ( .A(\D_cache/cache[2][23] ), .B(n4259), .S0(net112415), .Y(
        \D_cache/n1610 ) );
  MX2XL U10169 ( .A(\D_cache/cache[1][23] ), .B(n4259), .S0(net112537), .Y(
        \D_cache/n1611 ) );
  MX2XL U10170 ( .A(\D_cache/cache[0][23] ), .B(n4259), .S0(net112639), .Y(
        \D_cache/n1612 ) );
  MX2XL U10171 ( .A(\D_cache/cache[6][22] ), .B(n4260), .S0(net112005), .Y(
        \D_cache/n1614 ) );
  MX2XL U10172 ( .A(\D_cache/cache[5][22] ), .B(n4260), .S0(net112125), .Y(
        \D_cache/n1615 ) );
  MX2XL U10173 ( .A(\D_cache/cache[4][22] ), .B(n4260), .S0(net112211), .Y(
        \D_cache/n1616 ) );
  MX2XL U10174 ( .A(\D_cache/cache[3][22] ), .B(n4260), .S0(net112289), .Y(
        \D_cache/n1617 ) );
  MX2XL U10175 ( .A(\D_cache/cache[2][22] ), .B(n4260), .S0(net112415), .Y(
        \D_cache/n1618 ) );
  MX2XL U10176 ( .A(\D_cache/cache[1][22] ), .B(n4260), .S0(net112537), .Y(
        \D_cache/n1619 ) );
  MX2XL U10177 ( .A(\D_cache/cache[0][22] ), .B(n4260), .S0(net112639), .Y(
        \D_cache/n1620 ) );
  MX2XL U10178 ( .A(\D_cache/cache[6][21] ), .B(n10534), .S0(net111995), .Y(
        \D_cache/n1622 ) );
  MX2XL U10179 ( .A(\D_cache/cache[5][21] ), .B(n10534), .S0(net112125), .Y(
        \D_cache/n1623 ) );
  MX2XL U10180 ( .A(\D_cache/cache[4][21] ), .B(n10534), .S0(net112211), .Y(
        \D_cache/n1624 ) );
  MX2XL U10181 ( .A(\D_cache/cache[3][21] ), .B(n10534), .S0(net112289), .Y(
        \D_cache/n1625 ) );
  MX2XL U10182 ( .A(\D_cache/cache[2][21] ), .B(n10534), .S0(net112405), .Y(
        \D_cache/n1626 ) );
  MX2XL U10183 ( .A(\D_cache/cache[1][21] ), .B(n10534), .S0(net112537), .Y(
        \D_cache/n1627 ) );
  MX2XL U10184 ( .A(\D_cache/cache[0][21] ), .B(n10534), .S0(net112639), .Y(
        \D_cache/n1628 ) );
  MX2XL U10185 ( .A(\D_cache/cache[6][20] ), .B(n10522), .S0(net111991), .Y(
        \D_cache/n1630 ) );
  MX2XL U10186 ( .A(\D_cache/cache[5][20] ), .B(n10522), .S0(net112115), .Y(
        \D_cache/n1631 ) );
  MX2XL U10187 ( .A(\D_cache/cache[4][20] ), .B(n10522), .S0(net112197), .Y(
        \D_cache/n1632 ) );
  MX2XL U10188 ( .A(\D_cache/cache[3][20] ), .B(n10522), .S0(net112279), .Y(
        \D_cache/n1633 ) );
  MX2XL U10189 ( .A(\D_cache/cache[2][20] ), .B(n10522), .S0(net112403), .Y(
        \D_cache/n1634 ) );
  MX2XL U10190 ( .A(\D_cache/cache[1][20] ), .B(n10522), .S0(net112527), .Y(
        \D_cache/n1635 ) );
  MX2XL U10191 ( .A(\D_cache/cache[0][20] ), .B(n10522), .S0(net112629), .Y(
        \D_cache/n1636 ) );
  MX2XL U10192 ( .A(\D_cache/cache[6][19] ), .B(n4261), .S0(net111993), .Y(
        \D_cache/n1638 ) );
  MX2XL U10193 ( .A(\D_cache/cache[5][19] ), .B(n4261), .S0(net112117), .Y(
        \D_cache/n1639 ) );
  MX2XL U10194 ( .A(\D_cache/cache[4][19] ), .B(n4261), .S0(net112199), .Y(
        \D_cache/n1640 ) );
  MX2XL U10195 ( .A(\D_cache/cache[3][19] ), .B(n4261), .S0(net112281), .Y(
        \D_cache/n1641 ) );
  MX2XL U10196 ( .A(\D_cache/cache[2][19] ), .B(n4261), .S0(net112405), .Y(
        \D_cache/n1642 ) );
  MX2XL U10197 ( .A(\D_cache/cache[1][19] ), .B(n4261), .S0(net112529), .Y(
        \D_cache/n1643 ) );
  MX2XL U10198 ( .A(\D_cache/cache[0][19] ), .B(n4261), .S0(net112631), .Y(
        \D_cache/n1644 ) );
  MX2XL U10199 ( .A(\D_cache/cache[6][18] ), .B(n4262), .S0(net111989), .Y(
        \D_cache/n1646 ) );
  MX2XL U10200 ( .A(\D_cache/cache[5][18] ), .B(n4262), .S0(net112123), .Y(
        \D_cache/n1647 ) );
  MX2XL U10201 ( .A(\D_cache/cache[4][18] ), .B(n4262), .S0(net112211), .Y(
        \D_cache/n1648 ) );
  MX2XL U10202 ( .A(\D_cache/cache[3][18] ), .B(n4262), .S0(net112285), .Y(
        \D_cache/n1649 ) );
  MX2XL U10203 ( .A(\D_cache/cache[2][18] ), .B(n4262), .S0(net112409), .Y(
        \D_cache/n1650 ) );
  MX2XL U10204 ( .A(\D_cache/cache[1][18] ), .B(n4262), .S0(net112533), .Y(
        \D_cache/n1651 ) );
  MX2XL U10205 ( .A(\D_cache/cache[0][18] ), .B(n4262), .S0(net112635), .Y(
        \D_cache/n1652 ) );
  MX2XL U10206 ( .A(\D_cache/cache[6][17] ), .B(n10597), .S0(net112003), .Y(
        \D_cache/n1654 ) );
  MX2XL U10207 ( .A(\D_cache/cache[5][17] ), .B(n10597), .S0(net112127), .Y(
        \D_cache/n1655 ) );
  MX2XL U10208 ( .A(\D_cache/cache[4][17] ), .B(n10597), .S0(net112197), .Y(
        \D_cache/n1656 ) );
  MX2XL U10209 ( .A(\D_cache/cache[3][17] ), .B(n10597), .S0(net112291), .Y(
        \D_cache/n1657 ) );
  MX2XL U10210 ( .A(\D_cache/cache[2][17] ), .B(n10597), .S0(net112415), .Y(
        \D_cache/n1658 ) );
  MX2XL U10211 ( .A(\D_cache/cache[1][17] ), .B(n10597), .S0(net112539), .Y(
        \D_cache/n1659 ) );
  MX2XL U10212 ( .A(\D_cache/cache[0][17] ), .B(n10597), .S0(net112641), .Y(
        \D_cache/n1660 ) );
  MX2XL U10213 ( .A(\D_cache/cache[6][16] ), .B(n4263), .S0(net111989), .Y(
        \D_cache/n1662 ) );
  MX2XL U10214 ( .A(\D_cache/cache[5][16] ), .B(n4263), .S0(net112113), .Y(
        \D_cache/n1663 ) );
  MX2XL U10215 ( .A(\D_cache/cache[4][16] ), .B(n4263), .S0(net112195), .Y(
        \D_cache/n1664 ) );
  MX2XL U10216 ( .A(\D_cache/cache[3][16] ), .B(n4263), .S0(net112277), .Y(
        \D_cache/n1665 ) );
  MX2XL U10217 ( .A(\D_cache/cache[2][16] ), .B(n4263), .S0(net112401), .Y(
        \D_cache/n1666 ) );
  MX2XL U10218 ( .A(\D_cache/cache[1][16] ), .B(n4263), .S0(net112525), .Y(
        \D_cache/n1667 ) );
  MX2XL U10219 ( .A(\D_cache/cache[0][16] ), .B(n4263), .S0(net112627), .Y(
        \D_cache/n1668 ) );
  MX2XL U10220 ( .A(\D_cache/cache[6][15] ), .B(n10188), .S0(net111995), .Y(
        \D_cache/n1670 ) );
  MX2XL U10221 ( .A(\D_cache/cache[5][15] ), .B(n10188), .S0(net112119), .Y(
        \D_cache/n1671 ) );
  MX2XL U10222 ( .A(\D_cache/cache[4][15] ), .B(n10188), .S0(net112201), .Y(
        \D_cache/n1672 ) );
  MX2XL U10223 ( .A(\D_cache/cache[3][15] ), .B(n10188), .S0(net112283), .Y(
        \D_cache/n1673 ) );
  MX2XL U10224 ( .A(\D_cache/cache[2][15] ), .B(n10188), .S0(net112405), .Y(
        \D_cache/n1674 ) );
  MX2XL U10225 ( .A(\D_cache/cache[1][15] ), .B(n10188), .S0(net112531), .Y(
        \D_cache/n1675 ) );
  MX2XL U10226 ( .A(\D_cache/cache[0][15] ), .B(n10188), .S0(net112633), .Y(
        \D_cache/n1676 ) );
  MX2XL U10227 ( .A(\D_cache/cache[6][14] ), .B(n10437), .S0(net111989), .Y(
        \D_cache/n1678 ) );
  MX2XL U10228 ( .A(\D_cache/cache[5][14] ), .B(n10437), .S0(net112113), .Y(
        \D_cache/n1679 ) );
  MX2XL U10229 ( .A(\D_cache/cache[4][14] ), .B(n10437), .S0(net112195), .Y(
        \D_cache/n1680 ) );
  MX2XL U10230 ( .A(\D_cache/cache[3][14] ), .B(n10437), .S0(net112277), .Y(
        \D_cache/n1681 ) );
  MX2XL U10231 ( .A(\D_cache/cache[2][14] ), .B(n10437), .S0(net112405), .Y(
        \D_cache/n1682 ) );
  MX2XL U10232 ( .A(\D_cache/cache[1][14] ), .B(n10437), .S0(net112525), .Y(
        \D_cache/n1683 ) );
  MX2XL U10233 ( .A(\D_cache/cache[6][10] ), .B(n4264), .S0(net112003), .Y(
        \D_cache/n1710 ) );
  MX2XL U10234 ( .A(\D_cache/cache[5][10] ), .B(n4264), .S0(net112127), .Y(
        \D_cache/n1711 ) );
  MX2XL U10235 ( .A(\D_cache/cache[4][10] ), .B(n4264), .S0(net112197), .Y(
        \D_cache/n1712 ) );
  MX2XL U10236 ( .A(\D_cache/cache[3][10] ), .B(n4264), .S0(net112291), .Y(
        \D_cache/n1713 ) );
  MX2XL U10237 ( .A(\D_cache/cache[2][10] ), .B(n4264), .S0(net112415), .Y(
        \D_cache/n1714 ) );
  MX2XL U10238 ( .A(\D_cache/cache[1][10] ), .B(n4264), .S0(net112539), .Y(
        \D_cache/n1715 ) );
  MX2XL U10239 ( .A(\D_cache/cache[0][10] ), .B(n4264), .S0(net112641), .Y(
        \D_cache/n1716 ) );
  MX2XL U10240 ( .A(\D_cache/cache[6][9] ), .B(n10767), .S0(net112011), .Y(
        \D_cache/n1718 ) );
  MX2XL U10241 ( .A(\D_cache/cache[5][9] ), .B(n10767), .S0(net112121), .Y(
        \D_cache/n1719 ) );
  MX2XL U10242 ( .A(\D_cache/cache[3][9] ), .B(n10767), .S0(net112293), .Y(
        \D_cache/n1721 ) );
  MX2XL U10243 ( .A(\D_cache/cache[2][9] ), .B(n10767), .S0(net112423), .Y(
        \D_cache/n1722 ) );
  MX2XL U10244 ( .A(\D_cache/cache[1][9] ), .B(n10767), .S0(net112547), .Y(
        \D_cache/n1723 ) );
  MX2XL U10245 ( .A(\D_cache/cache[0][9] ), .B(n10767), .S0(net112649), .Y(
        \D_cache/n1724 ) );
  MX2XL U10246 ( .A(\D_cache/cache[6][7] ), .B(n4265), .S0(net112009), .Y(
        \D_cache/n1734 ) );
  MX2XL U10247 ( .A(\D_cache/cache[5][7] ), .B(n4265), .S0(net112121), .Y(
        \D_cache/n1735 ) );
  MX2XL U10248 ( .A(\D_cache/cache[4][7] ), .B(n4265), .S0(net112215), .Y(
        \D_cache/n1736 ) );
  MX2XL U10249 ( .A(\D_cache/cache[3][7] ), .B(n4265), .S0(net112281), .Y(
        \D_cache/n1737 ) );
  MX2XL U10250 ( .A(\D_cache/cache[2][7] ), .B(n4265), .S0(net112417), .Y(
        \D_cache/n1738 ) );
  MX2XL U10251 ( .A(\D_cache/cache[1][7] ), .B(n4265), .S0(net112545), .Y(
        \D_cache/n1739 ) );
  MX2XL U10252 ( .A(\D_cache/cache[0][7] ), .B(n4265), .S0(net112647), .Y(
        \D_cache/n1740 ) );
  MX2XL U10253 ( .A(\D_cache/cache[6][6] ), .B(n4247), .S0(net111993), .Y(
        \D_cache/n1742 ) );
  MX2XL U10254 ( .A(\D_cache/cache[5][6] ), .B(n4247), .S0(net112117), .Y(
        \D_cache/n1743 ) );
  MX2XL U10255 ( .A(\D_cache/cache[4][6] ), .B(n4247), .S0(net112199), .Y(
        \D_cache/n1744 ) );
  MX2XL U10256 ( .A(\D_cache/cache[3][6] ), .B(n4247), .S0(net112281), .Y(
        \D_cache/n1745 ) );
  MX2XL U10257 ( .A(\D_cache/cache[2][6] ), .B(n4247), .S0(net112401), .Y(
        \D_cache/n1746 ) );
  MX2XL U10258 ( .A(\D_cache/cache[1][6] ), .B(n4247), .S0(net112529), .Y(
        \D_cache/n1747 ) );
  MX2XL U10259 ( .A(\D_cache/cache[0][6] ), .B(n4247), .S0(net112631), .Y(
        \D_cache/n1748 ) );
  MX2XL U10260 ( .A(\D_cache/cache[6][4] ), .B(n4248), .S0(net112005), .Y(
        \D_cache/n1758 ) );
  MX2XL U10261 ( .A(\D_cache/cache[5][4] ), .B(n4248), .S0(net112129), .Y(
        \D_cache/n1759 ) );
  MX2XL U10262 ( .A(\D_cache/cache[4][4] ), .B(n4248), .S0(net112211), .Y(
        \D_cache/n1760 ) );
  MX2XL U10263 ( .A(\D_cache/cache[3][4] ), .B(n4248), .S0(net112293), .Y(
        \D_cache/n1761 ) );
  MX2XL U10264 ( .A(\D_cache/cache[2][4] ), .B(n4248), .S0(net112417), .Y(
        \D_cache/n1762 ) );
  MX2XL U10265 ( .A(\D_cache/cache[1][4] ), .B(n4248), .S0(net112529), .Y(
        \D_cache/n1763 ) );
  MX2XL U10266 ( .A(\D_cache/cache[0][4] ), .B(n4248), .S0(net112631), .Y(
        \D_cache/n1764 ) );
  MX2XL U10267 ( .A(\D_cache/cache[6][3] ), .B(n10509), .S0(net111991), .Y(
        \D_cache/n1766 ) );
  MX2XL U10268 ( .A(\D_cache/cache[5][3] ), .B(n10509), .S0(net112115), .Y(
        \D_cache/n1767 ) );
  MX2XL U10269 ( .A(\D_cache/cache[4][3] ), .B(n10509), .S0(net112197), .Y(
        \D_cache/n1768 ) );
  MX2XL U10270 ( .A(\D_cache/cache[3][3] ), .B(n10509), .S0(net112279), .Y(
        \D_cache/n1769 ) );
  MX2XL U10271 ( .A(\D_cache/cache[2][3] ), .B(n10509), .S0(net112403), .Y(
        \D_cache/n1770 ) );
  MX2XL U10272 ( .A(\D_cache/cache[1][3] ), .B(n10509), .S0(net112541), .Y(
        \D_cache/n1771 ) );
  MX2XL U10273 ( .A(\D_cache/cache[0][3] ), .B(n10509), .S0(net112631), .Y(
        \D_cache/n1772 ) );
  MX2XL U10274 ( .A(\D_cache/cache[6][94] ), .B(n4283), .S0(net112009), .Y(
        \D_cache/n1038 ) );
  MX2XL U10275 ( .A(\D_cache/cache[5][94] ), .B(n4283), .S0(net112123), .Y(
        \D_cache/n1039 ) );
  MX2XL U10276 ( .A(\D_cache/cache[4][94] ), .B(n4283), .S0(net112215), .Y(
        \D_cache/n1040 ) );
  MX2XL U10277 ( .A(\D_cache/cache[3][94] ), .B(n4283), .S0(net112279), .Y(
        \D_cache/n1041 ) );
  MX2XL U10278 ( .A(\D_cache/cache[2][94] ), .B(n4283), .S0(net112419), .Y(
        \D_cache/n1042 ) );
  MX2XL U10279 ( .A(\D_cache/cache[1][94] ), .B(n4283), .S0(net112545), .Y(
        \D_cache/n1043 ) );
  MX2XL U10280 ( .A(\D_cache/cache[0][94] ), .B(n4283), .S0(net112647), .Y(
        \D_cache/n1044 ) );
  MX2XL U10281 ( .A(\D_cache/cache[6][93] ), .B(n4284), .S0(net111991), .Y(
        \D_cache/n1046 ) );
  MX2XL U10282 ( .A(\D_cache/cache[5][93] ), .B(n4284), .S0(net112115), .Y(
        \D_cache/n1047 ) );
  MX2XL U10283 ( .A(\D_cache/cache[4][93] ), .B(n4284), .S0(net112197), .Y(
        \D_cache/n1048 ) );
  MX2XL U10284 ( .A(\D_cache/cache[3][93] ), .B(n4284), .S0(net112279), .Y(
        \D_cache/n1049 ) );
  MX2XL U10285 ( .A(\D_cache/cache[2][93] ), .B(n4284), .S0(net112403), .Y(
        \D_cache/n1050 ) );
  MX2XL U10286 ( .A(\D_cache/cache[1][93] ), .B(n4284), .S0(net112527), .Y(
        \D_cache/n1051 ) );
  MX2XL U10287 ( .A(\D_cache/cache[0][93] ), .B(n4284), .S0(net112629), .Y(
        \D_cache/n1052 ) );
  MX2XL U10288 ( .A(\D_cache/cache[6][92] ), .B(n4285), .S0(net111995), .Y(
        \D_cache/n1054 ) );
  MX2XL U10289 ( .A(\D_cache/cache[5][92] ), .B(n4285), .S0(net112119), .Y(
        \D_cache/n1055 ) );
  MX2XL U10290 ( .A(\D_cache/cache[4][92] ), .B(n4285), .S0(net112201), .Y(
        \D_cache/n1056 ) );
  MX2XL U10291 ( .A(\D_cache/cache[3][92] ), .B(n4285), .S0(net112283), .Y(
        \D_cache/n1057 ) );
  MX2XL U10292 ( .A(\D_cache/cache[2][92] ), .B(n4285), .S0(net112401), .Y(
        \D_cache/n1058 ) );
  MX2XL U10293 ( .A(\D_cache/cache[1][92] ), .B(n4285), .S0(net112531), .Y(
        \D_cache/n1059 ) );
  MX2XL U10294 ( .A(\D_cache/cache[0][92] ), .B(n4285), .S0(net112633), .Y(
        \D_cache/n1060 ) );
  MX2XL U10295 ( .A(\D_cache/cache[6][91] ), .B(n4286), .S0(net111991), .Y(
        \D_cache/n1062 ) );
  MX2XL U10296 ( .A(\D_cache/cache[5][91] ), .B(n4286), .S0(net112115), .Y(
        \D_cache/n1063 ) );
  MX2XL U10297 ( .A(\D_cache/cache[4][91] ), .B(n4286), .S0(net112197), .Y(
        \D_cache/n1064 ) );
  MX2XL U10298 ( .A(\D_cache/cache[3][91] ), .B(n4286), .S0(net112279), .Y(
        \D_cache/n1065 ) );
  MX2XL U10299 ( .A(\D_cache/cache[2][91] ), .B(n4286), .S0(net112403), .Y(
        \D_cache/n1066 ) );
  MX2XL U10300 ( .A(\D_cache/cache[1][91] ), .B(n4286), .S0(net112527), .Y(
        \D_cache/n1067 ) );
  MX2XL U10301 ( .A(\D_cache/cache[0][91] ), .B(n4286), .S0(net112629), .Y(
        \D_cache/n1068 ) );
  MX2XL U10302 ( .A(\D_cache/cache[6][90] ), .B(n4287), .S0(net111993), .Y(
        \D_cache/n1070 ) );
  MX2XL U10303 ( .A(\D_cache/cache[5][90] ), .B(n4287), .S0(net112117), .Y(
        \D_cache/n1071 ) );
  MX2XL U10304 ( .A(\D_cache/cache[4][90] ), .B(n4287), .S0(net112199), .Y(
        \D_cache/n1072 ) );
  MX2XL U10305 ( .A(\D_cache/cache[3][90] ), .B(n4287), .S0(net112281), .Y(
        \D_cache/n1073 ) );
  MX2XL U10306 ( .A(\D_cache/cache[2][90] ), .B(n4287), .S0(net112405), .Y(
        \D_cache/n1074 ) );
  MX2XL U10307 ( .A(\D_cache/cache[1][90] ), .B(n4287), .S0(net112529), .Y(
        \D_cache/n1075 ) );
  MX2XL U10308 ( .A(\D_cache/cache[0][90] ), .B(n4287), .S0(net112627), .Y(
        \D_cache/n1076 ) );
  MX2XL U10309 ( .A(\D_cache/cache[6][89] ), .B(n4288), .S0(net111989), .Y(
        \D_cache/n1078 ) );
  MX2XL U10310 ( .A(\D_cache/cache[5][89] ), .B(n4288), .S0(net112113), .Y(
        \D_cache/n1079 ) );
  MX2XL U10311 ( .A(\D_cache/cache[4][89] ), .B(n4288), .S0(net112195), .Y(
        \D_cache/n1080 ) );
  MX2XL U10312 ( .A(\D_cache/cache[3][89] ), .B(n4288), .S0(net112277), .Y(
        \D_cache/n1081 ) );
  MX2XL U10313 ( .A(\D_cache/cache[2][89] ), .B(n4288), .S0(net112401), .Y(
        \D_cache/n1082 ) );
  MX2XL U10314 ( .A(\D_cache/cache[1][89] ), .B(n4288), .S0(net112525), .Y(
        \D_cache/n1083 ) );
  MX2XL U10315 ( .A(\D_cache/cache[0][89] ), .B(n4288), .S0(net112627), .Y(
        \D_cache/n1084 ) );
  MX2XL U10316 ( .A(\D_cache/cache[6][88] ), .B(n4289), .S0(net112003), .Y(
        \D_cache/n1086 ) );
  MX2XL U10317 ( .A(\D_cache/cache[5][88] ), .B(n4289), .S0(net112127), .Y(
        \D_cache/n1087 ) );
  MX2XL U10318 ( .A(\D_cache/cache[4][88] ), .B(n4289), .S0(net112195), .Y(
        \D_cache/n1088 ) );
  MX2XL U10319 ( .A(\D_cache/cache[3][88] ), .B(n4289), .S0(net112291), .Y(
        \D_cache/n1089 ) );
  MX2XL U10320 ( .A(\D_cache/cache[2][88] ), .B(n4289), .S0(net112415), .Y(
        \D_cache/n1090 ) );
  MX2XL U10321 ( .A(\D_cache/cache[1][88] ), .B(n4289), .S0(net112539), .Y(
        \D_cache/n1091 ) );
  MX2XL U10322 ( .A(\D_cache/cache[0][88] ), .B(n4289), .S0(net112641), .Y(
        \D_cache/n1092 ) );
  MX2XL U10323 ( .A(\D_cache/cache[6][87] ), .B(n4290), .S0(net112003), .Y(
        \D_cache/n1094 ) );
  MX2XL U10324 ( .A(\D_cache/cache[5][87] ), .B(n4290), .S0(net112127), .Y(
        \D_cache/n1095 ) );
  MX2XL U10325 ( .A(\D_cache/cache[4][87] ), .B(n4290), .S0(net112199), .Y(
        \D_cache/n1096 ) );
  MX2XL U10326 ( .A(\D_cache/cache[3][87] ), .B(n4290), .S0(net112291), .Y(
        \D_cache/n1097 ) );
  MX2XL U10327 ( .A(\D_cache/cache[2][87] ), .B(n4290), .S0(net112415), .Y(
        \D_cache/n1098 ) );
  MX2XL U10328 ( .A(\D_cache/cache[1][87] ), .B(n4290), .S0(net112539), .Y(
        \D_cache/n1099 ) );
  MX2XL U10329 ( .A(\D_cache/cache[0][87] ), .B(n4290), .S0(net112641), .Y(
        \D_cache/n1100 ) );
  MX2XL U10330 ( .A(\D_cache/cache[6][86] ), .B(n4291), .S0(net111991), .Y(
        \D_cache/n1102 ) );
  MX2XL U10331 ( .A(\D_cache/cache[5][86] ), .B(n4291), .S0(net112125), .Y(
        \D_cache/n1103 ) );
  MX2XL U10332 ( .A(\D_cache/cache[4][86] ), .B(n4291), .S0(net112211), .Y(
        \D_cache/n1104 ) );
  MX2XL U10333 ( .A(\D_cache/cache[3][86] ), .B(n4291), .S0(net112289), .Y(
        \D_cache/n1105 ) );
  MX2XL U10334 ( .A(\D_cache/cache[2][86] ), .B(n4291), .S0(net112415), .Y(
        \D_cache/n1106 ) );
  MX2XL U10335 ( .A(\D_cache/cache[1][86] ), .B(n4291), .S0(net112537), .Y(
        \D_cache/n1107 ) );
  MX2XL U10336 ( .A(\D_cache/cache[0][86] ), .B(n4291), .S0(net112639), .Y(
        \D_cache/n1108 ) );
  MX2XL U10337 ( .A(\D_cache/cache[6][85] ), .B(n4292), .S0(net112005), .Y(
        \D_cache/n1110 ) );
  MX2XL U10338 ( .A(\D_cache/cache[5][85] ), .B(n4292), .S0(net112125), .Y(
        \D_cache/n1111 ) );
  MX2XL U10339 ( .A(\D_cache/cache[4][85] ), .B(n4292), .S0(net112211), .Y(
        \D_cache/n1112 ) );
  MX2XL U10340 ( .A(\D_cache/cache[3][85] ), .B(n4292), .S0(net112289), .Y(
        \D_cache/n1113 ) );
  MX2XL U10341 ( .A(\D_cache/cache[2][85] ), .B(n4292), .S0(net112423), .Y(
        \D_cache/n1114 ) );
  MX2XL U10342 ( .A(\D_cache/cache[1][85] ), .B(n4292), .S0(net112537), .Y(
        \D_cache/n1115 ) );
  MX2XL U10343 ( .A(\D_cache/cache[0][85] ), .B(n4292), .S0(net112639), .Y(
        \D_cache/n1116 ) );
  MX2XL U10344 ( .A(\D_cache/cache[6][84] ), .B(n4293), .S0(net111993), .Y(
        \D_cache/n1118 ) );
  MX2XL U10345 ( .A(\D_cache/cache[5][84] ), .B(n4293), .S0(net112125), .Y(
        \D_cache/n1119 ) );
  MX2XL U10346 ( .A(\D_cache/cache[4][84] ), .B(n4293), .S0(net112211), .Y(
        \D_cache/n1120 ) );
  MX2XL U10347 ( .A(\D_cache/cache[3][84] ), .B(n4293), .S0(net112289), .Y(
        \D_cache/n1121 ) );
  MX2XL U10348 ( .A(\D_cache/cache[2][84] ), .B(n4293), .S0(net112411), .Y(
        \D_cache/n1122 ) );
  MX2XL U10349 ( .A(\D_cache/cache[1][84] ), .B(n4293), .S0(net112537), .Y(
        \D_cache/n1123 ) );
  MX2XL U10350 ( .A(\D_cache/cache[0][84] ), .B(n4293), .S0(net112639), .Y(
        \D_cache/n1124 ) );
  MX2XL U10351 ( .A(\D_cache/cache[6][83] ), .B(n4294), .S0(net111993), .Y(
        \D_cache/n1126 ) );
  MX2XL U10352 ( .A(\D_cache/cache[5][83] ), .B(n4294), .S0(net112117), .Y(
        \D_cache/n1127 ) );
  MX2XL U10353 ( .A(\D_cache/cache[4][83] ), .B(n4294), .S0(net112199), .Y(
        \D_cache/n1128 ) );
  MX2XL U10354 ( .A(\D_cache/cache[3][83] ), .B(n4294), .S0(net112281), .Y(
        \D_cache/n1129 ) );
  MX2XL U10355 ( .A(\D_cache/cache[2][83] ), .B(n4294), .S0(net112401), .Y(
        \D_cache/n1130 ) );
  MX2XL U10356 ( .A(\D_cache/cache[1][83] ), .B(n4294), .S0(net112531), .Y(
        \D_cache/n1131 ) );
  MX2XL U10357 ( .A(\D_cache/cache[0][83] ), .B(n4294), .S0(net112633), .Y(
        \D_cache/n1132 ) );
  MX2XL U10358 ( .A(\D_cache/cache[6][82] ), .B(n4295), .S0(net111999), .Y(
        \D_cache/n1134 ) );
  MX2XL U10359 ( .A(\D_cache/cache[5][82] ), .B(n4295), .S0(net112123), .Y(
        \D_cache/n1135 ) );
  MX2XL U10360 ( .A(\D_cache/cache[4][82] ), .B(n4295), .S0(net112195), .Y(
        \D_cache/n1136 ) );
  MX2XL U10361 ( .A(\D_cache/cache[3][82] ), .B(n4295), .S0(net112285), .Y(
        \D_cache/n1137 ) );
  MX2XL U10362 ( .A(\D_cache/cache[2][82] ), .B(n4295), .S0(net112409), .Y(
        \D_cache/n1138 ) );
  MX2XL U10363 ( .A(\D_cache/cache[1][82] ), .B(n4295), .S0(net112533), .Y(
        \D_cache/n1139 ) );
  MX2XL U10364 ( .A(\D_cache/cache[0][82] ), .B(n4295), .S0(net112635), .Y(
        \D_cache/n1140 ) );
  MX2XL U10365 ( .A(\D_cache/cache[6][81] ), .B(n10606), .S0(net112011), .Y(
        \D_cache/n1142 ) );
  MX2XL U10366 ( .A(\D_cache/cache[5][81] ), .B(n10606), .S0(net112125), .Y(
        \D_cache/n1143 ) );
  MX2XL U10367 ( .A(\D_cache/cache[4][81] ), .B(n10606), .S0(net112213), .Y(
        \D_cache/n1144 ) );
  MX2XL U10368 ( .A(\D_cache/cache[3][81] ), .B(n10606), .S0(net112289), .Y(
        \D_cache/n1145 ) );
  MX2XL U10369 ( .A(\D_cache/cache[2][81] ), .B(n10606), .S0(net112403), .Y(
        \D_cache/n1146 ) );
  MX2XL U10370 ( .A(\D_cache/cache[1][81] ), .B(n10606), .S0(net112537), .Y(
        \D_cache/n1147 ) );
  MX2XL U10371 ( .A(\D_cache/cache[0][81] ), .B(n10606), .S0(net112639), .Y(
        \D_cache/n1148 ) );
  MX2XL U10372 ( .A(\D_cache/cache[6][80] ), .B(n4296), .S0(net111989), .Y(
        \D_cache/n1150 ) );
  MX2XL U10373 ( .A(\D_cache/cache[5][80] ), .B(n4296), .S0(net112113), .Y(
        \D_cache/n1151 ) );
  MX2XL U10374 ( .A(\D_cache/cache[4][80] ), .B(n4296), .S0(net112195), .Y(
        \D_cache/n1152 ) );
  MX2XL U10375 ( .A(\D_cache/cache[3][80] ), .B(n4296), .S0(net112277), .Y(
        \D_cache/n1153 ) );
  MX2XL U10376 ( .A(\D_cache/cache[2][80] ), .B(n4296), .S0(net112405), .Y(
        \D_cache/n1154 ) );
  MX2XL U10377 ( .A(\D_cache/cache[1][80] ), .B(n4296), .S0(net112525), .Y(
        \D_cache/n1155 ) );
  MX2XL U10378 ( .A(\D_cache/cache[0][80] ), .B(n4296), .S0(net112637), .Y(
        \D_cache/n1156 ) );
  MX2XL U10379 ( .A(\D_cache/cache[6][79] ), .B(n4297), .S0(net111995), .Y(
        \D_cache/n1158 ) );
  MX2XL U10380 ( .A(\D_cache/cache[5][79] ), .B(n4297), .S0(net112119), .Y(
        \D_cache/n1159 ) );
  MX2XL U10381 ( .A(\D_cache/cache[4][79] ), .B(n4297), .S0(net112201), .Y(
        \D_cache/n1160 ) );
  MX2XL U10382 ( .A(\D_cache/cache[3][79] ), .B(n4297), .S0(net112283), .Y(
        \D_cache/n1161 ) );
  MX2XL U10383 ( .A(\D_cache/cache[2][79] ), .B(n4297), .S0(net112405), .Y(
        \D_cache/n1162 ) );
  MX2XL U10384 ( .A(\D_cache/cache[1][79] ), .B(n4297), .S0(net112531), .Y(
        \D_cache/n1163 ) );
  MX2XL U10385 ( .A(\D_cache/cache[0][79] ), .B(n4297), .S0(net112633), .Y(
        \D_cache/n1164 ) );
  MX2XL U10386 ( .A(\D_cache/cache[6][78] ), .B(n4298), .S0(net111989), .Y(
        \D_cache/n1166 ) );
  MX2XL U10387 ( .A(\D_cache/cache[5][78] ), .B(n4298), .S0(net112113), .Y(
        \D_cache/n1167 ) );
  MX2XL U10388 ( .A(\D_cache/cache[4][78] ), .B(n4298), .S0(net112195), .Y(
        \D_cache/n1168 ) );
  MX2XL U10389 ( .A(\D_cache/cache[3][78] ), .B(n4298), .S0(net112277), .Y(
        \D_cache/n1169 ) );
  MX2XL U10390 ( .A(\D_cache/cache[2][78] ), .B(n4298), .S0(net112401), .Y(
        \D_cache/n1170 ) );
  MX2XL U10391 ( .A(\D_cache/cache[1][78] ), .B(n4298), .S0(net112525), .Y(
        \D_cache/n1171 ) );
  MX2XL U10392 ( .A(\D_cache/cache[0][78] ), .B(n4298), .S0(net112627), .Y(
        \D_cache/n1172 ) );
  MX2XL U10393 ( .A(\D_cache/cache[6][74] ), .B(n10594), .S0(net112003), .Y(
        \D_cache/n1198 ) );
  MX2XL U10394 ( .A(\D_cache/cache[5][74] ), .B(n10594), .S0(net112127), .Y(
        \D_cache/n1199 ) );
  MX2XL U10395 ( .A(\D_cache/cache[4][74] ), .B(n10594), .S0(net112201), .Y(
        \D_cache/n1200 ) );
  MX2XL U10396 ( .A(\D_cache/cache[3][74] ), .B(n10594), .S0(net112291), .Y(
        \D_cache/n1201 ) );
  MX2XL U10397 ( .A(\D_cache/cache[2][74] ), .B(n10594), .S0(net112415), .Y(
        \D_cache/n1202 ) );
  MX2XL U10398 ( .A(\D_cache/cache[1][74] ), .B(n10594), .S0(net112539), .Y(
        \D_cache/n1203 ) );
  MX2XL U10399 ( .A(\D_cache/cache[0][74] ), .B(n10594), .S0(net112641), .Y(
        \D_cache/n1204 ) );
  MX2XL U10400 ( .A(\D_cache/cache[6][73] ), .B(n4299), .S0(net112011), .Y(
        \D_cache/n1206 ) );
  MX2XL U10401 ( .A(\D_cache/cache[5][73] ), .B(n4299), .S0(net112121), .Y(
        \D_cache/n1207 ) );
  MX2XL U10402 ( .A(\D_cache/cache[3][73] ), .B(n4299), .S0(net112295), .Y(
        \D_cache/n1209 ) );
  MX2XL U10403 ( .A(\D_cache/cache[2][73] ), .B(n4299), .S0(net112423), .Y(
        \D_cache/n1210 ) );
  MX2XL U10404 ( .A(\D_cache/cache[1][73] ), .B(n4299), .S0(net112547), .Y(
        \D_cache/n1211 ) );
  MX2XL U10405 ( .A(\D_cache/cache[0][73] ), .B(n4299), .S0(net112649), .Y(
        \D_cache/n1212 ) );
  MX2XL U10406 ( .A(\D_cache/cache[6][71] ), .B(n4300), .S0(net112009), .Y(
        \D_cache/n1222 ) );
  MX2XL U10407 ( .A(\D_cache/cache[5][71] ), .B(n4300), .S0(net112121), .Y(
        \D_cache/n1223 ) );
  MX2XL U10408 ( .A(\D_cache/cache[4][71] ), .B(n4300), .S0(net112215), .Y(
        \D_cache/n1224 ) );
  MX2XL U10409 ( .A(\D_cache/cache[3][71] ), .B(n4300), .S0(net112295), .Y(
        \D_cache/n1225 ) );
  MX2XL U10410 ( .A(\D_cache/cache[2][71] ), .B(n4300), .S0(net112417), .Y(
        \D_cache/n1226 ) );
  MX2XL U10411 ( .A(\D_cache/cache[1][71] ), .B(n4300), .S0(net112545), .Y(
        \D_cache/n1227 ) );
  MX2XL U10412 ( .A(\D_cache/cache[0][71] ), .B(n4300), .S0(net112647), .Y(
        \D_cache/n1228 ) );
  MX2XL U10413 ( .A(\D_cache/cache[6][70] ), .B(n4282), .S0(net111993), .Y(
        \D_cache/n1230 ) );
  MX2XL U10414 ( .A(\D_cache/cache[5][70] ), .B(n4282), .S0(net112117), .Y(
        \D_cache/n1231 ) );
  MX2XL U10415 ( .A(\D_cache/cache[4][70] ), .B(n4282), .S0(net112199), .Y(
        \D_cache/n1232 ) );
  MX2XL U10416 ( .A(\D_cache/cache[3][70] ), .B(n4282), .S0(net112281), .Y(
        \D_cache/n1233 ) );
  MX2XL U10417 ( .A(\D_cache/cache[2][70] ), .B(n4282), .S0(net112401), .Y(
        \D_cache/n1234 ) );
  MX2XL U10418 ( .A(\D_cache/cache[1][70] ), .B(n4282), .S0(net112529), .Y(
        \D_cache/n1235 ) );
  MX2XL U10419 ( .A(\D_cache/cache[0][70] ), .B(n4282), .S0(net112631), .Y(
        \D_cache/n1236 ) );
  MX2XL U10420 ( .A(\D_cache/cache[6][69] ), .B(n4301), .S0(net112011), .Y(
        \D_cache/n1238 ) );
  MX2XL U10421 ( .A(\D_cache/cache[5][69] ), .B(n4301), .S0(net112123), .Y(
        \D_cache/n1239 ) );
  MX2XL U10422 ( .A(\D_cache/cache[3][69] ), .B(n4301), .S0(net112289), .Y(
        \D_cache/n1241 ) );
  MX2XL U10423 ( .A(\D_cache/cache[2][69] ), .B(n4301), .S0(net112423), .Y(
        \D_cache/n1242 ) );
  MX2XL U10424 ( .A(\D_cache/cache[1][69] ), .B(n4301), .S0(net112547), .Y(
        \D_cache/n1243 ) );
  MX2XL U10425 ( .A(\D_cache/cache[0][69] ), .B(n4301), .S0(net112649), .Y(
        \D_cache/n1244 ) );
  MX2XL U10426 ( .A(\D_cache/cache[6][68] ), .B(n4251), .S0(net111993), .Y(
        \D_cache/n1246 ) );
  MX2XL U10427 ( .A(\D_cache/cache[5][68] ), .B(n4251), .S0(net112117), .Y(
        \D_cache/n1247 ) );
  MX2XL U10428 ( .A(\D_cache/cache[4][68] ), .B(n4251), .S0(net112199), .Y(
        \D_cache/n1248 ) );
  MX2XL U10429 ( .A(\D_cache/cache[3][68] ), .B(n4251), .S0(net112281), .Y(
        \D_cache/n1249 ) );
  MX2XL U10430 ( .A(\D_cache/cache[2][68] ), .B(n4251), .S0(net112405), .Y(
        \D_cache/n1250 ) );
  MX2XL U10431 ( .A(\D_cache/cache[1][68] ), .B(n4251), .S0(net112529), .Y(
        \D_cache/n1251 ) );
  MX2XL U10432 ( .A(\D_cache/cache[0][68] ), .B(n4251), .S0(net112631), .Y(
        \D_cache/n1252 ) );
  MX2XL U10433 ( .A(\D_cache/cache[6][67] ), .B(n4302), .S0(net111991), .Y(
        \D_cache/n1254 ) );
  MX2XL U10434 ( .A(\D_cache/cache[5][67] ), .B(n4302), .S0(net112115), .Y(
        \D_cache/n1255 ) );
  MX2XL U10435 ( .A(\D_cache/cache[4][67] ), .B(n4302), .S0(net112197), .Y(
        \D_cache/n1256 ) );
  MX2XL U10436 ( .A(\D_cache/cache[3][67] ), .B(n4302), .S0(net112279), .Y(
        \D_cache/n1257 ) );
  MX2XL U10437 ( .A(\D_cache/cache[2][67] ), .B(n4302), .S0(net112403), .Y(
        \D_cache/n1258 ) );
  MX2XL U10438 ( .A(\D_cache/cache[1][67] ), .B(n4302), .S0(net112527), .Y(
        \D_cache/n1259 ) );
  MX2XL U10439 ( .A(\D_cache/cache[0][67] ), .B(n4302), .S0(net112629), .Y(
        \D_cache/n1260 ) );
  MX2XL U10440 ( .A(\D_cache/cache[6][126] ), .B(n4303), .S0(net112009), .Y(
        \D_cache/n782 ) );
  MX2XL U10441 ( .A(\D_cache/cache[5][126] ), .B(n4303), .S0(net112123), .Y(
        \D_cache/n783 ) );
  MX2XL U10442 ( .A(\D_cache/cache[4][126] ), .B(n4303), .S0(net112215), .Y(
        \D_cache/n784 ) );
  MX2XL U10443 ( .A(\D_cache/cache[3][126] ), .B(n4303), .S0(net112293), .Y(
        \D_cache/n785 ) );
  MX2XL U10444 ( .A(\D_cache/cache[2][126] ), .B(n4303), .S0(net112419), .Y(
        \D_cache/n786 ) );
  MX2XL U10445 ( .A(\D_cache/cache[1][126] ), .B(n4303), .S0(net112545), .Y(
        \D_cache/n787 ) );
  MX2XL U10446 ( .A(\D_cache/cache[0][126] ), .B(n4303), .S0(net112647), .Y(
        \D_cache/n788 ) );
  MX2XL U10447 ( .A(\D_cache/cache[6][125] ), .B(n4304), .S0(net111991), .Y(
        \D_cache/n790 ) );
  MX2XL U10448 ( .A(\D_cache/cache[5][125] ), .B(n4304), .S0(net112115), .Y(
        \D_cache/n791 ) );
  MX2XL U10449 ( .A(\D_cache/cache[4][125] ), .B(n4304), .S0(net112197), .Y(
        \D_cache/n792 ) );
  MX2XL U10450 ( .A(\D_cache/cache[3][125] ), .B(n4304), .S0(net112279), .Y(
        \D_cache/n793 ) );
  MX2XL U10451 ( .A(\D_cache/cache[2][125] ), .B(n4304), .S0(net112403), .Y(
        \D_cache/n794 ) );
  MX2XL U10452 ( .A(\D_cache/cache[1][125] ), .B(n4304), .S0(net112527), .Y(
        \D_cache/n795 ) );
  MX2XL U10453 ( .A(\D_cache/cache[0][125] ), .B(n4304), .S0(net112629), .Y(
        \D_cache/n796 ) );
  MX2XL U10454 ( .A(\D_cache/cache[6][124] ), .B(n10403), .S0(net111995), .Y(
        \D_cache/n798 ) );
  MX2XL U10455 ( .A(\D_cache/cache[5][124] ), .B(n10403), .S0(net112119), .Y(
        \D_cache/n799 ) );
  MX2XL U10456 ( .A(\D_cache/cache[4][124] ), .B(n10403), .S0(net112201), .Y(
        \D_cache/n800 ) );
  MX2XL U10457 ( .A(\D_cache/cache[3][124] ), .B(n10403), .S0(net112283), .Y(
        \D_cache/n801 ) );
  MX2XL U10458 ( .A(\D_cache/cache[2][124] ), .B(n10403), .S0(net112401), .Y(
        \D_cache/n802 ) );
  MX2XL U10459 ( .A(\D_cache/cache[1][124] ), .B(n10403), .S0(net112531), .Y(
        \D_cache/n803 ) );
  MX2XL U10460 ( .A(\D_cache/cache[0][124] ), .B(n10403), .S0(net112633), .Y(
        \D_cache/n804 ) );
  MX2XL U10461 ( .A(\D_cache/cache[6][123] ), .B(n4305), .S0(net111991), .Y(
        \D_cache/n806 ) );
  MX2XL U10462 ( .A(\D_cache/cache[5][123] ), .B(n4305), .S0(net112115), .Y(
        \D_cache/n807 ) );
  MX2XL U10463 ( .A(\D_cache/cache[4][123] ), .B(n4305), .S0(net112197), .Y(
        \D_cache/n808 ) );
  MX2XL U10464 ( .A(\D_cache/cache[3][123] ), .B(n4305), .S0(net112279), .Y(
        \D_cache/n809 ) );
  MX2XL U10465 ( .A(\D_cache/cache[2][123] ), .B(n4305), .S0(net112403), .Y(
        \D_cache/n810 ) );
  MX2XL U10466 ( .A(\D_cache/cache[1][123] ), .B(n4305), .S0(net112527), .Y(
        \D_cache/n811 ) );
  MX2XL U10467 ( .A(\D_cache/cache[0][123] ), .B(n4305), .S0(net112629), .Y(
        \D_cache/n812 ) );
  MX2XL U10468 ( .A(\D_cache/cache[6][122] ), .B(n4306), .S0(net111995), .Y(
        \D_cache/n814 ) );
  MX2XL U10469 ( .A(\D_cache/cache[5][122] ), .B(n4306), .S0(net112119), .Y(
        \D_cache/n815 ) );
  MX2XL U10470 ( .A(\D_cache/cache[4][122] ), .B(n4306), .S0(net112201), .Y(
        \D_cache/n816 ) );
  MX2XL U10471 ( .A(\D_cache/cache[3][122] ), .B(n4306), .S0(net112283), .Y(
        \D_cache/n817 ) );
  MX2XL U10472 ( .A(\D_cache/cache[2][122] ), .B(n4306), .S0(net112405), .Y(
        \D_cache/n818 ) );
  MX2XL U10473 ( .A(\D_cache/cache[1][122] ), .B(n4306), .S0(net112529), .Y(
        \D_cache/n819 ) );
  MX2XL U10474 ( .A(\D_cache/cache[0][122] ), .B(n4306), .S0(net112631), .Y(
        \D_cache/n820 ) );
  MX2XL U10475 ( .A(\D_cache/cache[6][121] ), .B(n4307), .S0(net111989), .Y(
        \D_cache/n822 ) );
  MX2XL U10476 ( .A(\D_cache/cache[5][121] ), .B(n4307), .S0(net112113), .Y(
        \D_cache/n823 ) );
  MX2XL U10477 ( .A(\D_cache/cache[4][121] ), .B(n4307), .S0(net112195), .Y(
        \D_cache/n824 ) );
  MX2XL U10478 ( .A(\D_cache/cache[3][121] ), .B(n4307), .S0(net112277), .Y(
        \D_cache/n825 ) );
  MX2XL U10479 ( .A(\D_cache/cache[2][121] ), .B(n4307), .S0(net112405), .Y(
        \D_cache/n826 ) );
  MX2XL U10480 ( .A(\D_cache/cache[1][121] ), .B(n4307), .S0(net112525), .Y(
        \D_cache/n827 ) );
  MX2XL U10481 ( .A(\D_cache/cache[0][121] ), .B(n4307), .S0(net112627), .Y(
        \D_cache/n828 ) );
  MX2XL U10482 ( .A(\D_cache/cache[6][120] ), .B(n4308), .S0(net112003), .Y(
        \D_cache/n830 ) );
  MX2XL U10483 ( .A(\D_cache/cache[5][120] ), .B(n4308), .S0(net112127), .Y(
        \D_cache/n831 ) );
  MX2XL U10484 ( .A(\D_cache/cache[4][120] ), .B(n4308), .S0(net112211), .Y(
        \D_cache/n832 ) );
  MX2XL U10485 ( .A(\D_cache/cache[3][120] ), .B(n4308), .S0(net112291), .Y(
        \D_cache/n833 ) );
  MX2XL U10486 ( .A(\D_cache/cache[2][120] ), .B(n4308), .S0(net112415), .Y(
        \D_cache/n834 ) );
  MX2XL U10487 ( .A(\D_cache/cache[1][120] ), .B(n4308), .S0(net112539), .Y(
        \D_cache/n835 ) );
  MX2XL U10488 ( .A(\D_cache/cache[0][120] ), .B(n4308), .S0(net112641), .Y(
        \D_cache/n836 ) );
  MX2XL U10489 ( .A(\D_cache/cache[6][119] ), .B(n4309), .S0(net111999), .Y(
        \D_cache/n838 ) );
  MX2XL U10490 ( .A(\D_cache/cache[5][119] ), .B(n4309), .S0(net112123), .Y(
        \D_cache/n839 ) );
  MX2XL U10491 ( .A(\D_cache/cache[4][119] ), .B(n4309), .S0(net112215), .Y(
        \D_cache/n840 ) );
  MX2XL U10492 ( .A(\D_cache/cache[3][119] ), .B(n4309), .S0(net112279), .Y(
        \D_cache/n841 ) );
  MX2XL U10493 ( .A(\D_cache/cache[2][119] ), .B(n4309), .S0(net112411), .Y(
        \D_cache/n842 ) );
  MX2XL U10494 ( .A(\D_cache/cache[1][119] ), .B(n4309), .S0(net112535), .Y(
        \D_cache/n843 ) );
  MX2XL U10495 ( .A(\D_cache/cache[0][119] ), .B(n4309), .S0(net112637), .Y(
        \D_cache/n844 ) );
  MX2XL U10496 ( .A(\D_cache/cache[6][118] ), .B(n4310), .S0(net112005), .Y(
        \D_cache/n846 ) );
  MX2XL U10497 ( .A(\D_cache/cache[5][118] ), .B(n4310), .S0(net112125), .Y(
        \D_cache/n847 ) );
  MX2XL U10498 ( .A(\D_cache/cache[4][118] ), .B(n4310), .S0(net112213), .Y(
        \D_cache/n848 ) );
  MX2XL U10499 ( .A(\D_cache/cache[3][118] ), .B(n4310), .S0(net112289), .Y(
        \D_cache/n849 ) );
  MX2XL U10500 ( .A(\D_cache/cache[2][118] ), .B(n4310), .S0(net112411), .Y(
        \D_cache/n850 ) );
  MX2XL U10501 ( .A(\D_cache/cache[1][118] ), .B(n4310), .S0(net112537), .Y(
        \D_cache/n851 ) );
  MX2XL U10502 ( .A(\D_cache/cache[0][118] ), .B(n4310), .S0(net112639), .Y(
        \D_cache/n852 ) );
  MX2XL U10503 ( .A(\D_cache/cache[6][117] ), .B(n4311), .S0(net112003), .Y(
        \D_cache/n854 ) );
  MX2XL U10504 ( .A(\D_cache/cache[5][117] ), .B(n4311), .S0(net112125), .Y(
        \D_cache/n855 ) );
  MX2XL U10505 ( .A(\D_cache/cache[4][117] ), .B(n4311), .S0(net112213), .Y(
        \D_cache/n856 ) );
  MX2XL U10506 ( .A(\D_cache/cache[3][117] ), .B(n4311), .S0(net112289), .Y(
        \D_cache/n857 ) );
  MX2XL U10507 ( .A(\D_cache/cache[2][117] ), .B(n4311), .S0(net112403), .Y(
        \D_cache/n858 ) );
  MX2XL U10508 ( .A(\D_cache/cache[1][117] ), .B(n4311), .S0(net112537), .Y(
        \D_cache/n859 ) );
  MX2XL U10509 ( .A(\D_cache/cache[0][117] ), .B(n4311), .S0(net112639), .Y(
        \D_cache/n860 ) );
  MX2XL U10510 ( .A(\D_cache/cache[6][116] ), .B(n4312), .S0(net112003), .Y(
        \D_cache/n862 ) );
  MX2XL U10511 ( .A(\D_cache/cache[5][116] ), .B(n4312), .S0(net112125), .Y(
        \D_cache/n863 ) );
  MX2XL U10512 ( .A(\D_cache/cache[4][116] ), .B(n4312), .S0(net112213), .Y(
        \D_cache/n864 ) );
  MX2XL U10513 ( .A(\D_cache/cache[3][116] ), .B(n4312), .S0(net112289), .Y(
        \D_cache/n865 ) );
  MX2XL U10514 ( .A(\D_cache/cache[2][116] ), .B(n4312), .S0(net112411), .Y(
        \D_cache/n866 ) );
  MX2XL U10515 ( .A(\D_cache/cache[1][116] ), .B(n4312), .S0(net112537), .Y(
        \D_cache/n867 ) );
  MX2XL U10516 ( .A(\D_cache/cache[0][116] ), .B(n4312), .S0(net112639), .Y(
        \D_cache/n868 ) );
  MX2XL U10517 ( .A(\D_cache/cache[6][115] ), .B(n10180), .S0(net111993), .Y(
        \D_cache/n870 ) );
  MX2XL U10518 ( .A(\D_cache/cache[5][115] ), .B(n10180), .S0(net112117), .Y(
        \D_cache/n871 ) );
  MX2XL U10519 ( .A(\D_cache/cache[4][115] ), .B(n10180), .S0(net112199), .Y(
        \D_cache/n872 ) );
  MX2XL U10520 ( .A(\D_cache/cache[3][115] ), .B(n10180), .S0(net112281), .Y(
        \D_cache/n873 ) );
  MX2XL U10521 ( .A(\D_cache/cache[2][115] ), .B(n10180), .S0(net112401), .Y(
        \D_cache/n874 ) );
  MX2XL U10522 ( .A(\D_cache/cache[1][115] ), .B(n10180), .S0(net112529), .Y(
        \D_cache/n875 ) );
  MX2XL U10523 ( .A(\D_cache/cache[0][115] ), .B(n10180), .S0(net112633), .Y(
        \D_cache/n876 ) );
  MX2XL U10524 ( .A(\D_cache/cache[6][114] ), .B(n4313), .S0(net112009), .Y(
        \D_cache/n878 ) );
  MX2XL U10525 ( .A(\D_cache/cache[5][114] ), .B(n4313), .S0(net112121), .Y(
        \D_cache/n879 ) );
  MX2XL U10526 ( .A(\D_cache/cache[4][114] ), .B(n4313), .S0(net112199), .Y(
        \D_cache/n880 ) );
  MX2XL U10527 ( .A(\D_cache/cache[3][114] ), .B(n4313), .S0(net112285), .Y(
        \D_cache/n881 ) );
  MX2XL U10528 ( .A(\D_cache/cache[2][114] ), .B(n4313), .S0(net112409), .Y(
        \D_cache/n882 ) );
  MX2XL U10529 ( .A(\D_cache/cache[1][114] ), .B(n4313), .S0(net112533), .Y(
        \D_cache/n883 ) );
  MX2XL U10530 ( .A(\D_cache/cache[0][114] ), .B(n4313), .S0(net112635), .Y(
        \D_cache/n884 ) );
  MX2XL U10531 ( .A(\D_cache/cache[6][113] ), .B(n4314), .S0(net112003), .Y(
        \D_cache/n886 ) );
  MX2XL U10532 ( .A(\D_cache/cache[5][113] ), .B(n4314), .S0(net112127), .Y(
        \D_cache/n887 ) );
  MX2XL U10533 ( .A(\D_cache/cache[4][113] ), .B(n4314), .S0(net112215), .Y(
        \D_cache/n888 ) );
  MX2XL U10534 ( .A(\D_cache/cache[3][113] ), .B(n4314), .S0(net112291), .Y(
        \D_cache/n889 ) );
  MX2XL U10535 ( .A(\D_cache/cache[2][113] ), .B(n4314), .S0(net112415), .Y(
        \D_cache/n890 ) );
  MX2XL U10536 ( .A(\D_cache/cache[1][113] ), .B(n4314), .S0(net112539), .Y(
        \D_cache/n891 ) );
  MX2XL U10537 ( .A(\D_cache/cache[0][113] ), .B(n4314), .S0(net112641), .Y(
        \D_cache/n892 ) );
  MX2XL U10538 ( .A(\D_cache/cache[6][112] ), .B(n4315), .S0(net111989), .Y(
        \D_cache/n894 ) );
  MX2XL U10539 ( .A(\D_cache/cache[5][112] ), .B(n4315), .S0(net112113), .Y(
        \D_cache/n895 ) );
  MX2XL U10540 ( .A(\D_cache/cache[4][112] ), .B(n4315), .S0(net112195), .Y(
        \D_cache/n896 ) );
  MX2XL U10541 ( .A(\D_cache/cache[3][112] ), .B(n4315), .S0(net112277), .Y(
        \D_cache/n897 ) );
  MX2XL U10542 ( .A(\D_cache/cache[2][112] ), .B(n4315), .S0(net112401), .Y(
        \D_cache/n898 ) );
  MX2XL U10543 ( .A(\D_cache/cache[1][112] ), .B(n4315), .S0(net112525), .Y(
        \D_cache/n899 ) );
  MX2XL U10544 ( .A(\D_cache/cache[0][112] ), .B(n4315), .S0(net112627), .Y(
        \D_cache/n900 ) );
  MX2XL U10545 ( .A(\D_cache/cache[6][111] ), .B(n10194), .S0(net111995), .Y(
        \D_cache/n902 ) );
  MX2XL U10546 ( .A(\D_cache/cache[5][111] ), .B(n10194), .S0(net112119), .Y(
        \D_cache/n903 ) );
  MX2XL U10547 ( .A(\D_cache/cache[4][111] ), .B(n10194), .S0(net112201), .Y(
        \D_cache/n904 ) );
  MX2XL U10548 ( .A(\D_cache/cache[3][111] ), .B(n10194), .S0(net112283), .Y(
        \D_cache/n905 ) );
  MX2XL U10549 ( .A(\D_cache/cache[2][111] ), .B(n10194), .S0(net112401), .Y(
        \D_cache/n906 ) );
  MX2XL U10550 ( .A(\D_cache/cache[1][111] ), .B(n10194), .S0(net112531), .Y(
        \D_cache/n907 ) );
  MX2XL U10551 ( .A(\D_cache/cache[0][111] ), .B(n10194), .S0(net112633), .Y(
        \D_cache/n908 ) );
  MX2XL U10552 ( .A(\D_cache/cache[6][110] ), .B(n10443), .S0(net111989), .Y(
        \D_cache/n910 ) );
  MX2XL U10553 ( .A(\D_cache/cache[5][110] ), .B(n10443), .S0(net112113), .Y(
        \D_cache/n911 ) );
  MX2XL U10554 ( .A(\D_cache/cache[4][110] ), .B(n10443), .S0(net112195), .Y(
        \D_cache/n912 ) );
  MX2XL U10555 ( .A(\D_cache/cache[3][110] ), .B(n10443), .S0(net112277), .Y(
        \D_cache/n913 ) );
  MX2XL U10556 ( .A(\D_cache/cache[2][110] ), .B(n10443), .S0(net112405), .Y(
        \D_cache/n914 ) );
  MX2XL U10557 ( .A(\D_cache/cache[1][110] ), .B(n10443), .S0(net112525), .Y(
        \D_cache/n915 ) );
  MX2XL U10558 ( .A(\D_cache/cache[0][110] ), .B(n10443), .S0(net112627), .Y(
        \D_cache/n916 ) );
  MX2XL U10559 ( .A(\D_cache/cache[6][106] ), .B(n10591), .S0(net112003), .Y(
        \D_cache/n942 ) );
  MX2XL U10560 ( .A(\D_cache/cache[5][106] ), .B(n10591), .S0(net112127), .Y(
        \D_cache/n943 ) );
  MX2XL U10561 ( .A(\D_cache/cache[4][106] ), .B(n10591), .S0(net112199), .Y(
        \D_cache/n944 ) );
  MX2XL U10562 ( .A(\D_cache/cache[3][106] ), .B(n10591), .S0(net112291), .Y(
        \D_cache/n945 ) );
  MX2XL U10563 ( .A(\D_cache/cache[2][106] ), .B(n10591), .S0(net112415), .Y(
        \D_cache/n946 ) );
  MX2XL U10564 ( .A(\D_cache/cache[1][106] ), .B(n10591), .S0(net112539), .Y(
        \D_cache/n947 ) );
  MX2XL U10565 ( .A(\D_cache/cache[0][106] ), .B(n10591), .S0(net112641), .Y(
        \D_cache/n948 ) );
  MX2XL U10566 ( .A(\D_cache/cache[6][105] ), .B(n4316), .S0(net112011), .Y(
        \D_cache/n950 ) );
  MX2XL U10567 ( .A(\D_cache/cache[5][105] ), .B(n4316), .S0(net112121), .Y(
        \D_cache/n951 ) );
  MX2XL U10568 ( .A(\D_cache/cache[4][105] ), .B(n4316), .S0(net112211), .Y(
        \D_cache/n952 ) );
  MX2XL U10569 ( .A(\D_cache/cache[3][105] ), .B(n4316), .S0(net112291), .Y(
        \D_cache/n953 ) );
  MX2XL U10570 ( .A(\D_cache/cache[2][105] ), .B(n4316), .S0(net112423), .Y(
        \D_cache/n954 ) );
  MX2XL U10571 ( .A(\D_cache/cache[1][105] ), .B(n4316), .S0(net112547), .Y(
        \D_cache/n955 ) );
  MX2XL U10572 ( .A(\D_cache/cache[0][105] ), .B(n4316), .S0(net112649), .Y(
        \D_cache/n956 ) );
  MX2XL U10573 ( .A(\D_cache/cache[6][103] ), .B(n10746), .S0(net112009), .Y(
        \D_cache/n966 ) );
  MX2XL U10574 ( .A(\D_cache/cache[5][103] ), .B(n10746), .S0(net112123), .Y(
        \D_cache/n967 ) );
  MX2XL U10575 ( .A(\D_cache/cache[4][103] ), .B(n10746), .S0(net112215), .Y(
        \D_cache/n968 ) );
  MX2XL U10576 ( .A(\D_cache/cache[3][103] ), .B(n10746), .S0(net112277), .Y(
        \D_cache/n969 ) );
  MX2XL U10577 ( .A(\D_cache/cache[2][103] ), .B(n10746), .S0(net112417), .Y(
        \D_cache/n970 ) );
  MX2XL U10578 ( .A(\D_cache/cache[1][103] ), .B(n10746), .S0(net112545), .Y(
        \D_cache/n971 ) );
  MX2XL U10579 ( .A(\D_cache/cache[0][103] ), .B(n10746), .S0(net112647), .Y(
        \D_cache/n972 ) );
  MX2XL U10580 ( .A(\D_cache/cache[6][102] ), .B(n10169), .S0(net111993), .Y(
        \D_cache/n974 ) );
  MX2XL U10581 ( .A(\D_cache/cache[5][102] ), .B(n10169), .S0(net112117), .Y(
        \D_cache/n975 ) );
  MX2XL U10582 ( .A(\D_cache/cache[4][102] ), .B(n10169), .S0(net112199), .Y(
        \D_cache/n976 ) );
  MX2XL U10583 ( .A(\D_cache/cache[3][102] ), .B(n10169), .S0(net112281), .Y(
        \D_cache/n977 ) );
  MX2XL U10584 ( .A(\D_cache/cache[2][102] ), .B(n10169), .S0(net112405), .Y(
        \D_cache/n978 ) );
  MX2XL U10585 ( .A(\D_cache/cache[1][102] ), .B(n10169), .S0(net112529), .Y(
        \D_cache/n979 ) );
  MX2XL U10586 ( .A(\D_cache/cache[0][102] ), .B(n10169), .S0(net112631), .Y(
        \D_cache/n980 ) );
  MX2XL U10587 ( .A(\D_cache/cache[6][101] ), .B(n10760), .S0(net112011), .Y(
        \D_cache/n982 ) );
  MX2XL U10588 ( .A(\D_cache/cache[5][101] ), .B(n10760), .S0(net112123), .Y(
        \D_cache/n983 ) );
  MX2XL U10589 ( .A(\D_cache/cache[4][101] ), .B(n10760), .S0(net112211), .Y(
        \D_cache/n984 ) );
  MX2XL U10590 ( .A(\D_cache/cache[3][101] ), .B(n10760), .S0(net112295), .Y(
        \D_cache/n985 ) );
  MX2XL U10591 ( .A(\D_cache/cache[2][101] ), .B(n10760), .S0(net112423), .Y(
        \D_cache/n986 ) );
  MX2XL U10592 ( .A(\D_cache/cache[1][101] ), .B(n10760), .S0(net112547), .Y(
        \D_cache/n987 ) );
  MX2XL U10593 ( .A(\D_cache/cache[0][101] ), .B(n10760), .S0(net112649), .Y(
        \D_cache/n988 ) );
  MX2XL U10594 ( .A(\D_cache/cache[6][100] ), .B(n4252), .S0(net111993), .Y(
        \D_cache/n990 ) );
  MX2XL U10595 ( .A(\D_cache/cache[5][100] ), .B(n4252), .S0(net112117), .Y(
        \D_cache/n991 ) );
  MX2XL U10596 ( .A(\D_cache/cache[4][100] ), .B(n4252), .S0(net112199), .Y(
        \D_cache/n992 ) );
  MX2XL U10597 ( .A(\D_cache/cache[3][100] ), .B(n4252), .S0(net112281), .Y(
        \D_cache/n993 ) );
  MX2XL U10598 ( .A(\D_cache/cache[2][100] ), .B(n4252), .S0(net112405), .Y(
        \D_cache/n994 ) );
  MX2XL U10599 ( .A(\D_cache/cache[1][100] ), .B(n4252), .S0(net112529), .Y(
        \D_cache/n995 ) );
  MX2XL U10600 ( .A(\D_cache/cache[0][100] ), .B(n4252), .S0(net112631), .Y(
        \D_cache/n996 ) );
  MX2XL U10601 ( .A(\D_cache/cache[6][99] ), .B(n4317), .S0(net111991), .Y(
        \D_cache/n998 ) );
  MX2XL U10602 ( .A(\D_cache/cache[5][99] ), .B(n4317), .S0(net112115), .Y(
        \D_cache/n999 ) );
  MX2XL U10603 ( .A(\D_cache/cache[4][99] ), .B(n4317), .S0(net112197), .Y(
        \D_cache/n1000 ) );
  MX2XL U10604 ( .A(\D_cache/cache[3][99] ), .B(n4317), .S0(net112279), .Y(
        \D_cache/n1001 ) );
  MX2XL U10605 ( .A(\D_cache/cache[2][99] ), .B(n4317), .S0(net112403), .Y(
        \D_cache/n1002 ) );
  MX2XL U10606 ( .A(\D_cache/cache[1][99] ), .B(n4317), .S0(net112527), .Y(
        \D_cache/n1003 ) );
  MX2XL U10607 ( .A(\D_cache/cache[0][99] ), .B(n4317), .S0(net112629), .Y(
        \D_cache/n1004 ) );
  MX2XL U10608 ( .A(\D_cache/cache[6][45] ), .B(n4236), .S0(net112005), .Y(
        \D_cache/n1430 ) );
  MX2XL U10609 ( .A(\D_cache/cache[5][45] ), .B(n4236), .S0(net112129), .Y(
        \D_cache/n1431 ) );
  MX2XL U10610 ( .A(\D_cache/cache[4][45] ), .B(n4236), .S0(net112211), .Y(
        \D_cache/n1432 ) );
  MX2XL U10611 ( .A(\D_cache/cache[3][45] ), .B(n4236), .S0(net112293), .Y(
        \D_cache/n1433 ) );
  MX2XL U10612 ( .A(\D_cache/cache[2][45] ), .B(n4236), .S0(net112417), .Y(
        \D_cache/n1434 ) );
  MX2XL U10613 ( .A(\D_cache/cache[1][45] ), .B(n4236), .S0(net112541), .Y(
        \D_cache/n1435 ) );
  MX2XL U10614 ( .A(\D_cache/cache[0][45] ), .B(n4236), .S0(net112643), .Y(
        \D_cache/n1436 ) );
  MX2XL U10615 ( .A(\D_cache/cache[6][44] ), .B(n10794), .S0(net112009), .Y(
        \D_cache/n1438 ) );
  MX2XL U10616 ( .A(\D_cache/cache[5][44] ), .B(n10794), .S0(net112121), .Y(
        \D_cache/n1439 ) );
  MX2XL U10617 ( .A(\D_cache/cache[4][44] ), .B(n10794), .S0(net112215), .Y(
        \D_cache/n1440 ) );
  MX2XL U10618 ( .A(\D_cache/cache[3][44] ), .B(n10794), .S0(net112281), .Y(
        \D_cache/n1441 ) );
  MX2XL U10619 ( .A(\D_cache/cache[2][44] ), .B(n10794), .S0(net112419), .Y(
        \D_cache/n1442 ) );
  MX2XL U10620 ( .A(\D_cache/cache[1][44] ), .B(n10794), .S0(net112545), .Y(
        \D_cache/n1443 ) );
  MX2XL U10621 ( .A(\D_cache/cache[0][44] ), .B(n10794), .S0(net112647), .Y(
        \D_cache/n1444 ) );
  MX2XL U10622 ( .A(\D_cache/cache[6][43] ), .B(n4239), .S0(net112011), .Y(
        \D_cache/n1446 ) );
  MX2XL U10623 ( .A(\D_cache/cache[5][43] ), .B(n4239), .S0(net112123), .Y(
        \D_cache/n1447 ) );
  MX2XL U10624 ( .A(\D_cache/cache[4][43] ), .B(n4239), .S0(net112211), .Y(
        \D_cache/n1448 ) );
  MX2XL U10625 ( .A(\D_cache/cache[3][43] ), .B(n4239), .S0(net112289), .Y(
        \D_cache/n1449 ) );
  MX2XL U10626 ( .A(\D_cache/cache[2][43] ), .B(n4239), .S0(net112423), .Y(
        \D_cache/n1450 ) );
  MX2XL U10627 ( .A(\D_cache/cache[1][43] ), .B(n4239), .S0(net112547), .Y(
        \D_cache/n1451 ) );
  MX2XL U10628 ( .A(\D_cache/cache[0][43] ), .B(n4239), .S0(net112649), .Y(
        \D_cache/n1452 ) );
  MX2XL U10629 ( .A(\D_cache/cache[6][40] ), .B(n4237), .S0(net112005), .Y(
        \D_cache/n1470 ) );
  MX2XL U10630 ( .A(\D_cache/cache[5][40] ), .B(n4237), .S0(net112129), .Y(
        \D_cache/n1471 ) );
  MX2XL U10631 ( .A(\D_cache/cache[4][40] ), .B(n4237), .S0(net112211), .Y(
        \D_cache/n1472 ) );
  MX2XL U10632 ( .A(\D_cache/cache[3][40] ), .B(n4237), .S0(net112293), .Y(
        \D_cache/n1473 ) );
  MX2XL U10633 ( .A(\D_cache/cache[2][40] ), .B(n4237), .S0(net112417), .Y(
        \D_cache/n1474 ) );
  MX2XL U10634 ( .A(\D_cache/cache[1][40] ), .B(n4237), .S0(net112541), .Y(
        \D_cache/n1475 ) );
  MX2XL U10635 ( .A(\D_cache/cache[0][40] ), .B(n4237), .S0(net112643), .Y(
        \D_cache/n1476 ) );
  MX2XL U10636 ( .A(\D_cache/cache[6][34] ), .B(n4240), .S0(net111995), .Y(
        \D_cache/n1518 ) );
  MX2XL U10637 ( .A(\D_cache/cache[5][34] ), .B(n4240), .S0(net112131), .Y(
        \D_cache/n1519 ) );
  MX2XL U10638 ( .A(\D_cache/cache[4][34] ), .B(n4240), .S0(net112213), .Y(
        \D_cache/n1520 ) );
  MX2XL U10639 ( .A(\D_cache/cache[3][34] ), .B(n4240), .S0(net112295), .Y(
        \D_cache/n1521 ) );
  MX2XL U10640 ( .A(\D_cache/cache[2][34] ), .B(n4240), .S0(net112419), .Y(
        \D_cache/n1522 ) );
  MX2XL U10641 ( .A(\D_cache/cache[1][34] ), .B(n4240), .S0(net112543), .Y(
        \D_cache/n1523 ) );
  MX2XL U10642 ( .A(\D_cache/cache[0][34] ), .B(n4240), .S0(net112645), .Y(
        \D_cache/n1524 ) );
  MX2XL U10643 ( .A(\D_cache/cache[6][33] ), .B(n4238), .S0(net112005), .Y(
        \D_cache/n1526 ) );
  MX2XL U10644 ( .A(\D_cache/cache[5][33] ), .B(n4238), .S0(net112129), .Y(
        \D_cache/n1527 ) );
  MX2XL U10645 ( .A(\D_cache/cache[4][33] ), .B(n4238), .S0(net112211), .Y(
        \D_cache/n1528 ) );
  MX2XL U10646 ( .A(\D_cache/cache[3][33] ), .B(n4238), .S0(net112293), .Y(
        \D_cache/n1529 ) );
  MX2XL U10647 ( .A(\D_cache/cache[2][33] ), .B(n4238), .S0(net112417), .Y(
        \D_cache/n1530 ) );
  MX2XL U10648 ( .A(\D_cache/cache[1][33] ), .B(n4238), .S0(net112541), .Y(
        \D_cache/n1531 ) );
  MX2XL U10649 ( .A(\D_cache/cache[0][33] ), .B(n4238), .S0(net112643), .Y(
        \D_cache/n1532 ) );
  MX2XL U10650 ( .A(\D_cache/cache[6][32] ), .B(n10856), .S0(net111993), .Y(
        \D_cache/n1534 ) );
  MX2XL U10651 ( .A(\D_cache/cache[5][32] ), .B(n10856), .S0(net112131), .Y(
        \D_cache/n1535 ) );
  MX2XL U10652 ( .A(\D_cache/cache[4][32] ), .B(n10856), .S0(net112211), .Y(
        \D_cache/n1536 ) );
  MX2XL U10653 ( .A(\D_cache/cache[3][32] ), .B(n10856), .S0(net112295), .Y(
        \D_cache/n1537 ) );
  MX2XL U10654 ( .A(\D_cache/cache[2][32] ), .B(n10856), .S0(net112419), .Y(
        \D_cache/n1538 ) );
  MX2XL U10655 ( .A(\D_cache/cache[1][32] ), .B(n10856), .S0(net112543), .Y(
        \D_cache/n1539 ) );
  MX2XL U10656 ( .A(\D_cache/cache[0][32] ), .B(n10856), .S0(net112645), .Y(
        \D_cache/n1540 ) );
  MX2XL U10657 ( .A(\D_cache/cache[6][13] ), .B(n4232), .S0(net112005), .Y(
        \D_cache/n1686 ) );
  MX2XL U10658 ( .A(\D_cache/cache[5][13] ), .B(n4232), .S0(net112129), .Y(
        \D_cache/n1687 ) );
  MX2XL U10659 ( .A(\D_cache/cache[4][13] ), .B(n4232), .S0(net112211), .Y(
        \D_cache/n1688 ) );
  MX2XL U10660 ( .A(\D_cache/cache[3][13] ), .B(n4232), .S0(net112293), .Y(
        \D_cache/n1689 ) );
  MX2XL U10661 ( .A(\D_cache/cache[2][13] ), .B(n4232), .S0(net112417), .Y(
        \D_cache/n1690 ) );
  MX2XL U10662 ( .A(\D_cache/cache[1][13] ), .B(n4232), .S0(net112541), .Y(
        \D_cache/n1691 ) );
  MX2XL U10663 ( .A(\D_cache/cache[0][13] ), .B(n4232), .S0(net112643), .Y(
        \D_cache/n1692 ) );
  MX2XL U10664 ( .A(\D_cache/cache[6][12] ), .B(n4233), .S0(net112011), .Y(
        \D_cache/n1694 ) );
  MX2XL U10665 ( .A(\D_cache/cache[5][12] ), .B(n4233), .S0(net112121), .Y(
        \D_cache/n1695 ) );
  MX2XL U10666 ( .A(\D_cache/cache[4][12] ), .B(n4233), .S0(net112211), .Y(
        \D_cache/n1696 ) );
  MX2XL U10667 ( .A(\D_cache/cache[3][12] ), .B(n4233), .S0(net112291), .Y(
        \D_cache/n1697 ) );
  MX2XL U10668 ( .A(\D_cache/cache[2][12] ), .B(n4233), .S0(net112423), .Y(
        \D_cache/n1698 ) );
  MX2XL U10669 ( .A(\D_cache/cache[1][12] ), .B(n4233), .S0(net112547), .Y(
        \D_cache/n1699 ) );
  MX2XL U10670 ( .A(\D_cache/cache[0][12] ), .B(n4233), .S0(net112649), .Y(
        \D_cache/n1700 ) );
  MX2XL U10671 ( .A(\D_cache/cache[6][11] ), .B(n4234), .S0(net112011), .Y(
        \D_cache/n1702 ) );
  MX2XL U10672 ( .A(\D_cache/cache[5][11] ), .B(n4234), .S0(net112123), .Y(
        \D_cache/n1703 ) );
  MX2XL U10673 ( .A(\D_cache/cache[4][11] ), .B(n4234), .S0(net112211), .Y(
        \D_cache/n1704 ) );
  MX2XL U10674 ( .A(\D_cache/cache[3][11] ), .B(n4234), .S0(net112289), .Y(
        \D_cache/n1705 ) );
  MX2XL U10675 ( .A(\D_cache/cache[2][11] ), .B(n4234), .S0(net112423), .Y(
        \D_cache/n1706 ) );
  MX2XL U10676 ( .A(\D_cache/cache[1][11] ), .B(n4234), .S0(net112547), .Y(
        \D_cache/n1707 ) );
  MX2XL U10677 ( .A(\D_cache/cache[0][11] ), .B(n4234), .S0(net112649), .Y(
        \D_cache/n1708 ) );
  MX2XL U10678 ( .A(\D_cache/cache[6][8] ), .B(n10819), .S0(net112005), .Y(
        \D_cache/n1726 ) );
  MX2XL U10679 ( .A(\D_cache/cache[5][8] ), .B(n10819), .S0(net112129), .Y(
        \D_cache/n1727 ) );
  MX2XL U10680 ( .A(\D_cache/cache[4][8] ), .B(n10819), .S0(net112211), .Y(
        \D_cache/n1728 ) );
  MX2XL U10681 ( .A(\D_cache/cache[3][8] ), .B(n10819), .S0(net112293), .Y(
        \D_cache/n1729 ) );
  MX2XL U10682 ( .A(\D_cache/cache[2][8] ), .B(n10819), .S0(net112417), .Y(
        \D_cache/n1730 ) );
  MX2XL U10683 ( .A(\D_cache/cache[1][8] ), .B(n10819), .S0(net112541), .Y(
        \D_cache/n1731 ) );
  MX2XL U10684 ( .A(\D_cache/cache[0][8] ), .B(n10819), .S0(net112643), .Y(
        \D_cache/n1732 ) );
  MX2XL U10685 ( .A(\D_cache/cache[6][2] ), .B(n4235), .S0(net112009), .Y(
        \D_cache/n1774 ) );
  MX2XL U10686 ( .A(\D_cache/cache[5][2] ), .B(n4235), .S0(net112131), .Y(
        \D_cache/n1775 ) );
  MX2XL U10687 ( .A(\D_cache/cache[4][2] ), .B(n4235), .S0(net112213), .Y(
        \D_cache/n1776 ) );
  MX2XL U10688 ( .A(\D_cache/cache[3][2] ), .B(n4235), .S0(net112295), .Y(
        \D_cache/n1777 ) );
  MX2XL U10689 ( .A(\D_cache/cache[2][2] ), .B(n4235), .S0(net112419), .Y(
        \D_cache/n1778 ) );
  MX2XL U10690 ( .A(\D_cache/cache[1][2] ), .B(n4235), .S0(net112543), .Y(
        \D_cache/n1779 ) );
  MX2XL U10691 ( .A(\D_cache/cache[0][2] ), .B(n4235), .S0(net112645), .Y(
        \D_cache/n1780 ) );
  MX2XL U10692 ( .A(\D_cache/cache[6][1] ), .B(n10840), .S0(net112005), .Y(
        \D_cache/n1782 ) );
  MX2XL U10693 ( .A(\D_cache/cache[5][1] ), .B(n10840), .S0(net112129), .Y(
        \D_cache/n1783 ) );
  MX2XL U10694 ( .A(\D_cache/cache[4][1] ), .B(n10840), .S0(net112211), .Y(
        \D_cache/n1784 ) );
  MX2XL U10695 ( .A(\D_cache/cache[3][1] ), .B(n10840), .S0(net112293), .Y(
        \D_cache/n1785 ) );
  MX2XL U10696 ( .A(\D_cache/cache[2][1] ), .B(n10840), .S0(net112417), .Y(
        \D_cache/n1786 ) );
  MX2XL U10697 ( .A(\D_cache/cache[1][1] ), .B(n10840), .S0(net112541), .Y(
        \D_cache/n1787 ) );
  MX2XL U10698 ( .A(\D_cache/cache[0][1] ), .B(n10840), .S0(net112643), .Y(
        \D_cache/n1788 ) );
  MX2XL U10699 ( .A(\D_cache/cache[6][0] ), .B(n10853), .S0(net111995), .Y(
        \D_cache/n1789 ) );
  MX2XL U10700 ( .A(\D_cache/cache[5][0] ), .B(n10853), .S0(net112131), .Y(
        \D_cache/n1790 ) );
  MX2XL U10701 ( .A(\D_cache/cache[4][0] ), .B(n10853), .S0(net112211), .Y(
        \D_cache/n1791 ) );
  MX2XL U10702 ( .A(\D_cache/cache[3][0] ), .B(n10853), .S0(net112295), .Y(
        \D_cache/n1792 ) );
  MX2XL U10703 ( .A(\D_cache/cache[2][0] ), .B(n10853), .S0(net112419), .Y(
        \D_cache/n1793 ) );
  MX2XL U10704 ( .A(\D_cache/cache[1][0] ), .B(n10853), .S0(net112543), .Y(
        \D_cache/n1794 ) );
  MX2XL U10705 ( .A(\D_cache/cache[0][0] ), .B(n10853), .S0(net112645), .Y(
        \D_cache/n1795 ) );
  MX2XL U10706 ( .A(\D_cache/cache[6][95] ), .B(n4245), .S0(net111993), .Y(
        \D_cache/n1030 ) );
  MX2XL U10707 ( .A(\D_cache/cache[5][95] ), .B(n4245), .S0(net112123), .Y(
        \D_cache/n1031 ) );
  MX2XL U10708 ( .A(\D_cache/cache[4][95] ), .B(n4245), .S0(net112201), .Y(
        \D_cache/n1032 ) );
  MX2XL U10709 ( .A(\D_cache/cache[3][95] ), .B(n4245), .S0(net112285), .Y(
        \D_cache/n1033 ) );
  MX2XL U10710 ( .A(\D_cache/cache[2][95] ), .B(n4245), .S0(net112409), .Y(
        \D_cache/n1034 ) );
  MX2XL U10711 ( .A(\D_cache/cache[1][95] ), .B(n4245), .S0(net112533), .Y(
        \D_cache/n1035 ) );
  MX2XL U10712 ( .A(\D_cache/cache[0][95] ), .B(n4245), .S0(net112635), .Y(
        \D_cache/n1036 ) );
  MX2XL U10713 ( .A(\D_cache/cache[6][77] ), .B(n4241), .S0(net112005), .Y(
        \D_cache/n1174 ) );
  MX2XL U10714 ( .A(\D_cache/cache[5][77] ), .B(n4241), .S0(net112129), .Y(
        \D_cache/n1175 ) );
  MX2XL U10715 ( .A(\D_cache/cache[4][77] ), .B(n4241), .S0(net112211), .Y(
        \D_cache/n1176 ) );
  MX2XL U10716 ( .A(\D_cache/cache[3][77] ), .B(n4241), .S0(net112293), .Y(
        \D_cache/n1177 ) );
  MX2XL U10717 ( .A(\D_cache/cache[2][77] ), .B(n4241), .S0(net112417), .Y(
        \D_cache/n1178 ) );
  MX2XL U10718 ( .A(\D_cache/cache[1][77] ), .B(n4241), .S0(net112541), .Y(
        \D_cache/n1179 ) );
  MX2XL U10719 ( .A(\D_cache/cache[0][77] ), .B(n4241), .S0(net112643), .Y(
        \D_cache/n1180 ) );
  MX2XL U10720 ( .A(\D_cache/cache[6][76] ), .B(n10800), .S0(net112005), .Y(
        \D_cache/n1182 ) );
  MX2XL U10721 ( .A(\D_cache/cache[5][76] ), .B(n10800), .S0(net112129), .Y(
        \D_cache/n1183 ) );
  MX2XL U10722 ( .A(\D_cache/cache[4][76] ), .B(n10800), .S0(net112211), .Y(
        \D_cache/n1184 ) );
  MX2XL U10723 ( .A(\D_cache/cache[3][76] ), .B(n10800), .S0(net112293), .Y(
        \D_cache/n1185 ) );
  MX2XL U10724 ( .A(\D_cache/cache[2][76] ), .B(n10800), .S0(net112417), .Y(
        \D_cache/n1186 ) );
  MX2XL U10725 ( .A(\D_cache/cache[1][76] ), .B(n10800), .S0(net112541), .Y(
        \D_cache/n1187 ) );
  MX2XL U10726 ( .A(\D_cache/cache[0][76] ), .B(n10800), .S0(net112643), .Y(
        \D_cache/n1188 ) );
  MX2XL U10727 ( .A(\D_cache/cache[6][75] ), .B(n4244), .S0(net112011), .Y(
        \D_cache/n1190 ) );
  MX2XL U10728 ( .A(\D_cache/cache[5][75] ), .B(n4244), .S0(net112121), .Y(
        \D_cache/n1191 ) );
  MX2XL U10729 ( .A(\D_cache/cache[4][75] ), .B(n4244), .S0(net112211), .Y(
        \D_cache/n1192 ) );
  MX2XL U10730 ( .A(\D_cache/cache[3][75] ), .B(n4244), .S0(net112291), .Y(
        \D_cache/n1193 ) );
  MX2XL U10731 ( .A(\D_cache/cache[2][75] ), .B(n4244), .S0(net112423), .Y(
        \D_cache/n1194 ) );
  MX2XL U10732 ( .A(\D_cache/cache[1][75] ), .B(n4244), .S0(net112547), .Y(
        \D_cache/n1195 ) );
  MX2XL U10733 ( .A(\D_cache/cache[0][75] ), .B(n4244), .S0(net112649), .Y(
        \D_cache/n1196 ) );
  MX2XL U10734 ( .A(\D_cache/cache[6][72] ), .B(n4242), .S0(net112005), .Y(
        \D_cache/n1214 ) );
  MX2XL U10735 ( .A(\D_cache/cache[5][72] ), .B(n4242), .S0(net112129), .Y(
        \D_cache/n1215 ) );
  MX2XL U10736 ( .A(\D_cache/cache[4][72] ), .B(n4242), .S0(net112211), .Y(
        \D_cache/n1216 ) );
  MX2XL U10737 ( .A(\D_cache/cache[3][72] ), .B(n4242), .S0(net112293), .Y(
        \D_cache/n1217 ) );
  MX2XL U10738 ( .A(\D_cache/cache[2][72] ), .B(n4242), .S0(net112417), .Y(
        \D_cache/n1218 ) );
  MX2XL U10739 ( .A(\D_cache/cache[1][72] ), .B(n4242), .S0(net112541), .Y(
        \D_cache/n1219 ) );
  MX2XL U10740 ( .A(\D_cache/cache[0][72] ), .B(n4242), .S0(net112643), .Y(
        \D_cache/n1220 ) );
  MX2XL U10741 ( .A(\D_cache/cache[6][66] ), .B(n4246), .S0(net112005), .Y(
        \D_cache/n1262 ) );
  MX2XL U10742 ( .A(\D_cache/cache[5][66] ), .B(n4246), .S0(net112131), .Y(
        \D_cache/n1263 ) );
  MX2XL U10743 ( .A(\D_cache/cache[4][66] ), .B(n4246), .S0(net112213), .Y(
        \D_cache/n1264 ) );
  MX2XL U10744 ( .A(\D_cache/cache[3][66] ), .B(n4246), .S0(net112295), .Y(
        \D_cache/n1265 ) );
  MX2XL U10745 ( .A(\D_cache/cache[2][66] ), .B(n4246), .S0(net112419), .Y(
        \D_cache/n1266 ) );
  MX2XL U10746 ( .A(\D_cache/cache[1][66] ), .B(n4246), .S0(net112543), .Y(
        \D_cache/n1267 ) );
  MX2XL U10747 ( .A(\D_cache/cache[0][66] ), .B(n4246), .S0(net112645), .Y(
        \D_cache/n1268 ) );
  MX2XL U10748 ( .A(\D_cache/cache[6][65] ), .B(n4243), .S0(net111991), .Y(
        \D_cache/n1270 ) );
  MX2XL U10749 ( .A(\D_cache/cache[5][65] ), .B(n4243), .S0(net112131), .Y(
        \D_cache/n1271 ) );
  MX2XL U10750 ( .A(\D_cache/cache[4][65] ), .B(n4243), .S0(net112213), .Y(
        \D_cache/n1272 ) );
  MX2XL U10751 ( .A(\D_cache/cache[3][65] ), .B(n4243), .S0(net112295), .Y(
        \D_cache/n1273 ) );
  MX2XL U10752 ( .A(\D_cache/cache[2][65] ), .B(n4243), .S0(net112419), .Y(
        \D_cache/n1274 ) );
  MX2XL U10753 ( .A(\D_cache/cache[1][65] ), .B(n4243), .S0(net112543), .Y(
        \D_cache/n1275 ) );
  MX2XL U10754 ( .A(\D_cache/cache[0][65] ), .B(n4243), .S0(net112645), .Y(
        \D_cache/n1276 ) );
  MX2XL U10755 ( .A(\D_cache/cache[6][64] ), .B(n10862), .S0(net111993), .Y(
        \D_cache/n1278 ) );
  MX2XL U10756 ( .A(\D_cache/cache[5][64] ), .B(n10862), .S0(net112131), .Y(
        \D_cache/n1279 ) );
  MX2XL U10757 ( .A(\D_cache/cache[4][64] ), .B(n10862), .S0(net112211), .Y(
        \D_cache/n1280 ) );
  MX2XL U10758 ( .A(\D_cache/cache[3][64] ), .B(n10862), .S0(net112295), .Y(
        \D_cache/n1281 ) );
  MX2XL U10759 ( .A(\D_cache/cache[2][64] ), .B(n10862), .S0(net112419), .Y(
        \D_cache/n1282 ) );
  MX2XL U10760 ( .A(\D_cache/cache[1][64] ), .B(n10862), .S0(net112543), .Y(
        \D_cache/n1283 ) );
  MX2XL U10761 ( .A(\D_cache/cache[0][64] ), .B(n10862), .S0(net112645), .Y(
        \D_cache/n1284 ) );
  MX2XL U10762 ( .A(\D_cache/cache[6][109] ), .B(n10809), .S0(net112005), .Y(
        \D_cache/n918 ) );
  MX2XL U10763 ( .A(\D_cache/cache[5][109] ), .B(n10809), .S0(net112129), .Y(
        \D_cache/n919 ) );
  MX2XL U10764 ( .A(\D_cache/cache[4][109] ), .B(n10809), .S0(net112211), .Y(
        \D_cache/n920 ) );
  MX2XL U10765 ( .A(\D_cache/cache[3][109] ), .B(n10809), .S0(net112293), .Y(
        \D_cache/n921 ) );
  MX2XL U10766 ( .A(\D_cache/cache[2][109] ), .B(n10809), .S0(net112417), .Y(
        \D_cache/n922 ) );
  MX2XL U10767 ( .A(\D_cache/cache[1][109] ), .B(n10809), .S0(net112541), .Y(
        \D_cache/n923 ) );
  MX2XL U10768 ( .A(\D_cache/cache[0][109] ), .B(n10809), .S0(net112643), .Y(
        \D_cache/n924 ) );
  MX2XL U10769 ( .A(\D_cache/cache[6][108] ), .B(n10797), .S0(net112005), .Y(
        \D_cache/n926 ) );
  MX2XL U10770 ( .A(\D_cache/cache[5][108] ), .B(n10797), .S0(net112129), .Y(
        \D_cache/n927 ) );
  MX2XL U10771 ( .A(\D_cache/cache[4][108] ), .B(n10797), .S0(net112211), .Y(
        \D_cache/n928 ) );
  MX2XL U10772 ( .A(\D_cache/cache[3][108] ), .B(n10797), .S0(net112293), .Y(
        \D_cache/n929 ) );
  MX2XL U10773 ( .A(\D_cache/cache[2][108] ), .B(n10797), .S0(net112417), .Y(
        \D_cache/n930 ) );
  MX2XL U10774 ( .A(\D_cache/cache[1][108] ), .B(n10797), .S0(net112541), .Y(
        \D_cache/n931 ) );
  MX2XL U10775 ( .A(\D_cache/cache[6][107] ), .B(n10785), .S0(net112011), .Y(
        \D_cache/n934 ) );
  MX2XL U10776 ( .A(\D_cache/cache[5][107] ), .B(n10785), .S0(net112121), .Y(
        \D_cache/n935 ) );
  MX2XL U10777 ( .A(\D_cache/cache[3][107] ), .B(n10785), .S0(net112293), .Y(
        \D_cache/n937 ) );
  MX2XL U10778 ( .A(\D_cache/cache[2][107] ), .B(n10785), .S0(net112423), .Y(
        \D_cache/n938 ) );
  MX2XL U10779 ( .A(\D_cache/cache[1][107] ), .B(n10785), .S0(net112547), .Y(
        \D_cache/n939 ) );
  MX2XL U10780 ( .A(\D_cache/cache[0][107] ), .B(n10785), .S0(net112649), .Y(
        \D_cache/n940 ) );
  MX2XL U10781 ( .A(\D_cache/cache[6][104] ), .B(n10825), .S0(net112005), .Y(
        \D_cache/n958 ) );
  MX2XL U10782 ( .A(\D_cache/cache[5][104] ), .B(n10825), .S0(net112129), .Y(
        \D_cache/n959 ) );
  MX2XL U10783 ( .A(\D_cache/cache[4][104] ), .B(n10825), .S0(net112211), .Y(
        \D_cache/n960 ) );
  MX2XL U10784 ( .A(\D_cache/cache[3][104] ), .B(n10825), .S0(net112293), .Y(
        \D_cache/n961 ) );
  MX2XL U10785 ( .A(\D_cache/cache[2][104] ), .B(n10825), .S0(net112417), .Y(
        \D_cache/n962 ) );
  MX2XL U10786 ( .A(\D_cache/cache[1][104] ), .B(n10825), .S0(net112541), .Y(
        \D_cache/n963 ) );
  MX2XL U10787 ( .A(\D_cache/cache[0][104] ), .B(n10825), .S0(net112643), .Y(
        \D_cache/n964 ) );
  MX2XL U10788 ( .A(\D_cache/cache[6][98] ), .B(n11177), .S0(net112005), .Y(
        \D_cache/n1006 ) );
  MX2XL U10789 ( .A(\D_cache/cache[5][98] ), .B(n11177), .S0(net112131), .Y(
        \D_cache/n1007 ) );
  MX2XL U10790 ( .A(\D_cache/cache[4][98] ), .B(n11177), .S0(net112211), .Y(
        \D_cache/n1008 ) );
  MX2XL U10791 ( .A(\D_cache/cache[3][98] ), .B(n11177), .S0(net112295), .Y(
        \D_cache/n1009 ) );
  MX2XL U10792 ( .A(\D_cache/cache[2][98] ), .B(n11177), .S0(net112419), .Y(
        \D_cache/n1010 ) );
  MX2XL U10793 ( .A(\D_cache/cache[1][98] ), .B(n11177), .S0(net112543), .Y(
        \D_cache/n1011 ) );
  MX2XL U10794 ( .A(\D_cache/cache[0][98] ), .B(n11177), .S0(net112645), .Y(
        \D_cache/n1012 ) );
  MX2XL U10795 ( .A(\D_cache/cache[6][97] ), .B(n10846), .S0(net112003), .Y(
        \D_cache/n1014 ) );
  MX2XL U10796 ( .A(\D_cache/cache[5][97] ), .B(n10846), .S0(net112127), .Y(
        \D_cache/n1015 ) );
  MX2XL U10797 ( .A(\D_cache/cache[4][97] ), .B(n10846), .S0(net112201), .Y(
        \D_cache/n1016 ) );
  MX2XL U10798 ( .A(\D_cache/cache[3][97] ), .B(n10846), .S0(net112291), .Y(
        \D_cache/n1017 ) );
  MX2XL U10799 ( .A(\D_cache/cache[2][97] ), .B(n10846), .S0(net112415), .Y(
        \D_cache/n1018 ) );
  MX2XL U10800 ( .A(\D_cache/cache[1][97] ), .B(n10846), .S0(net112539), .Y(
        \D_cache/n1019 ) );
  MX2XL U10801 ( .A(\D_cache/cache[0][97] ), .B(n10846), .S0(net112641), .Y(
        \D_cache/n1020 ) );
  MX2XL U10802 ( .A(\D_cache/cache[6][96] ), .B(n10859), .S0(net111991), .Y(
        \D_cache/n1022 ) );
  MX2XL U10803 ( .A(\D_cache/cache[5][96] ), .B(n10859), .S0(net112131), .Y(
        \D_cache/n1023 ) );
  MX2XL U10804 ( .A(\D_cache/cache[4][96] ), .B(n10859), .S0(net112211), .Y(
        \D_cache/n1024 ) );
  MX2XL U10805 ( .A(\D_cache/cache[3][96] ), .B(n10859), .S0(net112295), .Y(
        \D_cache/n1025 ) );
  MX2XL U10806 ( .A(\D_cache/cache[2][96] ), .B(n10859), .S0(net112419), .Y(
        \D_cache/n1026 ) );
  MX2XL U10807 ( .A(\D_cache/cache[1][96] ), .B(n10859), .S0(net112543), .Y(
        \D_cache/n1027 ) );
  MX2XL U10808 ( .A(\D_cache/cache[0][96] ), .B(n10859), .S0(net112645), .Y(
        \D_cache/n1028 ) );
  OA22X1 U10809 ( .A0(\i_MIPS/Register/register[17][22] ), .A1(n4835), .B0(
        \i_MIPS/Register/register[25][22] ), .B1(n4831), .Y(n8000) );
  OA22X1 U10810 ( .A0(\i_MIPS/Register/register[17][16] ), .A1(n4835), .B0(
        \i_MIPS/Register/register[25][16] ), .B1(n4831), .Y(n8183) );
  OA22X1 U10811 ( .A0(\i_MIPS/Register/register[17][10] ), .A1(n4833), .B0(
        \i_MIPS/Register/register[25][10] ), .B1(n4830), .Y(n7223) );
  OA22XL U10812 ( .A0(net112673), .A1(n1581), .B0(net112571), .B1(n3194), .Y(
        net105008) );
  OA22XL U10813 ( .A0(net112673), .A1(n1582), .B0(net112571), .B1(n3195), .Y(
        net105020) );
  MXI2X1 U10814 ( .A(\i_MIPS/Pred_2bit/n1 ), .B(n4699), .S0(n4700), .Y(
        \i_MIPS/Pred_2bit/n7 ) );
  CLKMX2X2 U10815 ( .A(\D_cache/cache[7][153] ), .B(n10519), .S0(net111867), 
        .Y(\D_cache/n565 ) );
  CLKMX2X2 U10816 ( .A(\D_cache/cache[6][153] ), .B(n10519), .S0(net111991), 
        .Y(\D_cache/n566 ) );
  CLKMX2X2 U10817 ( .A(\D_cache/cache[5][153] ), .B(n10519), .S0(net112115), 
        .Y(\D_cache/n567 ) );
  CLKMX2X2 U10818 ( .A(\D_cache/cache[4][153] ), .B(n10519), .S0(net112197), 
        .Y(\D_cache/n568 ) );
  CLKMX2X2 U10819 ( .A(\D_cache/cache[3][153] ), .B(n10519), .S0(net112279), 
        .Y(\D_cache/n569 ) );
  CLKMX2X2 U10820 ( .A(\D_cache/cache[2][153] ), .B(n10519), .S0(net112403), 
        .Y(\D_cache/n570 ) );
  CLKMX2X2 U10821 ( .A(\D_cache/cache[1][153] ), .B(n10519), .S0(net112527), 
        .Y(\D_cache/n571 ) );
  CLKMX2X2 U10822 ( .A(\D_cache/cache[0][153] ), .B(n10519), .S0(net112643), 
        .Y(\D_cache/n572 ) );
  MXI2XL U10823 ( .A(n4705), .B(n10132), .S0(n5509), .Y(\i_MIPS/n475 ) );
  MXI2XL U10824 ( .A(n4715), .B(n10129), .S0(n5510), .Y(\i_MIPS/n473 ) );
  MX2XL U10825 ( .A(\i_MIPS/Reg_W[1] ), .B(n10131), .S0(n5511), .Y(
        \i_MIPS/n476 ) );
  MXI2X1 U10826 ( .A(n177), .B(\i_MIPS/n219 ), .S0(n5508), .Y(\i_MIPS/n505 )
         );
  MX2XL U10827 ( .A(\D_cache/cache[6][145] ), .B(n121), .S0(net111999), .Y(
        \D_cache/n630 ) );
  MX2XL U10828 ( .A(\D_cache/cache[5][145] ), .B(n121), .S0(net112121), .Y(
        \D_cache/n631 ) );
  MX2XL U10829 ( .A(\D_cache/cache[4][145] ), .B(n121), .S0(net112215), .Y(
        \D_cache/n632 ) );
  MX2XL U10830 ( .A(\D_cache/cache[3][145] ), .B(n121), .S0(net112281), .Y(
        \D_cache/n633 ) );
  MX2XL U10831 ( .A(\D_cache/cache[2][145] ), .B(n121), .S0(net112411), .Y(
        \D_cache/n634 ) );
  MX2XL U10832 ( .A(\D_cache/cache[1][145] ), .B(n121), .S0(net112535), .Y(
        \D_cache/n635 ) );
  MX2XL U10833 ( .A(\D_cache/cache[0][145] ), .B(n121), .S0(net112637), .Y(
        \D_cache/n636 ) );
  MX2XL U10834 ( .A(\D_cache/cache[7][130] ), .B(n131), .S0(net111885), .Y(
        \D_cache/n749 ) );
  MX2XL U10835 ( .A(\D_cache/cache[6][130] ), .B(n131), .S0(net112009), .Y(
        \D_cache/n750 ) );
  MX2XL U10836 ( .A(\D_cache/cache[5][130] ), .B(n131), .S0(net112121), .Y(
        \D_cache/n751 ) );
  MX2XL U10837 ( .A(\D_cache/cache[4][130] ), .B(n131), .S0(net112215), .Y(
        \D_cache/n752 ) );
  MX2XL U10838 ( .A(\D_cache/cache[3][130] ), .B(n131), .S0(net112279), .Y(
        \D_cache/n753 ) );
  MX2XL U10839 ( .A(\D_cache/cache[2][130] ), .B(n131), .S0(net112417), .Y(
        \D_cache/n754 ) );
  MX2XL U10840 ( .A(\D_cache/cache[1][130] ), .B(n131), .S0(net112545), .Y(
        \D_cache/n755 ) );
  MX2XL U10841 ( .A(\D_cache/cache[0][130] ), .B(n131), .S0(net112647), .Y(
        \D_cache/n756 ) );
  MX2XL U10842 ( .A(\D_cache/cache[6][143] ), .B(n143), .S0(net111995), .Y(
        \D_cache/n646 ) );
  MX2XL U10843 ( .A(\D_cache/cache[5][143] ), .B(n143), .S0(net112121), .Y(
        \D_cache/n647 ) );
  MX2XL U10844 ( .A(\D_cache/cache[4][143] ), .B(n143), .S0(net112197), .Y(
        \D_cache/n648 ) );
  MX2XL U10845 ( .A(\D_cache/cache[3][143] ), .B(n143), .S0(net112285), .Y(
        \D_cache/n649 ) );
  MX2XL U10846 ( .A(\D_cache/cache[2][143] ), .B(n143), .S0(net112409), .Y(
        \D_cache/n650 ) );
  MX2XL U10847 ( .A(\D_cache/cache[1][143] ), .B(n143), .S0(net112533), .Y(
        \D_cache/n651 ) );
  MX2XL U10848 ( .A(\D_cache/cache[0][143] ), .B(n143), .S0(net112635), .Y(
        \D_cache/n652 ) );
  MX2XL U10849 ( .A(\D_cache/cache[6][147] ), .B(n122), .S0(net111995), .Y(
        \D_cache/n614 ) );
  MX2XL U10850 ( .A(\D_cache/cache[5][147] ), .B(n122), .S0(net112119), .Y(
        \D_cache/n615 ) );
  MX2XL U10851 ( .A(\D_cache/cache[4][147] ), .B(n122), .S0(net112201), .Y(
        \D_cache/n616 ) );
  MX2XL U10852 ( .A(\D_cache/cache[3][147] ), .B(n122), .S0(net112283), .Y(
        \D_cache/n617 ) );
  MX2XL U10853 ( .A(\D_cache/cache[2][147] ), .B(n122), .S0(net112405), .Y(
        \D_cache/n618 ) );
  MX2XL U10854 ( .A(\D_cache/cache[1][147] ), .B(n122), .S0(net112531), .Y(
        \D_cache/n619 ) );
  MX2XL U10855 ( .A(\D_cache/cache[0][147] ), .B(n122), .S0(net112633), .Y(
        \D_cache/n620 ) );
  MX2XL U10856 ( .A(\D_cache/cache[7][131] ), .B(n134), .S0(net111885), .Y(
        \D_cache/n741 ) );
  MX2XL U10857 ( .A(\D_cache/cache[6][131] ), .B(n134), .S0(net112009), .Y(
        \D_cache/n742 ) );
  MX2XL U10858 ( .A(\D_cache/cache[5][131] ), .B(n134), .S0(net112123), .Y(
        \D_cache/n743 ) );
  MX2XL U10859 ( .A(\D_cache/cache[4][131] ), .B(n134), .S0(net112215), .Y(
        \D_cache/n744 ) );
  MX2XL U10860 ( .A(\D_cache/cache[3][131] ), .B(n134), .S0(net112295), .Y(
        \D_cache/n745 ) );
  MX2XL U10861 ( .A(\D_cache/cache[2][131] ), .B(n134), .S0(net112419), .Y(
        \D_cache/n746 ) );
  MX2XL U10862 ( .A(\D_cache/cache[1][131] ), .B(n134), .S0(net112545), .Y(
        \D_cache/n747 ) );
  MX2XL U10863 ( .A(\D_cache/cache[0][131] ), .B(n134), .S0(net112647), .Y(
        \D_cache/n748 ) );
  MX2XL U10864 ( .A(\D_cache/cache[6][129] ), .B(n137), .S0(net112009), .Y(
        \D_cache/n758 ) );
  MX2XL U10865 ( .A(\D_cache/cache[5][129] ), .B(n137), .S0(net112121), .Y(
        \D_cache/n759 ) );
  MX2XL U10866 ( .A(\D_cache/cache[4][129] ), .B(n137), .S0(net112215), .Y(
        \D_cache/n760 ) );
  MX2XL U10867 ( .A(\D_cache/cache[3][129] ), .B(n137), .S0(net112293), .Y(
        \D_cache/n761 ) );
  MX2XL U10868 ( .A(\D_cache/cache[2][129] ), .B(n137), .S0(net112417), .Y(
        \D_cache/n762 ) );
  MX2XL U10869 ( .A(\D_cache/cache[1][129] ), .B(n137), .S0(net112545), .Y(
        \D_cache/n763 ) );
  MX2XL U10870 ( .A(\D_cache/cache[0][129] ), .B(n137), .S0(net112647), .Y(
        \D_cache/n764 ) );
  MX2XL U10871 ( .A(\D_cache/cache[6][150] ), .B(n119), .S0(net111999), .Y(
        \D_cache/n590 ) );
  MX2XL U10872 ( .A(\D_cache/cache[5][150] ), .B(n119), .S0(net112123), .Y(
        \D_cache/n591 ) );
  MX2XL U10873 ( .A(\D_cache/cache[4][150] ), .B(n119), .S0(net112215), .Y(
        \D_cache/n592 ) );
  MX2XL U10874 ( .A(\D_cache/cache[3][150] ), .B(n119), .S0(net112279), .Y(
        \D_cache/n593 ) );
  MX2XL U10875 ( .A(\D_cache/cache[2][150] ), .B(n119), .S0(net112411), .Y(
        \D_cache/n594 ) );
  MX2XL U10876 ( .A(\D_cache/cache[1][150] ), .B(n119), .S0(net112535), .Y(
        \D_cache/n595 ) );
  MX2XL U10877 ( .A(\D_cache/cache[0][150] ), .B(n119), .S0(net112637), .Y(
        \D_cache/n596 ) );
  MX2XL U10878 ( .A(\D_cache/cache[6][141] ), .B(n125), .S0(net111989), .Y(
        \D_cache/n662 ) );
  MX2XL U10879 ( .A(\D_cache/cache[5][141] ), .B(n125), .S0(net112123), .Y(
        \D_cache/n663 ) );
  MX2XL U10880 ( .A(\D_cache/cache[4][141] ), .B(n125), .S0(net112211), .Y(
        \D_cache/n664 ) );
  MX2XL U10881 ( .A(\D_cache/cache[3][141] ), .B(n125), .S0(net112285), .Y(
        \D_cache/n665 ) );
  MX2XL U10882 ( .A(\D_cache/cache[2][141] ), .B(n125), .S0(net112409), .Y(
        \D_cache/n666 ) );
  MX2XL U10883 ( .A(\D_cache/cache[1][141] ), .B(n125), .S0(net112533), .Y(
        \D_cache/n667 ) );
  MX2XL U10884 ( .A(\D_cache/cache[0][141] ), .B(n125), .S0(net112635), .Y(
        \D_cache/n668 ) );
  MX2XL U10885 ( .A(\D_cache/cache[6][134] ), .B(n127), .S0(net111999), .Y(
        \D_cache/n718 ) );
  MX2XL U10886 ( .A(\D_cache/cache[5][134] ), .B(n127), .S0(net112121), .Y(
        \D_cache/n719 ) );
  MX2XL U10887 ( .A(\D_cache/cache[4][134] ), .B(n127), .S0(net112211), .Y(
        \D_cache/n720 ) );
  MX2XL U10888 ( .A(\D_cache/cache[3][134] ), .B(n127), .S0(net112277), .Y(
        \D_cache/n721 ) );
  MX2XL U10889 ( .A(\D_cache/cache[2][134] ), .B(n127), .S0(net112411), .Y(
        \D_cache/n722 ) );
  MX2XL U10890 ( .A(\D_cache/cache[1][134] ), .B(n127), .S0(net112535), .Y(
        \D_cache/n723 ) );
  MX2XL U10891 ( .A(\D_cache/cache[0][134] ), .B(n127), .S0(net112637), .Y(
        \D_cache/n724 ) );
  MX2XL U10892 ( .A(\D_cache/cache[6][149] ), .B(n120), .S0(net111999), .Y(
        \D_cache/n598 ) );
  MX2XL U10893 ( .A(\D_cache/cache[5][149] ), .B(n120), .S0(net112123), .Y(
        \D_cache/n599 ) );
  MX2XL U10894 ( .A(\D_cache/cache[4][149] ), .B(n120), .S0(net112195), .Y(
        \D_cache/n600 ) );
  MX2XL U10895 ( .A(\D_cache/cache[3][149] ), .B(n120), .S0(net112281), .Y(
        \D_cache/n601 ) );
  MX2XL U10896 ( .A(\D_cache/cache[2][149] ), .B(n120), .S0(net112411), .Y(
        \D_cache/n602 ) );
  MX2XL U10897 ( .A(\D_cache/cache[1][149] ), .B(n120), .S0(net112535), .Y(
        \D_cache/n603 ) );
  MX2XL U10898 ( .A(\D_cache/cache[0][149] ), .B(n120), .S0(net112637), .Y(
        \D_cache/n604 ) );
  MX2XL U10899 ( .A(\D_cache/cache[6][132] ), .B(n145), .S0(net111999), .Y(
        \D_cache/n734 ) );
  MX2XL U10900 ( .A(\D_cache/cache[5][132] ), .B(n145), .S0(net112121), .Y(
        \D_cache/n735 ) );
  MX2XL U10901 ( .A(\D_cache/cache[4][132] ), .B(n145), .S0(net112197), .Y(
        \D_cache/n736 ) );
  MX2XL U10902 ( .A(\D_cache/cache[3][132] ), .B(n145), .S0(net112279), .Y(
        \D_cache/n737 ) );
  MX2XL U10903 ( .A(\D_cache/cache[2][132] ), .B(n145), .S0(net112411), .Y(
        \D_cache/n738 ) );
  MX2XL U10904 ( .A(\D_cache/cache[1][132] ), .B(n145), .S0(net112535), .Y(
        \D_cache/n739 ) );
  MX2XL U10905 ( .A(\D_cache/cache[0][132] ), .B(n145), .S0(net112637), .Y(
        \D_cache/n740 ) );
  MX2XL U10906 ( .A(\D_cache/cache[6][151] ), .B(n132), .S0(net111995), .Y(
        \D_cache/n582 ) );
  MX2XL U10907 ( .A(\D_cache/cache[5][151] ), .B(n132), .S0(net112119), .Y(
        \D_cache/n583 ) );
  MX2XL U10908 ( .A(\D_cache/cache[4][151] ), .B(n132), .S0(net112201), .Y(
        \D_cache/n584 ) );
  MX2XL U10909 ( .A(\D_cache/cache[3][151] ), .B(n132), .S0(net112283), .Y(
        \D_cache/n585 ) );
  MX2XL U10910 ( .A(\D_cache/cache[2][151] ), .B(n132), .S0(net112405), .Y(
        \D_cache/n586 ) );
  MX2XL U10911 ( .A(\D_cache/cache[1][151] ), .B(n132), .S0(net112531), .Y(
        \D_cache/n587 ) );
  MX2XL U10912 ( .A(\D_cache/cache[0][151] ), .B(n132), .S0(net112633), .Y(
        \D_cache/n588 ) );
  MX2XL U10913 ( .A(\D_cache/cache[6][137] ), .B(n136), .S0(net111999), .Y(
        \D_cache/n694 ) );
  MX2XL U10914 ( .A(\D_cache/cache[5][137] ), .B(n136), .S0(net112123), .Y(
        \D_cache/n695 ) );
  MX2XL U10915 ( .A(\D_cache/cache[4][137] ), .B(n136), .S0(net112215), .Y(
        \D_cache/n696 ) );
  MX2XL U10916 ( .A(\D_cache/cache[3][137] ), .B(n136), .S0(net112277), .Y(
        \D_cache/n697 ) );
  MX2XL U10917 ( .A(\D_cache/cache[2][137] ), .B(n136), .S0(net112411), .Y(
        \D_cache/n698 ) );
  MX2XL U10918 ( .A(\D_cache/cache[1][137] ), .B(n136), .S0(net112535), .Y(
        \D_cache/n699 ) );
  MX2XL U10919 ( .A(\D_cache/cache[0][137] ), .B(n136), .S0(net112637), .Y(
        \D_cache/n700 ) );
  MX2XL U10920 ( .A(\D_cache/cache[6][135] ), .B(n130), .S0(net111999), .Y(
        \D_cache/n710 ) );
  MX2XL U10921 ( .A(\D_cache/cache[5][135] ), .B(n130), .S0(net112121), .Y(
        \D_cache/n711 ) );
  MX2XL U10922 ( .A(\D_cache/cache[4][135] ), .B(n130), .S0(net112201), .Y(
        \D_cache/n712 ) );
  MX2XL U10923 ( .A(\D_cache/cache[3][135] ), .B(n130), .S0(net112281), .Y(
        \D_cache/n713 ) );
  MX2XL U10924 ( .A(\D_cache/cache[2][135] ), .B(n130), .S0(net112411), .Y(
        \D_cache/n714 ) );
  MX2XL U10925 ( .A(\D_cache/cache[1][135] ), .B(n130), .S0(net112535), .Y(
        \D_cache/n715 ) );
  MX2XL U10926 ( .A(\D_cache/cache[0][135] ), .B(n130), .S0(net112637), .Y(
        \D_cache/n716 ) );
  MX2XL U10927 ( .A(\D_cache/cache[6][128] ), .B(n118), .S0(net111991), .Y(
        \D_cache/n766 ) );
  MX2XL U10928 ( .A(\D_cache/cache[5][128] ), .B(n118), .S0(net112123), .Y(
        \D_cache/n767 ) );
  MX2XL U10929 ( .A(\D_cache/cache[4][128] ), .B(n118), .S0(net112211), .Y(
        \D_cache/n768 ) );
  MX2XL U10930 ( .A(\D_cache/cache[3][128] ), .B(n118), .S0(net112285), .Y(
        \D_cache/n769 ) );
  MX2XL U10931 ( .A(\D_cache/cache[2][128] ), .B(n118), .S0(net112409), .Y(
        \D_cache/n770 ) );
  MX2XL U10932 ( .A(\D_cache/cache[1][128] ), .B(n118), .S0(net112533), .Y(
        \D_cache/n771 ) );
  MX2XL U10933 ( .A(\D_cache/cache[0][128] ), .B(n118), .S0(net112635), .Y(
        \D_cache/n772 ) );
  MX2XL U10934 ( .A(\D_cache/cache[6][148] ), .B(n144), .S0(net111999), .Y(
        \D_cache/n606 ) );
  MX2XL U10935 ( .A(\D_cache/cache[5][148] ), .B(n144), .S0(net112123), .Y(
        \D_cache/n607 ) );
  MX2XL U10936 ( .A(\D_cache/cache[4][148] ), .B(n144), .S0(net112199), .Y(
        \D_cache/n608 ) );
  MX2XL U10937 ( .A(\D_cache/cache[3][148] ), .B(n144), .S0(net112279), .Y(
        \D_cache/n609 ) );
  MX2XL U10938 ( .A(\D_cache/cache[2][148] ), .B(n144), .S0(net112411), .Y(
        \D_cache/n610 ) );
  MX2XL U10939 ( .A(\D_cache/cache[1][148] ), .B(n144), .S0(net112535), .Y(
        \D_cache/n611 ) );
  MX2XL U10940 ( .A(\D_cache/cache[0][148] ), .B(n144), .S0(net112637), .Y(
        \D_cache/n612 ) );
  MX2XL U10941 ( .A(\D_cache/cache[6][136] ), .B(n142), .S0(net111999), .Y(
        \D_cache/n702 ) );
  MX2XL U10942 ( .A(\D_cache/cache[5][136] ), .B(n142), .S0(net112121), .Y(
        \D_cache/n703 ) );
  MX2XL U10943 ( .A(\D_cache/cache[4][136] ), .B(n142), .S0(net112195), .Y(
        \D_cache/n704 ) );
  MX2XL U10944 ( .A(\D_cache/cache[3][136] ), .B(n142), .S0(net112285), .Y(
        \D_cache/n705 ) );
  MX2XL U10945 ( .A(\D_cache/cache[2][136] ), .B(n142), .S0(net112409), .Y(
        \D_cache/n706 ) );
  MX2XL U10946 ( .A(\D_cache/cache[1][136] ), .B(n142), .S0(net112533), .Y(
        \D_cache/n707 ) );
  MX2XL U10947 ( .A(\D_cache/cache[0][136] ), .B(n142), .S0(net112635), .Y(
        \D_cache/n708 ) );
  MX2XL U10948 ( .A(\i_MIPS/Reg_W[0] ), .B(n10133), .S0(n5509), .Y(
        \i_MIPS/n477 ) );
  MX2XL U10949 ( .A(\D_cache/cache[7][144] ), .B(n128), .S0(net111873), .Y(
        \D_cache/n637 ) );
  MX2XL U10950 ( .A(\D_cache/cache[6][144] ), .B(n128), .S0(net112009), .Y(
        \D_cache/n638 ) );
  MX2XL U10951 ( .A(\D_cache/cache[5][144] ), .B(n128), .S0(net112123), .Y(
        \D_cache/n639 ) );
  MX2XL U10952 ( .A(\D_cache/cache[4][144] ), .B(n128), .S0(net112199), .Y(
        \D_cache/n640 ) );
  MX2XL U10953 ( .A(\D_cache/cache[3][144] ), .B(n128), .S0(net112285), .Y(
        \D_cache/n641 ) );
  MX2XL U10954 ( .A(\D_cache/cache[2][144] ), .B(n128), .S0(net112409), .Y(
        \D_cache/n642 ) );
  MX2XL U10955 ( .A(\D_cache/cache[1][144] ), .B(n128), .S0(net112533), .Y(
        \D_cache/n643 ) );
  MX2XL U10956 ( .A(\D_cache/cache[0][144] ), .B(n128), .S0(net112635), .Y(
        \D_cache/n644 ) );
  MX2XL U10957 ( .A(\D_cache/cache[7][139] ), .B(n124), .S0(net111873), .Y(
        \D_cache/n677 ) );
  MX2XL U10958 ( .A(\D_cache/cache[6][139] ), .B(n124), .S0(net111993), .Y(
        \D_cache/n678 ) );
  MX2XL U10959 ( .A(\D_cache/cache[5][139] ), .B(n124), .S0(net112121), .Y(
        \D_cache/n679 ) );
  MX2XL U10960 ( .A(\D_cache/cache[4][139] ), .B(n124), .S0(net112201), .Y(
        \D_cache/n680 ) );
  MX2XL U10961 ( .A(\D_cache/cache[3][139] ), .B(n124), .S0(net112285), .Y(
        \D_cache/n681 ) );
  MX2XL U10962 ( .A(\D_cache/cache[2][139] ), .B(n124), .S0(net112409), .Y(
        \D_cache/n682 ) );
  MX2XL U10963 ( .A(\D_cache/cache[1][139] ), .B(n124), .S0(net112533), .Y(
        \D_cache/n683 ) );
  MX2XL U10964 ( .A(\D_cache/cache[0][139] ), .B(n124), .S0(net112635), .Y(
        \D_cache/n684 ) );
  MX2XL U10965 ( .A(\D_cache/cache[7][140] ), .B(n10622), .S0(net111873), .Y(
        \D_cache/n669 ) );
  MX2XL U10966 ( .A(\D_cache/cache[5][140] ), .B(n10622), .S0(net112123), .Y(
        \D_cache/n671 ) );
  MX2XL U10967 ( .A(\D_cache/cache[6][146] ), .B(n10669), .S0(net111999), .Y(
        \D_cache/n622 ) );
  MX2XL U10968 ( .A(\D_cache/cache[5][146] ), .B(n10669), .S0(net112121), .Y(
        \D_cache/n623 ) );
  MX2XL U10969 ( .A(\D_cache/cache[6][138] ), .B(n129), .S0(net111999), .Y(
        \D_cache/n686 ) );
  MX2XL U10970 ( .A(\D_cache/cache[5][138] ), .B(n129), .S0(net112123), .Y(
        \D_cache/n687 ) );
  MX2XL U10971 ( .A(\D_cache/cache[4][138] ), .B(n129), .S0(net112211), .Y(
        \D_cache/n688 ) );
  MX2XL U10972 ( .A(\D_cache/cache[3][138] ), .B(n129), .S0(net112293), .Y(
        \D_cache/n689 ) );
  MX2XL U10973 ( .A(\D_cache/cache[2][138] ), .B(n129), .S0(net112411), .Y(
        \D_cache/n690 ) );
  MX2XL U10974 ( .A(\D_cache/cache[1][138] ), .B(n129), .S0(net112535), .Y(
        \D_cache/n691 ) );
  MX2XL U10975 ( .A(\D_cache/cache[0][138] ), .B(n129), .S0(net112637), .Y(
        \D_cache/n692 ) );
  MX2XL U10976 ( .A(\D_cache/cache[6][133] ), .B(n123), .S0(net111999), .Y(
        \D_cache/n726 ) );
  MX2XL U10977 ( .A(\D_cache/cache[5][133] ), .B(n123), .S0(net112121), .Y(
        \D_cache/n727 ) );
  MX2XL U10978 ( .A(\D_cache/cache[4][133] ), .B(n123), .S0(net112195), .Y(
        \D_cache/n728 ) );
  MX2XL U10979 ( .A(\D_cache/cache[3][133] ), .B(n123), .S0(net112295), .Y(
        \D_cache/n729 ) );
  MX2XL U10980 ( .A(\D_cache/cache[2][133] ), .B(n123), .S0(net112411), .Y(
        \D_cache/n730 ) );
  MX2XL U10981 ( .A(\D_cache/cache[1][133] ), .B(n123), .S0(net112535), .Y(
        \D_cache/n731 ) );
  MX2XL U10982 ( .A(\D_cache/cache[0][133] ), .B(n123), .S0(net112637), .Y(
        \D_cache/n732 ) );
  CLKMX2X2 U10983 ( .A(\I_cache/cache[7][99] ), .B(n9517), .S0(n5372), .Y(
        n12024) );
  CLKMX2X2 U10984 ( .A(\I_cache/cache[6][99] ), .B(n9517), .S0(n5416), .Y(
        n12025) );
  CLKMX2X2 U10985 ( .A(\I_cache/cache[5][99] ), .B(n9517), .S0(n5285), .Y(
        n12026) );
  CLKMX2X2 U10986 ( .A(\I_cache/cache[4][99] ), .B(n9517), .S0(n5325), .Y(
        n12027) );
  CLKMX2X2 U10987 ( .A(\I_cache/cache[3][99] ), .B(n9517), .S0(n5193), .Y(
        n12028) );
  CLKMX2X2 U10988 ( .A(\I_cache/cache[2][99] ), .B(n9517), .S0(n5242), .Y(
        n12029) );
  CLKMX2X2 U10989 ( .A(\I_cache/cache[1][99] ), .B(n9517), .S0(n5111), .Y(
        n12030) );
  CLKMX2X2 U10990 ( .A(\I_cache/cache[0][99] ), .B(n9517), .S0(n5148), .Y(
        n12031) );
  MX2XL U10991 ( .A(\i_MIPS/ID_EX[56] ), .B(n4029), .S0(n5507), .Y(
        \i_MIPS/n407 ) );
  MX2XL U10992 ( .A(\D_cache/cache[6][142] ), .B(n10682), .S0(net112009), .Y(
        \D_cache/n654 ) );
  MX2XL U10993 ( .A(\D_cache/cache[5][142] ), .B(n10682), .S0(net112123), .Y(
        \D_cache/n655 ) );
  MX2XL U10994 ( .A(\D_cache/cache[4][142] ), .B(n10682), .S0(net112215), .Y(
        \D_cache/n656 ) );
  MX2XL U10995 ( .A(\D_cache/cache[3][142] ), .B(n10682), .S0(net112277), .Y(
        \D_cache/n657 ) );
  MX2XL U10996 ( .A(\D_cache/cache[2][142] ), .B(n10682), .S0(net112415), .Y(
        \D_cache/n658 ) );
  MX2XL U10997 ( .A(\D_cache/cache[1][142] ), .B(n10682), .S0(net112545), .Y(
        \D_cache/n659 ) );
  MX2XL U10998 ( .A(\D_cache/cache[0][142] ), .B(n10682), .S0(net112647), .Y(
        \D_cache/n660 ) );
  MX2XL U10999 ( .A(\I_cache/cache[4][138] ), .B(n10989), .S0(n5320), .Y(
        n11715) );
  MX2XL U11000 ( .A(\I_cache/cache[4][129] ), .B(n10995), .S0(n5321), .Y(
        n11787) );
  CLKMX2X2 U11001 ( .A(\I_cache/cache[7][127] ), .B(n11037), .S0(n5367), .Y(
        n11800) );
  CLKMX2X2 U11002 ( .A(\I_cache/cache[6][127] ), .B(n11037), .S0(n5411), .Y(
        n11801) );
  CLKMX2X2 U11003 ( .A(\I_cache/cache[5][127] ), .B(n11037), .S0(n5278), .Y(
        n11802) );
  CLKMX2X2 U11004 ( .A(\I_cache/cache[4][127] ), .B(n11037), .S0(n5320), .Y(
        n11803) );
  CLKMX2X2 U11005 ( .A(\I_cache/cache[3][127] ), .B(n11037), .S0(n5191), .Y(
        n11804) );
  CLKMX2X2 U11006 ( .A(\I_cache/cache[2][127] ), .B(n11037), .S0(n5233), .Y(
        n11805) );
  CLKMX2X2 U11007 ( .A(\I_cache/cache[1][127] ), .B(n11037), .S0(n5104), .Y(
        n11806) );
  CLKMX2X2 U11008 ( .A(\I_cache/cache[0][127] ), .B(n11037), .S0(n5146), .Y(
        n11807) );
  CLKMX2X2 U11009 ( .A(\I_cache/cache[7][126] ), .B(n9798), .S0(n5370), .Y(
        n11808) );
  CLKMX2X2 U11010 ( .A(\I_cache/cache[6][126] ), .B(n9798), .S0(n5414), .Y(
        n11809) );
  CLKMX2X2 U11011 ( .A(\I_cache/cache[5][126] ), .B(n9798), .S0(n5280), .Y(
        n11810) );
  CLKMX2X2 U11012 ( .A(\I_cache/cache[4][126] ), .B(n9798), .S0(n5323), .Y(
        n11811) );
  CLKMX2X2 U11013 ( .A(\I_cache/cache[3][126] ), .B(n9798), .S0(n5194), .Y(
        n11812) );
  CLKMX2X2 U11014 ( .A(\I_cache/cache[2][126] ), .B(n9798), .S0(n5236), .Y(
        n11813) );
  CLKMX2X2 U11015 ( .A(\I_cache/cache[1][126] ), .B(n9798), .S0(n5107), .Y(
        n11814) );
  CLKMX2X2 U11016 ( .A(\I_cache/cache[0][126] ), .B(n9798), .S0(n5149), .Y(
        n11815) );
  CLKMX2X2 U11017 ( .A(\I_cache/cache[7][125] ), .B(n11160), .S0(n5367), .Y(
        n11816) );
  CLKMX2X2 U11018 ( .A(\I_cache/cache[6][125] ), .B(n11160), .S0(n5411), .Y(
        n11817) );
  CLKMX2X2 U11019 ( .A(\I_cache/cache[5][125] ), .B(n11160), .S0(n5278), .Y(
        n11818) );
  CLKMX2X2 U11020 ( .A(\I_cache/cache[4][125] ), .B(n11160), .S0(n5320), .Y(
        n11819) );
  CLKMX2X2 U11021 ( .A(\I_cache/cache[3][125] ), .B(n11160), .S0(n5191), .Y(
        n11820) );
  CLKMX2X2 U11022 ( .A(\I_cache/cache[2][125] ), .B(n11160), .S0(n5233), .Y(
        n11821) );
  CLKMX2X2 U11023 ( .A(\I_cache/cache[1][125] ), .B(n11160), .S0(n5104), .Y(
        n11822) );
  CLKMX2X2 U11024 ( .A(\I_cache/cache[0][125] ), .B(n11160), .S0(n5146), .Y(
        n11823) );
  CLKMX2X2 U11025 ( .A(\I_cache/cache[7][124] ), .B(n9774), .S0(n5370), .Y(
        n11824) );
  CLKMX2X2 U11026 ( .A(\I_cache/cache[6][124] ), .B(n9774), .S0(n5414), .Y(
        n11825) );
  CLKMX2X2 U11027 ( .A(\I_cache/cache[5][124] ), .B(n9774), .S0(n5280), .Y(
        n11826) );
  CLKMX2X2 U11028 ( .A(\I_cache/cache[4][124] ), .B(n9774), .S0(n5323), .Y(
        n11827) );
  CLKMX2X2 U11029 ( .A(\I_cache/cache[3][124] ), .B(n9774), .S0(n5194), .Y(
        n11828) );
  CLKMX2X2 U11030 ( .A(\I_cache/cache[2][124] ), .B(n9774), .S0(n5236), .Y(
        n11829) );
  CLKMX2X2 U11031 ( .A(\I_cache/cache[1][124] ), .B(n9774), .S0(n5107), .Y(
        n11830) );
  CLKMX2X2 U11032 ( .A(\I_cache/cache[0][124] ), .B(n9774), .S0(n5149), .Y(
        n11831) );
  CLKMX2X2 U11033 ( .A(\I_cache/cache[7][123] ), .B(n9730), .S0(n5370), .Y(
        n11832) );
  CLKMX2X2 U11034 ( .A(\I_cache/cache[6][123] ), .B(n9730), .S0(n5414), .Y(
        n11833) );
  CLKMX2X2 U11035 ( .A(\I_cache/cache[5][123] ), .B(n9730), .S0(n5280), .Y(
        n11834) );
  CLKMX2X2 U11036 ( .A(\I_cache/cache[4][123] ), .B(n9730), .S0(n5323), .Y(
        n11835) );
  CLKMX2X2 U11037 ( .A(\I_cache/cache[3][123] ), .B(n9730), .S0(n5194), .Y(
        n11836) );
  CLKMX2X2 U11038 ( .A(\I_cache/cache[2][123] ), .B(n9730), .S0(n5236), .Y(
        n11837) );
  CLKMX2X2 U11039 ( .A(\I_cache/cache[1][123] ), .B(n9730), .S0(n5107), .Y(
        n11838) );
  CLKMX2X2 U11040 ( .A(\I_cache/cache[0][123] ), .B(n9730), .S0(n5149), .Y(
        n11839) );
  CLKMX2X2 U11041 ( .A(\I_cache/cache[7][122] ), .B(n9706), .S0(n5374), .Y(
        n11840) );
  CLKMX2X2 U11042 ( .A(\I_cache/cache[6][122] ), .B(n9706), .S0(n5419), .Y(
        n11841) );
  CLKMX2X2 U11043 ( .A(\I_cache/cache[5][122] ), .B(n9706), .S0(n5283), .Y(
        n11842) );
  CLKMX2X2 U11044 ( .A(\I_cache/cache[4][122] ), .B(n9706), .S0(n5327), .Y(
        n11843) );
  CLKMX2X2 U11045 ( .A(\I_cache/cache[3][122] ), .B(n9706), .S0(n5199), .Y(
        n11844) );
  CLKMX2X2 U11046 ( .A(\I_cache/cache[2][122] ), .B(n9706), .S0(n5241), .Y(
        n11845) );
  CLKMX2X2 U11047 ( .A(\I_cache/cache[1][122] ), .B(n9706), .S0(n5110), .Y(
        n11846) );
  CLKMX2X2 U11048 ( .A(\I_cache/cache[0][122] ), .B(n9706), .S0(n5154), .Y(
        n11847) );
  CLKMX2X2 U11049 ( .A(\I_cache/cache[6][121] ), .B(n10119), .S0(n5410), .Y(
        n11849) );
  CLKMX2X2 U11050 ( .A(\I_cache/cache[4][121] ), .B(n10119), .S0(n4679), .Y(
        n11851) );
  CLKMX2X2 U11051 ( .A(\I_cache/cache[3][121] ), .B(n10119), .S0(n5190), .Y(
        n11852) );
  CLKMX2X2 U11052 ( .A(\I_cache/cache[2][121] ), .B(n10119), .S0(n5235), .Y(
        n11853) );
  CLKMX2X2 U11053 ( .A(\I_cache/cache[1][121] ), .B(n10119), .S0(n5103), .Y(
        n11854) );
  CLKMX2X2 U11054 ( .A(\I_cache/cache[0][121] ), .B(n10119), .S0(n5145), .Y(
        n11855) );
  CLKMX2X2 U11055 ( .A(\I_cache/cache[7][120] ), .B(n9897), .S0(n5371), .Y(
        n11856) );
  CLKMX2X2 U11056 ( .A(\I_cache/cache[6][120] ), .B(n9897), .S0(n5415), .Y(
        n11857) );
  CLKMX2X2 U11057 ( .A(\I_cache/cache[5][120] ), .B(n9897), .S0(n5281), .Y(
        n11858) );
  CLKMX2X2 U11058 ( .A(\I_cache/cache[4][120] ), .B(n9897), .S0(n5324), .Y(
        n11859) );
  CLKMX2X2 U11059 ( .A(\I_cache/cache[3][120] ), .B(n9897), .S0(n5195), .Y(
        n11860) );
  CLKMX2X2 U11060 ( .A(\I_cache/cache[2][120] ), .B(n9897), .S0(n5237), .Y(
        n11861) );
  CLKMX2X2 U11061 ( .A(\I_cache/cache[1][120] ), .B(n9897), .S0(n5108), .Y(
        n11862) );
  CLKMX2X2 U11062 ( .A(\I_cache/cache[0][120] ), .B(n9897), .S0(n5150), .Y(
        n11863) );
  CLKMX2X2 U11063 ( .A(\I_cache/cache[7][119] ), .B(n9921), .S0(n5372), .Y(
        n11864) );
  CLKMX2X2 U11064 ( .A(\I_cache/cache[6][119] ), .B(n9921), .S0(n5416), .Y(
        n11865) );
  CLKMX2X2 U11065 ( .A(\I_cache/cache[5][119] ), .B(n9921), .S0(n5282), .Y(
        n11866) );
  CLKMX2X2 U11066 ( .A(\I_cache/cache[4][119] ), .B(n9921), .S0(n5325), .Y(
        n11867) );
  CLKMX2X2 U11067 ( .A(\I_cache/cache[3][119] ), .B(n9921), .S0(n5196), .Y(
        n11868) );
  CLKMX2X2 U11068 ( .A(\I_cache/cache[2][119] ), .B(n9921), .S0(n5238), .Y(
        n11869) );
  CLKMX2X2 U11069 ( .A(\I_cache/cache[1][119] ), .B(n9921), .S0(n5109), .Y(
        n11870) );
  CLKMX2X2 U11070 ( .A(\I_cache/cache[0][119] ), .B(n9921), .S0(n5151), .Y(
        n11871) );
  CLKMX2X2 U11071 ( .A(\I_cache/cache[7][118] ), .B(n9853), .S0(n5369), .Y(
        n11872) );
  CLKMX2X2 U11072 ( .A(\I_cache/cache[6][118] ), .B(n9853), .S0(n5413), .Y(
        n11873) );
  CLKMX2X2 U11073 ( .A(\I_cache/cache[5][118] ), .B(n9853), .S0(n5279), .Y(
        n11874) );
  CLKMX2X2 U11074 ( .A(\I_cache/cache[4][118] ), .B(n9853), .S0(n5322), .Y(
        n11875) );
  CLKMX2X2 U11075 ( .A(\I_cache/cache[3][118] ), .B(n9853), .S0(n5193), .Y(
        n11876) );
  CLKMX2X2 U11076 ( .A(\I_cache/cache[2][118] ), .B(n9853), .S0(n5235), .Y(
        n11877) );
  CLKMX2X2 U11077 ( .A(\I_cache/cache[1][118] ), .B(n9853), .S0(n5106), .Y(
        n11878) );
  CLKMX2X2 U11078 ( .A(\I_cache/cache[0][118] ), .B(n9853), .S0(n5148), .Y(
        n11879) );
  CLKMX2X2 U11079 ( .A(\I_cache/cache[7][117] ), .B(n9873), .S0(n5369), .Y(
        n11880) );
  CLKMX2X2 U11080 ( .A(\I_cache/cache[6][117] ), .B(n9873), .S0(n5413), .Y(
        n11881) );
  CLKMX2X2 U11081 ( .A(\I_cache/cache[5][117] ), .B(n9873), .S0(n5279), .Y(
        n11882) );
  CLKMX2X2 U11082 ( .A(\I_cache/cache[4][117] ), .B(n9873), .S0(n5322), .Y(
        n11883) );
  CLKMX2X2 U11083 ( .A(\I_cache/cache[3][117] ), .B(n9873), .S0(n5193), .Y(
        n11884) );
  CLKMX2X2 U11084 ( .A(\I_cache/cache[2][117] ), .B(n9873), .S0(n5235), .Y(
        n11885) );
  CLKMX2X2 U11085 ( .A(\I_cache/cache[1][117] ), .B(n9873), .S0(n5106), .Y(
        n11886) );
  CLKMX2X2 U11086 ( .A(\I_cache/cache[0][117] ), .B(n9873), .S0(n5148), .Y(
        n11887) );
  CLKMX2X2 U11087 ( .A(\I_cache/cache[7][116] ), .B(n10017), .S0(n5371), .Y(
        n11888) );
  CLKMX2X2 U11088 ( .A(\I_cache/cache[6][116] ), .B(n10017), .S0(n5415), .Y(
        n11889) );
  CLKMX2X2 U11089 ( .A(\I_cache/cache[5][116] ), .B(n10017), .S0(n5281), .Y(
        n11890) );
  CLKMX2X2 U11090 ( .A(\I_cache/cache[4][116] ), .B(n10017), .S0(n5324), .Y(
        n11891) );
  CLKMX2X2 U11091 ( .A(\I_cache/cache[3][116] ), .B(n10017), .S0(n5195), .Y(
        n11892) );
  CLKMX2X2 U11092 ( .A(\I_cache/cache[2][116] ), .B(n10017), .S0(n5237), .Y(
        n11893) );
  CLKMX2X2 U11093 ( .A(\I_cache/cache[1][116] ), .B(n10017), .S0(n5108), .Y(
        n11894) );
  CLKMX2X2 U11094 ( .A(\I_cache/cache[0][116] ), .B(n10017), .S0(n5150), .Y(
        n11895) );
  CLKMX2X2 U11095 ( .A(\I_cache/cache[7][115] ), .B(n9988), .S0(n5372), .Y(
        n11896) );
  CLKMX2X2 U11096 ( .A(\I_cache/cache[6][115] ), .B(n9988), .S0(n5416), .Y(
        n11897) );
  CLKMX2X2 U11097 ( .A(\I_cache/cache[5][115] ), .B(n9988), .S0(n5282), .Y(
        n11898) );
  CLKMX2X2 U11098 ( .A(\I_cache/cache[4][115] ), .B(n9988), .S0(n5325), .Y(
        n11899) );
  CLKMX2X2 U11099 ( .A(\I_cache/cache[3][115] ), .B(n9988), .S0(n5196), .Y(
        n11900) );
  CLKMX2X2 U11100 ( .A(\I_cache/cache[2][115] ), .B(n9988), .S0(n5238), .Y(
        n11901) );
  CLKMX2X2 U11101 ( .A(\I_cache/cache[1][115] ), .B(n9988), .S0(n5109), .Y(
        n11902) );
  CLKMX2X2 U11102 ( .A(\I_cache/cache[0][115] ), .B(n9988), .S0(n5151), .Y(
        n11903) );
  CLKMX2X2 U11103 ( .A(\I_cache/cache[7][114] ), .B(n10041), .S0(n5371), .Y(
        n11904) );
  CLKMX2X2 U11104 ( .A(\I_cache/cache[6][114] ), .B(n10041), .S0(n5415), .Y(
        n11905) );
  CLKMX2X2 U11105 ( .A(\I_cache/cache[5][114] ), .B(n10041), .S0(n5281), .Y(
        n11906) );
  CLKMX2X2 U11106 ( .A(\I_cache/cache[2][114] ), .B(n10041), .S0(n5237), .Y(
        n11909) );
  CLKMX2X2 U11107 ( .A(\I_cache/cache[1][114] ), .B(n10041), .S0(n5108), .Y(
        n11910) );
  CLKMX2X2 U11108 ( .A(\I_cache/cache[0][114] ), .B(n10041), .S0(n5150), .Y(
        n11911) );
  CLKMX2X2 U11109 ( .A(\I_cache/cache[7][113] ), .B(n11134), .S0(n5367), .Y(
        n11912) );
  CLKMX2X2 U11110 ( .A(\I_cache/cache[6][113] ), .B(n11134), .S0(n5411), .Y(
        n11913) );
  CLKMX2X2 U11111 ( .A(\I_cache/cache[5][113] ), .B(n11134), .S0(n5278), .Y(
        n11914) );
  CLKMX2X2 U11112 ( .A(\I_cache/cache[4][113] ), .B(n11134), .S0(n5320), .Y(
        n11915) );
  CLKMX2X2 U11113 ( .A(\I_cache/cache[3][113] ), .B(n11134), .S0(n5191), .Y(
        n11916) );
  CLKMX2X2 U11114 ( .A(\I_cache/cache[2][113] ), .B(n11134), .S0(n5233), .Y(
        n11917) );
  CLKMX2X2 U11115 ( .A(\I_cache/cache[1][113] ), .B(n11134), .S0(n5104), .Y(
        n11918) );
  CLKMX2X2 U11116 ( .A(\I_cache/cache[0][113] ), .B(n11134), .S0(n5146), .Y(
        n11919) );
  CLKMX2X2 U11117 ( .A(\I_cache/cache[6][112] ), .B(n10070), .S0(n5415), .Y(
        n11921) );
  CLKMX2X2 U11118 ( .A(\I_cache/cache[5][112] ), .B(n10070), .S0(n5281), .Y(
        n11922) );
  CLKMX2X2 U11119 ( .A(\I_cache/cache[4][112] ), .B(n10070), .S0(n5324), .Y(
        n11923) );
  CLKMX2X2 U11120 ( .A(\I_cache/cache[3][112] ), .B(n10070), .S0(n5195), .Y(
        n11924) );
  CLKMX2X2 U11121 ( .A(\I_cache/cache[2][112] ), .B(n10070), .S0(n5237), .Y(
        n11925) );
  CLKMX2X2 U11122 ( .A(\I_cache/cache[0][112] ), .B(n10070), .S0(n5150), .Y(
        n11927) );
  CLKMX2X2 U11123 ( .A(\I_cache/cache[7][110] ), .B(n9402), .S0(n5367), .Y(
        n11936) );
  CLKMX2X2 U11124 ( .A(\I_cache/cache[6][110] ), .B(n9402), .S0(n5418), .Y(
        n11937) );
  CLKMX2X2 U11125 ( .A(\I_cache/cache[5][110] ), .B(n9402), .S0(n5284), .Y(
        n11938) );
  CLKMX2X2 U11126 ( .A(\I_cache/cache[4][110] ), .B(n9402), .S0(n5326), .Y(
        n11939) );
  CLKMX2X2 U11127 ( .A(\I_cache/cache[3][110] ), .B(n9402), .S0(n5198), .Y(
        n11940) );
  CLKMX2X2 U11128 ( .A(\I_cache/cache[2][110] ), .B(n9402), .S0(n5240), .Y(
        n11941) );
  CLKMX2X2 U11129 ( .A(\I_cache/cache[1][110] ), .B(n9402), .S0(n5111), .Y(
        n11942) );
  CLKMX2X2 U11130 ( .A(\I_cache/cache[0][110] ), .B(n9402), .S0(n5153), .Y(
        n11943) );
  CLKMX2X2 U11131 ( .A(\I_cache/cache[7][109] ), .B(n9382), .S0(n5370), .Y(
        n11944) );
  CLKMX2X2 U11132 ( .A(\I_cache/cache[6][109] ), .B(n9382), .S0(n5418), .Y(
        n11945) );
  CLKMX2X2 U11133 ( .A(\I_cache/cache[5][109] ), .B(n9382), .S0(n5284), .Y(
        n11946) );
  CLKMX2X2 U11134 ( .A(\I_cache/cache[4][109] ), .B(n9382), .S0(n5322), .Y(
        n11947) );
  CLKMX2X2 U11135 ( .A(\I_cache/cache[3][109] ), .B(n9382), .S0(n5198), .Y(
        n11948) );
  CLKMX2X2 U11136 ( .A(\I_cache/cache[2][109] ), .B(n9382), .S0(n5240), .Y(
        n11949) );
  CLKMX2X2 U11137 ( .A(\I_cache/cache[1][109] ), .B(n9382), .S0(n5107), .Y(
        n11950) );
  CLKMX2X2 U11138 ( .A(\I_cache/cache[0][109] ), .B(n9382), .S0(n5153), .Y(
        n11951) );
  CLKMX2X2 U11139 ( .A(\I_cache/cache[6][108] ), .B(n10095), .S0(n5410), .Y(
        n11953) );
  CLKMX2X2 U11140 ( .A(\I_cache/cache[4][108] ), .B(n10095), .S0(n4698), .Y(
        n11955) );
  CLKMX2X2 U11141 ( .A(\I_cache/cache[3][108] ), .B(n10095), .S0(n5190), .Y(
        n11956) );
  CLKMX2X2 U11142 ( .A(\I_cache/cache[2][108] ), .B(n10095), .S0(n5235), .Y(
        n11957) );
  CLKMX2X2 U11143 ( .A(\I_cache/cache[1][108] ), .B(n10095), .S0(n5103), .Y(
        n11958) );
  CLKMX2X2 U11144 ( .A(\I_cache/cache[0][108] ), .B(n10095), .S0(n5145), .Y(
        n11959) );
  CLKMX2X2 U11145 ( .A(\I_cache/cache[7][107] ), .B(n9964), .S0(n5372), .Y(
        n11960) );
  CLKMX2X2 U11146 ( .A(\I_cache/cache[6][107] ), .B(n9964), .S0(n5416), .Y(
        n11961) );
  CLKMX2X2 U11147 ( .A(\I_cache/cache[5][107] ), .B(n9964), .S0(n5282), .Y(
        n11962) );
  CLKMX2X2 U11148 ( .A(\I_cache/cache[4][107] ), .B(n9964), .S0(n5325), .Y(
        n11963) );
  CLKMX2X2 U11149 ( .A(\I_cache/cache[3][107] ), .B(n9964), .S0(n5196), .Y(
        n11964) );
  CLKMX2X2 U11150 ( .A(\I_cache/cache[2][107] ), .B(n9964), .S0(n5238), .Y(
        n11965) );
  CLKMX2X2 U11151 ( .A(\I_cache/cache[1][107] ), .B(n9964), .S0(n5109), .Y(
        n11966) );
  CLKMX2X2 U11152 ( .A(\I_cache/cache[0][107] ), .B(n9964), .S0(n5151), .Y(
        n11967) );
  CLKMX2X2 U11153 ( .A(\I_cache/cache[7][106] ), .B(n9669), .S0(n5374), .Y(
        n11968) );
  CLKMX2X2 U11154 ( .A(\I_cache/cache[6][106] ), .B(n9669), .S0(n5419), .Y(
        n11969) );
  CLKMX2X2 U11155 ( .A(\I_cache/cache[5][106] ), .B(n9669), .S0(n5281), .Y(
        n11970) );
  CLKMX2X2 U11156 ( .A(\I_cache/cache[4][106] ), .B(n9669), .S0(n5327), .Y(
        n11971) );
  CLKMX2X2 U11157 ( .A(\I_cache/cache[3][106] ), .B(n9669), .S0(n5199), .Y(
        n11972) );
  CLKMX2X2 U11158 ( .A(\I_cache/cache[2][106] ), .B(n9669), .S0(n5241), .Y(
        n11973) );
  CLKMX2X2 U11159 ( .A(\I_cache/cache[1][106] ), .B(n9669), .S0(n5110), .Y(
        n11974) );
  CLKMX2X2 U11160 ( .A(\I_cache/cache[0][106] ), .B(n9669), .S0(n5154), .Y(
        n11975) );
  CLKMX2X2 U11161 ( .A(\I_cache/cache[7][105] ), .B(n9650), .S0(n5374), .Y(
        n11976) );
  CLKMX2X2 U11162 ( .A(\I_cache/cache[6][105] ), .B(n9650), .S0(n5419), .Y(
        n11977) );
  CLKMX2X2 U11163 ( .A(\I_cache/cache[4][105] ), .B(n9650), .S0(n5327), .Y(
        n11979) );
  CLKMX2X2 U11164 ( .A(\I_cache/cache[3][105] ), .B(n9650), .S0(n5199), .Y(
        n11980) );
  CLKMX2X2 U11165 ( .A(\I_cache/cache[2][105] ), .B(n9650), .S0(n5241), .Y(
        n11981) );
  CLKMX2X2 U11166 ( .A(\I_cache/cache[1][105] ), .B(n9650), .S0(n5110), .Y(
        n11982) );
  CLKMX2X2 U11167 ( .A(\I_cache/cache[0][105] ), .B(n9650), .S0(n5154), .Y(
        n11983) );
  CLKMX2X2 U11168 ( .A(\I_cache/cache[7][104] ), .B(n9426), .S0(n5373), .Y(
        n11984) );
  CLKMX2X2 U11169 ( .A(\I_cache/cache[6][104] ), .B(n9426), .S0(n5417), .Y(
        n11985) );
  CLKMX2X2 U11170 ( .A(\I_cache/cache[5][104] ), .B(n9426), .S0(n5283), .Y(
        n11986) );
  CLKMX2X2 U11171 ( .A(\I_cache/cache[3][104] ), .B(n9426), .S0(n5197), .Y(
        n11988) );
  CLKMX2X2 U11172 ( .A(\I_cache/cache[2][104] ), .B(n9426), .S0(n5239), .Y(
        n11989) );
  CLKMX2X2 U11173 ( .A(\I_cache/cache[1][104] ), .B(n9426), .S0(n5111), .Y(
        n11990) );
  CLKMX2X2 U11174 ( .A(\I_cache/cache[0][104] ), .B(n9426), .S0(n5152), .Y(
        n11991) );
  CLKMX2X2 U11175 ( .A(\I_cache/cache[7][103] ), .B(n9830), .S0(n5369), .Y(
        n11992) );
  CLKMX2X2 U11176 ( .A(\I_cache/cache[6][103] ), .B(n9830), .S0(n5413), .Y(
        n11993) );
  CLKMX2X2 U11177 ( .A(\I_cache/cache[5][103] ), .B(n9830), .S0(n5279), .Y(
        n11994) );
  CLKMX2X2 U11178 ( .A(\I_cache/cache[4][103] ), .B(n9830), .S0(n5322), .Y(
        n11995) );
  CLKMX2X2 U11179 ( .A(\I_cache/cache[3][103] ), .B(n9830), .S0(n5193), .Y(
        n11996) );
  CLKMX2X2 U11180 ( .A(\I_cache/cache[2][103] ), .B(n9830), .S0(n5235), .Y(
        n11997) );
  CLKMX2X2 U11181 ( .A(\I_cache/cache[1][103] ), .B(n9830), .S0(n5106), .Y(
        n11998) );
  CLKMX2X2 U11182 ( .A(\I_cache/cache[0][103] ), .B(n9830), .S0(n5148), .Y(
        n11999) );
  CLKMX2X2 U11183 ( .A(\I_cache/cache[7][102] ), .B(n9441), .S0(n5373), .Y(
        n12000) );
  CLKMX2X2 U11184 ( .A(\I_cache/cache[6][102] ), .B(n9441), .S0(n5417), .Y(
        n12001) );
  CLKMX2X2 U11185 ( .A(\I_cache/cache[5][102] ), .B(n9441), .S0(n5283), .Y(
        n12002) );
  CLKMX2X2 U11186 ( .A(\I_cache/cache[4][102] ), .B(n9441), .S0(n5326), .Y(
        n12003) );
  CLKMX2X2 U11187 ( .A(\I_cache/cache[3][102] ), .B(n9441), .S0(n5197), .Y(
        n12004) );
  CLKMX2X2 U11188 ( .A(\I_cache/cache[2][102] ), .B(n9441), .S0(n5239), .Y(
        n12005) );
  CLKMX2X2 U11189 ( .A(\I_cache/cache[1][102] ), .B(n9441), .S0(n5102), .Y(
        n12006) );
  CLKMX2X2 U11190 ( .A(\I_cache/cache[0][102] ), .B(n9441), .S0(n5152), .Y(
        n12007) );
  CLKMX2X2 U11191 ( .A(\I_cache/cache[7][101] ), .B(n9546), .S0(n5371), .Y(
        n12008) );
  CLKMX2X2 U11192 ( .A(\I_cache/cache[6][101] ), .B(n9546), .S0(n5419), .Y(
        n12009) );
  CLKMX2X2 U11193 ( .A(\I_cache/cache[5][101] ), .B(n9546), .S0(n4675), .Y(
        n12010) );
  CLKMX2X2 U11194 ( .A(\I_cache/cache[4][101] ), .B(n9546), .S0(n5327), .Y(
        n12011) );
  CLKMX2X2 U11195 ( .A(\I_cache/cache[3][101] ), .B(n9546), .S0(n5199), .Y(
        n12012) );
  CLKMX2X2 U11196 ( .A(\I_cache/cache[2][101] ), .B(n9546), .S0(n5235), .Y(
        n12013) );
  CLKMX2X2 U11197 ( .A(\I_cache/cache[1][101] ), .B(n9546), .S0(n5102), .Y(
        n12014) );
  CLKMX2X2 U11198 ( .A(\I_cache/cache[0][101] ), .B(n9546), .S0(n5150), .Y(
        n12015) );
  CLKMX2X2 U11199 ( .A(\I_cache/cache[7][100] ), .B(n9463), .S0(n5373), .Y(
        n12016) );
  CLKMX2X2 U11200 ( .A(\I_cache/cache[6][100] ), .B(n9463), .S0(n5417), .Y(
        n12017) );
  CLKMX2X2 U11201 ( .A(\I_cache/cache[5][100] ), .B(n9463), .S0(n5283), .Y(
        n12018) );
  CLKMX2X2 U11202 ( .A(\I_cache/cache[4][100] ), .B(n9463), .S0(n5326), .Y(
        n12019) );
  CLKMX2X2 U11203 ( .A(\I_cache/cache[3][100] ), .B(n9463), .S0(n5197), .Y(
        n12020) );
  CLKMX2X2 U11204 ( .A(\I_cache/cache[2][100] ), .B(n9463), .S0(n5239), .Y(
        n12021) );
  CLKMX2X2 U11205 ( .A(\I_cache/cache[1][100] ), .B(n9463), .S0(n5108), .Y(
        n12022) );
  CLKMX2X2 U11206 ( .A(\I_cache/cache[0][100] ), .B(n9463), .S0(n5152), .Y(
        n12023) );
  CLKMX2X2 U11207 ( .A(\I_cache/cache[7][98] ), .B(n9482), .S0(n5373), .Y(
        n12032) );
  CLKMX2X2 U11208 ( .A(\I_cache/cache[6][98] ), .B(n9482), .S0(n5417), .Y(
        n12033) );
  CLKMX2X2 U11209 ( .A(\I_cache/cache[5][98] ), .B(n9482), .S0(n5283), .Y(
        n12034) );
  CLKMX2X2 U11210 ( .A(\I_cache/cache[4][98] ), .B(n9482), .S0(n5326), .Y(
        n12035) );
  CLKMX2X2 U11211 ( .A(\I_cache/cache[3][98] ), .B(n9482), .S0(n5197), .Y(
        n12036) );
  CLKMX2X2 U11212 ( .A(\I_cache/cache[2][98] ), .B(n9482), .S0(n5239), .Y(
        n12037) );
  CLKMX2X2 U11213 ( .A(\I_cache/cache[1][98] ), .B(n9482), .S0(n5107), .Y(
        n12038) );
  CLKMX2X2 U11214 ( .A(\I_cache/cache[0][98] ), .B(n9482), .S0(n5152), .Y(
        n12039) );
  CLKMX2X2 U11215 ( .A(\I_cache/cache[6][97] ), .B(n9361), .S0(n5418), .Y(
        n12041) );
  CLKMX2X2 U11216 ( .A(\I_cache/cache[4][97] ), .B(n9361), .S0(n5327), .Y(
        n12043) );
  CLKMX2X2 U11217 ( .A(\I_cache/cache[3][97] ), .B(n9361), .S0(n5198), .Y(
        n12044) );
  CLKMX2X2 U11218 ( .A(\I_cache/cache[2][97] ), .B(n9361), .S0(n5240), .Y(
        n12045) );
  CLKMX2X2 U11219 ( .A(\I_cache/cache[1][97] ), .B(n9361), .S0(n5106), .Y(
        n12046) );
  CLKMX2X2 U11220 ( .A(\I_cache/cache[0][97] ), .B(n9361), .S0(n5153), .Y(
        n12047) );
  CLKMX2X2 U11221 ( .A(\I_cache/cache[7][96] ), .B(n9507), .S0(n5369), .Y(
        n12048) );
  CLKMX2X2 U11222 ( .A(\I_cache/cache[6][96] ), .B(n9507), .S0(n5417), .Y(
        n12049) );
  CLKMX2X2 U11223 ( .A(\I_cache/cache[5][96] ), .B(n9507), .S0(n5285), .Y(
        n12050) );
  CLKMX2X2 U11224 ( .A(\I_cache/cache[4][96] ), .B(n9507), .S0(n5325), .Y(
        n12051) );
  CLKMX2X2 U11225 ( .A(\I_cache/cache[3][96] ), .B(n9507), .S0(n5195), .Y(
        n12052) );
  CLKMX2X2 U11226 ( .A(\I_cache/cache[2][96] ), .B(n9507), .S0(n5242), .Y(
        n12053) );
  CLKMX2X2 U11227 ( .A(\I_cache/cache[1][96] ), .B(n9507), .S0(n5111), .Y(
        n12054) );
  CLKMX2X2 U11228 ( .A(\I_cache/cache[0][96] ), .B(n9507), .S0(n5148), .Y(
        n12055) );
  CLKMX2X2 U11229 ( .A(\I_cache/cache[7][95] ), .B(n11038), .S0(n5367), .Y(
        n12056) );
  CLKMX2X2 U11230 ( .A(\I_cache/cache[6][95] ), .B(n11038), .S0(n5411), .Y(
        n12057) );
  CLKMX2X2 U11231 ( .A(\I_cache/cache[5][95] ), .B(n11038), .S0(n5278), .Y(
        n12058) );
  CLKMX2X2 U11232 ( .A(\I_cache/cache[4][95] ), .B(n11038), .S0(n5320), .Y(
        n12059) );
  CLKMX2X2 U11233 ( .A(\I_cache/cache[3][95] ), .B(n11038), .S0(n5191), .Y(
        n12060) );
  CLKMX2X2 U11234 ( .A(\I_cache/cache[2][95] ), .B(n11038), .S0(n5233), .Y(
        n12061) );
  CLKMX2X2 U11235 ( .A(\I_cache/cache[1][95] ), .B(n11038), .S0(n5104), .Y(
        n12062) );
  CLKMX2X2 U11236 ( .A(\I_cache/cache[0][95] ), .B(n11038), .S0(n5146), .Y(
        n12063) );
  CLKMX2X2 U11237 ( .A(\I_cache/cache[7][94] ), .B(n9803), .S0(n5370), .Y(
        n12064) );
  CLKMX2X2 U11238 ( .A(\I_cache/cache[6][94] ), .B(n9803), .S0(n5414), .Y(
        n12065) );
  CLKMX2X2 U11239 ( .A(\I_cache/cache[5][94] ), .B(n9803), .S0(n5280), .Y(
        n12066) );
  CLKMX2X2 U11240 ( .A(\I_cache/cache[4][94] ), .B(n9803), .S0(n5323), .Y(
        n12067) );
  CLKMX2X2 U11241 ( .A(\I_cache/cache[3][94] ), .B(n9803), .S0(n5194), .Y(
        n12068) );
  CLKMX2X2 U11242 ( .A(\I_cache/cache[2][94] ), .B(n9803), .S0(n5236), .Y(
        n12069) );
  CLKMX2X2 U11243 ( .A(\I_cache/cache[1][94] ), .B(n9803), .S0(n5107), .Y(
        n12070) );
  CLKMX2X2 U11244 ( .A(\I_cache/cache[0][94] ), .B(n9803), .S0(n5149), .Y(
        n12071) );
  CLKMX2X2 U11245 ( .A(\I_cache/cache[7][93] ), .B(n11163), .S0(n5367), .Y(
        n12072) );
  CLKMX2X2 U11246 ( .A(\I_cache/cache[6][93] ), .B(n11163), .S0(n5411), .Y(
        n12073) );
  CLKMX2X2 U11247 ( .A(\I_cache/cache[5][93] ), .B(n11163), .S0(n5278), .Y(
        n12074) );
  CLKMX2X2 U11248 ( .A(\I_cache/cache[4][93] ), .B(n11163), .S0(n5320), .Y(
        n12075) );
  CLKMX2X2 U11249 ( .A(\I_cache/cache[3][93] ), .B(n11163), .S0(n5191), .Y(
        n12076) );
  CLKMX2X2 U11250 ( .A(\I_cache/cache[2][93] ), .B(n11163), .S0(n5233), .Y(
        n12077) );
  CLKMX2X2 U11251 ( .A(\I_cache/cache[1][93] ), .B(n11163), .S0(n5104), .Y(
        n12078) );
  CLKMX2X2 U11252 ( .A(\I_cache/cache[0][93] ), .B(n11163), .S0(n5146), .Y(
        n12079) );
  CLKMX2X2 U11253 ( .A(\I_cache/cache[7][92] ), .B(n9779), .S0(n5370), .Y(
        n12080) );
  CLKMX2X2 U11254 ( .A(\I_cache/cache[6][92] ), .B(n9779), .S0(n5414), .Y(
        n12081) );
  CLKMX2X2 U11255 ( .A(\I_cache/cache[5][92] ), .B(n9779), .S0(n5280), .Y(
        n12082) );
  CLKMX2X2 U11256 ( .A(\I_cache/cache[4][92] ), .B(n9779), .S0(n5323), .Y(
        n12083) );
  CLKMX2X2 U11257 ( .A(\I_cache/cache[3][92] ), .B(n9779), .S0(n5194), .Y(
        n12084) );
  CLKMX2X2 U11258 ( .A(\I_cache/cache[2][92] ), .B(n9779), .S0(n5236), .Y(
        n12085) );
  CLKMX2X2 U11259 ( .A(\I_cache/cache[1][92] ), .B(n9779), .S0(n5107), .Y(
        n12086) );
  CLKMX2X2 U11260 ( .A(\I_cache/cache[0][92] ), .B(n9779), .S0(n5149), .Y(
        n12087) );
  CLKMX2X2 U11261 ( .A(\I_cache/cache[7][91] ), .B(n9735), .S0(n5370), .Y(
        n12088) );
  CLKMX2X2 U11262 ( .A(\I_cache/cache[6][91] ), .B(n9735), .S0(n5414), .Y(
        n12089) );
  CLKMX2X2 U11263 ( .A(\I_cache/cache[5][91] ), .B(n9735), .S0(n5280), .Y(
        n12090) );
  CLKMX2X2 U11264 ( .A(\I_cache/cache[4][91] ), .B(n9735), .S0(n5323), .Y(
        n12091) );
  CLKMX2X2 U11265 ( .A(\I_cache/cache[3][91] ), .B(n9735), .S0(n5194), .Y(
        n12092) );
  CLKMX2X2 U11266 ( .A(\I_cache/cache[2][91] ), .B(n9735), .S0(n5236), .Y(
        n12093) );
  CLKMX2X2 U11267 ( .A(\I_cache/cache[1][91] ), .B(n9735), .S0(n5107), .Y(
        n12094) );
  CLKMX2X2 U11268 ( .A(\I_cache/cache[0][91] ), .B(n9735), .S0(n5149), .Y(
        n12095) );
  CLKMX2X2 U11269 ( .A(\I_cache/cache[7][90] ), .B(n9711), .S0(n5374), .Y(
        n12096) );
  CLKMX2X2 U11270 ( .A(\I_cache/cache[6][90] ), .B(n9711), .S0(n5419), .Y(
        n12097) );
  CLKMX2X2 U11271 ( .A(\I_cache/cache[3][90] ), .B(n9711), .S0(n5199), .Y(
        n12100) );
  CLKMX2X2 U11272 ( .A(\I_cache/cache[2][90] ), .B(n9711), .S0(n5241), .Y(
        n12101) );
  CLKMX2X2 U11273 ( .A(\I_cache/cache[1][90] ), .B(n9711), .S0(n5110), .Y(
        n12102) );
  CLKMX2X2 U11274 ( .A(\I_cache/cache[0][90] ), .B(n9711), .S0(n5154), .Y(
        n12103) );
  CLKMX2X2 U11275 ( .A(\I_cache/cache[7][89] ), .B(n10124), .S0(n5366), .Y(
        n12104) );
  CLKMX2X2 U11276 ( .A(\I_cache/cache[6][89] ), .B(n10124), .S0(n5410), .Y(
        n12105) );
  CLKMX2X2 U11277 ( .A(\I_cache/cache[5][89] ), .B(n10124), .S0(n5277), .Y(
        n12106) );
  CLKMX2X2 U11278 ( .A(\I_cache/cache[4][89] ), .B(n10124), .S0(n4678), .Y(
        n12107) );
  CLKMX2X2 U11279 ( .A(\I_cache/cache[3][89] ), .B(n10124), .S0(n5190), .Y(
        n12108) );
  CLKMX2X2 U11280 ( .A(\I_cache/cache[2][89] ), .B(n10124), .S0(n5233), .Y(
        n12109) );
  CLKMX2X2 U11281 ( .A(\I_cache/cache[1][89] ), .B(n10124), .S0(n5103), .Y(
        n12110) );
  CLKMX2X2 U11282 ( .A(\I_cache/cache[0][89] ), .B(n10124), .S0(n5145), .Y(
        n12111) );
  CLKMX2X2 U11283 ( .A(\I_cache/cache[7][88] ), .B(n9902), .S0(n5372), .Y(
        n12112) );
  CLKMX2X2 U11284 ( .A(\I_cache/cache[6][88] ), .B(n9902), .S0(n5416), .Y(
        n12113) );
  CLKMX2X2 U11285 ( .A(\I_cache/cache[5][88] ), .B(n9902), .S0(n5282), .Y(
        n12114) );
  CLKMX2X2 U11286 ( .A(\I_cache/cache[4][88] ), .B(n9902), .S0(n5325), .Y(
        n12115) );
  CLKMX2X2 U11287 ( .A(\I_cache/cache[3][88] ), .B(n9902), .S0(n5196), .Y(
        n12116) );
  CLKMX2X2 U11288 ( .A(\I_cache/cache[2][88] ), .B(n9902), .S0(n5238), .Y(
        n12117) );
  CLKMX2X2 U11289 ( .A(\I_cache/cache[1][88] ), .B(n9902), .S0(n5109), .Y(
        n12118) );
  CLKMX2X2 U11290 ( .A(\I_cache/cache[0][88] ), .B(n9902), .S0(n5151), .Y(
        n12119) );
  CLKMX2X2 U11291 ( .A(\I_cache/cache[7][87] ), .B(n9926), .S0(n5372), .Y(
        n12120) );
  CLKMX2X2 U11292 ( .A(\I_cache/cache[6][87] ), .B(n9926), .S0(n5416), .Y(
        n12121) );
  CLKMX2X2 U11293 ( .A(\I_cache/cache[5][87] ), .B(n9926), .S0(n5282), .Y(
        n12122) );
  CLKMX2X2 U11294 ( .A(\I_cache/cache[4][87] ), .B(n9926), .S0(n5325), .Y(
        n12123) );
  CLKMX2X2 U11295 ( .A(\I_cache/cache[3][87] ), .B(n9926), .S0(n5196), .Y(
        n12124) );
  CLKMX2X2 U11296 ( .A(\I_cache/cache[2][87] ), .B(n9926), .S0(n5238), .Y(
        n12125) );
  CLKMX2X2 U11297 ( .A(\I_cache/cache[1][87] ), .B(n9926), .S0(n5109), .Y(
        n12126) );
  CLKMX2X2 U11298 ( .A(\I_cache/cache[0][87] ), .B(n9926), .S0(n5151), .Y(
        n12127) );
  CLKMX2X2 U11299 ( .A(\I_cache/cache[7][86] ), .B(n9858), .S0(n5369), .Y(
        n12128) );
  CLKMX2X2 U11300 ( .A(\I_cache/cache[6][86] ), .B(n9858), .S0(n5413), .Y(
        n12129) );
  CLKMX2X2 U11301 ( .A(\I_cache/cache[5][86] ), .B(n9858), .S0(n5279), .Y(
        n12130) );
  CLKMX2X2 U11302 ( .A(\I_cache/cache[4][86] ), .B(n9858), .S0(n5322), .Y(
        n12131) );
  CLKMX2X2 U11303 ( .A(\I_cache/cache[3][86] ), .B(n9858), .S0(n5193), .Y(
        n12132) );
  CLKMX2X2 U11304 ( .A(\I_cache/cache[2][86] ), .B(n9858), .S0(n5235), .Y(
        n12133) );
  CLKMX2X2 U11305 ( .A(\I_cache/cache[1][86] ), .B(n9858), .S0(n5106), .Y(
        n12134) );
  CLKMX2X2 U11306 ( .A(\I_cache/cache[0][86] ), .B(n9858), .S0(n5148), .Y(
        n12135) );
  CLKMX2X2 U11307 ( .A(\I_cache/cache[7][85] ), .B(n9878), .S0(n5369), .Y(
        n12136) );
  CLKMX2X2 U11308 ( .A(\I_cache/cache[6][85] ), .B(n9878), .S0(n5413), .Y(
        n12137) );
  CLKMX2X2 U11309 ( .A(\I_cache/cache[5][85] ), .B(n9878), .S0(n5279), .Y(
        n12138) );
  CLKMX2X2 U11310 ( .A(\I_cache/cache[4][85] ), .B(n9878), .S0(n5322), .Y(
        n12139) );
  CLKMX2X2 U11311 ( .A(\I_cache/cache[3][85] ), .B(n9878), .S0(n5193), .Y(
        n12140) );
  CLKMX2X2 U11312 ( .A(\I_cache/cache[2][85] ), .B(n9878), .S0(n5235), .Y(
        n12141) );
  CLKMX2X2 U11313 ( .A(\I_cache/cache[1][85] ), .B(n9878), .S0(n5106), .Y(
        n12142) );
  CLKMX2X2 U11314 ( .A(\I_cache/cache[0][85] ), .B(n9878), .S0(n5148), .Y(
        n12143) );
  CLKMX2X2 U11315 ( .A(\I_cache/cache[7][84] ), .B(n10022), .S0(n5371), .Y(
        n12144) );
  CLKMX2X2 U11316 ( .A(\I_cache/cache[6][84] ), .B(n10022), .S0(n5415), .Y(
        n12145) );
  CLKMX2X2 U11317 ( .A(\I_cache/cache[5][84] ), .B(n10022), .S0(n5281), .Y(
        n12146) );
  CLKMX2X2 U11318 ( .A(\I_cache/cache[4][84] ), .B(n10022), .S0(n5324), .Y(
        n12147) );
  CLKMX2X2 U11319 ( .A(\I_cache/cache[3][84] ), .B(n10022), .S0(n5195), .Y(
        n12148) );
  CLKMX2X2 U11320 ( .A(\I_cache/cache[2][84] ), .B(n10022), .S0(n5237), .Y(
        n12149) );
  CLKMX2X2 U11321 ( .A(\I_cache/cache[1][84] ), .B(n10022), .S0(n5108), .Y(
        n12150) );
  CLKMX2X2 U11322 ( .A(\I_cache/cache[0][84] ), .B(n10022), .S0(n5150), .Y(
        n12151) );
  CLKMX2X2 U11323 ( .A(\I_cache/cache[7][83] ), .B(n9993), .S0(n5370), .Y(
        n12152) );
  CLKMX2X2 U11324 ( .A(\I_cache/cache[6][83] ), .B(n9993), .S0(n5414), .Y(
        n12153) );
  CLKMX2X2 U11325 ( .A(\I_cache/cache[5][83] ), .B(n9993), .S0(n5280), .Y(
        n12154) );
  CLKMX2X2 U11326 ( .A(\I_cache/cache[4][83] ), .B(n9993), .S0(n5323), .Y(
        n12155) );
  CLKMX2X2 U11327 ( .A(\I_cache/cache[3][83] ), .B(n9993), .S0(n5194), .Y(
        n12156) );
  CLKMX2X2 U11328 ( .A(\I_cache/cache[2][83] ), .B(n9993), .S0(n5236), .Y(
        n12157) );
  CLKMX2X2 U11329 ( .A(\I_cache/cache[1][83] ), .B(n9993), .S0(n5107), .Y(
        n12158) );
  CLKMX2X2 U11330 ( .A(\I_cache/cache[0][83] ), .B(n9993), .S0(n5149), .Y(
        n12159) );
  CLKMX2X2 U11331 ( .A(\I_cache/cache[6][82] ), .B(n10046), .S0(n5415), .Y(
        n12161) );
  CLKMX2X2 U11332 ( .A(\I_cache/cache[5][82] ), .B(n10046), .S0(n5281), .Y(
        n12162) );
  CLKMX2X2 U11333 ( .A(\I_cache/cache[4][82] ), .B(n10046), .S0(n5324), .Y(
        n12163) );
  CLKMX2X2 U11334 ( .A(\I_cache/cache[3][82] ), .B(n10046), .S0(n5195), .Y(
        n12164) );
  CLKMX2X2 U11335 ( .A(\I_cache/cache[2][82] ), .B(n10046), .S0(n5237), .Y(
        n12165) );
  CLKMX2X2 U11336 ( .A(\I_cache/cache[0][82] ), .B(n10046), .S0(n5150), .Y(
        n12167) );
  CLKMX2X2 U11337 ( .A(\I_cache/cache[7][81] ), .B(n11145), .S0(n5367), .Y(
        n12168) );
  CLKMX2X2 U11338 ( .A(\I_cache/cache[6][81] ), .B(n11145), .S0(n5411), .Y(
        n12169) );
  CLKMX2X2 U11339 ( .A(\I_cache/cache[5][81] ), .B(n11145), .S0(n5278), .Y(
        n12170) );
  CLKMX2X2 U11340 ( .A(\I_cache/cache[4][81] ), .B(n11145), .S0(n5320), .Y(
        n12171) );
  CLKMX2X2 U11341 ( .A(\I_cache/cache[3][81] ), .B(n11145), .S0(n5191), .Y(
        n12172) );
  CLKMX2X2 U11342 ( .A(\I_cache/cache[2][81] ), .B(n11145), .S0(n5233), .Y(
        n12173) );
  CLKMX2X2 U11343 ( .A(\I_cache/cache[1][81] ), .B(n11145), .S0(n5104), .Y(
        n12174) );
  CLKMX2X2 U11344 ( .A(\I_cache/cache[0][81] ), .B(n11145), .S0(n5146), .Y(
        n12175) );
  CLKMX2X2 U11345 ( .A(\I_cache/cache[6][80] ), .B(n10075), .S0(n5415), .Y(
        n12177) );
  CLKMX2X2 U11346 ( .A(\I_cache/cache[5][80] ), .B(n10075), .S0(n5281), .Y(
        n12178) );
  CLKMX2X2 U11347 ( .A(\I_cache/cache[4][80] ), .B(n10075), .S0(n5324), .Y(
        n12179) );
  CLKMX2X2 U11348 ( .A(\I_cache/cache[2][80] ), .B(n10075), .S0(n5237), .Y(
        n12181) );
  CLKMX2X2 U11349 ( .A(\I_cache/cache[1][80] ), .B(n10075), .S0(n5108), .Y(
        n12182) );
  CLKMX2X2 U11350 ( .A(\I_cache/cache[0][80] ), .B(n10075), .S0(n5150), .Y(
        n12183) );
  CLKMX2X2 U11351 ( .A(\I_cache/cache[7][78] ), .B(n9407), .S0(n5366), .Y(
        n12192) );
  CLKMX2X2 U11352 ( .A(\I_cache/cache[6][78] ), .B(n9407), .S0(n5418), .Y(
        n12193) );
  CLKMX2X2 U11353 ( .A(\I_cache/cache[5][78] ), .B(n9407), .S0(n5284), .Y(
        n12194) );
  CLKMX2X2 U11354 ( .A(\I_cache/cache[4][78] ), .B(n9407), .S0(n5326), .Y(
        n12195) );
  CLKMX2X2 U11355 ( .A(\I_cache/cache[3][78] ), .B(n9407), .S0(n5198), .Y(
        n12196) );
  CLKMX2X2 U11356 ( .A(\I_cache/cache[2][78] ), .B(n9407), .S0(n5240), .Y(
        n12197) );
  CLKMX2X2 U11357 ( .A(\I_cache/cache[1][78] ), .B(n9407), .S0(n5109), .Y(
        n12198) );
  CLKMX2X2 U11358 ( .A(\I_cache/cache[0][78] ), .B(n9407), .S0(n5153), .Y(
        n12199) );
  CLKMX2X2 U11359 ( .A(\I_cache/cache[7][77] ), .B(n9387), .S0(n5367), .Y(
        n12200) );
  CLKMX2X2 U11360 ( .A(\I_cache/cache[6][77] ), .B(n9387), .S0(n5418), .Y(
        n12201) );
  CLKMX2X2 U11361 ( .A(\I_cache/cache[5][77] ), .B(n9387), .S0(n5284), .Y(
        n12202) );
  CLKMX2X2 U11362 ( .A(\I_cache/cache[4][77] ), .B(n9387), .S0(n5322), .Y(
        n12203) );
  CLKMX2X2 U11363 ( .A(\I_cache/cache[3][77] ), .B(n9387), .S0(n5198), .Y(
        n12204) );
  CLKMX2X2 U11364 ( .A(\I_cache/cache[2][77] ), .B(n9387), .S0(n5240), .Y(
        n12205) );
  CLKMX2X2 U11365 ( .A(\I_cache/cache[1][77] ), .B(n9387), .S0(n5106), .Y(
        n12206) );
  CLKMX2X2 U11366 ( .A(\I_cache/cache[0][77] ), .B(n9387), .S0(n5153), .Y(
        n12207) );
  CLKMX2X2 U11367 ( .A(\I_cache/cache[7][76] ), .B(n10100), .S0(n5366), .Y(
        n12208) );
  CLKMX2X2 U11368 ( .A(\I_cache/cache[6][76] ), .B(n10100), .S0(n5410), .Y(
        n12209) );
  CLKMX2X2 U11369 ( .A(\I_cache/cache[4][76] ), .B(n10100), .S0(n4681), .Y(
        n12211) );
  CLKMX2X2 U11370 ( .A(\I_cache/cache[3][76] ), .B(n10100), .S0(n5190), .Y(
        n12212) );
  CLKMX2X2 U11371 ( .A(\I_cache/cache[2][76] ), .B(n10100), .S0(n5236), .Y(
        n12213) );
  CLKMX2X2 U11372 ( .A(\I_cache/cache[1][76] ), .B(n10100), .S0(n5103), .Y(
        n12214) );
  CLKMX2X2 U11373 ( .A(\I_cache/cache[0][76] ), .B(n10100), .S0(n5145), .Y(
        n12215) );
  CLKMX2X2 U11374 ( .A(\I_cache/cache[7][75] ), .B(n9969), .S0(n5372), .Y(
        n12216) );
  CLKMX2X2 U11375 ( .A(\I_cache/cache[6][75] ), .B(n9969), .S0(n5416), .Y(
        n12217) );
  CLKMX2X2 U11376 ( .A(\I_cache/cache[5][75] ), .B(n9969), .S0(n5282), .Y(
        n12218) );
  CLKMX2X2 U11377 ( .A(\I_cache/cache[4][75] ), .B(n9969), .S0(n5325), .Y(
        n12219) );
  CLKMX2X2 U11378 ( .A(\I_cache/cache[3][75] ), .B(n9969), .S0(n5196), .Y(
        n12220) );
  CLKMX2X2 U11379 ( .A(\I_cache/cache[2][75] ), .B(n9969), .S0(n5238), .Y(
        n12221) );
  CLKMX2X2 U11380 ( .A(\I_cache/cache[1][75] ), .B(n9969), .S0(n5109), .Y(
        n12222) );
  CLKMX2X2 U11381 ( .A(\I_cache/cache[0][75] ), .B(n9969), .S0(n5151), .Y(
        n12223) );
  CLKMX2X2 U11382 ( .A(\I_cache/cache[7][74] ), .B(n9673), .S0(n5374), .Y(
        n12224) );
  CLKMX2X2 U11383 ( .A(\I_cache/cache[6][74] ), .B(n9673), .S0(n5419), .Y(
        n12225) );
  CLKMX2X2 U11384 ( .A(\I_cache/cache[4][74] ), .B(n9673), .S0(n5327), .Y(
        n12227) );
  CLKMX2X2 U11385 ( .A(\I_cache/cache[3][74] ), .B(n9673), .S0(n5199), .Y(
        n12228) );
  CLKMX2X2 U11386 ( .A(\I_cache/cache[2][74] ), .B(n9673), .S0(n5241), .Y(
        n12229) );
  CLKMX2X2 U11387 ( .A(\I_cache/cache[1][74] ), .B(n9673), .S0(n5110), .Y(
        n12230) );
  CLKMX2X2 U11388 ( .A(\I_cache/cache[0][74] ), .B(n9673), .S0(n5154), .Y(
        n12231) );
  CLKMX2X2 U11389 ( .A(\I_cache/cache[7][73] ), .B(n9640), .S0(n5374), .Y(
        n12232) );
  CLKMX2X2 U11390 ( .A(\I_cache/cache[6][73] ), .B(n9640), .S0(n5419), .Y(
        n12233) );
  CLKMX2X2 U11391 ( .A(\I_cache/cache[4][73] ), .B(n9640), .S0(n5327), .Y(
        n12235) );
  CLKMX2X2 U11392 ( .A(\I_cache/cache[3][73] ), .B(n9640), .S0(n5199), .Y(
        n12236) );
  CLKMX2X2 U11393 ( .A(\I_cache/cache[2][73] ), .B(n9640), .S0(n5241), .Y(
        n12237) );
  CLKMX2X2 U11394 ( .A(\I_cache/cache[1][73] ), .B(n9640), .S0(n5110), .Y(
        n12238) );
  CLKMX2X2 U11395 ( .A(\I_cache/cache[0][73] ), .B(n9640), .S0(n5154), .Y(
        n12239) );
  CLKMX2X2 U11396 ( .A(\I_cache/cache[7][72] ), .B(n9416), .S0(n5372), .Y(
        n12240) );
  CLKMX2X2 U11397 ( .A(\I_cache/cache[6][72] ), .B(n9416), .S0(n5416), .Y(
        n12241) );
  CLKMX2X2 U11398 ( .A(\I_cache/cache[5][72] ), .B(n9416), .S0(n5282), .Y(
        n12242) );
  CLKMX2X2 U11399 ( .A(\I_cache/cache[4][72] ), .B(n9416), .S0(n5325), .Y(
        n12243) );
  CLKMX2X2 U11400 ( .A(\I_cache/cache[3][72] ), .B(n9416), .S0(n5196), .Y(
        n12244) );
  CLKMX2X2 U11401 ( .A(\I_cache/cache[2][72] ), .B(n9416), .S0(n5238), .Y(
        n12245) );
  CLKMX2X2 U11402 ( .A(\I_cache/cache[1][72] ), .B(n9416), .S0(n5109), .Y(
        n12246) );
  CLKMX2X2 U11403 ( .A(\I_cache/cache[0][72] ), .B(n9416), .S0(n5151), .Y(
        n12247) );
  CLKMX2X2 U11404 ( .A(\I_cache/cache[7][71] ), .B(n9820), .S0(n5368), .Y(
        n12248) );
  CLKMX2X2 U11405 ( .A(\I_cache/cache[6][71] ), .B(n9820), .S0(n5412), .Y(
        n12249) );
  CLKMX2X2 U11406 ( .A(\I_cache/cache[5][71] ), .B(n9820), .S0(n5282), .Y(
        n12250) );
  CLKMX2X2 U11407 ( .A(\I_cache/cache[4][71] ), .B(n9820), .S0(n5321), .Y(
        n12251) );
  CLKMX2X2 U11408 ( .A(\I_cache/cache[3][71] ), .B(n9820), .S0(n5192), .Y(
        n12252) );
  CLKMX2X2 U11409 ( .A(\I_cache/cache[2][71] ), .B(n9820), .S0(n5234), .Y(
        n12253) );
  CLKMX2X2 U11410 ( .A(\I_cache/cache[1][71] ), .B(n9820), .S0(n5105), .Y(
        n12254) );
  CLKMX2X2 U11411 ( .A(\I_cache/cache[0][71] ), .B(n9820), .S0(n5147), .Y(
        n12255) );
  CLKMX2X2 U11412 ( .A(\I_cache/cache[7][70] ), .B(n9450), .S0(n5373), .Y(
        n12256) );
  CLKMX2X2 U11413 ( .A(\I_cache/cache[6][70] ), .B(n9450), .S0(n5417), .Y(
        n12257) );
  CLKMX2X2 U11414 ( .A(\I_cache/cache[5][70] ), .B(n9450), .S0(n5283), .Y(
        n12258) );
  CLKMX2X2 U11415 ( .A(\I_cache/cache[4][70] ), .B(n9450), .S0(n5326), .Y(
        n12259) );
  CLKMX2X2 U11416 ( .A(\I_cache/cache[3][70] ), .B(n9450), .S0(n5197), .Y(
        n12260) );
  CLKMX2X2 U11417 ( .A(\I_cache/cache[2][70] ), .B(n9450), .S0(n5239), .Y(
        n12261) );
  CLKMX2X2 U11418 ( .A(\I_cache/cache[1][70] ), .B(n9450), .S0(n5111), .Y(
        n12262) );
  CLKMX2X2 U11419 ( .A(\I_cache/cache[0][70] ), .B(n9450), .S0(n5152), .Y(
        n12263) );
  CLKMX2X2 U11420 ( .A(\I_cache/cache[7][69] ), .B(n9537), .S0(n5374), .Y(
        n12264) );
  CLKMX2X2 U11421 ( .A(\I_cache/cache[6][69] ), .B(n9537), .S0(n5413), .Y(
        n12265) );
  CLKMX2X2 U11422 ( .A(\I_cache/cache[5][69] ), .B(n9537), .S0(n5285), .Y(
        n12266) );
  CLKMX2X2 U11423 ( .A(\I_cache/cache[4][69] ), .B(n9537), .S0(n5324), .Y(
        n12267) );
  CLKMX2X2 U11424 ( .A(\I_cache/cache[3][69] ), .B(n9537), .S0(n5199), .Y(
        n12268) );
  CLKMX2X2 U11425 ( .A(\I_cache/cache[2][69] ), .B(n9537), .S0(n5242), .Y(
        n12269) );
  CLKMX2X2 U11426 ( .A(\I_cache/cache[1][69] ), .B(n9537), .S0(n5111), .Y(
        n12270) );
  CLKMX2X2 U11427 ( .A(\I_cache/cache[0][69] ), .B(n9537), .S0(n5154), .Y(
        n12271) );
  CLKMX2X2 U11428 ( .A(\I_cache/cache[7][68] ), .B(n9472), .S0(n5373), .Y(
        n12272) );
  CLKMX2X2 U11429 ( .A(\I_cache/cache[6][68] ), .B(n9472), .S0(n5417), .Y(
        n12273) );
  CLKMX2X2 U11430 ( .A(\I_cache/cache[5][68] ), .B(n9472), .S0(n5283), .Y(
        n12274) );
  CLKMX2X2 U11431 ( .A(\I_cache/cache[4][68] ), .B(n9472), .S0(n5326), .Y(
        n12275) );
  CLKMX2X2 U11432 ( .A(\I_cache/cache[3][68] ), .B(n9472), .S0(n5197), .Y(
        n12276) );
  CLKMX2X2 U11433 ( .A(\I_cache/cache[2][68] ), .B(n9472), .S0(n5239), .Y(
        n12277) );
  CLKMX2X2 U11434 ( .A(\I_cache/cache[1][68] ), .B(n9472), .S0(n5102), .Y(
        n12278) );
  CLKMX2X2 U11435 ( .A(\I_cache/cache[0][68] ), .B(n9472), .S0(n5152), .Y(
        n12279) );
  CLKMX2X2 U11436 ( .A(\I_cache/cache[7][67] ), .B(n9527), .S0(n5373), .Y(
        n12280) );
  CLKMX2X2 U11437 ( .A(\I_cache/cache[6][67] ), .B(n9527), .S0(n5416), .Y(
        n12281) );
  CLKMX2X2 U11438 ( .A(\I_cache/cache[5][67] ), .B(n9527), .S0(n5285), .Y(
        n12282) );
  CLKMX2X2 U11439 ( .A(\I_cache/cache[4][67] ), .B(n9527), .S0(n5325), .Y(
        n12283) );
  CLKMX2X2 U11440 ( .A(\I_cache/cache[3][67] ), .B(n9527), .S0(n5193), .Y(
        n12284) );
  CLKMX2X2 U11441 ( .A(\I_cache/cache[2][67] ), .B(n9527), .S0(n5242), .Y(
        n12285) );
  CLKMX2X2 U11442 ( .A(\I_cache/cache[1][67] ), .B(n9527), .S0(n5111), .Y(
        n12286) );
  CLKMX2X2 U11443 ( .A(\I_cache/cache[0][67] ), .B(n9527), .S0(n5152), .Y(
        n12287) );
  CLKMX2X2 U11444 ( .A(\I_cache/cache[7][66] ), .B(n9492), .S0(n5371), .Y(
        n12288) );
  CLKMX2X2 U11445 ( .A(\I_cache/cache[6][66] ), .B(n9492), .S0(n5417), .Y(
        n12289) );
  CLKMX2X2 U11446 ( .A(\I_cache/cache[5][66] ), .B(n9492), .S0(n5285), .Y(
        n12290) );
  CLKMX2X2 U11447 ( .A(\I_cache/cache[4][66] ), .B(n9492), .S0(n5324), .Y(
        n12291) );
  CLKMX2X2 U11448 ( .A(\I_cache/cache[3][66] ), .B(n9492), .S0(n5195), .Y(
        n12292) );
  CLKMX2X2 U11449 ( .A(\I_cache/cache[2][66] ), .B(n9492), .S0(n5242), .Y(
        n12293) );
  CLKMX2X2 U11450 ( .A(\I_cache/cache[1][66] ), .B(n9492), .S0(n5111), .Y(
        n12294) );
  CLKMX2X2 U11451 ( .A(\I_cache/cache[0][66] ), .B(n9492), .S0(n5148), .Y(
        n12295) );
  CLKMX2X2 U11452 ( .A(\I_cache/cache[7][65] ), .B(n10999), .S0(n5368), .Y(
        n12296) );
  CLKMX2X2 U11453 ( .A(\I_cache/cache[6][65] ), .B(n10999), .S0(n5412), .Y(
        n12297) );
  CLKMX2X2 U11454 ( .A(\I_cache/cache[5][65] ), .B(n10999), .S0(n5277), .Y(
        n12298) );
  CLKMX2X2 U11455 ( .A(\I_cache/cache[4][65] ), .B(n10999), .S0(n5321), .Y(
        n12299) );
  CLKMX2X2 U11456 ( .A(\I_cache/cache[3][65] ), .B(n10999), .S0(n5192), .Y(
        n12300) );
  CLKMX2X2 U11457 ( .A(\I_cache/cache[2][65] ), .B(n10999), .S0(n5234), .Y(
        n12301) );
  CLKMX2X2 U11458 ( .A(\I_cache/cache[1][65] ), .B(n10999), .S0(n5105), .Y(
        n12302) );
  CLKMX2X2 U11459 ( .A(\I_cache/cache[0][65] ), .B(n10999), .S0(n5147), .Y(
        n12303) );
  CLKMX2X2 U11460 ( .A(\I_cache/cache[7][64] ), .B(n9683), .S0(n5374), .Y(
        n12304) );
  CLKMX2X2 U11461 ( .A(\I_cache/cache[6][64] ), .B(n9683), .S0(n5419), .Y(
        n12305) );
  CLKMX2X2 U11462 ( .A(\I_cache/cache[3][64] ), .B(n9683), .S0(n5199), .Y(
        n12308) );
  CLKMX2X2 U11463 ( .A(\I_cache/cache[2][64] ), .B(n9683), .S0(n5241), .Y(
        n12309) );
  CLKMX2X2 U11464 ( .A(\I_cache/cache[1][64] ), .B(n9683), .S0(n5110), .Y(
        n12310) );
  CLKMX2X2 U11465 ( .A(\I_cache/cache[0][64] ), .B(n9683), .S0(n5154), .Y(
        n12311) );
  CLKMX2X2 U11466 ( .A(\I_cache/cache[7][63] ), .B(n11036), .S0(n5368), .Y(
        n12312) );
  CLKMX2X2 U11467 ( .A(\I_cache/cache[6][63] ), .B(n11036), .S0(n5412), .Y(
        n12313) );
  CLKMX2X2 U11468 ( .A(\I_cache/cache[5][63] ), .B(n11036), .S0(n5284), .Y(
        n12314) );
  CLKMX2X2 U11469 ( .A(\I_cache/cache[4][63] ), .B(n11036), .S0(n5321), .Y(
        n12315) );
  CLKMX2X2 U11470 ( .A(\I_cache/cache[3][63] ), .B(n11036), .S0(n5192), .Y(
        n12316) );
  CLKMX2X2 U11471 ( .A(\I_cache/cache[2][63] ), .B(n11036), .S0(n5234), .Y(
        n12317) );
  CLKMX2X2 U11472 ( .A(\I_cache/cache[1][63] ), .B(n11036), .S0(n5105), .Y(
        n12318) );
  CLKMX2X2 U11473 ( .A(\I_cache/cache[0][63] ), .B(n11036), .S0(n5147), .Y(
        n12319) );
  CLKMX2X2 U11474 ( .A(\I_cache/cache[7][62] ), .B(n9793), .S0(n5370), .Y(
        n12320) );
  CLKMX2X2 U11475 ( .A(\I_cache/cache[6][62] ), .B(n9793), .S0(n5414), .Y(
        n12321) );
  CLKMX2X2 U11476 ( .A(\I_cache/cache[5][62] ), .B(n9793), .S0(n5280), .Y(
        n12322) );
  CLKMX2X2 U11477 ( .A(\I_cache/cache[4][62] ), .B(n9793), .S0(n5323), .Y(
        n12323) );
  CLKMX2X2 U11478 ( .A(\I_cache/cache[3][62] ), .B(n9793), .S0(n5194), .Y(
        n12324) );
  CLKMX2X2 U11479 ( .A(\I_cache/cache[2][62] ), .B(n9793), .S0(n5236), .Y(
        n12325) );
  CLKMX2X2 U11480 ( .A(\I_cache/cache[1][62] ), .B(n9793), .S0(n5107), .Y(
        n12326) );
  CLKMX2X2 U11481 ( .A(\I_cache/cache[0][62] ), .B(n9793), .S0(n5149), .Y(
        n12327) );
  CLKMX2X2 U11482 ( .A(\I_cache/cache[7][61] ), .B(n11159), .S0(n5367), .Y(
        n12328) );
  CLKMX2X2 U11483 ( .A(\I_cache/cache[6][61] ), .B(n11159), .S0(n5411), .Y(
        n12329) );
  CLKMX2X2 U11484 ( .A(\I_cache/cache[5][61] ), .B(n11159), .S0(n5278), .Y(
        n12330) );
  CLKMX2X2 U11485 ( .A(\I_cache/cache[4][61] ), .B(n11159), .S0(n5320), .Y(
        n12331) );
  CLKMX2X2 U11486 ( .A(\I_cache/cache[3][61] ), .B(n11159), .S0(n5191), .Y(
        n12332) );
  CLKMX2X2 U11487 ( .A(\I_cache/cache[2][61] ), .B(n11159), .S0(n5233), .Y(
        n12333) );
  CLKMX2X2 U11488 ( .A(\I_cache/cache[1][61] ), .B(n11159), .S0(n5104), .Y(
        n12334) );
  CLKMX2X2 U11489 ( .A(\I_cache/cache[0][61] ), .B(n11159), .S0(n5146), .Y(
        n12335) );
  CLKMX2X2 U11490 ( .A(\I_cache/cache[7][60] ), .B(n9769), .S0(n5370), .Y(
        n12336) );
  CLKMX2X2 U11491 ( .A(\I_cache/cache[6][60] ), .B(n9769), .S0(n5414), .Y(
        n12337) );
  CLKMX2X2 U11492 ( .A(\I_cache/cache[5][60] ), .B(n9769), .S0(n5280), .Y(
        n12338) );
  CLKMX2X2 U11493 ( .A(\I_cache/cache[4][60] ), .B(n9769), .S0(n5323), .Y(
        n12339) );
  CLKMX2X2 U11494 ( .A(\I_cache/cache[3][60] ), .B(n9769), .S0(n5194), .Y(
        n12340) );
  CLKMX2X2 U11495 ( .A(\I_cache/cache[2][60] ), .B(n9769), .S0(n5236), .Y(
        n12341) );
  CLKMX2X2 U11496 ( .A(\I_cache/cache[1][60] ), .B(n9769), .S0(n5107), .Y(
        n12342) );
  CLKMX2X2 U11497 ( .A(\I_cache/cache[0][60] ), .B(n9769), .S0(n5149), .Y(
        n12343) );
  CLKMX2X2 U11498 ( .A(\I_cache/cache[7][59] ), .B(n9725), .S0(n5369), .Y(
        n12344) );
  CLKMX2X2 U11499 ( .A(\I_cache/cache[6][59] ), .B(n9725), .S0(n5413), .Y(
        n12345) );
  CLKMX2X2 U11500 ( .A(\I_cache/cache[5][59] ), .B(n9725), .S0(n5279), .Y(
        n12346) );
  CLKMX2X2 U11501 ( .A(\I_cache/cache[4][59] ), .B(n9725), .S0(n5322), .Y(
        n12347) );
  CLKMX2X2 U11502 ( .A(\I_cache/cache[3][59] ), .B(n9725), .S0(n5193), .Y(
        n12348) );
  CLKMX2X2 U11503 ( .A(\I_cache/cache[2][59] ), .B(n9725), .S0(n5235), .Y(
        n12349) );
  CLKMX2X2 U11504 ( .A(\I_cache/cache[1][59] ), .B(n9725), .S0(n5106), .Y(
        n12350) );
  CLKMX2X2 U11505 ( .A(\I_cache/cache[0][59] ), .B(n9725), .S0(n5148), .Y(
        n12351) );
  CLKMX2X2 U11506 ( .A(\I_cache/cache[7][58] ), .B(n9701), .S0(n5374), .Y(
        n12352) );
  CLKMX2X2 U11507 ( .A(\I_cache/cache[6][58] ), .B(n9701), .S0(n5419), .Y(
        n12353) );
  CLKMX2X2 U11508 ( .A(\I_cache/cache[5][58] ), .B(n9701), .S0(n5282), .Y(
        n12354) );
  CLKMX2X2 U11509 ( .A(\I_cache/cache[4][58] ), .B(n9701), .S0(n5327), .Y(
        n12355) );
  CLKMX2X2 U11510 ( .A(\I_cache/cache[3][58] ), .B(n9701), .S0(n5199), .Y(
        n12356) );
  CLKMX2X2 U11511 ( .A(\I_cache/cache[2][58] ), .B(n9701), .S0(n5241), .Y(
        n12357) );
  CLKMX2X2 U11512 ( .A(\I_cache/cache[1][58] ), .B(n9701), .S0(n5110), .Y(
        n12358) );
  CLKMX2X2 U11513 ( .A(\I_cache/cache[0][58] ), .B(n9701), .S0(n5154), .Y(
        n12359) );
  CLKMX2X2 U11514 ( .A(\I_cache/cache[7][57] ), .B(n10114), .S0(n5366), .Y(
        n12360) );
  CLKMX2X2 U11515 ( .A(\I_cache/cache[6][57] ), .B(n10114), .S0(n5410), .Y(
        n12361) );
  CLKMX2X2 U11516 ( .A(\I_cache/cache[5][57] ), .B(n10114), .S0(n5277), .Y(
        n12362) );
  CLKMX2X2 U11517 ( .A(\I_cache/cache[4][57] ), .B(n10114), .S0(n4676), .Y(
        n12363) );
  CLKMX2X2 U11518 ( .A(\I_cache/cache[3][57] ), .B(n10114), .S0(n5190), .Y(
        n12364) );
  CLKMX2X2 U11519 ( .A(\I_cache/cache[2][57] ), .B(n10114), .S0(n5237), .Y(
        n12365) );
  CLKMX2X2 U11520 ( .A(\I_cache/cache[1][57] ), .B(n10114), .S0(n5103), .Y(
        n12366) );
  CLKMX2X2 U11521 ( .A(\I_cache/cache[0][57] ), .B(n10114), .S0(n5145), .Y(
        n12367) );
  CLKMX2X2 U11522 ( .A(\I_cache/cache[7][56] ), .B(n9892), .S0(n5369), .Y(
        n12368) );
  CLKMX2X2 U11523 ( .A(\I_cache/cache[6][56] ), .B(n9892), .S0(n5413), .Y(
        n12369) );
  CLKMX2X2 U11524 ( .A(\I_cache/cache[5][56] ), .B(n9892), .S0(n5279), .Y(
        n12370) );
  CLKMX2X2 U11525 ( .A(\I_cache/cache[4][56] ), .B(n9892), .S0(n5322), .Y(
        n12371) );
  CLKMX2X2 U11526 ( .A(\I_cache/cache[3][56] ), .B(n9892), .S0(n5193), .Y(
        n12372) );
  CLKMX2X2 U11527 ( .A(\I_cache/cache[2][56] ), .B(n9892), .S0(n5235), .Y(
        n12373) );
  CLKMX2X2 U11528 ( .A(\I_cache/cache[1][56] ), .B(n9892), .S0(n5106), .Y(
        n12374) );
  CLKMX2X2 U11529 ( .A(\I_cache/cache[0][56] ), .B(n9892), .S0(n5148), .Y(
        n12375) );
  CLKMX2X2 U11530 ( .A(\I_cache/cache[7][55] ), .B(n9916), .S0(n5372), .Y(
        n12376) );
  CLKMX2X2 U11531 ( .A(\I_cache/cache[6][55] ), .B(n9916), .S0(n5416), .Y(
        n12377) );
  CLKMX2X2 U11532 ( .A(\I_cache/cache[5][55] ), .B(n9916), .S0(n5282), .Y(
        n12378) );
  CLKMX2X2 U11533 ( .A(\I_cache/cache[4][55] ), .B(n9916), .S0(n5325), .Y(
        n12379) );
  CLKMX2X2 U11534 ( .A(\I_cache/cache[3][55] ), .B(n9916), .S0(n5196), .Y(
        n12380) );
  CLKMX2X2 U11535 ( .A(\I_cache/cache[2][55] ), .B(n9916), .S0(n5238), .Y(
        n12381) );
  CLKMX2X2 U11536 ( .A(\I_cache/cache[1][55] ), .B(n9916), .S0(n5109), .Y(
        n12382) );
  CLKMX2X2 U11537 ( .A(\I_cache/cache[0][55] ), .B(n9916), .S0(n5151), .Y(
        n12383) );
  CLKMX2X2 U11538 ( .A(\I_cache/cache[7][54] ), .B(n9848), .S0(n5369), .Y(
        n12384) );
  CLKMX2X2 U11539 ( .A(\I_cache/cache[6][54] ), .B(n9848), .S0(n5413), .Y(
        n12385) );
  CLKMX2X2 U11540 ( .A(\I_cache/cache[5][54] ), .B(n9848), .S0(n5279), .Y(
        n12386) );
  CLKMX2X2 U11541 ( .A(\I_cache/cache[4][54] ), .B(n9848), .S0(n5322), .Y(
        n12387) );
  CLKMX2X2 U11542 ( .A(\I_cache/cache[3][54] ), .B(n9848), .S0(n5193), .Y(
        n12388) );
  CLKMX2X2 U11543 ( .A(\I_cache/cache[2][54] ), .B(n9848), .S0(n5235), .Y(
        n12389) );
  CLKMX2X2 U11544 ( .A(\I_cache/cache[1][54] ), .B(n9848), .S0(n5106), .Y(
        n12390) );
  CLKMX2X2 U11545 ( .A(\I_cache/cache[0][54] ), .B(n9848), .S0(n5148), .Y(
        n12391) );
  CLKMX2X2 U11546 ( .A(\I_cache/cache[7][53] ), .B(n9868), .S0(n5369), .Y(
        n12392) );
  CLKMX2X2 U11547 ( .A(\I_cache/cache[6][53] ), .B(n9868), .S0(n5413), .Y(
        n12393) );
  CLKMX2X2 U11548 ( .A(\I_cache/cache[5][53] ), .B(n9868), .S0(n5279), .Y(
        n12394) );
  CLKMX2X2 U11549 ( .A(\I_cache/cache[4][53] ), .B(n9868), .S0(n5322), .Y(
        n12395) );
  CLKMX2X2 U11550 ( .A(\I_cache/cache[3][53] ), .B(n9868), .S0(n5193), .Y(
        n12396) );
  CLKMX2X2 U11551 ( .A(\I_cache/cache[2][53] ), .B(n9868), .S0(n5235), .Y(
        n12397) );
  CLKMX2X2 U11552 ( .A(\I_cache/cache[1][53] ), .B(n9868), .S0(n5106), .Y(
        n12398) );
  CLKMX2X2 U11553 ( .A(\I_cache/cache[0][53] ), .B(n9868), .S0(n5148), .Y(
        n12399) );
  CLKMX2X2 U11554 ( .A(\I_cache/cache[7][52] ), .B(n10012), .S0(n5371), .Y(
        n12400) );
  CLKMX2X2 U11555 ( .A(\I_cache/cache[6][52] ), .B(n10012), .S0(n5415), .Y(
        n12401) );
  CLKMX2X2 U11556 ( .A(\I_cache/cache[5][52] ), .B(n10012), .S0(n5281), .Y(
        n12402) );
  CLKMX2X2 U11557 ( .A(\I_cache/cache[4][52] ), .B(n10012), .S0(n5324), .Y(
        n12403) );
  CLKMX2X2 U11558 ( .A(\I_cache/cache[3][52] ), .B(n10012), .S0(n5195), .Y(
        n12404) );
  CLKMX2X2 U11559 ( .A(\I_cache/cache[2][52] ), .B(n10012), .S0(n5237), .Y(
        n12405) );
  CLKMX2X2 U11560 ( .A(\I_cache/cache[1][52] ), .B(n10012), .S0(n5108), .Y(
        n12406) );
  CLKMX2X2 U11561 ( .A(\I_cache/cache[0][52] ), .B(n10012), .S0(n5150), .Y(
        n12407) );
  CLKMX2X2 U11562 ( .A(\I_cache/cache[7][51] ), .B(n9983), .S0(n5372), .Y(
        n12408) );
  CLKMX2X2 U11563 ( .A(\I_cache/cache[6][51] ), .B(n9983), .S0(n5416), .Y(
        n12409) );
  CLKMX2X2 U11564 ( .A(\I_cache/cache[5][51] ), .B(n9983), .S0(n5282), .Y(
        n12410) );
  CLKMX2X2 U11565 ( .A(\I_cache/cache[4][51] ), .B(n9983), .S0(n5325), .Y(
        n12411) );
  CLKMX2X2 U11566 ( .A(\I_cache/cache[3][51] ), .B(n9983), .S0(n5196), .Y(
        n12412) );
  CLKMX2X2 U11567 ( .A(\I_cache/cache[2][51] ), .B(n9983), .S0(n5238), .Y(
        n12413) );
  CLKMX2X2 U11568 ( .A(\I_cache/cache[1][51] ), .B(n9983), .S0(n5109), .Y(
        n12414) );
  CLKMX2X2 U11569 ( .A(\I_cache/cache[0][51] ), .B(n9983), .S0(n5151), .Y(
        n12415) );
  CLKMX2X2 U11570 ( .A(\I_cache/cache[6][50] ), .B(n10036), .S0(n5415), .Y(
        n12417) );
  CLKMX2X2 U11571 ( .A(\I_cache/cache[5][50] ), .B(n10036), .S0(n5281), .Y(
        n12418) );
  CLKMX2X2 U11572 ( .A(\I_cache/cache[4][50] ), .B(n10036), .S0(n5324), .Y(
        n12419) );
  CLKMX2X2 U11573 ( .A(\I_cache/cache[2][50] ), .B(n10036), .S0(n5237), .Y(
        n12421) );
  CLKMX2X2 U11574 ( .A(\I_cache/cache[1][50] ), .B(n10036), .S0(n5108), .Y(
        n12422) );
  CLKMX2X2 U11575 ( .A(\I_cache/cache[0][50] ), .B(n10036), .S0(n5150), .Y(
        n12423) );
  CLKMX2X2 U11576 ( .A(\I_cache/cache[7][49] ), .B(n11129), .S0(n5367), .Y(
        n12424) );
  CLKMX2X2 U11577 ( .A(\I_cache/cache[6][49] ), .B(n11129), .S0(n5411), .Y(
        n12425) );
  CLKMX2X2 U11578 ( .A(\I_cache/cache[5][49] ), .B(n11129), .S0(n5278), .Y(
        n12426) );
  CLKMX2X2 U11579 ( .A(\I_cache/cache[4][49] ), .B(n11129), .S0(n5320), .Y(
        n12427) );
  CLKMX2X2 U11580 ( .A(\I_cache/cache[3][49] ), .B(n11129), .S0(n5191), .Y(
        n12428) );
  CLKMX2X2 U11581 ( .A(\I_cache/cache[2][49] ), .B(n11129), .S0(n5233), .Y(
        n12429) );
  CLKMX2X2 U11582 ( .A(\I_cache/cache[1][49] ), .B(n11129), .S0(n5104), .Y(
        n12430) );
  CLKMX2X2 U11583 ( .A(\I_cache/cache[0][49] ), .B(n11129), .S0(n5146), .Y(
        n12431) );
  CLKMX2X2 U11584 ( .A(\I_cache/cache[6][48] ), .B(n10065), .S0(n5415), .Y(
        n12433) );
  CLKMX2X2 U11585 ( .A(\I_cache/cache[5][48] ), .B(n10065), .S0(n5281), .Y(
        n12434) );
  CLKMX2X2 U11586 ( .A(\I_cache/cache[4][48] ), .B(n10065), .S0(n5324), .Y(
        n12435) );
  CLKMX2X2 U11587 ( .A(\I_cache/cache[2][48] ), .B(n10065), .S0(n5237), .Y(
        n12437) );
  CLKMX2X2 U11588 ( .A(\I_cache/cache[1][48] ), .B(n10065), .S0(n5108), .Y(
        n12438) );
  CLKMX2X2 U11589 ( .A(\I_cache/cache[0][48] ), .B(n10065), .S0(n5150), .Y(
        n12439) );
  CLKMX2X2 U11590 ( .A(\I_cache/cache[7][46] ), .B(n9397), .S0(n5368), .Y(
        n12448) );
  CLKMX2X2 U11591 ( .A(\I_cache/cache[6][46] ), .B(n9397), .S0(n5418), .Y(
        n12449) );
  CLKMX2X2 U11592 ( .A(\I_cache/cache[5][46] ), .B(n9397), .S0(n5284), .Y(
        n12450) );
  CLKMX2X2 U11593 ( .A(\I_cache/cache[4][46] ), .B(n9397), .S0(n5327), .Y(
        n12451) );
  CLKMX2X2 U11594 ( .A(\I_cache/cache[3][46] ), .B(n9397), .S0(n5198), .Y(
        n12452) );
  CLKMX2X2 U11595 ( .A(\I_cache/cache[2][46] ), .B(n9397), .S0(n5240), .Y(
        n12453) );
  CLKMX2X2 U11596 ( .A(\I_cache/cache[1][46] ), .B(n9397), .S0(n5110), .Y(
        n12454) );
  CLKMX2X2 U11597 ( .A(\I_cache/cache[0][46] ), .B(n9397), .S0(n5153), .Y(
        n12455) );
  CLKMX2X2 U11598 ( .A(\I_cache/cache[7][45] ), .B(n9377), .S0(n5366), .Y(
        n12456) );
  CLKMX2X2 U11599 ( .A(\I_cache/cache[6][45] ), .B(n9377), .S0(n5418), .Y(
        n12457) );
  CLKMX2X2 U11600 ( .A(\I_cache/cache[5][45] ), .B(n9377), .S0(n5284), .Y(
        n12458) );
  CLKMX2X2 U11601 ( .A(\I_cache/cache[4][45] ), .B(n9377), .S0(n5322), .Y(
        n12459) );
  CLKMX2X2 U11602 ( .A(\I_cache/cache[3][45] ), .B(n9377), .S0(n5198), .Y(
        n12460) );
  CLKMX2X2 U11603 ( .A(\I_cache/cache[2][45] ), .B(n9377), .S0(n5240), .Y(
        n12461) );
  CLKMX2X2 U11604 ( .A(\I_cache/cache[1][45] ), .B(n9377), .S0(n5102), .Y(
        n12462) );
  CLKMX2X2 U11605 ( .A(\I_cache/cache[0][45] ), .B(n9377), .S0(n5153), .Y(
        n12463) );
  CLKMX2X2 U11606 ( .A(\I_cache/cache[7][44] ), .B(n10090), .S0(n5366), .Y(
        n12464) );
  CLKMX2X2 U11607 ( .A(\I_cache/cache[6][44] ), .B(n10090), .S0(n5410), .Y(
        n12465) );
  CLKMX2X2 U11608 ( .A(\I_cache/cache[4][44] ), .B(n10090), .S0(n4679), .Y(
        n12467) );
  CLKMX2X2 U11609 ( .A(\I_cache/cache[3][44] ), .B(n10090), .S0(n5190), .Y(
        n12468) );
  CLKMX2X2 U11610 ( .A(\I_cache/cache[2][44] ), .B(n10090), .S0(n5234), .Y(
        n12469) );
  CLKMX2X2 U11611 ( .A(\I_cache/cache[1][44] ), .B(n10090), .S0(n5103), .Y(
        n12470) );
  CLKMX2X2 U11612 ( .A(\I_cache/cache[0][44] ), .B(n10090), .S0(n5145), .Y(
        n12471) );
  CLKMX2X2 U11613 ( .A(\I_cache/cache[7][43] ), .B(n9959), .S0(n5372), .Y(
        n12472) );
  CLKMX2X2 U11614 ( .A(\I_cache/cache[6][43] ), .B(n9959), .S0(n5416), .Y(
        n12473) );
  CLKMX2X2 U11615 ( .A(\I_cache/cache[5][43] ), .B(n9959), .S0(n5282), .Y(
        n12474) );
  CLKMX2X2 U11616 ( .A(\I_cache/cache[4][43] ), .B(n9959), .S0(n5325), .Y(
        n12475) );
  CLKMX2X2 U11617 ( .A(\I_cache/cache[3][43] ), .B(n9959), .S0(n5196), .Y(
        n12476) );
  CLKMX2X2 U11618 ( .A(\I_cache/cache[2][43] ), .B(n9959), .S0(n5238), .Y(
        n12477) );
  CLKMX2X2 U11619 ( .A(\I_cache/cache[1][43] ), .B(n9959), .S0(n5109), .Y(
        n12478) );
  CLKMX2X2 U11620 ( .A(\I_cache/cache[0][43] ), .B(n9959), .S0(n5151), .Y(
        n12479) );
  CLKMX2X2 U11621 ( .A(\I_cache/cache[7][42] ), .B(n9664), .S0(n5374), .Y(
        n12480) );
  CLKMX2X2 U11622 ( .A(\I_cache/cache[6][42] ), .B(n9664), .S0(n5419), .Y(
        n12481) );
  CLKMX2X2 U11623 ( .A(\I_cache/cache[5][42] ), .B(n9664), .S0(n5283), .Y(
        n12482) );
  CLKMX2X2 U11624 ( .A(\I_cache/cache[4][42] ), .B(n9664), .S0(n5327), .Y(
        n12483) );
  CLKMX2X2 U11625 ( .A(\I_cache/cache[3][42] ), .B(n9664), .S0(n5199), .Y(
        n12484) );
  CLKMX2X2 U11626 ( .A(\I_cache/cache[2][42] ), .B(n9664), .S0(n5241), .Y(
        n12485) );
  CLKMX2X2 U11627 ( .A(\I_cache/cache[1][42] ), .B(n9664), .S0(n5110), .Y(
        n12486) );
  CLKMX2X2 U11628 ( .A(\I_cache/cache[0][42] ), .B(n9664), .S0(n5154), .Y(
        n12487) );
  CLKMX2X2 U11629 ( .A(\I_cache/cache[7][41] ), .B(n9635), .S0(n5368), .Y(
        n12488) );
  CLKMX2X2 U11630 ( .A(\I_cache/cache[5][41] ), .B(n9635), .S0(n5284), .Y(
        n12490) );
  CLKMX2X2 U11631 ( .A(\I_cache/cache[4][41] ), .B(n9635), .S0(n4698), .Y(
        n12491) );
  CLKMX2X2 U11632 ( .A(\I_cache/cache[3][41] ), .B(n9635), .S0(n5198), .Y(
        n12492) );
  CLKMX2X2 U11633 ( .A(\I_cache/cache[2][41] ), .B(n9635), .S0(n5240), .Y(
        n12493) );
  CLKMX2X2 U11634 ( .A(\I_cache/cache[1][41] ), .B(n9635), .S0(n5109), .Y(
        n12494) );
  CLKMX2X2 U11635 ( .A(\I_cache/cache[0][41] ), .B(n9635), .S0(n5153), .Y(
        n12495) );
  CLKMX2X2 U11636 ( .A(\I_cache/cache[7][40] ), .B(n9412), .S0(n3617), .Y(
        n12496) );
  CLKMX2X2 U11637 ( .A(\I_cache/cache[6][40] ), .B(n9412), .S0(n5418), .Y(
        n12497) );
  CLKMX2X2 U11638 ( .A(\I_cache/cache[5][40] ), .B(n9412), .S0(n5284), .Y(
        n12498) );
  CLKMX2X2 U11639 ( .A(\I_cache/cache[4][40] ), .B(n9412), .S0(n4678), .Y(
        n12499) );
  CLKMX2X2 U11640 ( .A(\I_cache/cache[3][40] ), .B(n9412), .S0(n5198), .Y(
        n12500) );
  CLKMX2X2 U11641 ( .A(\I_cache/cache[2][40] ), .B(n9412), .S0(n5240), .Y(
        n12501) );
  CLKMX2X2 U11642 ( .A(\I_cache/cache[1][40] ), .B(n9412), .S0(n5106), .Y(
        n12502) );
  CLKMX2X2 U11643 ( .A(\I_cache/cache[0][40] ), .B(n9412), .S0(n5153), .Y(
        n12503) );
  CLKMX2X2 U11644 ( .A(\I_cache/cache[7][39] ), .B(n9815), .S0(n5370), .Y(
        n12504) );
  CLKMX2X2 U11645 ( .A(\I_cache/cache[6][39] ), .B(n9815), .S0(n5414), .Y(
        n12505) );
  CLKMX2X2 U11646 ( .A(\I_cache/cache[5][39] ), .B(n9815), .S0(n5280), .Y(
        n12506) );
  CLKMX2X2 U11647 ( .A(\I_cache/cache[4][39] ), .B(n9815), .S0(n5323), .Y(
        n12507) );
  CLKMX2X2 U11648 ( .A(\I_cache/cache[3][39] ), .B(n9815), .S0(n5194), .Y(
        n12508) );
  CLKMX2X2 U11649 ( .A(\I_cache/cache[2][39] ), .B(n9815), .S0(n5236), .Y(
        n12509) );
  CLKMX2X2 U11650 ( .A(\I_cache/cache[1][39] ), .B(n9815), .S0(n5107), .Y(
        n12510) );
  CLKMX2X2 U11651 ( .A(\I_cache/cache[0][39] ), .B(n9815), .S0(n5149), .Y(
        n12511) );
  CLKMX2X2 U11652 ( .A(\I_cache/cache[7][38] ), .B(n9446), .S0(n5373), .Y(
        n12512) );
  CLKMX2X2 U11653 ( .A(\I_cache/cache[6][38] ), .B(n9446), .S0(n5417), .Y(
        n12513) );
  CLKMX2X2 U11654 ( .A(\I_cache/cache[5][38] ), .B(n9446), .S0(n5283), .Y(
        n12514) );
  CLKMX2X2 U11655 ( .A(\I_cache/cache[4][38] ), .B(n9446), .S0(n5326), .Y(
        n12515) );
  CLKMX2X2 U11656 ( .A(\I_cache/cache[3][38] ), .B(n9446), .S0(n5197), .Y(
        n12516) );
  CLKMX2X2 U11657 ( .A(\I_cache/cache[2][38] ), .B(n9446), .S0(n5239), .Y(
        n12517) );
  CLKMX2X2 U11658 ( .A(\I_cache/cache[1][38] ), .B(n9446), .S0(n5108), .Y(
        n12518) );
  CLKMX2X2 U11659 ( .A(\I_cache/cache[0][38] ), .B(n9446), .S0(n5152), .Y(
        n12519) );
  CLKMX2X2 U11660 ( .A(\I_cache/cache[7][37] ), .B(n9532), .S0(n5372), .Y(
        n12520) );
  CLKMX2X2 U11661 ( .A(\I_cache/cache[6][37] ), .B(n9532), .S0(n5413), .Y(
        n12521) );
  CLKMX2X2 U11662 ( .A(\I_cache/cache[5][37] ), .B(n9532), .S0(n5285), .Y(
        n12522) );
  CLKMX2X2 U11663 ( .A(\I_cache/cache[4][37] ), .B(n9532), .S0(n5321), .Y(
        n12523) );
  CLKMX2X2 U11664 ( .A(\I_cache/cache[3][37] ), .B(n9532), .S0(n5197), .Y(
        n12524) );
  CLKMX2X2 U11665 ( .A(\I_cache/cache[2][37] ), .B(n9532), .S0(n5242), .Y(
        n12525) );
  CLKMX2X2 U11666 ( .A(\I_cache/cache[1][37] ), .B(n9532), .S0(n5111), .Y(
        n12526) );
  CLKMX2X2 U11667 ( .A(\I_cache/cache[0][37] ), .B(n9532), .S0(n5154), .Y(
        n12527) );
  CLKMX2X2 U11668 ( .A(\I_cache/cache[7][36] ), .B(n9468), .S0(n5373), .Y(
        n12528) );
  CLKMX2X2 U11669 ( .A(\I_cache/cache[6][36] ), .B(n9468), .S0(n5417), .Y(
        n12529) );
  CLKMX2X2 U11670 ( .A(\I_cache/cache[5][36] ), .B(n9468), .S0(n5283), .Y(
        n12530) );
  CLKMX2X2 U11671 ( .A(\I_cache/cache[4][36] ), .B(n9468), .S0(n5326), .Y(
        n12531) );
  CLKMX2X2 U11672 ( .A(\I_cache/cache[3][36] ), .B(n9468), .S0(n5197), .Y(
        n12532) );
  CLKMX2X2 U11673 ( .A(\I_cache/cache[2][36] ), .B(n9468), .S0(n5239), .Y(
        n12533) );
  CLKMX2X2 U11674 ( .A(\I_cache/cache[1][36] ), .B(n9468), .S0(n5107), .Y(
        n12534) );
  CLKMX2X2 U11675 ( .A(\I_cache/cache[0][36] ), .B(n9468), .S0(n5152), .Y(
        n12535) );
  CLKMX2X2 U11676 ( .A(\I_cache/cache[6][31] ), .B(n11035), .S0(n5412), .Y(
        n12569) );
  CLKMX2X2 U11677 ( .A(\I_cache/cache[4][31] ), .B(n11035), .S0(n5321), .Y(
        n12571) );
  CLKMX2X2 U11678 ( .A(\I_cache/cache[3][31] ), .B(n11035), .S0(n5192), .Y(
        n12572) );
  CLKMX2X2 U11679 ( .A(\I_cache/cache[2][31] ), .B(n11035), .S0(n5234), .Y(
        n12573) );
  CLKMX2X2 U11680 ( .A(\I_cache/cache[1][31] ), .B(n11035), .S0(n5105), .Y(
        n12574) );
  CLKMX2X2 U11681 ( .A(\I_cache/cache[0][31] ), .B(n11035), .S0(n5147), .Y(
        n12575) );
  CLKMX2X2 U11682 ( .A(\I_cache/cache[7][30] ), .B(n9788), .S0(n5370), .Y(
        n12576) );
  CLKMX2X2 U11683 ( .A(\I_cache/cache[6][30] ), .B(n9788), .S0(n5414), .Y(
        n12577) );
  CLKMX2X2 U11684 ( .A(\I_cache/cache[5][30] ), .B(n9788), .S0(n5280), .Y(
        n12578) );
  CLKMX2X2 U11685 ( .A(\I_cache/cache[4][30] ), .B(n9788), .S0(n5323), .Y(
        n12579) );
  CLKMX2X2 U11686 ( .A(\I_cache/cache[3][30] ), .B(n9788), .S0(n5194), .Y(
        n12580) );
  CLKMX2X2 U11687 ( .A(\I_cache/cache[2][30] ), .B(n9788), .S0(n5236), .Y(
        n12581) );
  CLKMX2X2 U11688 ( .A(\I_cache/cache[1][30] ), .B(n9788), .S0(n5107), .Y(
        n12582) );
  CLKMX2X2 U11689 ( .A(\I_cache/cache[0][30] ), .B(n9788), .S0(n5149), .Y(
        n12583) );
  CLKMX2X2 U11690 ( .A(\I_cache/cache[7][29] ), .B(n11158), .S0(n5367), .Y(
        n12584) );
  CLKMX2X2 U11691 ( .A(\I_cache/cache[6][29] ), .B(n11158), .S0(n5411), .Y(
        n12585) );
  CLKMX2X2 U11692 ( .A(\I_cache/cache[5][29] ), .B(n11158), .S0(n5278), .Y(
        n12586) );
  CLKMX2X2 U11693 ( .A(\I_cache/cache[4][29] ), .B(n11158), .S0(n5320), .Y(
        n12587) );
  CLKMX2X2 U11694 ( .A(\I_cache/cache[3][29] ), .B(n11158), .S0(n5191), .Y(
        n12588) );
  CLKMX2X2 U11695 ( .A(\I_cache/cache[2][29] ), .B(n11158), .S0(n5233), .Y(
        n12589) );
  CLKMX2X2 U11696 ( .A(\I_cache/cache[1][29] ), .B(n11158), .S0(n5104), .Y(
        n12590) );
  CLKMX2X2 U11697 ( .A(\I_cache/cache[0][29] ), .B(n11158), .S0(n5146), .Y(
        n12591) );
  CLKMX2X2 U11698 ( .A(\I_cache/cache[7][28] ), .B(n9764), .S0(n5370), .Y(
        n12592) );
  CLKMX2X2 U11699 ( .A(\I_cache/cache[6][28] ), .B(n9764), .S0(n5414), .Y(
        n12593) );
  CLKMX2X2 U11700 ( .A(\I_cache/cache[5][28] ), .B(n9764), .S0(n5280), .Y(
        n12594) );
  CLKMX2X2 U11701 ( .A(\I_cache/cache[4][28] ), .B(n9764), .S0(n5323), .Y(
        n12595) );
  CLKMX2X2 U11702 ( .A(\I_cache/cache[3][28] ), .B(n9764), .S0(n5194), .Y(
        n12596) );
  CLKMX2X2 U11703 ( .A(\I_cache/cache[2][28] ), .B(n9764), .S0(n5236), .Y(
        n12597) );
  CLKMX2X2 U11704 ( .A(\I_cache/cache[1][28] ), .B(n9764), .S0(n5107), .Y(
        n12598) );
  CLKMX2X2 U11705 ( .A(\I_cache/cache[0][28] ), .B(n9764), .S0(n5149), .Y(
        n12599) );
  CLKMX2X2 U11706 ( .A(\I_cache/cache[7][27] ), .B(n9720), .S0(n5369), .Y(
        n12600) );
  CLKMX2X2 U11707 ( .A(\I_cache/cache[6][27] ), .B(n9720), .S0(n5413), .Y(
        n12601) );
  CLKMX2X2 U11708 ( .A(\I_cache/cache[5][27] ), .B(n9720), .S0(n5279), .Y(
        n12602) );
  CLKMX2X2 U11709 ( .A(\I_cache/cache[4][27] ), .B(n9720), .S0(n5322), .Y(
        n12603) );
  CLKMX2X2 U11710 ( .A(\I_cache/cache[3][27] ), .B(n9720), .S0(n5193), .Y(
        n12604) );
  CLKMX2X2 U11711 ( .A(\I_cache/cache[2][27] ), .B(n9720), .S0(n5235), .Y(
        n12605) );
  CLKMX2X2 U11712 ( .A(\I_cache/cache[1][27] ), .B(n9720), .S0(n5106), .Y(
        n12606) );
  CLKMX2X2 U11713 ( .A(\I_cache/cache[0][27] ), .B(n9720), .S0(n5148), .Y(
        n12607) );
  CLKMX2X2 U11714 ( .A(\I_cache/cache[7][26] ), .B(n9696), .S0(n5374), .Y(
        n12608) );
  CLKMX2X2 U11715 ( .A(\I_cache/cache[6][26] ), .B(n9696), .S0(n5419), .Y(
        n12609) );
  CLKMX2X2 U11716 ( .A(\I_cache/cache[5][26] ), .B(n9696), .S0(n5281), .Y(
        n12610) );
  CLKMX2X2 U11717 ( .A(\I_cache/cache[4][26] ), .B(n9696), .S0(n5327), .Y(
        n12611) );
  CLKMX2X2 U11718 ( .A(\I_cache/cache[3][26] ), .B(n9696), .S0(n5199), .Y(
        n12612) );
  CLKMX2X2 U11719 ( .A(\I_cache/cache[2][26] ), .B(n9696), .S0(n5241), .Y(
        n12613) );
  CLKMX2X2 U11720 ( .A(\I_cache/cache[1][26] ), .B(n9696), .S0(n5110), .Y(
        n12614) );
  CLKMX2X2 U11721 ( .A(\I_cache/cache[0][26] ), .B(n9696), .S0(n5154), .Y(
        n12615) );
  CLKMX2X2 U11722 ( .A(\I_cache/cache[7][25] ), .B(n10109), .S0(n5366), .Y(
        n12616) );
  CLKMX2X2 U11723 ( .A(\I_cache/cache[6][25] ), .B(n10109), .S0(n5410), .Y(
        n12617) );
  CLKMX2X2 U11724 ( .A(\I_cache/cache[4][25] ), .B(n10109), .S0(n4680), .Y(
        n12619) );
  CLKMX2X2 U11725 ( .A(\I_cache/cache[3][25] ), .B(n10109), .S0(n5190), .Y(
        n12620) );
  CLKMX2X2 U11726 ( .A(\I_cache/cache[2][25] ), .B(n10109), .S0(n5238), .Y(
        n12621) );
  CLKMX2X2 U11727 ( .A(\I_cache/cache[1][25] ), .B(n10109), .S0(n5103), .Y(
        n12622) );
  CLKMX2X2 U11728 ( .A(\I_cache/cache[0][25] ), .B(n10109), .S0(n5145), .Y(
        n12623) );
  CLKMX2X2 U11729 ( .A(\I_cache/cache[7][24] ), .B(n9887), .S0(n5369), .Y(
        n12624) );
  CLKMX2X2 U11730 ( .A(\I_cache/cache[6][24] ), .B(n9887), .S0(n5413), .Y(
        n12625) );
  CLKMX2X2 U11731 ( .A(\I_cache/cache[5][24] ), .B(n9887), .S0(n5279), .Y(
        n12626) );
  CLKMX2X2 U11732 ( .A(\I_cache/cache[4][24] ), .B(n9887), .S0(n5322), .Y(
        n12627) );
  CLKMX2X2 U11733 ( .A(\I_cache/cache[3][24] ), .B(n9887), .S0(n5193), .Y(
        n12628) );
  CLKMX2X2 U11734 ( .A(\I_cache/cache[2][24] ), .B(n9887), .S0(n5235), .Y(
        n12629) );
  CLKMX2X2 U11735 ( .A(\I_cache/cache[1][24] ), .B(n9887), .S0(n5106), .Y(
        n12630) );
  CLKMX2X2 U11736 ( .A(\I_cache/cache[0][24] ), .B(n9887), .S0(n5148), .Y(
        n12631) );
  CLKMX2X2 U11737 ( .A(\I_cache/cache[7][23] ), .B(n9911), .S0(n5372), .Y(
        n12632) );
  CLKMX2X2 U11738 ( .A(\I_cache/cache[6][23] ), .B(n9911), .S0(n5416), .Y(
        n12633) );
  CLKMX2X2 U11739 ( .A(\I_cache/cache[5][23] ), .B(n9911), .S0(n5282), .Y(
        n12634) );
  CLKMX2X2 U11740 ( .A(\I_cache/cache[4][23] ), .B(n9911), .S0(n5325), .Y(
        n12635) );
  CLKMX2X2 U11741 ( .A(\I_cache/cache[3][23] ), .B(n9911), .S0(n5196), .Y(
        n12636) );
  CLKMX2X2 U11742 ( .A(\I_cache/cache[2][23] ), .B(n9911), .S0(n5238), .Y(
        n12637) );
  CLKMX2X2 U11743 ( .A(\I_cache/cache[1][23] ), .B(n9911), .S0(n5109), .Y(
        n12638) );
  CLKMX2X2 U11744 ( .A(\I_cache/cache[0][23] ), .B(n9911), .S0(n5151), .Y(
        n12639) );
  CLKMX2X2 U11745 ( .A(\I_cache/cache[7][22] ), .B(n9843), .S0(n5369), .Y(
        n12640) );
  CLKMX2X2 U11746 ( .A(\I_cache/cache[6][22] ), .B(n9843), .S0(n5413), .Y(
        n12641) );
  CLKMX2X2 U11747 ( .A(\I_cache/cache[5][22] ), .B(n9843), .S0(n5279), .Y(
        n12642) );
  CLKMX2X2 U11748 ( .A(\I_cache/cache[4][22] ), .B(n9843), .S0(n5322), .Y(
        n12643) );
  CLKMX2X2 U11749 ( .A(\I_cache/cache[3][22] ), .B(n9843), .S0(n5193), .Y(
        n12644) );
  CLKMX2X2 U11750 ( .A(\I_cache/cache[2][22] ), .B(n9843), .S0(n5235), .Y(
        n12645) );
  CLKMX2X2 U11751 ( .A(\I_cache/cache[1][22] ), .B(n9843), .S0(n5106), .Y(
        n12646) );
  CLKMX2X2 U11752 ( .A(\I_cache/cache[0][22] ), .B(n9843), .S0(n5148), .Y(
        n12647) );
  CLKMX2X2 U11753 ( .A(\I_cache/cache[7][21] ), .B(n9863), .S0(n5369), .Y(
        n12648) );
  CLKMX2X2 U11754 ( .A(\I_cache/cache[6][21] ), .B(n9863), .S0(n5413), .Y(
        n12649) );
  CLKMX2X2 U11755 ( .A(\I_cache/cache[5][21] ), .B(n9863), .S0(n5279), .Y(
        n12650) );
  CLKMX2X2 U11756 ( .A(\I_cache/cache[4][21] ), .B(n9863), .S0(n5322), .Y(
        n12651) );
  CLKMX2X2 U11757 ( .A(\I_cache/cache[3][21] ), .B(n9863), .S0(n5193), .Y(
        n12652) );
  CLKMX2X2 U11758 ( .A(\I_cache/cache[2][21] ), .B(n9863), .S0(n5235), .Y(
        n12653) );
  CLKMX2X2 U11759 ( .A(\I_cache/cache[1][21] ), .B(n9863), .S0(n5106), .Y(
        n12654) );
  CLKMX2X2 U11760 ( .A(\I_cache/cache[0][21] ), .B(n9863), .S0(n5148), .Y(
        n12655) );
  CLKMX2X2 U11761 ( .A(\I_cache/cache[7][20] ), .B(n10007), .S0(n5371), .Y(
        n12656) );
  CLKMX2X2 U11762 ( .A(\I_cache/cache[6][20] ), .B(n10007), .S0(n5415), .Y(
        n12657) );
  CLKMX2X2 U11763 ( .A(\I_cache/cache[5][20] ), .B(n10007), .S0(n5281), .Y(
        n12658) );
  CLKMX2X2 U11764 ( .A(\I_cache/cache[4][20] ), .B(n10007), .S0(n5324), .Y(
        n12659) );
  CLKMX2X2 U11765 ( .A(\I_cache/cache[3][20] ), .B(n10007), .S0(n5195), .Y(
        n12660) );
  CLKMX2X2 U11766 ( .A(\I_cache/cache[2][20] ), .B(n10007), .S0(n5237), .Y(
        n12661) );
  CLKMX2X2 U11767 ( .A(\I_cache/cache[1][20] ), .B(n10007), .S0(n5108), .Y(
        n12662) );
  CLKMX2X2 U11768 ( .A(\I_cache/cache[0][20] ), .B(n10007), .S0(n5150), .Y(
        n12663) );
  CLKMX2X2 U11769 ( .A(\I_cache/cache[7][19] ), .B(n9978), .S0(n5372), .Y(
        n12664) );
  CLKMX2X2 U11770 ( .A(\I_cache/cache[6][19] ), .B(n9978), .S0(n5416), .Y(
        n12665) );
  CLKMX2X2 U11771 ( .A(\I_cache/cache[5][19] ), .B(n9978), .S0(n5282), .Y(
        n12666) );
  CLKMX2X2 U11772 ( .A(\I_cache/cache[4][19] ), .B(n9978), .S0(n5325), .Y(
        n12667) );
  CLKMX2X2 U11773 ( .A(\I_cache/cache[3][19] ), .B(n9978), .S0(n5196), .Y(
        n12668) );
  CLKMX2X2 U11774 ( .A(\I_cache/cache[2][19] ), .B(n9978), .S0(n5238), .Y(
        n12669) );
  CLKMX2X2 U11775 ( .A(\I_cache/cache[1][19] ), .B(n9978), .S0(n5109), .Y(
        n12670) );
  CLKMX2X2 U11776 ( .A(\I_cache/cache[0][19] ), .B(n9978), .S0(n5151), .Y(
        n12671) );
  CLKMX2X2 U11777 ( .A(\I_cache/cache[7][18] ), .B(n10031), .S0(n5371), .Y(
        n12672) );
  CLKMX2X2 U11778 ( .A(\I_cache/cache[6][18] ), .B(n10031), .S0(n5415), .Y(
        n12673) );
  CLKMX2X2 U11779 ( .A(\I_cache/cache[5][18] ), .B(n10031), .S0(n5281), .Y(
        n12674) );
  CLKMX2X2 U11780 ( .A(\I_cache/cache[4][18] ), .B(n10031), .S0(n5324), .Y(
        n12675) );
  CLKMX2X2 U11781 ( .A(\I_cache/cache[3][18] ), .B(n10031), .S0(n5195), .Y(
        n12676) );
  CLKMX2X2 U11782 ( .A(\I_cache/cache[2][18] ), .B(n10031), .S0(n5237), .Y(
        n12677) );
  CLKMX2X2 U11783 ( .A(\I_cache/cache[1][18] ), .B(n10031), .S0(n5108), .Y(
        n12678) );
  CLKMX2X2 U11784 ( .A(\I_cache/cache[0][18] ), .B(n10031), .S0(n5150), .Y(
        n12679) );
  CLKMX2X2 U11785 ( .A(\I_cache/cache[7][17] ), .B(n11124), .S0(n5367), .Y(
        n12680) );
  CLKMX2X2 U11786 ( .A(\I_cache/cache[6][17] ), .B(n11124), .S0(n5411), .Y(
        n12681) );
  CLKMX2X2 U11787 ( .A(\I_cache/cache[5][17] ), .B(n11124), .S0(n5278), .Y(
        n12682) );
  CLKMX2X2 U11788 ( .A(\I_cache/cache[4][17] ), .B(n11124), .S0(n5320), .Y(
        n12683) );
  CLKMX2X2 U11789 ( .A(\I_cache/cache[3][17] ), .B(n11124), .S0(n5191), .Y(
        n12684) );
  CLKMX2X2 U11790 ( .A(\I_cache/cache[2][17] ), .B(n11124), .S0(n5233), .Y(
        n12685) );
  CLKMX2X2 U11791 ( .A(\I_cache/cache[1][17] ), .B(n11124), .S0(n5104), .Y(
        n12686) );
  CLKMX2X2 U11792 ( .A(\I_cache/cache[0][17] ), .B(n11124), .S0(n5146), .Y(
        n12687) );
  CLKMX2X2 U11793 ( .A(\I_cache/cache[7][16] ), .B(n10060), .S0(n5371), .Y(
        n12688) );
  CLKMX2X2 U11794 ( .A(\I_cache/cache[6][16] ), .B(n10060), .S0(n5415), .Y(
        n12689) );
  CLKMX2X2 U11795 ( .A(\I_cache/cache[5][16] ), .B(n10060), .S0(n5281), .Y(
        n12690) );
  CLKMX2X2 U11796 ( .A(\I_cache/cache[2][16] ), .B(n10060), .S0(n5237), .Y(
        n12693) );
  CLKMX2X2 U11797 ( .A(\I_cache/cache[1][16] ), .B(n10060), .S0(n5108), .Y(
        n12694) );
  CLKMX2X2 U11798 ( .A(\I_cache/cache[0][16] ), .B(n10060), .S0(n5150), .Y(
        n12695) );
  CLKMX2X2 U11799 ( .A(\I_cache/cache[3][6] ), .B(n9436), .S0(n5197), .Y(
        n12772) );
  CLKMX2X2 U11800 ( .A(\I_cache/cache[1][6] ), .B(n9436), .S0(n5103), .Y(
        n12774) );
  CLKMX2X2 U11801 ( .A(\I_cache/cache[4][1] ), .B(n9356), .S0(n4677), .Y(
        n12811) );
  MX2XL U11802 ( .A(\I_cache/cache[6][152] ), .B(n10977), .S0(n5410), .Y(
        n11601) );
  MX2XL U11803 ( .A(\I_cache/cache[5][152] ), .B(n10977), .S0(n5277), .Y(
        n11602) );
  MX2XL U11804 ( .A(\I_cache/cache[4][152] ), .B(n10977), .S0(n4698), .Y(
        n11603) );
  MX2XL U11805 ( .A(\I_cache/cache[3][152] ), .B(n10977), .S0(n5190), .Y(
        n11604) );
  MX2XL U11806 ( .A(\I_cache/cache[2][152] ), .B(n10977), .S0(n5234), .Y(
        n11605) );
  MX2XL U11807 ( .A(\I_cache/cache[1][152] ), .B(n10977), .S0(n5103), .Y(
        n11606) );
  MX2XL U11808 ( .A(\I_cache/cache[0][152] ), .B(n10977), .S0(n5145), .Y(
        n11607) );
  MX2XL U11809 ( .A(\I_cache/cache[5][151] ), .B(n3512), .S0(n5277), .Y(n11610) );
  MX2XL U11810 ( .A(\I_cache/cache[4][151] ), .B(n3512), .S0(n4679), .Y(n11611) );
  MX2XL U11811 ( .A(\I_cache/cache[2][151] ), .B(n3512), .S0(n5240), .Y(n11613) );
  MX2XL U11812 ( .A(\I_cache/cache[0][151] ), .B(n3512), .S0(n5145), .Y(n11615) );
  MX2XL U11813 ( .A(\I_cache/cache[5][150] ), .B(n10991), .S0(n5278), .Y(
        n11618) );
  MX2XL U11814 ( .A(\I_cache/cache[4][150] ), .B(n10991), .S0(n5323), .Y(
        n11619) );
  MX2XL U11815 ( .A(\I_cache/cache[6][149] ), .B(n10985), .S0(n5412), .Y(
        n11625) );
  MX2XL U11816 ( .A(\I_cache/cache[5][149] ), .B(n10985), .S0(n5280), .Y(
        n11626) );
  MX2XL U11817 ( .A(\I_cache/cache[4][149] ), .B(n10985), .S0(n5321), .Y(
        n11627) );
  MX2XL U11818 ( .A(\I_cache/cache[3][149] ), .B(n10985), .S0(n5190), .Y(
        n11628) );
  MX2XL U11819 ( .A(\I_cache/cache[2][149] ), .B(n10985), .S0(n5241), .Y(
        n11629) );
  MX2XL U11820 ( .A(\I_cache/cache[1][149] ), .B(n10985), .S0(n5102), .Y(
        n11630) );
  MX2XL U11821 ( .A(\I_cache/cache[0][149] ), .B(n10985), .S0(n5145), .Y(
        n11631) );
  MX2XL U11822 ( .A(\I_cache/cache[5][148] ), .B(n10983), .S0(n5277), .Y(
        n11634) );
  MX2XL U11823 ( .A(\I_cache/cache[4][148] ), .B(n10983), .S0(n4679), .Y(
        n11635) );
  MX2XL U11824 ( .A(\I_cache/cache[7][147] ), .B(n10984), .S0(n5373), .Y(
        n11640) );
  MX2XL U11825 ( .A(\I_cache/cache[6][147] ), .B(n10984), .S0(n5411), .Y(
        n11641) );
  MX2XL U11826 ( .A(\I_cache/cache[5][147] ), .B(n10984), .S0(n5278), .Y(
        n11642) );
  MX2XL U11827 ( .A(\I_cache/cache[4][147] ), .B(n10984), .S0(n5320), .Y(
        n11643) );
  MX2XL U11828 ( .A(\I_cache/cache[3][147] ), .B(n10984), .S0(n5197), .Y(
        n11644) );
  MX2XL U11829 ( .A(\I_cache/cache[2][147] ), .B(n10984), .S0(n5239), .Y(
        n11645) );
  MX2XL U11830 ( .A(\I_cache/cache[1][147] ), .B(n10984), .S0(n5102), .Y(
        n11646) );
  MX2XL U11831 ( .A(\I_cache/cache[0][147] ), .B(n10984), .S0(n5151), .Y(
        n11647) );
  MX2XL U11832 ( .A(\I_cache/cache[5][146] ), .B(n10992), .S0(n5280), .Y(
        n11650) );
  MX2XL U11833 ( .A(\I_cache/cache[4][146] ), .B(n10992), .S0(n5323), .Y(
        n11651) );
  MX2XL U11834 ( .A(\I_cache/cache[1][145] ), .B(n10990), .S0(n5102), .Y(
        n11662) );
  MX2XL U11835 ( .A(\I_cache/cache[0][145] ), .B(n10990), .S0(n5153), .Y(
        n11663) );
  MX2XL U11836 ( .A(\I_cache/cache[5][144] ), .B(n3514), .S0(n5277), .Y(n11666) );
  MX2XL U11837 ( .A(\I_cache/cache[4][144] ), .B(n3514), .S0(n4678), .Y(n11667) );
  MX2XL U11838 ( .A(\I_cache/cache[6][143] ), .B(n10996), .S0(n5412), .Y(
        n11673) );
  MX2XL U11839 ( .A(\I_cache/cache[5][143] ), .B(n10996), .S0(n5285), .Y(
        n11674) );
  MX2XL U11840 ( .A(\I_cache/cache[4][143] ), .B(n10996), .S0(n5321), .Y(
        n11675) );
  MX2XL U11841 ( .A(\I_cache/cache[3][143] ), .B(n10996), .S0(n5192), .Y(
        n11676) );
  MX2XL U11842 ( .A(\I_cache/cache[2][143] ), .B(n10996), .S0(n5234), .Y(
        n11677) );
  MX2XL U11843 ( .A(\I_cache/cache[1][143] ), .B(n10996), .S0(n5105), .Y(
        n11678) );
  MX2XL U11844 ( .A(\I_cache/cache[4][142] ), .B(n11034), .S0(n5321), .Y(
        n11683) );
  MX2XL U11845 ( .A(\I_cache/cache[3][142] ), .B(n11034), .S0(n5192), .Y(
        n11684) );
  MX2XL U11846 ( .A(\I_cache/cache[1][142] ), .B(n11034), .S0(n5105), .Y(
        n11686) );
  MX2XL U11847 ( .A(\I_cache/cache[6][140] ), .B(n11157), .S0(n5411), .Y(
        n11697) );
  MX2XL U11848 ( .A(\I_cache/cache[5][140] ), .B(n11157), .S0(n5278), .Y(
        n11698) );
  MX2XL U11849 ( .A(\I_cache/cache[4][140] ), .B(n11157), .S0(n5320), .Y(
        n11699) );
  MX2XL U11850 ( .A(\I_cache/cache[3][140] ), .B(n11157), .S0(n5191), .Y(
        n11700) );
  MX2XL U11851 ( .A(\I_cache/cache[1][140] ), .B(n11157), .S0(n5104), .Y(
        n11702) );
  CLKMX2X2 U11852 ( .A(\I_cache/cache[4][104] ), .B(n9426), .S0(n5326), .Y(
        n11987) );
  MX2XL U11853 ( .A(\I_cache/cache[7][141] ), .B(n10997), .S0(n5368), .Y(
        n11688) );
  MX2XL U11854 ( .A(\I_cache/cache[6][141] ), .B(n10997), .S0(n5412), .Y(
        n11689) );
  MX2XL U11855 ( .A(\I_cache/cache[5][141] ), .B(n10997), .S0(n5280), .Y(
        n11690) );
  MX2XL U11856 ( .A(\I_cache/cache[4][141] ), .B(n10997), .S0(n5321), .Y(
        n11691) );
  MX2XL U11857 ( .A(\I_cache/cache[3][141] ), .B(n10997), .S0(n5192), .Y(
        n11692) );
  MX2XL U11858 ( .A(\I_cache/cache[1][141] ), .B(n10997), .S0(n5105), .Y(
        n11694) );
  MX2XL U11859 ( .A(\I_cache/cache[5][139] ), .B(n10976), .S0(n5277), .Y(
        n11706) );
  MX2XL U11860 ( .A(\I_cache/cache[0][139] ), .B(n10976), .S0(n5145), .Y(
        n11711) );
  MX2XL U11861 ( .A(\I_cache/cache[5][138] ), .B(n10989), .S0(n5277), .Y(
        n11714) );
  MX2XL U11862 ( .A(\I_cache/cache[5][137] ), .B(n3510), .S0(n4675), .Y(n11722) );
  MX2XL U11863 ( .A(\I_cache/cache[4][137] ), .B(n3510), .S0(n5321), .Y(n11723) );
  MX2XL U11864 ( .A(\I_cache/cache[6][136] ), .B(n10980), .S0(n5414), .Y(
        n11729) );
  MX2XL U11865 ( .A(\I_cache/cache[5][136] ), .B(n10980), .S0(n5280), .Y(
        n11730) );
  MX2XL U11866 ( .A(\I_cache/cache[4][136] ), .B(n10980), .S0(n5323), .Y(
        n11731) );
  MX2XL U11867 ( .A(\I_cache/cache[3][136] ), .B(n10980), .S0(n5194), .Y(
        n11732) );
  MX2XL U11868 ( .A(\I_cache/cache[2][136] ), .B(n10980), .S0(n5236), .Y(
        n11733) );
  MX2XL U11869 ( .A(\I_cache/cache[1][136] ), .B(n10980), .S0(n5107), .Y(
        n11734) );
  MX2XL U11870 ( .A(\I_cache/cache[6][135] ), .B(n10981), .S0(n5415), .Y(
        n11737) );
  MX2XL U11871 ( .A(\I_cache/cache[5][135] ), .B(n10981), .S0(n4675), .Y(
        n11738) );
  MX2XL U11872 ( .A(\I_cache/cache[4][135] ), .B(n10981), .S0(n4678), .Y(
        n11739) );
  MX2XL U11873 ( .A(\I_cache/cache[3][135] ), .B(n10981), .S0(n5198), .Y(
        n11740) );
  MX2XL U11874 ( .A(\I_cache/cache[1][135] ), .B(n10981), .S0(n5102), .Y(
        n11742) );
  MX2XL U11875 ( .A(\I_cache/cache[5][134] ), .B(n10987), .S0(n4675), .Y(
        n11746) );
  MX2XL U11876 ( .A(\I_cache/cache[4][134] ), .B(n10987), .S0(n5320), .Y(
        n11747) );
  MX2XL U11877 ( .A(\I_cache/cache[5][133] ), .B(n10988), .S0(n4675), .Y(
        n11754) );
  MX2XL U11878 ( .A(\I_cache/cache[4][133] ), .B(n10988), .S0(n5323), .Y(
        n11755) );
  MX2XL U11879 ( .A(\I_cache/cache[5][131] ), .B(n10994), .S0(n5278), .Y(
        n11770) );
  MX2XL U11880 ( .A(\I_cache/cache[4][131] ), .B(n10994), .S0(n5320), .Y(
        n11771) );
  MX2XL U11881 ( .A(\I_cache/cache[5][130] ), .B(n10993), .S0(n5278), .Y(
        n11778) );
  MX2XL U11882 ( .A(\I_cache/cache[4][130] ), .B(n10993), .S0(n5320), .Y(
        n11779) );
  MX2XL U11883 ( .A(\I_cache/cache[6][129] ), .B(n10995), .S0(n5412), .Y(
        n11785) );
  MX2XL U11884 ( .A(\I_cache/cache[3][129] ), .B(n10995), .S0(n5192), .Y(
        n11788) );
  MX2XL U11885 ( .A(\I_cache/cache[2][129] ), .B(n10995), .S0(n5234), .Y(
        n11789) );
  MX2XL U11886 ( .A(\I_cache/cache[1][129] ), .B(n10995), .S0(n5105), .Y(
        n11790) );
  MX2XL U11887 ( .A(\I_cache/cache[0][129] ), .B(n10995), .S0(n5147), .Y(
        n11791) );
  CLKMX2X2 U11888 ( .A(\I_cache/cache[7][35] ), .B(n9522), .S0(n5369), .Y(
        n12536) );
  CLKMX2X2 U11889 ( .A(\I_cache/cache[6][35] ), .B(n9522), .S0(n5416), .Y(
        n12537) );
  CLKMX2X2 U11890 ( .A(\I_cache/cache[5][35] ), .B(n9522), .S0(n5285), .Y(
        n12538) );
  CLKMX2X2 U11891 ( .A(\I_cache/cache[4][35] ), .B(n9522), .S0(n5324), .Y(
        n12539) );
  CLKMX2X2 U11892 ( .A(\I_cache/cache[3][35] ), .B(n9522), .S0(n5199), .Y(
        n12540) );
  CLKMX2X2 U11893 ( .A(\I_cache/cache[2][35] ), .B(n9522), .S0(n5242), .Y(
        n12541) );
  CLKMX2X2 U11894 ( .A(\I_cache/cache[1][35] ), .B(n9522), .S0(n5111), .Y(
        n12542) );
  CLKMX2X2 U11895 ( .A(\I_cache/cache[0][35] ), .B(n9522), .S0(n5152), .Y(
        n12543) );
  CLKMX2X2 U11896 ( .A(\I_cache/cache[7][34] ), .B(n9487), .S0(n5374), .Y(
        n12544) );
  CLKMX2X2 U11897 ( .A(\I_cache/cache[6][34] ), .B(n9487), .S0(n5419), .Y(
        n12545) );
  CLKMX2X2 U11898 ( .A(\I_cache/cache[5][34] ), .B(n9487), .S0(n5285), .Y(
        n12546) );
  CLKMX2X2 U11899 ( .A(\I_cache/cache[4][34] ), .B(n9487), .S0(n5327), .Y(
        n12547) );
  CLKMX2X2 U11900 ( .A(\I_cache/cache[3][34] ), .B(n9487), .S0(n5199), .Y(
        n12548) );
  CLKMX2X2 U11901 ( .A(\I_cache/cache[2][34] ), .B(n9487), .S0(n5241), .Y(
        n12549) );
  CLKMX2X2 U11902 ( .A(\I_cache/cache[1][34] ), .B(n9487), .S0(n5110), .Y(
        n12550) );
  CLKMX2X2 U11903 ( .A(\I_cache/cache[0][34] ), .B(n9487), .S0(n5154), .Y(
        n12551) );
  CLKMX2X2 U11904 ( .A(\I_cache/cache[7][33] ), .B(n10998), .S0(n5368), .Y(
        n12552) );
  CLKMX2X2 U11905 ( .A(\I_cache/cache[6][33] ), .B(n10998), .S0(n5412), .Y(
        n12553) );
  CLKMX2X2 U11906 ( .A(\I_cache/cache[5][33] ), .B(n10998), .S0(n5280), .Y(
        n12554) );
  CLKMX2X2 U11907 ( .A(\I_cache/cache[4][33] ), .B(n10998), .S0(n5321), .Y(
        n12555) );
  CLKMX2X2 U11908 ( .A(\I_cache/cache[3][33] ), .B(n10998), .S0(n5192), .Y(
        n12556) );
  CLKMX2X2 U11909 ( .A(\I_cache/cache[2][33] ), .B(n10998), .S0(n5234), .Y(
        n12557) );
  CLKMX2X2 U11910 ( .A(\I_cache/cache[1][33] ), .B(n10998), .S0(n5105), .Y(
        n12558) );
  CLKMX2X2 U11911 ( .A(\I_cache/cache[0][33] ), .B(n10998), .S0(n5147), .Y(
        n12559) );
  CLKMX2X2 U11912 ( .A(\I_cache/cache[7][32] ), .B(n9502), .S0(n5374), .Y(
        n12560) );
  CLKMX2X2 U11913 ( .A(\I_cache/cache[6][32] ), .B(n9502), .S0(n5417), .Y(
        n12561) );
  CLKMX2X2 U11914 ( .A(\I_cache/cache[5][32] ), .B(n9502), .S0(n5285), .Y(
        n12562) );
  CLKMX2X2 U11915 ( .A(\I_cache/cache[4][32] ), .B(n9502), .S0(n4680), .Y(
        n12563) );
  CLKMX2X2 U11916 ( .A(\I_cache/cache[3][32] ), .B(n9502), .S0(n5196), .Y(
        n12564) );
  CLKMX2X2 U11917 ( .A(\I_cache/cache[2][32] ), .B(n9502), .S0(n5242), .Y(
        n12565) );
  CLKMX2X2 U11918 ( .A(\I_cache/cache[1][32] ), .B(n9502), .S0(n5111), .Y(
        n12566) );
  CLKMX2X2 U11919 ( .A(\I_cache/cache[0][32] ), .B(n9502), .S0(n5151), .Y(
        n12567) );
  CLKMX2X2 U11920 ( .A(\I_cache/cache[7][14] ), .B(n9392), .S0(n3617), .Y(
        n12704) );
  CLKMX2X2 U11921 ( .A(\I_cache/cache[6][14] ), .B(n9392), .S0(n5418), .Y(
        n12705) );
  CLKMX2X2 U11922 ( .A(\I_cache/cache[5][14] ), .B(n9392), .S0(n5284), .Y(
        n12706) );
  CLKMX2X2 U11923 ( .A(\I_cache/cache[4][14] ), .B(n9392), .S0(n4680), .Y(
        n12707) );
  CLKMX2X2 U11924 ( .A(\I_cache/cache[3][14] ), .B(n9392), .S0(n5198), .Y(
        n12708) );
  CLKMX2X2 U11925 ( .A(\I_cache/cache[2][14] ), .B(n9392), .S0(n5240), .Y(
        n12709) );
  CLKMX2X2 U11926 ( .A(\I_cache/cache[1][14] ), .B(n9392), .S0(n5110), .Y(
        n12710) );
  CLKMX2X2 U11927 ( .A(\I_cache/cache[0][14] ), .B(n9392), .S0(n5153), .Y(
        n12711) );
  CLKMX2X2 U11928 ( .A(\I_cache/cache[7][13] ), .B(n9372), .S0(n3617), .Y(
        n12712) );
  CLKMX2X2 U11929 ( .A(\I_cache/cache[6][13] ), .B(n9372), .S0(n5418), .Y(
        n12713) );
  CLKMX2X2 U11930 ( .A(\I_cache/cache[5][13] ), .B(n9372), .S0(n5284), .Y(
        n12714) );
  CLKMX2X2 U11931 ( .A(\I_cache/cache[4][13] ), .B(n9372), .S0(n4698), .Y(
        n12715) );
  CLKMX2X2 U11932 ( .A(\I_cache/cache[3][13] ), .B(n9372), .S0(n5198), .Y(
        n12716) );
  CLKMX2X2 U11933 ( .A(\I_cache/cache[2][13] ), .B(n9372), .S0(n5240), .Y(
        n12717) );
  CLKMX2X2 U11934 ( .A(\I_cache/cache[1][13] ), .B(n9372), .S0(n5102), .Y(
        n12718) );
  CLKMX2X2 U11935 ( .A(\I_cache/cache[0][13] ), .B(n9372), .S0(n5153), .Y(
        n12719) );
  CLKMX2X2 U11936 ( .A(\I_cache/cache[7][12] ), .B(n10085), .S0(n5366), .Y(
        n12720) );
  CLKMX2X2 U11937 ( .A(\I_cache/cache[6][12] ), .B(n10085), .S0(n5410), .Y(
        n12721) );
  CLKMX2X2 U11938 ( .A(\I_cache/cache[4][12] ), .B(n10085), .S0(n4681), .Y(
        n12723) );
  CLKMX2X2 U11939 ( .A(\I_cache/cache[3][12] ), .B(n10085), .S0(n5190), .Y(
        n12724) );
  CLKMX2X2 U11940 ( .A(\I_cache/cache[1][12] ), .B(n10085), .S0(n5103), .Y(
        n12726) );
  CLKMX2X2 U11941 ( .A(\I_cache/cache[0][12] ), .B(n10085), .S0(n5145), .Y(
        n12727) );
  CLKMX2X2 U11942 ( .A(\I_cache/cache[7][11] ), .B(n9954), .S0(n5372), .Y(
        n12728) );
  CLKMX2X2 U11943 ( .A(\I_cache/cache[6][11] ), .B(n9954), .S0(n5416), .Y(
        n12729) );
  CLKMX2X2 U11944 ( .A(\I_cache/cache[5][11] ), .B(n9954), .S0(n5282), .Y(
        n12730) );
  CLKMX2X2 U11945 ( .A(\I_cache/cache[4][11] ), .B(n9954), .S0(n5325), .Y(
        n12731) );
  CLKMX2X2 U11946 ( .A(\I_cache/cache[3][11] ), .B(n9954), .S0(n5196), .Y(
        n12732) );
  CLKMX2X2 U11947 ( .A(\I_cache/cache[2][11] ), .B(n9954), .S0(n5238), .Y(
        n12733) );
  CLKMX2X2 U11948 ( .A(\I_cache/cache[1][11] ), .B(n9954), .S0(n5109), .Y(
        n12734) );
  CLKMX2X2 U11949 ( .A(\I_cache/cache[0][11] ), .B(n9954), .S0(n5151), .Y(
        n12735) );
  CLKMX2X2 U11950 ( .A(\I_cache/cache[7][10] ), .B(n9659), .S0(n5374), .Y(
        n12736) );
  CLKMX2X2 U11951 ( .A(\I_cache/cache[6][10] ), .B(n9659), .S0(n5419), .Y(
        n12737) );
  CLKMX2X2 U11952 ( .A(\I_cache/cache[3][10] ), .B(n9659), .S0(n5199), .Y(
        n12740) );
  CLKMX2X2 U11953 ( .A(\I_cache/cache[2][10] ), .B(n9659), .S0(n5241), .Y(
        n12741) );
  CLKMX2X2 U11954 ( .A(\I_cache/cache[1][10] ), .B(n9659), .S0(n5110), .Y(
        n12742) );
  CLKMX2X2 U11955 ( .A(\I_cache/cache[0][10] ), .B(n9659), .S0(n5154), .Y(
        n12743) );
  CLKMX2X2 U11956 ( .A(\I_cache/cache[7][9] ), .B(n9645), .S0(n5374), .Y(
        n12744) );
  CLKMX2X2 U11957 ( .A(\I_cache/cache[6][9] ), .B(n9645), .S0(n5419), .Y(
        n12745) );
  CLKMX2X2 U11958 ( .A(\I_cache/cache[3][9] ), .B(n9645), .S0(n5199), .Y(
        n12748) );
  CLKMX2X2 U11959 ( .A(\I_cache/cache[2][9] ), .B(n9645), .S0(n5241), .Y(
        n12749) );
  CLKMX2X2 U11960 ( .A(\I_cache/cache[1][9] ), .B(n9645), .S0(n5110), .Y(
        n12750) );
  CLKMX2X2 U11961 ( .A(\I_cache/cache[0][9] ), .B(n9645), .S0(n5154), .Y(
        n12751) );
  CLKMX2X2 U11962 ( .A(\I_cache/cache[7][8] ), .B(n9421), .S0(n5373), .Y(
        n12752) );
  CLKMX2X2 U11963 ( .A(\I_cache/cache[6][8] ), .B(n9421), .S0(n5417), .Y(
        n12753) );
  CLKMX2X2 U11964 ( .A(\I_cache/cache[5][8] ), .B(n9421), .S0(n5283), .Y(
        n12754) );
  CLKMX2X2 U11965 ( .A(\I_cache/cache[4][8] ), .B(n9421), .S0(n5326), .Y(
        n12755) );
  CLKMX2X2 U11966 ( .A(\I_cache/cache[3][8] ), .B(n9421), .S0(n5197), .Y(
        n12756) );
  CLKMX2X2 U11967 ( .A(\I_cache/cache[2][8] ), .B(n9421), .S0(n5239), .Y(
        n12757) );
  CLKMX2X2 U11968 ( .A(\I_cache/cache[1][8] ), .B(n9421), .S0(n5111), .Y(
        n12758) );
  CLKMX2X2 U11969 ( .A(\I_cache/cache[0][8] ), .B(n9421), .S0(n5152), .Y(
        n12759) );
  CLKMX2X2 U11970 ( .A(\I_cache/cache[7][7] ), .B(n9825), .S0(n5368), .Y(
        n12760) );
  CLKMX2X2 U11971 ( .A(\I_cache/cache[6][7] ), .B(n9825), .S0(n5412), .Y(
        n12761) );
  CLKMX2X2 U11972 ( .A(\I_cache/cache[5][7] ), .B(n9825), .S0(n5285), .Y(
        n12762) );
  CLKMX2X2 U11973 ( .A(\I_cache/cache[4][7] ), .B(n9825), .S0(n5321), .Y(
        n12763) );
  CLKMX2X2 U11974 ( .A(\I_cache/cache[3][7] ), .B(n9825), .S0(n5192), .Y(
        n12764) );
  CLKMX2X2 U11975 ( .A(\I_cache/cache[2][7] ), .B(n9825), .S0(n5234), .Y(
        n12765) );
  CLKMX2X2 U11976 ( .A(\I_cache/cache[1][7] ), .B(n9825), .S0(n5105), .Y(
        n12766) );
  CLKMX2X2 U11977 ( .A(\I_cache/cache[0][7] ), .B(n9825), .S0(n5147), .Y(
        n12767) );
  CLKMX2X2 U11978 ( .A(\I_cache/cache[7][6] ), .B(n9436), .S0(n5373), .Y(
        n12768) );
  CLKMX2X2 U11979 ( .A(\I_cache/cache[6][6] ), .B(n9436), .S0(n5417), .Y(
        n12769) );
  CLKMX2X2 U11980 ( .A(\I_cache/cache[5][6] ), .B(n9436), .S0(n5283), .Y(
        n12770) );
  CLKMX2X2 U11981 ( .A(\I_cache/cache[4][6] ), .B(n9436), .S0(n5326), .Y(
        n12771) );
  CLKMX2X2 U11982 ( .A(\I_cache/cache[2][6] ), .B(n9436), .S0(n5239), .Y(
        n12773) );
  CLKMX2X2 U11983 ( .A(\I_cache/cache[0][6] ), .B(n9436), .S0(n5152), .Y(
        n12775) );
  CLKMX2X2 U11984 ( .A(\I_cache/cache[6][5] ), .B(n9541), .S0(n5419), .Y(
        n12777) );
  CLKMX2X2 U11985 ( .A(\I_cache/cache[4][5] ), .B(n9541), .S0(n5326), .Y(
        n12779) );
  CLKMX2X2 U11986 ( .A(\I_cache/cache[3][5] ), .B(n9541), .S0(n5193), .Y(
        n12780) );
  CLKMX2X2 U11987 ( .A(\I_cache/cache[2][5] ), .B(n9541), .S0(n5242), .Y(
        n12781) );
  CLKMX2X2 U11988 ( .A(\I_cache/cache[1][5] ), .B(n9541), .S0(n5111), .Y(
        n12782) );
  CLKMX2X2 U11989 ( .A(\I_cache/cache[0][5] ), .B(n9541), .S0(n5154), .Y(
        n12783) );
  CLKMX2X2 U11990 ( .A(\I_cache/cache[7][4] ), .B(n9458), .S0(n5373), .Y(
        n12784) );
  CLKMX2X2 U11991 ( .A(\I_cache/cache[6][4] ), .B(n9458), .S0(n5417), .Y(
        n12785) );
  CLKMX2X2 U11992 ( .A(\I_cache/cache[5][4] ), .B(n9458), .S0(n5283), .Y(
        n12786) );
  CLKMX2X2 U11993 ( .A(\I_cache/cache[4][4] ), .B(n9458), .S0(n5326), .Y(
        n12787) );
  CLKMX2X2 U11994 ( .A(\I_cache/cache[3][4] ), .B(n9458), .S0(n5197), .Y(
        n12788) );
  CLKMX2X2 U11995 ( .A(\I_cache/cache[2][4] ), .B(n9458), .S0(n5239), .Y(
        n12789) );
  CLKMX2X2 U11996 ( .A(\I_cache/cache[1][4] ), .B(n9458), .S0(n5108), .Y(
        n12790) );
  CLKMX2X2 U11997 ( .A(\I_cache/cache[0][4] ), .B(n9458), .S0(n5152), .Y(
        n12791) );
  CLKMX2X2 U11998 ( .A(\I_cache/cache[7][3] ), .B(n9512), .S0(n5371), .Y(
        n12792) );
  CLKMX2X2 U11999 ( .A(\I_cache/cache[6][3] ), .B(n9512), .S0(n5415), .Y(
        n12793) );
  CLKMX2X2 U12000 ( .A(\I_cache/cache[5][3] ), .B(n9512), .S0(n5285), .Y(
        n12794) );
  CLKMX2X2 U12001 ( .A(\I_cache/cache[4][3] ), .B(n9512), .S0(n5320), .Y(
        n12795) );
  CLKMX2X2 U12002 ( .A(\I_cache/cache[3][3] ), .B(n9512), .S0(n5195), .Y(
        n12796) );
  CLKMX2X2 U12003 ( .A(\I_cache/cache[2][3] ), .B(n9512), .S0(n5242), .Y(
        n12797) );
  CLKMX2X2 U12004 ( .A(\I_cache/cache[1][3] ), .B(n9512), .S0(n5111), .Y(
        n12798) );
  CLKMX2X2 U12005 ( .A(\I_cache/cache[0][3] ), .B(n9512), .S0(n5152), .Y(
        n12799) );
  CLKMX2X2 U12006 ( .A(\I_cache/cache[7][2] ), .B(n9477), .S0(n5373), .Y(
        n12800) );
  CLKMX2X2 U12007 ( .A(\I_cache/cache[6][2] ), .B(n9477), .S0(n5417), .Y(
        n12801) );
  CLKMX2X2 U12008 ( .A(\I_cache/cache[5][2] ), .B(n9477), .S0(n5283), .Y(
        n12802) );
  CLKMX2X2 U12009 ( .A(\I_cache/cache[4][2] ), .B(n9477), .S0(n5326), .Y(
        n12803) );
  CLKMX2X2 U12010 ( .A(\I_cache/cache[3][2] ), .B(n9477), .S0(n5197), .Y(
        n12804) );
  CLKMX2X2 U12011 ( .A(\I_cache/cache[2][2] ), .B(n9477), .S0(n5239), .Y(
        n12805) );
  CLKMX2X2 U12012 ( .A(\I_cache/cache[1][2] ), .B(n9477), .S0(n5103), .Y(
        n12806) );
  CLKMX2X2 U12013 ( .A(\I_cache/cache[0][2] ), .B(n9477), .S0(n5152), .Y(
        n12807) );
  CLKMX2X2 U12014 ( .A(\I_cache/cache[7][1] ), .B(n9356), .S0(n3617), .Y(
        n12808) );
  CLKMX2X2 U12015 ( .A(\I_cache/cache[6][1] ), .B(n9356), .S0(n5418), .Y(
        n12809) );
  CLKMX2X2 U12016 ( .A(\I_cache/cache[5][1] ), .B(n9356), .S0(n5284), .Y(
        n12810) );
  CLKMX2X2 U12017 ( .A(\I_cache/cache[3][1] ), .B(n9356), .S0(n5198), .Y(
        n12812) );
  CLKMX2X2 U12018 ( .A(\I_cache/cache[2][1] ), .B(n9356), .S0(n5240), .Y(
        n12813) );
  CLKMX2X2 U12019 ( .A(\I_cache/cache[1][1] ), .B(n9356), .S0(n5109), .Y(
        n12814) );
  CLKMX2X2 U12020 ( .A(\I_cache/cache[0][1] ), .B(n9356), .S0(n5153), .Y(
        n12815) );
  CLKMX2X2 U12021 ( .A(\I_cache/cache[7][0] ), .B(n9497), .S0(n5372), .Y(
        n12823) );
  CLKMX2X2 U12022 ( .A(\I_cache/cache[6][0] ), .B(n9497), .S0(n5413), .Y(
        n12816) );
  CLKMX2X2 U12023 ( .A(\I_cache/cache[5][0] ), .B(n9497), .S0(n5285), .Y(
        n12817) );
  CLKMX2X2 U12024 ( .A(\I_cache/cache[4][0] ), .B(n9497), .S0(n5323), .Y(
        n12818) );
  CLKMX2X2 U12025 ( .A(\I_cache/cache[3][0] ), .B(n9497), .S0(n5197), .Y(
        n12819) );
  CLKMX2X2 U12026 ( .A(\I_cache/cache[2][0] ), .B(n9497), .S0(n5242), .Y(
        n12820) );
  CLKMX2X2 U12027 ( .A(\I_cache/cache[1][0] ), .B(n9497), .S0(n5111), .Y(
        n12821) );
  CLKMX2X2 U12028 ( .A(\I_cache/cache[0][0] ), .B(n9497), .S0(n5151), .Y(
        n12822) );
  MX2XL U12029 ( .A(n3493), .B(net99009), .S0(n5507), .Y(\i_MIPS/n413 ) );
  MX2XL U12030 ( .A(n3494), .B(net98988), .S0(n5510), .Y(\i_MIPS/n411 ) );
  CLKMX2X2 U12031 ( .A(n9126), .B(\i_MIPS/Register/register[0][31] ), .S0(
        \i_MIPS/Register/n147 ), .Y(\i_MIPS/Register/n1139 ) );
  CLKMX2X2 U12032 ( .A(n5086), .B(\i_MIPS/Register/register[0][13] ), .S0(
        n5585), .Y(\i_MIPS/Register/n1121 ) );
  CLKMX2X2 U12033 ( .A(n5083), .B(\i_MIPS/Register/register[0][12] ), .S0(
        n5586), .Y(\i_MIPS/Register/n1120 ) );
  CLKMX2X2 U12034 ( .A(n5089), .B(\i_MIPS/Register/register[0][8] ), .S0(n5585), .Y(\i_MIPS/Register/n1116 ) );
  CLKMX2X2 U12035 ( .A(n5092), .B(\i_MIPS/Register/register[0][1] ), .S0(n5586), .Y(\i_MIPS/Register/n1109 ) );
  CLKMX2X2 U12036 ( .A(n5099), .B(\i_MIPS/Register/register[0][0] ), .S0(
        \i_MIPS/Register/n147 ), .Y(\i_MIPS/Register/n1108 ) );
  CLKMX2X2 U12037 ( .A(n5086), .B(\i_MIPS/Register/register[1][13] ), .S0(
        n5583), .Y(\i_MIPS/Register/n1089 ) );
  CLKMX2X2 U12038 ( .A(n5083), .B(\i_MIPS/Register/register[1][12] ), .S0(
        n5584), .Y(\i_MIPS/Register/n1088 ) );
  CLKMX2X2 U12039 ( .A(n5080), .B(\i_MIPS/Register/register[1][11] ), .S0(
        n5583), .Y(\i_MIPS/Register/n1087 ) );
  CLKMX2X2 U12040 ( .A(n5089), .B(\i_MIPS/Register/register[1][8] ), .S0(n5584), .Y(\i_MIPS/Register/n1084 ) );
  CLKMX2X2 U12041 ( .A(n5092), .B(\i_MIPS/Register/register[1][1] ), .S0(
        \i_MIPS/Register/n146 ), .Y(\i_MIPS/Register/n1077 ) );
  CLKMX2X2 U12042 ( .A(n5099), .B(\i_MIPS/Register/register[1][0] ), .S0(
        \i_MIPS/Register/n146 ), .Y(\i_MIPS/Register/n1076 ) );
  CLKMX2X2 U12043 ( .A(n5086), .B(\i_MIPS/Register/register[2][13] ), .S0(
        n5581), .Y(\i_MIPS/Register/n1057 ) );
  CLKMX2X2 U12044 ( .A(n5083), .B(\i_MIPS/Register/register[2][12] ), .S0(
        n5582), .Y(\i_MIPS/Register/n1056 ) );
  CLKMX2X2 U12045 ( .A(n5080), .B(\i_MIPS/Register/register[2][11] ), .S0(
        n5581), .Y(\i_MIPS/Register/n1055 ) );
  CLKMX2X2 U12046 ( .A(n5089), .B(\i_MIPS/Register/register[2][8] ), .S0(n5582), .Y(\i_MIPS/Register/n1052 ) );
  CLKMX2X2 U12047 ( .A(n5092), .B(\i_MIPS/Register/register[2][1] ), .S0(
        \i_MIPS/Register/n145 ), .Y(\i_MIPS/Register/n1045 ) );
  CLKMX2X2 U12048 ( .A(n5099), .B(\i_MIPS/Register/register[2][0] ), .S0(
        \i_MIPS/Register/n145 ), .Y(\i_MIPS/Register/n1044 ) );
  CLKMX2X2 U12049 ( .A(n5086), .B(\i_MIPS/Register/register[3][13] ), .S0(
        n5579), .Y(\i_MIPS/Register/n1025 ) );
  CLKMX2X2 U12050 ( .A(n5083), .B(\i_MIPS/Register/register[3][12] ), .S0(
        n5580), .Y(\i_MIPS/Register/n1024 ) );
  CLKMX2X2 U12051 ( .A(n5080), .B(\i_MIPS/Register/register[3][11] ), .S0(
        n5579), .Y(\i_MIPS/Register/n1023 ) );
  CLKMX2X2 U12052 ( .A(n5089), .B(\i_MIPS/Register/register[3][8] ), .S0(n5580), .Y(\i_MIPS/Register/n1020 ) );
  CLKMX2X2 U12053 ( .A(n5092), .B(\i_MIPS/Register/register[3][1] ), .S0(
        \i_MIPS/Register/n144 ), .Y(\i_MIPS/Register/n1013 ) );
  CLKMX2X2 U12054 ( .A(n5099), .B(\i_MIPS/Register/register[3][0] ), .S0(
        \i_MIPS/Register/n144 ), .Y(\i_MIPS/Register/n1012 ) );
  CLKMX2X2 U12055 ( .A(n5086), .B(\i_MIPS/Register/register[4][13] ), .S0(
        n5577), .Y(\i_MIPS/Register/n993 ) );
  CLKMX2X2 U12056 ( .A(n5083), .B(\i_MIPS/Register/register[4][12] ), .S0(
        n5578), .Y(\i_MIPS/Register/n992 ) );
  CLKMX2X2 U12057 ( .A(n5080), .B(\i_MIPS/Register/register[4][11] ), .S0(
        n5577), .Y(\i_MIPS/Register/n991 ) );
  CLKMX2X2 U12058 ( .A(n5089), .B(\i_MIPS/Register/register[4][8] ), .S0(n5578), .Y(\i_MIPS/Register/n988 ) );
  CLKMX2X2 U12059 ( .A(n5092), .B(\i_MIPS/Register/register[4][1] ), .S0(
        \i_MIPS/Register/n143 ), .Y(\i_MIPS/Register/n981 ) );
  CLKMX2X2 U12060 ( .A(n5099), .B(\i_MIPS/Register/register[4][0] ), .S0(
        \i_MIPS/Register/n143 ), .Y(\i_MIPS/Register/n980 ) );
  CLKMX2X2 U12061 ( .A(n5086), .B(\i_MIPS/Register/register[5][13] ), .S0(
        n5575), .Y(\i_MIPS/Register/n961 ) );
  CLKMX2X2 U12062 ( .A(n5083), .B(\i_MIPS/Register/register[5][12] ), .S0(
        n5576), .Y(\i_MIPS/Register/n960 ) );
  CLKMX2X2 U12063 ( .A(n5080), .B(\i_MIPS/Register/register[5][11] ), .S0(
        n5575), .Y(\i_MIPS/Register/n959 ) );
  CLKMX2X2 U12064 ( .A(n5089), .B(\i_MIPS/Register/register[5][8] ), .S0(n5576), .Y(\i_MIPS/Register/n956 ) );
  CLKMX2X2 U12065 ( .A(n5092), .B(\i_MIPS/Register/register[5][1] ), .S0(
        \i_MIPS/Register/n142 ), .Y(\i_MIPS/Register/n949 ) );
  CLKMX2X2 U12066 ( .A(n5099), .B(\i_MIPS/Register/register[5][0] ), .S0(
        \i_MIPS/Register/n142 ), .Y(\i_MIPS/Register/n948 ) );
  CLKMX2X2 U12067 ( .A(n5086), .B(\i_MIPS/Register/register[6][13] ), .S0(
        n5573), .Y(\i_MIPS/Register/n929 ) );
  CLKMX2X2 U12068 ( .A(n5083), .B(\i_MIPS/Register/register[6][12] ), .S0(
        n5574), .Y(\i_MIPS/Register/n928 ) );
  CLKMX2X2 U12069 ( .A(n5080), .B(\i_MIPS/Register/register[6][11] ), .S0(
        n5573), .Y(\i_MIPS/Register/n927 ) );
  CLKMX2X2 U12070 ( .A(n5089), .B(\i_MIPS/Register/register[6][8] ), .S0(n5574), .Y(\i_MIPS/Register/n924 ) );
  CLKMX2X2 U12071 ( .A(n5092), .B(\i_MIPS/Register/register[6][1] ), .S0(
        \i_MIPS/Register/n141 ), .Y(\i_MIPS/Register/n917 ) );
  CLKMX2X2 U12072 ( .A(n5099), .B(\i_MIPS/Register/register[6][0] ), .S0(
        \i_MIPS/Register/n141 ), .Y(\i_MIPS/Register/n916 ) );
  CLKMX2X2 U12073 ( .A(n5087), .B(\i_MIPS/Register/register[7][13] ), .S0(
        n5571), .Y(\i_MIPS/Register/n897 ) );
  CLKMX2X2 U12074 ( .A(n5084), .B(\i_MIPS/Register/register[7][12] ), .S0(
        n5572), .Y(\i_MIPS/Register/n896 ) );
  CLKMX2X2 U12075 ( .A(n5081), .B(\i_MIPS/Register/register[7][11] ), .S0(
        n5571), .Y(\i_MIPS/Register/n895 ) );
  CLKMX2X2 U12076 ( .A(n5090), .B(\i_MIPS/Register/register[7][8] ), .S0(n5572), .Y(\i_MIPS/Register/n892 ) );
  CLKMX2X2 U12077 ( .A(n5093), .B(\i_MIPS/Register/register[7][1] ), .S0(
        \i_MIPS/Register/n139 ), .Y(\i_MIPS/Register/n885 ) );
  CLKMX2X2 U12078 ( .A(n5100), .B(\i_MIPS/Register/register[7][0] ), .S0(
        \i_MIPS/Register/n139 ), .Y(\i_MIPS/Register/n884 ) );
  CLKMX2X2 U12079 ( .A(n5086), .B(\i_MIPS/Register/register[8][13] ), .S0(
        n5569), .Y(\i_MIPS/Register/n865 ) );
  CLKMX2X2 U12080 ( .A(n5083), .B(\i_MIPS/Register/register[8][12] ), .S0(
        n5570), .Y(\i_MIPS/Register/n864 ) );
  CLKMX2X2 U12081 ( .A(n5080), .B(\i_MIPS/Register/register[8][11] ), .S0(
        n5569), .Y(\i_MIPS/Register/n863 ) );
  CLKMX2X2 U12082 ( .A(n5089), .B(\i_MIPS/Register/register[8][8] ), .S0(n5570), .Y(\i_MIPS/Register/n860 ) );
  CLKMX2X2 U12083 ( .A(n5092), .B(\i_MIPS/Register/register[8][1] ), .S0(
        \i_MIPS/Register/n138 ), .Y(\i_MIPS/Register/n853 ) );
  CLKMX2X2 U12084 ( .A(n5099), .B(\i_MIPS/Register/register[8][0] ), .S0(
        \i_MIPS/Register/n138 ), .Y(\i_MIPS/Register/n852 ) );
  CLKMX2X2 U12085 ( .A(n5086), .B(\i_MIPS/Register/register[9][13] ), .S0(
        n5567), .Y(\i_MIPS/Register/n833 ) );
  CLKMX2X2 U12086 ( .A(n5083), .B(\i_MIPS/Register/register[9][12] ), .S0(
        n5568), .Y(\i_MIPS/Register/n832 ) );
  CLKMX2X2 U12087 ( .A(n5080), .B(\i_MIPS/Register/register[9][11] ), .S0(
        n5567), .Y(\i_MIPS/Register/n831 ) );
  CLKMX2X2 U12088 ( .A(n5089), .B(\i_MIPS/Register/register[9][8] ), .S0(n5568), .Y(\i_MIPS/Register/n828 ) );
  CLKMX2X2 U12089 ( .A(n5092), .B(\i_MIPS/Register/register[9][1] ), .S0(
        \i_MIPS/Register/n137 ), .Y(\i_MIPS/Register/n821 ) );
  CLKMX2X2 U12090 ( .A(n5099), .B(\i_MIPS/Register/register[9][0] ), .S0(
        \i_MIPS/Register/n137 ), .Y(\i_MIPS/Register/n820 ) );
  CLKMX2X2 U12091 ( .A(n5086), .B(\i_MIPS/Register/register[10][13] ), .S0(
        n5565), .Y(\i_MIPS/Register/n801 ) );
  CLKMX2X2 U12092 ( .A(n5083), .B(\i_MIPS/Register/register[10][12] ), .S0(
        n5566), .Y(\i_MIPS/Register/n800 ) );
  CLKMX2X2 U12093 ( .A(n5080), .B(\i_MIPS/Register/register[10][11] ), .S0(
        n5565), .Y(\i_MIPS/Register/n799 ) );
  CLKMX2X2 U12094 ( .A(n5089), .B(\i_MIPS/Register/register[10][8] ), .S0(
        n5566), .Y(\i_MIPS/Register/n796 ) );
  CLKMX2X2 U12095 ( .A(n5092), .B(\i_MIPS/Register/register[10][1] ), .S0(
        \i_MIPS/Register/n136 ), .Y(\i_MIPS/Register/n789 ) );
  CLKMX2X2 U12096 ( .A(n5099), .B(\i_MIPS/Register/register[10][0] ), .S0(
        \i_MIPS/Register/n136 ), .Y(\i_MIPS/Register/n788 ) );
  CLKMX2X2 U12097 ( .A(n5087), .B(\i_MIPS/Register/register[11][13] ), .S0(
        n5563), .Y(\i_MIPS/Register/n769 ) );
  CLKMX2X2 U12098 ( .A(n5084), .B(\i_MIPS/Register/register[11][12] ), .S0(
        n5564), .Y(\i_MIPS/Register/n768 ) );
  CLKMX2X2 U12099 ( .A(n5081), .B(\i_MIPS/Register/register[11][11] ), .S0(
        n5563), .Y(\i_MIPS/Register/n767 ) );
  CLKMX2X2 U12100 ( .A(n5090), .B(\i_MIPS/Register/register[11][8] ), .S0(
        n5564), .Y(\i_MIPS/Register/n764 ) );
  CLKMX2X2 U12101 ( .A(n5093), .B(\i_MIPS/Register/register[11][1] ), .S0(
        \i_MIPS/Register/n135 ), .Y(\i_MIPS/Register/n757 ) );
  CLKMX2X2 U12102 ( .A(n5099), .B(\i_MIPS/Register/register[11][0] ), .S0(
        \i_MIPS/Register/n135 ), .Y(\i_MIPS/Register/n756 ) );
  CLKMX2X2 U12103 ( .A(n5086), .B(\i_MIPS/Register/register[12][13] ), .S0(
        n5561), .Y(\i_MIPS/Register/n737 ) );
  CLKMX2X2 U12104 ( .A(n5083), .B(\i_MIPS/Register/register[12][12] ), .S0(
        n5562), .Y(\i_MIPS/Register/n736 ) );
  CLKMX2X2 U12105 ( .A(n5080), .B(\i_MIPS/Register/register[12][11] ), .S0(
        n5561), .Y(\i_MIPS/Register/n735 ) );
  CLKMX2X2 U12106 ( .A(n5089), .B(\i_MIPS/Register/register[12][8] ), .S0(
        n5562), .Y(\i_MIPS/Register/n732 ) );
  CLKMX2X2 U12107 ( .A(n5092), .B(\i_MIPS/Register/register[12][1] ), .S0(
        \i_MIPS/Register/n134 ), .Y(\i_MIPS/Register/n725 ) );
  CLKMX2X2 U12108 ( .A(n5099), .B(\i_MIPS/Register/register[12][0] ), .S0(
        \i_MIPS/Register/n134 ), .Y(\i_MIPS/Register/n724 ) );
  CLKMX2X2 U12109 ( .A(n5086), .B(\i_MIPS/Register/register[13][13] ), .S0(
        n5559), .Y(\i_MIPS/Register/n705 ) );
  CLKMX2X2 U12110 ( .A(n5083), .B(\i_MIPS/Register/register[13][12] ), .S0(
        n5560), .Y(\i_MIPS/Register/n704 ) );
  CLKMX2X2 U12111 ( .A(n5080), .B(\i_MIPS/Register/register[13][11] ), .S0(
        n5559), .Y(\i_MIPS/Register/n703 ) );
  CLKMX2X2 U12112 ( .A(n5089), .B(\i_MIPS/Register/register[13][8] ), .S0(
        n5560), .Y(\i_MIPS/Register/n700 ) );
  CLKMX2X2 U12113 ( .A(n5092), .B(\i_MIPS/Register/register[13][1] ), .S0(
        \i_MIPS/Register/n133 ), .Y(\i_MIPS/Register/n693 ) );
  CLKMX2X2 U12114 ( .A(n5099), .B(\i_MIPS/Register/register[13][0] ), .S0(
        \i_MIPS/Register/n133 ), .Y(\i_MIPS/Register/n692 ) );
  CLKMX2X2 U12115 ( .A(n5086), .B(\i_MIPS/Register/register[14][13] ), .S0(
        n5557), .Y(\i_MIPS/Register/n673 ) );
  CLKMX2X2 U12116 ( .A(n5083), .B(\i_MIPS/Register/register[14][12] ), .S0(
        n5558), .Y(\i_MIPS/Register/n672 ) );
  CLKMX2X2 U12117 ( .A(n5080), .B(\i_MIPS/Register/register[14][11] ), .S0(
        n5557), .Y(\i_MIPS/Register/n671 ) );
  CLKMX2X2 U12118 ( .A(n5089), .B(\i_MIPS/Register/register[14][8] ), .S0(
        n5558), .Y(\i_MIPS/Register/n668 ) );
  CLKMX2X2 U12119 ( .A(n5092), .B(\i_MIPS/Register/register[14][1] ), .S0(
        \i_MIPS/Register/n132 ), .Y(\i_MIPS/Register/n661 ) );
  CLKMX2X2 U12120 ( .A(n5099), .B(\i_MIPS/Register/register[14][0] ), .S0(
        \i_MIPS/Register/n132 ), .Y(\i_MIPS/Register/n660 ) );
  CLKMX2X2 U12121 ( .A(n5087), .B(\i_MIPS/Register/register[15][13] ), .S0(
        n5555), .Y(\i_MIPS/Register/n641 ) );
  CLKMX2X2 U12122 ( .A(n5084), .B(\i_MIPS/Register/register[15][12] ), .S0(
        n5556), .Y(\i_MIPS/Register/n640 ) );
  CLKMX2X2 U12123 ( .A(n5081), .B(\i_MIPS/Register/register[15][11] ), .S0(
        n5555), .Y(\i_MIPS/Register/n639 ) );
  CLKMX2X2 U12124 ( .A(n5090), .B(\i_MIPS/Register/register[15][8] ), .S0(
        n5556), .Y(\i_MIPS/Register/n636 ) );
  CLKMX2X2 U12125 ( .A(n5093), .B(\i_MIPS/Register/register[15][1] ), .S0(
        \i_MIPS/Register/n130 ), .Y(\i_MIPS/Register/n629 ) );
  CLKMX2X2 U12126 ( .A(n5100), .B(\i_MIPS/Register/register[15][0] ), .S0(
        \i_MIPS/Register/n130 ), .Y(\i_MIPS/Register/n628 ) );
  CLKMX2X2 U12127 ( .A(n5087), .B(\i_MIPS/Register/register[16][13] ), .S0(
        n5553), .Y(\i_MIPS/Register/n609 ) );
  CLKMX2X2 U12128 ( .A(n5084), .B(\i_MIPS/Register/register[16][12] ), .S0(
        n5554), .Y(\i_MIPS/Register/n608 ) );
  CLKMX2X2 U12129 ( .A(n5081), .B(\i_MIPS/Register/register[16][11] ), .S0(
        n5553), .Y(\i_MIPS/Register/n607 ) );
  CLKMX2X2 U12130 ( .A(n5090), .B(\i_MIPS/Register/register[16][8] ), .S0(
        n5554), .Y(\i_MIPS/Register/n604 ) );
  CLKMX2X2 U12131 ( .A(n5093), .B(\i_MIPS/Register/register[16][1] ), .S0(
        \i_MIPS/Register/n129 ), .Y(\i_MIPS/Register/n597 ) );
  CLKMX2X2 U12132 ( .A(n5100), .B(\i_MIPS/Register/register[16][0] ), .S0(
        \i_MIPS/Register/n129 ), .Y(\i_MIPS/Register/n596 ) );
  CLKMX2X2 U12133 ( .A(n5087), .B(\i_MIPS/Register/register[17][13] ), .S0(
        n5551), .Y(\i_MIPS/Register/n577 ) );
  CLKMX2X2 U12134 ( .A(n5084), .B(\i_MIPS/Register/register[17][12] ), .S0(
        n5552), .Y(\i_MIPS/Register/n576 ) );
  CLKMX2X2 U12135 ( .A(n5081), .B(\i_MIPS/Register/register[17][11] ), .S0(
        n5551), .Y(\i_MIPS/Register/n575 ) );
  CLKMX2X2 U12136 ( .A(n5090), .B(\i_MIPS/Register/register[17][8] ), .S0(
        n5552), .Y(\i_MIPS/Register/n572 ) );
  CLKMX2X2 U12137 ( .A(n5093), .B(\i_MIPS/Register/register[17][1] ), .S0(
        \i_MIPS/Register/n128 ), .Y(\i_MIPS/Register/n565 ) );
  CLKMX2X2 U12138 ( .A(n5100), .B(\i_MIPS/Register/register[17][0] ), .S0(
        \i_MIPS/Register/n128 ), .Y(\i_MIPS/Register/n564 ) );
  CLKMX2X2 U12139 ( .A(n5087), .B(\i_MIPS/Register/register[18][13] ), .S0(
        n5549), .Y(\i_MIPS/Register/n545 ) );
  CLKMX2X2 U12140 ( .A(n5084), .B(\i_MIPS/Register/register[18][12] ), .S0(
        n5550), .Y(\i_MIPS/Register/n544 ) );
  CLKMX2X2 U12141 ( .A(n5081), .B(\i_MIPS/Register/register[18][11] ), .S0(
        n5549), .Y(\i_MIPS/Register/n543 ) );
  CLKMX2X2 U12142 ( .A(n5090), .B(\i_MIPS/Register/register[18][8] ), .S0(
        n5550), .Y(\i_MIPS/Register/n540 ) );
  CLKMX2X2 U12143 ( .A(n5093), .B(\i_MIPS/Register/register[18][1] ), .S0(
        \i_MIPS/Register/n127 ), .Y(\i_MIPS/Register/n533 ) );
  CLKMX2X2 U12144 ( .A(n5100), .B(\i_MIPS/Register/register[18][0] ), .S0(
        \i_MIPS/Register/n127 ), .Y(\i_MIPS/Register/n532 ) );
  CLKMX2X2 U12145 ( .A(n5086), .B(\i_MIPS/Register/register[19][13] ), .S0(
        n5547), .Y(\i_MIPS/Register/n513 ) );
  CLKMX2X2 U12146 ( .A(n5083), .B(\i_MIPS/Register/register[19][12] ), .S0(
        n5548), .Y(\i_MIPS/Register/n512 ) );
  CLKMX2X2 U12147 ( .A(n5081), .B(\i_MIPS/Register/register[19][11] ), .S0(
        \i_MIPS/Register/n126 ), .Y(\i_MIPS/Register/n511 ) );
  CLKMX2X2 U12148 ( .A(n5089), .B(\i_MIPS/Register/register[19][8] ), .S0(
        n5547), .Y(\i_MIPS/Register/n508 ) );
  CLKMX2X2 U12149 ( .A(n5093), .B(\i_MIPS/Register/register[19][1] ), .S0(
        n5548), .Y(\i_MIPS/Register/n501 ) );
  CLKMX2X2 U12150 ( .A(n5100), .B(\i_MIPS/Register/register[19][0] ), .S0(
        \i_MIPS/Register/n126 ), .Y(\i_MIPS/Register/n500 ) );
  CLKMX2X2 U12151 ( .A(n5087), .B(\i_MIPS/Register/register[20][13] ), .S0(
        n5545), .Y(\i_MIPS/Register/n481 ) );
  CLKMX2X2 U12152 ( .A(n5084), .B(\i_MIPS/Register/register[20][12] ), .S0(
        n5546), .Y(\i_MIPS/Register/n480 ) );
  CLKMX2X2 U12153 ( .A(n5081), .B(\i_MIPS/Register/register[20][11] ), .S0(
        n5545), .Y(\i_MIPS/Register/n479 ) );
  CLKMX2X2 U12154 ( .A(n5090), .B(\i_MIPS/Register/register[20][8] ), .S0(
        n5546), .Y(\i_MIPS/Register/n476 ) );
  CLKMX2X2 U12155 ( .A(n5093), .B(\i_MIPS/Register/register[20][1] ), .S0(
        \i_MIPS/Register/n125 ), .Y(\i_MIPS/Register/n469 ) );
  CLKMX2X2 U12156 ( .A(n5100), .B(\i_MIPS/Register/register[20][0] ), .S0(
        \i_MIPS/Register/n125 ), .Y(\i_MIPS/Register/n468 ) );
  CLKMX2X2 U12157 ( .A(n5087), .B(\i_MIPS/Register/register[21][13] ), .S0(
        n5544), .Y(\i_MIPS/Register/n449 ) );
  CLKMX2X2 U12158 ( .A(n5084), .B(\i_MIPS/Register/register[21][12] ), .S0(
        n5543), .Y(\i_MIPS/Register/n448 ) );
  CLKMX2X2 U12159 ( .A(n5080), .B(\i_MIPS/Register/register[21][11] ), .S0(
        \i_MIPS/Register/n124 ), .Y(\i_MIPS/Register/n447 ) );
  CLKMX2X2 U12160 ( .A(n5090), .B(\i_MIPS/Register/register[21][8] ), .S0(
        n5544), .Y(\i_MIPS/Register/n444 ) );
  CLKMX2X2 U12161 ( .A(n5093), .B(\i_MIPS/Register/register[21][1] ), .S0(
        \i_MIPS/Register/n124 ), .Y(\i_MIPS/Register/n437 ) );
  CLKMX2X2 U12162 ( .A(n5100), .B(\i_MIPS/Register/register[21][0] ), .S0(
        n5543), .Y(\i_MIPS/Register/n436 ) );
  CLKMX2X2 U12163 ( .A(n5087), .B(\i_MIPS/Register/register[22][13] ), .S0(
        n5541), .Y(\i_MIPS/Register/n417 ) );
  CLKMX2X2 U12164 ( .A(n5084), .B(\i_MIPS/Register/register[22][12] ), .S0(
        n5542), .Y(\i_MIPS/Register/n416 ) );
  CLKMX2X2 U12165 ( .A(n5081), .B(\i_MIPS/Register/register[22][11] ), .S0(
        n5541), .Y(\i_MIPS/Register/n415 ) );
  CLKMX2X2 U12166 ( .A(n5090), .B(\i_MIPS/Register/register[22][8] ), .S0(
        n5542), .Y(\i_MIPS/Register/n412 ) );
  CLKMX2X2 U12167 ( .A(n5093), .B(\i_MIPS/Register/register[22][1] ), .S0(
        \i_MIPS/Register/n123 ), .Y(\i_MIPS/Register/n405 ) );
  CLKMX2X2 U12168 ( .A(n5100), .B(\i_MIPS/Register/register[22][0] ), .S0(
        \i_MIPS/Register/n123 ), .Y(\i_MIPS/Register/n404 ) );
  CLKMX2X2 U12169 ( .A(n5086), .B(\i_MIPS/Register/register[23][13] ), .S0(
        n5539), .Y(\i_MIPS/Register/n385 ) );
  CLKMX2X2 U12170 ( .A(n5083), .B(\i_MIPS/Register/register[23][12] ), .S0(
        n5540), .Y(\i_MIPS/Register/n384 ) );
  CLKMX2X2 U12171 ( .A(n5080), .B(\i_MIPS/Register/register[23][11] ), .S0(
        \i_MIPS/Register/n121 ), .Y(\i_MIPS/Register/n383 ) );
  CLKMX2X2 U12172 ( .A(n5089), .B(\i_MIPS/Register/register[23][8] ), .S0(
        n5539), .Y(\i_MIPS/Register/n380 ) );
  CLKMX2X2 U12173 ( .A(n5092), .B(\i_MIPS/Register/register[23][1] ), .S0(
        n5540), .Y(\i_MIPS/Register/n373 ) );
  CLKMX2X2 U12174 ( .A(n5099), .B(\i_MIPS/Register/register[23][0] ), .S0(
        \i_MIPS/Register/n121 ), .Y(\i_MIPS/Register/n372 ) );
  CLKMX2X2 U12175 ( .A(n5087), .B(\i_MIPS/Register/register[24][13] ), .S0(
        n5537), .Y(\i_MIPS/Register/n353 ) );
  CLKMX2X2 U12176 ( .A(n5084), .B(\i_MIPS/Register/register[24][12] ), .S0(
        n5538), .Y(\i_MIPS/Register/n352 ) );
  CLKMX2X2 U12177 ( .A(n5081), .B(\i_MIPS/Register/register[24][11] ), .S0(
        n5537), .Y(\i_MIPS/Register/n351 ) );
  CLKMX2X2 U12178 ( .A(n5090), .B(\i_MIPS/Register/register[24][8] ), .S0(
        n5538), .Y(\i_MIPS/Register/n348 ) );
  CLKMX2X2 U12179 ( .A(n5093), .B(\i_MIPS/Register/register[24][1] ), .S0(
        \i_MIPS/Register/n118 ), .Y(\i_MIPS/Register/n341 ) );
  CLKMX2X2 U12180 ( .A(n5100), .B(\i_MIPS/Register/register[24][0] ), .S0(
        \i_MIPS/Register/n118 ), .Y(\i_MIPS/Register/n340 ) );
  CLKMX2X2 U12181 ( .A(n5087), .B(\i_MIPS/Register/register[25][13] ), .S0(
        n5535), .Y(\i_MIPS/Register/n321 ) );
  CLKMX2X2 U12182 ( .A(n5084), .B(\i_MIPS/Register/register[25][12] ), .S0(
        n5536), .Y(\i_MIPS/Register/n320 ) );
  CLKMX2X2 U12183 ( .A(n5081), .B(\i_MIPS/Register/register[25][11] ), .S0(
        n5535), .Y(\i_MIPS/Register/n319 ) );
  CLKMX2X2 U12184 ( .A(n5090), .B(\i_MIPS/Register/register[25][8] ), .S0(
        n5536), .Y(\i_MIPS/Register/n316 ) );
  CLKMX2X2 U12185 ( .A(n5093), .B(\i_MIPS/Register/register[25][1] ), .S0(
        \i_MIPS/Register/n116 ), .Y(\i_MIPS/Register/n309 ) );
  CLKMX2X2 U12186 ( .A(n5100), .B(\i_MIPS/Register/register[25][0] ), .S0(
        \i_MIPS/Register/n116 ), .Y(\i_MIPS/Register/n308 ) );
  CLKMX2X2 U12187 ( .A(n5087), .B(\i_MIPS/Register/register[26][13] ), .S0(
        n5533), .Y(\i_MIPS/Register/n289 ) );
  CLKMX2X2 U12188 ( .A(n5084), .B(\i_MIPS/Register/register[26][12] ), .S0(
        n5534), .Y(\i_MIPS/Register/n288 ) );
  CLKMX2X2 U12189 ( .A(n5081), .B(\i_MIPS/Register/register[26][11] ), .S0(
        n5533), .Y(\i_MIPS/Register/n287 ) );
  CLKMX2X2 U12190 ( .A(n5090), .B(\i_MIPS/Register/register[26][8] ), .S0(
        n5534), .Y(\i_MIPS/Register/n284 ) );
  CLKMX2X2 U12191 ( .A(n5093), .B(\i_MIPS/Register/register[26][1] ), .S0(
        \i_MIPS/Register/n114 ), .Y(\i_MIPS/Register/n277 ) );
  CLKMX2X2 U12192 ( .A(n5100), .B(\i_MIPS/Register/register[26][0] ), .S0(
        \i_MIPS/Register/n114 ), .Y(\i_MIPS/Register/n276 ) );
  CLKMX2X2 U12193 ( .A(n5087), .B(\i_MIPS/Register/register[27][13] ), .S0(
        n5531), .Y(\i_MIPS/Register/n257 ) );
  CLKMX2X2 U12194 ( .A(n5084), .B(\i_MIPS/Register/register[27][12] ), .S0(
        n5532), .Y(\i_MIPS/Register/n256 ) );
  CLKMX2X2 U12195 ( .A(n5081), .B(\i_MIPS/Register/register[27][11] ), .S0(
        \i_MIPS/Register/n112 ), .Y(\i_MIPS/Register/n255 ) );
  CLKMX2X2 U12196 ( .A(n5090), .B(\i_MIPS/Register/register[27][8] ), .S0(
        n5531), .Y(\i_MIPS/Register/n252 ) );
  CLKMX2X2 U12197 ( .A(n5093), .B(\i_MIPS/Register/register[27][1] ), .S0(
        n5532), .Y(\i_MIPS/Register/n245 ) );
  CLKMX2X2 U12198 ( .A(n5100), .B(\i_MIPS/Register/register[27][0] ), .S0(
        \i_MIPS/Register/n112 ), .Y(\i_MIPS/Register/n244 ) );
  CLKMX2X2 U12199 ( .A(n5087), .B(\i_MIPS/Register/register[28][13] ), .S0(
        n5529), .Y(\i_MIPS/Register/n225 ) );
  CLKMX2X2 U12200 ( .A(n5084), .B(\i_MIPS/Register/register[28][12] ), .S0(
        n5530), .Y(\i_MIPS/Register/n224 ) );
  CLKMX2X2 U12201 ( .A(n5081), .B(\i_MIPS/Register/register[28][11] ), .S0(
        n5529), .Y(\i_MIPS/Register/n223 ) );
  CLKMX2X2 U12202 ( .A(n5090), .B(\i_MIPS/Register/register[28][8] ), .S0(
        n5530), .Y(\i_MIPS/Register/n220 ) );
  CLKMX2X2 U12203 ( .A(n5093), .B(\i_MIPS/Register/register[28][1] ), .S0(
        \i_MIPS/Register/n110 ), .Y(\i_MIPS/Register/n213 ) );
  CLKMX2X2 U12204 ( .A(n5100), .B(\i_MIPS/Register/register[28][0] ), .S0(
        \i_MIPS/Register/n110 ), .Y(\i_MIPS/Register/n212 ) );
  CLKMX2X2 U12205 ( .A(n5086), .B(\i_MIPS/Register/register[29][13] ), .S0(
        n5527), .Y(\i_MIPS/Register/n193 ) );
  CLKMX2X2 U12206 ( .A(n5083), .B(\i_MIPS/Register/register[29][12] ), .S0(
        n5528), .Y(\i_MIPS/Register/n192 ) );
  CLKMX2X2 U12207 ( .A(n5080), .B(\i_MIPS/Register/register[29][11] ), .S0(
        \i_MIPS/Register/n108 ), .Y(\i_MIPS/Register/n191 ) );
  CLKMX2X2 U12208 ( .A(n5089), .B(\i_MIPS/Register/register[29][8] ), .S0(
        n5527), .Y(\i_MIPS/Register/n188 ) );
  CLKMX2X2 U12209 ( .A(n5092), .B(\i_MIPS/Register/register[29][1] ), .S0(
        n5528), .Y(\i_MIPS/Register/n181 ) );
  CLKMX2X2 U12210 ( .A(n5099), .B(\i_MIPS/Register/register[29][0] ), .S0(
        \i_MIPS/Register/n108 ), .Y(\i_MIPS/Register/n180 ) );
  CLKMX2X2 U12211 ( .A(n5087), .B(\i_MIPS/Register/register[30][13] ), .S0(
        n5525), .Y(\i_MIPS/Register/n161 ) );
  CLKMX2X2 U12212 ( .A(n5084), .B(\i_MIPS/Register/register[30][12] ), .S0(
        n5526), .Y(\i_MIPS/Register/n160 ) );
  CLKMX2X2 U12213 ( .A(n5081), .B(\i_MIPS/Register/register[30][11] ), .S0(
        n5525), .Y(\i_MIPS/Register/n159 ) );
  CLKMX2X2 U12214 ( .A(n5090), .B(\i_MIPS/Register/register[30][8] ), .S0(
        n5526), .Y(\i_MIPS/Register/n156 ) );
  CLKMX2X2 U12215 ( .A(n5093), .B(\i_MIPS/Register/register[30][1] ), .S0(
        \i_MIPS/Register/n106 ), .Y(\i_MIPS/Register/n149 ) );
  CLKMX2X2 U12216 ( .A(n5100), .B(\i_MIPS/Register/register[30][0] ), .S0(
        \i_MIPS/Register/n106 ), .Y(\i_MIPS/Register/n148 ) );
  MXI2X1 U12217 ( .A(n4707), .B(\i_MIPS/n221 ), .S0(n5511), .Y(\i_MIPS/n503 )
         );
  CLKMX2X2 U12218 ( .A(n5036), .B(\i_MIPS/Register/register[0][20] ), .S0(
        n5585), .Y(\i_MIPS/Register/n1128 ) );
  CLKMX2X2 U12219 ( .A(n5006), .B(\i_MIPS/Register/register[0][4] ), .S0(n5585), .Y(\i_MIPS/Register/n1112 ) );
  CLKMX2X2 U12220 ( .A(n5071), .B(\i_MIPS/Register/register[0][2] ), .S0(n5586), .Y(\i_MIPS/Register/n1110 ) );
  CLKMX2X2 U12221 ( .A(n5036), .B(\i_MIPS/Register/register[1][20] ), .S0(
        n5583), .Y(\i_MIPS/Register/n1096 ) );
  CLKMX2X2 U12222 ( .A(n5006), .B(\i_MIPS/Register/register[1][4] ), .S0(n5583), .Y(\i_MIPS/Register/n1080 ) );
  CLKMX2X2 U12223 ( .A(n5071), .B(\i_MIPS/Register/register[1][2] ), .S0(n5584), .Y(\i_MIPS/Register/n1078 ) );
  CLKMX2X2 U12224 ( .A(n5036), .B(\i_MIPS/Register/register[2][20] ), .S0(
        n5581), .Y(\i_MIPS/Register/n1064 ) );
  CLKMX2X2 U12225 ( .A(n5006), .B(\i_MIPS/Register/register[2][4] ), .S0(n5581), .Y(\i_MIPS/Register/n1048 ) );
  CLKMX2X2 U12226 ( .A(n5071), .B(\i_MIPS/Register/register[2][2] ), .S0(n5582), .Y(\i_MIPS/Register/n1046 ) );
  CLKMX2X2 U12227 ( .A(n5036), .B(\i_MIPS/Register/register[3][20] ), .S0(
        n5579), .Y(\i_MIPS/Register/n1032 ) );
  CLKMX2X2 U12228 ( .A(n5006), .B(\i_MIPS/Register/register[3][4] ), .S0(n5579), .Y(\i_MIPS/Register/n1016 ) );
  CLKMX2X2 U12229 ( .A(n5071), .B(\i_MIPS/Register/register[3][2] ), .S0(n5580), .Y(\i_MIPS/Register/n1014 ) );
  CLKMX2X2 U12230 ( .A(n5036), .B(\i_MIPS/Register/register[4][20] ), .S0(
        n5577), .Y(\i_MIPS/Register/n1000 ) );
  CLKMX2X2 U12231 ( .A(n5006), .B(\i_MIPS/Register/register[4][4] ), .S0(n5577), .Y(\i_MIPS/Register/n984 ) );
  CLKMX2X2 U12232 ( .A(n5071), .B(\i_MIPS/Register/register[4][2] ), .S0(n5578), .Y(\i_MIPS/Register/n982 ) );
  CLKMX2X2 U12233 ( .A(n5036), .B(\i_MIPS/Register/register[5][20] ), .S0(
        n5575), .Y(\i_MIPS/Register/n968 ) );
  CLKMX2X2 U12234 ( .A(n5006), .B(\i_MIPS/Register/register[5][4] ), .S0(n5575), .Y(\i_MIPS/Register/n952 ) );
  CLKMX2X2 U12235 ( .A(n5071), .B(\i_MIPS/Register/register[5][2] ), .S0(n5576), .Y(\i_MIPS/Register/n950 ) );
  CLKMX2X2 U12236 ( .A(n5036), .B(\i_MIPS/Register/register[6][20] ), .S0(
        n5573), .Y(\i_MIPS/Register/n936 ) );
  CLKMX2X2 U12237 ( .A(n5006), .B(\i_MIPS/Register/register[6][4] ), .S0(n5573), .Y(\i_MIPS/Register/n920 ) );
  CLKMX2X2 U12238 ( .A(n5071), .B(\i_MIPS/Register/register[6][2] ), .S0(n5574), .Y(\i_MIPS/Register/n918 ) );
  CLKMX2X2 U12239 ( .A(n5037), .B(\i_MIPS/Register/register[7][20] ), .S0(
        n5571), .Y(\i_MIPS/Register/n904 ) );
  CLKMX2X2 U12240 ( .A(n5007), .B(\i_MIPS/Register/register[7][4] ), .S0(n5571), .Y(\i_MIPS/Register/n888 ) );
  CLKMX2X2 U12241 ( .A(n5072), .B(\i_MIPS/Register/register[7][2] ), .S0(n5572), .Y(\i_MIPS/Register/n886 ) );
  CLKMX2X2 U12242 ( .A(n5036), .B(\i_MIPS/Register/register[8][20] ), .S0(
        n5569), .Y(\i_MIPS/Register/n872 ) );
  CLKMX2X2 U12243 ( .A(n5006), .B(\i_MIPS/Register/register[8][4] ), .S0(n5569), .Y(\i_MIPS/Register/n856 ) );
  CLKMX2X2 U12244 ( .A(n5071), .B(\i_MIPS/Register/register[8][2] ), .S0(n5570), .Y(\i_MIPS/Register/n854 ) );
  CLKMX2X2 U12245 ( .A(n5036), .B(\i_MIPS/Register/register[9][20] ), .S0(
        n5567), .Y(\i_MIPS/Register/n840 ) );
  CLKMX2X2 U12246 ( .A(n5006), .B(\i_MIPS/Register/register[9][4] ), .S0(n5567), .Y(\i_MIPS/Register/n824 ) );
  CLKMX2X2 U12247 ( .A(n5071), .B(\i_MIPS/Register/register[9][2] ), .S0(n5568), .Y(\i_MIPS/Register/n822 ) );
  CLKMX2X2 U12248 ( .A(n5036), .B(\i_MIPS/Register/register[10][20] ), .S0(
        n5565), .Y(\i_MIPS/Register/n808 ) );
  CLKMX2X2 U12249 ( .A(n5006), .B(\i_MIPS/Register/register[10][4] ), .S0(
        n5565), .Y(\i_MIPS/Register/n792 ) );
  CLKMX2X2 U12250 ( .A(n5071), .B(\i_MIPS/Register/register[10][2] ), .S0(
        n5566), .Y(\i_MIPS/Register/n790 ) );
  CLKMX2X2 U12251 ( .A(n5036), .B(\i_MIPS/Register/register[11][20] ), .S0(
        n5563), .Y(\i_MIPS/Register/n776 ) );
  CLKMX2X2 U12252 ( .A(n5007), .B(\i_MIPS/Register/register[11][4] ), .S0(
        n5563), .Y(\i_MIPS/Register/n760 ) );
  CLKMX2X2 U12253 ( .A(n5072), .B(\i_MIPS/Register/register[11][2] ), .S0(
        n5564), .Y(\i_MIPS/Register/n758 ) );
  CLKMX2X2 U12254 ( .A(n5036), .B(\i_MIPS/Register/register[12][20] ), .S0(
        n5561), .Y(\i_MIPS/Register/n744 ) );
  CLKMX2X2 U12255 ( .A(n5006), .B(\i_MIPS/Register/register[12][4] ), .S0(
        n5561), .Y(\i_MIPS/Register/n728 ) );
  CLKMX2X2 U12256 ( .A(n5071), .B(\i_MIPS/Register/register[12][2] ), .S0(
        n5562), .Y(\i_MIPS/Register/n726 ) );
  CLKMX2X2 U12257 ( .A(n5036), .B(\i_MIPS/Register/register[13][20] ), .S0(
        n5559), .Y(\i_MIPS/Register/n712 ) );
  CLKMX2X2 U12258 ( .A(n5006), .B(\i_MIPS/Register/register[13][4] ), .S0(
        n5559), .Y(\i_MIPS/Register/n696 ) );
  CLKMX2X2 U12259 ( .A(n5071), .B(\i_MIPS/Register/register[13][2] ), .S0(
        n5560), .Y(\i_MIPS/Register/n694 ) );
  CLKMX2X2 U12260 ( .A(n5036), .B(\i_MIPS/Register/register[14][20] ), .S0(
        n5557), .Y(\i_MIPS/Register/n680 ) );
  CLKMX2X2 U12261 ( .A(n5006), .B(\i_MIPS/Register/register[14][4] ), .S0(
        n5557), .Y(\i_MIPS/Register/n664 ) );
  CLKMX2X2 U12262 ( .A(n5071), .B(\i_MIPS/Register/register[14][2] ), .S0(
        n5558), .Y(\i_MIPS/Register/n662 ) );
  CLKMX2X2 U12263 ( .A(n5037), .B(\i_MIPS/Register/register[15][20] ), .S0(
        n5555), .Y(\i_MIPS/Register/n648 ) );
  CLKMX2X2 U12264 ( .A(n5007), .B(\i_MIPS/Register/register[15][4] ), .S0(
        n5555), .Y(\i_MIPS/Register/n632 ) );
  CLKMX2X2 U12265 ( .A(n5072), .B(\i_MIPS/Register/register[15][2] ), .S0(
        n5556), .Y(\i_MIPS/Register/n630 ) );
  CLKMX2X2 U12266 ( .A(n5037), .B(\i_MIPS/Register/register[16][20] ), .S0(
        n5553), .Y(\i_MIPS/Register/n616 ) );
  CLKMX2X2 U12267 ( .A(n5007), .B(\i_MIPS/Register/register[16][4] ), .S0(
        n5553), .Y(\i_MIPS/Register/n600 ) );
  CLKMX2X2 U12268 ( .A(n5072), .B(\i_MIPS/Register/register[16][2] ), .S0(
        n5554), .Y(\i_MIPS/Register/n598 ) );
  CLKMX2X2 U12269 ( .A(n5037), .B(\i_MIPS/Register/register[17][20] ), .S0(
        n5551), .Y(\i_MIPS/Register/n584 ) );
  CLKMX2X2 U12270 ( .A(n5007), .B(\i_MIPS/Register/register[17][4] ), .S0(
        n5551), .Y(\i_MIPS/Register/n568 ) );
  CLKMX2X2 U12271 ( .A(n5072), .B(\i_MIPS/Register/register[17][2] ), .S0(
        n5552), .Y(\i_MIPS/Register/n566 ) );
  CLKMX2X2 U12272 ( .A(n5037), .B(\i_MIPS/Register/register[18][20] ), .S0(
        n5549), .Y(\i_MIPS/Register/n552 ) );
  CLKMX2X2 U12273 ( .A(n5007), .B(\i_MIPS/Register/register[18][4] ), .S0(
        n5549), .Y(\i_MIPS/Register/n536 ) );
  CLKMX2X2 U12274 ( .A(n5072), .B(\i_MIPS/Register/register[18][2] ), .S0(
        n5550), .Y(\i_MIPS/Register/n534 ) );
  CLKMX2X2 U12275 ( .A(n5037), .B(\i_MIPS/Register/register[19][20] ), .S0(
        n5547), .Y(\i_MIPS/Register/n520 ) );
  CLKMX2X2 U12276 ( .A(n5007), .B(\i_MIPS/Register/register[19][4] ), .S0(
        n5547), .Y(\i_MIPS/Register/n504 ) );
  CLKMX2X2 U12277 ( .A(n5037), .B(\i_MIPS/Register/register[20][20] ), .S0(
        n5545), .Y(\i_MIPS/Register/n488 ) );
  CLKMX2X2 U12278 ( .A(n5007), .B(\i_MIPS/Register/register[20][4] ), .S0(
        n5545), .Y(\i_MIPS/Register/n472 ) );
  CLKMX2X2 U12279 ( .A(n5072), .B(\i_MIPS/Register/register[20][2] ), .S0(
        n5546), .Y(\i_MIPS/Register/n470 ) );
  CLKMX2X2 U12280 ( .A(n5037), .B(\i_MIPS/Register/register[21][20] ), .S0(
        n5543), .Y(\i_MIPS/Register/n456 ) );
  CLKMX2X2 U12281 ( .A(n5007), .B(\i_MIPS/Register/register[21][4] ), .S0(
        n5543), .Y(\i_MIPS/Register/n440 ) );
  CLKMX2X2 U12282 ( .A(n5037), .B(\i_MIPS/Register/register[22][20] ), .S0(
        n5541), .Y(\i_MIPS/Register/n424 ) );
  CLKMX2X2 U12283 ( .A(n5006), .B(\i_MIPS/Register/register[22][4] ), .S0(
        n5541), .Y(\i_MIPS/Register/n408 ) );
  CLKMX2X2 U12284 ( .A(n5072), .B(\i_MIPS/Register/register[22][2] ), .S0(
        n5542), .Y(\i_MIPS/Register/n406 ) );
  CLKMX2X2 U12285 ( .A(n5036), .B(\i_MIPS/Register/register[23][20] ), .S0(
        n5539), .Y(\i_MIPS/Register/n392 ) );
  CLKMX2X2 U12286 ( .A(n5007), .B(\i_MIPS/Register/register[23][4] ), .S0(
        n5539), .Y(\i_MIPS/Register/n376 ) );
  CLKMX2X2 U12287 ( .A(n5037), .B(\i_MIPS/Register/register[24][20] ), .S0(
        n5537), .Y(\i_MIPS/Register/n360 ) );
  CLKMX2X2 U12288 ( .A(n5007), .B(\i_MIPS/Register/register[24][4] ), .S0(
        n5537), .Y(\i_MIPS/Register/n344 ) );
  CLKMX2X2 U12289 ( .A(n5072), .B(\i_MIPS/Register/register[24][2] ), .S0(
        n5538), .Y(\i_MIPS/Register/n342 ) );
  CLKMX2X2 U12290 ( .A(n5037), .B(\i_MIPS/Register/register[25][20] ), .S0(
        n5535), .Y(\i_MIPS/Register/n328 ) );
  CLKMX2X2 U12291 ( .A(n5006), .B(\i_MIPS/Register/register[25][4] ), .S0(
        n5535), .Y(\i_MIPS/Register/n312 ) );
  CLKMX2X2 U12292 ( .A(n5072), .B(\i_MIPS/Register/register[25][2] ), .S0(
        n5536), .Y(\i_MIPS/Register/n310 ) );
  CLKMX2X2 U12293 ( .A(n5037), .B(\i_MIPS/Register/register[26][20] ), .S0(
        n5533), .Y(\i_MIPS/Register/n296 ) );
  CLKMX2X2 U12294 ( .A(n5007), .B(\i_MIPS/Register/register[26][4] ), .S0(
        n5533), .Y(\i_MIPS/Register/n280 ) );
  CLKMX2X2 U12295 ( .A(n5072), .B(\i_MIPS/Register/register[26][2] ), .S0(
        n5534), .Y(\i_MIPS/Register/n278 ) );
  CLKMX2X2 U12296 ( .A(n5037), .B(\i_MIPS/Register/register[27][20] ), .S0(
        n5531), .Y(\i_MIPS/Register/n264 ) );
  CLKMX2X2 U12297 ( .A(n5007), .B(\i_MIPS/Register/register[27][4] ), .S0(
        n5531), .Y(\i_MIPS/Register/n248 ) );
  CLKMX2X2 U12298 ( .A(n5037), .B(\i_MIPS/Register/register[28][20] ), .S0(
        n5529), .Y(\i_MIPS/Register/n232 ) );
  CLKMX2X2 U12299 ( .A(n5006), .B(\i_MIPS/Register/register[28][4] ), .S0(
        n5529), .Y(\i_MIPS/Register/n216 ) );
  CLKMX2X2 U12300 ( .A(n5072), .B(\i_MIPS/Register/register[28][2] ), .S0(
        n5530), .Y(\i_MIPS/Register/n214 ) );
  CLKMX2X2 U12301 ( .A(n5036), .B(\i_MIPS/Register/register[29][20] ), .S0(
        n5527), .Y(\i_MIPS/Register/n200 ) );
  CLKMX2X2 U12302 ( .A(n5007), .B(\i_MIPS/Register/register[29][4] ), .S0(
        n5527), .Y(\i_MIPS/Register/n184 ) );
  CLKMX2X2 U12303 ( .A(n5037), .B(\i_MIPS/Register/register[30][20] ), .S0(
        n5525), .Y(\i_MIPS/Register/n168 ) );
  CLKMX2X2 U12304 ( .A(n5007), .B(\i_MIPS/Register/register[30][4] ), .S0(
        n5525), .Y(\i_MIPS/Register/n152 ) );
  CLKMX2X2 U12305 ( .A(n5072), .B(\i_MIPS/Register/register[30][2] ), .S0(
        n5526), .Y(\i_MIPS/Register/n150 ) );
  CLKMX2X2 U12306 ( .A(n5065), .B(\i_MIPS/Register/register[0][30] ), .S0(
        n5586), .Y(\i_MIPS/Register/n1138 ) );
  CLKMX2X2 U12307 ( .A(n5033), .B(\i_MIPS/Register/register[0][29] ), .S0(
        n5585), .Y(\i_MIPS/Register/n1137 ) );
  CLKMX2X2 U12308 ( .A(n5012), .B(\i_MIPS/Register/register[0][28] ), .S0(
        n5585), .Y(\i_MIPS/Register/n1136 ) );
  CLKMX2X2 U12309 ( .A(n5030), .B(\i_MIPS/Register/register[0][27] ), .S0(
        n5585), .Y(\i_MIPS/Register/n1135 ) );
  CLKMX2X2 U12310 ( .A(n5015), .B(\i_MIPS/Register/register[0][26] ), .S0(
        n5585), .Y(\i_MIPS/Register/n1134 ) );
  CLKMX2X2 U12311 ( .A(n5021), .B(\i_MIPS/Register/register[0][25] ), .S0(
        n5585), .Y(\i_MIPS/Register/n1133 ) );
  CLKMX2X2 U12312 ( .A(n5048), .B(\i_MIPS/Register/register[0][24] ), .S0(
        n5586), .Y(\i_MIPS/Register/n1132 ) );
  CLKMX2X2 U12313 ( .A(n5045), .B(\i_MIPS/Register/register[0][23] ), .S0(
        n5586), .Y(\i_MIPS/Register/n1131 ) );
  CLKMX2X2 U12314 ( .A(n5042), .B(\i_MIPS/Register/register[0][22] ), .S0(
        n5586), .Y(\i_MIPS/Register/n1130 ) );
  CLKMX2X2 U12315 ( .A(n5039), .B(\i_MIPS/Register/register[0][21] ), .S0(
        n5586), .Y(\i_MIPS/Register/n1129 ) );
  CLKMX2X2 U12316 ( .A(n5009), .B(\i_MIPS/Register/register[0][19] ), .S0(
        n5585), .Y(\i_MIPS/Register/n1127 ) );
  CLKMX2X2 U12317 ( .A(n5057), .B(\i_MIPS/Register/register[0][18] ), .S0(
        n5586), .Y(\i_MIPS/Register/n1126 ) );
  CLKMX2X2 U12318 ( .A(n5054), .B(\i_MIPS/Register/register[0][17] ), .S0(
        n5586), .Y(\i_MIPS/Register/n1125 ) );
  CLKMX2X2 U12319 ( .A(n5027), .B(\i_MIPS/Register/register[0][16] ), .S0(
        n5585), .Y(\i_MIPS/Register/n1124 ) );
  CLKMX2X2 U12320 ( .A(n5018), .B(\i_MIPS/Register/register[0][15] ), .S0(
        n5585), .Y(\i_MIPS/Register/n1123 ) );
  CLKMX2X2 U12321 ( .A(n5024), .B(\i_MIPS/Register/register[0][14] ), .S0(
        n5585), .Y(\i_MIPS/Register/n1122 ) );
  CLKMX2X2 U12322 ( .A(n5080), .B(\i_MIPS/Register/register[0][11] ), .S0(
        n5586), .Y(\i_MIPS/Register/n1119 ) );
  CLKMX2X2 U12323 ( .A(n5051), .B(\i_MIPS/Register/register[0][10] ), .S0(
        n5586), .Y(\i_MIPS/Register/n1118 ) );
  CLKMX2X2 U12324 ( .A(n5077), .B(\i_MIPS/Register/register[0][9] ), .S0(n5586), .Y(\i_MIPS/Register/n1117 ) );
  CLKMX2X2 U12325 ( .A(n5068), .B(\i_MIPS/Register/register[0][7] ), .S0(n5586), .Y(\i_MIPS/Register/n1115 ) );
  CLKMX2X2 U12326 ( .A(net111835), .B(\i_MIPS/Register/register[0][6] ), .S0(
        n5585), .Y(\i_MIPS/Register/n1114 ) );
  CLKMX2X2 U12327 ( .A(n5075), .B(\i_MIPS/Register/register[0][5] ), .S0(n5586), .Y(\i_MIPS/Register/n1113 ) );
  CLKMX2X2 U12328 ( .A(n5003), .B(\i_MIPS/Register/register[0][3] ), .S0(n5585), .Y(\i_MIPS/Register/n1111 ) );
  CLKMX2X2 U12329 ( .A(n5500), .B(\i_MIPS/Register/register[1][31] ), .S0(
        n5583), .Y(\i_MIPS/Register/n1107 ) );
  CLKMX2X2 U12330 ( .A(n5065), .B(\i_MIPS/Register/register[1][30] ), .S0(
        n5584), .Y(\i_MIPS/Register/n1106 ) );
  CLKMX2X2 U12331 ( .A(n5033), .B(\i_MIPS/Register/register[1][29] ), .S0(
        n5584), .Y(\i_MIPS/Register/n1105 ) );
  CLKMX2X2 U12332 ( .A(n5012), .B(\i_MIPS/Register/register[1][28] ), .S0(
        n5583), .Y(\i_MIPS/Register/n1104 ) );
  CLKMX2X2 U12333 ( .A(n5030), .B(\i_MIPS/Register/register[1][27] ), .S0(
        n5584), .Y(\i_MIPS/Register/n1103 ) );
  CLKMX2X2 U12334 ( .A(n5015), .B(\i_MIPS/Register/register[1][26] ), .S0(
        n5583), .Y(\i_MIPS/Register/n1102 ) );
  CLKMX2X2 U12335 ( .A(n5021), .B(\i_MIPS/Register/register[1][25] ), .S0(
        n5583), .Y(\i_MIPS/Register/n1101 ) );
  CLKMX2X2 U12336 ( .A(n5048), .B(\i_MIPS/Register/register[1][24] ), .S0(
        n5584), .Y(\i_MIPS/Register/n1100 ) );
  CLKMX2X2 U12337 ( .A(n5045), .B(\i_MIPS/Register/register[1][23] ), .S0(
        n5584), .Y(\i_MIPS/Register/n1099 ) );
  CLKMX2X2 U12338 ( .A(n5042), .B(\i_MIPS/Register/register[1][22] ), .S0(
        n5584), .Y(\i_MIPS/Register/n1098 ) );
  CLKMX2X2 U12339 ( .A(n5039), .B(\i_MIPS/Register/register[1][21] ), .S0(
        n5584), .Y(\i_MIPS/Register/n1097 ) );
  CLKMX2X2 U12340 ( .A(n5009), .B(\i_MIPS/Register/register[1][19] ), .S0(
        n5583), .Y(\i_MIPS/Register/n1095 ) );
  CLKMX2X2 U12341 ( .A(n5057), .B(\i_MIPS/Register/register[1][18] ), .S0(
        n5584), .Y(\i_MIPS/Register/n1094 ) );
  CLKMX2X2 U12342 ( .A(n5054), .B(\i_MIPS/Register/register[1][17] ), .S0(
        n5584), .Y(\i_MIPS/Register/n1093 ) );
  CLKMX2X2 U12343 ( .A(n5027), .B(\i_MIPS/Register/register[1][16] ), .S0(
        n5583), .Y(\i_MIPS/Register/n1092 ) );
  CLKMX2X2 U12344 ( .A(n5018), .B(\i_MIPS/Register/register[1][15] ), .S0(
        n5583), .Y(\i_MIPS/Register/n1091 ) );
  CLKMX2X2 U12345 ( .A(n5024), .B(\i_MIPS/Register/register[1][14] ), .S0(
        n5583), .Y(\i_MIPS/Register/n1090 ) );
  CLKMX2X2 U12346 ( .A(n5051), .B(\i_MIPS/Register/register[1][10] ), .S0(
        n5584), .Y(\i_MIPS/Register/n1086 ) );
  CLKMX2X2 U12347 ( .A(n5077), .B(\i_MIPS/Register/register[1][9] ), .S0(n5584), .Y(\i_MIPS/Register/n1085 ) );
  CLKMX2X2 U12348 ( .A(n5068), .B(\i_MIPS/Register/register[1][7] ), .S0(n5584), .Y(\i_MIPS/Register/n1083 ) );
  CLKMX2X2 U12349 ( .A(net111835), .B(\i_MIPS/Register/register[1][6] ), .S0(
        n5583), .Y(\i_MIPS/Register/n1082 ) );
  CLKMX2X2 U12350 ( .A(n5074), .B(\i_MIPS/Register/register[1][5] ), .S0(n5583), .Y(\i_MIPS/Register/n1081 ) );
  CLKMX2X2 U12351 ( .A(n5003), .B(\i_MIPS/Register/register[1][3] ), .S0(n5583), .Y(\i_MIPS/Register/n1079 ) );
  CLKMX2X2 U12352 ( .A(n5500), .B(\i_MIPS/Register/register[2][31] ), .S0(
        n5581), .Y(\i_MIPS/Register/n1075 ) );
  CLKMX2X2 U12353 ( .A(n5065), .B(\i_MIPS/Register/register[2][30] ), .S0(
        n5582), .Y(\i_MIPS/Register/n1074 ) );
  CLKMX2X2 U12354 ( .A(n5033), .B(\i_MIPS/Register/register[2][29] ), .S0(
        n5582), .Y(\i_MIPS/Register/n1073 ) );
  CLKMX2X2 U12355 ( .A(n5012), .B(\i_MIPS/Register/register[2][28] ), .S0(
        n5581), .Y(\i_MIPS/Register/n1072 ) );
  CLKMX2X2 U12356 ( .A(n5030), .B(\i_MIPS/Register/register[2][27] ), .S0(
        n5582), .Y(\i_MIPS/Register/n1071 ) );
  CLKMX2X2 U12357 ( .A(n5015), .B(\i_MIPS/Register/register[2][26] ), .S0(
        n5581), .Y(\i_MIPS/Register/n1070 ) );
  CLKMX2X2 U12358 ( .A(n5021), .B(\i_MIPS/Register/register[2][25] ), .S0(
        n5581), .Y(\i_MIPS/Register/n1069 ) );
  CLKMX2X2 U12359 ( .A(n5048), .B(\i_MIPS/Register/register[2][24] ), .S0(
        n5582), .Y(\i_MIPS/Register/n1068 ) );
  CLKMX2X2 U12360 ( .A(n5045), .B(\i_MIPS/Register/register[2][23] ), .S0(
        n5582), .Y(\i_MIPS/Register/n1067 ) );
  CLKMX2X2 U12361 ( .A(n5042), .B(\i_MIPS/Register/register[2][22] ), .S0(
        n5582), .Y(\i_MIPS/Register/n1066 ) );
  CLKMX2X2 U12362 ( .A(n5039), .B(\i_MIPS/Register/register[2][21] ), .S0(
        n5582), .Y(\i_MIPS/Register/n1065 ) );
  CLKMX2X2 U12363 ( .A(n5009), .B(\i_MIPS/Register/register[2][19] ), .S0(
        n5581), .Y(\i_MIPS/Register/n1063 ) );
  CLKMX2X2 U12364 ( .A(n5057), .B(\i_MIPS/Register/register[2][18] ), .S0(
        n5582), .Y(\i_MIPS/Register/n1062 ) );
  CLKMX2X2 U12365 ( .A(n5054), .B(\i_MIPS/Register/register[2][17] ), .S0(
        n5582), .Y(\i_MIPS/Register/n1061 ) );
  CLKMX2X2 U12366 ( .A(n5027), .B(\i_MIPS/Register/register[2][16] ), .S0(
        n5581), .Y(\i_MIPS/Register/n1060 ) );
  CLKMX2X2 U12367 ( .A(n5018), .B(\i_MIPS/Register/register[2][15] ), .S0(
        n5581), .Y(\i_MIPS/Register/n1059 ) );
  CLKMX2X2 U12368 ( .A(n5024), .B(\i_MIPS/Register/register[2][14] ), .S0(
        n5581), .Y(\i_MIPS/Register/n1058 ) );
  CLKMX2X2 U12369 ( .A(n5051), .B(\i_MIPS/Register/register[2][10] ), .S0(
        n5582), .Y(\i_MIPS/Register/n1054 ) );
  CLKMX2X2 U12370 ( .A(n5077), .B(\i_MIPS/Register/register[2][9] ), .S0(n5582), .Y(\i_MIPS/Register/n1053 ) );
  CLKMX2X2 U12371 ( .A(n5068), .B(\i_MIPS/Register/register[2][7] ), .S0(n5582), .Y(\i_MIPS/Register/n1051 ) );
  CLKMX2X2 U12372 ( .A(net111835), .B(\i_MIPS/Register/register[2][6] ), .S0(
        n5581), .Y(\i_MIPS/Register/n1050 ) );
  CLKMX2X2 U12373 ( .A(n5074), .B(\i_MIPS/Register/register[2][5] ), .S0(n5581), .Y(\i_MIPS/Register/n1049 ) );
  CLKMX2X2 U12374 ( .A(n5003), .B(\i_MIPS/Register/register[2][3] ), .S0(n5581), .Y(\i_MIPS/Register/n1047 ) );
  CLKMX2X2 U12375 ( .A(n5500), .B(\i_MIPS/Register/register[3][31] ), .S0(
        n5579), .Y(\i_MIPS/Register/n1043 ) );
  CLKMX2X2 U12376 ( .A(n5065), .B(\i_MIPS/Register/register[3][30] ), .S0(
        n5580), .Y(\i_MIPS/Register/n1042 ) );
  CLKMX2X2 U12377 ( .A(n5033), .B(\i_MIPS/Register/register[3][29] ), .S0(
        n5580), .Y(\i_MIPS/Register/n1041 ) );
  CLKMX2X2 U12378 ( .A(n5012), .B(\i_MIPS/Register/register[3][28] ), .S0(
        n5579), .Y(\i_MIPS/Register/n1040 ) );
  CLKMX2X2 U12379 ( .A(n5030), .B(\i_MIPS/Register/register[3][27] ), .S0(
        n5580), .Y(\i_MIPS/Register/n1039 ) );
  CLKMX2X2 U12380 ( .A(n5015), .B(\i_MIPS/Register/register[3][26] ), .S0(
        n5579), .Y(\i_MIPS/Register/n1038 ) );
  CLKMX2X2 U12381 ( .A(n5021), .B(\i_MIPS/Register/register[3][25] ), .S0(
        n5579), .Y(\i_MIPS/Register/n1037 ) );
  CLKMX2X2 U12382 ( .A(n5048), .B(\i_MIPS/Register/register[3][24] ), .S0(
        n5580), .Y(\i_MIPS/Register/n1036 ) );
  CLKMX2X2 U12383 ( .A(n5045), .B(\i_MIPS/Register/register[3][23] ), .S0(
        n5580), .Y(\i_MIPS/Register/n1035 ) );
  CLKMX2X2 U12384 ( .A(n5042), .B(\i_MIPS/Register/register[3][22] ), .S0(
        n5580), .Y(\i_MIPS/Register/n1034 ) );
  CLKMX2X2 U12385 ( .A(n5039), .B(\i_MIPS/Register/register[3][21] ), .S0(
        n5580), .Y(\i_MIPS/Register/n1033 ) );
  CLKMX2X2 U12386 ( .A(n5009), .B(\i_MIPS/Register/register[3][19] ), .S0(
        n5579), .Y(\i_MIPS/Register/n1031 ) );
  CLKMX2X2 U12387 ( .A(n5057), .B(\i_MIPS/Register/register[3][18] ), .S0(
        n5580), .Y(\i_MIPS/Register/n1030 ) );
  CLKMX2X2 U12388 ( .A(n5054), .B(\i_MIPS/Register/register[3][17] ), .S0(
        n5580), .Y(\i_MIPS/Register/n1029 ) );
  CLKMX2X2 U12389 ( .A(n5027), .B(\i_MIPS/Register/register[3][16] ), .S0(
        n5579), .Y(\i_MIPS/Register/n1028 ) );
  CLKMX2X2 U12390 ( .A(n5018), .B(\i_MIPS/Register/register[3][15] ), .S0(
        n5579), .Y(\i_MIPS/Register/n1027 ) );
  CLKMX2X2 U12391 ( .A(n5024), .B(\i_MIPS/Register/register[3][14] ), .S0(
        n5579), .Y(\i_MIPS/Register/n1026 ) );
  CLKMX2X2 U12392 ( .A(n5051), .B(\i_MIPS/Register/register[3][10] ), .S0(
        n5580), .Y(\i_MIPS/Register/n1022 ) );
  CLKMX2X2 U12393 ( .A(n5077), .B(\i_MIPS/Register/register[3][9] ), .S0(n5580), .Y(\i_MIPS/Register/n1021 ) );
  CLKMX2X2 U12394 ( .A(n5068), .B(\i_MIPS/Register/register[3][7] ), .S0(n5580), .Y(\i_MIPS/Register/n1019 ) );
  CLKMX2X2 U12395 ( .A(net111835), .B(\i_MIPS/Register/register[3][6] ), .S0(
        n5579), .Y(\i_MIPS/Register/n1018 ) );
  CLKMX2X2 U12396 ( .A(n5074), .B(\i_MIPS/Register/register[3][5] ), .S0(n5579), .Y(\i_MIPS/Register/n1017 ) );
  CLKMX2X2 U12397 ( .A(n5003), .B(\i_MIPS/Register/register[3][3] ), .S0(n5579), .Y(\i_MIPS/Register/n1015 ) );
  CLKMX2X2 U12398 ( .A(n5500), .B(\i_MIPS/Register/register[4][31] ), .S0(
        n5577), .Y(\i_MIPS/Register/n1011 ) );
  CLKMX2X2 U12399 ( .A(n5065), .B(\i_MIPS/Register/register[4][30] ), .S0(
        n5578), .Y(\i_MIPS/Register/n1010 ) );
  CLKMX2X2 U12400 ( .A(n5033), .B(\i_MIPS/Register/register[4][29] ), .S0(
        n5578), .Y(\i_MIPS/Register/n1009 ) );
  CLKMX2X2 U12401 ( .A(n5012), .B(\i_MIPS/Register/register[4][28] ), .S0(
        n5577), .Y(\i_MIPS/Register/n1008 ) );
  CLKMX2X2 U12402 ( .A(n5030), .B(\i_MIPS/Register/register[4][27] ), .S0(
        n5578), .Y(\i_MIPS/Register/n1007 ) );
  CLKMX2X2 U12403 ( .A(n5015), .B(\i_MIPS/Register/register[4][26] ), .S0(
        n5577), .Y(\i_MIPS/Register/n1006 ) );
  CLKMX2X2 U12404 ( .A(n5021), .B(\i_MIPS/Register/register[4][25] ), .S0(
        n5577), .Y(\i_MIPS/Register/n1005 ) );
  CLKMX2X2 U12405 ( .A(n5048), .B(\i_MIPS/Register/register[4][24] ), .S0(
        n5578), .Y(\i_MIPS/Register/n1004 ) );
  CLKMX2X2 U12406 ( .A(n5045), .B(\i_MIPS/Register/register[4][23] ), .S0(
        n5578), .Y(\i_MIPS/Register/n1003 ) );
  CLKMX2X2 U12407 ( .A(n5042), .B(\i_MIPS/Register/register[4][22] ), .S0(
        n5578), .Y(\i_MIPS/Register/n1002 ) );
  CLKMX2X2 U12408 ( .A(n5039), .B(\i_MIPS/Register/register[4][21] ), .S0(
        n5578), .Y(\i_MIPS/Register/n1001 ) );
  CLKMX2X2 U12409 ( .A(n5009), .B(\i_MIPS/Register/register[4][19] ), .S0(
        n5577), .Y(\i_MIPS/Register/n999 ) );
  CLKMX2X2 U12410 ( .A(n5057), .B(\i_MIPS/Register/register[4][18] ), .S0(
        n5578), .Y(\i_MIPS/Register/n998 ) );
  CLKMX2X2 U12411 ( .A(n5054), .B(\i_MIPS/Register/register[4][17] ), .S0(
        n5578), .Y(\i_MIPS/Register/n997 ) );
  CLKMX2X2 U12412 ( .A(n5027), .B(\i_MIPS/Register/register[4][16] ), .S0(
        n5577), .Y(\i_MIPS/Register/n996 ) );
  CLKMX2X2 U12413 ( .A(n5018), .B(\i_MIPS/Register/register[4][15] ), .S0(
        n5577), .Y(\i_MIPS/Register/n995 ) );
  CLKMX2X2 U12414 ( .A(n5024), .B(\i_MIPS/Register/register[4][14] ), .S0(
        n5577), .Y(\i_MIPS/Register/n994 ) );
  CLKMX2X2 U12415 ( .A(n5051), .B(\i_MIPS/Register/register[4][10] ), .S0(
        n5578), .Y(\i_MIPS/Register/n990 ) );
  CLKMX2X2 U12416 ( .A(n5077), .B(\i_MIPS/Register/register[4][9] ), .S0(n5578), .Y(\i_MIPS/Register/n989 ) );
  CLKMX2X2 U12417 ( .A(n5068), .B(\i_MIPS/Register/register[4][7] ), .S0(n5578), .Y(\i_MIPS/Register/n987 ) );
  CLKMX2X2 U12418 ( .A(net111835), .B(\i_MIPS/Register/register[4][6] ), .S0(
        n5577), .Y(\i_MIPS/Register/n986 ) );
  CLKMX2X2 U12419 ( .A(n5074), .B(\i_MIPS/Register/register[4][5] ), .S0(n5577), .Y(\i_MIPS/Register/n985 ) );
  CLKMX2X2 U12420 ( .A(n5003), .B(\i_MIPS/Register/register[4][3] ), .S0(n5577), .Y(\i_MIPS/Register/n983 ) );
  CLKMX2X2 U12421 ( .A(n5500), .B(\i_MIPS/Register/register[5][31] ), .S0(
        n5575), .Y(\i_MIPS/Register/n979 ) );
  CLKMX2X2 U12422 ( .A(n5065), .B(\i_MIPS/Register/register[5][30] ), .S0(
        n5576), .Y(\i_MIPS/Register/n978 ) );
  CLKMX2X2 U12423 ( .A(n5033), .B(\i_MIPS/Register/register[5][29] ), .S0(
        n5576), .Y(\i_MIPS/Register/n977 ) );
  CLKMX2X2 U12424 ( .A(n5012), .B(\i_MIPS/Register/register[5][28] ), .S0(
        n5575), .Y(\i_MIPS/Register/n976 ) );
  CLKMX2X2 U12425 ( .A(n5030), .B(\i_MIPS/Register/register[5][27] ), .S0(
        n5576), .Y(\i_MIPS/Register/n975 ) );
  CLKMX2X2 U12426 ( .A(n5015), .B(\i_MIPS/Register/register[5][26] ), .S0(
        n5575), .Y(\i_MIPS/Register/n974 ) );
  CLKMX2X2 U12427 ( .A(n5021), .B(\i_MIPS/Register/register[5][25] ), .S0(
        n5575), .Y(\i_MIPS/Register/n973 ) );
  CLKMX2X2 U12428 ( .A(n5048), .B(\i_MIPS/Register/register[5][24] ), .S0(
        n5576), .Y(\i_MIPS/Register/n972 ) );
  CLKMX2X2 U12429 ( .A(n5045), .B(\i_MIPS/Register/register[5][23] ), .S0(
        n5576), .Y(\i_MIPS/Register/n971 ) );
  CLKMX2X2 U12430 ( .A(n5042), .B(\i_MIPS/Register/register[5][22] ), .S0(
        n5576), .Y(\i_MIPS/Register/n970 ) );
  CLKMX2X2 U12431 ( .A(n5039), .B(\i_MIPS/Register/register[5][21] ), .S0(
        n5576), .Y(\i_MIPS/Register/n969 ) );
  CLKMX2X2 U12432 ( .A(n5009), .B(\i_MIPS/Register/register[5][19] ), .S0(
        n5575), .Y(\i_MIPS/Register/n967 ) );
  CLKMX2X2 U12433 ( .A(n5057), .B(\i_MIPS/Register/register[5][18] ), .S0(
        n5576), .Y(\i_MIPS/Register/n966 ) );
  CLKMX2X2 U12434 ( .A(n5054), .B(\i_MIPS/Register/register[5][17] ), .S0(
        n5576), .Y(\i_MIPS/Register/n965 ) );
  CLKMX2X2 U12435 ( .A(n5027), .B(\i_MIPS/Register/register[5][16] ), .S0(
        n5575), .Y(\i_MIPS/Register/n964 ) );
  CLKMX2X2 U12436 ( .A(n5018), .B(\i_MIPS/Register/register[5][15] ), .S0(
        n5575), .Y(\i_MIPS/Register/n963 ) );
  CLKMX2X2 U12437 ( .A(n5024), .B(\i_MIPS/Register/register[5][14] ), .S0(
        n5575), .Y(\i_MIPS/Register/n962 ) );
  CLKMX2X2 U12438 ( .A(n5051), .B(\i_MIPS/Register/register[5][10] ), .S0(
        n5576), .Y(\i_MIPS/Register/n958 ) );
  CLKMX2X2 U12439 ( .A(n5077), .B(\i_MIPS/Register/register[5][9] ), .S0(n5576), .Y(\i_MIPS/Register/n957 ) );
  CLKMX2X2 U12440 ( .A(n5068), .B(\i_MIPS/Register/register[5][7] ), .S0(n5576), .Y(\i_MIPS/Register/n955 ) );
  CLKMX2X2 U12441 ( .A(net111835), .B(\i_MIPS/Register/register[5][6] ), .S0(
        n5575), .Y(\i_MIPS/Register/n954 ) );
  CLKMX2X2 U12442 ( .A(n5074), .B(\i_MIPS/Register/register[5][5] ), .S0(n5575), .Y(\i_MIPS/Register/n953 ) );
  CLKMX2X2 U12443 ( .A(n5003), .B(\i_MIPS/Register/register[5][3] ), .S0(n5575), .Y(\i_MIPS/Register/n951 ) );
  CLKMX2X2 U12444 ( .A(n5500), .B(\i_MIPS/Register/register[6][31] ), .S0(
        n5573), .Y(\i_MIPS/Register/n947 ) );
  CLKMX2X2 U12445 ( .A(n5065), .B(\i_MIPS/Register/register[6][30] ), .S0(
        n5574), .Y(\i_MIPS/Register/n946 ) );
  CLKMX2X2 U12446 ( .A(n5033), .B(\i_MIPS/Register/register[6][29] ), .S0(
        n5574), .Y(\i_MIPS/Register/n945 ) );
  CLKMX2X2 U12447 ( .A(n5012), .B(\i_MIPS/Register/register[6][28] ), .S0(
        n5573), .Y(\i_MIPS/Register/n944 ) );
  CLKMX2X2 U12448 ( .A(n5030), .B(\i_MIPS/Register/register[6][27] ), .S0(
        n5574), .Y(\i_MIPS/Register/n943 ) );
  CLKMX2X2 U12449 ( .A(n5015), .B(\i_MIPS/Register/register[6][26] ), .S0(
        n5573), .Y(\i_MIPS/Register/n942 ) );
  CLKMX2X2 U12450 ( .A(n5021), .B(\i_MIPS/Register/register[6][25] ), .S0(
        n5573), .Y(\i_MIPS/Register/n941 ) );
  CLKMX2X2 U12451 ( .A(n5048), .B(\i_MIPS/Register/register[6][24] ), .S0(
        n5574), .Y(\i_MIPS/Register/n940 ) );
  CLKMX2X2 U12452 ( .A(n5045), .B(\i_MIPS/Register/register[6][23] ), .S0(
        n5574), .Y(\i_MIPS/Register/n939 ) );
  CLKMX2X2 U12453 ( .A(n5042), .B(\i_MIPS/Register/register[6][22] ), .S0(
        n5574), .Y(\i_MIPS/Register/n938 ) );
  CLKMX2X2 U12454 ( .A(n5039), .B(\i_MIPS/Register/register[6][21] ), .S0(
        n5574), .Y(\i_MIPS/Register/n937 ) );
  CLKMX2X2 U12455 ( .A(n5009), .B(\i_MIPS/Register/register[6][19] ), .S0(
        n5573), .Y(\i_MIPS/Register/n935 ) );
  CLKMX2X2 U12456 ( .A(n5057), .B(\i_MIPS/Register/register[6][18] ), .S0(
        n5574), .Y(\i_MIPS/Register/n934 ) );
  CLKMX2X2 U12457 ( .A(n5054), .B(\i_MIPS/Register/register[6][17] ), .S0(
        n5574), .Y(\i_MIPS/Register/n933 ) );
  CLKMX2X2 U12458 ( .A(n5027), .B(\i_MIPS/Register/register[6][16] ), .S0(
        n5573), .Y(\i_MIPS/Register/n932 ) );
  CLKMX2X2 U12459 ( .A(n5018), .B(\i_MIPS/Register/register[6][15] ), .S0(
        n5573), .Y(\i_MIPS/Register/n931 ) );
  CLKMX2X2 U12460 ( .A(n5024), .B(\i_MIPS/Register/register[6][14] ), .S0(
        n5573), .Y(\i_MIPS/Register/n930 ) );
  CLKMX2X2 U12461 ( .A(n5051), .B(\i_MIPS/Register/register[6][10] ), .S0(
        n5574), .Y(\i_MIPS/Register/n926 ) );
  CLKMX2X2 U12462 ( .A(n5077), .B(\i_MIPS/Register/register[6][9] ), .S0(n5574), .Y(\i_MIPS/Register/n925 ) );
  CLKMX2X2 U12463 ( .A(n5068), .B(\i_MIPS/Register/register[6][7] ), .S0(n5574), .Y(\i_MIPS/Register/n923 ) );
  CLKMX2X2 U12464 ( .A(net111835), .B(\i_MIPS/Register/register[6][6] ), .S0(
        n5573), .Y(\i_MIPS/Register/n922 ) );
  CLKMX2X2 U12465 ( .A(n5074), .B(\i_MIPS/Register/register[6][5] ), .S0(n5573), .Y(\i_MIPS/Register/n921 ) );
  CLKMX2X2 U12466 ( .A(n5003), .B(\i_MIPS/Register/register[6][3] ), .S0(n5573), .Y(\i_MIPS/Register/n919 ) );
  CLKMX2X2 U12467 ( .A(n5500), .B(\i_MIPS/Register/register[7][31] ), .S0(
        n5571), .Y(\i_MIPS/Register/n915 ) );
  CLKMX2X2 U12468 ( .A(n5066), .B(\i_MIPS/Register/register[7][30] ), .S0(
        n5572), .Y(\i_MIPS/Register/n914 ) );
  CLKMX2X2 U12469 ( .A(n5034), .B(\i_MIPS/Register/register[7][29] ), .S0(
        n5572), .Y(\i_MIPS/Register/n913 ) );
  CLKMX2X2 U12470 ( .A(n5013), .B(\i_MIPS/Register/register[7][28] ), .S0(
        n5571), .Y(\i_MIPS/Register/n912 ) );
  CLKMX2X2 U12471 ( .A(n5031), .B(\i_MIPS/Register/register[7][27] ), .S0(
        n5572), .Y(\i_MIPS/Register/n911 ) );
  CLKMX2X2 U12472 ( .A(n5016), .B(\i_MIPS/Register/register[7][26] ), .S0(
        n5571), .Y(\i_MIPS/Register/n910 ) );
  CLKMX2X2 U12473 ( .A(n5022), .B(\i_MIPS/Register/register[7][25] ), .S0(
        n5571), .Y(\i_MIPS/Register/n909 ) );
  CLKMX2X2 U12474 ( .A(n5049), .B(\i_MIPS/Register/register[7][24] ), .S0(
        n5572), .Y(\i_MIPS/Register/n908 ) );
  CLKMX2X2 U12475 ( .A(n5046), .B(\i_MIPS/Register/register[7][23] ), .S0(
        n5572), .Y(\i_MIPS/Register/n907 ) );
  CLKMX2X2 U12476 ( .A(n5043), .B(\i_MIPS/Register/register[7][22] ), .S0(
        n5572), .Y(\i_MIPS/Register/n906 ) );
  CLKMX2X2 U12477 ( .A(n5040), .B(\i_MIPS/Register/register[7][21] ), .S0(
        n5572), .Y(\i_MIPS/Register/n905 ) );
  CLKMX2X2 U12478 ( .A(n5010), .B(\i_MIPS/Register/register[7][19] ), .S0(
        n5571), .Y(\i_MIPS/Register/n903 ) );
  CLKMX2X2 U12479 ( .A(n5058), .B(\i_MIPS/Register/register[7][18] ), .S0(
        n5572), .Y(\i_MIPS/Register/n902 ) );
  CLKMX2X2 U12480 ( .A(n5055), .B(\i_MIPS/Register/register[7][17] ), .S0(
        n5572), .Y(\i_MIPS/Register/n901 ) );
  CLKMX2X2 U12481 ( .A(n5028), .B(\i_MIPS/Register/register[7][16] ), .S0(
        n5571), .Y(\i_MIPS/Register/n900 ) );
  CLKMX2X2 U12482 ( .A(n5019), .B(\i_MIPS/Register/register[7][15] ), .S0(
        n5571), .Y(\i_MIPS/Register/n899 ) );
  CLKMX2X2 U12483 ( .A(n5025), .B(\i_MIPS/Register/register[7][14] ), .S0(
        n5571), .Y(\i_MIPS/Register/n898 ) );
  CLKMX2X2 U12484 ( .A(n5052), .B(\i_MIPS/Register/register[7][10] ), .S0(
        n5572), .Y(\i_MIPS/Register/n894 ) );
  CLKMX2X2 U12485 ( .A(n5078), .B(\i_MIPS/Register/register[7][9] ), .S0(n5572), .Y(\i_MIPS/Register/n893 ) );
  CLKMX2X2 U12486 ( .A(n5069), .B(\i_MIPS/Register/register[7][7] ), .S0(n5572), .Y(\i_MIPS/Register/n891 ) );
  CLKMX2X2 U12487 ( .A(net111837), .B(\i_MIPS/Register/register[7][6] ), .S0(
        n5571), .Y(\i_MIPS/Register/n890 ) );
  CLKMX2X2 U12488 ( .A(n5074), .B(\i_MIPS/Register/register[7][5] ), .S0(n5571), .Y(\i_MIPS/Register/n889 ) );
  CLKMX2X2 U12489 ( .A(n5004), .B(\i_MIPS/Register/register[7][3] ), .S0(n5571), .Y(\i_MIPS/Register/n887 ) );
  CLKMX2X2 U12490 ( .A(n5500), .B(\i_MIPS/Register/register[8][31] ), .S0(
        n5569), .Y(\i_MIPS/Register/n883 ) );
  CLKMX2X2 U12491 ( .A(n5065), .B(\i_MIPS/Register/register[8][30] ), .S0(
        n5570), .Y(\i_MIPS/Register/n882 ) );
  CLKMX2X2 U12492 ( .A(n5033), .B(\i_MIPS/Register/register[8][29] ), .S0(
        n5570), .Y(\i_MIPS/Register/n881 ) );
  CLKMX2X2 U12493 ( .A(n5012), .B(\i_MIPS/Register/register[8][28] ), .S0(
        n5569), .Y(\i_MIPS/Register/n880 ) );
  CLKMX2X2 U12494 ( .A(n5030), .B(\i_MIPS/Register/register[8][27] ), .S0(
        n5570), .Y(\i_MIPS/Register/n879 ) );
  CLKMX2X2 U12495 ( .A(n5015), .B(\i_MIPS/Register/register[8][26] ), .S0(
        n5569), .Y(\i_MIPS/Register/n878 ) );
  CLKMX2X2 U12496 ( .A(n5021), .B(\i_MIPS/Register/register[8][25] ), .S0(
        n5569), .Y(\i_MIPS/Register/n877 ) );
  CLKMX2X2 U12497 ( .A(n5048), .B(\i_MIPS/Register/register[8][24] ), .S0(
        n5570), .Y(\i_MIPS/Register/n876 ) );
  CLKMX2X2 U12498 ( .A(n5045), .B(\i_MIPS/Register/register[8][23] ), .S0(
        n5570), .Y(\i_MIPS/Register/n875 ) );
  CLKMX2X2 U12499 ( .A(n5042), .B(\i_MIPS/Register/register[8][22] ), .S0(
        n5570), .Y(\i_MIPS/Register/n874 ) );
  CLKMX2X2 U12500 ( .A(n5039), .B(\i_MIPS/Register/register[8][21] ), .S0(
        n5570), .Y(\i_MIPS/Register/n873 ) );
  CLKMX2X2 U12501 ( .A(n5009), .B(\i_MIPS/Register/register[8][19] ), .S0(
        n5569), .Y(\i_MIPS/Register/n871 ) );
  CLKMX2X2 U12502 ( .A(n5057), .B(\i_MIPS/Register/register[8][18] ), .S0(
        n5570), .Y(\i_MIPS/Register/n870 ) );
  CLKMX2X2 U12503 ( .A(n5054), .B(\i_MIPS/Register/register[8][17] ), .S0(
        n5570), .Y(\i_MIPS/Register/n869 ) );
  CLKMX2X2 U12504 ( .A(n5027), .B(\i_MIPS/Register/register[8][16] ), .S0(
        n5569), .Y(\i_MIPS/Register/n868 ) );
  CLKMX2X2 U12505 ( .A(n5018), .B(\i_MIPS/Register/register[8][15] ), .S0(
        n5569), .Y(\i_MIPS/Register/n867 ) );
  CLKMX2X2 U12506 ( .A(n5024), .B(\i_MIPS/Register/register[8][14] ), .S0(
        n5569), .Y(\i_MIPS/Register/n866 ) );
  CLKMX2X2 U12507 ( .A(n5051), .B(\i_MIPS/Register/register[8][10] ), .S0(
        n5570), .Y(\i_MIPS/Register/n862 ) );
  CLKMX2X2 U12508 ( .A(n5077), .B(\i_MIPS/Register/register[8][9] ), .S0(n5570), .Y(\i_MIPS/Register/n861 ) );
  CLKMX2X2 U12509 ( .A(n5068), .B(\i_MIPS/Register/register[8][7] ), .S0(n5570), .Y(\i_MIPS/Register/n859 ) );
  CLKMX2X2 U12510 ( .A(net111835), .B(\i_MIPS/Register/register[8][6] ), .S0(
        n5569), .Y(\i_MIPS/Register/n858 ) );
  CLKMX2X2 U12511 ( .A(n5074), .B(\i_MIPS/Register/register[8][5] ), .S0(n5569), .Y(\i_MIPS/Register/n857 ) );
  CLKMX2X2 U12512 ( .A(n5003), .B(\i_MIPS/Register/register[8][3] ), .S0(n5569), .Y(\i_MIPS/Register/n855 ) );
  CLKMX2X2 U12513 ( .A(n5500), .B(\i_MIPS/Register/register[9][31] ), .S0(
        n5567), .Y(\i_MIPS/Register/n851 ) );
  CLKMX2X2 U12514 ( .A(n5065), .B(\i_MIPS/Register/register[9][30] ), .S0(
        n5568), .Y(\i_MIPS/Register/n850 ) );
  CLKMX2X2 U12515 ( .A(n5033), .B(\i_MIPS/Register/register[9][29] ), .S0(
        n5568), .Y(\i_MIPS/Register/n849 ) );
  CLKMX2X2 U12516 ( .A(n5012), .B(\i_MIPS/Register/register[9][28] ), .S0(
        n5567), .Y(\i_MIPS/Register/n848 ) );
  CLKMX2X2 U12517 ( .A(n5030), .B(\i_MIPS/Register/register[9][27] ), .S0(
        n5568), .Y(\i_MIPS/Register/n847 ) );
  CLKMX2X2 U12518 ( .A(n5015), .B(\i_MIPS/Register/register[9][26] ), .S0(
        n5567), .Y(\i_MIPS/Register/n846 ) );
  CLKMX2X2 U12519 ( .A(n5021), .B(\i_MIPS/Register/register[9][25] ), .S0(
        n5567), .Y(\i_MIPS/Register/n845 ) );
  CLKMX2X2 U12520 ( .A(n5048), .B(\i_MIPS/Register/register[9][24] ), .S0(
        n5568), .Y(\i_MIPS/Register/n844 ) );
  CLKMX2X2 U12521 ( .A(n5045), .B(\i_MIPS/Register/register[9][23] ), .S0(
        n5568), .Y(\i_MIPS/Register/n843 ) );
  CLKMX2X2 U12522 ( .A(n5042), .B(\i_MIPS/Register/register[9][22] ), .S0(
        n5568), .Y(\i_MIPS/Register/n842 ) );
  CLKMX2X2 U12523 ( .A(n5039), .B(\i_MIPS/Register/register[9][21] ), .S0(
        n5568), .Y(\i_MIPS/Register/n841 ) );
  CLKMX2X2 U12524 ( .A(n5009), .B(\i_MIPS/Register/register[9][19] ), .S0(
        n5567), .Y(\i_MIPS/Register/n839 ) );
  CLKMX2X2 U12525 ( .A(n5057), .B(\i_MIPS/Register/register[9][18] ), .S0(
        n5568), .Y(\i_MIPS/Register/n838 ) );
  CLKMX2X2 U12526 ( .A(n5054), .B(\i_MIPS/Register/register[9][17] ), .S0(
        n5568), .Y(\i_MIPS/Register/n837 ) );
  CLKMX2X2 U12527 ( .A(n5027), .B(\i_MIPS/Register/register[9][16] ), .S0(
        n5567), .Y(\i_MIPS/Register/n836 ) );
  CLKMX2X2 U12528 ( .A(n5018), .B(\i_MIPS/Register/register[9][15] ), .S0(
        n5567), .Y(\i_MIPS/Register/n835 ) );
  CLKMX2X2 U12529 ( .A(n5024), .B(\i_MIPS/Register/register[9][14] ), .S0(
        n5567), .Y(\i_MIPS/Register/n834 ) );
  CLKMX2X2 U12530 ( .A(n5051), .B(\i_MIPS/Register/register[9][10] ), .S0(
        n5568), .Y(\i_MIPS/Register/n830 ) );
  CLKMX2X2 U12531 ( .A(n5077), .B(\i_MIPS/Register/register[9][9] ), .S0(n5568), .Y(\i_MIPS/Register/n829 ) );
  CLKMX2X2 U12532 ( .A(n5068), .B(\i_MIPS/Register/register[9][7] ), .S0(n5568), .Y(\i_MIPS/Register/n827 ) );
  CLKMX2X2 U12533 ( .A(net111835), .B(\i_MIPS/Register/register[9][6] ), .S0(
        n5567), .Y(\i_MIPS/Register/n826 ) );
  CLKMX2X2 U12534 ( .A(n5074), .B(\i_MIPS/Register/register[9][5] ), .S0(n5567), .Y(\i_MIPS/Register/n825 ) );
  CLKMX2X2 U12535 ( .A(n5003), .B(\i_MIPS/Register/register[9][3] ), .S0(n5567), .Y(\i_MIPS/Register/n823 ) );
  CLKMX2X2 U12536 ( .A(n5500), .B(\i_MIPS/Register/register[10][31] ), .S0(
        n5565), .Y(\i_MIPS/Register/n819 ) );
  CLKMX2X2 U12537 ( .A(n5065), .B(\i_MIPS/Register/register[10][30] ), .S0(
        n5566), .Y(\i_MIPS/Register/n818 ) );
  CLKMX2X2 U12538 ( .A(n5033), .B(\i_MIPS/Register/register[10][29] ), .S0(
        n5566), .Y(\i_MIPS/Register/n817 ) );
  CLKMX2X2 U12539 ( .A(n5012), .B(\i_MIPS/Register/register[10][28] ), .S0(
        n5565), .Y(\i_MIPS/Register/n816 ) );
  CLKMX2X2 U12540 ( .A(n5030), .B(\i_MIPS/Register/register[10][27] ), .S0(
        n5566), .Y(\i_MIPS/Register/n815 ) );
  CLKMX2X2 U12541 ( .A(n5015), .B(\i_MIPS/Register/register[10][26] ), .S0(
        n5565), .Y(\i_MIPS/Register/n814 ) );
  CLKMX2X2 U12542 ( .A(n5021), .B(\i_MIPS/Register/register[10][25] ), .S0(
        n5565), .Y(\i_MIPS/Register/n813 ) );
  CLKMX2X2 U12543 ( .A(n5048), .B(\i_MIPS/Register/register[10][24] ), .S0(
        n5566), .Y(\i_MIPS/Register/n812 ) );
  CLKMX2X2 U12544 ( .A(n5045), .B(\i_MIPS/Register/register[10][23] ), .S0(
        n5566), .Y(\i_MIPS/Register/n811 ) );
  CLKMX2X2 U12545 ( .A(n5042), .B(\i_MIPS/Register/register[10][22] ), .S0(
        n5566), .Y(\i_MIPS/Register/n810 ) );
  CLKMX2X2 U12546 ( .A(n5039), .B(\i_MIPS/Register/register[10][21] ), .S0(
        n5566), .Y(\i_MIPS/Register/n809 ) );
  CLKMX2X2 U12547 ( .A(n5009), .B(\i_MIPS/Register/register[10][19] ), .S0(
        n5565), .Y(\i_MIPS/Register/n807 ) );
  CLKMX2X2 U12548 ( .A(n5057), .B(\i_MIPS/Register/register[10][18] ), .S0(
        n5566), .Y(\i_MIPS/Register/n806 ) );
  CLKMX2X2 U12549 ( .A(n5054), .B(\i_MIPS/Register/register[10][17] ), .S0(
        n5566), .Y(\i_MIPS/Register/n805 ) );
  CLKMX2X2 U12550 ( .A(n5027), .B(\i_MIPS/Register/register[10][16] ), .S0(
        n5565), .Y(\i_MIPS/Register/n804 ) );
  CLKMX2X2 U12551 ( .A(n5018), .B(\i_MIPS/Register/register[10][15] ), .S0(
        n5565), .Y(\i_MIPS/Register/n803 ) );
  CLKMX2X2 U12552 ( .A(n5024), .B(\i_MIPS/Register/register[10][14] ), .S0(
        n5565), .Y(\i_MIPS/Register/n802 ) );
  CLKMX2X2 U12553 ( .A(n5051), .B(\i_MIPS/Register/register[10][10] ), .S0(
        n5566), .Y(\i_MIPS/Register/n798 ) );
  CLKMX2X2 U12554 ( .A(n5077), .B(\i_MIPS/Register/register[10][9] ), .S0(
        n5566), .Y(\i_MIPS/Register/n797 ) );
  CLKMX2X2 U12555 ( .A(n5068), .B(\i_MIPS/Register/register[10][7] ), .S0(
        n5566), .Y(\i_MIPS/Register/n795 ) );
  CLKMX2X2 U12556 ( .A(net111835), .B(\i_MIPS/Register/register[10][6] ), .S0(
        n5565), .Y(\i_MIPS/Register/n794 ) );
  CLKMX2X2 U12557 ( .A(n5074), .B(\i_MIPS/Register/register[10][5] ), .S0(
        n5565), .Y(\i_MIPS/Register/n793 ) );
  CLKMX2X2 U12558 ( .A(n5003), .B(\i_MIPS/Register/register[10][3] ), .S0(
        n5565), .Y(\i_MIPS/Register/n791 ) );
  CLKMX2X2 U12559 ( .A(n5500), .B(\i_MIPS/Register/register[11][31] ), .S0(
        n5563), .Y(\i_MIPS/Register/n787 ) );
  CLKMX2X2 U12560 ( .A(n5066), .B(\i_MIPS/Register/register[11][30] ), .S0(
        n5564), .Y(\i_MIPS/Register/n786 ) );
  CLKMX2X2 U12561 ( .A(n5034), .B(\i_MIPS/Register/register[11][29] ), .S0(
        n5564), .Y(\i_MIPS/Register/n785 ) );
  CLKMX2X2 U12562 ( .A(n5013), .B(\i_MIPS/Register/register[11][28] ), .S0(
        n5563), .Y(\i_MIPS/Register/n784 ) );
  CLKMX2X2 U12563 ( .A(n5031), .B(\i_MIPS/Register/register[11][27] ), .S0(
        n5564), .Y(\i_MIPS/Register/n783 ) );
  CLKMX2X2 U12564 ( .A(n5016), .B(\i_MIPS/Register/register[11][26] ), .S0(
        n5563), .Y(\i_MIPS/Register/n782 ) );
  CLKMX2X2 U12565 ( .A(n5022), .B(\i_MIPS/Register/register[11][25] ), .S0(
        n5563), .Y(\i_MIPS/Register/n781 ) );
  CLKMX2X2 U12566 ( .A(n5049), .B(\i_MIPS/Register/register[11][24] ), .S0(
        n5564), .Y(\i_MIPS/Register/n780 ) );
  CLKMX2X2 U12567 ( .A(n5046), .B(\i_MIPS/Register/register[11][23] ), .S0(
        n5564), .Y(\i_MIPS/Register/n779 ) );
  CLKMX2X2 U12568 ( .A(n5043), .B(\i_MIPS/Register/register[11][22] ), .S0(
        n5564), .Y(\i_MIPS/Register/n778 ) );
  CLKMX2X2 U12569 ( .A(n5040), .B(\i_MIPS/Register/register[11][21] ), .S0(
        n5564), .Y(\i_MIPS/Register/n777 ) );
  CLKMX2X2 U12570 ( .A(n5010), .B(\i_MIPS/Register/register[11][19] ), .S0(
        n5563), .Y(\i_MIPS/Register/n775 ) );
  CLKMX2X2 U12571 ( .A(n5058), .B(\i_MIPS/Register/register[11][18] ), .S0(
        n5564), .Y(\i_MIPS/Register/n774 ) );
  CLKMX2X2 U12572 ( .A(n5055), .B(\i_MIPS/Register/register[11][17] ), .S0(
        n5564), .Y(\i_MIPS/Register/n773 ) );
  CLKMX2X2 U12573 ( .A(n5028), .B(\i_MIPS/Register/register[11][16] ), .S0(
        n5563), .Y(\i_MIPS/Register/n772 ) );
  CLKMX2X2 U12574 ( .A(n5018), .B(\i_MIPS/Register/register[11][15] ), .S0(
        n5563), .Y(\i_MIPS/Register/n771 ) );
  CLKMX2X2 U12575 ( .A(n5025), .B(\i_MIPS/Register/register[11][14] ), .S0(
        n5563), .Y(\i_MIPS/Register/n770 ) );
  CLKMX2X2 U12576 ( .A(n5052), .B(\i_MIPS/Register/register[11][10] ), .S0(
        n5564), .Y(\i_MIPS/Register/n766 ) );
  CLKMX2X2 U12577 ( .A(n5078), .B(\i_MIPS/Register/register[11][9] ), .S0(
        n5564), .Y(\i_MIPS/Register/n765 ) );
  CLKMX2X2 U12578 ( .A(n5069), .B(\i_MIPS/Register/register[11][7] ), .S0(
        n5564), .Y(\i_MIPS/Register/n763 ) );
  CLKMX2X2 U12579 ( .A(net111837), .B(\i_MIPS/Register/register[11][6] ), .S0(
        n5563), .Y(\i_MIPS/Register/n762 ) );
  CLKMX2X2 U12580 ( .A(n5074), .B(\i_MIPS/Register/register[11][5] ), .S0(
        n5563), .Y(\i_MIPS/Register/n761 ) );
  CLKMX2X2 U12581 ( .A(n5004), .B(\i_MIPS/Register/register[11][3] ), .S0(
        n5563), .Y(\i_MIPS/Register/n759 ) );
  CLKMX2X2 U12582 ( .A(n5500), .B(\i_MIPS/Register/register[12][31] ), .S0(
        n5561), .Y(\i_MIPS/Register/n755 ) );
  CLKMX2X2 U12583 ( .A(n5065), .B(\i_MIPS/Register/register[12][30] ), .S0(
        n5562), .Y(\i_MIPS/Register/n754 ) );
  CLKMX2X2 U12584 ( .A(n5033), .B(\i_MIPS/Register/register[12][29] ), .S0(
        n5562), .Y(\i_MIPS/Register/n753 ) );
  CLKMX2X2 U12585 ( .A(n5012), .B(\i_MIPS/Register/register[12][28] ), .S0(
        n5561), .Y(\i_MIPS/Register/n752 ) );
  CLKMX2X2 U12586 ( .A(n5030), .B(\i_MIPS/Register/register[12][27] ), .S0(
        n5562), .Y(\i_MIPS/Register/n751 ) );
  CLKMX2X2 U12587 ( .A(n5015), .B(\i_MIPS/Register/register[12][26] ), .S0(
        n5561), .Y(\i_MIPS/Register/n750 ) );
  CLKMX2X2 U12588 ( .A(n5021), .B(\i_MIPS/Register/register[12][25] ), .S0(
        n5561), .Y(\i_MIPS/Register/n749 ) );
  CLKMX2X2 U12589 ( .A(n5048), .B(\i_MIPS/Register/register[12][24] ), .S0(
        n5562), .Y(\i_MIPS/Register/n748 ) );
  CLKMX2X2 U12590 ( .A(n5045), .B(\i_MIPS/Register/register[12][23] ), .S0(
        n5562), .Y(\i_MIPS/Register/n747 ) );
  CLKMX2X2 U12591 ( .A(n5042), .B(\i_MIPS/Register/register[12][22] ), .S0(
        n5562), .Y(\i_MIPS/Register/n746 ) );
  CLKMX2X2 U12592 ( .A(n5039), .B(\i_MIPS/Register/register[12][21] ), .S0(
        n5562), .Y(\i_MIPS/Register/n745 ) );
  CLKMX2X2 U12593 ( .A(n5009), .B(\i_MIPS/Register/register[12][19] ), .S0(
        n5561), .Y(\i_MIPS/Register/n743 ) );
  CLKMX2X2 U12594 ( .A(n5057), .B(\i_MIPS/Register/register[12][18] ), .S0(
        n5562), .Y(\i_MIPS/Register/n742 ) );
  CLKMX2X2 U12595 ( .A(n5054), .B(\i_MIPS/Register/register[12][17] ), .S0(
        n5562), .Y(\i_MIPS/Register/n741 ) );
  CLKMX2X2 U12596 ( .A(n5027), .B(\i_MIPS/Register/register[12][16] ), .S0(
        n5561), .Y(\i_MIPS/Register/n740 ) );
  CLKMX2X2 U12597 ( .A(n5018), .B(\i_MIPS/Register/register[12][15] ), .S0(
        n5561), .Y(\i_MIPS/Register/n739 ) );
  CLKMX2X2 U12598 ( .A(n5024), .B(\i_MIPS/Register/register[12][14] ), .S0(
        n5561), .Y(\i_MIPS/Register/n738 ) );
  CLKMX2X2 U12599 ( .A(n5051), .B(\i_MIPS/Register/register[12][10] ), .S0(
        n5562), .Y(\i_MIPS/Register/n734 ) );
  CLKMX2X2 U12600 ( .A(n5077), .B(\i_MIPS/Register/register[12][9] ), .S0(
        n5562), .Y(\i_MIPS/Register/n733 ) );
  CLKMX2X2 U12601 ( .A(n5068), .B(\i_MIPS/Register/register[12][7] ), .S0(
        n5562), .Y(\i_MIPS/Register/n731 ) );
  CLKMX2X2 U12602 ( .A(net111835), .B(\i_MIPS/Register/register[12][6] ), .S0(
        n5561), .Y(\i_MIPS/Register/n730 ) );
  CLKMX2X2 U12603 ( .A(n5074), .B(\i_MIPS/Register/register[12][5] ), .S0(
        n5561), .Y(\i_MIPS/Register/n729 ) );
  CLKMX2X2 U12604 ( .A(n5003), .B(\i_MIPS/Register/register[12][3] ), .S0(
        n5561), .Y(\i_MIPS/Register/n727 ) );
  CLKMX2X2 U12605 ( .A(n5500), .B(\i_MIPS/Register/register[13][31] ), .S0(
        n5559), .Y(\i_MIPS/Register/n723 ) );
  CLKMX2X2 U12606 ( .A(n5065), .B(\i_MIPS/Register/register[13][30] ), .S0(
        n5560), .Y(\i_MIPS/Register/n722 ) );
  CLKMX2X2 U12607 ( .A(n5033), .B(\i_MIPS/Register/register[13][29] ), .S0(
        n5560), .Y(\i_MIPS/Register/n721 ) );
  CLKMX2X2 U12608 ( .A(n5012), .B(\i_MIPS/Register/register[13][28] ), .S0(
        n5559), .Y(\i_MIPS/Register/n720 ) );
  CLKMX2X2 U12609 ( .A(n5030), .B(\i_MIPS/Register/register[13][27] ), .S0(
        n5560), .Y(\i_MIPS/Register/n719 ) );
  CLKMX2X2 U12610 ( .A(n5015), .B(\i_MIPS/Register/register[13][26] ), .S0(
        n5559), .Y(\i_MIPS/Register/n718 ) );
  CLKMX2X2 U12611 ( .A(n5021), .B(\i_MIPS/Register/register[13][25] ), .S0(
        n5559), .Y(\i_MIPS/Register/n717 ) );
  CLKMX2X2 U12612 ( .A(n5048), .B(\i_MIPS/Register/register[13][24] ), .S0(
        n5560), .Y(\i_MIPS/Register/n716 ) );
  CLKMX2X2 U12613 ( .A(n5045), .B(\i_MIPS/Register/register[13][23] ), .S0(
        n5560), .Y(\i_MIPS/Register/n715 ) );
  CLKMX2X2 U12614 ( .A(n5042), .B(\i_MIPS/Register/register[13][22] ), .S0(
        n5560), .Y(\i_MIPS/Register/n714 ) );
  CLKMX2X2 U12615 ( .A(n5039), .B(\i_MIPS/Register/register[13][21] ), .S0(
        n5560), .Y(\i_MIPS/Register/n713 ) );
  CLKMX2X2 U12616 ( .A(n5009), .B(\i_MIPS/Register/register[13][19] ), .S0(
        n5559), .Y(\i_MIPS/Register/n711 ) );
  CLKMX2X2 U12617 ( .A(n5057), .B(\i_MIPS/Register/register[13][18] ), .S0(
        n5560), .Y(\i_MIPS/Register/n710 ) );
  CLKMX2X2 U12618 ( .A(n5054), .B(\i_MIPS/Register/register[13][17] ), .S0(
        n5560), .Y(\i_MIPS/Register/n709 ) );
  CLKMX2X2 U12619 ( .A(n5027), .B(\i_MIPS/Register/register[13][16] ), .S0(
        n5559), .Y(\i_MIPS/Register/n708 ) );
  CLKMX2X2 U12620 ( .A(n5018), .B(\i_MIPS/Register/register[13][15] ), .S0(
        n5559), .Y(\i_MIPS/Register/n707 ) );
  CLKMX2X2 U12621 ( .A(n5024), .B(\i_MIPS/Register/register[13][14] ), .S0(
        n5559), .Y(\i_MIPS/Register/n706 ) );
  CLKMX2X2 U12622 ( .A(n5051), .B(\i_MIPS/Register/register[13][10] ), .S0(
        n5560), .Y(\i_MIPS/Register/n702 ) );
  CLKMX2X2 U12623 ( .A(n5077), .B(\i_MIPS/Register/register[13][9] ), .S0(
        n5560), .Y(\i_MIPS/Register/n701 ) );
  CLKMX2X2 U12624 ( .A(n5068), .B(\i_MIPS/Register/register[13][7] ), .S0(
        n5560), .Y(\i_MIPS/Register/n699 ) );
  CLKMX2X2 U12625 ( .A(net111835), .B(\i_MIPS/Register/register[13][6] ), .S0(
        n5559), .Y(\i_MIPS/Register/n698 ) );
  CLKMX2X2 U12626 ( .A(n5074), .B(\i_MIPS/Register/register[13][5] ), .S0(
        n5559), .Y(\i_MIPS/Register/n697 ) );
  CLKMX2X2 U12627 ( .A(n5003), .B(\i_MIPS/Register/register[13][3] ), .S0(
        n5559), .Y(\i_MIPS/Register/n695 ) );
  CLKMX2X2 U12628 ( .A(n5500), .B(\i_MIPS/Register/register[14][31] ), .S0(
        n5557), .Y(\i_MIPS/Register/n691 ) );
  CLKMX2X2 U12629 ( .A(n5065), .B(\i_MIPS/Register/register[14][30] ), .S0(
        n5558), .Y(\i_MIPS/Register/n690 ) );
  CLKMX2X2 U12630 ( .A(n5033), .B(\i_MIPS/Register/register[14][29] ), .S0(
        n5558), .Y(\i_MIPS/Register/n689 ) );
  CLKMX2X2 U12631 ( .A(n5012), .B(\i_MIPS/Register/register[14][28] ), .S0(
        n5557), .Y(\i_MIPS/Register/n688 ) );
  CLKMX2X2 U12632 ( .A(n5030), .B(\i_MIPS/Register/register[14][27] ), .S0(
        n5558), .Y(\i_MIPS/Register/n687 ) );
  CLKMX2X2 U12633 ( .A(n5015), .B(\i_MIPS/Register/register[14][26] ), .S0(
        n5557), .Y(\i_MIPS/Register/n686 ) );
  CLKMX2X2 U12634 ( .A(n5021), .B(\i_MIPS/Register/register[14][25] ), .S0(
        n5557), .Y(\i_MIPS/Register/n685 ) );
  CLKMX2X2 U12635 ( .A(n5048), .B(\i_MIPS/Register/register[14][24] ), .S0(
        n5558), .Y(\i_MIPS/Register/n684 ) );
  CLKMX2X2 U12636 ( .A(n5045), .B(\i_MIPS/Register/register[14][23] ), .S0(
        n5558), .Y(\i_MIPS/Register/n683 ) );
  CLKMX2X2 U12637 ( .A(n5042), .B(\i_MIPS/Register/register[14][22] ), .S0(
        n5558), .Y(\i_MIPS/Register/n682 ) );
  CLKMX2X2 U12638 ( .A(n5039), .B(\i_MIPS/Register/register[14][21] ), .S0(
        n5558), .Y(\i_MIPS/Register/n681 ) );
  CLKMX2X2 U12639 ( .A(n5009), .B(\i_MIPS/Register/register[14][19] ), .S0(
        n5557), .Y(\i_MIPS/Register/n679 ) );
  CLKMX2X2 U12640 ( .A(n5057), .B(\i_MIPS/Register/register[14][18] ), .S0(
        n5558), .Y(\i_MIPS/Register/n678 ) );
  CLKMX2X2 U12641 ( .A(n5054), .B(\i_MIPS/Register/register[14][17] ), .S0(
        n5558), .Y(\i_MIPS/Register/n677 ) );
  CLKMX2X2 U12642 ( .A(n5027), .B(\i_MIPS/Register/register[14][16] ), .S0(
        n5557), .Y(\i_MIPS/Register/n676 ) );
  CLKMX2X2 U12643 ( .A(n5018), .B(\i_MIPS/Register/register[14][15] ), .S0(
        n5557), .Y(\i_MIPS/Register/n675 ) );
  CLKMX2X2 U12644 ( .A(n5024), .B(\i_MIPS/Register/register[14][14] ), .S0(
        n5557), .Y(\i_MIPS/Register/n674 ) );
  CLKMX2X2 U12645 ( .A(n5051), .B(\i_MIPS/Register/register[14][10] ), .S0(
        n5558), .Y(\i_MIPS/Register/n670 ) );
  CLKMX2X2 U12646 ( .A(n5077), .B(\i_MIPS/Register/register[14][9] ), .S0(
        n5558), .Y(\i_MIPS/Register/n669 ) );
  CLKMX2X2 U12647 ( .A(n5068), .B(\i_MIPS/Register/register[14][7] ), .S0(
        n5558), .Y(\i_MIPS/Register/n667 ) );
  CLKMX2X2 U12648 ( .A(net111835), .B(\i_MIPS/Register/register[14][6] ), .S0(
        n5557), .Y(\i_MIPS/Register/n666 ) );
  CLKMX2X2 U12649 ( .A(n5074), .B(\i_MIPS/Register/register[14][5] ), .S0(
        n5557), .Y(\i_MIPS/Register/n665 ) );
  CLKMX2X2 U12650 ( .A(n5003), .B(\i_MIPS/Register/register[14][3] ), .S0(
        n5557), .Y(\i_MIPS/Register/n663 ) );
  CLKMX2X2 U12651 ( .A(n11217), .B(\i_MIPS/Register/register[15][31] ), .S0(
        n5555), .Y(\i_MIPS/Register/n659 ) );
  CLKMX2X2 U12652 ( .A(n5066), .B(\i_MIPS/Register/register[15][30] ), .S0(
        n5556), .Y(\i_MIPS/Register/n658 ) );
  CLKMX2X2 U12653 ( .A(n5034), .B(\i_MIPS/Register/register[15][29] ), .S0(
        n5556), .Y(\i_MIPS/Register/n657 ) );
  CLKMX2X2 U12654 ( .A(n5013), .B(\i_MIPS/Register/register[15][28] ), .S0(
        n5555), .Y(\i_MIPS/Register/n656 ) );
  CLKMX2X2 U12655 ( .A(n5031), .B(\i_MIPS/Register/register[15][27] ), .S0(
        n5556), .Y(\i_MIPS/Register/n655 ) );
  CLKMX2X2 U12656 ( .A(n5016), .B(\i_MIPS/Register/register[15][26] ), .S0(
        n5555), .Y(\i_MIPS/Register/n654 ) );
  CLKMX2X2 U12657 ( .A(n5022), .B(\i_MIPS/Register/register[15][25] ), .S0(
        n5555), .Y(\i_MIPS/Register/n653 ) );
  CLKMX2X2 U12658 ( .A(n5049), .B(\i_MIPS/Register/register[15][24] ), .S0(
        n5556), .Y(\i_MIPS/Register/n652 ) );
  CLKMX2X2 U12659 ( .A(n5046), .B(\i_MIPS/Register/register[15][23] ), .S0(
        n5556), .Y(\i_MIPS/Register/n651 ) );
  CLKMX2X2 U12660 ( .A(n5043), .B(\i_MIPS/Register/register[15][22] ), .S0(
        n5556), .Y(\i_MIPS/Register/n650 ) );
  CLKMX2X2 U12661 ( .A(n5040), .B(\i_MIPS/Register/register[15][21] ), .S0(
        n5556), .Y(\i_MIPS/Register/n649 ) );
  CLKMX2X2 U12662 ( .A(n5010), .B(\i_MIPS/Register/register[15][19] ), .S0(
        n5555), .Y(\i_MIPS/Register/n647 ) );
  CLKMX2X2 U12663 ( .A(n5058), .B(\i_MIPS/Register/register[15][18] ), .S0(
        n5556), .Y(\i_MIPS/Register/n646 ) );
  CLKMX2X2 U12664 ( .A(n5055), .B(\i_MIPS/Register/register[15][17] ), .S0(
        n5556), .Y(\i_MIPS/Register/n645 ) );
  CLKMX2X2 U12665 ( .A(n5028), .B(\i_MIPS/Register/register[15][16] ), .S0(
        n5555), .Y(\i_MIPS/Register/n644 ) );
  CLKMX2X2 U12666 ( .A(n5019), .B(\i_MIPS/Register/register[15][15] ), .S0(
        n5555), .Y(\i_MIPS/Register/n643 ) );
  CLKMX2X2 U12667 ( .A(n5025), .B(\i_MIPS/Register/register[15][14] ), .S0(
        n5555), .Y(\i_MIPS/Register/n642 ) );
  CLKMX2X2 U12668 ( .A(n5052), .B(\i_MIPS/Register/register[15][10] ), .S0(
        n5556), .Y(\i_MIPS/Register/n638 ) );
  CLKMX2X2 U12669 ( .A(n5078), .B(\i_MIPS/Register/register[15][9] ), .S0(
        n5556), .Y(\i_MIPS/Register/n637 ) );
  CLKMX2X2 U12670 ( .A(n5069), .B(\i_MIPS/Register/register[15][7] ), .S0(
        n5556), .Y(\i_MIPS/Register/n635 ) );
  CLKMX2X2 U12671 ( .A(net111837), .B(\i_MIPS/Register/register[15][6] ), .S0(
        n5555), .Y(\i_MIPS/Register/n634 ) );
  CLKMX2X2 U12672 ( .A(n5074), .B(\i_MIPS/Register/register[15][5] ), .S0(
        n5555), .Y(\i_MIPS/Register/n633 ) );
  CLKMX2X2 U12673 ( .A(n5004), .B(\i_MIPS/Register/register[15][3] ), .S0(
        n5555), .Y(\i_MIPS/Register/n631 ) );
  CLKMX2X2 U12674 ( .A(n11217), .B(\i_MIPS/Register/register[16][31] ), .S0(
        n5553), .Y(\i_MIPS/Register/n627 ) );
  CLKMX2X2 U12675 ( .A(n5066), .B(\i_MIPS/Register/register[16][30] ), .S0(
        n5554), .Y(\i_MIPS/Register/n626 ) );
  CLKMX2X2 U12676 ( .A(n5034), .B(\i_MIPS/Register/register[16][29] ), .S0(
        n5554), .Y(\i_MIPS/Register/n625 ) );
  CLKMX2X2 U12677 ( .A(n5013), .B(\i_MIPS/Register/register[16][28] ), .S0(
        n5553), .Y(\i_MIPS/Register/n624 ) );
  CLKMX2X2 U12678 ( .A(n5031), .B(\i_MIPS/Register/register[16][27] ), .S0(
        n5554), .Y(\i_MIPS/Register/n623 ) );
  CLKMX2X2 U12679 ( .A(n5016), .B(\i_MIPS/Register/register[16][26] ), .S0(
        n5553), .Y(\i_MIPS/Register/n622 ) );
  CLKMX2X2 U12680 ( .A(n5022), .B(\i_MIPS/Register/register[16][25] ), .S0(
        n5553), .Y(\i_MIPS/Register/n621 ) );
  CLKMX2X2 U12681 ( .A(n5049), .B(\i_MIPS/Register/register[16][24] ), .S0(
        n5554), .Y(\i_MIPS/Register/n620 ) );
  CLKMX2X2 U12682 ( .A(n5046), .B(\i_MIPS/Register/register[16][23] ), .S0(
        n5554), .Y(\i_MIPS/Register/n619 ) );
  CLKMX2X2 U12683 ( .A(n5043), .B(\i_MIPS/Register/register[16][22] ), .S0(
        n5554), .Y(\i_MIPS/Register/n618 ) );
  CLKMX2X2 U12684 ( .A(n5040), .B(\i_MIPS/Register/register[16][21] ), .S0(
        n5554), .Y(\i_MIPS/Register/n617 ) );
  CLKMX2X2 U12685 ( .A(n5010), .B(\i_MIPS/Register/register[16][19] ), .S0(
        n5553), .Y(\i_MIPS/Register/n615 ) );
  CLKMX2X2 U12686 ( .A(n5058), .B(\i_MIPS/Register/register[16][18] ), .S0(
        n5554), .Y(\i_MIPS/Register/n614 ) );
  CLKMX2X2 U12687 ( .A(n5055), .B(\i_MIPS/Register/register[16][17] ), .S0(
        n5554), .Y(\i_MIPS/Register/n613 ) );
  CLKMX2X2 U12688 ( .A(n5028), .B(\i_MIPS/Register/register[16][16] ), .S0(
        n5553), .Y(\i_MIPS/Register/n612 ) );
  CLKMX2X2 U12689 ( .A(n5019), .B(\i_MIPS/Register/register[16][15] ), .S0(
        n5553), .Y(\i_MIPS/Register/n611 ) );
  CLKMX2X2 U12690 ( .A(n5025), .B(\i_MIPS/Register/register[16][14] ), .S0(
        n5553), .Y(\i_MIPS/Register/n610 ) );
  CLKMX2X2 U12691 ( .A(n5052), .B(\i_MIPS/Register/register[16][10] ), .S0(
        n5554), .Y(\i_MIPS/Register/n606 ) );
  CLKMX2X2 U12692 ( .A(n5078), .B(\i_MIPS/Register/register[16][9] ), .S0(
        n5554), .Y(\i_MIPS/Register/n605 ) );
  CLKMX2X2 U12693 ( .A(n5069), .B(\i_MIPS/Register/register[16][7] ), .S0(
        n5554), .Y(\i_MIPS/Register/n603 ) );
  CLKMX2X2 U12694 ( .A(net111837), .B(\i_MIPS/Register/register[16][6] ), .S0(
        n5553), .Y(\i_MIPS/Register/n602 ) );
  CLKMX2X2 U12695 ( .A(n5074), .B(\i_MIPS/Register/register[16][5] ), .S0(
        n5553), .Y(\i_MIPS/Register/n601 ) );
  CLKMX2X2 U12696 ( .A(n5004), .B(\i_MIPS/Register/register[16][3] ), .S0(
        n5553), .Y(\i_MIPS/Register/n599 ) );
  CLKMX2X2 U12697 ( .A(n11217), .B(\i_MIPS/Register/register[17][31] ), .S0(
        n5551), .Y(\i_MIPS/Register/n595 ) );
  CLKMX2X2 U12698 ( .A(n5066), .B(\i_MIPS/Register/register[17][30] ), .S0(
        n5552), .Y(\i_MIPS/Register/n594 ) );
  CLKMX2X2 U12699 ( .A(n5034), .B(\i_MIPS/Register/register[17][29] ), .S0(
        n5552), .Y(\i_MIPS/Register/n593 ) );
  CLKMX2X2 U12700 ( .A(n5013), .B(\i_MIPS/Register/register[17][28] ), .S0(
        n5551), .Y(\i_MIPS/Register/n592 ) );
  CLKMX2X2 U12701 ( .A(n5031), .B(\i_MIPS/Register/register[17][27] ), .S0(
        n5552), .Y(\i_MIPS/Register/n591 ) );
  CLKMX2X2 U12702 ( .A(n5016), .B(\i_MIPS/Register/register[17][26] ), .S0(
        n5551), .Y(\i_MIPS/Register/n590 ) );
  CLKMX2X2 U12703 ( .A(n5022), .B(\i_MIPS/Register/register[17][25] ), .S0(
        n5551), .Y(\i_MIPS/Register/n589 ) );
  CLKMX2X2 U12704 ( .A(n5049), .B(\i_MIPS/Register/register[17][24] ), .S0(
        n5552), .Y(\i_MIPS/Register/n588 ) );
  CLKMX2X2 U12705 ( .A(n5046), .B(\i_MIPS/Register/register[17][23] ), .S0(
        n5552), .Y(\i_MIPS/Register/n587 ) );
  CLKMX2X2 U12706 ( .A(n5043), .B(\i_MIPS/Register/register[17][22] ), .S0(
        n5552), .Y(\i_MIPS/Register/n586 ) );
  CLKMX2X2 U12707 ( .A(n5040), .B(\i_MIPS/Register/register[17][21] ), .S0(
        n5552), .Y(\i_MIPS/Register/n585 ) );
  CLKMX2X2 U12708 ( .A(n5010), .B(\i_MIPS/Register/register[17][19] ), .S0(
        n5551), .Y(\i_MIPS/Register/n583 ) );
  CLKMX2X2 U12709 ( .A(n5058), .B(\i_MIPS/Register/register[17][18] ), .S0(
        n5552), .Y(\i_MIPS/Register/n582 ) );
  CLKMX2X2 U12710 ( .A(n5055), .B(\i_MIPS/Register/register[17][17] ), .S0(
        n5552), .Y(\i_MIPS/Register/n581 ) );
  CLKMX2X2 U12711 ( .A(n5028), .B(\i_MIPS/Register/register[17][16] ), .S0(
        n5551), .Y(\i_MIPS/Register/n580 ) );
  CLKMX2X2 U12712 ( .A(n5019), .B(\i_MIPS/Register/register[17][15] ), .S0(
        n5551), .Y(\i_MIPS/Register/n579 ) );
  CLKMX2X2 U12713 ( .A(n5025), .B(\i_MIPS/Register/register[17][14] ), .S0(
        n5551), .Y(\i_MIPS/Register/n578 ) );
  CLKMX2X2 U12714 ( .A(n5052), .B(\i_MIPS/Register/register[17][10] ), .S0(
        n5552), .Y(\i_MIPS/Register/n574 ) );
  CLKMX2X2 U12715 ( .A(n5078), .B(\i_MIPS/Register/register[17][9] ), .S0(
        n5552), .Y(\i_MIPS/Register/n573 ) );
  CLKMX2X2 U12716 ( .A(n5069), .B(\i_MIPS/Register/register[17][7] ), .S0(
        n5552), .Y(\i_MIPS/Register/n571 ) );
  CLKMX2X2 U12717 ( .A(net111837), .B(\i_MIPS/Register/register[17][6] ), .S0(
        n5551), .Y(\i_MIPS/Register/n570 ) );
  CLKMX2X2 U12718 ( .A(n5074), .B(\i_MIPS/Register/register[17][5] ), .S0(
        n5551), .Y(\i_MIPS/Register/n569 ) );
  CLKMX2X2 U12719 ( .A(n5004), .B(\i_MIPS/Register/register[17][3] ), .S0(
        n5551), .Y(\i_MIPS/Register/n567 ) );
  CLKMX2X2 U12720 ( .A(n11217), .B(\i_MIPS/Register/register[18][31] ), .S0(
        n5549), .Y(\i_MIPS/Register/n563 ) );
  CLKMX2X2 U12721 ( .A(n5066), .B(\i_MIPS/Register/register[18][30] ), .S0(
        n5550), .Y(\i_MIPS/Register/n562 ) );
  CLKMX2X2 U12722 ( .A(n5034), .B(\i_MIPS/Register/register[18][29] ), .S0(
        n5550), .Y(\i_MIPS/Register/n561 ) );
  CLKMX2X2 U12723 ( .A(n5013), .B(\i_MIPS/Register/register[18][28] ), .S0(
        n5549), .Y(\i_MIPS/Register/n560 ) );
  CLKMX2X2 U12724 ( .A(n5031), .B(\i_MIPS/Register/register[18][27] ), .S0(
        n5550), .Y(\i_MIPS/Register/n559 ) );
  CLKMX2X2 U12725 ( .A(n5016), .B(\i_MIPS/Register/register[18][26] ), .S0(
        n5549), .Y(\i_MIPS/Register/n558 ) );
  CLKMX2X2 U12726 ( .A(n5022), .B(\i_MIPS/Register/register[18][25] ), .S0(
        n5549), .Y(\i_MIPS/Register/n557 ) );
  CLKMX2X2 U12727 ( .A(n5049), .B(\i_MIPS/Register/register[18][24] ), .S0(
        n5550), .Y(\i_MIPS/Register/n556 ) );
  CLKMX2X2 U12728 ( .A(n5046), .B(\i_MIPS/Register/register[18][23] ), .S0(
        n5550), .Y(\i_MIPS/Register/n555 ) );
  CLKMX2X2 U12729 ( .A(n5043), .B(\i_MIPS/Register/register[18][22] ), .S0(
        n5550), .Y(\i_MIPS/Register/n554 ) );
  CLKMX2X2 U12730 ( .A(n5040), .B(\i_MIPS/Register/register[18][21] ), .S0(
        n5550), .Y(\i_MIPS/Register/n553 ) );
  CLKMX2X2 U12731 ( .A(n5010), .B(\i_MIPS/Register/register[18][19] ), .S0(
        n5549), .Y(\i_MIPS/Register/n551 ) );
  CLKMX2X2 U12732 ( .A(n5058), .B(\i_MIPS/Register/register[18][18] ), .S0(
        n5550), .Y(\i_MIPS/Register/n550 ) );
  CLKMX2X2 U12733 ( .A(n5055), .B(\i_MIPS/Register/register[18][17] ), .S0(
        n5550), .Y(\i_MIPS/Register/n549 ) );
  CLKMX2X2 U12734 ( .A(n5028), .B(\i_MIPS/Register/register[18][16] ), .S0(
        n5549), .Y(\i_MIPS/Register/n548 ) );
  CLKMX2X2 U12735 ( .A(n5019), .B(\i_MIPS/Register/register[18][15] ), .S0(
        n5549), .Y(\i_MIPS/Register/n547 ) );
  CLKMX2X2 U12736 ( .A(n5025), .B(\i_MIPS/Register/register[18][14] ), .S0(
        n5549), .Y(\i_MIPS/Register/n546 ) );
  CLKMX2X2 U12737 ( .A(n5052), .B(\i_MIPS/Register/register[18][10] ), .S0(
        n5550), .Y(\i_MIPS/Register/n542 ) );
  CLKMX2X2 U12738 ( .A(n5078), .B(\i_MIPS/Register/register[18][9] ), .S0(
        n5550), .Y(\i_MIPS/Register/n541 ) );
  CLKMX2X2 U12739 ( .A(n5069), .B(\i_MIPS/Register/register[18][7] ), .S0(
        n5550), .Y(\i_MIPS/Register/n539 ) );
  CLKMX2X2 U12740 ( .A(net111837), .B(\i_MIPS/Register/register[18][6] ), .S0(
        n5549), .Y(\i_MIPS/Register/n538 ) );
  CLKMX2X2 U12741 ( .A(n10764), .B(\i_MIPS/Register/register[18][5] ), .S0(
        n5549), .Y(\i_MIPS/Register/n537 ) );
  CLKMX2X2 U12742 ( .A(n5004), .B(\i_MIPS/Register/register[18][3] ), .S0(
        n5549), .Y(\i_MIPS/Register/n535 ) );
  CLKMX2X2 U12743 ( .A(n5500), .B(\i_MIPS/Register/register[19][31] ), .S0(
        n5547), .Y(\i_MIPS/Register/n531 ) );
  CLKMX2X2 U12744 ( .A(n5066), .B(\i_MIPS/Register/register[19][30] ), .S0(
        n5548), .Y(\i_MIPS/Register/n530 ) );
  CLKMX2X2 U12745 ( .A(n5033), .B(\i_MIPS/Register/register[19][29] ), .S0(
        n5548), .Y(\i_MIPS/Register/n529 ) );
  CLKMX2X2 U12746 ( .A(n5012), .B(\i_MIPS/Register/register[19][28] ), .S0(
        n5547), .Y(\i_MIPS/Register/n528 ) );
  CLKMX2X2 U12747 ( .A(n5030), .B(\i_MIPS/Register/register[19][27] ), .S0(
        n5548), .Y(\i_MIPS/Register/n527 ) );
  CLKMX2X2 U12748 ( .A(n5016), .B(\i_MIPS/Register/register[19][26] ), .S0(
        n5547), .Y(\i_MIPS/Register/n526 ) );
  CLKMX2X2 U12749 ( .A(n5021), .B(\i_MIPS/Register/register[19][25] ), .S0(
        n5547), .Y(\i_MIPS/Register/n525 ) );
  CLKMX2X2 U12750 ( .A(n5048), .B(\i_MIPS/Register/register[19][24] ), .S0(
        n5548), .Y(\i_MIPS/Register/n524 ) );
  CLKMX2X2 U12751 ( .A(n5045), .B(\i_MIPS/Register/register[19][23] ), .S0(
        n5548), .Y(\i_MIPS/Register/n523 ) );
  CLKMX2X2 U12752 ( .A(n5042), .B(\i_MIPS/Register/register[19][22] ), .S0(
        n5548), .Y(\i_MIPS/Register/n522 ) );
  CLKMX2X2 U12753 ( .A(n5040), .B(\i_MIPS/Register/register[19][21] ), .S0(
        n5548), .Y(\i_MIPS/Register/n521 ) );
  CLKMX2X2 U12754 ( .A(n5010), .B(\i_MIPS/Register/register[19][19] ), .S0(
        n5547), .Y(\i_MIPS/Register/n519 ) );
  CLKMX2X2 U12755 ( .A(n5058), .B(\i_MIPS/Register/register[19][18] ), .S0(
        n5548), .Y(\i_MIPS/Register/n518 ) );
  CLKMX2X2 U12756 ( .A(n5054), .B(\i_MIPS/Register/register[19][17] ), .S0(
        n5548), .Y(\i_MIPS/Register/n517 ) );
  CLKMX2X2 U12757 ( .A(n5027), .B(\i_MIPS/Register/register[19][16] ), .S0(
        n5547), .Y(\i_MIPS/Register/n516 ) );
  CLKMX2X2 U12758 ( .A(n5019), .B(\i_MIPS/Register/register[19][15] ), .S0(
        n5547), .Y(\i_MIPS/Register/n515 ) );
  CLKMX2X2 U12759 ( .A(n5024), .B(\i_MIPS/Register/register[19][14] ), .S0(
        n5547), .Y(\i_MIPS/Register/n514 ) );
  CLKMX2X2 U12760 ( .A(n5051), .B(\i_MIPS/Register/register[19][10] ), .S0(
        n5548), .Y(\i_MIPS/Register/n510 ) );
  CLKMX2X2 U12761 ( .A(n5077), .B(\i_MIPS/Register/register[19][9] ), .S0(
        n5548), .Y(\i_MIPS/Register/n509 ) );
  CLKMX2X2 U12762 ( .A(n5068), .B(\i_MIPS/Register/register[19][7] ), .S0(
        n5548), .Y(\i_MIPS/Register/n507 ) );
  CLKMX2X2 U12763 ( .A(net111835), .B(\i_MIPS/Register/register[19][6] ), .S0(
        n5547), .Y(\i_MIPS/Register/n506 ) );
  CLKMX2X2 U12764 ( .A(n5075), .B(\i_MIPS/Register/register[19][5] ), .S0(
        n5547), .Y(\i_MIPS/Register/n505 ) );
  CLKMX2X2 U12765 ( .A(n5003), .B(\i_MIPS/Register/register[19][3] ), .S0(
        n5547), .Y(\i_MIPS/Register/n503 ) );
  CLKMX2X2 U12766 ( .A(n5072), .B(\i_MIPS/Register/register[19][2] ), .S0(
        n5548), .Y(\i_MIPS/Register/n502 ) );
  CLKMX2X2 U12767 ( .A(n11217), .B(\i_MIPS/Register/register[20][31] ), .S0(
        n5545), .Y(\i_MIPS/Register/n499 ) );
  CLKMX2X2 U12768 ( .A(n5066), .B(\i_MIPS/Register/register[20][30] ), .S0(
        n5546), .Y(\i_MIPS/Register/n498 ) );
  CLKMX2X2 U12769 ( .A(n5034), .B(\i_MIPS/Register/register[20][29] ), .S0(
        n5546), .Y(\i_MIPS/Register/n497 ) );
  CLKMX2X2 U12770 ( .A(n5013), .B(\i_MIPS/Register/register[20][28] ), .S0(
        n5545), .Y(\i_MIPS/Register/n496 ) );
  CLKMX2X2 U12771 ( .A(n5031), .B(\i_MIPS/Register/register[20][27] ), .S0(
        n5546), .Y(\i_MIPS/Register/n495 ) );
  CLKMX2X2 U12772 ( .A(n5016), .B(\i_MIPS/Register/register[20][26] ), .S0(
        n5545), .Y(\i_MIPS/Register/n494 ) );
  CLKMX2X2 U12773 ( .A(n5022), .B(\i_MIPS/Register/register[20][25] ), .S0(
        n5545), .Y(\i_MIPS/Register/n493 ) );
  CLKMX2X2 U12774 ( .A(n5049), .B(\i_MIPS/Register/register[20][24] ), .S0(
        n5546), .Y(\i_MIPS/Register/n492 ) );
  CLKMX2X2 U12775 ( .A(n5046), .B(\i_MIPS/Register/register[20][23] ), .S0(
        n5546), .Y(\i_MIPS/Register/n491 ) );
  CLKMX2X2 U12776 ( .A(n5043), .B(\i_MIPS/Register/register[20][22] ), .S0(
        n5546), .Y(\i_MIPS/Register/n490 ) );
  CLKMX2X2 U12777 ( .A(n5040), .B(\i_MIPS/Register/register[20][21] ), .S0(
        n5546), .Y(\i_MIPS/Register/n489 ) );
  CLKMX2X2 U12778 ( .A(n5010), .B(\i_MIPS/Register/register[20][19] ), .S0(
        n5545), .Y(\i_MIPS/Register/n487 ) );
  CLKMX2X2 U12779 ( .A(n5058), .B(\i_MIPS/Register/register[20][18] ), .S0(
        n5546), .Y(\i_MIPS/Register/n486 ) );
  CLKMX2X2 U12780 ( .A(n5055), .B(\i_MIPS/Register/register[20][17] ), .S0(
        n5546), .Y(\i_MIPS/Register/n485 ) );
  CLKMX2X2 U12781 ( .A(n5028), .B(\i_MIPS/Register/register[20][16] ), .S0(
        n5545), .Y(\i_MIPS/Register/n484 ) );
  CLKMX2X2 U12782 ( .A(n5019), .B(\i_MIPS/Register/register[20][15] ), .S0(
        n5545), .Y(\i_MIPS/Register/n483 ) );
  CLKMX2X2 U12783 ( .A(n5025), .B(\i_MIPS/Register/register[20][14] ), .S0(
        n5545), .Y(\i_MIPS/Register/n482 ) );
  CLKMX2X2 U12784 ( .A(n5052), .B(\i_MIPS/Register/register[20][10] ), .S0(
        n5546), .Y(\i_MIPS/Register/n478 ) );
  CLKMX2X2 U12785 ( .A(n5078), .B(\i_MIPS/Register/register[20][9] ), .S0(
        n5546), .Y(\i_MIPS/Register/n477 ) );
  CLKMX2X2 U12786 ( .A(n5069), .B(\i_MIPS/Register/register[20][7] ), .S0(
        n5546), .Y(\i_MIPS/Register/n475 ) );
  CLKMX2X2 U12787 ( .A(net111837), .B(\i_MIPS/Register/register[20][6] ), .S0(
        n5545), .Y(\i_MIPS/Register/n474 ) );
  CLKMX2X2 U12788 ( .A(n10764), .B(\i_MIPS/Register/register[20][5] ), .S0(
        n5545), .Y(\i_MIPS/Register/n473 ) );
  CLKMX2X2 U12789 ( .A(n5004), .B(\i_MIPS/Register/register[20][3] ), .S0(
        n5545), .Y(\i_MIPS/Register/n471 ) );
  CLKMX2X2 U12790 ( .A(n11217), .B(\i_MIPS/Register/register[21][31] ), .S0(
        n5543), .Y(\i_MIPS/Register/n467 ) );
  CLKMX2X2 U12791 ( .A(n5066), .B(\i_MIPS/Register/register[21][30] ), .S0(
        n5544), .Y(\i_MIPS/Register/n466 ) );
  CLKMX2X2 U12792 ( .A(n5034), .B(\i_MIPS/Register/register[21][29] ), .S0(
        n5544), .Y(\i_MIPS/Register/n465 ) );
  CLKMX2X2 U12793 ( .A(n5013), .B(\i_MIPS/Register/register[21][28] ), .S0(
        n5543), .Y(\i_MIPS/Register/n464 ) );
  CLKMX2X2 U12794 ( .A(n5031), .B(\i_MIPS/Register/register[21][27] ), .S0(
        n5544), .Y(\i_MIPS/Register/n463 ) );
  CLKMX2X2 U12795 ( .A(n5015), .B(\i_MIPS/Register/register[21][26] ), .S0(
        n5543), .Y(\i_MIPS/Register/n462 ) );
  CLKMX2X2 U12796 ( .A(n5022), .B(\i_MIPS/Register/register[21][25] ), .S0(
        n5543), .Y(\i_MIPS/Register/n461 ) );
  CLKMX2X2 U12797 ( .A(n5049), .B(\i_MIPS/Register/register[21][24] ), .S0(
        n5544), .Y(\i_MIPS/Register/n460 ) );
  CLKMX2X2 U12798 ( .A(n5046), .B(\i_MIPS/Register/register[21][23] ), .S0(
        n5544), .Y(\i_MIPS/Register/n459 ) );
  CLKMX2X2 U12799 ( .A(n5043), .B(\i_MIPS/Register/register[21][22] ), .S0(
        n5544), .Y(\i_MIPS/Register/n458 ) );
  CLKMX2X2 U12800 ( .A(n5039), .B(\i_MIPS/Register/register[21][21] ), .S0(
        n5544), .Y(\i_MIPS/Register/n457 ) );
  CLKMX2X2 U12801 ( .A(n5009), .B(\i_MIPS/Register/register[21][19] ), .S0(
        n5543), .Y(\i_MIPS/Register/n455 ) );
  CLKMX2X2 U12802 ( .A(n5057), .B(\i_MIPS/Register/register[21][18] ), .S0(
        n5544), .Y(\i_MIPS/Register/n454 ) );
  CLKMX2X2 U12803 ( .A(n5055), .B(\i_MIPS/Register/register[21][17] ), .S0(
        n5544), .Y(\i_MIPS/Register/n453 ) );
  CLKMX2X2 U12804 ( .A(n5028), .B(\i_MIPS/Register/register[21][16] ), .S0(
        n5543), .Y(\i_MIPS/Register/n452 ) );
  CLKMX2X2 U12805 ( .A(n5019), .B(\i_MIPS/Register/register[21][15] ), .S0(
        n5543), .Y(\i_MIPS/Register/n451 ) );
  CLKMX2X2 U12806 ( .A(n5025), .B(\i_MIPS/Register/register[21][14] ), .S0(
        n5543), .Y(\i_MIPS/Register/n450 ) );
  CLKMX2X2 U12807 ( .A(n5052), .B(\i_MIPS/Register/register[21][10] ), .S0(
        n5544), .Y(\i_MIPS/Register/n446 ) );
  CLKMX2X2 U12808 ( .A(n5078), .B(\i_MIPS/Register/register[21][9] ), .S0(
        n5544), .Y(\i_MIPS/Register/n445 ) );
  CLKMX2X2 U12809 ( .A(n5069), .B(\i_MIPS/Register/register[21][7] ), .S0(
        n5544), .Y(\i_MIPS/Register/n443 ) );
  CLKMX2X2 U12810 ( .A(net111837), .B(\i_MIPS/Register/register[21][6] ), .S0(
        n5543), .Y(\i_MIPS/Register/n442 ) );
  CLKMX2X2 U12811 ( .A(n10764), .B(\i_MIPS/Register/register[21][5] ), .S0(
        n5543), .Y(\i_MIPS/Register/n441 ) );
  CLKMX2X2 U12812 ( .A(n5004), .B(\i_MIPS/Register/register[21][3] ), .S0(
        n5543), .Y(\i_MIPS/Register/n439 ) );
  CLKMX2X2 U12813 ( .A(n5071), .B(\i_MIPS/Register/register[21][2] ), .S0(
        n5544), .Y(\i_MIPS/Register/n438 ) );
  CLKMX2X2 U12814 ( .A(n11217), .B(\i_MIPS/Register/register[22][31] ), .S0(
        n5541), .Y(\i_MIPS/Register/n435 ) );
  CLKMX2X2 U12815 ( .A(n5066), .B(\i_MIPS/Register/register[22][30] ), .S0(
        n5542), .Y(\i_MIPS/Register/n434 ) );
  CLKMX2X2 U12816 ( .A(n5034), .B(\i_MIPS/Register/register[22][29] ), .S0(
        n5542), .Y(\i_MIPS/Register/n433 ) );
  CLKMX2X2 U12817 ( .A(n5013), .B(\i_MIPS/Register/register[22][28] ), .S0(
        n5541), .Y(\i_MIPS/Register/n432 ) );
  CLKMX2X2 U12818 ( .A(n5031), .B(\i_MIPS/Register/register[22][27] ), .S0(
        n5542), .Y(\i_MIPS/Register/n431 ) );
  CLKMX2X2 U12819 ( .A(n5016), .B(\i_MIPS/Register/register[22][26] ), .S0(
        n5541), .Y(\i_MIPS/Register/n430 ) );
  CLKMX2X2 U12820 ( .A(n5022), .B(\i_MIPS/Register/register[22][25] ), .S0(
        n5541), .Y(\i_MIPS/Register/n429 ) );
  CLKMX2X2 U12821 ( .A(n5049), .B(\i_MIPS/Register/register[22][24] ), .S0(
        n5542), .Y(\i_MIPS/Register/n428 ) );
  CLKMX2X2 U12822 ( .A(n5046), .B(\i_MIPS/Register/register[22][23] ), .S0(
        n5542), .Y(\i_MIPS/Register/n427 ) );
  CLKMX2X2 U12823 ( .A(n5043), .B(\i_MIPS/Register/register[22][22] ), .S0(
        n5542), .Y(\i_MIPS/Register/n426 ) );
  CLKMX2X2 U12824 ( .A(n5040), .B(\i_MIPS/Register/register[22][21] ), .S0(
        n5542), .Y(\i_MIPS/Register/n425 ) );
  CLKMX2X2 U12825 ( .A(n5010), .B(\i_MIPS/Register/register[22][19] ), .S0(
        n5541), .Y(\i_MIPS/Register/n423 ) );
  CLKMX2X2 U12826 ( .A(n5058), .B(\i_MIPS/Register/register[22][18] ), .S0(
        n5542), .Y(\i_MIPS/Register/n422 ) );
  CLKMX2X2 U12827 ( .A(n5055), .B(\i_MIPS/Register/register[22][17] ), .S0(
        n5542), .Y(\i_MIPS/Register/n421 ) );
  CLKMX2X2 U12828 ( .A(n5028), .B(\i_MIPS/Register/register[22][16] ), .S0(
        n5541), .Y(\i_MIPS/Register/n420 ) );
  CLKMX2X2 U12829 ( .A(n5019), .B(\i_MIPS/Register/register[22][15] ), .S0(
        n5541), .Y(\i_MIPS/Register/n419 ) );
  CLKMX2X2 U12830 ( .A(n5025), .B(\i_MIPS/Register/register[22][14] ), .S0(
        n5541), .Y(\i_MIPS/Register/n418 ) );
  CLKMX2X2 U12831 ( .A(n5052), .B(\i_MIPS/Register/register[22][10] ), .S0(
        n5542), .Y(\i_MIPS/Register/n414 ) );
  CLKMX2X2 U12832 ( .A(n5078), .B(\i_MIPS/Register/register[22][9] ), .S0(
        n5542), .Y(\i_MIPS/Register/n413 ) );
  CLKMX2X2 U12833 ( .A(n5069), .B(\i_MIPS/Register/register[22][7] ), .S0(
        n5542), .Y(\i_MIPS/Register/n411 ) );
  CLKMX2X2 U12834 ( .A(net111837), .B(\i_MIPS/Register/register[22][6] ), .S0(
        n5541), .Y(\i_MIPS/Register/n410 ) );
  CLKMX2X2 U12835 ( .A(n10764), .B(\i_MIPS/Register/register[22][5] ), .S0(
        n5541), .Y(\i_MIPS/Register/n409 ) );
  CLKMX2X2 U12836 ( .A(n5004), .B(\i_MIPS/Register/register[22][3] ), .S0(
        n5541), .Y(\i_MIPS/Register/n407 ) );
  CLKMX2X2 U12837 ( .A(n5500), .B(\i_MIPS/Register/register[23][31] ), .S0(
        n5539), .Y(\i_MIPS/Register/n403 ) );
  CLKMX2X2 U12838 ( .A(n5066), .B(\i_MIPS/Register/register[23][30] ), .S0(
        n5540), .Y(\i_MIPS/Register/n402 ) );
  CLKMX2X2 U12839 ( .A(n5033), .B(\i_MIPS/Register/register[23][29] ), .S0(
        n5540), .Y(\i_MIPS/Register/n401 ) );
  CLKMX2X2 U12840 ( .A(n5012), .B(\i_MIPS/Register/register[23][28] ), .S0(
        n5539), .Y(\i_MIPS/Register/n400 ) );
  CLKMX2X2 U12841 ( .A(n5030), .B(\i_MIPS/Register/register[23][27] ), .S0(
        n5540), .Y(\i_MIPS/Register/n399 ) );
  CLKMX2X2 U12842 ( .A(n5016), .B(\i_MIPS/Register/register[23][26] ), .S0(
        n5539), .Y(\i_MIPS/Register/n398 ) );
  CLKMX2X2 U12843 ( .A(n5021), .B(\i_MIPS/Register/register[23][25] ), .S0(
        n5539), .Y(\i_MIPS/Register/n397 ) );
  CLKMX2X2 U12844 ( .A(n5048), .B(\i_MIPS/Register/register[23][24] ), .S0(
        n5540), .Y(\i_MIPS/Register/n396 ) );
  CLKMX2X2 U12845 ( .A(n5045), .B(\i_MIPS/Register/register[23][23] ), .S0(
        n5540), .Y(\i_MIPS/Register/n395 ) );
  CLKMX2X2 U12846 ( .A(n5042), .B(\i_MIPS/Register/register[23][22] ), .S0(
        n5540), .Y(\i_MIPS/Register/n394 ) );
  CLKMX2X2 U12847 ( .A(n5040), .B(\i_MIPS/Register/register[23][21] ), .S0(
        n5540), .Y(\i_MIPS/Register/n393 ) );
  CLKMX2X2 U12848 ( .A(n5010), .B(\i_MIPS/Register/register[23][19] ), .S0(
        n5539), .Y(\i_MIPS/Register/n391 ) );
  CLKMX2X2 U12849 ( .A(n5058), .B(\i_MIPS/Register/register[23][18] ), .S0(
        n5540), .Y(\i_MIPS/Register/n390 ) );
  CLKMX2X2 U12850 ( .A(n5054), .B(\i_MIPS/Register/register[23][17] ), .S0(
        n5540), .Y(\i_MIPS/Register/n389 ) );
  CLKMX2X2 U12851 ( .A(n5027), .B(\i_MIPS/Register/register[23][16] ), .S0(
        n5539), .Y(\i_MIPS/Register/n388 ) );
  CLKMX2X2 U12852 ( .A(n5018), .B(\i_MIPS/Register/register[23][15] ), .S0(
        n5539), .Y(\i_MIPS/Register/n387 ) );
  CLKMX2X2 U12853 ( .A(n5024), .B(\i_MIPS/Register/register[23][14] ), .S0(
        n5539), .Y(\i_MIPS/Register/n386 ) );
  CLKMX2X2 U12854 ( .A(n5051), .B(\i_MIPS/Register/register[23][10] ), .S0(
        n5540), .Y(\i_MIPS/Register/n382 ) );
  CLKMX2X2 U12855 ( .A(n5077), .B(\i_MIPS/Register/register[23][9] ), .S0(
        n5540), .Y(\i_MIPS/Register/n381 ) );
  CLKMX2X2 U12856 ( .A(n5068), .B(\i_MIPS/Register/register[23][7] ), .S0(
        n5540), .Y(\i_MIPS/Register/n379 ) );
  CLKMX2X2 U12857 ( .A(net111835), .B(\i_MIPS/Register/register[23][6] ), .S0(
        n5539), .Y(\i_MIPS/Register/n378 ) );
  CLKMX2X2 U12858 ( .A(n5075), .B(\i_MIPS/Register/register[23][5] ), .S0(
        n5539), .Y(\i_MIPS/Register/n377 ) );
  CLKMX2X2 U12859 ( .A(n5003), .B(\i_MIPS/Register/register[23][3] ), .S0(
        n5539), .Y(\i_MIPS/Register/n375 ) );
  CLKMX2X2 U12860 ( .A(n5072), .B(\i_MIPS/Register/register[23][2] ), .S0(
        n5540), .Y(\i_MIPS/Register/n374 ) );
  CLKMX2X2 U12861 ( .A(n11217), .B(\i_MIPS/Register/register[24][31] ), .S0(
        n5537), .Y(\i_MIPS/Register/n371 ) );
  CLKMX2X2 U12862 ( .A(n5066), .B(\i_MIPS/Register/register[24][30] ), .S0(
        n5538), .Y(\i_MIPS/Register/n370 ) );
  CLKMX2X2 U12863 ( .A(n5034), .B(\i_MIPS/Register/register[24][29] ), .S0(
        n5538), .Y(\i_MIPS/Register/n369 ) );
  CLKMX2X2 U12864 ( .A(n5013), .B(\i_MIPS/Register/register[24][28] ), .S0(
        n5537), .Y(\i_MIPS/Register/n368 ) );
  CLKMX2X2 U12865 ( .A(n5031), .B(\i_MIPS/Register/register[24][27] ), .S0(
        n5538), .Y(\i_MIPS/Register/n367 ) );
  CLKMX2X2 U12866 ( .A(n5016), .B(\i_MIPS/Register/register[24][26] ), .S0(
        n5537), .Y(\i_MIPS/Register/n366 ) );
  CLKMX2X2 U12867 ( .A(n5022), .B(\i_MIPS/Register/register[24][25] ), .S0(
        n5537), .Y(\i_MIPS/Register/n365 ) );
  CLKMX2X2 U12868 ( .A(n5049), .B(\i_MIPS/Register/register[24][24] ), .S0(
        n5538), .Y(\i_MIPS/Register/n364 ) );
  CLKMX2X2 U12869 ( .A(n5046), .B(\i_MIPS/Register/register[24][23] ), .S0(
        n5538), .Y(\i_MIPS/Register/n363 ) );
  CLKMX2X2 U12870 ( .A(n5043), .B(\i_MIPS/Register/register[24][22] ), .S0(
        n5538), .Y(\i_MIPS/Register/n362 ) );
  CLKMX2X2 U12871 ( .A(n5040), .B(\i_MIPS/Register/register[24][21] ), .S0(
        n5538), .Y(\i_MIPS/Register/n361 ) );
  CLKMX2X2 U12872 ( .A(n5010), .B(\i_MIPS/Register/register[24][19] ), .S0(
        n5537), .Y(\i_MIPS/Register/n359 ) );
  CLKMX2X2 U12873 ( .A(n5058), .B(\i_MIPS/Register/register[24][18] ), .S0(
        n5538), .Y(\i_MIPS/Register/n358 ) );
  CLKMX2X2 U12874 ( .A(n5055), .B(\i_MIPS/Register/register[24][17] ), .S0(
        n5538), .Y(\i_MIPS/Register/n357 ) );
  CLKMX2X2 U12875 ( .A(n5028), .B(\i_MIPS/Register/register[24][16] ), .S0(
        n5537), .Y(\i_MIPS/Register/n356 ) );
  CLKMX2X2 U12876 ( .A(n5019), .B(\i_MIPS/Register/register[24][15] ), .S0(
        n5537), .Y(\i_MIPS/Register/n355 ) );
  CLKMX2X2 U12877 ( .A(n5025), .B(\i_MIPS/Register/register[24][14] ), .S0(
        n5537), .Y(\i_MIPS/Register/n354 ) );
  CLKMX2X2 U12878 ( .A(n5052), .B(\i_MIPS/Register/register[24][10] ), .S0(
        n5538), .Y(\i_MIPS/Register/n350 ) );
  CLKMX2X2 U12879 ( .A(n5078), .B(\i_MIPS/Register/register[24][9] ), .S0(
        n5538), .Y(\i_MIPS/Register/n349 ) );
  CLKMX2X2 U12880 ( .A(n5069), .B(\i_MIPS/Register/register[24][7] ), .S0(
        n5538), .Y(\i_MIPS/Register/n347 ) );
  CLKMX2X2 U12881 ( .A(net111837), .B(\i_MIPS/Register/register[24][6] ), .S0(
        n5537), .Y(\i_MIPS/Register/n346 ) );
  CLKMX2X2 U12882 ( .A(n10764), .B(\i_MIPS/Register/register[24][5] ), .S0(
        n5537), .Y(\i_MIPS/Register/n345 ) );
  CLKMX2X2 U12883 ( .A(n5004), .B(\i_MIPS/Register/register[24][3] ), .S0(
        n5537), .Y(\i_MIPS/Register/n343 ) );
  CLKMX2X2 U12884 ( .A(n11217), .B(\i_MIPS/Register/register[25][31] ), .S0(
        n5535), .Y(\i_MIPS/Register/n339 ) );
  CLKMX2X2 U12885 ( .A(n5066), .B(\i_MIPS/Register/register[25][30] ), .S0(
        n5536), .Y(\i_MIPS/Register/n338 ) );
  CLKMX2X2 U12886 ( .A(n5034), .B(\i_MIPS/Register/register[25][29] ), .S0(
        n5536), .Y(\i_MIPS/Register/n337 ) );
  CLKMX2X2 U12887 ( .A(n5013), .B(\i_MIPS/Register/register[25][28] ), .S0(
        n5535), .Y(\i_MIPS/Register/n336 ) );
  CLKMX2X2 U12888 ( .A(n5031), .B(\i_MIPS/Register/register[25][27] ), .S0(
        n5536), .Y(\i_MIPS/Register/n335 ) );
  CLKMX2X2 U12889 ( .A(n5016), .B(\i_MIPS/Register/register[25][26] ), .S0(
        n5535), .Y(\i_MIPS/Register/n334 ) );
  CLKMX2X2 U12890 ( .A(n5022), .B(\i_MIPS/Register/register[25][25] ), .S0(
        n5535), .Y(\i_MIPS/Register/n333 ) );
  CLKMX2X2 U12891 ( .A(n5049), .B(\i_MIPS/Register/register[25][24] ), .S0(
        n5536), .Y(\i_MIPS/Register/n332 ) );
  CLKMX2X2 U12892 ( .A(n5046), .B(\i_MIPS/Register/register[25][23] ), .S0(
        n5536), .Y(\i_MIPS/Register/n331 ) );
  CLKMX2X2 U12893 ( .A(n5043), .B(\i_MIPS/Register/register[25][22] ), .S0(
        n5536), .Y(\i_MIPS/Register/n330 ) );
  CLKMX2X2 U12894 ( .A(n5040), .B(\i_MIPS/Register/register[25][21] ), .S0(
        n5536), .Y(\i_MIPS/Register/n329 ) );
  CLKMX2X2 U12895 ( .A(n5010), .B(\i_MIPS/Register/register[25][19] ), .S0(
        n5535), .Y(\i_MIPS/Register/n327 ) );
  CLKMX2X2 U12896 ( .A(n5058), .B(\i_MIPS/Register/register[25][18] ), .S0(
        n5536), .Y(\i_MIPS/Register/n326 ) );
  CLKMX2X2 U12897 ( .A(n5055), .B(\i_MIPS/Register/register[25][17] ), .S0(
        n5536), .Y(\i_MIPS/Register/n325 ) );
  CLKMX2X2 U12898 ( .A(n5028), .B(\i_MIPS/Register/register[25][16] ), .S0(
        n5535), .Y(\i_MIPS/Register/n324 ) );
  CLKMX2X2 U12899 ( .A(n5019), .B(\i_MIPS/Register/register[25][15] ), .S0(
        n5535), .Y(\i_MIPS/Register/n323 ) );
  CLKMX2X2 U12900 ( .A(n5025), .B(\i_MIPS/Register/register[25][14] ), .S0(
        n5535), .Y(\i_MIPS/Register/n322 ) );
  CLKMX2X2 U12901 ( .A(n5052), .B(\i_MIPS/Register/register[25][10] ), .S0(
        n5536), .Y(\i_MIPS/Register/n318 ) );
  CLKMX2X2 U12902 ( .A(n5078), .B(\i_MIPS/Register/register[25][9] ), .S0(
        n5536), .Y(\i_MIPS/Register/n317 ) );
  CLKMX2X2 U12903 ( .A(n5069), .B(\i_MIPS/Register/register[25][7] ), .S0(
        n5536), .Y(\i_MIPS/Register/n315 ) );
  CLKMX2X2 U12904 ( .A(net111837), .B(\i_MIPS/Register/register[25][6] ), .S0(
        n5535), .Y(\i_MIPS/Register/n314 ) );
  CLKMX2X2 U12905 ( .A(n10764), .B(\i_MIPS/Register/register[25][5] ), .S0(
        n5535), .Y(\i_MIPS/Register/n313 ) );
  CLKMX2X2 U12906 ( .A(n5004), .B(\i_MIPS/Register/register[25][3] ), .S0(
        n5535), .Y(\i_MIPS/Register/n311 ) );
  CLKMX2X2 U12907 ( .A(n11217), .B(\i_MIPS/Register/register[26][31] ), .S0(
        n5533), .Y(\i_MIPS/Register/n307 ) );
  CLKMX2X2 U12908 ( .A(n5066), .B(\i_MIPS/Register/register[26][30] ), .S0(
        n5534), .Y(\i_MIPS/Register/n306 ) );
  CLKMX2X2 U12909 ( .A(n5034), .B(\i_MIPS/Register/register[26][29] ), .S0(
        n5534), .Y(\i_MIPS/Register/n305 ) );
  CLKMX2X2 U12910 ( .A(n5013), .B(\i_MIPS/Register/register[26][28] ), .S0(
        n5533), .Y(\i_MIPS/Register/n304 ) );
  CLKMX2X2 U12911 ( .A(n5031), .B(\i_MIPS/Register/register[26][27] ), .S0(
        n5534), .Y(\i_MIPS/Register/n303 ) );
  CLKMX2X2 U12912 ( .A(n5016), .B(\i_MIPS/Register/register[26][26] ), .S0(
        n5533), .Y(\i_MIPS/Register/n302 ) );
  CLKMX2X2 U12913 ( .A(n5022), .B(\i_MIPS/Register/register[26][25] ), .S0(
        n5533), .Y(\i_MIPS/Register/n301 ) );
  CLKMX2X2 U12914 ( .A(n5049), .B(\i_MIPS/Register/register[26][24] ), .S0(
        n5534), .Y(\i_MIPS/Register/n300 ) );
  CLKMX2X2 U12915 ( .A(n5046), .B(\i_MIPS/Register/register[26][23] ), .S0(
        n5534), .Y(\i_MIPS/Register/n299 ) );
  CLKMX2X2 U12916 ( .A(n5043), .B(\i_MIPS/Register/register[26][22] ), .S0(
        n5534), .Y(\i_MIPS/Register/n298 ) );
  CLKMX2X2 U12917 ( .A(n5040), .B(\i_MIPS/Register/register[26][21] ), .S0(
        n5534), .Y(\i_MIPS/Register/n297 ) );
  CLKMX2X2 U12918 ( .A(n5010), .B(\i_MIPS/Register/register[26][19] ), .S0(
        n5533), .Y(\i_MIPS/Register/n295 ) );
  CLKMX2X2 U12919 ( .A(n5058), .B(\i_MIPS/Register/register[26][18] ), .S0(
        n5534), .Y(\i_MIPS/Register/n294 ) );
  CLKMX2X2 U12920 ( .A(n5055), .B(\i_MIPS/Register/register[26][17] ), .S0(
        n5534), .Y(\i_MIPS/Register/n293 ) );
  CLKMX2X2 U12921 ( .A(n5028), .B(\i_MIPS/Register/register[26][16] ), .S0(
        n5533), .Y(\i_MIPS/Register/n292 ) );
  CLKMX2X2 U12922 ( .A(n5019), .B(\i_MIPS/Register/register[26][15] ), .S0(
        n5533), .Y(\i_MIPS/Register/n291 ) );
  CLKMX2X2 U12923 ( .A(n5025), .B(\i_MIPS/Register/register[26][14] ), .S0(
        n5533), .Y(\i_MIPS/Register/n290 ) );
  CLKMX2X2 U12924 ( .A(n5052), .B(\i_MIPS/Register/register[26][10] ), .S0(
        n5534), .Y(\i_MIPS/Register/n286 ) );
  CLKMX2X2 U12925 ( .A(n5078), .B(\i_MIPS/Register/register[26][9] ), .S0(
        n5534), .Y(\i_MIPS/Register/n285 ) );
  CLKMX2X2 U12926 ( .A(n5069), .B(\i_MIPS/Register/register[26][7] ), .S0(
        n5534), .Y(\i_MIPS/Register/n283 ) );
  CLKMX2X2 U12927 ( .A(net111837), .B(\i_MIPS/Register/register[26][6] ), .S0(
        n5533), .Y(\i_MIPS/Register/n282 ) );
  CLKMX2X2 U12928 ( .A(n10764), .B(\i_MIPS/Register/register[26][5] ), .S0(
        n5533), .Y(\i_MIPS/Register/n281 ) );
  CLKMX2X2 U12929 ( .A(n5004), .B(\i_MIPS/Register/register[26][3] ), .S0(
        n5533), .Y(\i_MIPS/Register/n279 ) );
  CLKMX2X2 U12930 ( .A(n5500), .B(\i_MIPS/Register/register[27][31] ), .S0(
        n5531), .Y(\i_MIPS/Register/n275 ) );
  CLKMX2X2 U12931 ( .A(n5066), .B(\i_MIPS/Register/register[27][30] ), .S0(
        n5532), .Y(\i_MIPS/Register/n274 ) );
  CLKMX2X2 U12932 ( .A(n5034), .B(\i_MIPS/Register/register[27][29] ), .S0(
        n5532), .Y(\i_MIPS/Register/n273 ) );
  CLKMX2X2 U12933 ( .A(n5013), .B(\i_MIPS/Register/register[27][28] ), .S0(
        n5531), .Y(\i_MIPS/Register/n272 ) );
  CLKMX2X2 U12934 ( .A(n5031), .B(\i_MIPS/Register/register[27][27] ), .S0(
        n5532), .Y(\i_MIPS/Register/n271 ) );
  CLKMX2X2 U12935 ( .A(n5015), .B(\i_MIPS/Register/register[27][26] ), .S0(
        n5531), .Y(\i_MIPS/Register/n270 ) );
  CLKMX2X2 U12936 ( .A(n5022), .B(\i_MIPS/Register/register[27][25] ), .S0(
        n5531), .Y(\i_MIPS/Register/n269 ) );
  CLKMX2X2 U12937 ( .A(n5049), .B(\i_MIPS/Register/register[27][24] ), .S0(
        n5532), .Y(\i_MIPS/Register/n268 ) );
  CLKMX2X2 U12938 ( .A(n5046), .B(\i_MIPS/Register/register[27][23] ), .S0(
        n5532), .Y(\i_MIPS/Register/n267 ) );
  CLKMX2X2 U12939 ( .A(n5043), .B(\i_MIPS/Register/register[27][22] ), .S0(
        n5532), .Y(\i_MIPS/Register/n266 ) );
  CLKMX2X2 U12940 ( .A(n5039), .B(\i_MIPS/Register/register[27][21] ), .S0(
        n5532), .Y(\i_MIPS/Register/n265 ) );
  CLKMX2X2 U12941 ( .A(n5009), .B(\i_MIPS/Register/register[27][19] ), .S0(
        n5531), .Y(\i_MIPS/Register/n263 ) );
  CLKMX2X2 U12942 ( .A(n5057), .B(\i_MIPS/Register/register[27][18] ), .S0(
        n5532), .Y(\i_MIPS/Register/n262 ) );
  CLKMX2X2 U12943 ( .A(n5055), .B(\i_MIPS/Register/register[27][17] ), .S0(
        n5532), .Y(\i_MIPS/Register/n261 ) );
  CLKMX2X2 U12944 ( .A(n5028), .B(\i_MIPS/Register/register[27][16] ), .S0(
        n5531), .Y(\i_MIPS/Register/n260 ) );
  CLKMX2X2 U12945 ( .A(n5019), .B(\i_MIPS/Register/register[27][15] ), .S0(
        n5531), .Y(\i_MIPS/Register/n259 ) );
  CLKMX2X2 U12946 ( .A(n5025), .B(\i_MIPS/Register/register[27][14] ), .S0(
        n5531), .Y(\i_MIPS/Register/n258 ) );
  CLKMX2X2 U12947 ( .A(n5052), .B(\i_MIPS/Register/register[27][10] ), .S0(
        n5532), .Y(\i_MIPS/Register/n254 ) );
  CLKMX2X2 U12948 ( .A(n5078), .B(\i_MIPS/Register/register[27][9] ), .S0(
        n5532), .Y(\i_MIPS/Register/n253 ) );
  CLKMX2X2 U12949 ( .A(n5069), .B(\i_MIPS/Register/register[27][7] ), .S0(
        n5532), .Y(\i_MIPS/Register/n251 ) );
  CLKMX2X2 U12950 ( .A(net111837), .B(\i_MIPS/Register/register[27][6] ), .S0(
        n5531), .Y(\i_MIPS/Register/n250 ) );
  CLKMX2X2 U12951 ( .A(n5075), .B(\i_MIPS/Register/register[27][5] ), .S0(
        n5531), .Y(\i_MIPS/Register/n249 ) );
  CLKMX2X2 U12952 ( .A(n5004), .B(\i_MIPS/Register/register[27][3] ), .S0(
        n5531), .Y(\i_MIPS/Register/n247 ) );
  CLKMX2X2 U12953 ( .A(n5071), .B(\i_MIPS/Register/register[27][2] ), .S0(
        n5532), .Y(\i_MIPS/Register/n246 ) );
  CLKMX2X2 U12954 ( .A(n11217), .B(\i_MIPS/Register/register[28][31] ), .S0(
        n5529), .Y(\i_MIPS/Register/n243 ) );
  CLKMX2X2 U12955 ( .A(n5066), .B(\i_MIPS/Register/register[28][30] ), .S0(
        n5530), .Y(\i_MIPS/Register/n242 ) );
  CLKMX2X2 U12956 ( .A(n5034), .B(\i_MIPS/Register/register[28][29] ), .S0(
        n5530), .Y(\i_MIPS/Register/n241 ) );
  CLKMX2X2 U12957 ( .A(n5013), .B(\i_MIPS/Register/register[28][28] ), .S0(
        n5529), .Y(\i_MIPS/Register/n240 ) );
  CLKMX2X2 U12958 ( .A(n5031), .B(\i_MIPS/Register/register[28][27] ), .S0(
        n5530), .Y(\i_MIPS/Register/n239 ) );
  CLKMX2X2 U12959 ( .A(n5016), .B(\i_MIPS/Register/register[28][26] ), .S0(
        n5529), .Y(\i_MIPS/Register/n238 ) );
  CLKMX2X2 U12960 ( .A(n5022), .B(\i_MIPS/Register/register[28][25] ), .S0(
        n5529), .Y(\i_MIPS/Register/n237 ) );
  CLKMX2X2 U12961 ( .A(n5049), .B(\i_MIPS/Register/register[28][24] ), .S0(
        n5530), .Y(\i_MIPS/Register/n236 ) );
  CLKMX2X2 U12962 ( .A(n5046), .B(\i_MIPS/Register/register[28][23] ), .S0(
        n5530), .Y(\i_MIPS/Register/n235 ) );
  CLKMX2X2 U12963 ( .A(n5043), .B(\i_MIPS/Register/register[28][22] ), .S0(
        n5530), .Y(\i_MIPS/Register/n234 ) );
  CLKMX2X2 U12964 ( .A(n5040), .B(\i_MIPS/Register/register[28][21] ), .S0(
        n5530), .Y(\i_MIPS/Register/n233 ) );
  CLKMX2X2 U12965 ( .A(n5010), .B(\i_MIPS/Register/register[28][19] ), .S0(
        n5529), .Y(\i_MIPS/Register/n231 ) );
  CLKMX2X2 U12966 ( .A(n5058), .B(\i_MIPS/Register/register[28][18] ), .S0(
        n5530), .Y(\i_MIPS/Register/n230 ) );
  CLKMX2X2 U12967 ( .A(n5055), .B(\i_MIPS/Register/register[28][17] ), .S0(
        n5530), .Y(\i_MIPS/Register/n229 ) );
  CLKMX2X2 U12968 ( .A(n5028), .B(\i_MIPS/Register/register[28][16] ), .S0(
        n5529), .Y(\i_MIPS/Register/n228 ) );
  CLKMX2X2 U12969 ( .A(n5019), .B(\i_MIPS/Register/register[28][15] ), .S0(
        n5529), .Y(\i_MIPS/Register/n227 ) );
  CLKMX2X2 U12970 ( .A(n5025), .B(\i_MIPS/Register/register[28][14] ), .S0(
        n5529), .Y(\i_MIPS/Register/n226 ) );
  CLKMX2X2 U12971 ( .A(n5052), .B(\i_MIPS/Register/register[28][10] ), .S0(
        n5530), .Y(\i_MIPS/Register/n222 ) );
  CLKMX2X2 U12972 ( .A(n5078), .B(\i_MIPS/Register/register[28][9] ), .S0(
        n5530), .Y(\i_MIPS/Register/n221 ) );
  CLKMX2X2 U12973 ( .A(n5069), .B(\i_MIPS/Register/register[28][7] ), .S0(
        n5530), .Y(\i_MIPS/Register/n219 ) );
  CLKMX2X2 U12974 ( .A(net111837), .B(\i_MIPS/Register/register[28][6] ), .S0(
        n5529), .Y(\i_MIPS/Register/n218 ) );
  CLKMX2X2 U12975 ( .A(n10764), .B(\i_MIPS/Register/register[28][5] ), .S0(
        n5529), .Y(\i_MIPS/Register/n217 ) );
  CLKMX2X2 U12976 ( .A(n5004), .B(\i_MIPS/Register/register[28][3] ), .S0(
        n5529), .Y(\i_MIPS/Register/n215 ) );
  CLKMX2X2 U12977 ( .A(n9126), .B(\i_MIPS/Register/register[29][31] ), .S0(
        n5527), .Y(\i_MIPS/Register/n211 ) );
  CLKMX2X2 U12978 ( .A(n5066), .B(\i_MIPS/Register/register[29][30] ), .S0(
        n5528), .Y(\i_MIPS/Register/n210 ) );
  CLKMX2X2 U12979 ( .A(n5033), .B(\i_MIPS/Register/register[29][29] ), .S0(
        n5528), .Y(\i_MIPS/Register/n209 ) );
  CLKMX2X2 U12980 ( .A(n5012), .B(\i_MIPS/Register/register[29][28] ), .S0(
        n5527), .Y(\i_MIPS/Register/n208 ) );
  CLKMX2X2 U12981 ( .A(n5030), .B(\i_MIPS/Register/register[29][27] ), .S0(
        n5528), .Y(\i_MIPS/Register/n207 ) );
  CLKMX2X2 U12982 ( .A(n5016), .B(\i_MIPS/Register/register[29][26] ), .S0(
        n5527), .Y(\i_MIPS/Register/n206 ) );
  CLKMX2X2 U12983 ( .A(n5021), .B(\i_MIPS/Register/register[29][25] ), .S0(
        n5527), .Y(\i_MIPS/Register/n205 ) );
  CLKMX2X2 U12984 ( .A(n5048), .B(\i_MIPS/Register/register[29][24] ), .S0(
        n5528), .Y(\i_MIPS/Register/n204 ) );
  CLKMX2X2 U12985 ( .A(n5045), .B(\i_MIPS/Register/register[29][23] ), .S0(
        n5528), .Y(\i_MIPS/Register/n203 ) );
  CLKMX2X2 U12986 ( .A(n5042), .B(\i_MIPS/Register/register[29][22] ), .S0(
        n5528), .Y(\i_MIPS/Register/n202 ) );
  CLKMX2X2 U12987 ( .A(n5040), .B(\i_MIPS/Register/register[29][21] ), .S0(
        n5528), .Y(\i_MIPS/Register/n201 ) );
  CLKMX2X2 U12988 ( .A(n5010), .B(\i_MIPS/Register/register[29][19] ), .S0(
        n5527), .Y(\i_MIPS/Register/n199 ) );
  CLKMX2X2 U12989 ( .A(n5058), .B(\i_MIPS/Register/register[29][18] ), .S0(
        n5528), .Y(\i_MIPS/Register/n198 ) );
  CLKMX2X2 U12990 ( .A(n5054), .B(\i_MIPS/Register/register[29][17] ), .S0(
        n5528), .Y(\i_MIPS/Register/n197 ) );
  CLKMX2X2 U12991 ( .A(n5027), .B(\i_MIPS/Register/register[29][16] ), .S0(
        n5527), .Y(\i_MIPS/Register/n196 ) );
  CLKMX2X2 U12992 ( .A(n5018), .B(\i_MIPS/Register/register[29][15] ), .S0(
        n5527), .Y(\i_MIPS/Register/n195 ) );
  CLKMX2X2 U12993 ( .A(n5024), .B(\i_MIPS/Register/register[29][14] ), .S0(
        n5527), .Y(\i_MIPS/Register/n194 ) );
  CLKMX2X2 U12994 ( .A(n5051), .B(\i_MIPS/Register/register[29][10] ), .S0(
        n5528), .Y(\i_MIPS/Register/n190 ) );
  CLKMX2X2 U12995 ( .A(n5077), .B(\i_MIPS/Register/register[29][9] ), .S0(
        n5528), .Y(\i_MIPS/Register/n189 ) );
  CLKMX2X2 U12996 ( .A(n5068), .B(\i_MIPS/Register/register[29][7] ), .S0(
        n5528), .Y(\i_MIPS/Register/n187 ) );
  CLKMX2X2 U12997 ( .A(net111835), .B(\i_MIPS/Register/register[29][6] ), .S0(
        n5527), .Y(\i_MIPS/Register/n186 ) );
  CLKMX2X2 U12998 ( .A(n5075), .B(\i_MIPS/Register/register[29][5] ), .S0(
        n5527), .Y(\i_MIPS/Register/n185 ) );
  CLKMX2X2 U12999 ( .A(n5003), .B(\i_MIPS/Register/register[29][3] ), .S0(
        n5527), .Y(\i_MIPS/Register/n183 ) );
  CLKMX2X2 U13000 ( .A(n5072), .B(\i_MIPS/Register/register[29][2] ), .S0(
        n5528), .Y(\i_MIPS/Register/n182 ) );
  CLKMX2X2 U13001 ( .A(n5500), .B(\i_MIPS/Register/register[30][31] ), .S0(
        n5525), .Y(\i_MIPS/Register/n179 ) );
  CLKMX2X2 U13002 ( .A(n5066), .B(\i_MIPS/Register/register[30][30] ), .S0(
        n5526), .Y(\i_MIPS/Register/n178 ) );
  CLKMX2X2 U13003 ( .A(n5034), .B(\i_MIPS/Register/register[30][29] ), .S0(
        n5526), .Y(\i_MIPS/Register/n177 ) );
  CLKMX2X2 U13004 ( .A(n5013), .B(\i_MIPS/Register/register[30][28] ), .S0(
        n5525), .Y(\i_MIPS/Register/n176 ) );
  CLKMX2X2 U13005 ( .A(n5031), .B(\i_MIPS/Register/register[30][27] ), .S0(
        n5526), .Y(\i_MIPS/Register/n175 ) );
  CLKMX2X2 U13006 ( .A(n5016), .B(\i_MIPS/Register/register[30][26] ), .S0(
        n5525), .Y(\i_MIPS/Register/n174 ) );
  CLKMX2X2 U13007 ( .A(n5022), .B(\i_MIPS/Register/register[30][25] ), .S0(
        n5525), .Y(\i_MIPS/Register/n173 ) );
  CLKMX2X2 U13008 ( .A(n5049), .B(\i_MIPS/Register/register[30][24] ), .S0(
        n5526), .Y(\i_MIPS/Register/n172 ) );
  CLKMX2X2 U13009 ( .A(n5046), .B(\i_MIPS/Register/register[30][23] ), .S0(
        n5526), .Y(\i_MIPS/Register/n171 ) );
  CLKMX2X2 U13010 ( .A(n5043), .B(\i_MIPS/Register/register[30][22] ), .S0(
        n5526), .Y(\i_MIPS/Register/n170 ) );
  CLKMX2X2 U13011 ( .A(n5040), .B(\i_MIPS/Register/register[30][21] ), .S0(
        n5526), .Y(\i_MIPS/Register/n169 ) );
  CLKMX2X2 U13012 ( .A(n5010), .B(\i_MIPS/Register/register[30][19] ), .S0(
        n5525), .Y(\i_MIPS/Register/n167 ) );
  CLKMX2X2 U13013 ( .A(n5058), .B(\i_MIPS/Register/register[30][18] ), .S0(
        n5526), .Y(\i_MIPS/Register/n166 ) );
  CLKMX2X2 U13014 ( .A(n5055), .B(\i_MIPS/Register/register[30][17] ), .S0(
        n5526), .Y(\i_MIPS/Register/n165 ) );
  CLKMX2X2 U13015 ( .A(n5028), .B(\i_MIPS/Register/register[30][16] ), .S0(
        n5525), .Y(\i_MIPS/Register/n164 ) );
  CLKMX2X2 U13016 ( .A(n5019), .B(\i_MIPS/Register/register[30][15] ), .S0(
        n5525), .Y(\i_MIPS/Register/n163 ) );
  CLKMX2X2 U13017 ( .A(n5025), .B(\i_MIPS/Register/register[30][14] ), .S0(
        n5525), .Y(\i_MIPS/Register/n162 ) );
  CLKMX2X2 U13018 ( .A(n5052), .B(\i_MIPS/Register/register[30][10] ), .S0(
        n5526), .Y(\i_MIPS/Register/n158 ) );
  CLKMX2X2 U13019 ( .A(n5078), .B(\i_MIPS/Register/register[30][9] ), .S0(
        n5526), .Y(\i_MIPS/Register/n157 ) );
  CLKMX2X2 U13020 ( .A(n5069), .B(\i_MIPS/Register/register[30][7] ), .S0(
        n5526), .Y(\i_MIPS/Register/n155 ) );
  CLKMX2X2 U13021 ( .A(net111837), .B(\i_MIPS/Register/register[30][6] ), .S0(
        n5525), .Y(\i_MIPS/Register/n154 ) );
  CLKMX2X2 U13022 ( .A(n10764), .B(\i_MIPS/Register/register[30][5] ), .S0(
        n5525), .Y(\i_MIPS/Register/n153 ) );
  CLKMX2X2 U13023 ( .A(n5004), .B(\i_MIPS/Register/register[30][3] ), .S0(
        n5525), .Y(\i_MIPS/Register/n151 ) );
  CLKINVX1 U13024 ( .A(\i_MIPS/n255 ), .Y(n10461) );
  MX2XL U13025 ( .A(n3708), .B(\i_MIPS/Sign_Extend_ID[3] ), .S0(n5507), .Y(
        \i_MIPS/n509 ) );
  MX2XL U13026 ( .A(n5589), .B(\i_MIPS/Sign_Extend_ID[8] ), .S0(n5507), .Y(
        \i_MIPS/n504 ) );
  MXI2X1 U13027 ( .A(n4710), .B(n4711), .S0(n5507), .Y(\i_MIPS/n469 ) );
  AND2XL U13028 ( .A(net98970), .B(net98971), .Y(n4711) );
  CLKMX2X2 U13029 ( .A(\i_MIPS/ID_EX[41] ), .B(n10850), .S0(n5507), .Y(
        \i_MIPS/n437 ) );
  NAND3BXL U13030 ( .AN(net98897), .B(net98898), .C(net98899), .Y(n10850) );
  INVXL U13031 ( .A(net98900), .Y(net98897) );
  MX2XL U13032 ( .A(\i_MIPS/ID_EX[73] ), .B(\i_MIPS/Sign_Extend_ID[0] ), .S0(
        n5508), .Y(\i_MIPS/n512 ) );
  MX2XL U13033 ( .A(n3768), .B(\i_MIPS/Sign_Extend_ID[1] ), .S0(n5508), .Y(
        \i_MIPS/n511 ) );
  MX2XL U13034 ( .A(n3700), .B(\i_MIPS/Sign_Extend_ID[4] ), .S0(n5508), .Y(
        \i_MIPS/n508 ) );
  MX2XL U13035 ( .A(\i_MIPS/ID_EX[78] ), .B(\i_MIPS/Sign_Extend_ID[5] ), .S0(
        n5508), .Y(\i_MIPS/n507 ) );
  MX2XL U13036 ( .A(n12951), .B(n4066), .S0(n5509), .Y(\i_MIPS/n450 ) );
  MX2XL U13037 ( .A(n12945), .B(net99605), .S0(n5509), .Y(\i_MIPS/n444 ) );
  CLKINVX1 U13038 ( .A(\i_MIPS/Control_ID/n10 ), .Y(n10002) );
  AO22X1 U13039 ( .A0(\i_MIPS/control_out[7] ), .A1(net110227), .B0(
        \i_MIPS/ALUOp[1] ), .B1(n5516), .Y(\i_MIPS/n471 ) );
  AO22XL U13040 ( .A0(net110227), .A1(n11167), .B0(n5517), .B1(n4413), .Y(
        \i_MIPS/n472 ) );
  OAI31XL U13041 ( .A0(n11166), .A1(\i_MIPS/IR_ID[30] ), .A2(
        \i_MIPS/IR_ID[27] ), .B0(\i_MIPS/Control_ID/n15 ), .Y(n11167) );
  NAND3BX1 U13042 ( .AN(n11165), .B(\i_MIPS/IR_ID[28] ), .C(\i_MIPS/n328 ), 
        .Y(n11166) );
  AO22XL U13043 ( .A0(n173), .A1(n11019), .B0(net113592), .B1(n10051), .Y(
        \i_MIPS/N73 ) );
  CLKINVX1 U13044 ( .A(\i_MIPS/n316 ), .Y(n10051) );
  AO22XL U13045 ( .A0(n174), .A1(n11218), .B0(net113592), .B1(
        \i_MIPS/IR_ID[17] ), .Y(\i_MIPS/N72 ) );
  CLKINVX1 U13046 ( .A(\i_MIPS/n312 ), .Y(n10080) );
  AO22X1 U13047 ( .A0(\i_MIPS/control_out[0] ), .A1(net110227), .B0(n5512), 
        .B1(\i_MIPS/ID_EX_0 ), .Y(\i_MIPS/n528 ) );
  NAND3BX1 U13048 ( .AN(\i_MIPS/control_out[7] ), .B(n5522), .C(
        \i_MIPS/Control_ID/n12 ), .Y(\i_MIPS/control_out[0] ) );
  AO21XL U13049 ( .A0(\i_MIPS/ID_EX[99] ), .A1(n5516), .B0(n4499), .Y(
        \i_MIPS/n486 ) );
  OAI2BB1XL U13050 ( .A0N(n5514), .A1N(n3507), .B0(n11200), .Y(\i_MIPS/n480 )
         );
  AO21XL U13051 ( .A0(n5513), .A1(n3504), .B0(n4588), .Y(\i_MIPS/n527 ) );
  XOR2XL U13052 ( .A(n6291), .B(\i_MIPS/IR_ID[19] ), .Y(n6204) );
  XOR2XL U13053 ( .A(n10129), .B(net108963), .Y(n6203) );
  AND3X2 U13054 ( .A(\i_MIPS/Register/n120 ), .B(n4715), .C(\i_MIPS/Reg_W[3] ), 
        .Y(\i_MIPS/Register/n131 ) );
  AND3X2 U13055 ( .A(\i_MIPS/Register/n120 ), .B(n4716), .C(\i_MIPS/Reg_W[4] ), 
        .Y(\i_MIPS/Register/n122 ) );
  AND3X2 U13056 ( .A(\i_MIPS/Register/n120 ), .B(\i_MIPS/Reg_W[3] ), .C(
        \i_MIPS/Reg_W[4] ), .Y(\i_MIPS/Register/n104 ) );
  XOR2XL U13057 ( .A(\i_MIPS/n313 ), .B(\i_MIPS/IR_ID[16] ), .Y(n5941) );
  XOR2XL U13058 ( .A(\i_MIPS/n317 ), .B(\i_MIPS/IR_ID[18] ), .Y(n5942) );
  XOR2XL U13059 ( .A(\i_MIPS/n228 ), .B(\i_MIPS/ID_EX[111] ), .Y(n5943) );
  XOR2XL U13060 ( .A(\i_MIPS/n230 ), .B(\i_MIPS/ID_EX[113] ), .Y(n5944) );
  NAND3BX1 U13061 ( .AN(\i_MIPS/IR_ID[28] ), .B(\i_MIPS/n328 ), .C(
        \i_MIPS/n330 ), .Y(n9808) );
  NOR2X1 U13062 ( .A(\i_MIPS/Sign_Extend_ID[0] ), .B(
        \i_MIPS/Sign_Extend_ID[5] ), .Y(net101971) );
  NOR2X1 U13063 ( .A(\i_MIPS/Sign_Extend_ID[2] ), .B(
        \i_MIPS/Sign_Extend_ID[4] ), .Y(net101973) );
  NOR2BX1 U13064 ( .AN(\i_MIPS/Sign_Extend_ID[3] ), .B(\i_MIPS/Control_ID/n10 ), .Y(net101970) );
  AND2X2 U13065 ( .A(\i_MIPS/IR_ID[27] ), .B(\i_MIPS/IR_ID[26] ), .Y(n4717) );
  CLKINVX1 U13066 ( .A(mem_ready_D), .Y(n11548) );
  CLKBUFX3 U13067 ( .A(\i_MIPS/IR_ID[25] ), .Y(n5588) );
  CLKBUFX3 U13068 ( .A(mem_ready_I), .Y(n4793) );
  NAND3BX1 U13069 ( .AN(n9691), .B(\i_MIPS/IR_ID[29] ), .C(n9690), .Y(
        \i_MIPS/Control_ID/n15 ) );
  AOI2BB1X1 U13070 ( .A0N(\i_MIPS/n322 ), .A1N(\i_MIPS/n332 ), .B0(
        \i_MIPS/IR_ID[30] ), .Y(n9690) );
  XOR2X1 U13071 ( .A(n9689), .B(n9688), .Y(n9691) );
  NAND2X1 U13072 ( .A(\i_MIPS/IR_ID[28] ), .B(\i_MIPS/n324 ), .Y(n9689) );
  NAND2X1 U13073 ( .A(\i_MIPS/IR_ID[31] ), .B(n4637), .Y(
        \i_MIPS/Control_ID/n12 ) );
  MX2XL U13074 ( .A(n12941), .B(n3651), .S0(n5508), .Y(\i_MIPS/n440 ) );
  NAND2X1 U13075 ( .A(n8144), .B(n8143), .Y(n8158) );
  MX2XL U13076 ( .A(n12946), .B(n3995), .S0(n5510), .Y(\i_MIPS/n445 ) );
  INVXL U13077 ( .A(n6598), .Y(n6346) );
  NAND2XL U13078 ( .A(n6602), .B(n6598), .Y(n6251) );
  MX2XL U13079 ( .A(n3743), .B(n152), .S0(n5510), .Y(\i_MIPS/n417 ) );
  NAND2XL U13080 ( .A(n7622), .B(n8714), .Y(n7623) );
  MX2XL U13081 ( .A(n12942), .B(n3528), .S0(n5508), .Y(\i_MIPS/n441 ) );
  NAND2X1 U13082 ( .A(n8524), .B(n8071), .Y(n7802) );
  MX2XL U13083 ( .A(n3501), .B(n4030), .S0(n5507), .Y(\i_MIPS/n377 ) );
  NAND2XL U13084 ( .A(n3796), .B(n3744), .Y(n7278) );
  MX2XL U13085 ( .A(n12944), .B(n10407), .S0(n5509), .Y(\i_MIPS/n443 ) );
  MX2XL U13086 ( .A(n3503), .B(net99624), .S0(n5506), .Y(\i_MIPS/n385 ) );
  MX2XL U13087 ( .A(DCACHE_addr[1]), .B(net99078), .S0(n5511), .Y(
        \i_MIPS/n466 ) );
  NAND3BX4 U13088 ( .AN(n4549), .B(n9613), .C(n9614), .Y(n11053) );
  XOR2X4 U13089 ( .A(n11382), .B(ICACHE_addr[23]), .Y(n9550) );
  XOR2X4 U13090 ( .A(n11383), .B(ICACHE_addr[24]), .Y(n9552) );
  NAND2XL U13091 ( .A(n7856), .B(n7777), .Y(n7714) );
  MX2XL U13092 ( .A(DCACHE_addr[21]), .B(net99384), .S0(n5507), .Y(
        \i_MIPS/n446 ) );
  OAI221XL U13093 ( .A0(net103390), .A1(net112707), .B0(net103391), .B1(
        net112721), .C0(net103392), .Y(n4747) );
  MX2XL U13094 ( .A(DCACHE_addr[16]), .B(n166), .S0(n5509), .Y(\i_MIPS/n451 )
         );
  INVX12 U13095 ( .A(n4748), .Y(DCACHE_addr[10]) );
  INVX12 U13096 ( .A(n4752), .Y(DCACHE_addr[15]) );
  INVX12 U13097 ( .A(n4754), .Y(DCACHE_addr[23]) );
  INVX12 U13098 ( .A(n4756), .Y(DCACHE_addr[19]) );
  INVX8 U13099 ( .A(n11228), .Y(n11229) );
  XOR2X4 U13100 ( .A(n11370), .B(ICACHE_addr[11]), .Y(n9335) );
  NAND2X1 U13101 ( .A(n10658), .B(n3774), .Y(n11534) );
  NAND2X1 U13102 ( .A(n10653), .B(n1637), .Y(n11537) );
  NAND2X1 U13103 ( .A(n10645), .B(n10644), .Y(n11538) );
  NAND2XL U13104 ( .A(n9620), .B(n3692), .Y(n9621) );
  XOR2X1 U13105 ( .A(n3819), .B(ICACHE_addr[0]), .Y(n11183) );
  XOR2X4 U13106 ( .A(n11381), .B(ICACHE_addr[22]), .Y(n9581) );
  NAND4X8 U13107 ( .A(n5948), .B(n5947), .C(n5946), .D(n5945), .Y(n11389) );
  XOR2X4 U13108 ( .A(n11375), .B(ICACHE_addr[16]), .Y(n9571) );
  AO21X4 U13109 ( .A0(n10830), .A1(n10829), .B0(net113077), .Y(n7671) );
  MX2XL U13110 ( .A(n3495), .B(net99378), .S0(n5510), .Y(\i_MIPS/n391 ) );
  XOR2X4 U13111 ( .A(n11380), .B(ICACHE_addr[21]), .Y(n9573) );
  AND2XL U13112 ( .A(n10151), .B(n11168), .Y(n4783) );
  CLKMX2X2 U13113 ( .A(n3488), .B(n4747), .S0(n5507), .Y(\i_MIPS/n387 ) );
  NAND2X1 U13114 ( .A(n12951), .B(net113089), .Y(n10185) );
  NAND2BX4 U13115 ( .AN(n9178), .B(n9177), .Y(n9263) );
  XOR2X4 U13116 ( .A(n11371), .B(ICACHE_addr[12]), .Y(n9569) );
  OAI221X4 U13117 ( .A0(n3609), .A1(n10504), .B0(n10503), .B1(n10502), .C0(
        n10501), .Y(n10717) );
  XOR2X4 U13118 ( .A(n11376), .B(ICACHE_addr[17]), .Y(n9574) );
  NAND2X8 U13119 ( .A(n9133), .B(\i_MIPS/ID_EX[83] ), .Y(n8726) );
  OA22X4 U13120 ( .A0(net112425), .A1(n2353), .B0(net112301), .B1(n851), .Y(
        n5947) );
  OA22X4 U13121 ( .A0(net112231), .A1(n2354), .B0(net112159), .B1(n852), .Y(
        n5946) );
  OA22X4 U13122 ( .A0(net112071), .A1(n2355), .B0(net111889), .B1(n853), .Y(
        n5945) );
  OA22X4 U13123 ( .A0(n5421), .A1(n1605), .B0(n5375), .B1(n3269), .Y(n5949) );
  OA22X4 U13124 ( .A0(n5421), .A1(n427), .B0(n5377), .B1(n3270), .Y(n5954) );
  OA22X4 U13125 ( .A0(n5334), .A1(n3285), .B0(n5317), .B1(n1625), .Y(n5962) );
  OA22X4 U13126 ( .A0(n5422), .A1(n3308), .B0(n5379), .B1(n408), .Y(n5965) );
  OA22X4 U13127 ( .A0(n5423), .A1(n3235), .B0(n5379), .B1(n1597), .Y(n5967) );
  OA22X4 U13128 ( .A0(n5426), .A1(n428), .B0(n5382), .B1(n3271), .Y(n5977) );
  OA22X4 U13129 ( .A0(n5427), .A1(n1606), .B0(n5385), .B1(n3272), .Y(n5979) );
  OA22X4 U13130 ( .A0(n5248), .A1(n3236), .B0(n5203), .B1(n1598), .Y(n5983) );
  OA22X4 U13131 ( .A0(n3611), .A1(n1607), .B0(n5383), .B1(n3273), .Y(n5981) );
  OA22X4 U13132 ( .A0(n5163), .A1(n1979), .B0(n5120), .B1(n412), .Y(n6010) );
  OA22X4 U13133 ( .A0(n5333), .A1(n3286), .B0(n5290), .B1(n1626), .Y(n6008) );
  OA22X4 U13134 ( .A0(n5428), .A1(n1980), .B0(n5384), .B1(n413), .Y(n6007) );
  OA22X4 U13135 ( .A0(n5163), .A1(n1981), .B0(n5120), .B1(n414), .Y(n6018) );
  OA22X4 U13136 ( .A0(n5249), .A1(n1982), .B0(n5204), .B1(n415), .Y(n6017) );
  OA22X4 U13137 ( .A0(n5428), .A1(n1983), .B0(n5384), .B1(n416), .Y(n6015) );
  OA22X4 U13138 ( .A0(n5163), .A1(n1984), .B0(n5120), .B1(n417), .Y(n6023) );
  OA22X4 U13139 ( .A0(n5249), .A1(n1985), .B0(n5204), .B1(n418), .Y(n6022) );
  OA22X4 U13140 ( .A0(n5428), .A1(n1986), .B0(n5384), .B1(n419), .Y(n6020) );
  OAI221X2 U13141 ( .A0(n6173), .A1(\i_MIPS/n335 ), .B0(n5498), .B1(n11389), 
        .C0(n6172), .Y(net98375) );
  OAI31X2 U13142 ( .A0(n6200), .A1(n10133), .A2(n10131), .B0(\i_MIPS/ID_EX_0 ), 
        .Y(n6201) );
  NAND4BBX4 U13143 ( .AN(n6206), .BN(n6205), .C(\i_MIPS/EX_MEM_0 ), .D(
        net112721), .Y(net101983) );
  AO22X4 U13144 ( .A0(n5595), .A1(n10837), .B0(n5593), .B1(n3768), .Y(n6234)
         );
  CLKINVX3 U13145 ( .A(\i_MIPS/ID_EX[83] ), .Y(n7698) );
  NAND4BBX4 U13146 ( .AN(n6304), .BN(n6303), .C(\i_MIPS/EX_MEM_0 ), .D(n6302), 
        .Y(net102088) );
  AO22X4 U13147 ( .A0(net102300), .A1(n6325), .B0(net113039), .B1(net99016), 
        .Y(net107168) );
  AOI2BB1X2 U13148 ( .A0N(n6651), .A1N(n9156), .B0(n8339), .Y(n6418) );
  NAND2X2 U13149 ( .A(\i_MIPS/ALUin1[16] ), .B(n6573), .Y(n8151) );
  NAND2X2 U13150 ( .A(\i_MIPS/ALUin1[25] ), .B(n6591), .Y(n8435) );
  NAND2X2 U13151 ( .A(\i_MIPS/ALUin1[24] ), .B(n6592), .Y(n8901) );
  OAI211X2 U13152 ( .A0(n4007), .A1(n6769), .B0(n6606), .C0(n6607), .Y(n6608)
         );
  OAI211X2 U13153 ( .A0(n6611), .A1(n3624), .B0(n6608), .C0(n6609), .Y(n8644)
         );
  AO22X4 U13154 ( .A0(n6623), .A1(n4434), .B0(n6622), .B1(n3826), .Y(n8152) );
  AOI211X2 U13155 ( .A0(n6631), .A1(n6630), .B0(n6629), .C0(n6628), .Y(n6647)
         );
  AO21X4 U13156 ( .A0(net99060), .A1(net99061), .B0(net112727), .Y(net106272)
         );
  AO21X4 U13157 ( .A0(n6929), .A1(n6928), .B0(n6932), .Y(n6938) );
  AO21X4 U13158 ( .A0(net99977), .A1(net99978), .B0(net112727), .Y(net105931)
         );
  AO21X4 U13159 ( .A0(net99108), .A1(net99109), .B0(net112727), .Y(net105152)
         );
  AO21X4 U13160 ( .A0(n10830), .A1(n10829), .B0(net112729), .Y(net104869) );
  NAND4BX2 U13161 ( .AN(n9149), .B(n9148), .C(n9147), .D(n9146), .Y(n9188) );
  AOI2BB1X2 U13162 ( .A0N(n4563), .A1N(n9152), .B0(n9151), .Y(n9159) );
  NAND3BX2 U13163 ( .AN(net113919), .B(net113083), .C(n4601), .Y(n9253) );
  AO21X4 U13164 ( .A0(n10696), .A1(n10695), .B0(net112731), .Y(n9325) );
  AO21X4 U13165 ( .A0(n4778), .A1(n10147), .B0(n10145), .Y(n11201) );
  AO21X4 U13166 ( .A0(n4778), .A1(n10146), .B0(n10145), .Y(n11205) );
  CLKINVX3 U13167 ( .A(n10158), .Y(n10160) );
  NAND4X2 U13168 ( .A(n11039), .B(\i_MIPS/Pred_2bit/current_state[1] ), .C(
        n11040), .D(n4511), .Y(n10389) );
  NAND2BX4 U13169 ( .AN(n10252), .B(n10255), .Y(net98429) );
  CLKINVX3 U13170 ( .A(n10720), .Y(n10724) );
  NAND3BX2 U13171 ( .AN(n10933), .B(n10932), .C(n10931), .Y(\i_MIPS/PC/n50 )
         );
  AOI2BB2X2 U13172 ( .B0(\i_MIPS/IF_ID[70] ), .B1(n149), .A0N(net110191), 
        .A1N(\i_MIPS/n185 ), .Y(n11054) );
endmodule

