
module CHIP ( clk, rst_n, mem_read_D, mem_write_D, mem_addr_D, mem_wdata_D, 
        mem_rdata_D, mem_ready_D, mem_read_I, mem_write_I, mem_addr_I, 
        mem_wdata_I, mem_rdata_I, mem_ready_I, DCACHE_addr, DCACHE_wdata, 
        DCACHE_wen );
  output [31:4] mem_addr_D;
  output [127:0] mem_wdata_D;
  input [127:0] mem_rdata_D;
  output [31:4] mem_addr_I;
  output [127:0] mem_wdata_I;
  input [127:0] mem_rdata_I;
  output [29:0] DCACHE_addr;
  output [31:0] DCACHE_wdata;
  input clk, rst_n, mem_ready_D, mem_ready_I;
  output mem_read_D, mem_write_D, mem_read_I, mem_write_I, DCACHE_wen;
  wire   n12846, n12847, n12848, n12849, n12850, n12851, n12852, n12853,
         n12854, n12855, n12856, n12857, n12858, n12859, n12860, n12861,
         n12862, n12863, n12864, n12865, n12866, n12867, n12868, n12869,
         n12870, n12871, n12872, n12873, n12874, n12875, n12876, n12877,
         n12878, n12879, n12880, n12881, n12882, n12883, n12884, n12885,
         n12886, n12887, n12888, n12889, n12890, n12891, n12892, n12893,
         n12894, n12895, n12896, n12897, n12898, n12899, n12900, n12901,
         n12902, n12903, n12904, n12905, n12906, n12907, n12908, n12909,
         n12910, n12911, n12912, n12913, n12914, n12915, n12916, n12917,
         n12918, n12919, n12920, n12921, n12922, n12923, n12924, n12925,
         n12926, n12927, n12928, n12929, n12930, n12931, n12932, n12933,
         n12934, n12935, n12936, n12937, n12938, n12939, n12940, n12941,
         n12942, n12943, n12944, n12945, n12946, n12947, n12948, n12949,
         n12950, n12951, n12952, n12953, n12954, n12955, n12956, n12957,
         n12958, n12959, n12960, n12961, n12962, n12963, n12964, n12965,
         n12966, n12967, n12968, n12969, n12970, n12971, n12972, n12973,
         n12974, n12975, n12976, n12977, n12978, n12979, n12980, n12981,
         n12982, n12983, n12984, n12985, n12986, n12987, n12988, n12989,
         n12990, n12991, n12992, n12993, n12994, n12995, n12996, n12997,
         n12998, n12999, n13000, n13001, n13002, n13003, n13004, n13005,
         n13006, n13007, n13008, n13009, n13010, n13011, n13012, n13013,
         DCACHE_ren, \i_MIPS/n525 , \i_MIPS/n524 , \i_MIPS/n523 ,
         \i_MIPS/n522 , \i_MIPS/n521 , \i_MIPS/n520 , \i_MIPS/n519 ,
         \i_MIPS/n518 , \i_MIPS/n517 , \i_MIPS/n516 , \i_MIPS/n515 ,
         \i_MIPS/n514 , \i_MIPS/n513 , \i_MIPS/n512 , \i_MIPS/n511 ,
         \i_MIPS/n510 , \i_MIPS/n509 , \i_MIPS/n508 , \i_MIPS/n507 ,
         \i_MIPS/n506 , \i_MIPS/n505 , \i_MIPS/n504 , \i_MIPS/n503 ,
         \i_MIPS/n502 , \i_MIPS/n501 , \i_MIPS/n500 , \i_MIPS/n499 ,
         \i_MIPS/n498 , \i_MIPS/n497 , \i_MIPS/n496 , \i_MIPS/n493 ,
         \i_MIPS/n492 , \i_MIPS/n491 , \i_MIPS/n490 , \i_MIPS/n489 ,
         \i_MIPS/n488 , \i_MIPS/n487 , \i_MIPS/n486 , \i_MIPS/n485 ,
         \i_MIPS/n484 , \i_MIPS/n483 , \i_MIPS/n482 , \i_MIPS/n481 ,
         \i_MIPS/n480 , \i_MIPS/n479 , \i_MIPS/n478 , \i_MIPS/n477 ,
         \i_MIPS/n476 , \i_MIPS/n475 , \i_MIPS/n474 , \i_MIPS/n473 ,
         \i_MIPS/n472 , \i_MIPS/n471 , \i_MIPS/n470 , \i_MIPS/n469 ,
         \i_MIPS/n468 , \i_MIPS/n467 , \i_MIPS/n466 , \i_MIPS/n465 ,
         \i_MIPS/n464 , \i_MIPS/n463 , \i_MIPS/n462 , \i_MIPS/n461 ,
         \i_MIPS/n460 , \i_MIPS/n459 , \i_MIPS/n458 , \i_MIPS/n457 ,
         \i_MIPS/n456 , \i_MIPS/n455 , \i_MIPS/n454 , \i_MIPS/n453 ,
         \i_MIPS/n452 , \i_MIPS/n451 , \i_MIPS/n450 , \i_MIPS/n449 ,
         \i_MIPS/n448 , \i_MIPS/n447 , \i_MIPS/n446 , \i_MIPS/n445 ,
         \i_MIPS/n444 , \i_MIPS/n443 , \i_MIPS/n442 , \i_MIPS/n441 ,
         \i_MIPS/n440 , \i_MIPS/n439 , \i_MIPS/n438 , \i_MIPS/n437 ,
         \i_MIPS/n436 , \i_MIPS/n435 , \i_MIPS/n434 , \i_MIPS/n433 ,
         \i_MIPS/n432 , \i_MIPS/n431 , \i_MIPS/n430 , \i_MIPS/n429 ,
         \i_MIPS/n428 , \i_MIPS/n427 , \i_MIPS/n426 , \i_MIPS/n425 ,
         \i_MIPS/n424 , \i_MIPS/n423 , \i_MIPS/n422 , \i_MIPS/n421 ,
         \i_MIPS/n420 , \i_MIPS/n419 , \i_MIPS/n418 , \i_MIPS/n417 ,
         \i_MIPS/n416 , \i_MIPS/n415 , \i_MIPS/n414 , \i_MIPS/n413 ,
         \i_MIPS/n412 , \i_MIPS/n411 , \i_MIPS/n410 , \i_MIPS/n409 ,
         \i_MIPS/n408 , \i_MIPS/n407 , \i_MIPS/n406 , \i_MIPS/n405 ,
         \i_MIPS/n404 , \i_MIPS/n403 , \i_MIPS/n402 , \i_MIPS/n401 ,
         \i_MIPS/n400 , \i_MIPS/n399 , \i_MIPS/n398 , \i_MIPS/n397 ,
         \i_MIPS/n396 , \i_MIPS/n395 , \i_MIPS/n394 , \i_MIPS/n393 ,
         \i_MIPS/n392 , \i_MIPS/n391 , \i_MIPS/n390 , \i_MIPS/n389 ,
         \i_MIPS/n388 , \i_MIPS/n387 , \i_MIPS/n386 , \i_MIPS/n385 ,
         \i_MIPS/n384 , \i_MIPS/n383 , \i_MIPS/n382 , \i_MIPS/n381 ,
         \i_MIPS/n380 , \i_MIPS/n379 , \i_MIPS/n378 , \i_MIPS/n377 ,
         \i_MIPS/n376 , \i_MIPS/n375 , \i_MIPS/n374 , \i_MIPS/n373 ,
         \i_MIPS/n372 , \i_MIPS/n371 , \i_MIPS/n370 , \i_MIPS/n369 ,
         \i_MIPS/n368 , \i_MIPS/n367 , \i_MIPS/n366 , \i_MIPS/n365 ,
         \i_MIPS/n364 , \i_MIPS/n363 , \i_MIPS/n362 , \i_MIPS/n361 ,
         \i_MIPS/n360 , \i_MIPS/n359 , \i_MIPS/n358 , \i_MIPS/n357 ,
         \i_MIPS/n356 , \i_MIPS/n355 , \i_MIPS/n354 , \i_MIPS/n353 ,
         \i_MIPS/n352 , \i_MIPS/n351 , \i_MIPS/n350 , \i_MIPS/n349 ,
         \i_MIPS/n348 , \i_MIPS/n347 , \i_MIPS/n346 , \i_MIPS/n345 ,
         \i_MIPS/n344 , \i_MIPS/n343 , \i_MIPS/n342 , \i_MIPS/n341 ,
         \i_MIPS/n340 , \i_MIPS/n339 , \i_MIPS/n338 , \i_MIPS/n337 ,
         \i_MIPS/n336 , \i_MIPS/n335 , \i_MIPS/n334 , \i_MIPS/n333 ,
         \i_MIPS/n332 , \i_MIPS/n331 , \i_MIPS/n330 , \i_MIPS/n329 ,
         \i_MIPS/n328 , \i_MIPS/n327 , \i_MIPS/n326 , \i_MIPS/n325 ,
         \i_MIPS/n324 , \i_MIPS/n323 , \i_MIPS/n322 , \i_MIPS/n321 ,
         \i_MIPS/n320 , \i_MIPS/n319 , \i_MIPS/n318 , \i_MIPS/n317 ,
         \i_MIPS/n316 , \i_MIPS/n315 , \i_MIPS/n314 , \i_MIPS/n313 ,
         \i_MIPS/n312 , \i_MIPS/n311 , \i_MIPS/n310 , \i_MIPS/n309 ,
         \i_MIPS/n308 , \i_MIPS/n307 , \i_MIPS/n306 , \i_MIPS/n305 ,
         \i_MIPS/n304 , \i_MIPS/n303 , \i_MIPS/n302 , \i_MIPS/n301 ,
         \i_MIPS/n300 , \i_MIPS/n299 , \i_MIPS/n297 , \i_MIPS/n296 ,
         \i_MIPS/n287 , \i_MIPS/n271 , \i_MIPS/n270 , \i_MIPS/n269 ,
         \i_MIPS/n268 , \i_MIPS/n267 , \i_MIPS/n266 , \i_MIPS/n265 ,
         \i_MIPS/n264 , \i_MIPS/n263 , \i_MIPS/n262 , \i_MIPS/n261 ,
         \i_MIPS/n260 , \i_MIPS/n259 , \i_MIPS/n258 , \i_MIPS/n257 ,
         \i_MIPS/n256 , \i_MIPS/n255 , \i_MIPS/n254 , \i_MIPS/n253 ,
         \i_MIPS/n252 , \i_MIPS/n251 , \i_MIPS/n250 , \i_MIPS/n249 ,
         \i_MIPS/n248 , \i_MIPS/n247 , \i_MIPS/n246 , \i_MIPS/n245 ,
         \i_MIPS/n243 , \i_MIPS/n242 , \i_MIPS/n241 , \i_MIPS/n240 ,
         \i_MIPS/n239 , \i_MIPS/n237 , \i_MIPS/n236 , \i_MIPS/n235 ,
         \i_MIPS/n234 , \i_MIPS/n233 , \i_MIPS/n232 , \i_MIPS/n231 ,
         \i_MIPS/n230 , \i_MIPS/n229 , \i_MIPS/n228 , \i_MIPS/n227 ,
         \i_MIPS/n226 , \i_MIPS/n225 , \i_MIPS/n223 , \i_MIPS/n222 ,
         \i_MIPS/n221 , \i_MIPS/n220 , \i_MIPS/n219 , \i_MIPS/n218 ,
         \i_MIPS/n217 , \i_MIPS/n216 , \i_MIPS/n215 , \i_MIPS/n214 ,
         \i_MIPS/n213 , \i_MIPS/n212 , \i_MIPS/n211 , \i_MIPS/n210 ,
         \i_MIPS/n209 , \i_MIPS/n208 , \i_MIPS/n207 , \i_MIPS/n206 ,
         \i_MIPS/n205 , \i_MIPS/n204 , \i_MIPS/n203 , \i_MIPS/n202 ,
         \i_MIPS/n201 , \i_MIPS/n200 , \i_MIPS/n199 , \i_MIPS/n198 ,
         \i_MIPS/n197 , \i_MIPS/n196 , \i_MIPS/n195 , \i_MIPS/n194 ,
         \i_MIPS/n193 , \i_MIPS/n192 , \i_MIPS/n191 , \i_MIPS/n190 ,
         \i_MIPS/n189 , \i_MIPS/n188 , \i_MIPS/n187 , \i_MIPS/n186 ,
         \i_MIPS/n185 , \i_MIPS/n184 , \i_MIPS/n183 , \i_MIPS/n182 ,
         \i_MIPS/n181 , \i_MIPS/n180 , \i_MIPS/n179 , \i_MIPS/n178 ,
         \i_MIPS/n177 , \i_MIPS/n176 , \i_MIPS/n175 , \i_MIPS/n174 ,
         \i_MIPS/n173 , \i_MIPS/n172 , \i_MIPS/n171 , \i_MIPS/n170 ,
         \i_MIPS/n169 , \i_MIPS/n168 , \i_MIPS/n167 , \i_MIPS/n166 ,
         \i_MIPS/n165 , \i_MIPS/n164 , \i_MIPS/n163 , \i_MIPS/n162 ,
         \i_MIPS/n161 , \i_MIPS/n160 , \i_MIPS/n159 , \i_MIPS/n158 ,
         \i_MIPS/n157 , \i_MIPS/n156 , \i_MIPS/n155 , \i_MIPS/n154 ,
         \i_MIPS/n153 , \i_MIPS/N80 , \i_MIPS/N79 , \i_MIPS/N78 , \i_MIPS/N77 ,
         \i_MIPS/N76 , \i_MIPS/N75 , \i_MIPS/N74 , \i_MIPS/N73 , \i_MIPS/N72 ,
         \i_MIPS/N71 , \i_MIPS/N70 , \i_MIPS/N69 , \i_MIPS/N68 , \i_MIPS/N67 ,
         \i_MIPS/N66 , \i_MIPS/N65 , \i_MIPS/N64 , \i_MIPS/N63 , \i_MIPS/N62 ,
         \i_MIPS/N61 , \i_MIPS/N60 , \i_MIPS/N59 , \i_MIPS/N58 , \i_MIPS/N57 ,
         \i_MIPS/N56 , \i_MIPS/N55 , \i_MIPS/N54 , \i_MIPS/N53 , \i_MIPS/N52 ,
         \i_MIPS/N51 , \i_MIPS/N50 , \i_MIPS/N49 , \i_MIPS/N48 , \i_MIPS/N47 ,
         \i_MIPS/N46 , \i_MIPS/N45 , \i_MIPS/N44 , \i_MIPS/N43 , \i_MIPS/N42 ,
         \i_MIPS/N41 , \i_MIPS/N40 , \i_MIPS/N39 , \i_MIPS/N38 , \i_MIPS/N37 ,
         \i_MIPS/N36 , \i_MIPS/N35 , \i_MIPS/N34 , \i_MIPS/N33 , \i_MIPS/N32 ,
         \i_MIPS/N31 , \i_MIPS/N30 , \i_MIPS/N29 , \i_MIPS/N28 , \i_MIPS/N27 ,
         \i_MIPS/N26 , \i_MIPS/N25 , \i_MIPS/N24 , \i_MIPS/N23 , \i_MIPS/N22 ,
         \i_MIPS/N21 , \i_MIPS/N20 , \i_MIPS/N19 , \i_MIPS/N18 , \i_MIPS/N17 ,
         \i_MIPS/ALUin1[30] , \i_MIPS/ALUin1[29] , \i_MIPS/ALUin1[28] ,
         \i_MIPS/ALUin1[27] , \i_MIPS/ALUin1[26] , \i_MIPS/ALUin1[25] ,
         \i_MIPS/ALUin1[24] , \i_MIPS/ALUin1[23] , \i_MIPS/ALUin1[22] ,
         \i_MIPS/ALUin1[21] , \i_MIPS/ALUin1[20] , \i_MIPS/ALUin1[19] ,
         \i_MIPS/ALUin1[18] , \i_MIPS/ALUin1[17] , \i_MIPS/ALUin1[16] ,
         \i_MIPS/ALUin1[15] , \i_MIPS/ALUin1[14] , \i_MIPS/ALUin1[13] ,
         \i_MIPS/ALUin1[12] , \i_MIPS/ALUin1[11] , \i_MIPS/ALUin1[10] ,
         \i_MIPS/ALUin1[9] , \i_MIPS/ALUin1[8] , \i_MIPS/ALUin1[7] ,
         \i_MIPS/ALUin1[6] , \i_MIPS/ALUin1[5] , \i_MIPS/ALUin1[4] ,
         \i_MIPS/ALUin1[3] , \i_MIPS/ALUin1[2] , \i_MIPS/ALUin1[1] ,
         \i_MIPS/ALUin1[0] , \i_MIPS/ALUOp[1] , \i_MIPS/EX_MEM_0 ,
         \i_MIPS/EX_MEM_1 , \i_MIPS/EX_MEM[5] , \i_MIPS/EX_MEM[6] ,
         \i_MIPS/EX_MEM_74 , \i_MIPS/ID_EX_0 , \i_MIPS/ID_EX_3 ,
         \i_MIPS/ID_EX_5 , \i_MIPS/ID_EX[43] , \i_MIPS/ID_EX[47] ,
         \i_MIPS/ID_EX[48] , \i_MIPS/ID_EX[50] , \i_MIPS/ID_EX[63] ,
         \i_MIPS/ID_EX[64] , \i_MIPS/ID_EX[65] , \i_MIPS/ID_EX[66] ,
         \i_MIPS/ID_EX[67] , \i_MIPS/ID_EX[68] , \i_MIPS/ID_EX[69] ,
         \i_MIPS/ID_EX[70] , \i_MIPS/ID_EX[71] , \i_MIPS/ID_EX[74] ,
         \i_MIPS/ID_EX[76] , \i_MIPS/ID_EX[78] , \i_MIPS/ID_EX[81] ,
         \i_MIPS/ID_EX[83] , \i_MIPS/ID_EX[84] , \i_MIPS/ID_EX[85] ,
         \i_MIPS/ID_EX[86] , \i_MIPS/ID_EX[87] , \i_MIPS/ID_EX[88] ,
         \i_MIPS/ID_EX[89] , \i_MIPS/ID_EX[90] , \i_MIPS/ID_EX[91] ,
         \i_MIPS/ID_EX[92] , \i_MIPS/ID_EX[93] , \i_MIPS/ID_EX[94] ,
         \i_MIPS/ID_EX[95] , \i_MIPS/ID_EX[96] , \i_MIPS/ID_EX[97] ,
         \i_MIPS/ID_EX[98] , \i_MIPS/ID_EX[99] , \i_MIPS/ID_EX[100] ,
         \i_MIPS/ID_EX[101] , \i_MIPS/ID_EX[102] , \i_MIPS/ID_EX[103] ,
         \i_MIPS/ID_EX[104] , \i_MIPS/ID_EX[105] , \i_MIPS/ID_EX[106] ,
         \i_MIPS/ID_EX[107] , \i_MIPS/ID_EX[111] , \i_MIPS/ID_EX[112] ,
         \i_MIPS/ID_EX[113] , \i_MIPS/ID_EX[114] , \i_MIPS/ID_EX[115] ,
         \i_MIPS/control_out[7] , \i_MIPS/control_out[6] ,
         \i_MIPS/control_out[0] , \i_MIPS/Reg_W[0] , \i_MIPS/Reg_W[1] ,
         \i_MIPS/Reg_W[2] , \i_MIPS/Reg_W[3] , \i_MIPS/Reg_W[4] ,
         \i_MIPS/PC_o[1] , \i_MIPS/PC_add4[0] , \i_MIPS/jump_addr[18] ,
         \i_MIPS/jump_addr[22] , \i_MIPS/jump_addr[23] ,
         \i_MIPS/jump_addr[26] , \i_MIPS/jump_addr[28] ,
         \i_MIPS/jump_addr[29] , \i_MIPS/jump_addr[30] ,
         \i_MIPS/jump_addr[31] , \i_MIPS/IR[31] , \i_MIPS/IR[30] ,
         \i_MIPS/IR[29] , \i_MIPS/IR[28] , \i_MIPS/IR[27] , \i_MIPS/IR[26] ,
         \i_MIPS/Sign_Extend[0] , \i_MIPS/Sign_Extend[1] ,
         \i_MIPS/Sign_Extend[2] , \i_MIPS/Sign_Extend[3] ,
         \i_MIPS/Sign_Extend[5] , \i_MIPS/Sign_Extend[8] ,
         \i_MIPS/Sign_Extend[9] , \i_MIPS/Sign_Extend[10] ,
         \i_MIPS/Sign_Extend[11] , \i_MIPS/Sign_Extend[12] ,
         \i_MIPS/Sign_Extend[13] , \i_MIPS/Sign_Extend[14] ,
         \i_MIPS/Sign_Extend[31] , \i_MIPS/IF_ID[2] , \i_MIPS/IF_ID[3] ,
         \i_MIPS/IF_ID[4] , \i_MIPS/IF_ID[5] , \i_MIPS/IF_ID[6] ,
         \i_MIPS/IF_ID[7] , \i_MIPS/IF_ID[8] , \i_MIPS/IF_ID[9] ,
         \i_MIPS/IF_ID[10] , \i_MIPS/IF_ID[11] , \i_MIPS/IF_ID[12] ,
         \i_MIPS/IF_ID[13] , \i_MIPS/IF_ID[14] , \i_MIPS/IF_ID[15] ,
         \i_MIPS/IF_ID[16] , \i_MIPS/IF_ID[17] , \i_MIPS/IF_ID[18] ,
         \i_MIPS/IF_ID[19] , \i_MIPS/IF_ID[20] , \i_MIPS/IF_ID[21] ,
         \i_MIPS/IF_ID[22] , \i_MIPS/IF_ID[23] , \i_MIPS/IF_ID[24] ,
         \i_MIPS/IF_ID[25] , \i_MIPS/IF_ID[26] , \i_MIPS/IF_ID[27] ,
         \D_cache/n1796 , \D_cache/n1795 , \D_cache/n1794 , \D_cache/n1793 ,
         \D_cache/n1792 , \D_cache/n1791 , \D_cache/n1790 , \D_cache/n1789 ,
         \D_cache/n1788 , \D_cache/n1787 , \D_cache/n1786 , \D_cache/n1785 ,
         \D_cache/n1784 , \D_cache/n1783 , \D_cache/n1782 , \D_cache/n1781 ,
         \D_cache/n1780 , \D_cache/n1779 , \D_cache/n1778 , \D_cache/n1777 ,
         \D_cache/n1776 , \D_cache/n1775 , \D_cache/n1774 , \D_cache/n1773 ,
         \D_cache/n1772 , \D_cache/n1771 , \D_cache/n1770 , \D_cache/n1769 ,
         \D_cache/n1768 , \D_cache/n1767 , \D_cache/n1766 , \D_cache/n1765 ,
         \D_cache/n1764 , \D_cache/n1763 , \D_cache/n1762 , \D_cache/n1761 ,
         \D_cache/n1760 , \D_cache/n1759 , \D_cache/n1758 , \D_cache/n1757 ,
         \D_cache/n1756 , \D_cache/n1755 , \D_cache/n1754 , \D_cache/n1753 ,
         \D_cache/n1752 , \D_cache/n1751 , \D_cache/n1750 , \D_cache/n1749 ,
         \D_cache/n1748 , \D_cache/n1747 , \D_cache/n1746 , \D_cache/n1745 ,
         \D_cache/n1744 , \D_cache/n1743 , \D_cache/n1742 , \D_cache/n1741 ,
         \D_cache/n1740 , \D_cache/n1739 , \D_cache/n1738 , \D_cache/n1737 ,
         \D_cache/n1736 , \D_cache/n1735 , \D_cache/n1734 , \D_cache/n1733 ,
         \D_cache/n1732 , \D_cache/n1731 , \D_cache/n1730 , \D_cache/n1729 ,
         \D_cache/n1728 , \D_cache/n1727 , \D_cache/n1726 , \D_cache/n1725 ,
         \D_cache/n1724 , \D_cache/n1723 , \D_cache/n1722 , \D_cache/n1721 ,
         \D_cache/n1720 , \D_cache/n1719 , \D_cache/n1718 , \D_cache/n1717 ,
         \D_cache/n1716 , \D_cache/n1715 , \D_cache/n1714 , \D_cache/n1713 ,
         \D_cache/n1712 , \D_cache/n1711 , \D_cache/n1710 , \D_cache/n1709 ,
         \D_cache/n1708 , \D_cache/n1707 , \D_cache/n1706 , \D_cache/n1705 ,
         \D_cache/n1704 , \D_cache/n1703 , \D_cache/n1702 , \D_cache/n1701 ,
         \D_cache/n1700 , \D_cache/n1699 , \D_cache/n1698 , \D_cache/n1697 ,
         \D_cache/n1696 , \D_cache/n1695 , \D_cache/n1694 , \D_cache/n1693 ,
         \D_cache/n1692 , \D_cache/n1691 , \D_cache/n1690 , \D_cache/n1689 ,
         \D_cache/n1688 , \D_cache/n1687 , \D_cache/n1686 , \D_cache/n1685 ,
         \D_cache/n1684 , \D_cache/n1683 , \D_cache/n1682 , \D_cache/n1681 ,
         \D_cache/n1680 , \D_cache/n1679 , \D_cache/n1678 , \D_cache/n1677 ,
         \D_cache/n1676 , \D_cache/n1675 , \D_cache/n1674 , \D_cache/n1673 ,
         \D_cache/n1672 , \D_cache/n1671 , \D_cache/n1670 , \D_cache/n1669 ,
         \D_cache/n1668 , \D_cache/n1667 , \D_cache/n1666 , \D_cache/n1665 ,
         \D_cache/n1664 , \D_cache/n1663 , \D_cache/n1662 , \D_cache/n1661 ,
         \D_cache/n1660 , \D_cache/n1659 , \D_cache/n1658 , \D_cache/n1657 ,
         \D_cache/n1656 , \D_cache/n1655 , \D_cache/n1654 , \D_cache/n1653 ,
         \D_cache/n1652 , \D_cache/n1651 , \D_cache/n1650 , \D_cache/n1649 ,
         \D_cache/n1648 , \D_cache/n1647 , \D_cache/n1646 , \D_cache/n1645 ,
         \D_cache/n1644 , \D_cache/n1643 , \D_cache/n1642 , \D_cache/n1641 ,
         \D_cache/n1640 , \D_cache/n1639 , \D_cache/n1638 , \D_cache/n1637 ,
         \D_cache/n1636 , \D_cache/n1635 , \D_cache/n1634 , \D_cache/n1633 ,
         \D_cache/n1632 , \D_cache/n1631 , \D_cache/n1630 , \D_cache/n1629 ,
         \D_cache/n1628 , \D_cache/n1627 , \D_cache/n1626 , \D_cache/n1625 ,
         \D_cache/n1624 , \D_cache/n1623 , \D_cache/n1622 , \D_cache/n1621 ,
         \D_cache/n1620 , \D_cache/n1619 , \D_cache/n1618 , \D_cache/n1617 ,
         \D_cache/n1616 , \D_cache/n1615 , \D_cache/n1614 , \D_cache/n1613 ,
         \D_cache/n1612 , \D_cache/n1611 , \D_cache/n1610 , \D_cache/n1609 ,
         \D_cache/n1608 , \D_cache/n1607 , \D_cache/n1606 , \D_cache/n1605 ,
         \D_cache/n1604 , \D_cache/n1603 , \D_cache/n1602 , \D_cache/n1601 ,
         \D_cache/n1600 , \D_cache/n1599 , \D_cache/n1598 , \D_cache/n1597 ,
         \D_cache/n1596 , \D_cache/n1595 , \D_cache/n1594 , \D_cache/n1593 ,
         \D_cache/n1592 , \D_cache/n1591 , \D_cache/n1590 , \D_cache/n1589 ,
         \D_cache/n1588 , \D_cache/n1587 , \D_cache/n1586 , \D_cache/n1585 ,
         \D_cache/n1584 , \D_cache/n1583 , \D_cache/n1582 , \D_cache/n1581 ,
         \D_cache/n1580 , \D_cache/n1579 , \D_cache/n1578 , \D_cache/n1577 ,
         \D_cache/n1576 , \D_cache/n1575 , \D_cache/n1574 , \D_cache/n1573 ,
         \D_cache/n1572 , \D_cache/n1571 , \D_cache/n1570 , \D_cache/n1569 ,
         \D_cache/n1568 , \D_cache/n1567 , \D_cache/n1566 , \D_cache/n1565 ,
         \D_cache/n1564 , \D_cache/n1563 , \D_cache/n1562 , \D_cache/n1561 ,
         \D_cache/n1560 , \D_cache/n1559 , \D_cache/n1558 , \D_cache/n1557 ,
         \D_cache/n1556 , \D_cache/n1555 , \D_cache/n1554 , \D_cache/n1553 ,
         \D_cache/n1552 , \D_cache/n1551 , \D_cache/n1550 , \D_cache/n1549 ,
         \D_cache/n1548 , \D_cache/n1547 , \D_cache/n1546 , \D_cache/n1545 ,
         \D_cache/n1544 , \D_cache/n1543 , \D_cache/n1542 , \D_cache/n1541 ,
         \D_cache/n1540 , \D_cache/n1539 , \D_cache/n1538 , \D_cache/n1537 ,
         \D_cache/n1536 , \D_cache/n1535 , \D_cache/n1534 , \D_cache/n1533 ,
         \D_cache/n1532 , \D_cache/n1531 , \D_cache/n1530 , \D_cache/n1529 ,
         \D_cache/n1528 , \D_cache/n1527 , \D_cache/n1526 , \D_cache/n1525 ,
         \D_cache/n1524 , \D_cache/n1523 , \D_cache/n1522 , \D_cache/n1521 ,
         \D_cache/n1520 , \D_cache/n1519 , \D_cache/n1518 , \D_cache/n1517 ,
         \D_cache/n1516 , \D_cache/n1515 , \D_cache/n1514 , \D_cache/n1513 ,
         \D_cache/n1512 , \D_cache/n1511 , \D_cache/n1510 , \D_cache/n1509 ,
         \D_cache/n1508 , \D_cache/n1507 , \D_cache/n1506 , \D_cache/n1505 ,
         \D_cache/n1504 , \D_cache/n1503 , \D_cache/n1502 , \D_cache/n1501 ,
         \D_cache/n1500 , \D_cache/n1499 , \D_cache/n1498 , \D_cache/n1497 ,
         \D_cache/n1496 , \D_cache/n1495 , \D_cache/n1494 , \D_cache/n1493 ,
         \D_cache/n1492 , \D_cache/n1491 , \D_cache/n1490 , \D_cache/n1489 ,
         \D_cache/n1488 , \D_cache/n1487 , \D_cache/n1486 , \D_cache/n1485 ,
         \D_cache/n1484 , \D_cache/n1483 , \D_cache/n1482 , \D_cache/n1481 ,
         \D_cache/n1480 , \D_cache/n1479 , \D_cache/n1478 , \D_cache/n1477 ,
         \D_cache/n1476 , \D_cache/n1475 , \D_cache/n1474 , \D_cache/n1473 ,
         \D_cache/n1472 , \D_cache/n1471 , \D_cache/n1470 , \D_cache/n1469 ,
         \D_cache/n1468 , \D_cache/n1467 , \D_cache/n1466 , \D_cache/n1465 ,
         \D_cache/n1464 , \D_cache/n1463 , \D_cache/n1462 , \D_cache/n1461 ,
         \D_cache/n1460 , \D_cache/n1459 , \D_cache/n1458 , \D_cache/n1457 ,
         \D_cache/n1456 , \D_cache/n1455 , \D_cache/n1454 , \D_cache/n1453 ,
         \D_cache/n1452 , \D_cache/n1451 , \D_cache/n1450 , \D_cache/n1449 ,
         \D_cache/n1448 , \D_cache/n1447 , \D_cache/n1446 , \D_cache/n1445 ,
         \D_cache/n1444 , \D_cache/n1443 , \D_cache/n1442 , \D_cache/n1441 ,
         \D_cache/n1440 , \D_cache/n1439 , \D_cache/n1438 , \D_cache/n1437 ,
         \D_cache/n1436 , \D_cache/n1435 , \D_cache/n1434 , \D_cache/n1433 ,
         \D_cache/n1432 , \D_cache/n1431 , \D_cache/n1430 , \D_cache/n1429 ,
         \D_cache/n1428 , \D_cache/n1427 , \D_cache/n1426 , \D_cache/n1425 ,
         \D_cache/n1424 , \D_cache/n1423 , \D_cache/n1422 , \D_cache/n1421 ,
         \D_cache/n1420 , \D_cache/n1419 , \D_cache/n1418 , \D_cache/n1417 ,
         \D_cache/n1416 , \D_cache/n1415 , \D_cache/n1414 , \D_cache/n1413 ,
         \D_cache/n1412 , \D_cache/n1411 , \D_cache/n1410 , \D_cache/n1409 ,
         \D_cache/n1408 , \D_cache/n1407 , \D_cache/n1406 , \D_cache/n1405 ,
         \D_cache/n1404 , \D_cache/n1403 , \D_cache/n1402 , \D_cache/n1401 ,
         \D_cache/n1400 , \D_cache/n1399 , \D_cache/n1398 , \D_cache/n1397 ,
         \D_cache/n1396 , \D_cache/n1395 , \D_cache/n1394 , \D_cache/n1393 ,
         \D_cache/n1392 , \D_cache/n1391 , \D_cache/n1390 , \D_cache/n1389 ,
         \D_cache/n1388 , \D_cache/n1387 , \D_cache/n1386 , \D_cache/n1385 ,
         \D_cache/n1384 , \D_cache/n1383 , \D_cache/n1382 , \D_cache/n1381 ,
         \D_cache/n1380 , \D_cache/n1379 , \D_cache/n1378 , \D_cache/n1377 ,
         \D_cache/n1376 , \D_cache/n1375 , \D_cache/n1374 , \D_cache/n1373 ,
         \D_cache/n1372 , \D_cache/n1371 , \D_cache/n1370 , \D_cache/n1369 ,
         \D_cache/n1368 , \D_cache/n1367 , \D_cache/n1366 , \D_cache/n1365 ,
         \D_cache/n1364 , \D_cache/n1363 , \D_cache/n1362 , \D_cache/n1361 ,
         \D_cache/n1360 , \D_cache/n1359 , \D_cache/n1358 , \D_cache/n1357 ,
         \D_cache/n1356 , \D_cache/n1355 , \D_cache/n1354 , \D_cache/n1353 ,
         \D_cache/n1352 , \D_cache/n1351 , \D_cache/n1350 , \D_cache/n1349 ,
         \D_cache/n1348 , \D_cache/n1347 , \D_cache/n1346 , \D_cache/n1345 ,
         \D_cache/n1344 , \D_cache/n1343 , \D_cache/n1342 , \D_cache/n1341 ,
         \D_cache/n1340 , \D_cache/n1339 , \D_cache/n1338 , \D_cache/n1337 ,
         \D_cache/n1336 , \D_cache/n1335 , \D_cache/n1334 , \D_cache/n1333 ,
         \D_cache/n1332 , \D_cache/n1331 , \D_cache/n1330 , \D_cache/n1329 ,
         \D_cache/n1328 , \D_cache/n1327 , \D_cache/n1326 , \D_cache/n1325 ,
         \D_cache/n1324 , \D_cache/n1323 , \D_cache/n1322 , \D_cache/n1321 ,
         \D_cache/n1320 , \D_cache/n1319 , \D_cache/n1318 , \D_cache/n1317 ,
         \D_cache/n1316 , \D_cache/n1315 , \D_cache/n1314 , \D_cache/n1313 ,
         \D_cache/n1312 , \D_cache/n1311 , \D_cache/n1310 , \D_cache/n1309 ,
         \D_cache/n1308 , \D_cache/n1307 , \D_cache/n1306 , \D_cache/n1305 ,
         \D_cache/n1304 , \D_cache/n1303 , \D_cache/n1302 , \D_cache/n1301 ,
         \D_cache/n1300 , \D_cache/n1299 , \D_cache/n1298 , \D_cache/n1297 ,
         \D_cache/n1296 , \D_cache/n1295 , \D_cache/n1294 , \D_cache/n1293 ,
         \D_cache/n1292 , \D_cache/n1291 , \D_cache/n1290 , \D_cache/n1289 ,
         \D_cache/n1288 , \D_cache/n1287 , \D_cache/n1286 , \D_cache/n1285 ,
         \D_cache/n1284 , \D_cache/n1283 , \D_cache/n1282 , \D_cache/n1281 ,
         \D_cache/n1280 , \D_cache/n1279 , \D_cache/n1278 , \D_cache/n1277 ,
         \D_cache/n1276 , \D_cache/n1275 , \D_cache/n1274 , \D_cache/n1273 ,
         \D_cache/n1272 , \D_cache/n1271 , \D_cache/n1270 , \D_cache/n1269 ,
         \D_cache/n1268 , \D_cache/n1267 , \D_cache/n1266 , \D_cache/n1265 ,
         \D_cache/n1264 , \D_cache/n1263 , \D_cache/n1262 , \D_cache/n1261 ,
         \D_cache/n1260 , \D_cache/n1259 , \D_cache/n1258 , \D_cache/n1257 ,
         \D_cache/n1256 , \D_cache/n1255 , \D_cache/n1254 , \D_cache/n1253 ,
         \D_cache/n1252 , \D_cache/n1251 , \D_cache/n1250 , \D_cache/n1249 ,
         \D_cache/n1248 , \D_cache/n1247 , \D_cache/n1246 , \D_cache/n1245 ,
         \D_cache/n1244 , \D_cache/n1243 , \D_cache/n1242 , \D_cache/n1241 ,
         \D_cache/n1240 , \D_cache/n1239 , \D_cache/n1238 , \D_cache/n1237 ,
         \D_cache/n1236 , \D_cache/n1235 , \D_cache/n1234 , \D_cache/n1233 ,
         \D_cache/n1232 , \D_cache/n1231 , \D_cache/n1230 , \D_cache/n1229 ,
         \D_cache/n1228 , \D_cache/n1227 , \D_cache/n1226 , \D_cache/n1225 ,
         \D_cache/n1224 , \D_cache/n1223 , \D_cache/n1222 , \D_cache/n1221 ,
         \D_cache/n1220 , \D_cache/n1219 , \D_cache/n1218 , \D_cache/n1217 ,
         \D_cache/n1216 , \D_cache/n1215 , \D_cache/n1214 , \D_cache/n1213 ,
         \D_cache/n1212 , \D_cache/n1211 , \D_cache/n1210 , \D_cache/n1209 ,
         \D_cache/n1208 , \D_cache/n1207 , \D_cache/n1206 , \D_cache/n1205 ,
         \D_cache/n1204 , \D_cache/n1203 , \D_cache/n1202 , \D_cache/n1201 ,
         \D_cache/n1200 , \D_cache/n1199 , \D_cache/n1198 , \D_cache/n1197 ,
         \D_cache/n1196 , \D_cache/n1195 , \D_cache/n1194 , \D_cache/n1193 ,
         \D_cache/n1192 , \D_cache/n1191 , \D_cache/n1190 , \D_cache/n1189 ,
         \D_cache/n1188 , \D_cache/n1187 , \D_cache/n1186 , \D_cache/n1185 ,
         \D_cache/n1184 , \D_cache/n1183 , \D_cache/n1182 , \D_cache/n1181 ,
         \D_cache/n1180 , \D_cache/n1179 , \D_cache/n1178 , \D_cache/n1177 ,
         \D_cache/n1176 , \D_cache/n1175 , \D_cache/n1174 , \D_cache/n1173 ,
         \D_cache/n1172 , \D_cache/n1171 , \D_cache/n1170 , \D_cache/n1169 ,
         \D_cache/n1168 , \D_cache/n1167 , \D_cache/n1166 , \D_cache/n1165 ,
         \D_cache/n1164 , \D_cache/n1163 , \D_cache/n1162 , \D_cache/n1161 ,
         \D_cache/n1160 , \D_cache/n1159 , \D_cache/n1158 , \D_cache/n1157 ,
         \D_cache/n1156 , \D_cache/n1155 , \D_cache/n1154 , \D_cache/n1153 ,
         \D_cache/n1152 , \D_cache/n1151 , \D_cache/n1150 , \D_cache/n1149 ,
         \D_cache/n1148 , \D_cache/n1147 , \D_cache/n1146 , \D_cache/n1145 ,
         \D_cache/n1144 , \D_cache/n1143 , \D_cache/n1142 , \D_cache/n1141 ,
         \D_cache/n1140 , \D_cache/n1139 , \D_cache/n1138 , \D_cache/n1137 ,
         \D_cache/n1136 , \D_cache/n1135 , \D_cache/n1134 , \D_cache/n1133 ,
         \D_cache/n1132 , \D_cache/n1131 , \D_cache/n1130 , \D_cache/n1129 ,
         \D_cache/n1128 , \D_cache/n1127 , \D_cache/n1126 , \D_cache/n1125 ,
         \D_cache/n1124 , \D_cache/n1123 , \D_cache/n1122 , \D_cache/n1121 ,
         \D_cache/n1120 , \D_cache/n1119 , \D_cache/n1118 , \D_cache/n1117 ,
         \D_cache/n1116 , \D_cache/n1115 , \D_cache/n1114 , \D_cache/n1113 ,
         \D_cache/n1112 , \D_cache/n1111 , \D_cache/n1110 , \D_cache/n1109 ,
         \D_cache/n1108 , \D_cache/n1107 , \D_cache/n1106 , \D_cache/n1105 ,
         \D_cache/n1104 , \D_cache/n1103 , \D_cache/n1102 , \D_cache/n1101 ,
         \D_cache/n1100 , \D_cache/n1099 , \D_cache/n1098 , \D_cache/n1097 ,
         \D_cache/n1096 , \D_cache/n1095 , \D_cache/n1094 , \D_cache/n1093 ,
         \D_cache/n1092 , \D_cache/n1091 , \D_cache/n1090 , \D_cache/n1089 ,
         \D_cache/n1088 , \D_cache/n1087 , \D_cache/n1086 , \D_cache/n1085 ,
         \D_cache/n1084 , \D_cache/n1083 , \D_cache/n1082 , \D_cache/n1081 ,
         \D_cache/n1080 , \D_cache/n1079 , \D_cache/n1078 , \D_cache/n1077 ,
         \D_cache/n1076 , \D_cache/n1075 , \D_cache/n1074 , \D_cache/n1073 ,
         \D_cache/n1072 , \D_cache/n1071 , \D_cache/n1070 , \D_cache/n1069 ,
         \D_cache/n1068 , \D_cache/n1067 , \D_cache/n1066 , \D_cache/n1065 ,
         \D_cache/n1064 , \D_cache/n1063 , \D_cache/n1062 , \D_cache/n1061 ,
         \D_cache/n1060 , \D_cache/n1059 , \D_cache/n1058 , \D_cache/n1057 ,
         \D_cache/n1056 , \D_cache/n1055 , \D_cache/n1054 , \D_cache/n1053 ,
         \D_cache/n1052 , \D_cache/n1051 , \D_cache/n1050 , \D_cache/n1049 ,
         \D_cache/n1048 , \D_cache/n1047 , \D_cache/n1046 , \D_cache/n1045 ,
         \D_cache/n1044 , \D_cache/n1043 , \D_cache/n1042 , \D_cache/n1041 ,
         \D_cache/n1040 , \D_cache/n1039 , \D_cache/n1038 , \D_cache/n1037 ,
         \D_cache/n1036 , \D_cache/n1035 , \D_cache/n1034 , \D_cache/n1033 ,
         \D_cache/n1032 , \D_cache/n1031 , \D_cache/n1030 , \D_cache/n1029 ,
         \D_cache/n1028 , \D_cache/n1027 , \D_cache/n1026 , \D_cache/n1025 ,
         \D_cache/n1024 , \D_cache/n1023 , \D_cache/n1022 , \D_cache/n1021 ,
         \D_cache/n1020 , \D_cache/n1019 , \D_cache/n1018 , \D_cache/n1017 ,
         \D_cache/n1016 , \D_cache/n1015 , \D_cache/n1014 , \D_cache/n1013 ,
         \D_cache/n1012 , \D_cache/n1011 , \D_cache/n1010 , \D_cache/n1009 ,
         \D_cache/n1008 , \D_cache/n1007 , \D_cache/n1006 , \D_cache/n1005 ,
         \D_cache/n1004 , \D_cache/n1003 , \D_cache/n1002 , \D_cache/n1001 ,
         \D_cache/n1000 , \D_cache/n999 , \D_cache/n998 , \D_cache/n997 ,
         \D_cache/n996 , \D_cache/n995 , \D_cache/n994 , \D_cache/n993 ,
         \D_cache/n992 , \D_cache/n991 , \D_cache/n990 , \D_cache/n989 ,
         \D_cache/n988 , \D_cache/n987 , \D_cache/n986 , \D_cache/n985 ,
         \D_cache/n984 , \D_cache/n983 , \D_cache/n982 , \D_cache/n981 ,
         \D_cache/n980 , \D_cache/n979 , \D_cache/n978 , \D_cache/n977 ,
         \D_cache/n976 , \D_cache/n975 , \D_cache/n974 , \D_cache/n973 ,
         \D_cache/n972 , \D_cache/n971 , \D_cache/n970 , \D_cache/n969 ,
         \D_cache/n968 , \D_cache/n967 , \D_cache/n966 , \D_cache/n965 ,
         \D_cache/n964 , \D_cache/n963 , \D_cache/n962 , \D_cache/n961 ,
         \D_cache/n960 , \D_cache/n959 , \D_cache/n958 , \D_cache/n957 ,
         \D_cache/n956 , \D_cache/n955 , \D_cache/n954 , \D_cache/n953 ,
         \D_cache/n952 , \D_cache/n951 , \D_cache/n950 , \D_cache/n949 ,
         \D_cache/n948 , \D_cache/n947 , \D_cache/n946 , \D_cache/n945 ,
         \D_cache/n944 , \D_cache/n943 , \D_cache/n942 , \D_cache/n941 ,
         \D_cache/n940 , \D_cache/n939 , \D_cache/n938 , \D_cache/n937 ,
         \D_cache/n936 , \D_cache/n935 , \D_cache/n934 , \D_cache/n933 ,
         \D_cache/n932 , \D_cache/n931 , \D_cache/n930 , \D_cache/n929 ,
         \D_cache/n928 , \D_cache/n927 , \D_cache/n926 , \D_cache/n925 ,
         \D_cache/n924 , \D_cache/n923 , \D_cache/n922 , \D_cache/n921 ,
         \D_cache/n920 , \D_cache/n919 , \D_cache/n918 , \D_cache/n917 ,
         \D_cache/n916 , \D_cache/n915 , \D_cache/n914 , \D_cache/n913 ,
         \D_cache/n912 , \D_cache/n911 , \D_cache/n910 , \D_cache/n909 ,
         \D_cache/n908 , \D_cache/n907 , \D_cache/n906 , \D_cache/n905 ,
         \D_cache/n904 , \D_cache/n903 , \D_cache/n902 , \D_cache/n901 ,
         \D_cache/n900 , \D_cache/n899 , \D_cache/n898 , \D_cache/n897 ,
         \D_cache/n896 , \D_cache/n895 , \D_cache/n894 , \D_cache/n893 ,
         \D_cache/n892 , \D_cache/n891 , \D_cache/n890 , \D_cache/n889 ,
         \D_cache/n888 , \D_cache/n887 , \D_cache/n886 , \D_cache/n885 ,
         \D_cache/n884 , \D_cache/n883 , \D_cache/n882 , \D_cache/n881 ,
         \D_cache/n880 , \D_cache/n879 , \D_cache/n878 , \D_cache/n877 ,
         \D_cache/n876 , \D_cache/n875 , \D_cache/n874 , \D_cache/n873 ,
         \D_cache/n872 , \D_cache/n871 , \D_cache/n870 , \D_cache/n869 ,
         \D_cache/n868 , \D_cache/n867 , \D_cache/n866 , \D_cache/n865 ,
         \D_cache/n864 , \D_cache/n863 , \D_cache/n862 , \D_cache/n861 ,
         \D_cache/n860 , \D_cache/n859 , \D_cache/n858 , \D_cache/n857 ,
         \D_cache/n856 , \D_cache/n855 , \D_cache/n854 , \D_cache/n853 ,
         \D_cache/n852 , \D_cache/n851 , \D_cache/n850 , \D_cache/n849 ,
         \D_cache/n848 , \D_cache/n847 , \D_cache/n846 , \D_cache/n845 ,
         \D_cache/n844 , \D_cache/n843 , \D_cache/n842 , \D_cache/n841 ,
         \D_cache/n840 , \D_cache/n839 , \D_cache/n838 , \D_cache/n837 ,
         \D_cache/n836 , \D_cache/n835 , \D_cache/n834 , \D_cache/n833 ,
         \D_cache/n832 , \D_cache/n831 , \D_cache/n830 , \D_cache/n829 ,
         \D_cache/n828 , \D_cache/n827 , \D_cache/n826 , \D_cache/n825 ,
         \D_cache/n824 , \D_cache/n823 , \D_cache/n822 , \D_cache/n821 ,
         \D_cache/n820 , \D_cache/n819 , \D_cache/n818 , \D_cache/n817 ,
         \D_cache/n816 , \D_cache/n815 , \D_cache/n814 , \D_cache/n813 ,
         \D_cache/n812 , \D_cache/n811 , \D_cache/n810 , \D_cache/n809 ,
         \D_cache/n808 , \D_cache/n807 , \D_cache/n806 , \D_cache/n805 ,
         \D_cache/n804 , \D_cache/n803 , \D_cache/n802 , \D_cache/n801 ,
         \D_cache/n800 , \D_cache/n799 , \D_cache/n798 , \D_cache/n797 ,
         \D_cache/n796 , \D_cache/n795 , \D_cache/n794 , \D_cache/n793 ,
         \D_cache/n792 , \D_cache/n791 , \D_cache/n790 , \D_cache/n789 ,
         \D_cache/n788 , \D_cache/n787 , \D_cache/n786 , \D_cache/n785 ,
         \D_cache/n784 , \D_cache/n783 , \D_cache/n782 , \D_cache/n781 ,
         \D_cache/n780 , \D_cache/n779 , \D_cache/n778 , \D_cache/n777 ,
         \D_cache/n776 , \D_cache/n775 , \D_cache/n774 , \D_cache/n773 ,
         \D_cache/n772 , \D_cache/n771 , \D_cache/n770 , \D_cache/n769 ,
         \D_cache/n768 , \D_cache/n767 , \D_cache/n766 , \D_cache/n765 ,
         \D_cache/n764 , \D_cache/n763 , \D_cache/n762 , \D_cache/n761 ,
         \D_cache/n760 , \D_cache/n759 , \D_cache/n758 , \D_cache/n757 ,
         \D_cache/n756 , \D_cache/n755 , \D_cache/n754 , \D_cache/n753 ,
         \D_cache/n752 , \D_cache/n751 , \D_cache/n750 , \D_cache/n749 ,
         \D_cache/n748 , \D_cache/n747 , \D_cache/n746 , \D_cache/n745 ,
         \D_cache/n744 , \D_cache/n743 , \D_cache/n742 , \D_cache/n741 ,
         \D_cache/n740 , \D_cache/n739 , \D_cache/n738 , \D_cache/n737 ,
         \D_cache/n736 , \D_cache/n735 , \D_cache/n734 , \D_cache/n733 ,
         \D_cache/n732 , \D_cache/n731 , \D_cache/n730 , \D_cache/n729 ,
         \D_cache/n728 , \D_cache/n727 , \D_cache/n726 , \D_cache/n725 ,
         \D_cache/n724 , \D_cache/n723 , \D_cache/n722 , \D_cache/n721 ,
         \D_cache/n720 , \D_cache/n719 , \D_cache/n718 , \D_cache/n717 ,
         \D_cache/n716 , \D_cache/n715 , \D_cache/n714 , \D_cache/n713 ,
         \D_cache/n712 , \D_cache/n711 , \D_cache/n710 , \D_cache/n709 ,
         \D_cache/n708 , \D_cache/n707 , \D_cache/n706 , \D_cache/n705 ,
         \D_cache/n704 , \D_cache/n703 , \D_cache/n702 , \D_cache/n701 ,
         \D_cache/n700 , \D_cache/n699 , \D_cache/n698 , \D_cache/n697 ,
         \D_cache/n696 , \D_cache/n695 , \D_cache/n694 , \D_cache/n693 ,
         \D_cache/n692 , \D_cache/n691 , \D_cache/n690 , \D_cache/n689 ,
         \D_cache/n688 , \D_cache/n687 , \D_cache/n686 , \D_cache/n685 ,
         \D_cache/n684 , \D_cache/n683 , \D_cache/n682 , \D_cache/n681 ,
         \D_cache/n680 , \D_cache/n679 , \D_cache/n678 , \D_cache/n677 ,
         \D_cache/n676 , \D_cache/n675 , \D_cache/n674 , \D_cache/n673 ,
         \D_cache/n672 , \D_cache/n671 , \D_cache/n670 , \D_cache/n669 ,
         \D_cache/n668 , \D_cache/n667 , \D_cache/n666 , \D_cache/n665 ,
         \D_cache/n664 , \D_cache/n663 , \D_cache/n662 , \D_cache/n661 ,
         \D_cache/n660 , \D_cache/n659 , \D_cache/n658 , \D_cache/n657 ,
         \D_cache/n656 , \D_cache/n655 , \D_cache/n654 , \D_cache/n653 ,
         \D_cache/n652 , \D_cache/n651 , \D_cache/n650 , \D_cache/n649 ,
         \D_cache/n648 , \D_cache/n647 , \D_cache/n646 , \D_cache/n645 ,
         \D_cache/n644 , \D_cache/n643 , \D_cache/n642 , \D_cache/n641 ,
         \D_cache/n640 , \D_cache/n639 , \D_cache/n638 , \D_cache/n637 ,
         \D_cache/n636 , \D_cache/n635 , \D_cache/n634 , \D_cache/n633 ,
         \D_cache/n632 , \D_cache/n631 , \D_cache/n630 , \D_cache/n629 ,
         \D_cache/n628 , \D_cache/n627 , \D_cache/n626 , \D_cache/n625 ,
         \D_cache/n624 , \D_cache/n623 , \D_cache/n622 , \D_cache/n621 ,
         \D_cache/n620 , \D_cache/n619 , \D_cache/n618 , \D_cache/n617 ,
         \D_cache/n616 , \D_cache/n615 , \D_cache/n614 , \D_cache/n613 ,
         \D_cache/n612 , \D_cache/n611 , \D_cache/n610 , \D_cache/n609 ,
         \D_cache/n608 , \D_cache/n607 , \D_cache/n606 , \D_cache/n605 ,
         \D_cache/n604 , \D_cache/n603 , \D_cache/n602 , \D_cache/n601 ,
         \D_cache/n600 , \D_cache/n599 , \D_cache/n598 , \D_cache/n597 ,
         \D_cache/n596 , \D_cache/n595 , \D_cache/n594 , \D_cache/n593 ,
         \D_cache/n592 , \D_cache/n591 , \D_cache/n590 , \D_cache/n589 ,
         \D_cache/n588 , \D_cache/n587 , \D_cache/n586 , \D_cache/n585 ,
         \D_cache/n584 , \D_cache/n583 , \D_cache/n582 , \D_cache/n581 ,
         \D_cache/n580 , \D_cache/n579 , \D_cache/n578 , \D_cache/n577 ,
         \D_cache/n576 , \D_cache/n575 , \D_cache/n574 , \D_cache/n573 ,
         \D_cache/n572 , \D_cache/n571 , \D_cache/n570 , \D_cache/n569 ,
         \D_cache/n568 , \D_cache/n567 , \D_cache/n566 , \D_cache/n565 ,
         \D_cache/n564 , \D_cache/n563 , \D_cache/n562 , \D_cache/n561 ,
         \D_cache/n560 , \D_cache/n559 , \D_cache/n558 , \D_cache/n557 ,
         \D_cache/cache[7][0] , \D_cache/cache[7][1] , \D_cache/cache[7][2] ,
         \D_cache/cache[7][3] , \D_cache/cache[7][4] , \D_cache/cache[7][5] ,
         \D_cache/cache[7][6] , \D_cache/cache[7][7] , \D_cache/cache[7][8] ,
         \D_cache/cache[7][9] , \D_cache/cache[7][10] , \D_cache/cache[7][11] ,
         \D_cache/cache[7][12] , \D_cache/cache[7][13] ,
         \D_cache/cache[7][14] , \D_cache/cache[7][15] ,
         \D_cache/cache[7][16] , \D_cache/cache[7][17] ,
         \D_cache/cache[7][18] , \D_cache/cache[7][19] ,
         \D_cache/cache[7][20] , \D_cache/cache[7][21] ,
         \D_cache/cache[7][22] , \D_cache/cache[7][23] ,
         \D_cache/cache[7][24] , \D_cache/cache[7][25] ,
         \D_cache/cache[7][26] , \D_cache/cache[7][27] ,
         \D_cache/cache[7][28] , \D_cache/cache[7][29] ,
         \D_cache/cache[7][30] , \D_cache/cache[7][31] ,
         \D_cache/cache[7][32] , \D_cache/cache[7][33] ,
         \D_cache/cache[7][34] , \D_cache/cache[7][35] ,
         \D_cache/cache[7][36] , \D_cache/cache[7][37] ,
         \D_cache/cache[7][38] , \D_cache/cache[7][39] ,
         \D_cache/cache[7][40] , \D_cache/cache[7][41] ,
         \D_cache/cache[7][42] , \D_cache/cache[7][43] ,
         \D_cache/cache[7][44] , \D_cache/cache[7][45] ,
         \D_cache/cache[7][46] , \D_cache/cache[7][47] ,
         \D_cache/cache[7][48] , \D_cache/cache[7][49] ,
         \D_cache/cache[7][50] , \D_cache/cache[7][51] ,
         \D_cache/cache[7][52] , \D_cache/cache[7][53] ,
         \D_cache/cache[7][54] , \D_cache/cache[7][55] ,
         \D_cache/cache[7][56] , \D_cache/cache[7][57] ,
         \D_cache/cache[7][58] , \D_cache/cache[7][59] ,
         \D_cache/cache[7][60] , \D_cache/cache[7][61] ,
         \D_cache/cache[7][62] , \D_cache/cache[7][63] ,
         \D_cache/cache[7][64] , \D_cache/cache[7][65] ,
         \D_cache/cache[7][66] , \D_cache/cache[7][67] ,
         \D_cache/cache[7][68] , \D_cache/cache[7][69] ,
         \D_cache/cache[7][70] , \D_cache/cache[7][71] ,
         \D_cache/cache[7][72] , \D_cache/cache[7][73] ,
         \D_cache/cache[7][74] , \D_cache/cache[7][75] ,
         \D_cache/cache[7][76] , \D_cache/cache[7][77] ,
         \D_cache/cache[7][78] , \D_cache/cache[7][79] ,
         \D_cache/cache[7][80] , \D_cache/cache[7][81] ,
         \D_cache/cache[7][82] , \D_cache/cache[7][83] ,
         \D_cache/cache[7][84] , \D_cache/cache[7][85] ,
         \D_cache/cache[7][86] , \D_cache/cache[7][87] ,
         \D_cache/cache[7][88] , \D_cache/cache[7][89] ,
         \D_cache/cache[7][90] , \D_cache/cache[7][91] ,
         \D_cache/cache[7][92] , \D_cache/cache[7][93] ,
         \D_cache/cache[7][94] , \D_cache/cache[7][95] ,
         \D_cache/cache[7][96] , \D_cache/cache[7][97] ,
         \D_cache/cache[7][98] , \D_cache/cache[7][99] ,
         \D_cache/cache[7][100] , \D_cache/cache[7][101] ,
         \D_cache/cache[7][102] , \D_cache/cache[7][103] ,
         \D_cache/cache[7][104] , \D_cache/cache[7][105] ,
         \D_cache/cache[7][106] , \D_cache/cache[7][107] ,
         \D_cache/cache[7][108] , \D_cache/cache[7][109] ,
         \D_cache/cache[7][110] , \D_cache/cache[7][111] ,
         \D_cache/cache[7][112] , \D_cache/cache[7][113] ,
         \D_cache/cache[7][114] , \D_cache/cache[7][115] ,
         \D_cache/cache[7][116] , \D_cache/cache[7][117] ,
         \D_cache/cache[7][118] , \D_cache/cache[7][119] ,
         \D_cache/cache[7][120] , \D_cache/cache[7][121] ,
         \D_cache/cache[7][122] , \D_cache/cache[7][123] ,
         \D_cache/cache[7][124] , \D_cache/cache[7][125] ,
         \D_cache/cache[7][126] , \D_cache/cache[7][127] ,
         \D_cache/cache[7][128] , \D_cache/cache[7][129] ,
         \D_cache/cache[7][130] , \D_cache/cache[7][131] ,
         \D_cache/cache[7][132] , \D_cache/cache[7][133] ,
         \D_cache/cache[7][134] , \D_cache/cache[7][135] ,
         \D_cache/cache[7][136] , \D_cache/cache[7][137] ,
         \D_cache/cache[7][138] , \D_cache/cache[7][139] ,
         \D_cache/cache[7][140] , \D_cache/cache[7][141] ,
         \D_cache/cache[7][142] , \D_cache/cache[7][143] ,
         \D_cache/cache[7][144] , \D_cache/cache[7][145] ,
         \D_cache/cache[7][146] , \D_cache/cache[7][147] ,
         \D_cache/cache[7][148] , \D_cache/cache[7][149] ,
         \D_cache/cache[7][150] , \D_cache/cache[7][151] ,
         \D_cache/cache[7][152] , \D_cache/cache[7][153] ,
         \D_cache/cache[7][154] , \D_cache/cache[6][0] , \D_cache/cache[6][1] ,
         \D_cache/cache[6][2] , \D_cache/cache[6][3] , \D_cache/cache[6][4] ,
         \D_cache/cache[6][5] , \D_cache/cache[6][6] , \D_cache/cache[6][7] ,
         \D_cache/cache[6][8] , \D_cache/cache[6][9] , \D_cache/cache[6][10] ,
         \D_cache/cache[6][11] , \D_cache/cache[6][12] ,
         \D_cache/cache[6][13] , \D_cache/cache[6][14] ,
         \D_cache/cache[6][15] , \D_cache/cache[6][16] ,
         \D_cache/cache[6][17] , \D_cache/cache[6][18] ,
         \D_cache/cache[6][19] , \D_cache/cache[6][20] ,
         \D_cache/cache[6][21] , \D_cache/cache[6][22] ,
         \D_cache/cache[6][23] , \D_cache/cache[6][24] ,
         \D_cache/cache[6][25] , \D_cache/cache[6][26] ,
         \D_cache/cache[6][27] , \D_cache/cache[6][28] ,
         \D_cache/cache[6][29] , \D_cache/cache[6][30] ,
         \D_cache/cache[6][31] , \D_cache/cache[6][32] ,
         \D_cache/cache[6][33] , \D_cache/cache[6][34] ,
         \D_cache/cache[6][35] , \D_cache/cache[6][36] ,
         \D_cache/cache[6][37] , \D_cache/cache[6][38] ,
         \D_cache/cache[6][39] , \D_cache/cache[6][40] ,
         \D_cache/cache[6][41] , \D_cache/cache[6][42] ,
         \D_cache/cache[6][43] , \D_cache/cache[6][44] ,
         \D_cache/cache[6][45] , \D_cache/cache[6][46] ,
         \D_cache/cache[6][47] , \D_cache/cache[6][48] ,
         \D_cache/cache[6][49] , \D_cache/cache[6][50] ,
         \D_cache/cache[6][51] , \D_cache/cache[6][52] ,
         \D_cache/cache[6][53] , \D_cache/cache[6][54] ,
         \D_cache/cache[6][55] , \D_cache/cache[6][56] ,
         \D_cache/cache[6][57] , \D_cache/cache[6][58] ,
         \D_cache/cache[6][59] , \D_cache/cache[6][60] ,
         \D_cache/cache[6][61] , \D_cache/cache[6][62] ,
         \D_cache/cache[6][63] , \D_cache/cache[6][64] ,
         \D_cache/cache[6][65] , \D_cache/cache[6][66] ,
         \D_cache/cache[6][67] , \D_cache/cache[6][68] ,
         \D_cache/cache[6][69] , \D_cache/cache[6][70] ,
         \D_cache/cache[6][71] , \D_cache/cache[6][72] ,
         \D_cache/cache[6][73] , \D_cache/cache[6][74] ,
         \D_cache/cache[6][75] , \D_cache/cache[6][76] ,
         \D_cache/cache[6][77] , \D_cache/cache[6][78] ,
         \D_cache/cache[6][79] , \D_cache/cache[6][80] ,
         \D_cache/cache[6][81] , \D_cache/cache[6][82] ,
         \D_cache/cache[6][83] , \D_cache/cache[6][84] ,
         \D_cache/cache[6][85] , \D_cache/cache[6][86] ,
         \D_cache/cache[6][87] , \D_cache/cache[6][88] ,
         \D_cache/cache[6][89] , \D_cache/cache[6][90] ,
         \D_cache/cache[6][91] , \D_cache/cache[6][92] ,
         \D_cache/cache[6][93] , \D_cache/cache[6][94] ,
         \D_cache/cache[6][95] , \D_cache/cache[6][96] ,
         \D_cache/cache[6][97] , \D_cache/cache[6][98] ,
         \D_cache/cache[6][99] , \D_cache/cache[6][100] ,
         \D_cache/cache[6][101] , \D_cache/cache[6][102] ,
         \D_cache/cache[6][103] , \D_cache/cache[6][104] ,
         \D_cache/cache[6][105] , \D_cache/cache[6][106] ,
         \D_cache/cache[6][107] , \D_cache/cache[6][108] ,
         \D_cache/cache[6][109] , \D_cache/cache[6][110] ,
         \D_cache/cache[6][111] , \D_cache/cache[6][112] ,
         \D_cache/cache[6][113] , \D_cache/cache[6][114] ,
         \D_cache/cache[6][115] , \D_cache/cache[6][116] ,
         \D_cache/cache[6][117] , \D_cache/cache[6][118] ,
         \D_cache/cache[6][119] , \D_cache/cache[6][120] ,
         \D_cache/cache[6][121] , \D_cache/cache[6][122] ,
         \D_cache/cache[6][123] , \D_cache/cache[6][124] ,
         \D_cache/cache[6][125] , \D_cache/cache[6][126] ,
         \D_cache/cache[6][127] , \D_cache/cache[6][128] ,
         \D_cache/cache[6][129] , \D_cache/cache[6][130] ,
         \D_cache/cache[6][131] , \D_cache/cache[6][132] ,
         \D_cache/cache[6][133] , \D_cache/cache[6][134] ,
         \D_cache/cache[6][135] , \D_cache/cache[6][136] ,
         \D_cache/cache[6][137] , \D_cache/cache[6][138] ,
         \D_cache/cache[6][139] , \D_cache/cache[6][140] ,
         \D_cache/cache[6][141] , \D_cache/cache[6][142] ,
         \D_cache/cache[6][143] , \D_cache/cache[6][144] ,
         \D_cache/cache[6][145] , \D_cache/cache[6][146] ,
         \D_cache/cache[6][147] , \D_cache/cache[6][148] ,
         \D_cache/cache[6][149] , \D_cache/cache[6][150] ,
         \D_cache/cache[6][151] , \D_cache/cache[6][152] ,
         \D_cache/cache[6][153] , \D_cache/cache[6][154] ,
         \D_cache/cache[5][0] , \D_cache/cache[5][1] , \D_cache/cache[5][2] ,
         \D_cache/cache[5][3] , \D_cache/cache[5][4] , \D_cache/cache[5][5] ,
         \D_cache/cache[5][6] , \D_cache/cache[5][7] , \D_cache/cache[5][8] ,
         \D_cache/cache[5][9] , \D_cache/cache[5][10] , \D_cache/cache[5][11] ,
         \D_cache/cache[5][12] , \D_cache/cache[5][13] ,
         \D_cache/cache[5][14] , \D_cache/cache[5][15] ,
         \D_cache/cache[5][16] , \D_cache/cache[5][17] ,
         \D_cache/cache[5][18] , \D_cache/cache[5][19] ,
         \D_cache/cache[5][20] , \D_cache/cache[5][21] ,
         \D_cache/cache[5][22] , \D_cache/cache[5][23] ,
         \D_cache/cache[5][24] , \D_cache/cache[5][25] ,
         \D_cache/cache[5][26] , \D_cache/cache[5][27] ,
         \D_cache/cache[5][28] , \D_cache/cache[5][29] ,
         \D_cache/cache[5][30] , \D_cache/cache[5][31] ,
         \D_cache/cache[5][32] , \D_cache/cache[5][33] ,
         \D_cache/cache[5][34] , \D_cache/cache[5][35] ,
         \D_cache/cache[5][36] , \D_cache/cache[5][37] ,
         \D_cache/cache[5][38] , \D_cache/cache[5][39] ,
         \D_cache/cache[5][40] , \D_cache/cache[5][41] ,
         \D_cache/cache[5][42] , \D_cache/cache[5][43] ,
         \D_cache/cache[5][44] , \D_cache/cache[5][45] ,
         \D_cache/cache[5][46] , \D_cache/cache[5][47] ,
         \D_cache/cache[5][48] , \D_cache/cache[5][49] ,
         \D_cache/cache[5][50] , \D_cache/cache[5][51] ,
         \D_cache/cache[5][52] , \D_cache/cache[5][53] ,
         \D_cache/cache[5][54] , \D_cache/cache[5][55] ,
         \D_cache/cache[5][56] , \D_cache/cache[5][57] ,
         \D_cache/cache[5][58] , \D_cache/cache[5][59] ,
         \D_cache/cache[5][60] , \D_cache/cache[5][61] ,
         \D_cache/cache[5][62] , \D_cache/cache[5][63] ,
         \D_cache/cache[5][64] , \D_cache/cache[5][65] ,
         \D_cache/cache[5][66] , \D_cache/cache[5][67] ,
         \D_cache/cache[5][68] , \D_cache/cache[5][69] ,
         \D_cache/cache[5][70] , \D_cache/cache[5][71] ,
         \D_cache/cache[5][72] , \D_cache/cache[5][73] ,
         \D_cache/cache[5][74] , \D_cache/cache[5][75] ,
         \D_cache/cache[5][76] , \D_cache/cache[5][77] ,
         \D_cache/cache[5][78] , \D_cache/cache[5][79] ,
         \D_cache/cache[5][80] , \D_cache/cache[5][81] ,
         \D_cache/cache[5][82] , \D_cache/cache[5][83] ,
         \D_cache/cache[5][84] , \D_cache/cache[5][85] ,
         \D_cache/cache[5][86] , \D_cache/cache[5][87] ,
         \D_cache/cache[5][88] , \D_cache/cache[5][89] ,
         \D_cache/cache[5][90] , \D_cache/cache[5][91] ,
         \D_cache/cache[5][92] , \D_cache/cache[5][93] ,
         \D_cache/cache[5][94] , \D_cache/cache[5][95] ,
         \D_cache/cache[5][96] , \D_cache/cache[5][97] ,
         \D_cache/cache[5][98] , \D_cache/cache[5][99] ,
         \D_cache/cache[5][100] , \D_cache/cache[5][101] ,
         \D_cache/cache[5][102] , \D_cache/cache[5][103] ,
         \D_cache/cache[5][104] , \D_cache/cache[5][105] ,
         \D_cache/cache[5][106] , \D_cache/cache[5][107] ,
         \D_cache/cache[5][108] , \D_cache/cache[5][109] ,
         \D_cache/cache[5][110] , \D_cache/cache[5][111] ,
         \D_cache/cache[5][112] , \D_cache/cache[5][113] ,
         \D_cache/cache[5][114] , \D_cache/cache[5][115] ,
         \D_cache/cache[5][116] , \D_cache/cache[5][117] ,
         \D_cache/cache[5][118] , \D_cache/cache[5][119] ,
         \D_cache/cache[5][120] , \D_cache/cache[5][121] ,
         \D_cache/cache[5][122] , \D_cache/cache[5][123] ,
         \D_cache/cache[5][124] , \D_cache/cache[5][125] ,
         \D_cache/cache[5][126] , \D_cache/cache[5][127] ,
         \D_cache/cache[5][128] , \D_cache/cache[5][129] ,
         \D_cache/cache[5][130] , \D_cache/cache[5][131] ,
         \D_cache/cache[5][132] , \D_cache/cache[5][133] ,
         \D_cache/cache[5][134] , \D_cache/cache[5][135] ,
         \D_cache/cache[5][136] , \D_cache/cache[5][137] ,
         \D_cache/cache[5][138] , \D_cache/cache[5][139] ,
         \D_cache/cache[5][140] , \D_cache/cache[5][141] ,
         \D_cache/cache[5][142] , \D_cache/cache[5][143] ,
         \D_cache/cache[5][144] , \D_cache/cache[5][145] ,
         \D_cache/cache[5][146] , \D_cache/cache[5][147] ,
         \D_cache/cache[5][148] , \D_cache/cache[5][149] ,
         \D_cache/cache[5][150] , \D_cache/cache[5][151] ,
         \D_cache/cache[5][152] , \D_cache/cache[5][153] ,
         \D_cache/cache[5][154] , \D_cache/cache[4][0] , \D_cache/cache[4][1] ,
         \D_cache/cache[4][2] , \D_cache/cache[4][3] , \D_cache/cache[4][4] ,
         \D_cache/cache[4][5] , \D_cache/cache[4][6] , \D_cache/cache[4][7] ,
         \D_cache/cache[4][8] , \D_cache/cache[4][9] , \D_cache/cache[4][10] ,
         \D_cache/cache[4][11] , \D_cache/cache[4][12] ,
         \D_cache/cache[4][13] , \D_cache/cache[4][14] ,
         \D_cache/cache[4][15] , \D_cache/cache[4][16] ,
         \D_cache/cache[4][17] , \D_cache/cache[4][18] ,
         \D_cache/cache[4][19] , \D_cache/cache[4][20] ,
         \D_cache/cache[4][21] , \D_cache/cache[4][22] ,
         \D_cache/cache[4][23] , \D_cache/cache[4][24] ,
         \D_cache/cache[4][25] , \D_cache/cache[4][26] ,
         \D_cache/cache[4][27] , \D_cache/cache[4][28] ,
         \D_cache/cache[4][29] , \D_cache/cache[4][30] ,
         \D_cache/cache[4][31] , \D_cache/cache[4][32] ,
         \D_cache/cache[4][33] , \D_cache/cache[4][34] ,
         \D_cache/cache[4][35] , \D_cache/cache[4][36] ,
         \D_cache/cache[4][37] , \D_cache/cache[4][38] ,
         \D_cache/cache[4][39] , \D_cache/cache[4][40] ,
         \D_cache/cache[4][41] , \D_cache/cache[4][42] ,
         \D_cache/cache[4][43] , \D_cache/cache[4][44] ,
         \D_cache/cache[4][45] , \D_cache/cache[4][46] ,
         \D_cache/cache[4][47] , \D_cache/cache[4][48] ,
         \D_cache/cache[4][49] , \D_cache/cache[4][50] ,
         \D_cache/cache[4][51] , \D_cache/cache[4][52] ,
         \D_cache/cache[4][53] , \D_cache/cache[4][54] ,
         \D_cache/cache[4][55] , \D_cache/cache[4][56] ,
         \D_cache/cache[4][57] , \D_cache/cache[4][58] ,
         \D_cache/cache[4][59] , \D_cache/cache[4][60] ,
         \D_cache/cache[4][61] , \D_cache/cache[4][62] ,
         \D_cache/cache[4][63] , \D_cache/cache[4][64] ,
         \D_cache/cache[4][65] , \D_cache/cache[4][66] ,
         \D_cache/cache[4][67] , \D_cache/cache[4][68] ,
         \D_cache/cache[4][69] , \D_cache/cache[4][70] ,
         \D_cache/cache[4][71] , \D_cache/cache[4][72] ,
         \D_cache/cache[4][73] , \D_cache/cache[4][74] ,
         \D_cache/cache[4][75] , \D_cache/cache[4][76] ,
         \D_cache/cache[4][77] , \D_cache/cache[4][78] ,
         \D_cache/cache[4][79] , \D_cache/cache[4][80] ,
         \D_cache/cache[4][81] , \D_cache/cache[4][82] ,
         \D_cache/cache[4][83] , \D_cache/cache[4][84] ,
         \D_cache/cache[4][85] , \D_cache/cache[4][86] ,
         \D_cache/cache[4][87] , \D_cache/cache[4][88] ,
         \D_cache/cache[4][89] , \D_cache/cache[4][90] ,
         \D_cache/cache[4][91] , \D_cache/cache[4][92] ,
         \D_cache/cache[4][93] , \D_cache/cache[4][94] ,
         \D_cache/cache[4][95] , \D_cache/cache[4][96] ,
         \D_cache/cache[4][97] , \D_cache/cache[4][98] ,
         \D_cache/cache[4][99] , \D_cache/cache[4][100] ,
         \D_cache/cache[4][101] , \D_cache/cache[4][102] ,
         \D_cache/cache[4][103] , \D_cache/cache[4][104] ,
         \D_cache/cache[4][105] , \D_cache/cache[4][106] ,
         \D_cache/cache[4][107] , \D_cache/cache[4][108] ,
         \D_cache/cache[4][109] , \D_cache/cache[4][110] ,
         \D_cache/cache[4][111] , \D_cache/cache[4][112] ,
         \D_cache/cache[4][113] , \D_cache/cache[4][114] ,
         \D_cache/cache[4][115] , \D_cache/cache[4][116] ,
         \D_cache/cache[4][117] , \D_cache/cache[4][118] ,
         \D_cache/cache[4][119] , \D_cache/cache[4][120] ,
         \D_cache/cache[4][121] , \D_cache/cache[4][122] ,
         \D_cache/cache[4][123] , \D_cache/cache[4][124] ,
         \D_cache/cache[4][125] , \D_cache/cache[4][126] ,
         \D_cache/cache[4][127] , \D_cache/cache[4][128] ,
         \D_cache/cache[4][129] , \D_cache/cache[4][130] ,
         \D_cache/cache[4][131] , \D_cache/cache[4][132] ,
         \D_cache/cache[4][133] , \D_cache/cache[4][134] ,
         \D_cache/cache[4][135] , \D_cache/cache[4][136] ,
         \D_cache/cache[4][137] , \D_cache/cache[4][138] ,
         \D_cache/cache[4][139] , \D_cache/cache[4][140] ,
         \D_cache/cache[4][141] , \D_cache/cache[4][142] ,
         \D_cache/cache[4][143] , \D_cache/cache[4][144] ,
         \D_cache/cache[4][145] , \D_cache/cache[4][146] ,
         \D_cache/cache[4][147] , \D_cache/cache[4][148] ,
         \D_cache/cache[4][149] , \D_cache/cache[4][150] ,
         \D_cache/cache[4][151] , \D_cache/cache[4][152] ,
         \D_cache/cache[4][153] , \D_cache/cache[4][154] ,
         \D_cache/cache[3][0] , \D_cache/cache[3][1] , \D_cache/cache[3][2] ,
         \D_cache/cache[3][3] , \D_cache/cache[3][4] , \D_cache/cache[3][5] ,
         \D_cache/cache[3][6] , \D_cache/cache[3][7] , \D_cache/cache[3][8] ,
         \D_cache/cache[3][9] , \D_cache/cache[3][10] , \D_cache/cache[3][11] ,
         \D_cache/cache[3][12] , \D_cache/cache[3][13] ,
         \D_cache/cache[3][14] , \D_cache/cache[3][15] ,
         \D_cache/cache[3][16] , \D_cache/cache[3][17] ,
         \D_cache/cache[3][18] , \D_cache/cache[3][19] ,
         \D_cache/cache[3][20] , \D_cache/cache[3][21] ,
         \D_cache/cache[3][22] , \D_cache/cache[3][23] ,
         \D_cache/cache[3][24] , \D_cache/cache[3][25] ,
         \D_cache/cache[3][26] , \D_cache/cache[3][27] ,
         \D_cache/cache[3][28] , \D_cache/cache[3][29] ,
         \D_cache/cache[3][30] , \D_cache/cache[3][31] ,
         \D_cache/cache[3][32] , \D_cache/cache[3][33] ,
         \D_cache/cache[3][34] , \D_cache/cache[3][35] ,
         \D_cache/cache[3][36] , \D_cache/cache[3][37] ,
         \D_cache/cache[3][38] , \D_cache/cache[3][39] ,
         \D_cache/cache[3][40] , \D_cache/cache[3][41] ,
         \D_cache/cache[3][42] , \D_cache/cache[3][43] ,
         \D_cache/cache[3][44] , \D_cache/cache[3][45] ,
         \D_cache/cache[3][46] , \D_cache/cache[3][47] ,
         \D_cache/cache[3][48] , \D_cache/cache[3][49] ,
         \D_cache/cache[3][50] , \D_cache/cache[3][51] ,
         \D_cache/cache[3][52] , \D_cache/cache[3][53] ,
         \D_cache/cache[3][54] , \D_cache/cache[3][55] ,
         \D_cache/cache[3][56] , \D_cache/cache[3][57] ,
         \D_cache/cache[3][58] , \D_cache/cache[3][59] ,
         \D_cache/cache[3][60] , \D_cache/cache[3][61] ,
         \D_cache/cache[3][62] , \D_cache/cache[3][63] ,
         \D_cache/cache[3][64] , \D_cache/cache[3][65] ,
         \D_cache/cache[3][66] , \D_cache/cache[3][67] ,
         \D_cache/cache[3][68] , \D_cache/cache[3][69] ,
         \D_cache/cache[3][70] , \D_cache/cache[3][71] ,
         \D_cache/cache[3][72] , \D_cache/cache[3][73] ,
         \D_cache/cache[3][74] , \D_cache/cache[3][75] ,
         \D_cache/cache[3][76] , \D_cache/cache[3][77] ,
         \D_cache/cache[3][78] , \D_cache/cache[3][79] ,
         \D_cache/cache[3][80] , \D_cache/cache[3][81] ,
         \D_cache/cache[3][82] , \D_cache/cache[3][83] ,
         \D_cache/cache[3][84] , \D_cache/cache[3][85] ,
         \D_cache/cache[3][86] , \D_cache/cache[3][87] ,
         \D_cache/cache[3][88] , \D_cache/cache[3][89] ,
         \D_cache/cache[3][90] , \D_cache/cache[3][91] ,
         \D_cache/cache[3][92] , \D_cache/cache[3][93] ,
         \D_cache/cache[3][94] , \D_cache/cache[3][95] ,
         \D_cache/cache[3][96] , \D_cache/cache[3][97] ,
         \D_cache/cache[3][98] , \D_cache/cache[3][99] ,
         \D_cache/cache[3][100] , \D_cache/cache[3][101] ,
         \D_cache/cache[3][102] , \D_cache/cache[3][103] ,
         \D_cache/cache[3][104] , \D_cache/cache[3][105] ,
         \D_cache/cache[3][106] , \D_cache/cache[3][107] ,
         \D_cache/cache[3][108] , \D_cache/cache[3][109] ,
         \D_cache/cache[3][110] , \D_cache/cache[3][111] ,
         \D_cache/cache[3][112] , \D_cache/cache[3][113] ,
         \D_cache/cache[3][114] , \D_cache/cache[3][115] ,
         \D_cache/cache[3][116] , \D_cache/cache[3][117] ,
         \D_cache/cache[3][118] , \D_cache/cache[3][119] ,
         \D_cache/cache[3][120] , \D_cache/cache[3][121] ,
         \D_cache/cache[3][122] , \D_cache/cache[3][123] ,
         \D_cache/cache[3][124] , \D_cache/cache[3][125] ,
         \D_cache/cache[3][126] , \D_cache/cache[3][127] ,
         \D_cache/cache[3][128] , \D_cache/cache[3][129] ,
         \D_cache/cache[3][130] , \D_cache/cache[3][131] ,
         \D_cache/cache[3][132] , \D_cache/cache[3][133] ,
         \D_cache/cache[3][134] , \D_cache/cache[3][135] ,
         \D_cache/cache[3][136] , \D_cache/cache[3][137] ,
         \D_cache/cache[3][138] , \D_cache/cache[3][139] ,
         \D_cache/cache[3][140] , \D_cache/cache[3][141] ,
         \D_cache/cache[3][142] , \D_cache/cache[3][143] ,
         \D_cache/cache[3][144] , \D_cache/cache[3][145] ,
         \D_cache/cache[3][146] , \D_cache/cache[3][147] ,
         \D_cache/cache[3][148] , \D_cache/cache[3][149] ,
         \D_cache/cache[3][150] , \D_cache/cache[3][151] ,
         \D_cache/cache[3][152] , \D_cache/cache[3][153] ,
         \D_cache/cache[3][154] , \D_cache/cache[2][0] , \D_cache/cache[2][1] ,
         \D_cache/cache[2][2] , \D_cache/cache[2][3] , \D_cache/cache[2][4] ,
         \D_cache/cache[2][5] , \D_cache/cache[2][6] , \D_cache/cache[2][7] ,
         \D_cache/cache[2][8] , \D_cache/cache[2][9] , \D_cache/cache[2][10] ,
         \D_cache/cache[2][11] , \D_cache/cache[2][12] ,
         \D_cache/cache[2][13] , \D_cache/cache[2][14] ,
         \D_cache/cache[2][15] , \D_cache/cache[2][16] ,
         \D_cache/cache[2][17] , \D_cache/cache[2][18] ,
         \D_cache/cache[2][19] , \D_cache/cache[2][20] ,
         \D_cache/cache[2][21] , \D_cache/cache[2][22] ,
         \D_cache/cache[2][23] , \D_cache/cache[2][24] ,
         \D_cache/cache[2][25] , \D_cache/cache[2][26] ,
         \D_cache/cache[2][27] , \D_cache/cache[2][28] ,
         \D_cache/cache[2][29] , \D_cache/cache[2][30] ,
         \D_cache/cache[2][31] , \D_cache/cache[2][32] ,
         \D_cache/cache[2][33] , \D_cache/cache[2][34] ,
         \D_cache/cache[2][35] , \D_cache/cache[2][36] ,
         \D_cache/cache[2][37] , \D_cache/cache[2][38] ,
         \D_cache/cache[2][39] , \D_cache/cache[2][40] ,
         \D_cache/cache[2][41] , \D_cache/cache[2][42] ,
         \D_cache/cache[2][43] , \D_cache/cache[2][44] ,
         \D_cache/cache[2][45] , \D_cache/cache[2][46] ,
         \D_cache/cache[2][47] , \D_cache/cache[2][48] ,
         \D_cache/cache[2][49] , \D_cache/cache[2][50] ,
         \D_cache/cache[2][51] , \D_cache/cache[2][52] ,
         \D_cache/cache[2][53] , \D_cache/cache[2][54] ,
         \D_cache/cache[2][55] , \D_cache/cache[2][56] ,
         \D_cache/cache[2][57] , \D_cache/cache[2][58] ,
         \D_cache/cache[2][59] , \D_cache/cache[2][60] ,
         \D_cache/cache[2][61] , \D_cache/cache[2][62] ,
         \D_cache/cache[2][63] , \D_cache/cache[2][64] ,
         \D_cache/cache[2][65] , \D_cache/cache[2][66] ,
         \D_cache/cache[2][67] , \D_cache/cache[2][68] ,
         \D_cache/cache[2][69] , \D_cache/cache[2][70] ,
         \D_cache/cache[2][71] , \D_cache/cache[2][72] ,
         \D_cache/cache[2][73] , \D_cache/cache[2][74] ,
         \D_cache/cache[2][75] , \D_cache/cache[2][76] ,
         \D_cache/cache[2][77] , \D_cache/cache[2][78] ,
         \D_cache/cache[2][79] , \D_cache/cache[2][80] ,
         \D_cache/cache[2][81] , \D_cache/cache[2][82] ,
         \D_cache/cache[2][83] , \D_cache/cache[2][84] ,
         \D_cache/cache[2][85] , \D_cache/cache[2][86] ,
         \D_cache/cache[2][87] , \D_cache/cache[2][88] ,
         \D_cache/cache[2][89] , \D_cache/cache[2][90] ,
         \D_cache/cache[2][91] , \D_cache/cache[2][92] ,
         \D_cache/cache[2][93] , \D_cache/cache[2][94] ,
         \D_cache/cache[2][95] , \D_cache/cache[2][96] ,
         \D_cache/cache[2][97] , \D_cache/cache[2][98] ,
         \D_cache/cache[2][99] , \D_cache/cache[2][100] ,
         \D_cache/cache[2][101] , \D_cache/cache[2][102] ,
         \D_cache/cache[2][103] , \D_cache/cache[2][104] ,
         \D_cache/cache[2][105] , \D_cache/cache[2][106] ,
         \D_cache/cache[2][107] , \D_cache/cache[2][108] ,
         \D_cache/cache[2][109] , \D_cache/cache[2][110] ,
         \D_cache/cache[2][111] , \D_cache/cache[2][112] ,
         \D_cache/cache[2][113] , \D_cache/cache[2][114] ,
         \D_cache/cache[2][115] , \D_cache/cache[2][116] ,
         \D_cache/cache[2][117] , \D_cache/cache[2][118] ,
         \D_cache/cache[2][119] , \D_cache/cache[2][120] ,
         \D_cache/cache[2][121] , \D_cache/cache[2][122] ,
         \D_cache/cache[2][123] , \D_cache/cache[2][124] ,
         \D_cache/cache[2][125] , \D_cache/cache[2][126] ,
         \D_cache/cache[2][127] , \D_cache/cache[2][128] ,
         \D_cache/cache[2][129] , \D_cache/cache[2][130] ,
         \D_cache/cache[2][131] , \D_cache/cache[2][132] ,
         \D_cache/cache[2][133] , \D_cache/cache[2][134] ,
         \D_cache/cache[2][135] , \D_cache/cache[2][136] ,
         \D_cache/cache[2][137] , \D_cache/cache[2][138] ,
         \D_cache/cache[2][139] , \D_cache/cache[2][140] ,
         \D_cache/cache[2][141] , \D_cache/cache[2][142] ,
         \D_cache/cache[2][143] , \D_cache/cache[2][144] ,
         \D_cache/cache[2][145] , \D_cache/cache[2][146] ,
         \D_cache/cache[2][147] , \D_cache/cache[2][148] ,
         \D_cache/cache[2][149] , \D_cache/cache[2][150] ,
         \D_cache/cache[2][151] , \D_cache/cache[2][152] ,
         \D_cache/cache[2][153] , \D_cache/cache[2][154] ,
         \D_cache/cache[1][0] , \D_cache/cache[1][1] , \D_cache/cache[1][2] ,
         \D_cache/cache[1][3] , \D_cache/cache[1][4] , \D_cache/cache[1][5] ,
         \D_cache/cache[1][6] , \D_cache/cache[1][7] , \D_cache/cache[1][8] ,
         \D_cache/cache[1][9] , \D_cache/cache[1][10] , \D_cache/cache[1][11] ,
         \D_cache/cache[1][12] , \D_cache/cache[1][13] ,
         \D_cache/cache[1][14] , \D_cache/cache[1][15] ,
         \D_cache/cache[1][16] , \D_cache/cache[1][17] ,
         \D_cache/cache[1][18] , \D_cache/cache[1][19] ,
         \D_cache/cache[1][20] , \D_cache/cache[1][21] ,
         \D_cache/cache[1][22] , \D_cache/cache[1][23] ,
         \D_cache/cache[1][24] , \D_cache/cache[1][25] ,
         \D_cache/cache[1][26] , \D_cache/cache[1][27] ,
         \D_cache/cache[1][28] , \D_cache/cache[1][29] ,
         \D_cache/cache[1][30] , \D_cache/cache[1][31] ,
         \D_cache/cache[1][32] , \D_cache/cache[1][33] ,
         \D_cache/cache[1][34] , \D_cache/cache[1][35] ,
         \D_cache/cache[1][36] , \D_cache/cache[1][37] ,
         \D_cache/cache[1][38] , \D_cache/cache[1][39] ,
         \D_cache/cache[1][40] , \D_cache/cache[1][41] ,
         \D_cache/cache[1][42] , \D_cache/cache[1][43] ,
         \D_cache/cache[1][44] , \D_cache/cache[1][45] ,
         \D_cache/cache[1][46] , \D_cache/cache[1][47] ,
         \D_cache/cache[1][48] , \D_cache/cache[1][49] ,
         \D_cache/cache[1][50] , \D_cache/cache[1][51] ,
         \D_cache/cache[1][52] , \D_cache/cache[1][53] ,
         \D_cache/cache[1][54] , \D_cache/cache[1][55] ,
         \D_cache/cache[1][56] , \D_cache/cache[1][57] ,
         \D_cache/cache[1][58] , \D_cache/cache[1][59] ,
         \D_cache/cache[1][60] , \D_cache/cache[1][61] ,
         \D_cache/cache[1][62] , \D_cache/cache[1][63] ,
         \D_cache/cache[1][64] , \D_cache/cache[1][65] ,
         \D_cache/cache[1][66] , \D_cache/cache[1][67] ,
         \D_cache/cache[1][68] , \D_cache/cache[1][69] ,
         \D_cache/cache[1][70] , \D_cache/cache[1][71] ,
         \D_cache/cache[1][72] , \D_cache/cache[1][73] ,
         \D_cache/cache[1][74] , \D_cache/cache[1][75] ,
         \D_cache/cache[1][76] , \D_cache/cache[1][77] ,
         \D_cache/cache[1][78] , \D_cache/cache[1][79] ,
         \D_cache/cache[1][80] , \D_cache/cache[1][81] ,
         \D_cache/cache[1][82] , \D_cache/cache[1][83] ,
         \D_cache/cache[1][84] , \D_cache/cache[1][85] ,
         \D_cache/cache[1][86] , \D_cache/cache[1][87] ,
         \D_cache/cache[1][88] , \D_cache/cache[1][89] ,
         \D_cache/cache[1][90] , \D_cache/cache[1][91] ,
         \D_cache/cache[1][92] , \D_cache/cache[1][93] ,
         \D_cache/cache[1][94] , \D_cache/cache[1][95] ,
         \D_cache/cache[1][96] , \D_cache/cache[1][97] ,
         \D_cache/cache[1][98] , \D_cache/cache[1][99] ,
         \D_cache/cache[1][100] , \D_cache/cache[1][101] ,
         \D_cache/cache[1][102] , \D_cache/cache[1][103] ,
         \D_cache/cache[1][104] , \D_cache/cache[1][105] ,
         \D_cache/cache[1][106] , \D_cache/cache[1][107] ,
         \D_cache/cache[1][108] , \D_cache/cache[1][109] ,
         \D_cache/cache[1][110] , \D_cache/cache[1][111] ,
         \D_cache/cache[1][112] , \D_cache/cache[1][113] ,
         \D_cache/cache[1][114] , \D_cache/cache[1][115] ,
         \D_cache/cache[1][116] , \D_cache/cache[1][117] ,
         \D_cache/cache[1][118] , \D_cache/cache[1][119] ,
         \D_cache/cache[1][120] , \D_cache/cache[1][121] ,
         \D_cache/cache[1][122] , \D_cache/cache[1][123] ,
         \D_cache/cache[1][124] , \D_cache/cache[1][125] ,
         \D_cache/cache[1][126] , \D_cache/cache[1][127] ,
         \D_cache/cache[1][128] , \D_cache/cache[1][129] ,
         \D_cache/cache[1][130] , \D_cache/cache[1][131] ,
         \D_cache/cache[1][132] , \D_cache/cache[1][133] ,
         \D_cache/cache[1][134] , \D_cache/cache[1][135] ,
         \D_cache/cache[1][136] , \D_cache/cache[1][137] ,
         \D_cache/cache[1][138] , \D_cache/cache[1][139] ,
         \D_cache/cache[1][140] , \D_cache/cache[1][141] ,
         \D_cache/cache[1][142] , \D_cache/cache[1][143] ,
         \D_cache/cache[1][144] , \D_cache/cache[1][145] ,
         \D_cache/cache[1][146] , \D_cache/cache[1][147] ,
         \D_cache/cache[1][148] , \D_cache/cache[1][149] ,
         \D_cache/cache[1][150] , \D_cache/cache[1][151] ,
         \D_cache/cache[1][152] , \D_cache/cache[1][153] ,
         \D_cache/cache[1][154] , \D_cache/cache[0][0] , \D_cache/cache[0][1] ,
         \D_cache/cache[0][2] , \D_cache/cache[0][3] , \D_cache/cache[0][4] ,
         \D_cache/cache[0][5] , \D_cache/cache[0][6] , \D_cache/cache[0][7] ,
         \D_cache/cache[0][8] , \D_cache/cache[0][9] , \D_cache/cache[0][10] ,
         \D_cache/cache[0][11] , \D_cache/cache[0][12] ,
         \D_cache/cache[0][13] , \D_cache/cache[0][14] ,
         \D_cache/cache[0][15] , \D_cache/cache[0][16] ,
         \D_cache/cache[0][17] , \D_cache/cache[0][18] ,
         \D_cache/cache[0][19] , \D_cache/cache[0][20] ,
         \D_cache/cache[0][21] , \D_cache/cache[0][22] ,
         \D_cache/cache[0][23] , \D_cache/cache[0][24] ,
         \D_cache/cache[0][25] , \D_cache/cache[0][26] ,
         \D_cache/cache[0][27] , \D_cache/cache[0][28] ,
         \D_cache/cache[0][29] , \D_cache/cache[0][30] ,
         \D_cache/cache[0][31] , \D_cache/cache[0][32] ,
         \D_cache/cache[0][33] , \D_cache/cache[0][34] ,
         \D_cache/cache[0][35] , \D_cache/cache[0][36] ,
         \D_cache/cache[0][37] , \D_cache/cache[0][38] ,
         \D_cache/cache[0][39] , \D_cache/cache[0][40] ,
         \D_cache/cache[0][41] , \D_cache/cache[0][42] ,
         \D_cache/cache[0][43] , \D_cache/cache[0][44] ,
         \D_cache/cache[0][45] , \D_cache/cache[0][46] ,
         \D_cache/cache[0][47] , \D_cache/cache[0][48] ,
         \D_cache/cache[0][49] , \D_cache/cache[0][50] ,
         \D_cache/cache[0][51] , \D_cache/cache[0][52] ,
         \D_cache/cache[0][53] , \D_cache/cache[0][54] ,
         \D_cache/cache[0][55] , \D_cache/cache[0][56] ,
         \D_cache/cache[0][57] , \D_cache/cache[0][58] ,
         \D_cache/cache[0][59] , \D_cache/cache[0][60] ,
         \D_cache/cache[0][61] , \D_cache/cache[0][62] ,
         \D_cache/cache[0][63] , \D_cache/cache[0][64] ,
         \D_cache/cache[0][65] , \D_cache/cache[0][66] ,
         \D_cache/cache[0][67] , \D_cache/cache[0][68] ,
         \D_cache/cache[0][69] , \D_cache/cache[0][70] ,
         \D_cache/cache[0][71] , \D_cache/cache[0][72] ,
         \D_cache/cache[0][73] , \D_cache/cache[0][74] ,
         \D_cache/cache[0][75] , \D_cache/cache[0][76] ,
         \D_cache/cache[0][77] , \D_cache/cache[0][78] ,
         \D_cache/cache[0][79] , \D_cache/cache[0][80] ,
         \D_cache/cache[0][81] , \D_cache/cache[0][82] ,
         \D_cache/cache[0][83] , \D_cache/cache[0][84] ,
         \D_cache/cache[0][85] , \D_cache/cache[0][86] ,
         \D_cache/cache[0][87] , \D_cache/cache[0][88] ,
         \D_cache/cache[0][89] , \D_cache/cache[0][90] ,
         \D_cache/cache[0][91] , \D_cache/cache[0][92] ,
         \D_cache/cache[0][93] , \D_cache/cache[0][94] ,
         \D_cache/cache[0][95] , \D_cache/cache[0][96] ,
         \D_cache/cache[0][97] , \D_cache/cache[0][98] ,
         \D_cache/cache[0][99] , \D_cache/cache[0][100] ,
         \D_cache/cache[0][101] , \D_cache/cache[0][102] ,
         \D_cache/cache[0][103] , \D_cache/cache[0][104] ,
         \D_cache/cache[0][105] , \D_cache/cache[0][106] ,
         \D_cache/cache[0][107] , \D_cache/cache[0][108] ,
         \D_cache/cache[0][109] , \D_cache/cache[0][110] ,
         \D_cache/cache[0][111] , \D_cache/cache[0][112] ,
         \D_cache/cache[0][113] , \D_cache/cache[0][114] ,
         \D_cache/cache[0][115] , \D_cache/cache[0][116] ,
         \D_cache/cache[0][117] , \D_cache/cache[0][118] ,
         \D_cache/cache[0][119] , \D_cache/cache[0][120] ,
         \D_cache/cache[0][121] , \D_cache/cache[0][122] ,
         \D_cache/cache[0][123] , \D_cache/cache[0][124] ,
         \D_cache/cache[0][125] , \D_cache/cache[0][126] ,
         \D_cache/cache[0][127] , \D_cache/cache[0][128] ,
         \D_cache/cache[0][129] , \D_cache/cache[0][130] ,
         \D_cache/cache[0][131] , \D_cache/cache[0][132] ,
         \D_cache/cache[0][133] , \D_cache/cache[0][134] ,
         \D_cache/cache[0][135] , \D_cache/cache[0][136] ,
         \D_cache/cache[0][137] , \D_cache/cache[0][138] ,
         \D_cache/cache[0][139] , \D_cache/cache[0][140] ,
         \D_cache/cache[0][141] , \D_cache/cache[0][142] ,
         \D_cache/cache[0][143] , \D_cache/cache[0][144] ,
         \D_cache/cache[0][145] , \D_cache/cache[0][146] ,
         \D_cache/cache[0][147] , \D_cache/cache[0][148] ,
         \D_cache/cache[0][149] , \D_cache/cache[0][150] ,
         \D_cache/cache[0][151] , \D_cache/cache[0][152] ,
         \D_cache/cache[0][153] , \D_cache/cache[0][154] , \i_MIPS/PC/n65 ,
         \i_MIPS/PC/n64 , \i_MIPS/PC/n63 , \i_MIPS/PC/n62 , \i_MIPS/PC/n61 ,
         \i_MIPS/PC/n60 , \i_MIPS/PC/n59 , \i_MIPS/PC/n58 , \i_MIPS/PC/n57 ,
         \i_MIPS/PC/n56 , \i_MIPS/PC/n55 , \i_MIPS/PC/n54 , \i_MIPS/PC/n53 ,
         \i_MIPS/PC/n52 , \i_MIPS/PC/n51 , \i_MIPS/PC/n50 , \i_MIPS/PC/n49 ,
         \i_MIPS/PC/n48 , \i_MIPS/PC/n47 , \i_MIPS/PC/n46 , \i_MIPS/PC/n45 ,
         \i_MIPS/PC/n44 , \i_MIPS/PC/n43 , \i_MIPS/PC/n42 , \i_MIPS/PC/n41 ,
         \i_MIPS/PC/n40 , \i_MIPS/PC/n39 , \i_MIPS/PC/n38 , \i_MIPS/PC/n37 ,
         \i_MIPS/PC/n36 , \i_MIPS/PC/n35 , \i_MIPS/PC/n34 , \i_MIPS/PC/n33 ,
         \i_MIPS/PC/n32 , \i_MIPS/PC/n31 , \i_MIPS/PC/n30 , \i_MIPS/PC/n29 ,
         \i_MIPS/PC/n28 , \i_MIPS/PC/n27 , \i_MIPS/PC/n26 , \i_MIPS/PC/n25 ,
         \i_MIPS/PC/n24 , \i_MIPS/PC/n23 , \i_MIPS/PC/n22 , \i_MIPS/PC/n21 ,
         \i_MIPS/PC/n20 , \i_MIPS/PC/n19 , \i_MIPS/PC/n18 , \i_MIPS/PC/n17 ,
         \i_MIPS/PC/n16 , \i_MIPS/PC/n15 , \i_MIPS/PC/n14 , \i_MIPS/PC/n13 ,
         \i_MIPS/PC/n12 , \i_MIPS/PC/n11 , \i_MIPS/PC/n10 , \i_MIPS/PC/n9 ,
         \i_MIPS/PC/n8 , \i_MIPS/PC/n7 , \i_MIPS/PC/n6 , \i_MIPS/PC/n5 ,
         \i_MIPS/PC/n4 , \i_MIPS/PC/n3 , \i_MIPS/PC/n2 ,
         \i_MIPS/Register/n1139 , \i_MIPS/Register/n1138 ,
         \i_MIPS/Register/n1137 , \i_MIPS/Register/n1136 ,
         \i_MIPS/Register/n1135 , \i_MIPS/Register/n1134 ,
         \i_MIPS/Register/n1133 , \i_MIPS/Register/n1132 ,
         \i_MIPS/Register/n1131 , \i_MIPS/Register/n1130 ,
         \i_MIPS/Register/n1129 , \i_MIPS/Register/n1128 ,
         \i_MIPS/Register/n1127 , \i_MIPS/Register/n1126 ,
         \i_MIPS/Register/n1125 , \i_MIPS/Register/n1124 ,
         \i_MIPS/Register/n1123 , \i_MIPS/Register/n1122 ,
         \i_MIPS/Register/n1121 , \i_MIPS/Register/n1120 ,
         \i_MIPS/Register/n1119 , \i_MIPS/Register/n1118 ,
         \i_MIPS/Register/n1117 , \i_MIPS/Register/n1116 ,
         \i_MIPS/Register/n1115 , \i_MIPS/Register/n1114 ,
         \i_MIPS/Register/n1113 , \i_MIPS/Register/n1112 ,
         \i_MIPS/Register/n1111 , \i_MIPS/Register/n1110 ,
         \i_MIPS/Register/n1109 , \i_MIPS/Register/n1108 ,
         \i_MIPS/Register/n1107 , \i_MIPS/Register/n1106 ,
         \i_MIPS/Register/n1105 , \i_MIPS/Register/n1104 ,
         \i_MIPS/Register/n1103 , \i_MIPS/Register/n1102 ,
         \i_MIPS/Register/n1101 , \i_MIPS/Register/n1100 ,
         \i_MIPS/Register/n1099 , \i_MIPS/Register/n1098 ,
         \i_MIPS/Register/n1097 , \i_MIPS/Register/n1096 ,
         \i_MIPS/Register/n1095 , \i_MIPS/Register/n1094 ,
         \i_MIPS/Register/n1093 , \i_MIPS/Register/n1092 ,
         \i_MIPS/Register/n1091 , \i_MIPS/Register/n1090 ,
         \i_MIPS/Register/n1089 , \i_MIPS/Register/n1088 ,
         \i_MIPS/Register/n1087 , \i_MIPS/Register/n1086 ,
         \i_MIPS/Register/n1085 , \i_MIPS/Register/n1084 ,
         \i_MIPS/Register/n1083 , \i_MIPS/Register/n1082 ,
         \i_MIPS/Register/n1081 , \i_MIPS/Register/n1080 ,
         \i_MIPS/Register/n1079 , \i_MIPS/Register/n1078 ,
         \i_MIPS/Register/n1077 , \i_MIPS/Register/n1076 ,
         \i_MIPS/Register/n1075 , \i_MIPS/Register/n1074 ,
         \i_MIPS/Register/n1073 , \i_MIPS/Register/n1072 ,
         \i_MIPS/Register/n1071 , \i_MIPS/Register/n1070 ,
         \i_MIPS/Register/n1069 , \i_MIPS/Register/n1068 ,
         \i_MIPS/Register/n1067 , \i_MIPS/Register/n1066 ,
         \i_MIPS/Register/n1065 , \i_MIPS/Register/n1064 ,
         \i_MIPS/Register/n1063 , \i_MIPS/Register/n1062 ,
         \i_MIPS/Register/n1061 , \i_MIPS/Register/n1060 ,
         \i_MIPS/Register/n1059 , \i_MIPS/Register/n1058 ,
         \i_MIPS/Register/n1057 , \i_MIPS/Register/n1056 ,
         \i_MIPS/Register/n1055 , \i_MIPS/Register/n1054 ,
         \i_MIPS/Register/n1053 , \i_MIPS/Register/n1052 ,
         \i_MIPS/Register/n1051 , \i_MIPS/Register/n1050 ,
         \i_MIPS/Register/n1049 , \i_MIPS/Register/n1048 ,
         \i_MIPS/Register/n1047 , \i_MIPS/Register/n1046 ,
         \i_MIPS/Register/n1045 , \i_MIPS/Register/n1044 ,
         \i_MIPS/Register/n1043 , \i_MIPS/Register/n1042 ,
         \i_MIPS/Register/n1041 , \i_MIPS/Register/n1040 ,
         \i_MIPS/Register/n1039 , \i_MIPS/Register/n1038 ,
         \i_MIPS/Register/n1037 , \i_MIPS/Register/n1036 ,
         \i_MIPS/Register/n1035 , \i_MIPS/Register/n1034 ,
         \i_MIPS/Register/n1033 , \i_MIPS/Register/n1032 ,
         \i_MIPS/Register/n1031 , \i_MIPS/Register/n1030 ,
         \i_MIPS/Register/n1029 , \i_MIPS/Register/n1028 ,
         \i_MIPS/Register/n1027 , \i_MIPS/Register/n1026 ,
         \i_MIPS/Register/n1025 , \i_MIPS/Register/n1024 ,
         \i_MIPS/Register/n1023 , \i_MIPS/Register/n1022 ,
         \i_MIPS/Register/n1021 , \i_MIPS/Register/n1020 ,
         \i_MIPS/Register/n1019 , \i_MIPS/Register/n1018 ,
         \i_MIPS/Register/n1017 , \i_MIPS/Register/n1016 ,
         \i_MIPS/Register/n1015 , \i_MIPS/Register/n1014 ,
         \i_MIPS/Register/n1013 , \i_MIPS/Register/n1012 ,
         \i_MIPS/Register/n1011 , \i_MIPS/Register/n1010 ,
         \i_MIPS/Register/n1009 , \i_MIPS/Register/n1008 ,
         \i_MIPS/Register/n1007 , \i_MIPS/Register/n1006 ,
         \i_MIPS/Register/n1005 , \i_MIPS/Register/n1004 ,
         \i_MIPS/Register/n1003 , \i_MIPS/Register/n1002 ,
         \i_MIPS/Register/n1001 , \i_MIPS/Register/n1000 ,
         \i_MIPS/Register/n999 , \i_MIPS/Register/n998 ,
         \i_MIPS/Register/n997 , \i_MIPS/Register/n996 ,
         \i_MIPS/Register/n995 , \i_MIPS/Register/n994 ,
         \i_MIPS/Register/n993 , \i_MIPS/Register/n992 ,
         \i_MIPS/Register/n991 , \i_MIPS/Register/n990 ,
         \i_MIPS/Register/n989 , \i_MIPS/Register/n988 ,
         \i_MIPS/Register/n987 , \i_MIPS/Register/n986 ,
         \i_MIPS/Register/n985 , \i_MIPS/Register/n984 ,
         \i_MIPS/Register/n983 , \i_MIPS/Register/n982 ,
         \i_MIPS/Register/n981 , \i_MIPS/Register/n980 ,
         \i_MIPS/Register/n979 , \i_MIPS/Register/n978 ,
         \i_MIPS/Register/n977 , \i_MIPS/Register/n976 ,
         \i_MIPS/Register/n975 , \i_MIPS/Register/n974 ,
         \i_MIPS/Register/n973 , \i_MIPS/Register/n972 ,
         \i_MIPS/Register/n971 , \i_MIPS/Register/n970 ,
         \i_MIPS/Register/n969 , \i_MIPS/Register/n968 ,
         \i_MIPS/Register/n967 , \i_MIPS/Register/n966 ,
         \i_MIPS/Register/n965 , \i_MIPS/Register/n964 ,
         \i_MIPS/Register/n963 , \i_MIPS/Register/n962 ,
         \i_MIPS/Register/n961 , \i_MIPS/Register/n960 ,
         \i_MIPS/Register/n959 , \i_MIPS/Register/n958 ,
         \i_MIPS/Register/n957 , \i_MIPS/Register/n956 ,
         \i_MIPS/Register/n955 , \i_MIPS/Register/n954 ,
         \i_MIPS/Register/n953 , \i_MIPS/Register/n952 ,
         \i_MIPS/Register/n951 , \i_MIPS/Register/n950 ,
         \i_MIPS/Register/n949 , \i_MIPS/Register/n948 ,
         \i_MIPS/Register/n947 , \i_MIPS/Register/n946 ,
         \i_MIPS/Register/n945 , \i_MIPS/Register/n944 ,
         \i_MIPS/Register/n943 , \i_MIPS/Register/n942 ,
         \i_MIPS/Register/n941 , \i_MIPS/Register/n940 ,
         \i_MIPS/Register/n939 , \i_MIPS/Register/n938 ,
         \i_MIPS/Register/n937 , \i_MIPS/Register/n936 ,
         \i_MIPS/Register/n935 , \i_MIPS/Register/n934 ,
         \i_MIPS/Register/n933 , \i_MIPS/Register/n932 ,
         \i_MIPS/Register/n931 , \i_MIPS/Register/n930 ,
         \i_MIPS/Register/n929 , \i_MIPS/Register/n928 ,
         \i_MIPS/Register/n927 , \i_MIPS/Register/n926 ,
         \i_MIPS/Register/n925 , \i_MIPS/Register/n924 ,
         \i_MIPS/Register/n923 , \i_MIPS/Register/n922 ,
         \i_MIPS/Register/n921 , \i_MIPS/Register/n920 ,
         \i_MIPS/Register/n919 , \i_MIPS/Register/n918 ,
         \i_MIPS/Register/n917 , \i_MIPS/Register/n916 ,
         \i_MIPS/Register/n915 , \i_MIPS/Register/n914 ,
         \i_MIPS/Register/n913 , \i_MIPS/Register/n912 ,
         \i_MIPS/Register/n911 , \i_MIPS/Register/n910 ,
         \i_MIPS/Register/n909 , \i_MIPS/Register/n908 ,
         \i_MIPS/Register/n907 , \i_MIPS/Register/n906 ,
         \i_MIPS/Register/n905 , \i_MIPS/Register/n904 ,
         \i_MIPS/Register/n903 , \i_MIPS/Register/n902 ,
         \i_MIPS/Register/n901 , \i_MIPS/Register/n900 ,
         \i_MIPS/Register/n899 , \i_MIPS/Register/n898 ,
         \i_MIPS/Register/n897 , \i_MIPS/Register/n896 ,
         \i_MIPS/Register/n895 , \i_MIPS/Register/n894 ,
         \i_MIPS/Register/n893 , \i_MIPS/Register/n892 ,
         \i_MIPS/Register/n891 , \i_MIPS/Register/n890 ,
         \i_MIPS/Register/n889 , \i_MIPS/Register/n888 ,
         \i_MIPS/Register/n887 , \i_MIPS/Register/n886 ,
         \i_MIPS/Register/n885 , \i_MIPS/Register/n884 ,
         \i_MIPS/Register/n883 , \i_MIPS/Register/n882 ,
         \i_MIPS/Register/n881 , \i_MIPS/Register/n880 ,
         \i_MIPS/Register/n879 , \i_MIPS/Register/n878 ,
         \i_MIPS/Register/n877 , \i_MIPS/Register/n876 ,
         \i_MIPS/Register/n875 , \i_MIPS/Register/n874 ,
         \i_MIPS/Register/n873 , \i_MIPS/Register/n872 ,
         \i_MIPS/Register/n871 , \i_MIPS/Register/n870 ,
         \i_MIPS/Register/n869 , \i_MIPS/Register/n868 ,
         \i_MIPS/Register/n867 , \i_MIPS/Register/n866 ,
         \i_MIPS/Register/n865 , \i_MIPS/Register/n864 ,
         \i_MIPS/Register/n863 , \i_MIPS/Register/n862 ,
         \i_MIPS/Register/n861 , \i_MIPS/Register/n860 ,
         \i_MIPS/Register/n859 , \i_MIPS/Register/n858 ,
         \i_MIPS/Register/n857 , \i_MIPS/Register/n856 ,
         \i_MIPS/Register/n855 , \i_MIPS/Register/n854 ,
         \i_MIPS/Register/n853 , \i_MIPS/Register/n852 ,
         \i_MIPS/Register/n851 , \i_MIPS/Register/n850 ,
         \i_MIPS/Register/n849 , \i_MIPS/Register/n848 ,
         \i_MIPS/Register/n847 , \i_MIPS/Register/n846 ,
         \i_MIPS/Register/n845 , \i_MIPS/Register/n844 ,
         \i_MIPS/Register/n843 , \i_MIPS/Register/n842 ,
         \i_MIPS/Register/n841 , \i_MIPS/Register/n840 ,
         \i_MIPS/Register/n839 , \i_MIPS/Register/n838 ,
         \i_MIPS/Register/n837 , \i_MIPS/Register/n836 ,
         \i_MIPS/Register/n835 , \i_MIPS/Register/n834 ,
         \i_MIPS/Register/n833 , \i_MIPS/Register/n832 ,
         \i_MIPS/Register/n831 , \i_MIPS/Register/n830 ,
         \i_MIPS/Register/n829 , \i_MIPS/Register/n828 ,
         \i_MIPS/Register/n827 , \i_MIPS/Register/n826 ,
         \i_MIPS/Register/n825 , \i_MIPS/Register/n824 ,
         \i_MIPS/Register/n823 , \i_MIPS/Register/n822 ,
         \i_MIPS/Register/n821 , \i_MIPS/Register/n820 ,
         \i_MIPS/Register/n819 , \i_MIPS/Register/n818 ,
         \i_MIPS/Register/n817 , \i_MIPS/Register/n816 ,
         \i_MIPS/Register/n815 , \i_MIPS/Register/n814 ,
         \i_MIPS/Register/n813 , \i_MIPS/Register/n812 ,
         \i_MIPS/Register/n811 , \i_MIPS/Register/n810 ,
         \i_MIPS/Register/n809 , \i_MIPS/Register/n808 ,
         \i_MIPS/Register/n807 , \i_MIPS/Register/n806 ,
         \i_MIPS/Register/n805 , \i_MIPS/Register/n804 ,
         \i_MIPS/Register/n803 , \i_MIPS/Register/n802 ,
         \i_MIPS/Register/n801 , \i_MIPS/Register/n800 ,
         \i_MIPS/Register/n799 , \i_MIPS/Register/n798 ,
         \i_MIPS/Register/n797 , \i_MIPS/Register/n796 ,
         \i_MIPS/Register/n795 , \i_MIPS/Register/n794 ,
         \i_MIPS/Register/n793 , \i_MIPS/Register/n792 ,
         \i_MIPS/Register/n791 , \i_MIPS/Register/n790 ,
         \i_MIPS/Register/n789 , \i_MIPS/Register/n788 ,
         \i_MIPS/Register/n787 , \i_MIPS/Register/n786 ,
         \i_MIPS/Register/n785 , \i_MIPS/Register/n784 ,
         \i_MIPS/Register/n783 , \i_MIPS/Register/n782 ,
         \i_MIPS/Register/n781 , \i_MIPS/Register/n780 ,
         \i_MIPS/Register/n779 , \i_MIPS/Register/n778 ,
         \i_MIPS/Register/n777 , \i_MIPS/Register/n776 ,
         \i_MIPS/Register/n775 , \i_MIPS/Register/n774 ,
         \i_MIPS/Register/n773 , \i_MIPS/Register/n772 ,
         \i_MIPS/Register/n771 , \i_MIPS/Register/n770 ,
         \i_MIPS/Register/n769 , \i_MIPS/Register/n768 ,
         \i_MIPS/Register/n767 , \i_MIPS/Register/n766 ,
         \i_MIPS/Register/n765 , \i_MIPS/Register/n764 ,
         \i_MIPS/Register/n763 , \i_MIPS/Register/n762 ,
         \i_MIPS/Register/n761 , \i_MIPS/Register/n760 ,
         \i_MIPS/Register/n759 , \i_MIPS/Register/n758 ,
         \i_MIPS/Register/n757 , \i_MIPS/Register/n756 ,
         \i_MIPS/Register/n755 , \i_MIPS/Register/n754 ,
         \i_MIPS/Register/n753 , \i_MIPS/Register/n752 ,
         \i_MIPS/Register/n751 , \i_MIPS/Register/n750 ,
         \i_MIPS/Register/n749 , \i_MIPS/Register/n748 ,
         \i_MIPS/Register/n747 , \i_MIPS/Register/n746 ,
         \i_MIPS/Register/n745 , \i_MIPS/Register/n744 ,
         \i_MIPS/Register/n743 , \i_MIPS/Register/n742 ,
         \i_MIPS/Register/n741 , \i_MIPS/Register/n740 ,
         \i_MIPS/Register/n739 , \i_MIPS/Register/n738 ,
         \i_MIPS/Register/n737 , \i_MIPS/Register/n736 ,
         \i_MIPS/Register/n735 , \i_MIPS/Register/n734 ,
         \i_MIPS/Register/n733 , \i_MIPS/Register/n732 ,
         \i_MIPS/Register/n731 , \i_MIPS/Register/n730 ,
         \i_MIPS/Register/n729 , \i_MIPS/Register/n728 ,
         \i_MIPS/Register/n727 , \i_MIPS/Register/n726 ,
         \i_MIPS/Register/n725 , \i_MIPS/Register/n724 ,
         \i_MIPS/Register/n723 , \i_MIPS/Register/n722 ,
         \i_MIPS/Register/n721 , \i_MIPS/Register/n720 ,
         \i_MIPS/Register/n719 , \i_MIPS/Register/n718 ,
         \i_MIPS/Register/n717 , \i_MIPS/Register/n716 ,
         \i_MIPS/Register/n715 , \i_MIPS/Register/n714 ,
         \i_MIPS/Register/n713 , \i_MIPS/Register/n712 ,
         \i_MIPS/Register/n711 , \i_MIPS/Register/n710 ,
         \i_MIPS/Register/n709 , \i_MIPS/Register/n708 ,
         \i_MIPS/Register/n707 , \i_MIPS/Register/n706 ,
         \i_MIPS/Register/n705 , \i_MIPS/Register/n704 ,
         \i_MIPS/Register/n703 , \i_MIPS/Register/n702 ,
         \i_MIPS/Register/n701 , \i_MIPS/Register/n700 ,
         \i_MIPS/Register/n699 , \i_MIPS/Register/n698 ,
         \i_MIPS/Register/n697 , \i_MIPS/Register/n696 ,
         \i_MIPS/Register/n695 , \i_MIPS/Register/n694 ,
         \i_MIPS/Register/n693 , \i_MIPS/Register/n692 ,
         \i_MIPS/Register/n691 , \i_MIPS/Register/n690 ,
         \i_MIPS/Register/n689 , \i_MIPS/Register/n688 ,
         \i_MIPS/Register/n687 , \i_MIPS/Register/n686 ,
         \i_MIPS/Register/n685 , \i_MIPS/Register/n684 ,
         \i_MIPS/Register/n683 , \i_MIPS/Register/n682 ,
         \i_MIPS/Register/n681 , \i_MIPS/Register/n680 ,
         \i_MIPS/Register/n679 , \i_MIPS/Register/n678 ,
         \i_MIPS/Register/n677 , \i_MIPS/Register/n676 ,
         \i_MIPS/Register/n675 , \i_MIPS/Register/n674 ,
         \i_MIPS/Register/n673 , \i_MIPS/Register/n672 ,
         \i_MIPS/Register/n671 , \i_MIPS/Register/n670 ,
         \i_MIPS/Register/n669 , \i_MIPS/Register/n668 ,
         \i_MIPS/Register/n667 , \i_MIPS/Register/n666 ,
         \i_MIPS/Register/n665 , \i_MIPS/Register/n664 ,
         \i_MIPS/Register/n663 , \i_MIPS/Register/n662 ,
         \i_MIPS/Register/n661 , \i_MIPS/Register/n660 ,
         \i_MIPS/Register/n659 , \i_MIPS/Register/n658 ,
         \i_MIPS/Register/n657 , \i_MIPS/Register/n656 ,
         \i_MIPS/Register/n655 , \i_MIPS/Register/n654 ,
         \i_MIPS/Register/n653 , \i_MIPS/Register/n652 ,
         \i_MIPS/Register/n651 , \i_MIPS/Register/n650 ,
         \i_MIPS/Register/n649 , \i_MIPS/Register/n648 ,
         \i_MIPS/Register/n647 , \i_MIPS/Register/n646 ,
         \i_MIPS/Register/n645 , \i_MIPS/Register/n644 ,
         \i_MIPS/Register/n643 , \i_MIPS/Register/n642 ,
         \i_MIPS/Register/n641 , \i_MIPS/Register/n640 ,
         \i_MIPS/Register/n639 , \i_MIPS/Register/n638 ,
         \i_MIPS/Register/n637 , \i_MIPS/Register/n636 ,
         \i_MIPS/Register/n635 , \i_MIPS/Register/n634 ,
         \i_MIPS/Register/n633 , \i_MIPS/Register/n632 ,
         \i_MIPS/Register/n631 , \i_MIPS/Register/n630 ,
         \i_MIPS/Register/n629 , \i_MIPS/Register/n628 ,
         \i_MIPS/Register/n627 , \i_MIPS/Register/n626 ,
         \i_MIPS/Register/n625 , \i_MIPS/Register/n624 ,
         \i_MIPS/Register/n623 , \i_MIPS/Register/n622 ,
         \i_MIPS/Register/n621 , \i_MIPS/Register/n620 ,
         \i_MIPS/Register/n619 , \i_MIPS/Register/n618 ,
         \i_MIPS/Register/n617 , \i_MIPS/Register/n616 ,
         \i_MIPS/Register/n615 , \i_MIPS/Register/n614 ,
         \i_MIPS/Register/n613 , \i_MIPS/Register/n612 ,
         \i_MIPS/Register/n611 , \i_MIPS/Register/n610 ,
         \i_MIPS/Register/n609 , \i_MIPS/Register/n608 ,
         \i_MIPS/Register/n607 , \i_MIPS/Register/n606 ,
         \i_MIPS/Register/n605 , \i_MIPS/Register/n604 ,
         \i_MIPS/Register/n603 , \i_MIPS/Register/n602 ,
         \i_MIPS/Register/n601 , \i_MIPS/Register/n600 ,
         \i_MIPS/Register/n599 , \i_MIPS/Register/n598 ,
         \i_MIPS/Register/n597 , \i_MIPS/Register/n596 ,
         \i_MIPS/Register/n595 , \i_MIPS/Register/n594 ,
         \i_MIPS/Register/n593 , \i_MIPS/Register/n592 ,
         \i_MIPS/Register/n591 , \i_MIPS/Register/n590 ,
         \i_MIPS/Register/n589 , \i_MIPS/Register/n588 ,
         \i_MIPS/Register/n587 , \i_MIPS/Register/n586 ,
         \i_MIPS/Register/n585 , \i_MIPS/Register/n584 ,
         \i_MIPS/Register/n583 , \i_MIPS/Register/n582 ,
         \i_MIPS/Register/n581 , \i_MIPS/Register/n580 ,
         \i_MIPS/Register/n579 , \i_MIPS/Register/n578 ,
         \i_MIPS/Register/n577 , \i_MIPS/Register/n576 ,
         \i_MIPS/Register/n575 , \i_MIPS/Register/n574 ,
         \i_MIPS/Register/n573 , \i_MIPS/Register/n572 ,
         \i_MIPS/Register/n571 , \i_MIPS/Register/n570 ,
         \i_MIPS/Register/n569 , \i_MIPS/Register/n568 ,
         \i_MIPS/Register/n567 , \i_MIPS/Register/n566 ,
         \i_MIPS/Register/n565 , \i_MIPS/Register/n564 ,
         \i_MIPS/Register/n563 , \i_MIPS/Register/n562 ,
         \i_MIPS/Register/n561 , \i_MIPS/Register/n560 ,
         \i_MIPS/Register/n559 , \i_MIPS/Register/n558 ,
         \i_MIPS/Register/n557 , \i_MIPS/Register/n556 ,
         \i_MIPS/Register/n555 , \i_MIPS/Register/n554 ,
         \i_MIPS/Register/n553 , \i_MIPS/Register/n552 ,
         \i_MIPS/Register/n551 , \i_MIPS/Register/n550 ,
         \i_MIPS/Register/n549 , \i_MIPS/Register/n548 ,
         \i_MIPS/Register/n547 , \i_MIPS/Register/n546 ,
         \i_MIPS/Register/n545 , \i_MIPS/Register/n544 ,
         \i_MIPS/Register/n543 , \i_MIPS/Register/n542 ,
         \i_MIPS/Register/n541 , \i_MIPS/Register/n540 ,
         \i_MIPS/Register/n539 , \i_MIPS/Register/n538 ,
         \i_MIPS/Register/n537 , \i_MIPS/Register/n536 ,
         \i_MIPS/Register/n535 , \i_MIPS/Register/n534 ,
         \i_MIPS/Register/n533 , \i_MIPS/Register/n532 ,
         \i_MIPS/Register/n531 , \i_MIPS/Register/n530 ,
         \i_MIPS/Register/n529 , \i_MIPS/Register/n528 ,
         \i_MIPS/Register/n527 , \i_MIPS/Register/n526 ,
         \i_MIPS/Register/n525 , \i_MIPS/Register/n524 ,
         \i_MIPS/Register/n523 , \i_MIPS/Register/n522 ,
         \i_MIPS/Register/n521 , \i_MIPS/Register/n520 ,
         \i_MIPS/Register/n519 , \i_MIPS/Register/n518 ,
         \i_MIPS/Register/n517 , \i_MIPS/Register/n516 ,
         \i_MIPS/Register/n515 , \i_MIPS/Register/n514 ,
         \i_MIPS/Register/n513 , \i_MIPS/Register/n512 ,
         \i_MIPS/Register/n511 , \i_MIPS/Register/n510 ,
         \i_MIPS/Register/n509 , \i_MIPS/Register/n508 ,
         \i_MIPS/Register/n507 , \i_MIPS/Register/n506 ,
         \i_MIPS/Register/n505 , \i_MIPS/Register/n504 ,
         \i_MIPS/Register/n503 , \i_MIPS/Register/n502 ,
         \i_MIPS/Register/n501 , \i_MIPS/Register/n500 ,
         \i_MIPS/Register/n499 , \i_MIPS/Register/n498 ,
         \i_MIPS/Register/n497 , \i_MIPS/Register/n496 ,
         \i_MIPS/Register/n495 , \i_MIPS/Register/n494 ,
         \i_MIPS/Register/n493 , \i_MIPS/Register/n492 ,
         \i_MIPS/Register/n491 , \i_MIPS/Register/n490 ,
         \i_MIPS/Register/n489 , \i_MIPS/Register/n488 ,
         \i_MIPS/Register/n487 , \i_MIPS/Register/n486 ,
         \i_MIPS/Register/n485 , \i_MIPS/Register/n484 ,
         \i_MIPS/Register/n483 , \i_MIPS/Register/n482 ,
         \i_MIPS/Register/n481 , \i_MIPS/Register/n480 ,
         \i_MIPS/Register/n479 , \i_MIPS/Register/n478 ,
         \i_MIPS/Register/n477 , \i_MIPS/Register/n476 ,
         \i_MIPS/Register/n475 , \i_MIPS/Register/n474 ,
         \i_MIPS/Register/n473 , \i_MIPS/Register/n472 ,
         \i_MIPS/Register/n471 , \i_MIPS/Register/n470 ,
         \i_MIPS/Register/n469 , \i_MIPS/Register/n468 ,
         \i_MIPS/Register/n467 , \i_MIPS/Register/n466 ,
         \i_MIPS/Register/n465 , \i_MIPS/Register/n464 ,
         \i_MIPS/Register/n463 , \i_MIPS/Register/n462 ,
         \i_MIPS/Register/n461 , \i_MIPS/Register/n460 ,
         \i_MIPS/Register/n459 , \i_MIPS/Register/n458 ,
         \i_MIPS/Register/n457 , \i_MIPS/Register/n456 ,
         \i_MIPS/Register/n455 , \i_MIPS/Register/n454 ,
         \i_MIPS/Register/n453 , \i_MIPS/Register/n452 ,
         \i_MIPS/Register/n451 , \i_MIPS/Register/n450 ,
         \i_MIPS/Register/n449 , \i_MIPS/Register/n448 ,
         \i_MIPS/Register/n447 , \i_MIPS/Register/n446 ,
         \i_MIPS/Register/n445 , \i_MIPS/Register/n444 ,
         \i_MIPS/Register/n443 , \i_MIPS/Register/n442 ,
         \i_MIPS/Register/n441 , \i_MIPS/Register/n440 ,
         \i_MIPS/Register/n439 , \i_MIPS/Register/n438 ,
         \i_MIPS/Register/n437 , \i_MIPS/Register/n436 ,
         \i_MIPS/Register/n435 , \i_MIPS/Register/n434 ,
         \i_MIPS/Register/n433 , \i_MIPS/Register/n432 ,
         \i_MIPS/Register/n431 , \i_MIPS/Register/n430 ,
         \i_MIPS/Register/n429 , \i_MIPS/Register/n428 ,
         \i_MIPS/Register/n427 , \i_MIPS/Register/n426 ,
         \i_MIPS/Register/n425 , \i_MIPS/Register/n424 ,
         \i_MIPS/Register/n423 , \i_MIPS/Register/n422 ,
         \i_MIPS/Register/n421 , \i_MIPS/Register/n420 ,
         \i_MIPS/Register/n419 , \i_MIPS/Register/n418 ,
         \i_MIPS/Register/n417 , \i_MIPS/Register/n416 ,
         \i_MIPS/Register/n415 , \i_MIPS/Register/n414 ,
         \i_MIPS/Register/n413 , \i_MIPS/Register/n412 ,
         \i_MIPS/Register/n411 , \i_MIPS/Register/n410 ,
         \i_MIPS/Register/n409 , \i_MIPS/Register/n408 ,
         \i_MIPS/Register/n407 , \i_MIPS/Register/n406 ,
         \i_MIPS/Register/n405 , \i_MIPS/Register/n404 ,
         \i_MIPS/Register/n403 , \i_MIPS/Register/n402 ,
         \i_MIPS/Register/n401 , \i_MIPS/Register/n400 ,
         \i_MIPS/Register/n399 , \i_MIPS/Register/n398 ,
         \i_MIPS/Register/n397 , \i_MIPS/Register/n396 ,
         \i_MIPS/Register/n395 , \i_MIPS/Register/n394 ,
         \i_MIPS/Register/n393 , \i_MIPS/Register/n392 ,
         \i_MIPS/Register/n391 , \i_MIPS/Register/n390 ,
         \i_MIPS/Register/n389 , \i_MIPS/Register/n388 ,
         \i_MIPS/Register/n387 , \i_MIPS/Register/n386 ,
         \i_MIPS/Register/n385 , \i_MIPS/Register/n384 ,
         \i_MIPS/Register/n383 , \i_MIPS/Register/n382 ,
         \i_MIPS/Register/n381 , \i_MIPS/Register/n380 ,
         \i_MIPS/Register/n379 , \i_MIPS/Register/n378 ,
         \i_MIPS/Register/n377 , \i_MIPS/Register/n376 ,
         \i_MIPS/Register/n375 , \i_MIPS/Register/n374 ,
         \i_MIPS/Register/n373 , \i_MIPS/Register/n372 ,
         \i_MIPS/Register/n371 , \i_MIPS/Register/n370 ,
         \i_MIPS/Register/n369 , \i_MIPS/Register/n368 ,
         \i_MIPS/Register/n367 , \i_MIPS/Register/n366 ,
         \i_MIPS/Register/n365 , \i_MIPS/Register/n364 ,
         \i_MIPS/Register/n363 , \i_MIPS/Register/n362 ,
         \i_MIPS/Register/n361 , \i_MIPS/Register/n360 ,
         \i_MIPS/Register/n359 , \i_MIPS/Register/n358 ,
         \i_MIPS/Register/n357 , \i_MIPS/Register/n356 ,
         \i_MIPS/Register/n355 , \i_MIPS/Register/n354 ,
         \i_MIPS/Register/n353 , \i_MIPS/Register/n352 ,
         \i_MIPS/Register/n351 , \i_MIPS/Register/n350 ,
         \i_MIPS/Register/n349 , \i_MIPS/Register/n348 ,
         \i_MIPS/Register/n347 , \i_MIPS/Register/n346 ,
         \i_MIPS/Register/n345 , \i_MIPS/Register/n344 ,
         \i_MIPS/Register/n343 , \i_MIPS/Register/n342 ,
         \i_MIPS/Register/n341 , \i_MIPS/Register/n340 ,
         \i_MIPS/Register/n339 , \i_MIPS/Register/n338 ,
         \i_MIPS/Register/n337 , \i_MIPS/Register/n336 ,
         \i_MIPS/Register/n335 , \i_MIPS/Register/n334 ,
         \i_MIPS/Register/n333 , \i_MIPS/Register/n332 ,
         \i_MIPS/Register/n331 , \i_MIPS/Register/n330 ,
         \i_MIPS/Register/n329 , \i_MIPS/Register/n328 ,
         \i_MIPS/Register/n327 , \i_MIPS/Register/n326 ,
         \i_MIPS/Register/n325 , \i_MIPS/Register/n324 ,
         \i_MIPS/Register/n323 , \i_MIPS/Register/n322 ,
         \i_MIPS/Register/n321 , \i_MIPS/Register/n320 ,
         \i_MIPS/Register/n319 , \i_MIPS/Register/n318 ,
         \i_MIPS/Register/n317 , \i_MIPS/Register/n316 ,
         \i_MIPS/Register/n315 , \i_MIPS/Register/n314 ,
         \i_MIPS/Register/n313 , \i_MIPS/Register/n312 ,
         \i_MIPS/Register/n311 , \i_MIPS/Register/n310 ,
         \i_MIPS/Register/n309 , \i_MIPS/Register/n308 ,
         \i_MIPS/Register/n307 , \i_MIPS/Register/n306 ,
         \i_MIPS/Register/n305 , \i_MIPS/Register/n304 ,
         \i_MIPS/Register/n303 , \i_MIPS/Register/n302 ,
         \i_MIPS/Register/n301 , \i_MIPS/Register/n300 ,
         \i_MIPS/Register/n299 , \i_MIPS/Register/n298 ,
         \i_MIPS/Register/n297 , \i_MIPS/Register/n296 ,
         \i_MIPS/Register/n295 , \i_MIPS/Register/n294 ,
         \i_MIPS/Register/n293 , \i_MIPS/Register/n292 ,
         \i_MIPS/Register/n291 , \i_MIPS/Register/n290 ,
         \i_MIPS/Register/n289 , \i_MIPS/Register/n288 ,
         \i_MIPS/Register/n287 , \i_MIPS/Register/n286 ,
         \i_MIPS/Register/n285 , \i_MIPS/Register/n284 ,
         \i_MIPS/Register/n283 , \i_MIPS/Register/n282 ,
         \i_MIPS/Register/n281 , \i_MIPS/Register/n280 ,
         \i_MIPS/Register/n279 , \i_MIPS/Register/n278 ,
         \i_MIPS/Register/n277 , \i_MIPS/Register/n276 ,
         \i_MIPS/Register/n275 , \i_MIPS/Register/n274 ,
         \i_MIPS/Register/n273 , \i_MIPS/Register/n272 ,
         \i_MIPS/Register/n271 , \i_MIPS/Register/n270 ,
         \i_MIPS/Register/n269 , \i_MIPS/Register/n268 ,
         \i_MIPS/Register/n267 , \i_MIPS/Register/n266 ,
         \i_MIPS/Register/n265 , \i_MIPS/Register/n264 ,
         \i_MIPS/Register/n263 , \i_MIPS/Register/n262 ,
         \i_MIPS/Register/n261 , \i_MIPS/Register/n260 ,
         \i_MIPS/Register/n259 , \i_MIPS/Register/n258 ,
         \i_MIPS/Register/n257 , \i_MIPS/Register/n256 ,
         \i_MIPS/Register/n255 , \i_MIPS/Register/n254 ,
         \i_MIPS/Register/n253 , \i_MIPS/Register/n252 ,
         \i_MIPS/Register/n251 , \i_MIPS/Register/n250 ,
         \i_MIPS/Register/n249 , \i_MIPS/Register/n248 ,
         \i_MIPS/Register/n247 , \i_MIPS/Register/n246 ,
         \i_MIPS/Register/n245 , \i_MIPS/Register/n244 ,
         \i_MIPS/Register/n243 , \i_MIPS/Register/n242 ,
         \i_MIPS/Register/n241 , \i_MIPS/Register/n240 ,
         \i_MIPS/Register/n239 , \i_MIPS/Register/n238 ,
         \i_MIPS/Register/n237 , \i_MIPS/Register/n236 ,
         \i_MIPS/Register/n235 , \i_MIPS/Register/n234 ,
         \i_MIPS/Register/n233 , \i_MIPS/Register/n232 ,
         \i_MIPS/Register/n231 , \i_MIPS/Register/n230 ,
         \i_MIPS/Register/n229 , \i_MIPS/Register/n228 ,
         \i_MIPS/Register/n227 , \i_MIPS/Register/n226 ,
         \i_MIPS/Register/n225 , \i_MIPS/Register/n224 ,
         \i_MIPS/Register/n223 , \i_MIPS/Register/n222 ,
         \i_MIPS/Register/n221 , \i_MIPS/Register/n220 ,
         \i_MIPS/Register/n219 , \i_MIPS/Register/n218 ,
         \i_MIPS/Register/n217 , \i_MIPS/Register/n216 ,
         \i_MIPS/Register/n215 , \i_MIPS/Register/n214 ,
         \i_MIPS/Register/n213 , \i_MIPS/Register/n212 ,
         \i_MIPS/Register/n211 , \i_MIPS/Register/n210 ,
         \i_MIPS/Register/n209 , \i_MIPS/Register/n208 ,
         \i_MIPS/Register/n207 , \i_MIPS/Register/n206 ,
         \i_MIPS/Register/n205 , \i_MIPS/Register/n204 ,
         \i_MIPS/Register/n203 , \i_MIPS/Register/n202 ,
         \i_MIPS/Register/n201 , \i_MIPS/Register/n200 ,
         \i_MIPS/Register/n199 , \i_MIPS/Register/n198 ,
         \i_MIPS/Register/n197 , \i_MIPS/Register/n196 ,
         \i_MIPS/Register/n195 , \i_MIPS/Register/n194 ,
         \i_MIPS/Register/n193 , \i_MIPS/Register/n192 ,
         \i_MIPS/Register/n191 , \i_MIPS/Register/n190 ,
         \i_MIPS/Register/n189 , \i_MIPS/Register/n188 ,
         \i_MIPS/Register/n187 , \i_MIPS/Register/n186 ,
         \i_MIPS/Register/n185 , \i_MIPS/Register/n184 ,
         \i_MIPS/Register/n183 , \i_MIPS/Register/n182 ,
         \i_MIPS/Register/n181 , \i_MIPS/Register/n180 ,
         \i_MIPS/Register/n179 , \i_MIPS/Register/n178 ,
         \i_MIPS/Register/n177 , \i_MIPS/Register/n176 ,
         \i_MIPS/Register/n175 , \i_MIPS/Register/n174 ,
         \i_MIPS/Register/n173 , \i_MIPS/Register/n172 ,
         \i_MIPS/Register/n171 , \i_MIPS/Register/n170 ,
         \i_MIPS/Register/n169 , \i_MIPS/Register/n168 ,
         \i_MIPS/Register/n167 , \i_MIPS/Register/n166 ,
         \i_MIPS/Register/n165 , \i_MIPS/Register/n164 ,
         \i_MIPS/Register/n163 , \i_MIPS/Register/n162 ,
         \i_MIPS/Register/n161 , \i_MIPS/Register/n160 ,
         \i_MIPS/Register/n159 , \i_MIPS/Register/n158 ,
         \i_MIPS/Register/n157 , \i_MIPS/Register/n156 ,
         \i_MIPS/Register/n155 , \i_MIPS/Register/n154 ,
         \i_MIPS/Register/n153 , \i_MIPS/Register/n152 ,
         \i_MIPS/Register/n151 , \i_MIPS/Register/n150 ,
         \i_MIPS/Register/n149 , \i_MIPS/Register/n148 ,
         \i_MIPS/Register/n147 , \i_MIPS/Register/n146 ,
         \i_MIPS/Register/n145 , \i_MIPS/Register/n144 ,
         \i_MIPS/Register/n143 , \i_MIPS/Register/n142 ,
         \i_MIPS/Register/n141 , \i_MIPS/Register/n140 ,
         \i_MIPS/Register/n139 , \i_MIPS/Register/n138 ,
         \i_MIPS/Register/n137 , \i_MIPS/Register/n136 ,
         \i_MIPS/Register/n135 , \i_MIPS/Register/n134 ,
         \i_MIPS/Register/n133 , \i_MIPS/Register/n132 ,
         \i_MIPS/Register/n131 , \i_MIPS/Register/n130 ,
         \i_MIPS/Register/n129 , \i_MIPS/Register/n128 ,
         \i_MIPS/Register/n127 , \i_MIPS/Register/n126 ,
         \i_MIPS/Register/n125 , \i_MIPS/Register/n124 ,
         \i_MIPS/Register/n123 , \i_MIPS/Register/n122 ,
         \i_MIPS/Register/n121 , \i_MIPS/Register/n120 ,
         \i_MIPS/Register/n119 , \i_MIPS/Register/n118 ,
         \i_MIPS/Register/n117 , \i_MIPS/Register/n116 ,
         \i_MIPS/Register/n115 , \i_MIPS/Register/n114 ,
         \i_MIPS/Register/n113 , \i_MIPS/Register/n112 ,
         \i_MIPS/Register/n111 , \i_MIPS/Register/n110 ,
         \i_MIPS/Register/n109 , \i_MIPS/Register/n108 ,
         \i_MIPS/Register/n107 , \i_MIPS/Register/n106 ,
         \i_MIPS/Register/n105 , \i_MIPS/Register/n104 ,
         \i_MIPS/Register/register[31][0] , \i_MIPS/Register/register[31][1] ,
         \i_MIPS/Register/register[31][2] , \i_MIPS/Register/register[31][3] ,
         \i_MIPS/Register/register[31][4] , \i_MIPS/Register/register[31][5] ,
         \i_MIPS/Register/register[31][6] , \i_MIPS/Register/register[31][7] ,
         \i_MIPS/Register/register[31][8] , \i_MIPS/Register/register[31][9] ,
         \i_MIPS/Register/register[31][10] ,
         \i_MIPS/Register/register[31][11] ,
         \i_MIPS/Register/register[31][12] ,
         \i_MIPS/Register/register[31][13] ,
         \i_MIPS/Register/register[31][15] ,
         \i_MIPS/Register/register[31][16] ,
         \i_MIPS/Register/register[31][17] ,
         \i_MIPS/Register/register[31][18] ,
         \i_MIPS/Register/register[31][19] ,
         \i_MIPS/Register/register[31][20] ,
         \i_MIPS/Register/register[31][21] ,
         \i_MIPS/Register/register[31][22] ,
         \i_MIPS/Register/register[31][23] ,
         \i_MIPS/Register/register[31][24] ,
         \i_MIPS/Register/register[31][25] ,
         \i_MIPS/Register/register[31][26] ,
         \i_MIPS/Register/register[31][27] ,
         \i_MIPS/Register/register[31][28] ,
         \i_MIPS/Register/register[31][29] , \i_MIPS/Register/register[30][0] ,
         \i_MIPS/Register/register[30][1] , \i_MIPS/Register/register[30][2] ,
         \i_MIPS/Register/register[30][3] , \i_MIPS/Register/register[30][4] ,
         \i_MIPS/Register/register[30][5] , \i_MIPS/Register/register[30][6] ,
         \i_MIPS/Register/register[30][7] , \i_MIPS/Register/register[30][8] ,
         \i_MIPS/Register/register[30][9] , \i_MIPS/Register/register[30][10] ,
         \i_MIPS/Register/register[30][11] ,
         \i_MIPS/Register/register[30][12] ,
         \i_MIPS/Register/register[30][13] ,
         \i_MIPS/Register/register[30][14] ,
         \i_MIPS/Register/register[30][15] ,
         \i_MIPS/Register/register[30][16] ,
         \i_MIPS/Register/register[30][17] ,
         \i_MIPS/Register/register[30][18] ,
         \i_MIPS/Register/register[30][19] ,
         \i_MIPS/Register/register[30][20] ,
         \i_MIPS/Register/register[30][21] ,
         \i_MIPS/Register/register[30][22] ,
         \i_MIPS/Register/register[30][23] ,
         \i_MIPS/Register/register[30][24] ,
         \i_MIPS/Register/register[30][25] ,
         \i_MIPS/Register/register[30][26] ,
         \i_MIPS/Register/register[30][27] ,
         \i_MIPS/Register/register[30][28] ,
         \i_MIPS/Register/register[30][29] ,
         \i_MIPS/Register/register[30][30] ,
         \i_MIPS/Register/register[30][31] , \i_MIPS/Register/register[29][0] ,
         \i_MIPS/Register/register[29][1] , \i_MIPS/Register/register[29][2] ,
         \i_MIPS/Register/register[29][3] , \i_MIPS/Register/register[29][4] ,
         \i_MIPS/Register/register[29][5] , \i_MIPS/Register/register[29][6] ,
         \i_MIPS/Register/register[29][7] , \i_MIPS/Register/register[29][8] ,
         \i_MIPS/Register/register[29][9] , \i_MIPS/Register/register[29][10] ,
         \i_MIPS/Register/register[29][11] ,
         \i_MIPS/Register/register[29][12] ,
         \i_MIPS/Register/register[29][13] ,
         \i_MIPS/Register/register[29][14] ,
         \i_MIPS/Register/register[29][15] ,
         \i_MIPS/Register/register[29][16] ,
         \i_MIPS/Register/register[29][17] ,
         \i_MIPS/Register/register[29][18] ,
         \i_MIPS/Register/register[29][19] ,
         \i_MIPS/Register/register[29][20] ,
         \i_MIPS/Register/register[29][21] ,
         \i_MIPS/Register/register[29][22] ,
         \i_MIPS/Register/register[29][23] ,
         \i_MIPS/Register/register[29][24] ,
         \i_MIPS/Register/register[29][25] ,
         \i_MIPS/Register/register[29][26] ,
         \i_MIPS/Register/register[29][27] ,
         \i_MIPS/Register/register[29][28] ,
         \i_MIPS/Register/register[29][29] ,
         \i_MIPS/Register/register[29][30] ,
         \i_MIPS/Register/register[29][31] , \i_MIPS/Register/register[28][0] ,
         \i_MIPS/Register/register[28][1] , \i_MIPS/Register/register[28][2] ,
         \i_MIPS/Register/register[28][3] , \i_MIPS/Register/register[28][4] ,
         \i_MIPS/Register/register[28][5] , \i_MIPS/Register/register[28][6] ,
         \i_MIPS/Register/register[28][7] , \i_MIPS/Register/register[28][8] ,
         \i_MIPS/Register/register[28][9] , \i_MIPS/Register/register[28][10] ,
         \i_MIPS/Register/register[28][11] ,
         \i_MIPS/Register/register[28][12] ,
         \i_MIPS/Register/register[28][13] ,
         \i_MIPS/Register/register[28][14] ,
         \i_MIPS/Register/register[28][15] ,
         \i_MIPS/Register/register[28][16] ,
         \i_MIPS/Register/register[28][17] ,
         \i_MIPS/Register/register[28][18] ,
         \i_MIPS/Register/register[28][19] ,
         \i_MIPS/Register/register[28][20] ,
         \i_MIPS/Register/register[28][21] ,
         \i_MIPS/Register/register[28][22] ,
         \i_MIPS/Register/register[28][23] ,
         \i_MIPS/Register/register[28][24] ,
         \i_MIPS/Register/register[28][25] ,
         \i_MIPS/Register/register[28][26] ,
         \i_MIPS/Register/register[28][27] ,
         \i_MIPS/Register/register[28][28] ,
         \i_MIPS/Register/register[28][29] ,
         \i_MIPS/Register/register[28][30] ,
         \i_MIPS/Register/register[28][31] , \i_MIPS/Register/register[27][0] ,
         \i_MIPS/Register/register[27][1] , \i_MIPS/Register/register[27][2] ,
         \i_MIPS/Register/register[27][3] , \i_MIPS/Register/register[27][4] ,
         \i_MIPS/Register/register[27][5] , \i_MIPS/Register/register[27][6] ,
         \i_MIPS/Register/register[27][7] , \i_MIPS/Register/register[27][8] ,
         \i_MIPS/Register/register[27][9] , \i_MIPS/Register/register[27][10] ,
         \i_MIPS/Register/register[27][11] ,
         \i_MIPS/Register/register[27][12] ,
         \i_MIPS/Register/register[27][13] ,
         \i_MIPS/Register/register[27][14] ,
         \i_MIPS/Register/register[27][15] ,
         \i_MIPS/Register/register[27][16] ,
         \i_MIPS/Register/register[27][17] ,
         \i_MIPS/Register/register[27][18] ,
         \i_MIPS/Register/register[27][19] ,
         \i_MIPS/Register/register[27][20] ,
         \i_MIPS/Register/register[27][21] ,
         \i_MIPS/Register/register[27][22] ,
         \i_MIPS/Register/register[27][23] ,
         \i_MIPS/Register/register[27][24] ,
         \i_MIPS/Register/register[27][25] ,
         \i_MIPS/Register/register[27][26] ,
         \i_MIPS/Register/register[27][27] ,
         \i_MIPS/Register/register[27][28] ,
         \i_MIPS/Register/register[27][29] ,
         \i_MIPS/Register/register[27][30] ,
         \i_MIPS/Register/register[27][31] , \i_MIPS/Register/register[26][0] ,
         \i_MIPS/Register/register[26][1] , \i_MIPS/Register/register[26][2] ,
         \i_MIPS/Register/register[26][3] , \i_MIPS/Register/register[26][4] ,
         \i_MIPS/Register/register[26][5] , \i_MIPS/Register/register[26][6] ,
         \i_MIPS/Register/register[26][7] , \i_MIPS/Register/register[26][8] ,
         \i_MIPS/Register/register[26][9] , \i_MIPS/Register/register[26][10] ,
         \i_MIPS/Register/register[26][11] ,
         \i_MIPS/Register/register[26][12] ,
         \i_MIPS/Register/register[26][13] ,
         \i_MIPS/Register/register[26][14] ,
         \i_MIPS/Register/register[26][15] ,
         \i_MIPS/Register/register[26][16] ,
         \i_MIPS/Register/register[26][17] ,
         \i_MIPS/Register/register[26][18] ,
         \i_MIPS/Register/register[26][19] ,
         \i_MIPS/Register/register[26][20] ,
         \i_MIPS/Register/register[26][21] ,
         \i_MIPS/Register/register[26][22] ,
         \i_MIPS/Register/register[26][23] ,
         \i_MIPS/Register/register[26][24] ,
         \i_MIPS/Register/register[26][25] ,
         \i_MIPS/Register/register[26][26] ,
         \i_MIPS/Register/register[26][27] ,
         \i_MIPS/Register/register[26][28] ,
         \i_MIPS/Register/register[26][29] ,
         \i_MIPS/Register/register[26][30] ,
         \i_MIPS/Register/register[26][31] , \i_MIPS/Register/register[25][0] ,
         \i_MIPS/Register/register[25][1] , \i_MIPS/Register/register[25][2] ,
         \i_MIPS/Register/register[25][3] , \i_MIPS/Register/register[25][4] ,
         \i_MIPS/Register/register[25][5] , \i_MIPS/Register/register[25][6] ,
         \i_MIPS/Register/register[25][7] , \i_MIPS/Register/register[25][8] ,
         \i_MIPS/Register/register[25][9] , \i_MIPS/Register/register[25][10] ,
         \i_MIPS/Register/register[25][11] ,
         \i_MIPS/Register/register[25][12] ,
         \i_MIPS/Register/register[25][13] ,
         \i_MIPS/Register/register[25][14] ,
         \i_MIPS/Register/register[25][15] ,
         \i_MIPS/Register/register[25][16] ,
         \i_MIPS/Register/register[25][17] ,
         \i_MIPS/Register/register[25][18] ,
         \i_MIPS/Register/register[25][19] ,
         \i_MIPS/Register/register[25][20] ,
         \i_MIPS/Register/register[25][21] ,
         \i_MIPS/Register/register[25][22] ,
         \i_MIPS/Register/register[25][23] ,
         \i_MIPS/Register/register[25][24] ,
         \i_MIPS/Register/register[25][25] ,
         \i_MIPS/Register/register[25][26] ,
         \i_MIPS/Register/register[25][27] ,
         \i_MIPS/Register/register[25][28] ,
         \i_MIPS/Register/register[25][29] ,
         \i_MIPS/Register/register[25][30] ,
         \i_MIPS/Register/register[25][31] , \i_MIPS/Register/register[24][0] ,
         \i_MIPS/Register/register[24][1] , \i_MIPS/Register/register[24][2] ,
         \i_MIPS/Register/register[24][3] , \i_MIPS/Register/register[24][4] ,
         \i_MIPS/Register/register[24][5] , \i_MIPS/Register/register[24][6] ,
         \i_MIPS/Register/register[24][7] , \i_MIPS/Register/register[24][8] ,
         \i_MIPS/Register/register[24][9] , \i_MIPS/Register/register[24][10] ,
         \i_MIPS/Register/register[24][11] ,
         \i_MIPS/Register/register[24][12] ,
         \i_MIPS/Register/register[24][13] ,
         \i_MIPS/Register/register[24][14] ,
         \i_MIPS/Register/register[24][15] ,
         \i_MIPS/Register/register[24][16] ,
         \i_MIPS/Register/register[24][17] ,
         \i_MIPS/Register/register[24][18] ,
         \i_MIPS/Register/register[24][19] ,
         \i_MIPS/Register/register[24][20] ,
         \i_MIPS/Register/register[24][21] ,
         \i_MIPS/Register/register[24][22] ,
         \i_MIPS/Register/register[24][23] ,
         \i_MIPS/Register/register[24][24] ,
         \i_MIPS/Register/register[24][25] ,
         \i_MIPS/Register/register[24][26] ,
         \i_MIPS/Register/register[24][27] ,
         \i_MIPS/Register/register[24][28] ,
         \i_MIPS/Register/register[24][29] ,
         \i_MIPS/Register/register[24][30] ,
         \i_MIPS/Register/register[24][31] , \i_MIPS/Register/register[23][0] ,
         \i_MIPS/Register/register[23][1] , \i_MIPS/Register/register[23][2] ,
         \i_MIPS/Register/register[23][3] , \i_MIPS/Register/register[23][4] ,
         \i_MIPS/Register/register[23][5] , \i_MIPS/Register/register[23][6] ,
         \i_MIPS/Register/register[23][7] , \i_MIPS/Register/register[23][8] ,
         \i_MIPS/Register/register[23][9] , \i_MIPS/Register/register[23][10] ,
         \i_MIPS/Register/register[23][11] ,
         \i_MIPS/Register/register[23][12] ,
         \i_MIPS/Register/register[23][13] ,
         \i_MIPS/Register/register[23][14] ,
         \i_MIPS/Register/register[23][15] ,
         \i_MIPS/Register/register[23][16] ,
         \i_MIPS/Register/register[23][17] ,
         \i_MIPS/Register/register[23][18] ,
         \i_MIPS/Register/register[23][19] ,
         \i_MIPS/Register/register[23][20] ,
         \i_MIPS/Register/register[23][21] ,
         \i_MIPS/Register/register[23][22] ,
         \i_MIPS/Register/register[23][23] ,
         \i_MIPS/Register/register[23][24] ,
         \i_MIPS/Register/register[23][25] ,
         \i_MIPS/Register/register[23][26] ,
         \i_MIPS/Register/register[23][27] ,
         \i_MIPS/Register/register[23][28] ,
         \i_MIPS/Register/register[23][29] ,
         \i_MIPS/Register/register[23][30] ,
         \i_MIPS/Register/register[23][31] , \i_MIPS/Register/register[22][0] ,
         \i_MIPS/Register/register[22][1] , \i_MIPS/Register/register[22][2] ,
         \i_MIPS/Register/register[22][3] , \i_MIPS/Register/register[22][4] ,
         \i_MIPS/Register/register[22][5] , \i_MIPS/Register/register[22][6] ,
         \i_MIPS/Register/register[22][7] , \i_MIPS/Register/register[22][8] ,
         \i_MIPS/Register/register[22][9] , \i_MIPS/Register/register[22][10] ,
         \i_MIPS/Register/register[22][11] ,
         \i_MIPS/Register/register[22][12] ,
         \i_MIPS/Register/register[22][13] ,
         \i_MIPS/Register/register[22][14] ,
         \i_MIPS/Register/register[22][15] ,
         \i_MIPS/Register/register[22][16] ,
         \i_MIPS/Register/register[22][17] ,
         \i_MIPS/Register/register[22][18] ,
         \i_MIPS/Register/register[22][19] ,
         \i_MIPS/Register/register[22][20] ,
         \i_MIPS/Register/register[22][21] ,
         \i_MIPS/Register/register[22][22] ,
         \i_MIPS/Register/register[22][23] ,
         \i_MIPS/Register/register[22][24] ,
         \i_MIPS/Register/register[22][25] ,
         \i_MIPS/Register/register[22][26] ,
         \i_MIPS/Register/register[22][27] ,
         \i_MIPS/Register/register[22][28] ,
         \i_MIPS/Register/register[22][29] ,
         \i_MIPS/Register/register[22][30] ,
         \i_MIPS/Register/register[22][31] , \i_MIPS/Register/register[21][0] ,
         \i_MIPS/Register/register[21][1] , \i_MIPS/Register/register[21][2] ,
         \i_MIPS/Register/register[21][3] , \i_MIPS/Register/register[21][4] ,
         \i_MIPS/Register/register[21][5] , \i_MIPS/Register/register[21][6] ,
         \i_MIPS/Register/register[21][7] , \i_MIPS/Register/register[21][8] ,
         \i_MIPS/Register/register[21][9] , \i_MIPS/Register/register[21][10] ,
         \i_MIPS/Register/register[21][11] ,
         \i_MIPS/Register/register[21][12] ,
         \i_MIPS/Register/register[21][13] ,
         \i_MIPS/Register/register[21][14] ,
         \i_MIPS/Register/register[21][15] ,
         \i_MIPS/Register/register[21][16] ,
         \i_MIPS/Register/register[21][17] ,
         \i_MIPS/Register/register[21][18] ,
         \i_MIPS/Register/register[21][19] ,
         \i_MIPS/Register/register[21][20] ,
         \i_MIPS/Register/register[21][21] ,
         \i_MIPS/Register/register[21][22] ,
         \i_MIPS/Register/register[21][23] ,
         \i_MIPS/Register/register[21][24] ,
         \i_MIPS/Register/register[21][25] ,
         \i_MIPS/Register/register[21][26] ,
         \i_MIPS/Register/register[21][27] ,
         \i_MIPS/Register/register[21][28] ,
         \i_MIPS/Register/register[21][29] ,
         \i_MIPS/Register/register[21][30] ,
         \i_MIPS/Register/register[21][31] , \i_MIPS/Register/register[20][0] ,
         \i_MIPS/Register/register[20][1] , \i_MIPS/Register/register[20][2] ,
         \i_MIPS/Register/register[20][3] , \i_MIPS/Register/register[20][4] ,
         \i_MIPS/Register/register[20][5] , \i_MIPS/Register/register[20][6] ,
         \i_MIPS/Register/register[20][7] , \i_MIPS/Register/register[20][8] ,
         \i_MIPS/Register/register[20][9] , \i_MIPS/Register/register[20][10] ,
         \i_MIPS/Register/register[20][11] ,
         \i_MIPS/Register/register[20][12] ,
         \i_MIPS/Register/register[20][13] ,
         \i_MIPS/Register/register[20][14] ,
         \i_MIPS/Register/register[20][15] ,
         \i_MIPS/Register/register[20][16] ,
         \i_MIPS/Register/register[20][17] ,
         \i_MIPS/Register/register[20][18] ,
         \i_MIPS/Register/register[20][19] ,
         \i_MIPS/Register/register[20][20] ,
         \i_MIPS/Register/register[20][21] ,
         \i_MIPS/Register/register[20][22] ,
         \i_MIPS/Register/register[20][23] ,
         \i_MIPS/Register/register[20][24] ,
         \i_MIPS/Register/register[20][25] ,
         \i_MIPS/Register/register[20][26] ,
         \i_MIPS/Register/register[20][27] ,
         \i_MIPS/Register/register[20][28] ,
         \i_MIPS/Register/register[20][29] ,
         \i_MIPS/Register/register[20][30] ,
         \i_MIPS/Register/register[20][31] , \i_MIPS/Register/register[19][0] ,
         \i_MIPS/Register/register[19][1] , \i_MIPS/Register/register[19][2] ,
         \i_MIPS/Register/register[19][3] , \i_MIPS/Register/register[19][4] ,
         \i_MIPS/Register/register[19][5] , \i_MIPS/Register/register[19][6] ,
         \i_MIPS/Register/register[19][7] , \i_MIPS/Register/register[19][8] ,
         \i_MIPS/Register/register[19][9] , \i_MIPS/Register/register[19][10] ,
         \i_MIPS/Register/register[19][11] ,
         \i_MIPS/Register/register[19][12] ,
         \i_MIPS/Register/register[19][13] ,
         \i_MIPS/Register/register[19][14] ,
         \i_MIPS/Register/register[19][15] ,
         \i_MIPS/Register/register[19][16] ,
         \i_MIPS/Register/register[19][17] ,
         \i_MIPS/Register/register[19][18] ,
         \i_MIPS/Register/register[19][19] ,
         \i_MIPS/Register/register[19][20] ,
         \i_MIPS/Register/register[19][21] ,
         \i_MIPS/Register/register[19][22] ,
         \i_MIPS/Register/register[19][23] ,
         \i_MIPS/Register/register[19][24] ,
         \i_MIPS/Register/register[19][25] ,
         \i_MIPS/Register/register[19][26] ,
         \i_MIPS/Register/register[19][27] ,
         \i_MIPS/Register/register[19][28] ,
         \i_MIPS/Register/register[19][29] ,
         \i_MIPS/Register/register[19][30] ,
         \i_MIPS/Register/register[19][31] , \i_MIPS/Register/register[18][0] ,
         \i_MIPS/Register/register[18][1] , \i_MIPS/Register/register[18][2] ,
         \i_MIPS/Register/register[18][3] , \i_MIPS/Register/register[18][4] ,
         \i_MIPS/Register/register[18][5] , \i_MIPS/Register/register[18][6] ,
         \i_MIPS/Register/register[18][7] , \i_MIPS/Register/register[18][8] ,
         \i_MIPS/Register/register[18][9] , \i_MIPS/Register/register[18][10] ,
         \i_MIPS/Register/register[18][11] ,
         \i_MIPS/Register/register[18][12] ,
         \i_MIPS/Register/register[18][13] ,
         \i_MIPS/Register/register[18][14] ,
         \i_MIPS/Register/register[18][15] ,
         \i_MIPS/Register/register[18][16] ,
         \i_MIPS/Register/register[18][17] ,
         \i_MIPS/Register/register[18][18] ,
         \i_MIPS/Register/register[18][19] ,
         \i_MIPS/Register/register[18][20] ,
         \i_MIPS/Register/register[18][21] ,
         \i_MIPS/Register/register[18][22] ,
         \i_MIPS/Register/register[18][23] ,
         \i_MIPS/Register/register[18][24] ,
         \i_MIPS/Register/register[18][25] ,
         \i_MIPS/Register/register[18][26] ,
         \i_MIPS/Register/register[18][27] ,
         \i_MIPS/Register/register[18][28] ,
         \i_MIPS/Register/register[18][29] ,
         \i_MIPS/Register/register[18][30] ,
         \i_MIPS/Register/register[18][31] , \i_MIPS/Register/register[17][0] ,
         \i_MIPS/Register/register[17][1] , \i_MIPS/Register/register[17][2] ,
         \i_MIPS/Register/register[17][3] , \i_MIPS/Register/register[17][4] ,
         \i_MIPS/Register/register[17][5] , \i_MIPS/Register/register[17][6] ,
         \i_MIPS/Register/register[17][7] , \i_MIPS/Register/register[17][8] ,
         \i_MIPS/Register/register[17][9] , \i_MIPS/Register/register[17][10] ,
         \i_MIPS/Register/register[17][11] ,
         \i_MIPS/Register/register[17][12] ,
         \i_MIPS/Register/register[17][13] ,
         \i_MIPS/Register/register[17][14] ,
         \i_MIPS/Register/register[17][15] ,
         \i_MIPS/Register/register[17][16] ,
         \i_MIPS/Register/register[17][17] ,
         \i_MIPS/Register/register[17][18] ,
         \i_MIPS/Register/register[17][19] ,
         \i_MIPS/Register/register[17][20] ,
         \i_MIPS/Register/register[17][21] ,
         \i_MIPS/Register/register[17][22] ,
         \i_MIPS/Register/register[17][23] ,
         \i_MIPS/Register/register[17][24] ,
         \i_MIPS/Register/register[17][25] ,
         \i_MIPS/Register/register[17][26] ,
         \i_MIPS/Register/register[17][27] ,
         \i_MIPS/Register/register[17][28] ,
         \i_MIPS/Register/register[17][29] ,
         \i_MIPS/Register/register[17][30] ,
         \i_MIPS/Register/register[17][31] , \i_MIPS/Register/register[16][0] ,
         \i_MIPS/Register/register[16][1] , \i_MIPS/Register/register[16][2] ,
         \i_MIPS/Register/register[16][3] , \i_MIPS/Register/register[16][4] ,
         \i_MIPS/Register/register[16][5] , \i_MIPS/Register/register[16][6] ,
         \i_MIPS/Register/register[16][7] , \i_MIPS/Register/register[16][8] ,
         \i_MIPS/Register/register[16][9] , \i_MIPS/Register/register[16][10] ,
         \i_MIPS/Register/register[16][11] ,
         \i_MIPS/Register/register[16][12] ,
         \i_MIPS/Register/register[16][13] ,
         \i_MIPS/Register/register[16][14] ,
         \i_MIPS/Register/register[16][15] ,
         \i_MIPS/Register/register[16][16] ,
         \i_MIPS/Register/register[16][17] ,
         \i_MIPS/Register/register[16][18] ,
         \i_MIPS/Register/register[16][19] ,
         \i_MIPS/Register/register[16][20] ,
         \i_MIPS/Register/register[16][21] ,
         \i_MIPS/Register/register[16][22] ,
         \i_MIPS/Register/register[16][23] ,
         \i_MIPS/Register/register[16][24] ,
         \i_MIPS/Register/register[16][25] ,
         \i_MIPS/Register/register[16][26] ,
         \i_MIPS/Register/register[16][27] ,
         \i_MIPS/Register/register[16][28] ,
         \i_MIPS/Register/register[16][29] ,
         \i_MIPS/Register/register[16][30] ,
         \i_MIPS/Register/register[16][31] , \i_MIPS/Register/register[15][0] ,
         \i_MIPS/Register/register[15][1] , \i_MIPS/Register/register[15][2] ,
         \i_MIPS/Register/register[15][3] , \i_MIPS/Register/register[15][4] ,
         \i_MIPS/Register/register[15][5] , \i_MIPS/Register/register[15][6] ,
         \i_MIPS/Register/register[15][7] , \i_MIPS/Register/register[15][8] ,
         \i_MIPS/Register/register[15][9] , \i_MIPS/Register/register[15][10] ,
         \i_MIPS/Register/register[15][11] ,
         \i_MIPS/Register/register[15][12] ,
         \i_MIPS/Register/register[15][13] ,
         \i_MIPS/Register/register[15][14] ,
         \i_MIPS/Register/register[15][15] ,
         \i_MIPS/Register/register[15][16] ,
         \i_MIPS/Register/register[15][17] ,
         \i_MIPS/Register/register[15][18] ,
         \i_MIPS/Register/register[15][19] ,
         \i_MIPS/Register/register[15][20] ,
         \i_MIPS/Register/register[15][21] ,
         \i_MIPS/Register/register[15][22] ,
         \i_MIPS/Register/register[15][23] ,
         \i_MIPS/Register/register[15][24] ,
         \i_MIPS/Register/register[15][25] ,
         \i_MIPS/Register/register[15][26] ,
         \i_MIPS/Register/register[15][27] ,
         \i_MIPS/Register/register[15][28] ,
         \i_MIPS/Register/register[15][29] ,
         \i_MIPS/Register/register[15][30] ,
         \i_MIPS/Register/register[15][31] , \i_MIPS/Register/register[14][0] ,
         \i_MIPS/Register/register[14][1] , \i_MIPS/Register/register[14][2] ,
         \i_MIPS/Register/register[14][3] , \i_MIPS/Register/register[14][4] ,
         \i_MIPS/Register/register[14][5] , \i_MIPS/Register/register[14][6] ,
         \i_MIPS/Register/register[14][7] , \i_MIPS/Register/register[14][8] ,
         \i_MIPS/Register/register[14][9] , \i_MIPS/Register/register[14][10] ,
         \i_MIPS/Register/register[14][11] ,
         \i_MIPS/Register/register[14][12] ,
         \i_MIPS/Register/register[14][13] ,
         \i_MIPS/Register/register[14][14] ,
         \i_MIPS/Register/register[14][15] ,
         \i_MIPS/Register/register[14][16] ,
         \i_MIPS/Register/register[14][17] ,
         \i_MIPS/Register/register[14][18] ,
         \i_MIPS/Register/register[14][19] ,
         \i_MIPS/Register/register[14][20] ,
         \i_MIPS/Register/register[14][21] ,
         \i_MIPS/Register/register[14][22] ,
         \i_MIPS/Register/register[14][23] ,
         \i_MIPS/Register/register[14][24] ,
         \i_MIPS/Register/register[14][25] ,
         \i_MIPS/Register/register[14][26] ,
         \i_MIPS/Register/register[14][27] ,
         \i_MIPS/Register/register[14][28] ,
         \i_MIPS/Register/register[14][29] ,
         \i_MIPS/Register/register[14][30] ,
         \i_MIPS/Register/register[14][31] , \i_MIPS/Register/register[13][0] ,
         \i_MIPS/Register/register[13][1] , \i_MIPS/Register/register[13][2] ,
         \i_MIPS/Register/register[13][3] , \i_MIPS/Register/register[13][4] ,
         \i_MIPS/Register/register[13][5] , \i_MIPS/Register/register[13][6] ,
         \i_MIPS/Register/register[13][7] , \i_MIPS/Register/register[13][8] ,
         \i_MIPS/Register/register[13][9] , \i_MIPS/Register/register[13][10] ,
         \i_MIPS/Register/register[13][11] ,
         \i_MIPS/Register/register[13][12] ,
         \i_MIPS/Register/register[13][13] ,
         \i_MIPS/Register/register[13][14] ,
         \i_MIPS/Register/register[13][15] ,
         \i_MIPS/Register/register[13][16] ,
         \i_MIPS/Register/register[13][17] ,
         \i_MIPS/Register/register[13][18] ,
         \i_MIPS/Register/register[13][19] ,
         \i_MIPS/Register/register[13][20] ,
         \i_MIPS/Register/register[13][21] ,
         \i_MIPS/Register/register[13][22] ,
         \i_MIPS/Register/register[13][23] ,
         \i_MIPS/Register/register[13][24] ,
         \i_MIPS/Register/register[13][25] ,
         \i_MIPS/Register/register[13][26] ,
         \i_MIPS/Register/register[13][27] ,
         \i_MIPS/Register/register[13][28] ,
         \i_MIPS/Register/register[13][29] ,
         \i_MIPS/Register/register[13][30] ,
         \i_MIPS/Register/register[13][31] , \i_MIPS/Register/register[12][0] ,
         \i_MIPS/Register/register[12][1] , \i_MIPS/Register/register[12][2] ,
         \i_MIPS/Register/register[12][3] , \i_MIPS/Register/register[12][4] ,
         \i_MIPS/Register/register[12][5] , \i_MIPS/Register/register[12][6] ,
         \i_MIPS/Register/register[12][7] , \i_MIPS/Register/register[12][8] ,
         \i_MIPS/Register/register[12][9] , \i_MIPS/Register/register[12][10] ,
         \i_MIPS/Register/register[12][11] ,
         \i_MIPS/Register/register[12][12] ,
         \i_MIPS/Register/register[12][13] ,
         \i_MIPS/Register/register[12][14] ,
         \i_MIPS/Register/register[12][15] ,
         \i_MIPS/Register/register[12][16] ,
         \i_MIPS/Register/register[12][17] ,
         \i_MIPS/Register/register[12][18] ,
         \i_MIPS/Register/register[12][19] ,
         \i_MIPS/Register/register[12][20] ,
         \i_MIPS/Register/register[12][21] ,
         \i_MIPS/Register/register[12][22] ,
         \i_MIPS/Register/register[12][23] ,
         \i_MIPS/Register/register[12][24] ,
         \i_MIPS/Register/register[12][25] ,
         \i_MIPS/Register/register[12][26] ,
         \i_MIPS/Register/register[12][27] ,
         \i_MIPS/Register/register[12][28] ,
         \i_MIPS/Register/register[12][29] ,
         \i_MIPS/Register/register[12][30] ,
         \i_MIPS/Register/register[12][31] , \i_MIPS/Register/register[11][0] ,
         \i_MIPS/Register/register[11][1] , \i_MIPS/Register/register[11][2] ,
         \i_MIPS/Register/register[11][3] , \i_MIPS/Register/register[11][4] ,
         \i_MIPS/Register/register[11][5] , \i_MIPS/Register/register[11][6] ,
         \i_MIPS/Register/register[11][7] , \i_MIPS/Register/register[11][8] ,
         \i_MIPS/Register/register[11][9] , \i_MIPS/Register/register[11][10] ,
         \i_MIPS/Register/register[11][11] ,
         \i_MIPS/Register/register[11][12] ,
         \i_MIPS/Register/register[11][13] ,
         \i_MIPS/Register/register[11][14] ,
         \i_MIPS/Register/register[11][15] ,
         \i_MIPS/Register/register[11][16] ,
         \i_MIPS/Register/register[11][17] ,
         \i_MIPS/Register/register[11][18] ,
         \i_MIPS/Register/register[11][19] ,
         \i_MIPS/Register/register[11][20] ,
         \i_MIPS/Register/register[11][21] ,
         \i_MIPS/Register/register[11][22] ,
         \i_MIPS/Register/register[11][23] ,
         \i_MIPS/Register/register[11][24] ,
         \i_MIPS/Register/register[11][25] ,
         \i_MIPS/Register/register[11][26] ,
         \i_MIPS/Register/register[11][27] ,
         \i_MIPS/Register/register[11][28] ,
         \i_MIPS/Register/register[11][29] ,
         \i_MIPS/Register/register[11][30] ,
         \i_MIPS/Register/register[11][31] , \i_MIPS/Register/register[10][0] ,
         \i_MIPS/Register/register[10][1] , \i_MIPS/Register/register[10][2] ,
         \i_MIPS/Register/register[10][3] , \i_MIPS/Register/register[10][4] ,
         \i_MIPS/Register/register[10][5] , \i_MIPS/Register/register[10][6] ,
         \i_MIPS/Register/register[10][7] , \i_MIPS/Register/register[10][8] ,
         \i_MIPS/Register/register[10][9] , \i_MIPS/Register/register[10][10] ,
         \i_MIPS/Register/register[10][11] ,
         \i_MIPS/Register/register[10][12] ,
         \i_MIPS/Register/register[10][13] ,
         \i_MIPS/Register/register[10][14] ,
         \i_MIPS/Register/register[10][15] ,
         \i_MIPS/Register/register[10][16] ,
         \i_MIPS/Register/register[10][17] ,
         \i_MIPS/Register/register[10][18] ,
         \i_MIPS/Register/register[10][19] ,
         \i_MIPS/Register/register[10][20] ,
         \i_MIPS/Register/register[10][21] ,
         \i_MIPS/Register/register[10][22] ,
         \i_MIPS/Register/register[10][23] ,
         \i_MIPS/Register/register[10][24] ,
         \i_MIPS/Register/register[10][25] ,
         \i_MIPS/Register/register[10][26] ,
         \i_MIPS/Register/register[10][27] ,
         \i_MIPS/Register/register[10][28] ,
         \i_MIPS/Register/register[10][29] ,
         \i_MIPS/Register/register[10][30] ,
         \i_MIPS/Register/register[10][31] , \i_MIPS/Register/register[9][0] ,
         \i_MIPS/Register/register[9][1] , \i_MIPS/Register/register[9][2] ,
         \i_MIPS/Register/register[9][3] , \i_MIPS/Register/register[9][4] ,
         \i_MIPS/Register/register[9][5] , \i_MIPS/Register/register[9][6] ,
         \i_MIPS/Register/register[9][7] , \i_MIPS/Register/register[9][8] ,
         \i_MIPS/Register/register[9][9] , \i_MIPS/Register/register[9][10] ,
         \i_MIPS/Register/register[9][11] , \i_MIPS/Register/register[9][12] ,
         \i_MIPS/Register/register[9][13] , \i_MIPS/Register/register[9][14] ,
         \i_MIPS/Register/register[9][15] , \i_MIPS/Register/register[9][16] ,
         \i_MIPS/Register/register[9][17] , \i_MIPS/Register/register[9][18] ,
         \i_MIPS/Register/register[9][19] , \i_MIPS/Register/register[9][20] ,
         \i_MIPS/Register/register[9][21] , \i_MIPS/Register/register[9][22] ,
         \i_MIPS/Register/register[9][23] , \i_MIPS/Register/register[9][24] ,
         \i_MIPS/Register/register[9][25] , \i_MIPS/Register/register[9][26] ,
         \i_MIPS/Register/register[9][27] , \i_MIPS/Register/register[9][28] ,
         \i_MIPS/Register/register[9][29] , \i_MIPS/Register/register[9][30] ,
         \i_MIPS/Register/register[9][31] , \i_MIPS/Register/register[8][0] ,
         \i_MIPS/Register/register[8][1] , \i_MIPS/Register/register[8][2] ,
         \i_MIPS/Register/register[8][3] , \i_MIPS/Register/register[8][4] ,
         \i_MIPS/Register/register[8][5] , \i_MIPS/Register/register[8][6] ,
         \i_MIPS/Register/register[8][7] , \i_MIPS/Register/register[8][8] ,
         \i_MIPS/Register/register[8][9] , \i_MIPS/Register/register[8][10] ,
         \i_MIPS/Register/register[8][11] , \i_MIPS/Register/register[8][12] ,
         \i_MIPS/Register/register[8][13] , \i_MIPS/Register/register[8][14] ,
         \i_MIPS/Register/register[8][15] , \i_MIPS/Register/register[8][16] ,
         \i_MIPS/Register/register[8][17] , \i_MIPS/Register/register[8][18] ,
         \i_MIPS/Register/register[8][19] , \i_MIPS/Register/register[8][20] ,
         \i_MIPS/Register/register[8][21] , \i_MIPS/Register/register[8][22] ,
         \i_MIPS/Register/register[8][23] , \i_MIPS/Register/register[8][24] ,
         \i_MIPS/Register/register[8][25] , \i_MIPS/Register/register[8][26] ,
         \i_MIPS/Register/register[8][27] , \i_MIPS/Register/register[8][28] ,
         \i_MIPS/Register/register[8][29] , \i_MIPS/Register/register[8][30] ,
         \i_MIPS/Register/register[8][31] , \i_MIPS/Register/register[7][0] ,
         \i_MIPS/Register/register[7][1] , \i_MIPS/Register/register[7][2] ,
         \i_MIPS/Register/register[7][3] , \i_MIPS/Register/register[7][4] ,
         \i_MIPS/Register/register[7][5] , \i_MIPS/Register/register[7][6] ,
         \i_MIPS/Register/register[7][7] , \i_MIPS/Register/register[7][8] ,
         \i_MIPS/Register/register[7][9] , \i_MIPS/Register/register[7][10] ,
         \i_MIPS/Register/register[7][11] , \i_MIPS/Register/register[7][12] ,
         \i_MIPS/Register/register[7][13] , \i_MIPS/Register/register[7][14] ,
         \i_MIPS/Register/register[7][15] , \i_MIPS/Register/register[7][16] ,
         \i_MIPS/Register/register[7][17] , \i_MIPS/Register/register[7][18] ,
         \i_MIPS/Register/register[7][19] , \i_MIPS/Register/register[7][20] ,
         \i_MIPS/Register/register[7][21] , \i_MIPS/Register/register[7][22] ,
         \i_MIPS/Register/register[7][23] , \i_MIPS/Register/register[7][24] ,
         \i_MIPS/Register/register[7][25] , \i_MIPS/Register/register[7][26] ,
         \i_MIPS/Register/register[7][27] , \i_MIPS/Register/register[7][28] ,
         \i_MIPS/Register/register[7][29] , \i_MIPS/Register/register[7][30] ,
         \i_MIPS/Register/register[7][31] , \i_MIPS/Register/register[6][0] ,
         \i_MIPS/Register/register[6][1] , \i_MIPS/Register/register[6][2] ,
         \i_MIPS/Register/register[6][3] , \i_MIPS/Register/register[6][4] ,
         \i_MIPS/Register/register[6][5] , \i_MIPS/Register/register[6][6] ,
         \i_MIPS/Register/register[6][7] , \i_MIPS/Register/register[6][8] ,
         \i_MIPS/Register/register[6][9] , \i_MIPS/Register/register[6][10] ,
         \i_MIPS/Register/register[6][11] , \i_MIPS/Register/register[6][12] ,
         \i_MIPS/Register/register[6][13] , \i_MIPS/Register/register[6][14] ,
         \i_MIPS/Register/register[6][15] , \i_MIPS/Register/register[6][16] ,
         \i_MIPS/Register/register[6][17] , \i_MIPS/Register/register[6][18] ,
         \i_MIPS/Register/register[6][19] , \i_MIPS/Register/register[6][20] ,
         \i_MIPS/Register/register[6][21] , \i_MIPS/Register/register[6][22] ,
         \i_MIPS/Register/register[6][23] , \i_MIPS/Register/register[6][24] ,
         \i_MIPS/Register/register[6][25] , \i_MIPS/Register/register[6][26] ,
         \i_MIPS/Register/register[6][27] , \i_MIPS/Register/register[6][28] ,
         \i_MIPS/Register/register[6][29] , \i_MIPS/Register/register[6][30] ,
         \i_MIPS/Register/register[6][31] , \i_MIPS/Register/register[5][0] ,
         \i_MIPS/Register/register[5][1] , \i_MIPS/Register/register[5][2] ,
         \i_MIPS/Register/register[5][3] , \i_MIPS/Register/register[5][4] ,
         \i_MIPS/Register/register[5][5] , \i_MIPS/Register/register[5][6] ,
         \i_MIPS/Register/register[5][7] , \i_MIPS/Register/register[5][8] ,
         \i_MIPS/Register/register[5][9] , \i_MIPS/Register/register[5][10] ,
         \i_MIPS/Register/register[5][11] , \i_MIPS/Register/register[5][12] ,
         \i_MIPS/Register/register[5][13] , \i_MIPS/Register/register[5][14] ,
         \i_MIPS/Register/register[5][15] , \i_MIPS/Register/register[5][16] ,
         \i_MIPS/Register/register[5][17] , \i_MIPS/Register/register[5][18] ,
         \i_MIPS/Register/register[5][19] , \i_MIPS/Register/register[5][20] ,
         \i_MIPS/Register/register[5][21] , \i_MIPS/Register/register[5][22] ,
         \i_MIPS/Register/register[5][23] , \i_MIPS/Register/register[5][24] ,
         \i_MIPS/Register/register[5][25] , \i_MIPS/Register/register[5][26] ,
         \i_MIPS/Register/register[5][27] , \i_MIPS/Register/register[5][28] ,
         \i_MIPS/Register/register[5][29] , \i_MIPS/Register/register[5][30] ,
         \i_MIPS/Register/register[5][31] , \i_MIPS/Register/register[4][0] ,
         \i_MIPS/Register/register[4][1] , \i_MIPS/Register/register[4][2] ,
         \i_MIPS/Register/register[4][3] , \i_MIPS/Register/register[4][4] ,
         \i_MIPS/Register/register[4][5] , \i_MIPS/Register/register[4][6] ,
         \i_MIPS/Register/register[4][7] , \i_MIPS/Register/register[4][8] ,
         \i_MIPS/Register/register[4][9] , \i_MIPS/Register/register[4][10] ,
         \i_MIPS/Register/register[4][11] , \i_MIPS/Register/register[4][12] ,
         \i_MIPS/Register/register[4][13] , \i_MIPS/Register/register[4][14] ,
         \i_MIPS/Register/register[4][15] , \i_MIPS/Register/register[4][16] ,
         \i_MIPS/Register/register[4][17] , \i_MIPS/Register/register[4][18] ,
         \i_MIPS/Register/register[4][19] , \i_MIPS/Register/register[4][20] ,
         \i_MIPS/Register/register[4][21] , \i_MIPS/Register/register[4][22] ,
         \i_MIPS/Register/register[4][23] , \i_MIPS/Register/register[4][24] ,
         \i_MIPS/Register/register[4][25] , \i_MIPS/Register/register[4][26] ,
         \i_MIPS/Register/register[4][27] , \i_MIPS/Register/register[4][28] ,
         \i_MIPS/Register/register[4][29] , \i_MIPS/Register/register[4][30] ,
         \i_MIPS/Register/register[4][31] , \i_MIPS/Register/register[3][0] ,
         \i_MIPS/Register/register[3][1] , \i_MIPS/Register/register[3][2] ,
         \i_MIPS/Register/register[3][3] , \i_MIPS/Register/register[3][4] ,
         \i_MIPS/Register/register[3][5] , \i_MIPS/Register/register[3][6] ,
         \i_MIPS/Register/register[3][7] , \i_MIPS/Register/register[3][8] ,
         \i_MIPS/Register/register[3][9] , \i_MIPS/Register/register[3][10] ,
         \i_MIPS/Register/register[3][11] , \i_MIPS/Register/register[3][12] ,
         \i_MIPS/Register/register[3][13] , \i_MIPS/Register/register[3][14] ,
         \i_MIPS/Register/register[3][15] , \i_MIPS/Register/register[3][16] ,
         \i_MIPS/Register/register[3][17] , \i_MIPS/Register/register[3][18] ,
         \i_MIPS/Register/register[3][19] , \i_MIPS/Register/register[3][20] ,
         \i_MIPS/Register/register[3][21] , \i_MIPS/Register/register[3][22] ,
         \i_MIPS/Register/register[3][23] , \i_MIPS/Register/register[3][24] ,
         \i_MIPS/Register/register[3][25] , \i_MIPS/Register/register[3][26] ,
         \i_MIPS/Register/register[3][27] , \i_MIPS/Register/register[3][28] ,
         \i_MIPS/Register/register[3][29] , \i_MIPS/Register/register[3][30] ,
         \i_MIPS/Register/register[3][31] , \i_MIPS/Register/register[2][0] ,
         \i_MIPS/Register/register[2][1] , \i_MIPS/Register/register[2][2] ,
         \i_MIPS/Register/register[2][3] , \i_MIPS/Register/register[2][4] ,
         \i_MIPS/Register/register[2][5] , \i_MIPS/Register/register[2][6] ,
         \i_MIPS/Register/register[2][7] , \i_MIPS/Register/register[2][8] ,
         \i_MIPS/Register/register[2][9] , \i_MIPS/Register/register[2][10] ,
         \i_MIPS/Register/register[2][11] , \i_MIPS/Register/register[2][12] ,
         \i_MIPS/Register/register[2][13] , \i_MIPS/Register/register[2][14] ,
         \i_MIPS/Register/register[2][15] , \i_MIPS/Register/register[2][16] ,
         \i_MIPS/Register/register[2][17] , \i_MIPS/Register/register[2][18] ,
         \i_MIPS/Register/register[2][19] , \i_MIPS/Register/register[2][20] ,
         \i_MIPS/Register/register[2][21] , \i_MIPS/Register/register[2][22] ,
         \i_MIPS/Register/register[2][23] , \i_MIPS/Register/register[2][24] ,
         \i_MIPS/Register/register[2][25] , \i_MIPS/Register/register[2][26] ,
         \i_MIPS/Register/register[2][27] , \i_MIPS/Register/register[2][28] ,
         \i_MIPS/Register/register[2][29] , \i_MIPS/Register/register[2][30] ,
         \i_MIPS/Register/register[2][31] , \i_MIPS/Register/register[1][0] ,
         \i_MIPS/Register/register[1][1] , \i_MIPS/Register/register[1][2] ,
         \i_MIPS/Register/register[1][3] , \i_MIPS/Register/register[1][4] ,
         \i_MIPS/Register/register[1][5] , \i_MIPS/Register/register[1][6] ,
         \i_MIPS/Register/register[1][7] , \i_MIPS/Register/register[1][8] ,
         \i_MIPS/Register/register[1][9] , \i_MIPS/Register/register[1][10] ,
         \i_MIPS/Register/register[1][11] , \i_MIPS/Register/register[1][12] ,
         \i_MIPS/Register/register[1][13] , \i_MIPS/Register/register[1][14] ,
         \i_MIPS/Register/register[1][15] , \i_MIPS/Register/register[1][16] ,
         \i_MIPS/Register/register[1][17] , \i_MIPS/Register/register[1][18] ,
         \i_MIPS/Register/register[1][19] , \i_MIPS/Register/register[1][20] ,
         \i_MIPS/Register/register[1][21] , \i_MIPS/Register/register[1][22] ,
         \i_MIPS/Register/register[1][23] , \i_MIPS/Register/register[1][24] ,
         \i_MIPS/Register/register[1][25] , \i_MIPS/Register/register[1][26] ,
         \i_MIPS/Register/register[1][27] , \i_MIPS/Register/register[1][28] ,
         \i_MIPS/Register/register[1][29] , \i_MIPS/Register/register[1][30] ,
         \i_MIPS/Register/register[1][31] , \i_MIPS/Register/register[0][0] ,
         \i_MIPS/Register/register[0][1] , \i_MIPS/Register/register[0][2] ,
         \i_MIPS/Register/register[0][3] , \i_MIPS/Register/register[0][4] ,
         \i_MIPS/Register/register[0][5] , \i_MIPS/Register/register[0][6] ,
         \i_MIPS/Register/register[0][7] , \i_MIPS/Register/register[0][8] ,
         \i_MIPS/Register/register[0][9] , \i_MIPS/Register/register[0][10] ,
         \i_MIPS/Register/register[0][11] , \i_MIPS/Register/register[0][12] ,
         \i_MIPS/Register/register[0][13] , \i_MIPS/Register/register[0][14] ,
         \i_MIPS/Register/register[0][15] , \i_MIPS/Register/register[0][16] ,
         \i_MIPS/Register/register[0][17] , \i_MIPS/Register/register[0][18] ,
         \i_MIPS/Register/register[0][19] , \i_MIPS/Register/register[0][20] ,
         \i_MIPS/Register/register[0][21] , \i_MIPS/Register/register[0][22] ,
         \i_MIPS/Register/register[0][23] , \i_MIPS/Register/register[0][24] ,
         \i_MIPS/Register/register[0][25] , \i_MIPS/Register/register[0][26] ,
         \i_MIPS/Register/register[0][27] , \i_MIPS/Register/register[0][28] ,
         \i_MIPS/Register/register[0][29] , \i_MIPS/Register/register[0][30] ,
         \i_MIPS/Register/register[0][31] , \i_MIPS/Control/n14 ,
         \i_MIPS/Control/n10 , \i_MIPS/Hazard_detection/n13 ,
         \i_MIPS/Hazard_detection/n12 , \i_MIPS/Hazard_detection/n11 ,
         \i_MIPS/Hazard_detection/n10 , \i_MIPS/Hazard_detection/n9 ,
         \i_MIPS/Hazard_detection/n8 , \i_MIPS/Hazard_detection/n7 ,
         \i_MIPS/Hazard_detection/n4 , \i_MIPS/forward_unit/n25 ,
         \i_MIPS/forward_unit/n10 , \i_MIPS/ALU_Control/n20 ,
         \i_MIPS/ALU_Control/n18 , \i_MIPS/ALU/N303 , \I_cache/cache[7][0] ,
         \I_cache/cache[7][1] , \I_cache/cache[7][2] , \I_cache/cache[7][3] ,
         \I_cache/cache[7][4] , \I_cache/cache[7][5] , \I_cache/cache[7][6] ,
         \I_cache/cache[7][7] , \I_cache/cache[7][8] , \I_cache/cache[7][9] ,
         \I_cache/cache[7][10] , \I_cache/cache[7][11] ,
         \I_cache/cache[7][12] , \I_cache/cache[7][13] ,
         \I_cache/cache[7][14] , \I_cache/cache[7][15] ,
         \I_cache/cache[7][16] , \I_cache/cache[7][17] ,
         \I_cache/cache[7][18] , \I_cache/cache[7][19] ,
         \I_cache/cache[7][20] , \I_cache/cache[7][21] ,
         \I_cache/cache[7][22] , \I_cache/cache[7][23] ,
         \I_cache/cache[7][24] , \I_cache/cache[7][25] ,
         \I_cache/cache[7][26] , \I_cache/cache[7][27] ,
         \I_cache/cache[7][28] , \I_cache/cache[7][29] ,
         \I_cache/cache[7][30] , \I_cache/cache[7][31] ,
         \I_cache/cache[7][32] , \I_cache/cache[7][33] ,
         \I_cache/cache[7][34] , \I_cache/cache[7][35] ,
         \I_cache/cache[7][36] , \I_cache/cache[7][37] ,
         \I_cache/cache[7][38] , \I_cache/cache[7][39] ,
         \I_cache/cache[7][40] , \I_cache/cache[7][41] ,
         \I_cache/cache[7][42] , \I_cache/cache[7][43] ,
         \I_cache/cache[7][44] , \I_cache/cache[7][45] ,
         \I_cache/cache[7][46] , \I_cache/cache[7][47] ,
         \I_cache/cache[7][48] , \I_cache/cache[7][49] ,
         \I_cache/cache[7][50] , \I_cache/cache[7][51] ,
         \I_cache/cache[7][52] , \I_cache/cache[7][53] ,
         \I_cache/cache[7][54] , \I_cache/cache[7][55] ,
         \I_cache/cache[7][56] , \I_cache/cache[7][57] ,
         \I_cache/cache[7][58] , \I_cache/cache[7][59] ,
         \I_cache/cache[7][60] , \I_cache/cache[7][61] ,
         \I_cache/cache[7][62] , \I_cache/cache[7][63] ,
         \I_cache/cache[7][64] , \I_cache/cache[7][65] ,
         \I_cache/cache[7][66] , \I_cache/cache[7][67] ,
         \I_cache/cache[7][68] , \I_cache/cache[7][69] ,
         \I_cache/cache[7][70] , \I_cache/cache[7][71] ,
         \I_cache/cache[7][72] , \I_cache/cache[7][73] ,
         \I_cache/cache[7][74] , \I_cache/cache[7][75] ,
         \I_cache/cache[7][76] , \I_cache/cache[7][77] ,
         \I_cache/cache[7][78] , \I_cache/cache[7][79] ,
         \I_cache/cache[7][80] , \I_cache/cache[7][81] ,
         \I_cache/cache[7][82] , \I_cache/cache[7][83] ,
         \I_cache/cache[7][84] , \I_cache/cache[7][85] ,
         \I_cache/cache[7][86] , \I_cache/cache[7][87] ,
         \I_cache/cache[7][88] , \I_cache/cache[7][89] ,
         \I_cache/cache[7][90] , \I_cache/cache[7][91] ,
         \I_cache/cache[7][92] , \I_cache/cache[7][93] ,
         \I_cache/cache[7][94] , \I_cache/cache[7][95] ,
         \I_cache/cache[7][96] , \I_cache/cache[7][97] ,
         \I_cache/cache[7][98] , \I_cache/cache[7][99] ,
         \I_cache/cache[7][100] , \I_cache/cache[7][101] ,
         \I_cache/cache[7][102] , \I_cache/cache[7][103] ,
         \I_cache/cache[7][104] , \I_cache/cache[7][105] ,
         \I_cache/cache[7][106] , \I_cache/cache[7][107] ,
         \I_cache/cache[7][108] , \I_cache/cache[7][109] ,
         \I_cache/cache[7][110] , \I_cache/cache[7][111] ,
         \I_cache/cache[7][112] , \I_cache/cache[7][113] ,
         \I_cache/cache[7][114] , \I_cache/cache[7][115] ,
         \I_cache/cache[7][116] , \I_cache/cache[7][117] ,
         \I_cache/cache[7][118] , \I_cache/cache[7][119] ,
         \I_cache/cache[7][120] , \I_cache/cache[7][121] ,
         \I_cache/cache[7][122] , \I_cache/cache[7][123] ,
         \I_cache/cache[7][124] , \I_cache/cache[7][125] ,
         \I_cache/cache[7][126] , \I_cache/cache[7][127] ,
         \I_cache/cache[7][128] , \I_cache/cache[7][129] ,
         \I_cache/cache[7][130] , \I_cache/cache[7][131] ,
         \I_cache/cache[7][132] , \I_cache/cache[7][133] ,
         \I_cache/cache[7][134] , \I_cache/cache[7][135] ,
         \I_cache/cache[7][136] , \I_cache/cache[7][137] ,
         \I_cache/cache[7][138] , \I_cache/cache[7][139] ,
         \I_cache/cache[7][140] , \I_cache/cache[7][141] ,
         \I_cache/cache[7][142] , \I_cache/cache[7][143] ,
         \I_cache/cache[7][144] , \I_cache/cache[7][145] ,
         \I_cache/cache[7][146] , \I_cache/cache[7][147] ,
         \I_cache/cache[7][148] , \I_cache/cache[7][149] ,
         \I_cache/cache[7][150] , \I_cache/cache[7][151] ,
         \I_cache/cache[7][152] , \I_cache/cache[7][153] ,
         \I_cache/cache[7][154] , \I_cache/cache[6][0] , \I_cache/cache[6][1] ,
         \I_cache/cache[6][2] , \I_cache/cache[6][3] , \I_cache/cache[6][4] ,
         \I_cache/cache[6][5] , \I_cache/cache[6][6] , \I_cache/cache[6][7] ,
         \I_cache/cache[6][8] , \I_cache/cache[6][9] , \I_cache/cache[6][10] ,
         \I_cache/cache[6][11] , \I_cache/cache[6][12] ,
         \I_cache/cache[6][13] , \I_cache/cache[6][14] ,
         \I_cache/cache[6][15] , \I_cache/cache[6][16] ,
         \I_cache/cache[6][17] , \I_cache/cache[6][18] ,
         \I_cache/cache[6][19] , \I_cache/cache[6][20] ,
         \I_cache/cache[6][21] , \I_cache/cache[6][22] ,
         \I_cache/cache[6][23] , \I_cache/cache[6][24] ,
         \I_cache/cache[6][25] , \I_cache/cache[6][26] ,
         \I_cache/cache[6][27] , \I_cache/cache[6][28] ,
         \I_cache/cache[6][29] , \I_cache/cache[6][30] ,
         \I_cache/cache[6][31] , \I_cache/cache[6][32] ,
         \I_cache/cache[6][33] , \I_cache/cache[6][34] ,
         \I_cache/cache[6][35] , \I_cache/cache[6][36] ,
         \I_cache/cache[6][37] , \I_cache/cache[6][38] ,
         \I_cache/cache[6][39] , \I_cache/cache[6][40] ,
         \I_cache/cache[6][41] , \I_cache/cache[6][42] ,
         \I_cache/cache[6][43] , \I_cache/cache[6][44] ,
         \I_cache/cache[6][45] , \I_cache/cache[6][46] ,
         \I_cache/cache[6][47] , \I_cache/cache[6][48] ,
         \I_cache/cache[6][49] , \I_cache/cache[6][50] ,
         \I_cache/cache[6][51] , \I_cache/cache[6][52] ,
         \I_cache/cache[6][53] , \I_cache/cache[6][54] ,
         \I_cache/cache[6][55] , \I_cache/cache[6][56] ,
         \I_cache/cache[6][57] , \I_cache/cache[6][58] ,
         \I_cache/cache[6][59] , \I_cache/cache[6][60] ,
         \I_cache/cache[6][61] , \I_cache/cache[6][62] ,
         \I_cache/cache[6][63] , \I_cache/cache[6][64] ,
         \I_cache/cache[6][65] , \I_cache/cache[6][66] ,
         \I_cache/cache[6][67] , \I_cache/cache[6][68] ,
         \I_cache/cache[6][69] , \I_cache/cache[6][70] ,
         \I_cache/cache[6][71] , \I_cache/cache[6][72] ,
         \I_cache/cache[6][73] , \I_cache/cache[6][74] ,
         \I_cache/cache[6][75] , \I_cache/cache[6][76] ,
         \I_cache/cache[6][77] , \I_cache/cache[6][78] ,
         \I_cache/cache[6][79] , \I_cache/cache[6][80] ,
         \I_cache/cache[6][81] , \I_cache/cache[6][82] ,
         \I_cache/cache[6][83] , \I_cache/cache[6][84] ,
         \I_cache/cache[6][85] , \I_cache/cache[6][86] ,
         \I_cache/cache[6][87] , \I_cache/cache[6][88] ,
         \I_cache/cache[6][89] , \I_cache/cache[6][90] ,
         \I_cache/cache[6][91] , \I_cache/cache[6][92] ,
         \I_cache/cache[6][93] , \I_cache/cache[6][94] ,
         \I_cache/cache[6][95] , \I_cache/cache[6][96] ,
         \I_cache/cache[6][97] , \I_cache/cache[6][98] ,
         \I_cache/cache[6][99] , \I_cache/cache[6][100] ,
         \I_cache/cache[6][101] , \I_cache/cache[6][102] ,
         \I_cache/cache[6][103] , \I_cache/cache[6][104] ,
         \I_cache/cache[6][105] , \I_cache/cache[6][106] ,
         \I_cache/cache[6][107] , \I_cache/cache[6][108] ,
         \I_cache/cache[6][109] , \I_cache/cache[6][110] ,
         \I_cache/cache[6][111] , \I_cache/cache[6][112] ,
         \I_cache/cache[6][113] , \I_cache/cache[6][114] ,
         \I_cache/cache[6][115] , \I_cache/cache[6][116] ,
         \I_cache/cache[6][117] , \I_cache/cache[6][118] ,
         \I_cache/cache[6][119] , \I_cache/cache[6][120] ,
         \I_cache/cache[6][121] , \I_cache/cache[6][122] ,
         \I_cache/cache[6][123] , \I_cache/cache[6][124] ,
         \I_cache/cache[6][125] , \I_cache/cache[6][126] ,
         \I_cache/cache[6][127] , \I_cache/cache[6][128] ,
         \I_cache/cache[6][129] , \I_cache/cache[6][130] ,
         \I_cache/cache[6][131] , \I_cache/cache[6][132] ,
         \I_cache/cache[6][133] , \I_cache/cache[6][134] ,
         \I_cache/cache[6][135] , \I_cache/cache[6][136] ,
         \I_cache/cache[6][137] , \I_cache/cache[6][138] ,
         \I_cache/cache[6][139] , \I_cache/cache[6][140] ,
         \I_cache/cache[6][141] , \I_cache/cache[6][142] ,
         \I_cache/cache[6][143] , \I_cache/cache[6][144] ,
         \I_cache/cache[6][145] , \I_cache/cache[6][146] ,
         \I_cache/cache[6][147] , \I_cache/cache[6][148] ,
         \I_cache/cache[6][149] , \I_cache/cache[6][150] ,
         \I_cache/cache[6][151] , \I_cache/cache[6][152] ,
         \I_cache/cache[6][153] , \I_cache/cache[6][154] ,
         \I_cache/cache[5][0] , \I_cache/cache[5][1] , \I_cache/cache[5][2] ,
         \I_cache/cache[5][3] , \I_cache/cache[5][4] , \I_cache/cache[5][5] ,
         \I_cache/cache[5][6] , \I_cache/cache[5][7] , \I_cache/cache[5][8] ,
         \I_cache/cache[5][9] , \I_cache/cache[5][10] , \I_cache/cache[5][11] ,
         \I_cache/cache[5][12] , \I_cache/cache[5][13] ,
         \I_cache/cache[5][14] , \I_cache/cache[5][15] ,
         \I_cache/cache[5][16] , \I_cache/cache[5][17] ,
         \I_cache/cache[5][18] , \I_cache/cache[5][19] ,
         \I_cache/cache[5][20] , \I_cache/cache[5][21] ,
         \I_cache/cache[5][22] , \I_cache/cache[5][23] ,
         \I_cache/cache[5][24] , \I_cache/cache[5][25] ,
         \I_cache/cache[5][26] , \I_cache/cache[5][27] ,
         \I_cache/cache[5][28] , \I_cache/cache[5][29] ,
         \I_cache/cache[5][30] , \I_cache/cache[5][31] ,
         \I_cache/cache[5][32] , \I_cache/cache[5][33] ,
         \I_cache/cache[5][34] , \I_cache/cache[5][35] ,
         \I_cache/cache[5][36] , \I_cache/cache[5][37] ,
         \I_cache/cache[5][38] , \I_cache/cache[5][39] ,
         \I_cache/cache[5][40] , \I_cache/cache[5][41] ,
         \I_cache/cache[5][42] , \I_cache/cache[5][43] ,
         \I_cache/cache[5][44] , \I_cache/cache[5][45] ,
         \I_cache/cache[5][46] , \I_cache/cache[5][47] ,
         \I_cache/cache[5][48] , \I_cache/cache[5][49] ,
         \I_cache/cache[5][50] , \I_cache/cache[5][51] ,
         \I_cache/cache[5][52] , \I_cache/cache[5][53] ,
         \I_cache/cache[5][54] , \I_cache/cache[5][55] ,
         \I_cache/cache[5][56] , \I_cache/cache[5][57] ,
         \I_cache/cache[5][58] , \I_cache/cache[5][59] ,
         \I_cache/cache[5][60] , \I_cache/cache[5][61] ,
         \I_cache/cache[5][62] , \I_cache/cache[5][63] ,
         \I_cache/cache[5][64] , \I_cache/cache[5][65] ,
         \I_cache/cache[5][66] , \I_cache/cache[5][67] ,
         \I_cache/cache[5][68] , \I_cache/cache[5][69] ,
         \I_cache/cache[5][70] , \I_cache/cache[5][71] ,
         \I_cache/cache[5][72] , \I_cache/cache[5][73] ,
         \I_cache/cache[5][74] , \I_cache/cache[5][75] ,
         \I_cache/cache[5][76] , \I_cache/cache[5][77] ,
         \I_cache/cache[5][78] , \I_cache/cache[5][79] ,
         \I_cache/cache[5][80] , \I_cache/cache[5][81] ,
         \I_cache/cache[5][82] , \I_cache/cache[5][83] ,
         \I_cache/cache[5][84] , \I_cache/cache[5][85] ,
         \I_cache/cache[5][86] , \I_cache/cache[5][87] ,
         \I_cache/cache[5][88] , \I_cache/cache[5][89] ,
         \I_cache/cache[5][90] , \I_cache/cache[5][91] ,
         \I_cache/cache[5][92] , \I_cache/cache[5][93] ,
         \I_cache/cache[5][94] , \I_cache/cache[5][95] ,
         \I_cache/cache[5][96] , \I_cache/cache[5][97] ,
         \I_cache/cache[5][98] , \I_cache/cache[5][99] ,
         \I_cache/cache[5][100] , \I_cache/cache[5][101] ,
         \I_cache/cache[5][102] , \I_cache/cache[5][103] ,
         \I_cache/cache[5][104] , \I_cache/cache[5][105] ,
         \I_cache/cache[5][106] , \I_cache/cache[5][107] ,
         \I_cache/cache[5][108] , \I_cache/cache[5][109] ,
         \I_cache/cache[5][110] , \I_cache/cache[5][111] ,
         \I_cache/cache[5][112] , \I_cache/cache[5][113] ,
         \I_cache/cache[5][114] , \I_cache/cache[5][115] ,
         \I_cache/cache[5][116] , \I_cache/cache[5][117] ,
         \I_cache/cache[5][118] , \I_cache/cache[5][119] ,
         \I_cache/cache[5][120] , \I_cache/cache[5][121] ,
         \I_cache/cache[5][122] , \I_cache/cache[5][123] ,
         \I_cache/cache[5][124] , \I_cache/cache[5][125] ,
         \I_cache/cache[5][126] , \I_cache/cache[5][127] ,
         \I_cache/cache[5][128] , \I_cache/cache[5][129] ,
         \I_cache/cache[5][130] , \I_cache/cache[5][131] ,
         \I_cache/cache[5][132] , \I_cache/cache[5][133] ,
         \I_cache/cache[5][134] , \I_cache/cache[5][135] ,
         \I_cache/cache[5][136] , \I_cache/cache[5][137] ,
         \I_cache/cache[5][138] , \I_cache/cache[5][139] ,
         \I_cache/cache[5][140] , \I_cache/cache[5][141] ,
         \I_cache/cache[5][142] , \I_cache/cache[5][143] ,
         \I_cache/cache[5][144] , \I_cache/cache[5][145] ,
         \I_cache/cache[5][146] , \I_cache/cache[5][147] ,
         \I_cache/cache[5][148] , \I_cache/cache[5][149] ,
         \I_cache/cache[5][150] , \I_cache/cache[5][151] ,
         \I_cache/cache[5][152] , \I_cache/cache[5][153] ,
         \I_cache/cache[5][154] , \I_cache/cache[4][0] , \I_cache/cache[4][1] ,
         \I_cache/cache[4][2] , \I_cache/cache[4][3] , \I_cache/cache[4][4] ,
         \I_cache/cache[4][5] , \I_cache/cache[4][6] , \I_cache/cache[4][7] ,
         \I_cache/cache[4][8] , \I_cache/cache[4][9] , \I_cache/cache[4][10] ,
         \I_cache/cache[4][11] , \I_cache/cache[4][12] ,
         \I_cache/cache[4][13] , \I_cache/cache[4][14] ,
         \I_cache/cache[4][15] , \I_cache/cache[4][16] ,
         \I_cache/cache[4][17] , \I_cache/cache[4][18] ,
         \I_cache/cache[4][19] , \I_cache/cache[4][20] ,
         \I_cache/cache[4][21] , \I_cache/cache[4][22] ,
         \I_cache/cache[4][23] , \I_cache/cache[4][24] ,
         \I_cache/cache[4][25] , \I_cache/cache[4][26] ,
         \I_cache/cache[4][27] , \I_cache/cache[4][28] ,
         \I_cache/cache[4][29] , \I_cache/cache[4][30] ,
         \I_cache/cache[4][31] , \I_cache/cache[4][32] ,
         \I_cache/cache[4][33] , \I_cache/cache[4][34] ,
         \I_cache/cache[4][35] , \I_cache/cache[4][36] ,
         \I_cache/cache[4][37] , \I_cache/cache[4][38] ,
         \I_cache/cache[4][39] , \I_cache/cache[4][40] ,
         \I_cache/cache[4][41] , \I_cache/cache[4][42] ,
         \I_cache/cache[4][43] , \I_cache/cache[4][44] ,
         \I_cache/cache[4][45] , \I_cache/cache[4][46] ,
         \I_cache/cache[4][47] , \I_cache/cache[4][48] ,
         \I_cache/cache[4][49] , \I_cache/cache[4][50] ,
         \I_cache/cache[4][51] , \I_cache/cache[4][52] ,
         \I_cache/cache[4][53] , \I_cache/cache[4][54] ,
         \I_cache/cache[4][55] , \I_cache/cache[4][56] ,
         \I_cache/cache[4][57] , \I_cache/cache[4][58] ,
         \I_cache/cache[4][59] , \I_cache/cache[4][60] ,
         \I_cache/cache[4][61] , \I_cache/cache[4][62] ,
         \I_cache/cache[4][63] , \I_cache/cache[4][64] ,
         \I_cache/cache[4][65] , \I_cache/cache[4][66] ,
         \I_cache/cache[4][67] , \I_cache/cache[4][68] ,
         \I_cache/cache[4][69] , \I_cache/cache[4][70] ,
         \I_cache/cache[4][71] , \I_cache/cache[4][72] ,
         \I_cache/cache[4][73] , \I_cache/cache[4][74] ,
         \I_cache/cache[4][75] , \I_cache/cache[4][76] ,
         \I_cache/cache[4][77] , \I_cache/cache[4][78] ,
         \I_cache/cache[4][79] , \I_cache/cache[4][80] ,
         \I_cache/cache[4][81] , \I_cache/cache[4][82] ,
         \I_cache/cache[4][83] , \I_cache/cache[4][84] ,
         \I_cache/cache[4][85] , \I_cache/cache[4][86] ,
         \I_cache/cache[4][87] , \I_cache/cache[4][88] ,
         \I_cache/cache[4][89] , \I_cache/cache[4][90] ,
         \I_cache/cache[4][91] , \I_cache/cache[4][92] ,
         \I_cache/cache[4][93] , \I_cache/cache[4][94] ,
         \I_cache/cache[4][95] , \I_cache/cache[4][96] ,
         \I_cache/cache[4][97] , \I_cache/cache[4][98] ,
         \I_cache/cache[4][99] , \I_cache/cache[4][100] ,
         \I_cache/cache[4][101] , \I_cache/cache[4][102] ,
         \I_cache/cache[4][103] , \I_cache/cache[4][104] ,
         \I_cache/cache[4][105] , \I_cache/cache[4][106] ,
         \I_cache/cache[4][107] , \I_cache/cache[4][108] ,
         \I_cache/cache[4][109] , \I_cache/cache[4][110] ,
         \I_cache/cache[4][111] , \I_cache/cache[4][112] ,
         \I_cache/cache[4][113] , \I_cache/cache[4][114] ,
         \I_cache/cache[4][115] , \I_cache/cache[4][116] ,
         \I_cache/cache[4][117] , \I_cache/cache[4][118] ,
         \I_cache/cache[4][119] , \I_cache/cache[4][120] ,
         \I_cache/cache[4][121] , \I_cache/cache[4][122] ,
         \I_cache/cache[4][123] , \I_cache/cache[4][124] ,
         \I_cache/cache[4][125] , \I_cache/cache[4][126] ,
         \I_cache/cache[4][127] , \I_cache/cache[4][128] ,
         \I_cache/cache[4][129] , \I_cache/cache[4][130] ,
         \I_cache/cache[4][131] , \I_cache/cache[4][132] ,
         \I_cache/cache[4][133] , \I_cache/cache[4][134] ,
         \I_cache/cache[4][135] , \I_cache/cache[4][136] ,
         \I_cache/cache[4][137] , \I_cache/cache[4][138] ,
         \I_cache/cache[4][139] , \I_cache/cache[4][140] ,
         \I_cache/cache[4][141] , \I_cache/cache[4][142] ,
         \I_cache/cache[4][143] , \I_cache/cache[4][144] ,
         \I_cache/cache[4][145] , \I_cache/cache[4][146] ,
         \I_cache/cache[4][147] , \I_cache/cache[4][148] ,
         \I_cache/cache[4][149] , \I_cache/cache[4][150] ,
         \I_cache/cache[4][151] , \I_cache/cache[4][152] ,
         \I_cache/cache[4][153] , \I_cache/cache[4][154] ,
         \I_cache/cache[3][0] , \I_cache/cache[3][1] , \I_cache/cache[3][2] ,
         \I_cache/cache[3][3] , \I_cache/cache[3][4] , \I_cache/cache[3][5] ,
         \I_cache/cache[3][6] , \I_cache/cache[3][7] , \I_cache/cache[3][8] ,
         \I_cache/cache[3][9] , \I_cache/cache[3][10] , \I_cache/cache[3][11] ,
         \I_cache/cache[3][12] , \I_cache/cache[3][13] ,
         \I_cache/cache[3][14] , \I_cache/cache[3][15] ,
         \I_cache/cache[3][16] , \I_cache/cache[3][17] ,
         \I_cache/cache[3][18] , \I_cache/cache[3][19] ,
         \I_cache/cache[3][20] , \I_cache/cache[3][21] ,
         \I_cache/cache[3][22] , \I_cache/cache[3][23] ,
         \I_cache/cache[3][24] , \I_cache/cache[3][25] ,
         \I_cache/cache[3][26] , \I_cache/cache[3][27] ,
         \I_cache/cache[3][28] , \I_cache/cache[3][29] ,
         \I_cache/cache[3][30] , \I_cache/cache[3][31] ,
         \I_cache/cache[3][32] , \I_cache/cache[3][33] ,
         \I_cache/cache[3][34] , \I_cache/cache[3][35] ,
         \I_cache/cache[3][36] , \I_cache/cache[3][37] ,
         \I_cache/cache[3][38] , \I_cache/cache[3][39] ,
         \I_cache/cache[3][40] , \I_cache/cache[3][41] ,
         \I_cache/cache[3][42] , \I_cache/cache[3][43] ,
         \I_cache/cache[3][44] , \I_cache/cache[3][45] ,
         \I_cache/cache[3][46] , \I_cache/cache[3][47] ,
         \I_cache/cache[3][48] , \I_cache/cache[3][49] ,
         \I_cache/cache[3][50] , \I_cache/cache[3][51] ,
         \I_cache/cache[3][52] , \I_cache/cache[3][53] ,
         \I_cache/cache[3][54] , \I_cache/cache[3][55] ,
         \I_cache/cache[3][56] , \I_cache/cache[3][57] ,
         \I_cache/cache[3][58] , \I_cache/cache[3][59] ,
         \I_cache/cache[3][60] , \I_cache/cache[3][61] ,
         \I_cache/cache[3][62] , \I_cache/cache[3][63] ,
         \I_cache/cache[3][64] , \I_cache/cache[3][65] ,
         \I_cache/cache[3][66] , \I_cache/cache[3][67] ,
         \I_cache/cache[3][68] , \I_cache/cache[3][69] ,
         \I_cache/cache[3][70] , \I_cache/cache[3][71] ,
         \I_cache/cache[3][72] , \I_cache/cache[3][73] ,
         \I_cache/cache[3][74] , \I_cache/cache[3][75] ,
         \I_cache/cache[3][76] , \I_cache/cache[3][77] ,
         \I_cache/cache[3][78] , \I_cache/cache[3][79] ,
         \I_cache/cache[3][80] , \I_cache/cache[3][81] ,
         \I_cache/cache[3][82] , \I_cache/cache[3][83] ,
         \I_cache/cache[3][84] , \I_cache/cache[3][85] ,
         \I_cache/cache[3][86] , \I_cache/cache[3][87] ,
         \I_cache/cache[3][88] , \I_cache/cache[3][89] ,
         \I_cache/cache[3][90] , \I_cache/cache[3][91] ,
         \I_cache/cache[3][92] , \I_cache/cache[3][93] ,
         \I_cache/cache[3][94] , \I_cache/cache[3][95] ,
         \I_cache/cache[3][96] , \I_cache/cache[3][97] ,
         \I_cache/cache[3][98] , \I_cache/cache[3][99] ,
         \I_cache/cache[3][100] , \I_cache/cache[3][101] ,
         \I_cache/cache[3][102] , \I_cache/cache[3][103] ,
         \I_cache/cache[3][104] , \I_cache/cache[3][105] ,
         \I_cache/cache[3][106] , \I_cache/cache[3][107] ,
         \I_cache/cache[3][108] , \I_cache/cache[3][109] ,
         \I_cache/cache[3][110] , \I_cache/cache[3][111] ,
         \I_cache/cache[3][112] , \I_cache/cache[3][113] ,
         \I_cache/cache[3][114] , \I_cache/cache[3][115] ,
         \I_cache/cache[3][116] , \I_cache/cache[3][117] ,
         \I_cache/cache[3][118] , \I_cache/cache[3][119] ,
         \I_cache/cache[3][120] , \I_cache/cache[3][121] ,
         \I_cache/cache[3][122] , \I_cache/cache[3][123] ,
         \I_cache/cache[3][124] , \I_cache/cache[3][125] ,
         \I_cache/cache[3][126] , \I_cache/cache[3][127] ,
         \I_cache/cache[3][128] , \I_cache/cache[3][129] ,
         \I_cache/cache[3][130] , \I_cache/cache[3][131] ,
         \I_cache/cache[3][132] , \I_cache/cache[3][133] ,
         \I_cache/cache[3][134] , \I_cache/cache[3][135] ,
         \I_cache/cache[3][136] , \I_cache/cache[3][137] ,
         \I_cache/cache[3][138] , \I_cache/cache[3][139] ,
         \I_cache/cache[3][140] , \I_cache/cache[3][141] ,
         \I_cache/cache[3][142] , \I_cache/cache[3][143] ,
         \I_cache/cache[3][144] , \I_cache/cache[3][145] ,
         \I_cache/cache[3][146] , \I_cache/cache[3][147] ,
         \I_cache/cache[3][148] , \I_cache/cache[3][149] ,
         \I_cache/cache[3][150] , \I_cache/cache[3][151] ,
         \I_cache/cache[3][152] , \I_cache/cache[3][153] ,
         \I_cache/cache[3][154] , \I_cache/cache[2][0] , \I_cache/cache[2][1] ,
         \I_cache/cache[2][2] , \I_cache/cache[2][3] , \I_cache/cache[2][4] ,
         \I_cache/cache[2][5] , \I_cache/cache[2][6] , \I_cache/cache[2][7] ,
         \I_cache/cache[2][8] , \I_cache/cache[2][9] , \I_cache/cache[2][10] ,
         \I_cache/cache[2][11] , \I_cache/cache[2][12] ,
         \I_cache/cache[2][13] , \I_cache/cache[2][14] ,
         \I_cache/cache[2][15] , \I_cache/cache[2][16] ,
         \I_cache/cache[2][17] , \I_cache/cache[2][18] ,
         \I_cache/cache[2][19] , \I_cache/cache[2][20] ,
         \I_cache/cache[2][21] , \I_cache/cache[2][22] ,
         \I_cache/cache[2][23] , \I_cache/cache[2][24] ,
         \I_cache/cache[2][25] , \I_cache/cache[2][26] ,
         \I_cache/cache[2][27] , \I_cache/cache[2][28] ,
         \I_cache/cache[2][29] , \I_cache/cache[2][30] ,
         \I_cache/cache[2][31] , \I_cache/cache[2][32] ,
         \I_cache/cache[2][33] , \I_cache/cache[2][34] ,
         \I_cache/cache[2][35] , \I_cache/cache[2][36] ,
         \I_cache/cache[2][37] , \I_cache/cache[2][38] ,
         \I_cache/cache[2][39] , \I_cache/cache[2][40] ,
         \I_cache/cache[2][41] , \I_cache/cache[2][42] ,
         \I_cache/cache[2][43] , \I_cache/cache[2][44] ,
         \I_cache/cache[2][45] , \I_cache/cache[2][46] ,
         \I_cache/cache[2][47] , \I_cache/cache[2][48] ,
         \I_cache/cache[2][49] , \I_cache/cache[2][50] ,
         \I_cache/cache[2][51] , \I_cache/cache[2][52] ,
         \I_cache/cache[2][53] , \I_cache/cache[2][54] ,
         \I_cache/cache[2][55] , \I_cache/cache[2][56] ,
         \I_cache/cache[2][57] , \I_cache/cache[2][58] ,
         \I_cache/cache[2][59] , \I_cache/cache[2][60] ,
         \I_cache/cache[2][61] , \I_cache/cache[2][62] ,
         \I_cache/cache[2][63] , \I_cache/cache[2][64] ,
         \I_cache/cache[2][65] , \I_cache/cache[2][66] ,
         \I_cache/cache[2][67] , \I_cache/cache[2][68] ,
         \I_cache/cache[2][69] , \I_cache/cache[2][70] ,
         \I_cache/cache[2][71] , \I_cache/cache[2][72] ,
         \I_cache/cache[2][73] , \I_cache/cache[2][74] ,
         \I_cache/cache[2][75] , \I_cache/cache[2][76] ,
         \I_cache/cache[2][77] , \I_cache/cache[2][78] ,
         \I_cache/cache[2][79] , \I_cache/cache[2][80] ,
         \I_cache/cache[2][81] , \I_cache/cache[2][82] ,
         \I_cache/cache[2][83] , \I_cache/cache[2][84] ,
         \I_cache/cache[2][85] , \I_cache/cache[2][86] ,
         \I_cache/cache[2][87] , \I_cache/cache[2][88] ,
         \I_cache/cache[2][89] , \I_cache/cache[2][90] ,
         \I_cache/cache[2][91] , \I_cache/cache[2][92] ,
         \I_cache/cache[2][93] , \I_cache/cache[2][94] ,
         \I_cache/cache[2][95] , \I_cache/cache[2][96] ,
         \I_cache/cache[2][97] , \I_cache/cache[2][98] ,
         \I_cache/cache[2][99] , \I_cache/cache[2][100] ,
         \I_cache/cache[2][101] , \I_cache/cache[2][102] ,
         \I_cache/cache[2][103] , \I_cache/cache[2][104] ,
         \I_cache/cache[2][105] , \I_cache/cache[2][106] ,
         \I_cache/cache[2][107] , \I_cache/cache[2][108] ,
         \I_cache/cache[2][109] , \I_cache/cache[2][110] ,
         \I_cache/cache[2][111] , \I_cache/cache[2][112] ,
         \I_cache/cache[2][113] , \I_cache/cache[2][114] ,
         \I_cache/cache[2][115] , \I_cache/cache[2][116] ,
         \I_cache/cache[2][117] , \I_cache/cache[2][118] ,
         \I_cache/cache[2][119] , \I_cache/cache[2][120] ,
         \I_cache/cache[2][121] , \I_cache/cache[2][122] ,
         \I_cache/cache[2][123] , \I_cache/cache[2][124] ,
         \I_cache/cache[2][125] , \I_cache/cache[2][126] ,
         \I_cache/cache[2][127] , \I_cache/cache[2][128] ,
         \I_cache/cache[2][129] , \I_cache/cache[2][130] ,
         \I_cache/cache[2][131] , \I_cache/cache[2][132] ,
         \I_cache/cache[2][133] , \I_cache/cache[2][134] ,
         \I_cache/cache[2][135] , \I_cache/cache[2][136] ,
         \I_cache/cache[2][137] , \I_cache/cache[2][138] ,
         \I_cache/cache[2][139] , \I_cache/cache[2][140] ,
         \I_cache/cache[2][141] , \I_cache/cache[2][142] ,
         \I_cache/cache[2][143] , \I_cache/cache[2][144] ,
         \I_cache/cache[2][145] , \I_cache/cache[2][146] ,
         \I_cache/cache[2][147] , \I_cache/cache[2][148] ,
         \I_cache/cache[2][149] , \I_cache/cache[2][150] ,
         \I_cache/cache[2][151] , \I_cache/cache[2][152] ,
         \I_cache/cache[2][153] , \I_cache/cache[2][154] ,
         \I_cache/cache[1][0] , \I_cache/cache[1][1] , \I_cache/cache[1][2] ,
         \I_cache/cache[1][3] , \I_cache/cache[1][4] , \I_cache/cache[1][5] ,
         \I_cache/cache[1][6] , \I_cache/cache[1][7] , \I_cache/cache[1][8] ,
         \I_cache/cache[1][9] , \I_cache/cache[1][10] , \I_cache/cache[1][11] ,
         \I_cache/cache[1][12] , \I_cache/cache[1][13] ,
         \I_cache/cache[1][14] , \I_cache/cache[1][15] ,
         \I_cache/cache[1][16] , \I_cache/cache[1][17] ,
         \I_cache/cache[1][18] , \I_cache/cache[1][19] ,
         \I_cache/cache[1][20] , \I_cache/cache[1][21] ,
         \I_cache/cache[1][22] , \I_cache/cache[1][23] ,
         \I_cache/cache[1][24] , \I_cache/cache[1][25] ,
         \I_cache/cache[1][26] , \I_cache/cache[1][27] ,
         \I_cache/cache[1][28] , \I_cache/cache[1][29] ,
         \I_cache/cache[1][30] , \I_cache/cache[1][31] ,
         \I_cache/cache[1][32] , \I_cache/cache[1][33] ,
         \I_cache/cache[1][34] , \I_cache/cache[1][35] ,
         \I_cache/cache[1][36] , \I_cache/cache[1][37] ,
         \I_cache/cache[1][38] , \I_cache/cache[1][39] ,
         \I_cache/cache[1][40] , \I_cache/cache[1][41] ,
         \I_cache/cache[1][42] , \I_cache/cache[1][43] ,
         \I_cache/cache[1][44] , \I_cache/cache[1][45] ,
         \I_cache/cache[1][46] , \I_cache/cache[1][47] ,
         \I_cache/cache[1][48] , \I_cache/cache[1][49] ,
         \I_cache/cache[1][50] , \I_cache/cache[1][51] ,
         \I_cache/cache[1][52] , \I_cache/cache[1][53] ,
         \I_cache/cache[1][54] , \I_cache/cache[1][55] ,
         \I_cache/cache[1][56] , \I_cache/cache[1][57] ,
         \I_cache/cache[1][58] , \I_cache/cache[1][59] ,
         \I_cache/cache[1][60] , \I_cache/cache[1][61] ,
         \I_cache/cache[1][62] , \I_cache/cache[1][63] ,
         \I_cache/cache[1][64] , \I_cache/cache[1][65] ,
         \I_cache/cache[1][66] , \I_cache/cache[1][67] ,
         \I_cache/cache[1][68] , \I_cache/cache[1][69] ,
         \I_cache/cache[1][70] , \I_cache/cache[1][71] ,
         \I_cache/cache[1][72] , \I_cache/cache[1][73] ,
         \I_cache/cache[1][74] , \I_cache/cache[1][75] ,
         \I_cache/cache[1][76] , \I_cache/cache[1][77] ,
         \I_cache/cache[1][78] , \I_cache/cache[1][79] ,
         \I_cache/cache[1][80] , \I_cache/cache[1][81] ,
         \I_cache/cache[1][82] , \I_cache/cache[1][83] ,
         \I_cache/cache[1][84] , \I_cache/cache[1][85] ,
         \I_cache/cache[1][86] , \I_cache/cache[1][87] ,
         \I_cache/cache[1][88] , \I_cache/cache[1][89] ,
         \I_cache/cache[1][90] , \I_cache/cache[1][91] ,
         \I_cache/cache[1][92] , \I_cache/cache[1][93] ,
         \I_cache/cache[1][94] , \I_cache/cache[1][95] ,
         \I_cache/cache[1][96] , \I_cache/cache[1][97] ,
         \I_cache/cache[1][98] , \I_cache/cache[1][99] ,
         \I_cache/cache[1][100] , \I_cache/cache[1][101] ,
         \I_cache/cache[1][102] , \I_cache/cache[1][103] ,
         \I_cache/cache[1][104] , \I_cache/cache[1][105] ,
         \I_cache/cache[1][106] , \I_cache/cache[1][107] ,
         \I_cache/cache[1][108] , \I_cache/cache[1][109] ,
         \I_cache/cache[1][110] , \I_cache/cache[1][111] ,
         \I_cache/cache[1][112] , \I_cache/cache[1][113] ,
         \I_cache/cache[1][114] , \I_cache/cache[1][115] ,
         \I_cache/cache[1][116] , \I_cache/cache[1][117] ,
         \I_cache/cache[1][118] , \I_cache/cache[1][119] ,
         \I_cache/cache[1][120] , \I_cache/cache[1][121] ,
         \I_cache/cache[1][122] , \I_cache/cache[1][123] ,
         \I_cache/cache[1][124] , \I_cache/cache[1][125] ,
         \I_cache/cache[1][126] , \I_cache/cache[1][127] ,
         \I_cache/cache[1][128] , \I_cache/cache[1][129] ,
         \I_cache/cache[1][130] , \I_cache/cache[1][131] ,
         \I_cache/cache[1][132] , \I_cache/cache[1][133] ,
         \I_cache/cache[1][134] , \I_cache/cache[1][135] ,
         \I_cache/cache[1][136] , \I_cache/cache[1][137] ,
         \I_cache/cache[1][138] , \I_cache/cache[1][139] ,
         \I_cache/cache[1][140] , \I_cache/cache[1][141] ,
         \I_cache/cache[1][142] , \I_cache/cache[1][143] ,
         \I_cache/cache[1][144] , \I_cache/cache[1][145] ,
         \I_cache/cache[1][146] , \I_cache/cache[1][147] ,
         \I_cache/cache[1][148] , \I_cache/cache[1][149] ,
         \I_cache/cache[1][150] , \I_cache/cache[1][151] ,
         \I_cache/cache[1][152] , \I_cache/cache[1][153] ,
         \I_cache/cache[1][154] , \I_cache/cache[0][0] , \I_cache/cache[0][1] ,
         \I_cache/cache[0][2] , \I_cache/cache[0][3] , \I_cache/cache[0][4] ,
         \I_cache/cache[0][5] , \I_cache/cache[0][6] , \I_cache/cache[0][7] ,
         \I_cache/cache[0][8] , \I_cache/cache[0][9] , \I_cache/cache[0][10] ,
         \I_cache/cache[0][11] , \I_cache/cache[0][12] ,
         \I_cache/cache[0][13] , \I_cache/cache[0][14] ,
         \I_cache/cache[0][15] , \I_cache/cache[0][16] ,
         \I_cache/cache[0][17] , \I_cache/cache[0][18] ,
         \I_cache/cache[0][19] , \I_cache/cache[0][20] ,
         \I_cache/cache[0][21] , \I_cache/cache[0][22] ,
         \I_cache/cache[0][23] , \I_cache/cache[0][24] ,
         \I_cache/cache[0][25] , \I_cache/cache[0][26] ,
         \I_cache/cache[0][27] , \I_cache/cache[0][28] ,
         \I_cache/cache[0][29] , \I_cache/cache[0][30] ,
         \I_cache/cache[0][31] , \I_cache/cache[0][32] ,
         \I_cache/cache[0][33] , \I_cache/cache[0][34] ,
         \I_cache/cache[0][35] , \I_cache/cache[0][36] ,
         \I_cache/cache[0][37] , \I_cache/cache[0][38] ,
         \I_cache/cache[0][39] , \I_cache/cache[0][40] ,
         \I_cache/cache[0][41] , \I_cache/cache[0][42] ,
         \I_cache/cache[0][43] , \I_cache/cache[0][44] ,
         \I_cache/cache[0][45] , \I_cache/cache[0][46] ,
         \I_cache/cache[0][47] , \I_cache/cache[0][48] ,
         \I_cache/cache[0][49] , \I_cache/cache[0][50] ,
         \I_cache/cache[0][51] , \I_cache/cache[0][52] ,
         \I_cache/cache[0][53] , \I_cache/cache[0][54] ,
         \I_cache/cache[0][55] , \I_cache/cache[0][56] ,
         \I_cache/cache[0][57] , \I_cache/cache[0][58] ,
         \I_cache/cache[0][59] , \I_cache/cache[0][60] ,
         \I_cache/cache[0][61] , \I_cache/cache[0][62] ,
         \I_cache/cache[0][63] , \I_cache/cache[0][64] ,
         \I_cache/cache[0][65] , \I_cache/cache[0][66] ,
         \I_cache/cache[0][67] , \I_cache/cache[0][68] ,
         \I_cache/cache[0][69] , \I_cache/cache[0][70] ,
         \I_cache/cache[0][71] , \I_cache/cache[0][72] ,
         \I_cache/cache[0][73] , \I_cache/cache[0][74] ,
         \I_cache/cache[0][75] , \I_cache/cache[0][76] ,
         \I_cache/cache[0][77] , \I_cache/cache[0][78] ,
         \I_cache/cache[0][79] , \I_cache/cache[0][80] ,
         \I_cache/cache[0][81] , \I_cache/cache[0][82] ,
         \I_cache/cache[0][83] , \I_cache/cache[0][84] ,
         \I_cache/cache[0][85] , \I_cache/cache[0][86] ,
         \I_cache/cache[0][87] , \I_cache/cache[0][88] ,
         \I_cache/cache[0][89] , \I_cache/cache[0][90] ,
         \I_cache/cache[0][91] , \I_cache/cache[0][92] ,
         \I_cache/cache[0][93] , \I_cache/cache[0][94] ,
         \I_cache/cache[0][95] , \I_cache/cache[0][96] ,
         \I_cache/cache[0][97] , \I_cache/cache[0][98] ,
         \I_cache/cache[0][99] , \I_cache/cache[0][100] ,
         \I_cache/cache[0][101] , \I_cache/cache[0][102] ,
         \I_cache/cache[0][103] , \I_cache/cache[0][104] ,
         \I_cache/cache[0][105] , \I_cache/cache[0][106] ,
         \I_cache/cache[0][107] , \I_cache/cache[0][108] ,
         \I_cache/cache[0][109] , \I_cache/cache[0][110] ,
         \I_cache/cache[0][111] , \I_cache/cache[0][112] ,
         \I_cache/cache[0][113] , \I_cache/cache[0][114] ,
         \I_cache/cache[0][115] , \I_cache/cache[0][116] ,
         \I_cache/cache[0][117] , \I_cache/cache[0][118] ,
         \I_cache/cache[0][119] , \I_cache/cache[0][120] ,
         \I_cache/cache[0][121] , \I_cache/cache[0][122] ,
         \I_cache/cache[0][123] , \I_cache/cache[0][124] ,
         \I_cache/cache[0][125] , \I_cache/cache[0][126] ,
         \I_cache/cache[0][127] , \I_cache/cache[0][128] ,
         \I_cache/cache[0][129] , \I_cache/cache[0][130] ,
         \I_cache/cache[0][131] , \I_cache/cache[0][132] ,
         \I_cache/cache[0][133] , \I_cache/cache[0][134] ,
         \I_cache/cache[0][135] , \I_cache/cache[0][136] ,
         \I_cache/cache[0][137] , \I_cache/cache[0][138] ,
         \I_cache/cache[0][139] , \I_cache/cache[0][140] ,
         \I_cache/cache[0][141] , \I_cache/cache[0][142] ,
         \I_cache/cache[0][143] , \I_cache/cache[0][144] ,
         \I_cache/cache[0][145] , \I_cache/cache[0][146] ,
         \I_cache/cache[0][147] , \I_cache/cache[0][148] ,
         \I_cache/cache[0][149] , \I_cache/cache[0][150] ,
         \I_cache/cache[0][151] , \I_cache/cache[0][152] ,
         \I_cache/cache[0][153] , \I_cache/cache[0][154] , net36572, net36639,
         net49779, net103753, net103785, net103817, net103849, net104166,
         net104168, net104171, net104172, net104173, net104343, net104367,
         net104503, net104691, net104698, net104699, net104700, net104721,
         net104725, net104752, net104754, net104755, net104765, net104791,
         net104792, net104793, net104794, net104801, net104828, net104830,
         net104861, net104866, net104867, net104868, net104884, net104889,
         net104890, net104891, net104905, net104906, net104915, net104916,
         net104917, net104918, net104934, net104939, net104940, net104941,
         net104957, net104962, net104963, net104964, net104980, net104985,
         net105003, net105008, net105009, net105010, net105071, net105075,
         net105076, net105077, net105093, net105105, net105110, net105111,
         net105112, net105119, net105120, net105121, net105137, net105142,
         net105143, net105160, net105165, net105166, net105167, net105179,
         net105195, net105227, net105232, net105233, net105234, net105236,
         net105250, net105255, net105256, net105264, net105265, net105266,
         net105269, net105283, net105288, net105289, net105290, net105311,
         net105312, net105313, net105329, net105334, net105335, net105336,
         net105364, net105375, net105376, net105396, net105412, net105423,
         net105424, net105425, net105430, net105433, net105434, net105435,
         net105436, net105447, net105448, net105449, net105462, net105463,
         net105477, net105479, net105490, net105491, net105492, net105506,
         net105517, net105531, net105549, net105567, net105662, net105663,
         net105731, net105732, net105746, net105751, net105752, net105753,
         net105756, net105764, net105783, net105798, net105820, net105834,
         net105835, net106031, net106037, net106038, net106040, net106041,
         net106290, net106297, net106298, net106301, net106596, net106602,
         net106603, net106674, net106675, net106679, net106680, net106681,
         net106682, net106692, net106693, net106694, net106695, net106705,
         net106706, net106707, net106708, net106718, net106719, net106720,
         net106721, net106819, net106822, net106828, net107119, net107120,
         net107123, net107134, net107135, net107138, net107141, net107167,
         net107168, net107169, net107170, net107195, net107196, net107210,
         net107217, net107218, net107224, net107228, net107230, net107389,
         net107404, net107411, net107517, net107518, net107519, net107606,
         net107607, net107615, net107617, net107619, net107621, net107652,
         net107656, net107657, net107659, net107661, net107665, net107680,
         net107688, net107689, net107696, net107828, net107841, net107854,
         net107855, net107856, net107857, net107858, net107943, net107977,
         net107987, net107988, net107991, net107992, net108003, net108004,
         net108005, net108010, net108012, net108101, net108148, net108149,
         net108150, net108151, net108160, net108161, net108162, net108249,
         net108281, net108284, net108285, net108290, net108297, net108299,
         net108300, net108306, net108308, net108310, net108323, net108412,
         net108490, net108491, net108492, net108579, net108622, net108623,
         net108624, net108625, net108631, net108632, net108640, net108641,
         net108642, net108729, net108779, net108781, net108787, net108846,
         net108847, net108851, net108852, net108853, net108854, net108868,
         net108869, net108873, net108874, net108876, net108893, net108894,
         net108895, net109040, net109042, net109129, net109168, net109172,
         net109176, net109179, net109196, net109201, net109202, net109203,
         net109359, net109360, net109447, net109496, net109510, net109511,
         net109512, net109513, net109519, net109527, net109528, net109529,
         net109616, net109661, net109666, net109673, net109674, net109675,
         net109762, net109839, net109840, net109841, net109965, net109989,
         net109990, net109991, net110129, net110131, net110147, net110227,
         net110406, net110423, net110424, net110429, net110470, net110473,
         net110569, net110602, net110640, net110642, net110729, net110798,
         net110799, net110800, net110928, net110932, net110953, net110954,
         net110955, net111041, net111128, net111129, net111130, net111216,
         net111249, net111256, net111262, net111276, net111277, net111278,
         net111364, net111413, net111416, net111421, net111422, net111423,
         net111509, net111572, net111580, net111581, net111582, net111710,
         net111723, net111724, net111762, net111763, net111764, net111930,
         net111931, net111932, net112118, net112119, net112120, net112214,
         net112219, net112328, net112329, net112330, net112392, net112393,
         net112410, net112414, net112417, net112418, net112425, net112446,
         net112449, net112512, net112534, net112544, net112549, net112555,
         net112585, net112586, net114073, net114065, net114081, net114079,
         net114087, net114085, net114341, net114331, net114325, net114319,
         net115799, net115797, net115795, net115793, net115791, net115789,
         net115813, net115811, net117631, net117625, net117623, net117643,
         net117641, net117639, net117637, net117635, net117647, net117667,
         net117665, net117663, net117661, net117659, net117657, net117655,
         net117653, net117681, net117675, net117673, net117685, net117683,
         net117697, net117695, net117691, net117703, net117719, net117715,
         net117713, net117711, net117709, net117727, net117723, net117741,
         net117733, net117731, net117747, net117745, net117743, net117751,
         net117759, net117757, net118217, net118215, net118223, net118227,
         net118225, net118239, net118237, net118235, net118233, net118243,
         net118241, net118255, net118253, net118263, net118261, net118259,
         net118275, net118273, net118271, net118269, net118267, net118281,
         net118291, net118289, net118297, net118295, net118321, net118319,
         net118315, net118313, net118311, net118307, net118305, net118303,
         net118347, net118345, net118343, net118341, net118339, net118337,
         net118335, net118331, net118329, net118327, net118369, net118367,
         net118365, net118359, net118357, net118355, net118353, net118351,
         net118395, net118381, net118379, net118375, net118417, net118415,
         net118413, net118409, net118407, net118405, net118403, net118401,
         net118399, net118441, net118439, net118431, net118429, net118425,
         net118423, net118467, net118457, net118455, net118453, net118451,
         net118491, net118487, net118483, net118481, net118479, net118477,
         net118475, net118473, net118581, net118584, net118592, net118597,
         net118601, net118926, net118925, net119021, net119020, net119018,
         net119104, net119263, net134069, net134375, net134414, net134445,
         net134673, net134679, net134680, net134681, net134682, net134683,
         net134684, net134685, net134686, net134710, net134815, net134876,
         net134907, net135423, net135522, net135551, net135772, net139718,
         net139719, net139756, net139765, net139774, net139775, net139776,
         net139777, net139778, net139810, net139838, net139849, net139850,
         net139859, net139860, net139862, net139863, net139864, net139865,
         net139866, net140147, net143504, net143503, net143507, net143506,
         net143514, net143513, net143525, net143524, net143548, net143547,
         net143556, net143555, net143858, net143857, net144187, net144227,
         net144224, net144236, net144667, net144666, net111716, net111668,
         net105582, net105581, net105257, net112413, net111270, net110430,
         net109668, net134145, net111570, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24,
         n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n170, n171, n172,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193, n194,
         n195, n196, n197, n198, n199, n200, n201, n202, n203, n204, n205,
         n206, n207, n208, n209, n210, n211, n212, n213, n214, n215, n216,
         n217, n218, n219, n220, n221, n222, n223, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n242, n243, n244, n245, n246, n247, n248, n249,
         n250, n251, n252, n253, n254, n255, n256, n257, n258, n259, n260,
         n261, n262, n263, n264, n265, n266, n267, n268, n269, n270, n271,
         n272, n273, n274, n275, n276, n277, n278, n279, n280, n281, n282,
         n283, n284, n285, n286, n287, n288, n289, n290, n291, n292, n293,
         n294, n295, n296, n297, n298, n299, n300, n301, n302, n303, n304,
         n305, n306, n307, n308, n309, n310, n311, n312, n313, n314, n315,
         n316, n317, n318, n319, n320, n321, n322, n323, n324, n325, n326,
         n327, n328, n329, n330, n331, n332, n333, n334, n335, n336, n337,
         n338, n339, n340, n341, n342, n343, n344, n345, n346, n347, n348,
         n349, n350, n351, n352, n353, n354, n355, n356, n357, n358, n359,
         n360, n361, n362, n363, n364, n365, n366, n367, n368, n369, n370,
         n371, n372, n373, n374, n375, n376, n377, n378, n379, n380, n381,
         n382, n383, n384, n385, n386, n387, n388, n389, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007,
         n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017,
         n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027,
         n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037,
         n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047,
         n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057,
         n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067,
         n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077,
         n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087,
         n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097,
         n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107,
         n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117,
         n1118, n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127,
         n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137,
         n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147,
         n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157,
         n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167,
         n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177,
         n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187,
         n1188, n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247,
         n1248, n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257,
         n1258, n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267,
         n1268, n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277,
         n1278, n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287,
         n1288, n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297,
         n1298, n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307,
         n1308, n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317,
         n1318, n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327,
         n1328, n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337,
         n1338, n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347,
         n1348, n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357,
         n1358, n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367,
         n1368, n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377,
         n1378, n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387,
         n1388, n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397,
         n1398, n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407,
         n1408, n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417,
         n1418, n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427,
         n1428, n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437,
         n1438, n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447,
         n1448, n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457,
         n1458, n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467,
         n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477,
         n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487,
         n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497,
         n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507,
         n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517,
         n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527,
         n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537,
         n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547,
         n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557,
         n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567,
         n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577,
         n1578, n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587,
         n1588, n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597,
         n1598, n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607,
         n1608, n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617,
         n1618, n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627,
         n1628, n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637,
         n1638, n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647,
         n1648, n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657,
         n1658, n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667,
         n1668, n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677,
         n1678, n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687,
         n1688, n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697,
         n1698, n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707,
         n1708, n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717,
         n1718, n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727,
         n1728, n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737,
         n1738, n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747,
         n1748, n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757,
         n1758, n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767,
         n1768, n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777,
         n1778, n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787,
         n1788, n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797,
         n1798, n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807,
         n1808, n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817,
         n1818, n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827,
         n1828, n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837,
         n1838, n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847,
         n1848, n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857,
         n1858, n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867,
         n1868, n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877,
         n1878, n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887,
         n1888, n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897,
         n1898, n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907,
         n1908, n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917,
         n1918, n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927,
         n1928, n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937,
         n1938, n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947,
         n1948, n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957,
         n1958, n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967,
         n1968, n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977,
         n1978, n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987,
         n1988, n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997,
         n1998, n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007,
         n2008, n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017,
         n2018, n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027,
         n2028, n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037,
         n2038, n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047,
         n2048, n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057,
         n2058, n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067,
         n2068, n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077,
         n2078, n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087,
         n2088, n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097,
         n2098, n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107,
         n2108, n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117,
         n2118, n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127,
         n2128, n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137,
         n2138, n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147,
         n2148, n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157,
         n2158, n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167,
         n2168, n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177,
         n2178, n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187,
         n2188, n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197,
         n2198, n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207,
         n2208, n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217,
         n2218, n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227,
         n2228, n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237,
         n2238, n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247,
         n2248, n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257,
         n2258, n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267,
         n2268, n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277,
         n2278, n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287,
         n2288, n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297,
         n2298, n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307,
         n2308, n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317,
         n2318, n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327,
         n2328, n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337,
         n2338, n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347,
         n2348, n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357,
         n2358, n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367,
         n2368, n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377,
         n2378, n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387,
         n2388, n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397,
         n2398, n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407,
         n2408, n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417,
         n2418, n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427,
         n2428, n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437,
         n2438, n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447,
         n2448, n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457,
         n2458, n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467,
         n2468, n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477,
         n2478, n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487,
         n2488, n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497,
         n2498, n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507,
         n2508, n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517,
         n2518, n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527,
         n2528, n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537,
         n2538, n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547,
         n2548, n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557,
         n2558, n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567,
         n2568, n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577,
         n2578, n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587,
         n2588, n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597,
         n2598, n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607,
         n2608, n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617,
         n2618, n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627,
         n2628, n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637,
         n2638, n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647,
         n2648, n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657,
         n2658, n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667,
         n2668, n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677,
         n2678, n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687,
         n2688, n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697,
         n2698, n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707,
         n2708, n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717,
         n2718, n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727,
         n2728, n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737,
         n2738, n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747,
         n2748, n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757,
         n2758, n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767,
         n2768, n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777,
         n2778, n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787,
         n2788, n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797,
         n2798, n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807,
         n2808, n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817,
         n2818, n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827,
         n2828, n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837,
         n2838, n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847,
         n2848, n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857,
         n2858, n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867,
         n2868, n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877,
         n2878, n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887,
         n2888, n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897,
         n2898, n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907,
         n2908, n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917,
         n2918, n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927,
         n2928, n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937,
         n2938, n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947,
         n2948, n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957,
         n2958, n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967,
         n2968, n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977,
         n2978, n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987,
         n2988, n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997,
         n2998, n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007,
         n3008, n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017,
         n3018, n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027,
         n3028, n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037,
         n3038, n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047,
         n3048, n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057,
         n3058, n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067,
         n3068, n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077,
         n3078, n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087,
         n3088, n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097,
         n3098, n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107,
         n3108, n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117,
         n3118, n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127,
         n3128, n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137,
         n3138, n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147,
         n3148, n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157,
         n3158, n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167,
         n3168, n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177,
         n3178, n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187,
         n3188, n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197,
         n3198, n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207,
         n3208, n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217,
         n3218, n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227,
         n3228, n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237,
         n3238, n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247,
         n3248, n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257,
         n3258, n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267,
         n3268, n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277,
         n3278, n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287,
         n3288, n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297,
         n3298, n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307,
         n3308, n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317,
         n3318, n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327,
         n3328, n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337,
         n3338, n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347,
         n3348, n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357,
         n3358, n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367,
         n3368, n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377,
         n3378, n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387,
         n3388, n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397,
         n3398, n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407,
         n3408, n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417,
         n3418, n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427,
         n3428, n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437,
         n3438, n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447,
         n3448, n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457,
         n3458, n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467,
         n3468, n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477,
         n3478, n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487,
         n3488, n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497,
         n3498, n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507,
         n3508, n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517,
         n3518, n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527,
         n3528, n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537,
         n3538, n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547,
         n3548, n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557,
         n3558, n3559, n3560, n3561, n3562, n3564, n3565, n3567, n3569, n3574,
         n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583, n3584,
         n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593, n3594,
         n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603, n3604,
         n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613, n3614,
         n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623, n3624,
         n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633, n3634,
         n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643, n3644,
         n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653, n3654,
         n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663, n3664,
         n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673, n3674,
         n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683, n3684,
         n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693, n3694,
         n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703, n3704,
         n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713, n3714,
         n3715, n3716, n3717, n3718, n3719, n3720, n3723, n3724, n3725, n3726,
         n3727, n3728, n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736,
         n3737, n3738, n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746,
         n3747, n3748, n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756,
         n3757, n3758, n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766,
         n3767, n3768, n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776,
         n3777, n3778, n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786,
         n3787, n3788, n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796,
         n3797, n3798, n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806,
         n3807, n3808, n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816,
         n3817, n3818, n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826,
         n3827, n3828, n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836,
         n3837, n3838, n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846,
         n3847, n3848, n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856,
         n3857, n3858, n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866,
         n3867, n3868, n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876,
         n3877, n3878, n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886,
         n3887, n3888, n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896,
         n3897, n3898, n3900, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3944, n3945, n3946, n3947, n3948, n3949,
         n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959,
         n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969,
         n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979,
         n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989,
         n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999,
         n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4053, n4054, n4055, n4056, n4057, n4059, n4060, n4064, n4065, n4066,
         n4067, n4068, n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076,
         n4077, n4078, n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086,
         n4087, n4088, n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096,
         n4097, n4098, n4099, n4100, n4101, n4103, n4105, n4106, n4107, n4109,
         n4111, n4113, n4115, n4117, n4119, n4121, n4123, n4125, n4127, n4129,
         n4131, n4133, n4135, n4137, n4139, n4141, n4143, n4145, n4147, n4149,
         n4151, n4153, n4155, n4157, n4159, n4161, n4163, n4165, n4167, n4169,
         n4171, n4173, n4175, n4177, n4179, n4181, n4183, n4185, n4187, n4189,
         n4191, n4193, n4195, n4197, n4199, n4201, n4203, n4205, n4207, n4209,
         n4211, n4213, n4215, n4217, n4219, n4221, n4223, n4225, n4227, n4229,
         n4231, n4233, n4235, n4237, n4239, n4241, n4243, n4245, n4247, n4249,
         n4251, n4253, n4255, n4257, n4259, n4261, n4263, n4265, n4267, n4269,
         n4271, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4511, n4512, n4513, n4514, n4515, n4516,
         n4517, n4518, n4519, n4520, n4521, n4522, n4523, n4525, n4526, n4527,
         n4528, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4581, n4617,
         n4618, n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627,
         n4628, n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637,
         n4638, n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647,
         n4648, n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657,
         n4658, n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667,
         n4668, n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677,
         n4678, n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687,
         n4688, n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697,
         n4698, n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707,
         n4708, n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717,
         n4718, n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727,
         n4728, n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737,
         n4738, n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747,
         n4748, n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757,
         n4758, n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767,
         n4768, n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777,
         n4778, n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787,
         n4788, n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797,
         n4798, n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807,
         n4808, n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817,
         n4818, n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827,
         n4828, n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837,
         n4838, n4840, n4842, n4844, n4846, n4848, n4850, n4852, n4854, n4856,
         n4858, n4875, n4877, n4882, n4883, n4893, n4902, n4907, n4920, n4922,
         n4929, n4932, n4933, n4935, n4936, n4937, n4938, n4939, n4941, n4943,
         n4944, n4954, n4971, n4973, n4974, n4975, n4976, n4978, n4979, n4980,
         n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990,
         n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000,
         n5001, n5002, n5003, n5004, n5005, n5006, n5008, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5021, n5023, n5024,
         n5026, n5027, n5028, n5031, n5032, n5033, n5035, n5037, n5038, n5039,
         n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049,
         n5050, n5051, n5052, n5053, n5055, n5056, n5057, n5058, n5059, n5060,
         n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070,
         n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080,
         n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090,
         n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100,
         n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110,
         n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120,
         n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130,
         n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140,
         n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150,
         n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160,
         n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170,
         n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180,
         n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190,
         n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200,
         n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210,
         n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220,
         n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230,
         n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240,
         n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250,
         n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260,
         n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270,
         n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280,
         n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290,
         n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300,
         n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310,
         n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320,
         n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330,
         n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340,
         n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350,
         n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360,
         n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370,
         n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380,
         n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390,
         n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400,
         n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410,
         n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420,
         n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430,
         n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440,
         n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450,
         n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460,
         n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470,
         n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480,
         n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490,
         n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500,
         n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510,
         n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520,
         n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530,
         n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540,
         n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550,
         n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560,
         n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570,
         n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580,
         n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590,
         n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600,
         n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610,
         n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620,
         n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630,
         n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640,
         n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650,
         n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660,
         n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670,
         n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680,
         n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690,
         n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700,
         n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710,
         n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720,
         n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730,
         n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740,
         n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750,
         n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760,
         n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770,
         n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780,
         n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790,
         n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800,
         n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810,
         n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820,
         n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830,
         n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840,
         n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850,
         n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860,
         n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870,
         n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880,
         n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890,
         n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900,
         n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910,
         n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920,
         n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930,
         n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940,
         n5941, n5942, n5943, n5944, n5945, n5947, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
         n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
         n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
         n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
         n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
         n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
         n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
         n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
         n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
         n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
         n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
         n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
         n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
         n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
         n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053,
         n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063,
         n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073,
         n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
         n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
         n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
         n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
         n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123,
         n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133,
         n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143,
         n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153,
         n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163,
         n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173,
         n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183,
         n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193,
         n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
         n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
         n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
         n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
         n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
         n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253,
         n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263,
         n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273,
         n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283,
         n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293,
         n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303,
         n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313,
         n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323,
         n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333,
         n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343,
         n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353,
         n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363,
         n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373,
         n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383,
         n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393,
         n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403,
         n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413,
         n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423,
         n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433,
         n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443,
         n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453,
         n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463,
         n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473,
         n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483,
         n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493,
         n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503,
         n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513,
         n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523,
         n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533,
         n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543,
         n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553,
         n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563,
         n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573,
         n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
         n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593,
         n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
         n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613,
         n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623,
         n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633,
         n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643,
         n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653,
         n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663,
         n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673,
         n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683,
         n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693,
         n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703,
         n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713,
         n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723,
         n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733,
         n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743,
         n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753,
         n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763,
         n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773,
         n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783,
         n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793,
         n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803,
         n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813,
         n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823,
         n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833,
         n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843,
         n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853,
         n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863,
         n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873,
         n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883,
         n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893,
         n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903,
         n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913,
         n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923,
         n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933,
         n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943,
         n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953,
         n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963,
         n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973,
         n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983,
         n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993,
         n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003,
         n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013,
         n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023,
         n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033,
         n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043,
         n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053,
         n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063,
         n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073,
         n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083,
         n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093,
         n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103,
         n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113,
         n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123,
         n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133,
         n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143,
         n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153,
         n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163,
         n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173,
         n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183,
         n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193,
         n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203,
         n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213,
         n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223,
         n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233,
         n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243,
         n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253,
         n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263,
         n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273,
         n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283,
         n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293,
         n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303,
         n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313,
         n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323,
         n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333,
         n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343,
         n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353,
         n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363,
         n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373,
         n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383,
         n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393,
         n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403,
         n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413,
         n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423,
         n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433,
         n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443,
         n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453,
         n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463,
         n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473,
         n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483,
         n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493,
         n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503,
         n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513,
         n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523,
         n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533,
         n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543,
         n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553,
         n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563,
         n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573,
         n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583,
         n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593,
         n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603,
         n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613,
         n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623,
         n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633,
         n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643,
         n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653,
         n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663,
         n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673,
         n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683,
         n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693,
         n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703,
         n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713,
         n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723,
         n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733,
         n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743,
         n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753,
         n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763,
         n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773,
         n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783,
         n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793,
         n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803,
         n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813,
         n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823,
         n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833,
         n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843,
         n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853,
         n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863,
         n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873,
         n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883,
         n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893,
         n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903,
         n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913,
         n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923,
         n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933,
         n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943,
         n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953,
         n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963,
         n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973,
         n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983,
         n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993,
         n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003,
         n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013,
         n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023,
         n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033,
         n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043,
         n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053,
         n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063,
         n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073,
         n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083,
         n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093,
         n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103,
         n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113,
         n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123,
         n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133,
         n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143,
         n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153,
         n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163,
         n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173,
         n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183,
         n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193,
         n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203,
         n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213,
         n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223,
         n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233,
         n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243,
         n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253,
         n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263,
         n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273,
         n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283,
         n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293,
         n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303,
         n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313,
         n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323,
         n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333,
         n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343,
         n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353,
         n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363,
         n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373,
         n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383,
         n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393,
         n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403,
         n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413,
         n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423,
         n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433,
         n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443,
         n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453,
         n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463,
         n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473,
         n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483,
         n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493,
         n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503,
         n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513,
         n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523,
         n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533,
         n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543,
         n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553,
         n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563,
         n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573,
         n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583,
         n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593,
         n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603,
         n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613,
         n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623,
         n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633,
         n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643,
         n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653,
         n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663,
         n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673,
         n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683,
         n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693,
         n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703,
         n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713,
         n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723,
         n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733,
         n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743,
         n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753,
         n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763,
         n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773,
         n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783,
         n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793,
         n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803,
         n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813,
         n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823,
         n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
         n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
         n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
         n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
         n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
         n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
         n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
         n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170,
         n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
         n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
         n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
         n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202,
         n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210,
         n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218,
         n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226,
         n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234,
         n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242,
         n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250,
         n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
         n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
         n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274,
         n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
         n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290,
         n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298,
         n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
         n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314,
         n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322,
         n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
         n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338,
         n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346,
         n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354,
         n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362,
         n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370,
         n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378,
         n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386,
         n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
         n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
         n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410,
         n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418,
         n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426,
         n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
         n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442,
         n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
         n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458,
         n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
         n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
         n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482,
         n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,
         n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
         n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506,
         n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514,
         n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522,
         n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530,
         n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538,
         n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546,
         n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554,
         n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562,
         n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570,
         n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578,
         n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586,
         n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594,
         n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602,
         n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610,
         n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618,
         n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626,
         n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634,
         n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642,
         n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650,
         n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658,
         n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666,
         n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674,
         n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682,
         n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690,
         n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698,
         n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706,
         n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714,
         n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722,
         n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730,
         n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738,
         n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746,
         n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754,
         n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762,
         n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770,
         n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778,
         n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786,
         n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794,
         n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802,
         n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810,
         n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818,
         n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826,
         n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834,
         n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842,
         n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850,
         n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858,
         n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866,
         n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874,
         n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882,
         n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890,
         n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898,
         n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906,
         n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914,
         n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922,
         n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930,
         n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938,
         n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946,
         n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954,
         n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962,
         n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970,
         n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978,
         n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986,
         n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994,
         n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002,
         n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010,
         n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018,
         n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026,
         n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034,
         n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042,
         n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050,
         n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058,
         n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066,
         n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074,
         n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082,
         n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090,
         n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098,
         n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106,
         n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114,
         n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122,
         n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130,
         n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138,
         n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146,
         n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154,
         n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162,
         n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170,
         n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178,
         n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186,
         n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194,
         n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202,
         n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210,
         n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218,
         n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226,
         n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234,
         n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242,
         n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250,
         n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258,
         n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266,
         n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274,
         n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282,
         n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290,
         n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298,
         n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306,
         n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314,
         n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322,
         n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330,
         n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338,
         n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346,
         n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354,
         n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362,
         n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370,
         n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378,
         n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386,
         n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394,
         n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402,
         n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410,
         n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418,
         n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426,
         n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434,
         n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442,
         n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450,
         n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458,
         n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466,
         n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474,
         n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482,
         n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490,
         n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498,
         n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506,
         n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514,
         n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522,
         n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530,
         n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538,
         n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546,
         n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554,
         n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562,
         n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570,
         n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578,
         n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586,
         n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594,
         n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602,
         n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610,
         n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618,
         n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626,
         n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634,
         n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642,
         n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650,
         n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658,
         n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666,
         n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674,
         n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682,
         n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690,
         n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698,
         n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706,
         n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714,
         n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722,
         n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730,
         n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738,
         n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746,
         n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754,
         n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762,
         n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770,
         n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778,
         n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786,
         n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794,
         n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802,
         n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810,
         n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818,
         n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826,
         n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834,
         n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842,
         n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850,
         n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858,
         n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866,
         n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874,
         n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882,
         n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890,
         n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898,
         n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906,
         n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914,
         n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922,
         n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930,
         n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938,
         n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946,
         n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954,
         n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962,
         n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970,
         n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978,
         n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986,
         n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994,
         n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002,
         n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010,
         n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018,
         n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026,
         n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034,
         n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042,
         n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050,
         n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058,
         n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066,
         n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074,
         n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082,
         n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090,
         n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098,
         n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106,
         n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114,
         n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122,
         n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130,
         n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138,
         n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146,
         n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154,
         n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162,
         n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170,
         n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178,
         n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186,
         n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194,
         n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202,
         n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210,
         n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218,
         n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226,
         n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234,
         n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242,
         n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250,
         n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258,
         n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266,
         n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274,
         n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282,
         n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290,
         n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298,
         n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306,
         n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314,
         n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322,
         n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330,
         n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338,
         n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346,
         n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354,
         n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362,
         n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370,
         n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378,
         n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386,
         n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394,
         n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402,
         n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410,
         n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418,
         n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426,
         n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434,
         n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442,
         n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450,
         n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458,
         n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466,
         n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474,
         n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482,
         n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490,
         n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498,
         n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506,
         n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514,
         n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522,
         n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530,
         n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538,
         n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546,
         n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554,
         n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562,
         n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570,
         n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578,
         n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586,
         n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594,
         n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602,
         n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610,
         n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618,
         n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626,
         n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634,
         n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642,
         n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650,
         n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658,
         n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666,
         n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674,
         n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682,
         n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690,
         n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698,
         n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706,
         n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714,
         n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722,
         n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730,
         n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738,
         n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746,
         n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754,
         n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762,
         n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770,
         n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778,
         n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786,
         n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794,
         n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802,
         n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810,
         n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818,
         n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826,
         n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834,
         n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842,
         n12843, n12844, n12845;
  wire   [29:0] ICACHE_addr;
  assign DCACHE_addr[13] = net118926;

  DFFRX4 \i_MIPS/EX_MEM_reg[9]  ( .D(\i_MIPS/n395 ), .CK(clk), .RN(n6322), .Q(
        n12979), .QN(n3930) );
  DFFRX4 \i_MIPS/ID_EX_reg[7]  ( .D(\i_MIPS/n401 ), .CK(clk), .RN(n6322), .Q(
        \i_MIPS/ALUOp[1] ), .QN(n3964) );
  DFFRX4 \i_MIPS/ID_EX_reg[5]  ( .D(\i_MIPS/n408 ), .CK(clk), .RN(n6321), .Q(
        \i_MIPS/ID_EX_5 ), .QN(n4790) );
  DFFRX4 \i_MIPS/ID_EX_reg[83]  ( .D(\i_MIPS/n438 ), .CK(clk), .RN(n6318), .Q(
        \i_MIPS/ID_EX[83] ), .QN(net134375) );
  DFFRX4 \i_MIPS/ID_EX_reg[81]  ( .D(\i_MIPS/n440 ), .CK(clk), .RN(n6318), .Q(
        \i_MIPS/ID_EX[81] ), .QN(n3903) );
  DFFRX4 \i_MIPS/ID_EX_reg[78]  ( .D(\i_MIPS/n443 ), .CK(clk), .RN(n6318), .Q(
        \i_MIPS/ID_EX[78] ), .QN(net134414) );
  DFFRX4 \i_MIPS/ID_EX_reg[76]  ( .D(\i_MIPS/n445 ), .CK(clk), .RN(n6317), .Q(
        \i_MIPS/ID_EX[76] ), .QN(n3908) );
  DFFRX4 \i_MIPS/ID_EX_reg[74]  ( .D(\i_MIPS/n447 ), .CK(clk), .RN(n6317), .Q(
        \i_MIPS/ID_EX[74] ), .QN(n4021) );
  DFFRX4 \i_MIPS/IF_ID_reg[34]  ( .D(\i_MIPS/N51 ), .CK(clk), .RN(n6317), .Q(
        \i_MIPS/Sign_Extend[2] ), .QN(\i_MIPS/n519 ) );
  DFFRX4 \i_MIPS/IF_ID_reg[48]  ( .D(\i_MIPS/N65 ), .CK(clk), .RN(n6316), .Q(
        \i_MIPS/jump_addr[18] ), .QN(\i_MIPS/n505 ) );
  DFFRX4 \i_MIPS/IF_ID_reg[49]  ( .D(\i_MIPS/N66 ), .CK(clk), .RN(n6316), .Q(
        n248), .QN(\i_MIPS/n504 ) );
  DFFRX4 \i_MIPS/IF_ID_reg[50]  ( .D(\i_MIPS/N67 ), .CK(clk), .RN(n6315), .QN(
        \i_MIPS/n503 ) );
  DFFRX4 \i_MIPS/IF_ID_reg[51]  ( .D(\i_MIPS/N68 ), .CK(clk), .RN(n6315), .QN(
        \i_MIPS/n502 ) );
  DFFRX4 \i_MIPS/IF_ID_reg[53]  ( .D(\i_MIPS/N70 ), .CK(clk), .RN(n6315), .Q(
        \i_MIPS/jump_addr[23] ), .QN(\i_MIPS/n500 ) );
  DFFRX4 \i_MIPS/IF_ID_reg[54]  ( .D(\i_MIPS/N71 ), .CK(clk), .RN(n6315), .Q(
        n254), .QN(\i_MIPS/n499 ) );
  DFFRX4 \i_MIPS/IF_ID_reg[55]  ( .D(\i_MIPS/N72 ), .CK(clk), .RN(n6315), .QN(
        \i_MIPS/n498 ) );
  DFFRX4 \i_MIPS/IF_ID_reg[56]  ( .D(\i_MIPS/N73 ), .CK(clk), .RN(n6315), .Q(
        \i_MIPS/jump_addr[26] ), .QN(\i_MIPS/n497 ) );
  DFFRX4 \i_MIPS/ID_EX_reg[40]  ( .D(\i_MIPS/n461 ), .CK(clk), .RN(n6314), .Q(
        \i_MIPS/ALU/N303 ), .QN(\i_MIPS/n270 ) );
  DFFRX4 \i_MIPS/ID_EX_reg[30]  ( .D(\i_MIPS/n471 ), .CK(clk), .RN(n6313), .Q(
        \i_MIPS/ALUin1[21] ), .QN(n345) );
  DFFRX4 \i_MIPS/ID_EX_reg[21]  ( .D(\i_MIPS/n480 ), .CK(clk), .RN(n6312), .Q(
        \i_MIPS/ALUin1[12] ), .QN(n1263) );
  DFFRX4 \i_MIPS/ID_EX_reg[20]  ( .D(\i_MIPS/n481 ), .CK(clk), .RN(n6312), .Q(
        \i_MIPS/ALUin1[11] ), .QN(n3744) );
  DFFRX4 \i_MIPS/ID_EX_reg[18]  ( .D(\i_MIPS/n483 ), .CK(clk), .RN(n6312), .Q(
        \i_MIPS/ALUin1[9] ), .QN(n2920) );
  DFFRX4 \i_MIPS/ID_EX_reg[17]  ( .D(\i_MIPS/n484 ), .CK(clk), .RN(n6312), .Q(
        \i_MIPS/ALUin1[8] ), .QN(n343) );
  DFFRX4 \i_MIPS/ID_EX_reg[15]  ( .D(\i_MIPS/n486 ), .CK(clk), .RN(n6312), .Q(
        \i_MIPS/ALUin1[6] ), .QN(n1302) );
  DFFRX4 \i_MIPS/ID_EX_reg[10]  ( .D(\i_MIPS/n491 ), .CK(clk), .RN(n6311), .Q(
        \i_MIPS/ALUin1[1] ), .QN(\i_MIPS/n300 ) );
  DFFRX4 \i_MIPS/PC/PC_o_reg[4]  ( .D(\i_MIPS/PC/n38 ), .CK(clk), .RN(n6311), 
        .Q(ICACHE_addr[2]), .QN(\i_MIPS/PC/n6 ) );
  DFFRX4 \i_MIPS/PC/PC_o_reg[5]  ( .D(\i_MIPS/PC/n39 ), .CK(clk), .RN(n6311), 
        .Q(ICACHE_addr[3]), .QN(\i_MIPS/PC/n7 ) );
  DFFRX4 \i_MIPS/PC/PC_o_reg[6]  ( .D(\i_MIPS/PC/n40 ), .CK(clk), .RN(n6311), 
        .Q(ICACHE_addr[4]), .QN(\i_MIPS/PC/n8 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[1]  ( .D(\i_MIPS/N18 ), .CK(clk), .RN(n6330), .QN(
        \i_MIPS/n154 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[0]  ( .D(\i_MIPS/N17 ), .CK(clk), .RN(n6330), .QN(
        \i_MIPS/n153 ) );
  DFFRX1 \i_MIPS/PC/PC_o_reg[0]  ( .D(\i_MIPS/PC/n34 ), .CK(clk), .RN(n6311), 
        .Q(\i_MIPS/PC_add4[0] ), .QN(\i_MIPS/PC/n2 ) );
  DFFRX1 \i_MIPS/PC/PC_o_reg[1]  ( .D(\i_MIPS/PC/n35 ), .CK(clk), .RN(n6311), 
        .Q(\i_MIPS/PC_o[1] ), .QN(\i_MIPS/PC/n3 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[31]  ( .D(\i_MIPS/N48 ), .CK(clk), .RN(n6332), .Q(
        \i_MIPS/jump_addr[31] ), .QN(\i_MIPS/n522 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[1]  ( .D(\i_MIPS/n457 ), .CK(clk), .RN(n6314), .QN(
        \i_MIPS/n267 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[28]  ( .D(\i_MIPS/N45 ), .CK(clk), .RN(n6332), .Q(
        \i_MIPS/jump_addr[28] ), .QN(\i_MIPS/n525 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[116]  ( .D(\i_MIPS/n460 ), .CK(clk), .RN(n6314), 
        .QN(\i_MIPS/n269 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[29]  ( .D(\i_MIPS/N46 ), .CK(clk), .RN(n6332), .Q(
        \i_MIPS/jump_addr[29] ), .QN(\i_MIPS/n524 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[4]  ( .D(\i_MIPS/n410 ), .CK(clk), .RN(n6321), .QN(
        \i_MIPS/n246 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[30]  ( .D(\i_MIPS/N47 ), .CK(clk), .RN(n6332), .Q(
        \i_MIPS/jump_addr[30] ), .QN(\i_MIPS/n523 ) );
  DFFRX1 \i_MIPS/Register/register_reg[31][30]  ( .D(n11542), .CK(clk), .RN(
        n6306), .QN(n352) );
  DFFRX1 \i_MIPS/EX_MEM_reg[74]  ( .D(\i_MIPS/n459 ), .CK(clk), .RN(n6314), 
        .Q(\i_MIPS/EX_MEM_74 ), .QN(\i_MIPS/n268 ) );
  DFFRX1 \i_MIPS/Register/register_reg[28][22]  ( .D(\i_MIPS/Register/n234 ), 
        .CK(clk), .RN(n6299), .Q(\i_MIPS/Register/register[28][22] ), .QN(n370) );
  DFFRX1 \i_MIPS/Register/register_reg[27][30]  ( .D(\i_MIPS/Register/n274 ), 
        .CK(clk), .RN(n6295), .Q(\i_MIPS/Register/register[27][30] ), .QN(n364) );
  DFFRX1 \i_MIPS/Register/register_reg[24][22]  ( .D(\i_MIPS/Register/n362 ), 
        .CK(clk), .RN(n6288), .Q(\i_MIPS/Register/register[24][22] ), .QN(n362) );
  DFFRX1 \i_MIPS/Register/register_reg[23][30]  ( .D(\i_MIPS/Register/n402 ), 
        .CK(clk), .RN(n6285), .Q(\i_MIPS/Register/register[23][30] ), .QN(
        n1992) );
  DFFRX1 \i_MIPS/Register/register_reg[20][22]  ( .D(\i_MIPS/Register/n490 ), 
        .CK(clk), .RN(n6277), .Q(\i_MIPS/Register/register[20][22] ), .QN(
        n1996) );
  DFFRX1 \i_MIPS/Register/register_reg[16][22]  ( .D(\i_MIPS/Register/n618 ), 
        .CK(clk), .RN(n6267), .Q(\i_MIPS/Register/register[16][22] ), .QN(
        n2000) );
  DFFRX1 \i_MIPS/Register/register_reg[15][30]  ( .D(\i_MIPS/Register/n658 ), 
        .CK(clk), .RN(n6263), .Q(\i_MIPS/Register/register[15][30] ), .QN(n243) );
  DFFRX1 \i_MIPS/Register/register_reg[15][31]  ( .D(\i_MIPS/Register/n659 ), 
        .CK(clk), .RN(n6263), .Q(\i_MIPS/Register/register[15][31] ), .QN(n369) );
  DFFRX1 \i_MIPS/Register/register_reg[12][22]  ( .D(\i_MIPS/Register/n746 ), 
        .CK(clk), .RN(n6256), .Q(\i_MIPS/Register/register[12][22] ), .QN(n371) );
  DFFRX1 \i_MIPS/Register/register_reg[11][30]  ( .D(\i_MIPS/Register/n786 ), 
        .CK(clk), .RN(n6253), .Q(\i_MIPS/Register/register[11][30] ), .QN(n365) );
  DFFRX1 \i_MIPS/Register/register_reg[8][22]  ( .D(\i_MIPS/Register/n874 ), 
        .CK(clk), .RN(n6245), .Q(\i_MIPS/Register/register[8][22] ), .QN(n361)
         );
  DFFRX1 \i_MIPS/Register/register_reg[7][30]  ( .D(\i_MIPS/Register/n914 ), 
        .CK(clk), .RN(n6242), .Q(\i_MIPS/Register/register[7][30] ), .QN(n1995) );
  DFFRX1 \i_MIPS/Register/register_reg[4][22]  ( .D(\i_MIPS/Register/n1002 ), 
        .CK(clk), .RN(n6235), .Q(\i_MIPS/Register/register[4][22] ), .QN(n1997) );
  DFFRX1 \i_MIPS/Register/register_reg[0][22]  ( .D(\i_MIPS/Register/n1130 ), 
        .CK(clk), .RN(n6224), .Q(\i_MIPS/Register/register[0][22] ), .QN(n1999) );
  DFFRX1 \i_MIPS/EX_MEM_reg[6]  ( .D(\i_MIPS/n398 ), .CK(clk), .RN(n6322), .Q(
        \i_MIPS/EX_MEM[6] ) );
  DFFRX1 \I_cache/cache_reg[0][0]  ( .D(n12844), .CK(clk), .RN(n6120), .Q(
        \I_cache/cache[0][0] ), .QN(n1439) );
  DFFRX1 \I_cache/cache_reg[1][0]  ( .D(n12843), .CK(clk), .RN(n6120), .Q(
        \I_cache/cache[1][0] ), .QN(n3126) );
  DFFRX1 \I_cache/cache_reg[2][0]  ( .D(n12842), .CK(clk), .RN(n6120), .Q(
        \I_cache/cache[2][0] ), .QN(n1441) );
  DFFRX1 \I_cache/cache_reg[3][0]  ( .D(n12841), .CK(clk), .RN(n6120), .Q(
        \I_cache/cache[3][0] ), .QN(n3128) );
  DFFRX1 \I_cache/cache_reg[4][0]  ( .D(n12840), .CK(clk), .RN(n6119), .Q(
        \I_cache/cache[4][0] ), .QN(n1440) );
  DFFRX1 \I_cache/cache_reg[0][1]  ( .D(n12837), .CK(clk), .RN(n6119), .Q(
        \I_cache/cache[0][1] ), .QN(n1511) );
  DFFRX1 \I_cache/cache_reg[1][1]  ( .D(n12836), .CK(clk), .RN(n6119), .Q(
        \I_cache/cache[1][1] ), .QN(n3198) );
  DFFRX1 \I_cache/cache_reg[2][1]  ( .D(n12835), .CK(clk), .RN(n6119), .Q(
        \I_cache/cache[2][1] ), .QN(n1513) );
  DFFRX1 \I_cache/cache_reg[3][1]  ( .D(n12834), .CK(clk), .RN(n6119), .Q(
        \I_cache/cache[3][1] ), .QN(n3200) );
  DFFRX1 \I_cache/cache_reg[4][1]  ( .D(n12833), .CK(clk), .RN(n6119), .Q(
        \I_cache/cache[4][1] ), .QN(n1512) );
  DFFRX1 \I_cache/cache_reg[0][2]  ( .D(n12829), .CK(clk), .RN(n6118), .Q(
        \I_cache/cache[0][2] ), .QN(n1508) );
  DFFRX1 \I_cache/cache_reg[1][2]  ( .D(n12828), .CK(clk), .RN(n6118), .Q(
        \I_cache/cache[1][2] ), .QN(n3195) );
  DFFRX1 \I_cache/cache_reg[2][2]  ( .D(n12827), .CK(clk), .RN(n6118), .Q(
        \I_cache/cache[2][2] ), .QN(n1510) );
  DFFRX1 \I_cache/cache_reg[3][2]  ( .D(n12826), .CK(clk), .RN(n6118), .Q(
        \I_cache/cache[3][2] ), .QN(n3197) );
  DFFRX1 \I_cache/cache_reg[4][2]  ( .D(n12825), .CK(clk), .RN(n6118), .Q(
        \I_cache/cache[4][2] ), .QN(n1509) );
  DFFRX1 \I_cache/cache_reg[0][3]  ( .D(n12821), .CK(clk), .RN(n6118), .Q(
        \I_cache/cache[0][3] ), .QN(n1505) );
  DFFRX1 \I_cache/cache_reg[1][3]  ( .D(n12820), .CK(clk), .RN(n6118), .Q(
        \I_cache/cache[1][3] ), .QN(n3192) );
  DFFRX1 \I_cache/cache_reg[2][3]  ( .D(n12819), .CK(clk), .RN(n6118), .Q(
        \I_cache/cache[2][3] ), .QN(n1507) );
  DFFRX1 \I_cache/cache_reg[3][3]  ( .D(n12818), .CK(clk), .RN(n6118), .Q(
        \I_cache/cache[3][3] ), .QN(n3194) );
  DFFRX1 \I_cache/cache_reg[4][3]  ( .D(n12817), .CK(clk), .RN(n6117), .Q(
        \I_cache/cache[4][3] ), .QN(n1506) );
  DFFRX1 \I_cache/cache_reg[0][4]  ( .D(n12813), .CK(clk), .RN(n6117), .Q(
        \I_cache/cache[0][4] ), .QN(n1502) );
  DFFRX1 \I_cache/cache_reg[1][4]  ( .D(n12812), .CK(clk), .RN(n6117), .Q(
        \I_cache/cache[1][4] ), .QN(n3189) );
  DFFRX1 \I_cache/cache_reg[2][4]  ( .D(n12811), .CK(clk), .RN(n6117), .Q(
        \I_cache/cache[2][4] ), .QN(n1504) );
  DFFRX1 \I_cache/cache_reg[3][4]  ( .D(n12810), .CK(clk), .RN(n6117), .Q(
        \I_cache/cache[3][4] ), .QN(n3191) );
  DFFRX1 \I_cache/cache_reg[4][4]  ( .D(n12809), .CK(clk), .RN(n6117), .Q(
        \I_cache/cache[4][4] ), .QN(n1503) );
  DFFRX1 \I_cache/cache_reg[0][5]  ( .D(n12805), .CK(clk), .RN(n6116), .Q(
        \I_cache/cache[0][5] ), .QN(n1499) );
  DFFRX1 \I_cache/cache_reg[1][5]  ( .D(n12804), .CK(clk), .RN(n6116), .Q(
        \I_cache/cache[1][5] ), .QN(n3186) );
  DFFRX1 \I_cache/cache_reg[2][5]  ( .D(n12803), .CK(clk), .RN(n6116), .Q(
        \I_cache/cache[2][5] ), .QN(n1501) );
  DFFRX1 \I_cache/cache_reg[3][5]  ( .D(n12802), .CK(clk), .RN(n6116), .Q(
        \I_cache/cache[3][5] ), .QN(n3188) );
  DFFRX1 \I_cache/cache_reg[4][5]  ( .D(n12801), .CK(clk), .RN(n6116), .Q(
        \I_cache/cache[4][5] ), .QN(n1500) );
  DFFRX1 \I_cache/cache_reg[0][6]  ( .D(n12797), .CK(clk), .RN(n6116), .Q(
        \I_cache/cache[0][6] ), .QN(n1496) );
  DFFRX1 \I_cache/cache_reg[1][6]  ( .D(n12796), .CK(clk), .RN(n6116), .Q(
        \I_cache/cache[1][6] ), .QN(n3183) );
  DFFRX1 \I_cache/cache_reg[2][6]  ( .D(n12795), .CK(clk), .RN(n6116), .Q(
        \I_cache/cache[2][6] ), .QN(n1498) );
  DFFRX1 \I_cache/cache_reg[3][6]  ( .D(n12794), .CK(clk), .RN(n6116), .Q(
        \I_cache/cache[3][6] ), .QN(n3185) );
  DFFRX1 \I_cache/cache_reg[4][6]  ( .D(n12793), .CK(clk), .RN(n6115), .Q(
        \I_cache/cache[4][6] ), .QN(n1497) );
  DFFRX1 \I_cache/cache_reg[0][7]  ( .D(n12789), .CK(clk), .RN(n6115), .Q(
        \I_cache/cache[0][7] ), .QN(n1493) );
  DFFRX1 \I_cache/cache_reg[1][7]  ( .D(n12788), .CK(clk), .RN(n6115), .Q(
        \I_cache/cache[1][7] ), .QN(n3180) );
  DFFRX1 \I_cache/cache_reg[2][7]  ( .D(n12787), .CK(clk), .RN(n6115), .Q(
        \I_cache/cache[2][7] ), .QN(n1495) );
  DFFRX1 \I_cache/cache_reg[3][7]  ( .D(n12786), .CK(clk), .RN(n6115), .Q(
        \I_cache/cache[3][7] ), .QN(n3182) );
  DFFRX1 \I_cache/cache_reg[4][7]  ( .D(n12785), .CK(clk), .RN(n6115), .Q(
        \I_cache/cache[4][7] ), .QN(n1494) );
  DFFRX1 \I_cache/cache_reg[0][8]  ( .D(n12781), .CK(clk), .RN(n6114), .Q(
        \I_cache/cache[0][8] ), .QN(n1490) );
  DFFRX1 \I_cache/cache_reg[1][8]  ( .D(n12780), .CK(clk), .RN(n6114), .Q(
        \I_cache/cache[1][8] ), .QN(n3177) );
  DFFRX1 \I_cache/cache_reg[2][8]  ( .D(n12779), .CK(clk), .RN(n6114), .Q(
        \I_cache/cache[2][8] ), .QN(n1492) );
  DFFRX1 \I_cache/cache_reg[3][8]  ( .D(n12778), .CK(clk), .RN(n6114), .Q(
        \I_cache/cache[3][8] ), .QN(n3179) );
  DFFRX1 \I_cache/cache_reg[4][8]  ( .D(n12777), .CK(clk), .RN(n6114), .Q(
        \I_cache/cache[4][8] ), .QN(n1491) );
  DFFRX1 \I_cache/cache_reg[0][9]  ( .D(n12773), .CK(clk), .RN(n6114), .Q(
        \I_cache/cache[0][9] ), .QN(n1487) );
  DFFRX1 \I_cache/cache_reg[1][9]  ( .D(n12772), .CK(clk), .RN(n6114), .Q(
        \I_cache/cache[1][9] ), .QN(n3174) );
  DFFRX1 \I_cache/cache_reg[2][9]  ( .D(n12771), .CK(clk), .RN(n6114), .Q(
        \I_cache/cache[2][9] ), .QN(n1489) );
  DFFRX1 \I_cache/cache_reg[3][9]  ( .D(n12770), .CK(clk), .RN(n6114), .Q(
        \I_cache/cache[3][9] ), .QN(n3176) );
  DFFRX1 \I_cache/cache_reg[4][9]  ( .D(n12769), .CK(clk), .RN(n6113), .Q(
        \I_cache/cache[4][9] ), .QN(n1488) );
  DFFRX1 \I_cache/cache_reg[0][10]  ( .D(n12765), .CK(clk), .RN(n6113), .Q(
        \I_cache/cache[0][10] ), .QN(n1484) );
  DFFRX1 \I_cache/cache_reg[1][10]  ( .D(n12764), .CK(clk), .RN(n6113), .Q(
        \I_cache/cache[1][10] ), .QN(n3171) );
  DFFRX1 \I_cache/cache_reg[2][10]  ( .D(n12763), .CK(clk), .RN(n6113), .Q(
        \I_cache/cache[2][10] ), .QN(n1486) );
  DFFRX1 \I_cache/cache_reg[3][10]  ( .D(n12762), .CK(clk), .RN(n6113), .Q(
        \I_cache/cache[3][10] ), .QN(n3173) );
  DFFRX1 \I_cache/cache_reg[4][10]  ( .D(n12761), .CK(clk), .RN(n6113), .Q(
        \I_cache/cache[4][10] ), .QN(n1485) );
  DFFRX1 \I_cache/cache_reg[0][11]  ( .D(n12757), .CK(clk), .RN(n6112), .Q(
        \I_cache/cache[0][11] ), .QN(n1481) );
  DFFRX1 \I_cache/cache_reg[1][11]  ( .D(n12756), .CK(clk), .RN(n6112), .Q(
        \I_cache/cache[1][11] ), .QN(n3168) );
  DFFRX1 \I_cache/cache_reg[2][11]  ( .D(n12755), .CK(clk), .RN(n6112), .Q(
        \I_cache/cache[2][11] ), .QN(n1483) );
  DFFRX1 \I_cache/cache_reg[3][11]  ( .D(n12754), .CK(clk), .RN(n6112), .Q(
        \I_cache/cache[3][11] ), .QN(n3170) );
  DFFRX1 \I_cache/cache_reg[4][11]  ( .D(n12753), .CK(clk), .RN(n6112), .Q(
        \I_cache/cache[4][11] ), .QN(n1482) );
  DFFRX1 \I_cache/cache_reg[0][12]  ( .D(n12749), .CK(clk), .RN(n6112), .Q(
        \I_cache/cache[0][12] ), .QN(n1478) );
  DFFRX1 \I_cache/cache_reg[1][12]  ( .D(n12748), .CK(clk), .RN(n6112), .Q(
        \I_cache/cache[1][12] ), .QN(n3165) );
  DFFRX1 \I_cache/cache_reg[2][12]  ( .D(n12747), .CK(clk), .RN(n6112), .Q(
        \I_cache/cache[2][12] ), .QN(n1480) );
  DFFRX1 \I_cache/cache_reg[3][12]  ( .D(n12746), .CK(clk), .RN(n6112), .Q(
        \I_cache/cache[3][12] ), .QN(n3167) );
  DFFRX1 \I_cache/cache_reg[4][12]  ( .D(n12745), .CK(clk), .RN(n6111), .Q(
        \I_cache/cache[4][12] ), .QN(n1479) );
  DFFRX1 \I_cache/cache_reg[0][13]  ( .D(n12741), .CK(clk), .RN(n6111), .Q(
        \I_cache/cache[0][13] ), .QN(n1475) );
  DFFRX1 \I_cache/cache_reg[1][13]  ( .D(n12740), .CK(clk), .RN(n6111), .Q(
        \I_cache/cache[1][13] ), .QN(n3162) );
  DFFRX1 \I_cache/cache_reg[2][13]  ( .D(n12739), .CK(clk), .RN(n6111), .Q(
        \I_cache/cache[2][13] ), .QN(n1477) );
  DFFRX1 \I_cache/cache_reg[3][13]  ( .D(n12738), .CK(clk), .RN(n6111), .Q(
        \I_cache/cache[3][13] ), .QN(n3164) );
  DFFRX1 \I_cache/cache_reg[4][13]  ( .D(n12737), .CK(clk), .RN(n6111), .Q(
        \I_cache/cache[4][13] ), .QN(n1476) );
  DFFRX1 \I_cache/cache_reg[0][14]  ( .D(n12733), .CK(clk), .RN(n6110), .Q(
        \I_cache/cache[0][14] ), .QN(n1472) );
  DFFRX1 \I_cache/cache_reg[1][14]  ( .D(n12732), .CK(clk), .RN(n6110), .Q(
        \I_cache/cache[1][14] ), .QN(n3159) );
  DFFRX1 \I_cache/cache_reg[2][14]  ( .D(n12731), .CK(clk), .RN(n6110), .Q(
        \I_cache/cache[2][14] ), .QN(n1474) );
  DFFRX1 \I_cache/cache_reg[3][14]  ( .D(n12730), .CK(clk), .RN(n6110), .Q(
        \I_cache/cache[3][14] ), .QN(n3161) );
  DFFRX1 \I_cache/cache_reg[4][14]  ( .D(n12729), .CK(clk), .RN(n6110), .Q(
        \I_cache/cache[4][14] ), .QN(n1473) );
  DFFRX1 \I_cache/cache_reg[0][15]  ( .D(n12725), .CK(clk), .RN(n6110), .Q(
        \I_cache/cache[0][15] ), .QN(n1469) );
  DFFRX1 \I_cache/cache_reg[1][15]  ( .D(n12724), .CK(clk), .RN(n6110), .Q(
        \I_cache/cache[1][15] ), .QN(n3156) );
  DFFRX1 \I_cache/cache_reg[2][15]  ( .D(n12723), .CK(clk), .RN(n6110), .Q(
        \I_cache/cache[2][15] ), .QN(n1471) );
  DFFRX1 \I_cache/cache_reg[3][15]  ( .D(n12722), .CK(clk), .RN(n6110), .Q(
        \I_cache/cache[3][15] ), .QN(n3158) );
  DFFRX1 \I_cache/cache_reg[4][15]  ( .D(n12721), .CK(clk), .RN(n6109), .Q(
        \I_cache/cache[4][15] ), .QN(n1470) );
  DFFRX1 \I_cache/cache_reg[0][16]  ( .D(n12717), .CK(clk), .RN(n6109), .Q(
        \I_cache/cache[0][16] ), .QN(n1466) );
  DFFRX1 \I_cache/cache_reg[1][16]  ( .D(n12716), .CK(clk), .RN(n6109), .Q(
        \I_cache/cache[1][16] ), .QN(n3153) );
  DFFRX1 \I_cache/cache_reg[2][16]  ( .D(n12715), .CK(clk), .RN(n6109), .Q(
        \I_cache/cache[2][16] ), .QN(n1468) );
  DFFRX1 \I_cache/cache_reg[3][16]  ( .D(n12714), .CK(clk), .RN(n6109), .Q(
        \I_cache/cache[3][16] ), .QN(n3155) );
  DFFRX1 \I_cache/cache_reg[4][16]  ( .D(n12713), .CK(clk), .RN(n6109), .Q(
        \I_cache/cache[4][16] ), .QN(n1467) );
  DFFRX1 \I_cache/cache_reg[0][17]  ( .D(n12709), .CK(clk), .RN(n6108), .Q(
        \I_cache/cache[0][17] ), .QN(n1463) );
  DFFRX1 \I_cache/cache_reg[1][17]  ( .D(n12708), .CK(clk), .RN(n6108), .Q(
        \I_cache/cache[1][17] ), .QN(n3150) );
  DFFRX1 \I_cache/cache_reg[2][17]  ( .D(n12707), .CK(clk), .RN(n6108), .Q(
        \I_cache/cache[2][17] ), .QN(n1465) );
  DFFRX1 \I_cache/cache_reg[3][17]  ( .D(n12706), .CK(clk), .RN(n6108), .Q(
        \I_cache/cache[3][17] ), .QN(n3152) );
  DFFRX1 \I_cache/cache_reg[4][17]  ( .D(n12705), .CK(clk), .RN(n6108), .Q(
        \I_cache/cache[4][17] ), .QN(n1464) );
  DFFRX1 \I_cache/cache_reg[0][18]  ( .D(n12701), .CK(clk), .RN(n6108), .Q(
        \I_cache/cache[0][18] ), .QN(n1460) );
  DFFRX1 \I_cache/cache_reg[1][18]  ( .D(n12700), .CK(clk), .RN(n6108), .Q(
        \I_cache/cache[1][18] ), .QN(n3147) );
  DFFRX1 \I_cache/cache_reg[2][18]  ( .D(n12699), .CK(clk), .RN(n6108), .Q(
        \I_cache/cache[2][18] ), .QN(n1462) );
  DFFRX1 \I_cache/cache_reg[3][18]  ( .D(n12698), .CK(clk), .RN(n6108), .Q(
        \I_cache/cache[3][18] ), .QN(n3149) );
  DFFRX1 \I_cache/cache_reg[4][18]  ( .D(n12697), .CK(clk), .RN(n6107), .Q(
        \I_cache/cache[4][18] ), .QN(n1461) );
  DFFRX1 \I_cache/cache_reg[0][19]  ( .D(n12693), .CK(clk), .RN(n6107), .Q(
        \I_cache/cache[0][19] ), .QN(n1596) );
  DFFRX1 \I_cache/cache_reg[1][19]  ( .D(n12692), .CK(clk), .RN(n6107), .Q(
        \I_cache/cache[1][19] ), .QN(n3283) );
  DFFRX1 \I_cache/cache_reg[2][19]  ( .D(n12691), .CK(clk), .RN(n6107), .Q(
        \I_cache/cache[2][19] ), .QN(n1598) );
  DFFRX1 \I_cache/cache_reg[3][19]  ( .D(n12690), .CK(clk), .RN(n6107), .Q(
        \I_cache/cache[3][19] ), .QN(n3285) );
  DFFRX1 \I_cache/cache_reg[4][19]  ( .D(n12689), .CK(clk), .RN(n6107), .Q(
        \I_cache/cache[4][19] ), .QN(n1597) );
  DFFRX1 \I_cache/cache_reg[0][20]  ( .D(n12685), .CK(clk), .RN(n6106), .Q(
        \I_cache/cache[0][20] ), .QN(n1457) );
  DFFRX1 \I_cache/cache_reg[1][20]  ( .D(n12684), .CK(clk), .RN(n6106), .Q(
        \I_cache/cache[1][20] ), .QN(n3144) );
  DFFRX1 \I_cache/cache_reg[2][20]  ( .D(n12683), .CK(clk), .RN(n6106), .Q(
        \I_cache/cache[2][20] ), .QN(n1459) );
  DFFRX1 \I_cache/cache_reg[3][20]  ( .D(n12682), .CK(clk), .RN(n6106), .Q(
        \I_cache/cache[3][20] ), .QN(n3146) );
  DFFRX1 \I_cache/cache_reg[4][20]  ( .D(n12681), .CK(clk), .RN(n6106), .Q(
        \I_cache/cache[4][20] ), .QN(n1458) );
  DFFRX1 \I_cache/cache_reg[0][21]  ( .D(n12677), .CK(clk), .RN(n6106), .Q(
        \I_cache/cache[0][21] ), .QN(n1454) );
  DFFRX1 \I_cache/cache_reg[1][21]  ( .D(n12676), .CK(clk), .RN(n6106), .Q(
        \I_cache/cache[1][21] ), .QN(n3141) );
  DFFRX1 \I_cache/cache_reg[2][21]  ( .D(n12675), .CK(clk), .RN(n6106), .Q(
        \I_cache/cache[2][21] ), .QN(n1456) );
  DFFRX1 \I_cache/cache_reg[3][21]  ( .D(n12674), .CK(clk), .RN(n6106), .Q(
        \I_cache/cache[3][21] ), .QN(n3143) );
  DFFRX1 \I_cache/cache_reg[4][21]  ( .D(n12673), .CK(clk), .RN(n6105), .Q(
        \I_cache/cache[4][21] ), .QN(n1455) );
  DFFRX1 \I_cache/cache_reg[0][22]  ( .D(n12669), .CK(clk), .RN(n6105), .Q(
        \I_cache/cache[0][22] ), .QN(n1451) );
  DFFRX1 \I_cache/cache_reg[1][22]  ( .D(n12668), .CK(clk), .RN(n6105), .Q(
        \I_cache/cache[1][22] ), .QN(n3138) );
  DFFRX1 \I_cache/cache_reg[2][22]  ( .D(n12667), .CK(clk), .RN(n6105), .Q(
        \I_cache/cache[2][22] ), .QN(n1453) );
  DFFRX1 \I_cache/cache_reg[3][22]  ( .D(n12666), .CK(clk), .RN(n6105), .Q(
        \I_cache/cache[3][22] ), .QN(n3140) );
  DFFRX1 \I_cache/cache_reg[4][22]  ( .D(n12665), .CK(clk), .RN(n6105), .Q(
        \I_cache/cache[4][22] ), .QN(n1452) );
  DFFRX1 \I_cache/cache_reg[0][23]  ( .D(n12661), .CK(clk), .RN(n6104), .Q(
        \I_cache/cache[0][23] ), .QN(n1448) );
  DFFRX1 \I_cache/cache_reg[1][23]  ( .D(n12660), .CK(clk), .RN(n6104), .Q(
        \I_cache/cache[1][23] ), .QN(n3135) );
  DFFRX1 \I_cache/cache_reg[2][23]  ( .D(n12659), .CK(clk), .RN(n6104), .Q(
        \I_cache/cache[2][23] ), .QN(n1450) );
  DFFRX1 \I_cache/cache_reg[3][23]  ( .D(n12658), .CK(clk), .RN(n6104), .Q(
        \I_cache/cache[3][23] ), .QN(n3137) );
  DFFRX1 \I_cache/cache_reg[4][23]  ( .D(n12657), .CK(clk), .RN(n6104), .Q(
        \I_cache/cache[4][23] ), .QN(n1449) );
  DFFRX1 \I_cache/cache_reg[0][24]  ( .D(n12653), .CK(clk), .RN(n6104), .Q(
        \I_cache/cache[0][24] ), .QN(n1445) );
  DFFRX1 \I_cache/cache_reg[1][24]  ( .D(n12652), .CK(clk), .RN(n6104), .Q(
        \I_cache/cache[1][24] ), .QN(n3132) );
  DFFRX1 \I_cache/cache_reg[2][24]  ( .D(n12651), .CK(clk), .RN(n6104), .Q(
        \I_cache/cache[2][24] ), .QN(n1447) );
  DFFRX1 \I_cache/cache_reg[3][24]  ( .D(n12650), .CK(clk), .RN(n6104), .Q(
        \I_cache/cache[3][24] ), .QN(n3134) );
  DFFRX1 \I_cache/cache_reg[4][24]  ( .D(n12649), .CK(clk), .RN(n6103), .Q(
        \I_cache/cache[4][24] ), .QN(n1446) );
  DFFRX1 \I_cache/cache_reg[0][25]  ( .D(n12645), .CK(clk), .RN(n6103), .Q(
        \I_cache/cache[0][25] ), .QN(n1442) );
  DFFRX1 \I_cache/cache_reg[1][25]  ( .D(n12644), .CK(clk), .RN(n6103), .Q(
        \I_cache/cache[1][25] ), .QN(n3129) );
  DFFRX1 \I_cache/cache_reg[2][25]  ( .D(n12643), .CK(clk), .RN(n6103), .Q(
        \I_cache/cache[2][25] ), .QN(n1444) );
  DFFRX1 \I_cache/cache_reg[3][25]  ( .D(n12642), .CK(clk), .RN(n6103), .Q(
        \I_cache/cache[3][25] ), .QN(n3131) );
  DFFRX1 \I_cache/cache_reg[4][25]  ( .D(n12641), .CK(clk), .RN(n6103), .Q(
        \I_cache/cache[4][25] ), .QN(n1443) );
  DFFRX1 \I_cache/cache_reg[0][26]  ( .D(n12637), .CK(clk), .RN(n6102), .Q(
        \I_cache/cache[0][26] ), .QN(n1526) );
  DFFRX1 \I_cache/cache_reg[1][26]  ( .D(n12636), .CK(clk), .RN(n6102), .Q(
        \I_cache/cache[1][26] ), .QN(n3213) );
  DFFRX1 \I_cache/cache_reg[2][26]  ( .D(n12635), .CK(clk), .RN(n6102), .Q(
        \I_cache/cache[2][26] ), .QN(n1528) );
  DFFRX1 \I_cache/cache_reg[3][26]  ( .D(n12634), .CK(clk), .RN(n6102), .Q(
        \I_cache/cache[3][26] ), .QN(n3215) );
  DFFRX1 \I_cache/cache_reg[4][26]  ( .D(n12633), .CK(clk), .RN(n6102), .Q(
        \I_cache/cache[4][26] ), .QN(n1527) );
  DFFRX1 \I_cache/cache_reg[0][27]  ( .D(n12629), .CK(clk), .RN(n6102), .Q(
        \I_cache/cache[0][27] ), .QN(n1523) );
  DFFRX1 \I_cache/cache_reg[1][27]  ( .D(n12628), .CK(clk), .RN(n6102), .Q(
        \I_cache/cache[1][27] ), .QN(n3210) );
  DFFRX1 \I_cache/cache_reg[2][27]  ( .D(n12627), .CK(clk), .RN(n6102), .Q(
        \I_cache/cache[2][27] ), .QN(n1525) );
  DFFRX1 \I_cache/cache_reg[3][27]  ( .D(n12626), .CK(clk), .RN(n6102), .Q(
        \I_cache/cache[3][27] ), .QN(n3212) );
  DFFRX1 \I_cache/cache_reg[4][27]  ( .D(n12625), .CK(clk), .RN(n6101), .Q(
        \I_cache/cache[4][27] ), .QN(n1524) );
  DFFRX1 \I_cache/cache_reg[0][28]  ( .D(n12621), .CK(clk), .RN(n6101), .Q(
        \I_cache/cache[0][28] ), .QN(n1520) );
  DFFRX1 \I_cache/cache_reg[1][28]  ( .D(n12620), .CK(clk), .RN(n6101), .Q(
        \I_cache/cache[1][28] ), .QN(n3207) );
  DFFRX1 \I_cache/cache_reg[2][28]  ( .D(n12619), .CK(clk), .RN(n6101), .Q(
        \I_cache/cache[2][28] ), .QN(n1522) );
  DFFRX1 \I_cache/cache_reg[3][28]  ( .D(n12618), .CK(clk), .RN(n6101), .Q(
        \I_cache/cache[3][28] ), .QN(n3209) );
  DFFRX1 \I_cache/cache_reg[4][28]  ( .D(n12617), .CK(clk), .RN(n6101), .Q(
        \I_cache/cache[4][28] ), .QN(n1521) );
  DFFRX1 \I_cache/cache_reg[0][29]  ( .D(n12613), .CK(clk), .RN(n6100), .Q(
        \I_cache/cache[0][29] ), .QN(n1517) );
  DFFRX1 \I_cache/cache_reg[1][29]  ( .D(n12612), .CK(clk), .RN(n6100), .Q(
        \I_cache/cache[1][29] ), .QN(n3204) );
  DFFRX1 \I_cache/cache_reg[2][29]  ( .D(n12611), .CK(clk), .RN(n6100), .Q(
        \I_cache/cache[2][29] ), .QN(n1519) );
  DFFRX1 \I_cache/cache_reg[3][29]  ( .D(n12610), .CK(clk), .RN(n6100), .Q(
        \I_cache/cache[3][29] ), .QN(n3206) );
  DFFRX1 \I_cache/cache_reg[4][29]  ( .D(n12609), .CK(clk), .RN(n6100), .Q(
        \I_cache/cache[4][29] ), .QN(n1518) );
  DFFRX1 \I_cache/cache_reg[0][30]  ( .D(n12605), .CK(clk), .RN(n6100), .Q(
        \I_cache/cache[0][30] ), .QN(n1514) );
  DFFRX1 \I_cache/cache_reg[1][30]  ( .D(n12604), .CK(clk), .RN(n6100), .Q(
        \I_cache/cache[1][30] ), .QN(n3201) );
  DFFRX1 \I_cache/cache_reg[2][30]  ( .D(n12603), .CK(clk), .RN(n6100), .Q(
        \I_cache/cache[2][30] ), .QN(n1516) );
  DFFRX1 \I_cache/cache_reg[3][30]  ( .D(n12602), .CK(clk), .RN(n6100), .Q(
        \I_cache/cache[3][30] ), .QN(n3203) );
  DFFRX1 \I_cache/cache_reg[4][30]  ( .D(n12601), .CK(clk), .RN(n6099), .Q(
        \I_cache/cache[4][30] ), .QN(n1515) );
  DFFRX1 \I_cache/cache_reg[0][31]  ( .D(n12597), .CK(clk), .RN(n6099), .Q(
        \I_cache/cache[0][31] ), .QN(n1591) );
  DFFRX1 \I_cache/cache_reg[1][31]  ( .D(n12596), .CK(clk), .RN(n6099), .Q(
        \I_cache/cache[1][31] ), .QN(n3278) );
  DFFRX1 \I_cache/cache_reg[2][31]  ( .D(n12595), .CK(clk), .RN(n6099), .Q(
        \I_cache/cache[2][31] ), .QN(n1589) );
  DFFRX1 \I_cache/cache_reg[3][31]  ( .D(n12594), .CK(clk), .RN(n6099), .Q(
        \I_cache/cache[3][31] ), .QN(n3276) );
  DFFRX1 \I_cache/cache_reg[4][31]  ( .D(n12593), .CK(clk), .RN(n6099), .Q(
        \I_cache/cache[4][31] ), .QN(n1592) );
  DFFRX1 \I_cache/cache_reg[5][31]  ( .D(n12592), .CK(clk), .RN(n6099), .Q(
        \I_cache/cache[5][31] ), .QN(n3279) );
  DFFRX1 \I_cache/cache_reg[6][31]  ( .D(n12591), .CK(clk), .RN(n6099), .Q(
        \I_cache/cache[6][31] ), .QN(n1590) );
  DFFRX1 \I_cache/cache_reg[7][31]  ( .D(n12590), .CK(clk), .RN(n6099), .Q(
        \I_cache/cache[7][31] ), .QN(n3277) );
  DFFRX1 \I_cache/cache_reg[0][32]  ( .D(n12589), .CK(clk), .RN(n6098), .Q(
        \I_cache/cache[0][32] ), .QN(n1692) );
  DFFRX1 \I_cache/cache_reg[1][32]  ( .D(n12588), .CK(clk), .RN(n6098), .Q(
        \I_cache/cache[1][32] ), .QN(n3380) );
  DFFRX1 \I_cache/cache_reg[2][32]  ( .D(n12587), .CK(clk), .RN(n6098), .Q(
        \I_cache/cache[2][32] ), .QN(n1694) );
  DFFRX1 \I_cache/cache_reg[0][33]  ( .D(n12581), .CK(clk), .RN(n6098), .Q(
        \I_cache/cache[0][33] ), .QN(n1764) );
  DFFRX1 \I_cache/cache_reg[1][33]  ( .D(n12580), .CK(clk), .RN(n6098), .Q(
        \I_cache/cache[1][33] ), .QN(n3452) );
  DFFRX1 \I_cache/cache_reg[2][33]  ( .D(n12579), .CK(clk), .RN(n6098), .Q(
        \I_cache/cache[2][33] ), .QN(n1766) );
  DFFRX1 \I_cache/cache_reg[0][34]  ( .D(n12573), .CK(clk), .RN(n6097), .Q(
        \I_cache/cache[0][34] ), .QN(n1761) );
  DFFRX1 \I_cache/cache_reg[1][34]  ( .D(n12572), .CK(clk), .RN(n6097), .Q(
        \I_cache/cache[1][34] ), .QN(n3449) );
  DFFRX1 \I_cache/cache_reg[2][34]  ( .D(n12571), .CK(clk), .RN(n6097), .Q(
        \I_cache/cache[2][34] ), .QN(n1763) );
  DFFRX1 \I_cache/cache_reg[0][35]  ( .D(n12565), .CK(clk), .RN(n6096), .Q(
        \I_cache/cache[0][35] ), .QN(n1758) );
  DFFRX1 \I_cache/cache_reg[1][35]  ( .D(n12564), .CK(clk), .RN(n6096), .Q(
        \I_cache/cache[1][35] ), .QN(n3446) );
  DFFRX1 \I_cache/cache_reg[2][35]  ( .D(n12563), .CK(clk), .RN(n6096), .Q(
        \I_cache/cache[2][35] ), .QN(n1760) );
  DFFRX1 \I_cache/cache_reg[0][36]  ( .D(n12557), .CK(clk), .RN(n6096), .Q(
        \I_cache/cache[0][36] ), .QN(n1755) );
  DFFRX1 \I_cache/cache_reg[1][36]  ( .D(n12556), .CK(clk), .RN(n6096), .Q(
        \I_cache/cache[1][36] ), .QN(n3443) );
  DFFRX1 \I_cache/cache_reg[2][36]  ( .D(n12555), .CK(clk), .RN(n6096), .Q(
        \I_cache/cache[2][36] ), .QN(n1757) );
  DFFRX1 \I_cache/cache_reg[0][37]  ( .D(n12549), .CK(clk), .RN(n6095), .Q(
        \I_cache/cache[0][37] ), .QN(n1752) );
  DFFRX1 \I_cache/cache_reg[1][37]  ( .D(n12548), .CK(clk), .RN(n6095), .Q(
        \I_cache/cache[1][37] ), .QN(n3440) );
  DFFRX1 \I_cache/cache_reg[2][37]  ( .D(n12547), .CK(clk), .RN(n6095), .Q(
        \I_cache/cache[2][37] ), .QN(n1754) );
  DFFRX1 \I_cache/cache_reg[0][38]  ( .D(n12541), .CK(clk), .RN(n6094), .Q(
        \I_cache/cache[0][38] ), .QN(n1749) );
  DFFRX1 \I_cache/cache_reg[1][38]  ( .D(n12540), .CK(clk), .RN(n6094), .Q(
        \I_cache/cache[1][38] ), .QN(n3437) );
  DFFRX1 \I_cache/cache_reg[2][38]  ( .D(n12539), .CK(clk), .RN(n6094), .Q(
        \I_cache/cache[2][38] ), .QN(n1751) );
  DFFRX1 \I_cache/cache_reg[0][39]  ( .D(n12533), .CK(clk), .RN(n6094), .Q(
        \I_cache/cache[0][39] ), .QN(n1746) );
  DFFRX1 \I_cache/cache_reg[1][39]  ( .D(n12532), .CK(clk), .RN(n6094), .Q(
        \I_cache/cache[1][39] ), .QN(n3434) );
  DFFRX1 \I_cache/cache_reg[2][39]  ( .D(n12531), .CK(clk), .RN(n6094), .Q(
        \I_cache/cache[2][39] ), .QN(n1748) );
  DFFRX1 \I_cache/cache_reg[0][40]  ( .D(n12525), .CK(clk), .RN(n6093), .Q(
        \I_cache/cache[0][40] ), .QN(n1743) );
  DFFRX1 \I_cache/cache_reg[1][40]  ( .D(n12524), .CK(clk), .RN(n6093), .Q(
        \I_cache/cache[1][40] ), .QN(n3431) );
  DFFRX1 \I_cache/cache_reg[2][40]  ( .D(n12523), .CK(clk), .RN(n6093), .Q(
        \I_cache/cache[2][40] ), .QN(n1745) );
  DFFRX1 \I_cache/cache_reg[0][41]  ( .D(n12517), .CK(clk), .RN(n6092), .Q(
        \I_cache/cache[0][41] ), .QN(n1740) );
  DFFRX1 \I_cache/cache_reg[1][41]  ( .D(n12516), .CK(clk), .RN(n6092), .Q(
        \I_cache/cache[1][41] ), .QN(n3428) );
  DFFRX1 \I_cache/cache_reg[2][41]  ( .D(n12515), .CK(clk), .RN(n6092), .Q(
        \I_cache/cache[2][41] ), .QN(n1742) );
  DFFRX1 \I_cache/cache_reg[0][42]  ( .D(n12509), .CK(clk), .RN(n6092), .Q(
        \I_cache/cache[0][42] ), .QN(n1737) );
  DFFRX1 \I_cache/cache_reg[1][42]  ( .D(n12508), .CK(clk), .RN(n6092), .Q(
        \I_cache/cache[1][42] ), .QN(n3425) );
  DFFRX1 \I_cache/cache_reg[2][42]  ( .D(n12507), .CK(clk), .RN(n6092), .Q(
        \I_cache/cache[2][42] ), .QN(n1739) );
  DFFRX1 \I_cache/cache_reg[0][43]  ( .D(n12501), .CK(clk), .RN(n6091), .Q(
        \I_cache/cache[0][43] ), .QN(n1734) );
  DFFRX1 \I_cache/cache_reg[1][43]  ( .D(n12500), .CK(clk), .RN(n6091), .Q(
        \I_cache/cache[1][43] ), .QN(n3422) );
  DFFRX1 \I_cache/cache_reg[2][43]  ( .D(n12499), .CK(clk), .RN(n6091), .Q(
        \I_cache/cache[2][43] ), .QN(n1736) );
  DFFRX1 \I_cache/cache_reg[0][44]  ( .D(n12493), .CK(clk), .RN(n6090), .Q(
        \I_cache/cache[0][44] ), .QN(n1731) );
  DFFRX1 \I_cache/cache_reg[1][44]  ( .D(n12492), .CK(clk), .RN(n6090), .Q(
        \I_cache/cache[1][44] ), .QN(n3419) );
  DFFRX1 \I_cache/cache_reg[2][44]  ( .D(n12491), .CK(clk), .RN(n6090), .Q(
        \I_cache/cache[2][44] ), .QN(n1733) );
  DFFRX1 \I_cache/cache_reg[0][45]  ( .D(n12485), .CK(clk), .RN(n6090), .Q(
        \I_cache/cache[0][45] ), .QN(n1728) );
  DFFRX1 \I_cache/cache_reg[1][45]  ( .D(n12484), .CK(clk), .RN(n6090), .Q(
        \I_cache/cache[1][45] ), .QN(n3416) );
  DFFRX1 \I_cache/cache_reg[2][45]  ( .D(n12483), .CK(clk), .RN(n6090), .Q(
        \I_cache/cache[2][45] ), .QN(n1730) );
  DFFRX1 \I_cache/cache_reg[0][46]  ( .D(n12477), .CK(clk), .RN(n6089), .Q(
        \I_cache/cache[0][46] ), .QN(n1725) );
  DFFRX1 \I_cache/cache_reg[1][46]  ( .D(n12476), .CK(clk), .RN(n6089), .Q(
        \I_cache/cache[1][46] ), .QN(n3413) );
  DFFRX1 \I_cache/cache_reg[2][46]  ( .D(n12475), .CK(clk), .RN(n6089), .Q(
        \I_cache/cache[2][46] ), .QN(n1727) );
  DFFRX1 \I_cache/cache_reg[0][47]  ( .D(n12469), .CK(clk), .RN(n6088), .Q(
        \I_cache/cache[0][47] ), .QN(n1722) );
  DFFRX1 \I_cache/cache_reg[1][47]  ( .D(n12468), .CK(clk), .RN(n6088), .Q(
        \I_cache/cache[1][47] ), .QN(n3410) );
  DFFRX1 \I_cache/cache_reg[2][47]  ( .D(n12467), .CK(clk), .RN(n6088), .Q(
        \I_cache/cache[2][47] ), .QN(n1724) );
  DFFRX1 \I_cache/cache_reg[0][48]  ( .D(n12461), .CK(clk), .RN(n6088), .Q(
        \I_cache/cache[0][48] ), .QN(n1719) );
  DFFRX1 \I_cache/cache_reg[1][48]  ( .D(n12460), .CK(clk), .RN(n6088), .Q(
        \I_cache/cache[1][48] ), .QN(n3407) );
  DFFRX1 \I_cache/cache_reg[2][48]  ( .D(n12459), .CK(clk), .RN(n6088), .Q(
        \I_cache/cache[2][48] ), .QN(n1721) );
  DFFRX1 \I_cache/cache_reg[0][49]  ( .D(n12453), .CK(clk), .RN(n6087), .Q(
        \I_cache/cache[0][49] ), .QN(n1716) );
  DFFRX1 \I_cache/cache_reg[1][49]  ( .D(n12452), .CK(clk), .RN(n6087), .Q(
        \I_cache/cache[1][49] ), .QN(n3404) );
  DFFRX1 \I_cache/cache_reg[2][49]  ( .D(n12451), .CK(clk), .RN(n6087), .Q(
        \I_cache/cache[2][49] ), .QN(n1718) );
  DFFRX1 \I_cache/cache_reg[0][50]  ( .D(n12445), .CK(clk), .RN(n6086), .Q(
        \I_cache/cache[0][50] ), .QN(n1713) );
  DFFRX1 \I_cache/cache_reg[1][50]  ( .D(n12444), .CK(clk), .RN(n6086), .Q(
        \I_cache/cache[1][50] ), .QN(n3401) );
  DFFRX1 \I_cache/cache_reg[2][50]  ( .D(n12443), .CK(clk), .RN(n6086), .Q(
        \I_cache/cache[2][50] ), .QN(n1715) );
  DFFRX1 \I_cache/cache_reg[0][51]  ( .D(n12437), .CK(clk), .RN(n6086), .Q(
        \I_cache/cache[0][51] ), .QN(n1851) );
  DFFRX1 \I_cache/cache_reg[1][51]  ( .D(n12436), .CK(clk), .RN(n6086), .Q(
        \I_cache/cache[1][51] ), .QN(n3538) );
  DFFRX1 \I_cache/cache_reg[2][51]  ( .D(n12435), .CK(clk), .RN(n6086), .Q(
        \I_cache/cache[2][51] ), .QN(n1853) );
  DFFRX1 \I_cache/cache_reg[0][52]  ( .D(n12429), .CK(clk), .RN(n6085), .Q(
        \I_cache/cache[0][52] ), .QN(n1710) );
  DFFRX1 \I_cache/cache_reg[1][52]  ( .D(n12428), .CK(clk), .RN(n6085), .Q(
        \I_cache/cache[1][52] ), .QN(n3398) );
  DFFRX1 \I_cache/cache_reg[2][52]  ( .D(n12427), .CK(clk), .RN(n6085), .Q(
        \I_cache/cache[2][52] ), .QN(n1712) );
  DFFRX1 \I_cache/cache_reg[0][53]  ( .D(n12421), .CK(clk), .RN(n6084), .Q(
        \I_cache/cache[0][53] ), .QN(n1707) );
  DFFRX1 \I_cache/cache_reg[1][53]  ( .D(n12420), .CK(clk), .RN(n6084), .Q(
        \I_cache/cache[1][53] ), .QN(n3395) );
  DFFRX1 \I_cache/cache_reg[2][53]  ( .D(n12419), .CK(clk), .RN(n6084), .Q(
        \I_cache/cache[2][53] ), .QN(n1709) );
  DFFRX1 \I_cache/cache_reg[0][54]  ( .D(n12413), .CK(clk), .RN(n6084), .Q(
        \I_cache/cache[0][54] ), .QN(n1704) );
  DFFRX1 \I_cache/cache_reg[1][54]  ( .D(n12412), .CK(clk), .RN(n6084), .Q(
        \I_cache/cache[1][54] ), .QN(n3392) );
  DFFRX1 \I_cache/cache_reg[2][54]  ( .D(n12411), .CK(clk), .RN(n6084), .Q(
        \I_cache/cache[2][54] ), .QN(n1706) );
  DFFRX1 \I_cache/cache_reg[0][55]  ( .D(n12405), .CK(clk), .RN(n6083), .Q(
        \I_cache/cache[0][55] ), .QN(n1701) );
  DFFRX1 \I_cache/cache_reg[1][55]  ( .D(n12404), .CK(clk), .RN(n6083), .Q(
        \I_cache/cache[1][55] ), .QN(n3389) );
  DFFRX1 \I_cache/cache_reg[2][55]  ( .D(n12403), .CK(clk), .RN(n6083), .Q(
        \I_cache/cache[2][55] ), .QN(n1703) );
  DFFRX1 \I_cache/cache_reg[0][56]  ( .D(n12397), .CK(clk), .RN(n6082), .Q(
        \I_cache/cache[0][56] ), .QN(n1698) );
  DFFRX1 \I_cache/cache_reg[1][56]  ( .D(n12396), .CK(clk), .RN(n6082), .Q(
        \I_cache/cache[1][56] ), .QN(n3386) );
  DFFRX1 \I_cache/cache_reg[2][56]  ( .D(n12395), .CK(clk), .RN(n6082), .Q(
        \I_cache/cache[2][56] ), .QN(n1700) );
  DFFRX1 \I_cache/cache_reg[0][57]  ( .D(n12389), .CK(clk), .RN(n6082), .Q(
        \I_cache/cache[0][57] ), .QN(n1695) );
  DFFRX1 \I_cache/cache_reg[1][57]  ( .D(n12388), .CK(clk), .RN(n6082), .Q(
        \I_cache/cache[1][57] ), .QN(n3383) );
  DFFRX1 \I_cache/cache_reg[2][57]  ( .D(n12387), .CK(clk), .RN(n6082), .Q(
        \I_cache/cache[2][57] ), .QN(n1697) );
  DFFRX1 \I_cache/cache_reg[0][58]  ( .D(n12381), .CK(clk), .RN(n6081), .Q(
        \I_cache/cache[0][58] ), .QN(n1782) );
  DFFRX1 \I_cache/cache_reg[1][58]  ( .D(n12380), .CK(clk), .RN(n6081), .Q(
        \I_cache/cache[1][58] ), .QN(n3470) );
  DFFRX1 \I_cache/cache_reg[2][58]  ( .D(n12379), .CK(clk), .RN(n6081), .Q(
        \I_cache/cache[2][58] ), .QN(n1784) );
  DFFRX1 \I_cache/cache_reg[0][59]  ( .D(n12373), .CK(clk), .RN(n6080), .Q(
        \I_cache/cache[0][59] ), .QN(n1779) );
  DFFRX1 \I_cache/cache_reg[1][59]  ( .D(n12372), .CK(clk), .RN(n6080), .Q(
        \I_cache/cache[1][59] ), .QN(n3467) );
  DFFRX1 \I_cache/cache_reg[2][59]  ( .D(n12371), .CK(clk), .RN(n6080), .Q(
        \I_cache/cache[2][59] ), .QN(n1781) );
  DFFRX1 \I_cache/cache_reg[0][60]  ( .D(n12365), .CK(clk), .RN(n6080), .Q(
        \I_cache/cache[0][60] ), .QN(n1776) );
  DFFRX1 \I_cache/cache_reg[1][60]  ( .D(n12364), .CK(clk), .RN(n6080), .Q(
        \I_cache/cache[1][60] ), .QN(n3464) );
  DFFRX1 \I_cache/cache_reg[2][60]  ( .D(n12363), .CK(clk), .RN(n6080), .Q(
        \I_cache/cache[2][60] ), .QN(n1778) );
  DFFRX1 \I_cache/cache_reg[0][61]  ( .D(n12357), .CK(clk), .RN(n6079), .Q(
        \I_cache/cache[0][61] ), .QN(n1773) );
  DFFRX1 \I_cache/cache_reg[1][61]  ( .D(n12356), .CK(clk), .RN(n6079), .Q(
        \I_cache/cache[1][61] ), .QN(n3461) );
  DFFRX1 \I_cache/cache_reg[2][61]  ( .D(n12355), .CK(clk), .RN(n6079), .Q(
        \I_cache/cache[2][61] ), .QN(n1775) );
  DFFRX1 \I_cache/cache_reg[0][62]  ( .D(n12349), .CK(clk), .RN(n6078), .Q(
        \I_cache/cache[0][62] ), .QN(n1770) );
  DFFRX1 \I_cache/cache_reg[1][62]  ( .D(n12348), .CK(clk), .RN(n6078), .Q(
        \I_cache/cache[1][62] ), .QN(n3458) );
  DFFRX1 \I_cache/cache_reg[2][62]  ( .D(n12347), .CK(clk), .RN(n6078), .Q(
        \I_cache/cache[2][62] ), .QN(n1772) );
  DFFRX1 \I_cache/cache_reg[0][63]  ( .D(n12341), .CK(clk), .RN(n6078), .Q(
        \I_cache/cache[0][63] ), .QN(n1767) );
  DFFRX1 \I_cache/cache_reg[1][63]  ( .D(n12340), .CK(clk), .RN(n6078), .Q(
        \I_cache/cache[1][63] ), .QN(n3455) );
  DFFRX1 \I_cache/cache_reg[2][63]  ( .D(n12339), .CK(clk), .RN(n6078), .Q(
        \I_cache/cache[2][63] ), .QN(n1769) );
  DFFRX1 \I_cache/cache_reg[0][64]  ( .D(n12333), .CK(clk), .RN(n6077), .Q(
        \I_cache/cache[0][64] ), .QN(n1601) );
  DFFRX1 \I_cache/cache_reg[1][64]  ( .D(n12332), .CK(clk), .RN(n6077), .Q(
        \I_cache/cache[1][64] ), .QN(n3289) );
  DFFRX1 \I_cache/cache_reg[2][64]  ( .D(n12331), .CK(clk), .RN(n6077), .Q(
        \I_cache/cache[2][64] ), .QN(n1603) );
  DFFRX1 \I_cache/cache_reg[0][65]  ( .D(n12325), .CK(clk), .RN(n6076), .Q(
        \I_cache/cache[0][65] ), .QN(n221) );
  DFFRX1 \I_cache/cache_reg[1][65]  ( .D(n12324), .CK(clk), .RN(n6076), .Q(
        \I_cache/cache[1][65] ), .QN(n1850) );
  DFFRX1 \I_cache/cache_reg[2][65]  ( .D(n12323), .CK(clk), .RN(n6076), .Q(
        \I_cache/cache[2][65] ), .QN(n1673) );
  DFFRX1 \I_cache/cache_reg[0][66]  ( .D(n12317), .CK(clk), .RN(n6076), .Q(
        \I_cache/cache[0][66] ), .QN(n1669) );
  DFFRX1 \I_cache/cache_reg[1][66]  ( .D(n12316), .CK(clk), .RN(n6076), .Q(
        \I_cache/cache[1][66] ), .QN(n3358) );
  DFFRX1 \I_cache/cache_reg[2][66]  ( .D(n12315), .CK(clk), .RN(n6076), .Q(
        \I_cache/cache[2][66] ), .QN(n1671) );
  DFFRX1 \I_cache/cache_reg[0][67]  ( .D(n12309), .CK(clk), .RN(n6075), .Q(
        \I_cache/cache[0][67] ), .QN(n1666) );
  DFFRX1 \I_cache/cache_reg[1][67]  ( .D(n12308), .CK(clk), .RN(n6075), .Q(
        \I_cache/cache[1][67] ), .QN(n3355) );
  DFFRX1 \I_cache/cache_reg[2][67]  ( .D(n12307), .CK(clk), .RN(n6075), .Q(
        \I_cache/cache[2][67] ), .QN(n1668) );
  DFFRX1 \I_cache/cache_reg[0][68]  ( .D(n12301), .CK(clk), .RN(n6074), .Q(
        \I_cache/cache[0][68] ), .QN(n1663) );
  DFFRX1 \I_cache/cache_reg[1][68]  ( .D(n12300), .CK(clk), .RN(n6074), .Q(
        \I_cache/cache[1][68] ), .QN(n3352) );
  DFFRX1 \I_cache/cache_reg[2][68]  ( .D(n12299), .CK(clk), .RN(n6074), .Q(
        \I_cache/cache[2][68] ), .QN(n1665) );
  DFFRX1 \I_cache/cache_reg[0][69]  ( .D(n12293), .CK(clk), .RN(n6074), .Q(
        \I_cache/cache[0][69] ), .QN(n1660) );
  DFFRX1 \I_cache/cache_reg[1][69]  ( .D(n12292), .CK(clk), .RN(n6074), .Q(
        \I_cache/cache[1][69] ), .QN(n3349) );
  DFFRX1 \I_cache/cache_reg[2][69]  ( .D(n12291), .CK(clk), .RN(n6074), .Q(
        \I_cache/cache[2][69] ), .QN(n1662) );
  DFFRX1 \I_cache/cache_reg[0][70]  ( .D(n12285), .CK(clk), .RN(n6073), .Q(
        \I_cache/cache[0][70] ), .QN(n1657) );
  DFFRX1 \I_cache/cache_reg[1][70]  ( .D(n12284), .CK(clk), .RN(n6073), .Q(
        \I_cache/cache[1][70] ), .QN(n3346) );
  DFFRX1 \I_cache/cache_reg[2][70]  ( .D(n12283), .CK(clk), .RN(n6073), .Q(
        \I_cache/cache[2][70] ), .QN(n1659) );
  DFFRX1 \I_cache/cache_reg[0][71]  ( .D(n12277), .CK(clk), .RN(n6072), .Q(
        \I_cache/cache[0][71] ), .QN(n1654) );
  DFFRX1 \I_cache/cache_reg[1][71]  ( .D(n12276), .CK(clk), .RN(n6072), .Q(
        \I_cache/cache[1][71] ), .QN(n3343) );
  DFFRX1 \I_cache/cache_reg[2][71]  ( .D(n12275), .CK(clk), .RN(n6072), .Q(
        \I_cache/cache[2][71] ), .QN(n1656) );
  DFFRX1 \I_cache/cache_reg[0][72]  ( .D(n12269), .CK(clk), .RN(n6072), .Q(
        \I_cache/cache[0][72] ), .QN(n1651) );
  DFFRX1 \I_cache/cache_reg[1][72]  ( .D(n12268), .CK(clk), .RN(n6072), .Q(
        \I_cache/cache[1][72] ), .QN(n3340) );
  DFFRX1 \I_cache/cache_reg[2][72]  ( .D(n12267), .CK(clk), .RN(n6072), .Q(
        \I_cache/cache[2][72] ), .QN(n1653) );
  DFFRX1 \I_cache/cache_reg[0][73]  ( .D(n12261), .CK(clk), .RN(n6071), .Q(
        \I_cache/cache[0][73] ), .QN(n1648) );
  DFFRX1 \I_cache/cache_reg[1][73]  ( .D(n12260), .CK(clk), .RN(n6071), .Q(
        \I_cache/cache[1][73] ), .QN(n3337) );
  DFFRX1 \I_cache/cache_reg[2][73]  ( .D(n12259), .CK(clk), .RN(n6071), .Q(
        \I_cache/cache[2][73] ), .QN(n1650) );
  DFFRX1 \I_cache/cache_reg[0][74]  ( .D(n12253), .CK(clk), .RN(n6070), .Q(
        \I_cache/cache[0][74] ), .QN(n1645) );
  DFFRX1 \I_cache/cache_reg[1][74]  ( .D(n12252), .CK(clk), .RN(n6070), .Q(
        \I_cache/cache[1][74] ), .QN(n3334) );
  DFFRX1 \I_cache/cache_reg[2][74]  ( .D(n12251), .CK(clk), .RN(n6070), .Q(
        \I_cache/cache[2][74] ), .QN(n1647) );
  DFFRX1 \I_cache/cache_reg[0][75]  ( .D(n12245), .CK(clk), .RN(n6070), .Q(
        \I_cache/cache[0][75] ), .QN(n1642) );
  DFFRX1 \I_cache/cache_reg[1][75]  ( .D(n12244), .CK(clk), .RN(n6070), .Q(
        \I_cache/cache[1][75] ), .QN(n3331) );
  DFFRX1 \I_cache/cache_reg[2][75]  ( .D(n12243), .CK(clk), .RN(n6070), .Q(
        \I_cache/cache[2][75] ), .QN(n1644) );
  DFFRX1 \I_cache/cache_reg[0][76]  ( .D(n12237), .CK(clk), .RN(n6069), .Q(
        \I_cache/cache[0][76] ), .QN(n1639) );
  DFFRX1 \I_cache/cache_reg[1][76]  ( .D(n12236), .CK(clk), .RN(n6069), .Q(
        \I_cache/cache[1][76] ), .QN(n3328) );
  DFFRX1 \I_cache/cache_reg[2][76]  ( .D(n12235), .CK(clk), .RN(n6069), .Q(
        \I_cache/cache[2][76] ), .QN(n1641) );
  DFFRX1 \I_cache/cache_reg[0][77]  ( .D(n12229), .CK(clk), .RN(n6068), .Q(
        \I_cache/cache[0][77] ), .QN(n1636) );
  DFFRX1 \I_cache/cache_reg[1][77]  ( .D(n12228), .CK(clk), .RN(n6068), .Q(
        \I_cache/cache[1][77] ), .QN(n3325) );
  DFFRX1 \I_cache/cache_reg[2][77]  ( .D(n12227), .CK(clk), .RN(n6068), .Q(
        \I_cache/cache[2][77] ), .QN(n1638) );
  DFFRX1 \I_cache/cache_reg[0][78]  ( .D(n12221), .CK(clk), .RN(n6068), .Q(
        \I_cache/cache[0][78] ), .QN(n1633) );
  DFFRX1 \I_cache/cache_reg[1][78]  ( .D(n12220), .CK(clk), .RN(n6068), .Q(
        \I_cache/cache[1][78] ), .QN(n3322) );
  DFFRX1 \I_cache/cache_reg[2][78]  ( .D(n12219), .CK(clk), .RN(n6068), .Q(
        \I_cache/cache[2][78] ), .QN(n1635) );
  DFFRX1 \I_cache/cache_reg[0][79]  ( .D(n12213), .CK(clk), .RN(n6067), .Q(
        \I_cache/cache[0][79] ), .QN(n1630) );
  DFFRX1 \I_cache/cache_reg[1][79]  ( .D(n12212), .CK(clk), .RN(n6067), .Q(
        \I_cache/cache[1][79] ), .QN(n3319) );
  DFFRX1 \I_cache/cache_reg[2][79]  ( .D(n12211), .CK(clk), .RN(n6067), .Q(
        \I_cache/cache[2][79] ), .QN(n1632) );
  DFFRX1 \I_cache/cache_reg[0][80]  ( .D(n12205), .CK(clk), .RN(n6066), .Q(
        \I_cache/cache[0][80] ), .QN(n1346) );
  DFFRX1 \I_cache/cache_reg[1][80]  ( .D(n12204), .CK(clk), .RN(n6066), .Q(
        \I_cache/cache[1][80] ), .QN(n3316) );
  DFFRX1 \I_cache/cache_reg[2][80]  ( .D(n12203), .CK(clk), .RN(n6066), .Q(
        \I_cache/cache[2][80] ), .QN(n1629) );
  DFFRX1 \I_cache/cache_reg[0][81]  ( .D(n12197), .CK(clk), .RN(n6066), .Q(
        \I_cache/cache[0][81] ), .QN(n1625) );
  DFFRX1 \I_cache/cache_reg[1][81]  ( .D(n12196), .CK(clk), .RN(n6066), .Q(
        \I_cache/cache[1][81] ), .QN(n3313) );
  DFFRX1 \I_cache/cache_reg[2][81]  ( .D(n12195), .CK(clk), .RN(n6066), .Q(
        \I_cache/cache[2][81] ), .QN(n1627) );
  DFFRX1 \I_cache/cache_reg[0][82]  ( .D(n12189), .CK(clk), .RN(n6065), .Q(
        \I_cache/cache[0][82] ), .QN(n1622) );
  DFFRX1 \I_cache/cache_reg[1][82]  ( .D(n12188), .CK(clk), .RN(n6065), .Q(
        \I_cache/cache[1][82] ), .QN(n3310) );
  DFFRX1 \I_cache/cache_reg[2][82]  ( .D(n12187), .CK(clk), .RN(n6065), .Q(
        \I_cache/cache[2][82] ), .QN(n1624) );
  DFFRX1 \I_cache/cache_reg[0][83]  ( .D(n12181), .CK(clk), .RN(n6064), .Q(
        \I_cache/cache[0][83] ), .QN(n1847) );
  DFFRX1 \I_cache/cache_reg[1][83]  ( .D(n12180), .CK(clk), .RN(n6064), .Q(
        \I_cache/cache[1][83] ), .QN(n3535) );
  DFFRX1 \I_cache/cache_reg[2][83]  ( .D(n12179), .CK(clk), .RN(n6064), .Q(
        \I_cache/cache[2][83] ), .QN(n1849) );
  DFFRX1 \I_cache/cache_reg[0][84]  ( .D(n12173), .CK(clk), .RN(n6064), .Q(
        \I_cache/cache[0][84] ), .QN(n1619) );
  DFFRX1 \I_cache/cache_reg[1][84]  ( .D(n12172), .CK(clk), .RN(n6064), .Q(
        \I_cache/cache[1][84] ), .QN(n3307) );
  DFFRX1 \I_cache/cache_reg[2][84]  ( .D(n12171), .CK(clk), .RN(n6064), .Q(
        \I_cache/cache[2][84] ), .QN(n1621) );
  DFFRX1 \I_cache/cache_reg[0][85]  ( .D(n12165), .CK(clk), .RN(n6063), .Q(
        \I_cache/cache[0][85] ), .QN(n1616) );
  DFFRX1 \I_cache/cache_reg[1][85]  ( .D(n12164), .CK(clk), .RN(n6063), .Q(
        \I_cache/cache[1][85] ), .QN(n3304) );
  DFFRX1 \I_cache/cache_reg[2][85]  ( .D(n12163), .CK(clk), .RN(n6063), .Q(
        \I_cache/cache[2][85] ), .QN(n1618) );
  DFFRX1 \I_cache/cache_reg[0][86]  ( .D(n12157), .CK(clk), .RN(n6062), .Q(
        \I_cache/cache[0][86] ), .QN(n1613) );
  DFFRX1 \I_cache/cache_reg[1][86]  ( .D(n12156), .CK(clk), .RN(n6062), .Q(
        \I_cache/cache[1][86] ), .QN(n3301) );
  DFFRX1 \I_cache/cache_reg[2][86]  ( .D(n12155), .CK(clk), .RN(n6062), .Q(
        \I_cache/cache[2][86] ), .QN(n1615) );
  DFFRX1 \I_cache/cache_reg[0][87]  ( .D(n12149), .CK(clk), .RN(n6062), .Q(
        \I_cache/cache[0][87] ), .QN(n1610) );
  DFFRX1 \I_cache/cache_reg[1][87]  ( .D(n12148), .CK(clk), .RN(n6062), .Q(
        \I_cache/cache[1][87] ), .QN(n3298) );
  DFFRX1 \I_cache/cache_reg[2][87]  ( .D(n12147), .CK(clk), .RN(n6062), .Q(
        \I_cache/cache[2][87] ), .QN(n1612) );
  DFFRX1 \I_cache/cache_reg[0][88]  ( .D(n12141), .CK(clk), .RN(n6061), .Q(
        \I_cache/cache[0][88] ), .QN(n1607) );
  DFFRX1 \I_cache/cache_reg[1][88]  ( .D(n12140), .CK(clk), .RN(n6061), .Q(
        \I_cache/cache[1][88] ), .QN(n3295) );
  DFFRX1 \I_cache/cache_reg[2][88]  ( .D(n12139), .CK(clk), .RN(n6061), .Q(
        \I_cache/cache[2][88] ), .QN(n1609) );
  DFFRX1 \I_cache/cache_reg[0][89]  ( .D(n12133), .CK(clk), .RN(n6060), .Q(
        \I_cache/cache[0][89] ), .QN(n1604) );
  DFFRX1 \I_cache/cache_reg[1][89]  ( .D(n12132), .CK(clk), .RN(n6060), .Q(
        \I_cache/cache[1][89] ), .QN(n3292) );
  DFFRX1 \I_cache/cache_reg[2][89]  ( .D(n12131), .CK(clk), .RN(n6060), .Q(
        \I_cache/cache[2][89] ), .QN(n1606) );
  DFFRX1 \I_cache/cache_reg[0][90]  ( .D(n12125), .CK(clk), .RN(n6060), .Q(
        \I_cache/cache[0][90] ), .QN(n1689) );
  DFFRX1 \I_cache/cache_reg[1][90]  ( .D(n12124), .CK(clk), .RN(n6060), .Q(
        \I_cache/cache[1][90] ), .QN(n3377) );
  DFFRX1 \I_cache/cache_reg[2][90]  ( .D(n12123), .CK(clk), .RN(n6060), .Q(
        \I_cache/cache[2][90] ), .QN(n1691) );
  DFFRX1 \I_cache/cache_reg[0][91]  ( .D(n12117), .CK(clk), .RN(n6059), .Q(
        \I_cache/cache[0][91] ), .QN(n1686) );
  DFFRX1 \I_cache/cache_reg[1][91]  ( .D(n12116), .CK(clk), .RN(n6059), .Q(
        \I_cache/cache[1][91] ), .QN(n3374) );
  DFFRX1 \I_cache/cache_reg[2][91]  ( .D(n12115), .CK(clk), .RN(n6059), .Q(
        \I_cache/cache[2][91] ), .QN(n1688) );
  DFFRX1 \I_cache/cache_reg[0][92]  ( .D(n12109), .CK(clk), .RN(n6058), .Q(
        \I_cache/cache[0][92] ), .QN(n1683) );
  DFFRX1 \I_cache/cache_reg[1][92]  ( .D(n12108), .CK(clk), .RN(n6058), .Q(
        \I_cache/cache[1][92] ), .QN(n3371) );
  DFFRX1 \I_cache/cache_reg[2][92]  ( .D(n12107), .CK(clk), .RN(n6058), .Q(
        \I_cache/cache[2][92] ), .QN(n1685) );
  DFFRX1 \I_cache/cache_reg[0][93]  ( .D(n12101), .CK(clk), .RN(n6058), .Q(
        \I_cache/cache[0][93] ), .QN(n1680) );
  DFFRX1 \I_cache/cache_reg[1][93]  ( .D(n12100), .CK(clk), .RN(n6058), .Q(
        \I_cache/cache[1][93] ), .QN(n3368) );
  DFFRX1 \I_cache/cache_reg[2][93]  ( .D(n12099), .CK(clk), .RN(n6058), .Q(
        \I_cache/cache[2][93] ), .QN(n1682) );
  DFFRX1 \I_cache/cache_reg[0][94]  ( .D(n12093), .CK(clk), .RN(n6057), .Q(
        \I_cache/cache[0][94] ), .QN(n1677) );
  DFFRX1 \I_cache/cache_reg[1][94]  ( .D(n12092), .CK(clk), .RN(n6057), .Q(
        \I_cache/cache[1][94] ), .QN(n3365) );
  DFFRX1 \I_cache/cache_reg[2][94]  ( .D(n12091), .CK(clk), .RN(n6057), .Q(
        \I_cache/cache[2][94] ), .QN(n1679) );
  DFFRX1 \I_cache/cache_reg[0][95]  ( .D(n12085), .CK(clk), .RN(n6056), .Q(
        \I_cache/cache[0][95] ), .QN(n1674) );
  DFFRX1 \I_cache/cache_reg[1][95]  ( .D(n12084), .CK(clk), .RN(n6056), .Q(
        \I_cache/cache[1][95] ), .QN(n3362) );
  DFFRX1 \I_cache/cache_reg[2][95]  ( .D(n12083), .CK(clk), .RN(n6056), .Q(
        \I_cache/cache[2][95] ), .QN(n1676) );
  DFFRX1 \I_cache/cache_reg[0][96]  ( .D(n12077), .CK(clk), .RN(n6056), .Q(
        \I_cache/cache[0][96] ), .QN(n1347) );
  DFFRX1 \I_cache/cache_reg[1][96]  ( .D(n12076), .CK(clk), .RN(n6056), .Q(
        \I_cache/cache[1][96] ), .QN(n3034) );
  DFFRX1 \I_cache/cache_reg[2][96]  ( .D(n12075), .CK(clk), .RN(n6056), .Q(
        \I_cache/cache[2][96] ), .QN(n1349) );
  DFFRX1 \I_cache/cache_reg[0][97]  ( .D(n12069), .CK(clk), .RN(n6055), .Q(
        \I_cache/cache[0][97] ), .QN(n1418) );
  DFFRX1 \I_cache/cache_reg[1][97]  ( .D(n12068), .CK(clk), .RN(n6055), .Q(
        \I_cache/cache[1][97] ), .QN(n3105) );
  DFFRX1 \I_cache/cache_reg[2][97]  ( .D(n12067), .CK(clk), .RN(n6055), .Q(
        \I_cache/cache[2][97] ), .QN(n1420) );
  DFFRX1 \I_cache/cache_reg[0][98]  ( .D(n12061), .CK(clk), .RN(n6054), .Q(
        \I_cache/cache[0][98] ), .QN(n1415) );
  DFFRX1 \I_cache/cache_reg[1][98]  ( .D(n12060), .CK(clk), .RN(n6054), .Q(
        \I_cache/cache[1][98] ), .QN(n3102) );
  DFFRX1 \I_cache/cache_reg[2][98]  ( .D(n12059), .CK(clk), .RN(n6054), .Q(
        \I_cache/cache[2][98] ), .QN(n1417) );
  DFFRX1 \I_cache/cache_reg[0][99]  ( .D(n12053), .CK(clk), .RN(n6054), .Q(
        \I_cache/cache[0][99] ), .QN(n1412) );
  DFFRX1 \I_cache/cache_reg[1][99]  ( .D(n12052), .CK(clk), .RN(n6054), .Q(
        \I_cache/cache[1][99] ), .QN(n3099) );
  DFFRX1 \I_cache/cache_reg[2][99]  ( .D(n12051), .CK(clk), .RN(n6054), .Q(
        \I_cache/cache[2][99] ), .QN(n1414) );
  DFFRX1 \I_cache/cache_reg[0][100]  ( .D(n12045), .CK(clk), .RN(n6053), .Q(
        \I_cache/cache[0][100] ), .QN(n1409) );
  DFFRX1 \I_cache/cache_reg[1][100]  ( .D(n12044), .CK(clk), .RN(n6053), .Q(
        \I_cache/cache[1][100] ), .QN(n3096) );
  DFFRX1 \I_cache/cache_reg[2][100]  ( .D(n12043), .CK(clk), .RN(n6053), .Q(
        \I_cache/cache[2][100] ), .QN(n1411) );
  DFFRX1 \I_cache/cache_reg[0][101]  ( .D(n12037), .CK(clk), .RN(n6052), .Q(
        \I_cache/cache[0][101] ), .QN(n1406) );
  DFFRX1 \I_cache/cache_reg[1][101]  ( .D(n12036), .CK(clk), .RN(n6052), .Q(
        \I_cache/cache[1][101] ), .QN(n3093) );
  DFFRX1 \I_cache/cache_reg[2][101]  ( .D(n12035), .CK(clk), .RN(n6052), .Q(
        \I_cache/cache[2][101] ), .QN(n1408) );
  DFFRX1 \I_cache/cache_reg[0][102]  ( .D(n12029), .CK(clk), .RN(n6052), .Q(
        \I_cache/cache[0][102] ), .QN(n1403) );
  DFFRX1 \I_cache/cache_reg[1][102]  ( .D(n12028), .CK(clk), .RN(n6052), .Q(
        \I_cache/cache[1][102] ), .QN(n3090) );
  DFFRX1 \I_cache/cache_reg[2][102]  ( .D(n12027), .CK(clk), .RN(n6052), .Q(
        \I_cache/cache[2][102] ), .QN(n1405) );
  DFFRX1 \I_cache/cache_reg[0][103]  ( .D(n12021), .CK(clk), .RN(n6051), .Q(
        \I_cache/cache[0][103] ), .QN(n1400) );
  DFFRX1 \I_cache/cache_reg[1][103]  ( .D(n12020), .CK(clk), .RN(n6051), .Q(
        \I_cache/cache[1][103] ), .QN(n3087) );
  DFFRX1 \I_cache/cache_reg[2][103]  ( .D(n12019), .CK(clk), .RN(n6051), .Q(
        \I_cache/cache[2][103] ), .QN(n1402) );
  DFFRX1 \I_cache/cache_reg[0][104]  ( .D(n12013), .CK(clk), .RN(n6050), .Q(
        \I_cache/cache[0][104] ), .QN(n1397) );
  DFFRX1 \I_cache/cache_reg[1][104]  ( .D(n12012), .CK(clk), .RN(n6050), .Q(
        \I_cache/cache[1][104] ), .QN(n3084) );
  DFFRX1 \I_cache/cache_reg[2][104]  ( .D(n12011), .CK(clk), .RN(n6050), .Q(
        \I_cache/cache[2][104] ), .QN(n1399) );
  DFFRX1 \I_cache/cache_reg[0][105]  ( .D(n12005), .CK(clk), .RN(n6050), .Q(
        \I_cache/cache[0][105] ), .QN(n1394) );
  DFFRX1 \I_cache/cache_reg[1][105]  ( .D(n12004), .CK(clk), .RN(n6050), .Q(
        \I_cache/cache[1][105] ), .QN(n3081) );
  DFFRX1 \I_cache/cache_reg[2][105]  ( .D(n12003), .CK(clk), .RN(n6050), .Q(
        \I_cache/cache[2][105] ), .QN(n1396) );
  DFFRX1 \I_cache/cache_reg[0][106]  ( .D(n11997), .CK(clk), .RN(n6049), .Q(
        \I_cache/cache[0][106] ), .QN(n1391) );
  DFFRX1 \I_cache/cache_reg[1][106]  ( .D(n11996), .CK(clk), .RN(n6049), .Q(
        \I_cache/cache[1][106] ), .QN(n3078) );
  DFFRX1 \I_cache/cache_reg[2][106]  ( .D(n11995), .CK(clk), .RN(n6049), .Q(
        \I_cache/cache[2][106] ), .QN(n1393) );
  DFFRX1 \I_cache/cache_reg[0][107]  ( .D(n11989), .CK(clk), .RN(n6048), .Q(
        \I_cache/cache[0][107] ), .QN(n1388) );
  DFFRX1 \I_cache/cache_reg[1][107]  ( .D(n11988), .CK(clk), .RN(n6048), .Q(
        \I_cache/cache[1][107] ), .QN(n3075) );
  DFFRX1 \I_cache/cache_reg[2][107]  ( .D(n11987), .CK(clk), .RN(n6048), .Q(
        \I_cache/cache[2][107] ), .QN(n1390) );
  DFFRX1 \I_cache/cache_reg[0][108]  ( .D(n11981), .CK(clk), .RN(n6048), .Q(
        \I_cache/cache[0][108] ), .QN(n1385) );
  DFFRX1 \I_cache/cache_reg[1][108]  ( .D(n11980), .CK(clk), .RN(n6048), .Q(
        \I_cache/cache[1][108] ), .QN(n3072) );
  DFFRX1 \I_cache/cache_reg[2][108]  ( .D(n11979), .CK(clk), .RN(n6048), .Q(
        \I_cache/cache[2][108] ), .QN(n1387) );
  DFFRX1 \I_cache/cache_reg[0][109]  ( .D(n11973), .CK(clk), .RN(n6047), .Q(
        \I_cache/cache[0][109] ), .QN(n1382) );
  DFFRX1 \I_cache/cache_reg[1][109]  ( .D(n11972), .CK(clk), .RN(n6047), .Q(
        \I_cache/cache[1][109] ), .QN(n3069) );
  DFFRX1 \I_cache/cache_reg[2][109]  ( .D(n11971), .CK(clk), .RN(n6047), .Q(
        \I_cache/cache[2][109] ), .QN(n1384) );
  DFFRX1 \I_cache/cache_reg[0][110]  ( .D(n11965), .CK(clk), .RN(n6046), .Q(
        \I_cache/cache[0][110] ), .QN(n1379) );
  DFFRX1 \I_cache/cache_reg[1][110]  ( .D(n11964), .CK(clk), .RN(n6046), .Q(
        \I_cache/cache[1][110] ), .QN(n3066) );
  DFFRX1 \I_cache/cache_reg[2][110]  ( .D(n11963), .CK(clk), .RN(n6046), .Q(
        \I_cache/cache[2][110] ), .QN(n1381) );
  DFFRX1 \I_cache/cache_reg[0][111]  ( .D(n11957), .CK(clk), .RN(n6046), .Q(
        \I_cache/cache[0][111] ), .QN(n1376) );
  DFFRX1 \I_cache/cache_reg[1][111]  ( .D(n11956), .CK(clk), .RN(n6046), .Q(
        \I_cache/cache[1][111] ), .QN(n3063) );
  DFFRX1 \I_cache/cache_reg[2][111]  ( .D(n11955), .CK(clk), .RN(n6046), .Q(
        \I_cache/cache[2][111] ), .QN(n1378) );
  DFFRX1 \I_cache/cache_reg[0][112]  ( .D(n11949), .CK(clk), .RN(n6045), .Q(
        \I_cache/cache[0][112] ), .QN(n1373) );
  DFFRX1 \I_cache/cache_reg[1][112]  ( .D(n11948), .CK(clk), .RN(n6045), .Q(
        \I_cache/cache[1][112] ), .QN(n3060) );
  DFFRX1 \I_cache/cache_reg[2][112]  ( .D(n11947), .CK(clk), .RN(n6045), .Q(
        \I_cache/cache[2][112] ), .QN(n1375) );
  DFFRX1 \I_cache/cache_reg[0][113]  ( .D(n11941), .CK(clk), .RN(n6044), .Q(
        \I_cache/cache[0][113] ), .QN(n3033) );
  DFFRX1 \I_cache/cache_reg[1][113]  ( .D(n11940), .CK(clk), .RN(n6044), .Q(
        \I_cache/cache[1][113] ), .QN(n1345) );
  DFFRX1 \I_cache/cache_reg[2][113]  ( .D(n11939), .CK(clk), .RN(n6044), .Q(
        \I_cache/cache[2][113] ), .QN(n1372) );
  DFFRX1 \I_cache/cache_reg[0][114]  ( .D(n11933), .CK(clk), .RN(n6044), .Q(
        \I_cache/cache[0][114] ), .QN(n1368) );
  DFFRX1 \I_cache/cache_reg[1][114]  ( .D(n11932), .CK(clk), .RN(n6044), .Q(
        \I_cache/cache[1][114] ), .QN(n3055) );
  DFFRX1 \I_cache/cache_reg[2][114]  ( .D(n11931), .CK(clk), .RN(n6044), .Q(
        \I_cache/cache[2][114] ), .QN(n1370) );
  DFFRX1 \I_cache/cache_reg[0][115]  ( .D(n11925), .CK(clk), .RN(n6043), .Q(
        \I_cache/cache[0][115] ), .QN(n1593) );
  DFFRX1 \I_cache/cache_reg[1][115]  ( .D(n11924), .CK(clk), .RN(n6043), .Q(
        \I_cache/cache[1][115] ), .QN(n3280) );
  DFFRX1 \I_cache/cache_reg[2][115]  ( .D(n11923), .CK(clk), .RN(n6043), .Q(
        \I_cache/cache[2][115] ), .QN(n1595) );
  DFFRX1 \I_cache/cache_reg[0][116]  ( .D(n11917), .CK(clk), .RN(n6042), .Q(
        \I_cache/cache[0][116] ), .QN(n1365) );
  DFFRX1 \I_cache/cache_reg[1][116]  ( .D(n11916), .CK(clk), .RN(n6042), .Q(
        \I_cache/cache[1][116] ), .QN(n3052) );
  DFFRX1 \I_cache/cache_reg[2][116]  ( .D(n11915), .CK(clk), .RN(n6042), .Q(
        \I_cache/cache[2][116] ), .QN(n1367) );
  DFFRX1 \I_cache/cache_reg[0][117]  ( .D(n11909), .CK(clk), .RN(n6042), .Q(
        \I_cache/cache[0][117] ), .QN(n1362) );
  DFFRX1 \I_cache/cache_reg[1][117]  ( .D(n11908), .CK(clk), .RN(n6042), .Q(
        \I_cache/cache[1][117] ), .QN(n3049) );
  DFFRX1 \I_cache/cache_reg[2][117]  ( .D(n11907), .CK(clk), .RN(n6042), .Q(
        \I_cache/cache[2][117] ), .QN(n1364) );
  DFFRX1 \I_cache/cache_reg[0][118]  ( .D(n11901), .CK(clk), .RN(n6041), .Q(
        \I_cache/cache[0][118] ), .QN(n1359) );
  DFFRX1 \I_cache/cache_reg[1][118]  ( .D(n11900), .CK(clk), .RN(n6041), .Q(
        \I_cache/cache[1][118] ), .QN(n3046) );
  DFFRX1 \I_cache/cache_reg[2][118]  ( .D(n11899), .CK(clk), .RN(n6041), .Q(
        \I_cache/cache[2][118] ), .QN(n1361) );
  DFFRX1 \I_cache/cache_reg[0][119]  ( .D(n11893), .CK(clk), .RN(n6040), .Q(
        \I_cache/cache[0][119] ), .QN(n1356) );
  DFFRX1 \I_cache/cache_reg[1][119]  ( .D(n11892), .CK(clk), .RN(n6040), .Q(
        \I_cache/cache[1][119] ), .QN(n3043) );
  DFFRX1 \I_cache/cache_reg[2][119]  ( .D(n11891), .CK(clk), .RN(n6040), .Q(
        \I_cache/cache[2][119] ), .QN(n1358) );
  DFFRX1 \I_cache/cache_reg[0][120]  ( .D(n11885), .CK(clk), .RN(n6040), .Q(
        \I_cache/cache[0][120] ), .QN(n1353) );
  DFFRX1 \I_cache/cache_reg[1][120]  ( .D(n11884), .CK(clk), .RN(n6040), .Q(
        \I_cache/cache[1][120] ), .QN(n3040) );
  DFFRX1 \I_cache/cache_reg[2][120]  ( .D(n11883), .CK(clk), .RN(n6040), .Q(
        \I_cache/cache[2][120] ), .QN(n1355) );
  DFFRX1 \I_cache/cache_reg[0][121]  ( .D(n11877), .CK(clk), .RN(n6039), .Q(
        \I_cache/cache[0][121] ), .QN(n1350) );
  DFFRX1 \I_cache/cache_reg[1][121]  ( .D(n11876), .CK(clk), .RN(n6039), .Q(
        \I_cache/cache[1][121] ), .QN(n3037) );
  DFFRX1 \I_cache/cache_reg[2][121]  ( .D(n11875), .CK(clk), .RN(n6039), .Q(
        \I_cache/cache[2][121] ), .QN(n1352) );
  DFFRX1 \I_cache/cache_reg[0][122]  ( .D(n11869), .CK(clk), .RN(n6038), .Q(
        \I_cache/cache[0][122] ), .QN(n1436) );
  DFFRX1 \I_cache/cache_reg[1][122]  ( .D(n11868), .CK(clk), .RN(n6038), .Q(
        \I_cache/cache[1][122] ), .QN(n3123) );
  DFFRX1 \I_cache/cache_reg[2][122]  ( .D(n11867), .CK(clk), .RN(n6038), .Q(
        \I_cache/cache[2][122] ), .QN(n1438) );
  DFFRX1 \I_cache/cache_reg[0][123]  ( .D(n11861), .CK(clk), .RN(n6038), .Q(
        \I_cache/cache[0][123] ), .QN(n1433) );
  DFFRX1 \I_cache/cache_reg[1][123]  ( .D(n11860), .CK(clk), .RN(n6038), .Q(
        \I_cache/cache[1][123] ), .QN(n3120) );
  DFFRX1 \I_cache/cache_reg[2][123]  ( .D(n11859), .CK(clk), .RN(n6038), .Q(
        \I_cache/cache[2][123] ), .QN(n1435) );
  DFFRX1 \I_cache/cache_reg[0][124]  ( .D(n11853), .CK(clk), .RN(n6037), .Q(
        \I_cache/cache[0][124] ), .QN(n1430) );
  DFFRX1 \I_cache/cache_reg[1][124]  ( .D(n11852), .CK(clk), .RN(n6037), .Q(
        \I_cache/cache[1][124] ), .QN(n3117) );
  DFFRX1 \I_cache/cache_reg[2][124]  ( .D(n11851), .CK(clk), .RN(n6037), .Q(
        \I_cache/cache[2][124] ), .QN(n1432) );
  DFFRX1 \I_cache/cache_reg[0][125]  ( .D(n11845), .CK(clk), .RN(n6036), .Q(
        \I_cache/cache[0][125] ), .QN(n1427) );
  DFFRX1 \I_cache/cache_reg[1][125]  ( .D(n11844), .CK(clk), .RN(n6036), .Q(
        \I_cache/cache[1][125] ), .QN(n3114) );
  DFFRX1 \I_cache/cache_reg[2][125]  ( .D(n11843), .CK(clk), .RN(n6036), .Q(
        \I_cache/cache[2][125] ), .QN(n1429) );
  DFFRX1 \I_cache/cache_reg[0][126]  ( .D(n11837), .CK(clk), .RN(n6036), .Q(
        \I_cache/cache[0][126] ), .QN(n1424) );
  DFFRX1 \I_cache/cache_reg[1][126]  ( .D(n11836), .CK(clk), .RN(n6036), .Q(
        \I_cache/cache[1][126] ), .QN(n3111) );
  DFFRX1 \I_cache/cache_reg[2][126]  ( .D(n11835), .CK(clk), .RN(n6036), .Q(
        \I_cache/cache[2][126] ), .QN(n1426) );
  DFFRX1 \I_cache/cache_reg[0][127]  ( .D(n11829), .CK(clk), .RN(n6035), .Q(
        \I_cache/cache[0][127] ), .QN(n1421) );
  DFFRX1 \I_cache/cache_reg[1][127]  ( .D(n11828), .CK(clk), .RN(n6035), .Q(
        \I_cache/cache[1][127] ), .QN(n3108) );
  DFFRX1 \I_cache/cache_reg[2][127]  ( .D(n11827), .CK(clk), .RN(n6035), .Q(
        \I_cache/cache[2][127] ), .QN(n1423) );
  DFFRX1 \i_MIPS/Register/register_reg[30][14]  ( .D(\i_MIPS/Register/n162 ), 
        .CK(clk), .RN(n6305), .Q(\i_MIPS/Register/register[30][14] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][30]  ( .D(\i_MIPS/Register/n178 ), 
        .CK(clk), .RN(n6303), .Q(\i_MIPS/Register/register[30][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][31]  ( .D(\i_MIPS/Register/n179 ), 
        .CK(clk), .RN(n6303), .Q(\i_MIPS/Register/register[30][31] ) );
  DFFRX1 \i_MIPS/Register/register_reg[28][14]  ( .D(\i_MIPS/Register/n226 ), 
        .CK(clk), .RN(n6299), .Q(\i_MIPS/Register/register[28][14] ) );
  DFFRX1 \i_MIPS/Register/register_reg[28][30]  ( .D(\i_MIPS/Register/n242 ), 
        .CK(clk), .RN(n6298), .Q(\i_MIPS/Register/register[28][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[28][31]  ( .D(\i_MIPS/Register/n243 ), 
        .CK(clk), .RN(n6298), .Q(\i_MIPS/Register/register[28][31] ) );
  DFFRX1 \i_MIPS/Register/register_reg[24][14]  ( .D(\i_MIPS/Register/n354 ), 
        .CK(clk), .RN(n6289), .Q(\i_MIPS/Register/register[24][14] ) );
  DFFRX1 \i_MIPS/Register/register_reg[24][30]  ( .D(\i_MIPS/Register/n370 ), 
        .CK(clk), .RN(n6287), .Q(\i_MIPS/Register/register[24][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[24][31]  ( .D(\i_MIPS/Register/n371 ), 
        .CK(clk), .RN(n6287), .Q(\i_MIPS/Register/register[24][31] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][14]  ( .D(\i_MIPS/Register/n674 ), 
        .CK(clk), .RN(n6262), .Q(\i_MIPS/Register/register[14][14] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][30]  ( .D(\i_MIPS/Register/n690 ), 
        .CK(clk), .RN(n6261), .Q(\i_MIPS/Register/register[14][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][31]  ( .D(\i_MIPS/Register/n691 ), 
        .CK(clk), .RN(n6261), .Q(\i_MIPS/Register/register[14][31] ) );
  DFFRX1 \i_MIPS/Register/register_reg[12][14]  ( .D(\i_MIPS/Register/n738 ), 
        .CK(clk), .RN(n6257), .Q(\i_MIPS/Register/register[12][14] ) );
  DFFRX1 \i_MIPS/Register/register_reg[12][30]  ( .D(\i_MIPS/Register/n754 ), 
        .CK(clk), .RN(n6255), .Q(\i_MIPS/Register/register[12][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[12][31]  ( .D(\i_MIPS/Register/n755 ), 
        .CK(clk), .RN(n6255), .Q(\i_MIPS/Register/register[12][31] ) );
  DFFRX1 \i_MIPS/Register/register_reg[8][14]  ( .D(\i_MIPS/Register/n866 ), 
        .CK(clk), .RN(n6246), .Q(\i_MIPS/Register/register[8][14] ) );
  DFFRX1 \i_MIPS/Register/register_reg[8][30]  ( .D(\i_MIPS/Register/n882 ), 
        .CK(clk), .RN(n6245), .Q(\i_MIPS/Register/register[8][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[8][31]  ( .D(\i_MIPS/Register/n883 ), 
        .CK(clk), .RN(n6245), .Q(\i_MIPS/Register/register[8][31] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][14]  ( .D(\i_MIPS/Register/n418 ), 
        .CK(clk), .RN(n6283), .Q(\i_MIPS/Register/register[22][14] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][15]  ( .D(\i_MIPS/Register/n419 ), 
        .CK(clk), .RN(n6283), .Q(\i_MIPS/Register/register[22][15] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][25]  ( .D(\i_MIPS/Register/n429 ), 
        .CK(clk), .RN(n6282), .Q(\i_MIPS/Register/register[22][25] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][30]  ( .D(\i_MIPS/Register/n434 ), 
        .CK(clk), .RN(n6282), .Q(\i_MIPS/Register/register[22][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][31]  ( .D(\i_MIPS/Register/n435 ), 
        .CK(clk), .RN(n6282), .Q(\i_MIPS/Register/register[22][31] ) );
  DFFRX1 \i_MIPS/Register/register_reg[21][22]  ( .D(\i_MIPS/Register/n458 ), 
        .CK(clk), .RN(n6280), .Q(\i_MIPS/Register/register[21][22] ) );
  DFFRX1 \i_MIPS/Register/register_reg[20][14]  ( .D(\i_MIPS/Register/n482 ), 
        .CK(clk), .RN(n6278), .Q(\i_MIPS/Register/register[20][14] ) );
  DFFRX1 \i_MIPS/Register/register_reg[20][30]  ( .D(\i_MIPS/Register/n498 ), 
        .CK(clk), .RN(n6277), .Q(\i_MIPS/Register/register[20][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[20][31]  ( .D(\i_MIPS/Register/n499 ), 
        .CK(clk), .RN(n6277), .Q(\i_MIPS/Register/register[20][31] ) );
  DFFRX1 \i_MIPS/Register/register_reg[19][22]  ( .D(\i_MIPS/Register/n522 ), 
        .CK(clk), .RN(n6275), .Q(\i_MIPS/Register/register[19][22] ) );
  DFFRX1 \i_MIPS/Register/register_reg[17][22]  ( .D(\i_MIPS/Register/n586 ), 
        .CK(clk), .RN(n6269), .Q(\i_MIPS/Register/register[17][22] ) );
  DFFRX1 \i_MIPS/Register/register_reg[16][14]  ( .D(\i_MIPS/Register/n610 ), 
        .CK(clk), .RN(n6267), .Q(\i_MIPS/Register/register[16][14] ) );
  DFFRX1 \i_MIPS/Register/register_reg[16][30]  ( .D(\i_MIPS/Register/n626 ), 
        .CK(clk), .RN(n6266), .Q(\i_MIPS/Register/register[16][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[16][31]  ( .D(\i_MIPS/Register/n627 ), 
        .CK(clk), .RN(n6266), .Q(\i_MIPS/Register/register[16][31] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][14]  ( .D(\i_MIPS/Register/n930 ), 
        .CK(clk), .RN(n6241), .Q(\i_MIPS/Register/register[6][14] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][15]  ( .D(\i_MIPS/Register/n931 ), 
        .CK(clk), .RN(n6241), .Q(\i_MIPS/Register/register[6][15] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][25]  ( .D(\i_MIPS/Register/n941 ), 
        .CK(clk), .RN(n6240), .Q(\i_MIPS/Register/register[6][25] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][30]  ( .D(\i_MIPS/Register/n946 ), 
        .CK(clk), .RN(n6239), .Q(\i_MIPS/Register/register[6][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][31]  ( .D(\i_MIPS/Register/n947 ), 
        .CK(clk), .RN(n6239), .Q(\i_MIPS/Register/register[6][31] ) );
  DFFRX1 \i_MIPS/Register/register_reg[5][22]  ( .D(\i_MIPS/Register/n970 ), 
        .CK(clk), .RN(n6237), .Q(\i_MIPS/Register/register[5][22] ) );
  DFFRX1 \i_MIPS/Register/register_reg[4][14]  ( .D(\i_MIPS/Register/n994 ), 
        .CK(clk), .RN(n6235), .Q(\i_MIPS/Register/register[4][14] ) );
  DFFRX1 \i_MIPS/Register/register_reg[4][30]  ( .D(\i_MIPS/Register/n1010 ), 
        .CK(clk), .RN(n6234), .Q(\i_MIPS/Register/register[4][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[4][31]  ( .D(\i_MIPS/Register/n1011 ), 
        .CK(clk), .RN(n6234), .Q(\i_MIPS/Register/register[4][31] ) );
  DFFRX1 \i_MIPS/Register/register_reg[3][22]  ( .D(\i_MIPS/Register/n1034 ), 
        .CK(clk), .RN(n6232), .Q(\i_MIPS/Register/register[3][22] ) );
  DFFRX1 \i_MIPS/Register/register_reg[1][22]  ( .D(\i_MIPS/Register/n1098 ), 
        .CK(clk), .RN(n6227), .Q(\i_MIPS/Register/register[1][22] ) );
  DFFRX1 \i_MIPS/Register/register_reg[0][14]  ( .D(\i_MIPS/Register/n1122 ), 
        .CK(clk), .RN(n6225), .Q(\i_MIPS/Register/register[0][14] ) );
  DFFRX1 \i_MIPS/Register/register_reg[0][30]  ( .D(\i_MIPS/Register/n1138 ), 
        .CK(clk), .RN(n6223), .Q(\i_MIPS/Register/register[0][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[0][31]  ( .D(\i_MIPS/Register/n1139 ), 
        .CK(clk), .RN(n6223), .Q(\i_MIPS/Register/register[0][31] ) );
  DFFRX1 \i_MIPS/Register/register_reg[28][2]  ( .D(\i_MIPS/Register/n214 ), 
        .CK(clk), .RN(n6300), .Q(\i_MIPS/Register/register[28][2] ), .QN(n287)
         );
  DFFRX1 \i_MIPS/Register/register_reg[28][15]  ( .D(\i_MIPS/Register/n227 ), 
        .CK(clk), .RN(n6299), .Q(\i_MIPS/Register/register[28][15] ), .QN(n269) );
  DFFRX1 \i_MIPS/Register/register_reg[28][24]  ( .D(\i_MIPS/Register/n236 ), 
        .CK(clk), .RN(n6298), .Q(\i_MIPS/Register/register[28][24] ), .QN(n303) );
  DFFRX1 \i_MIPS/Register/register_reg[28][25]  ( .D(\i_MIPS/Register/n237 ), 
        .CK(clk), .RN(n6298), .Q(\i_MIPS/Register/register[28][25] ), .QN(n301) );
  DFFRX1 \i_MIPS/Register/register_reg[28][28]  ( .D(\i_MIPS/Register/n240 ), 
        .CK(clk), .RN(n6298), .Q(\i_MIPS/Register/register[28][28] ), .QN(n899) );
  DFFRX1 \i_MIPS/Register/register_reg[28][29]  ( .D(\i_MIPS/Register/n241 ), 
        .CK(clk), .RN(n6298), .Q(\i_MIPS/Register/register[28][29] ), .QN(n286) );
  DFFRX1 \i_MIPS/Register/register_reg[24][15]  ( .D(\i_MIPS/Register/n355 ), 
        .CK(clk), .RN(n6289), .Q(\i_MIPS/Register/register[24][15] ), .QN(n187) );
  DFFRX1 \i_MIPS/Register/register_reg[24][24]  ( .D(\i_MIPS/Register/n364 ), 
        .CK(clk), .RN(n6288), .Q(\i_MIPS/Register/register[24][24] ), .QN(n215) );
  DFFRX1 \i_MIPS/Register/register_reg[24][25]  ( .D(\i_MIPS/Register/n365 ), 
        .CK(clk), .RN(n6288), .Q(\i_MIPS/Register/register[24][25] ), .QN(n182) );
  DFFRX1 \i_MIPS/Register/register_reg[12][2]  ( .D(\i_MIPS/Register/n726 ), 
        .CK(clk), .RN(n6258), .Q(\i_MIPS/Register/register[12][2] ), .QN(n292)
         );
  DFFRX1 \i_MIPS/Register/register_reg[12][15]  ( .D(\i_MIPS/Register/n739 ), 
        .CK(clk), .RN(n6257), .Q(\i_MIPS/Register/register[12][15] ), .QN(n268) );
  DFFRX1 \i_MIPS/Register/register_reg[12][24]  ( .D(\i_MIPS/Register/n748 ), 
        .CK(clk), .RN(n6256), .Q(\i_MIPS/Register/register[12][24] ), .QN(n220) );
  DFFRX1 \i_MIPS/Register/register_reg[12][25]  ( .D(\i_MIPS/Register/n749 ), 
        .CK(clk), .RN(n6256), .Q(\i_MIPS/Register/register[12][25] ), .QN(n302) );
  DFFRX1 \i_MIPS/Register/register_reg[12][28]  ( .D(\i_MIPS/Register/n752 ), 
        .CK(clk), .RN(n6255), .Q(\i_MIPS/Register/register[12][28] ), .QN(n902) );
  DFFRX1 \i_MIPS/Register/register_reg[12][29]  ( .D(\i_MIPS/Register/n753 ), 
        .CK(clk), .RN(n6255), .Q(\i_MIPS/Register/register[12][29] ), .QN(n291) );
  DFFRX1 \i_MIPS/Register/register_reg[8][15]  ( .D(\i_MIPS/Register/n867 ), 
        .CK(clk), .RN(n6246), .Q(\i_MIPS/Register/register[8][15] ), .QN(n186)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][24]  ( .D(\i_MIPS/Register/n876 ), 
        .CK(clk), .RN(n6245), .Q(\i_MIPS/Register/register[8][24] ), .QN(n219)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][25]  ( .D(\i_MIPS/Register/n877 ), 
        .CK(clk), .RN(n6245), .Q(\i_MIPS/Register/register[8][25] ), .QN(n214)
         );
  DFFRX1 \i_MIPS/Register/register_reg[20][15]  ( .D(\i_MIPS/Register/n483 ), 
        .CK(clk), .RN(n6278), .Q(\i_MIPS/Register/register[20][15] ), .QN(n914) );
  DFFRX1 \i_MIPS/Register/register_reg[4][15]  ( .D(\i_MIPS/Register/n995 ), 
        .CK(clk), .RN(n6235), .Q(\i_MIPS/Register/register[4][15] ), .QN(n913)
         );
  DFFRX1 \i_MIPS/IF_ID_reg[27]  ( .D(\i_MIPS/N44 ), .CK(clk), .RN(n6332), .Q(
        \i_MIPS/IF_ID[27] ), .QN(\i_MIPS/n180 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[26]  ( .D(\i_MIPS/N43 ), .CK(clk), .RN(n6332), .Q(
        \i_MIPS/IF_ID[26] ), .QN(\i_MIPS/n179 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[24]  ( .D(\i_MIPS/N41 ), .CK(clk), .RN(n6332), .Q(
        \i_MIPS/IF_ID[24] ), .QN(\i_MIPS/n177 ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][2]  ( .D(\i_MIPS/Register/n534 ), 
        .CK(clk), .RN(n6274), .Q(\i_MIPS/Register/register[18][2] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][6]  ( .D(\i_MIPS/Register/n538 ), 
        .CK(clk), .RN(n6273), .Q(\i_MIPS/Register/register[18][6] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][7]  ( .D(\i_MIPS/Register/n539 ), 
        .CK(clk), .RN(n6273), .Q(\i_MIPS/Register/register[18][7] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][9]  ( .D(\i_MIPS/Register/n541 ), 
        .CK(clk), .RN(n6273), .Q(\i_MIPS/Register/register[18][9] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][13]  ( .D(\i_MIPS/Register/n545 ), 
        .CK(clk), .RN(n6273), .Q(\i_MIPS/Register/register[18][13] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][14]  ( .D(\i_MIPS/Register/n546 ), 
        .CK(clk), .RN(n6273), .Q(\i_MIPS/Register/register[18][14] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][15]  ( .D(\i_MIPS/Register/n547 ), 
        .CK(clk), .RN(n6273), .Q(\i_MIPS/Register/register[18][15] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][22]  ( .D(\i_MIPS/Register/n554 ), 
        .CK(clk), .RN(n6272), .Q(\i_MIPS/Register/register[18][22] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][23]  ( .D(\i_MIPS/Register/n555 ), 
        .CK(clk), .RN(n6272), .Q(\i_MIPS/Register/register[18][23] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][24]  ( .D(\i_MIPS/Register/n556 ), 
        .CK(clk), .RN(n6272), .Q(\i_MIPS/Register/register[18][24] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][25]  ( .D(\i_MIPS/Register/n557 ), 
        .CK(clk), .RN(n6272), .Q(\i_MIPS/Register/register[18][25] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][26]  ( .D(\i_MIPS/Register/n558 ), 
        .CK(clk), .RN(n6272), .Q(\i_MIPS/Register/register[18][26] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][28]  ( .D(\i_MIPS/Register/n560 ), 
        .CK(clk), .RN(n6271), .Q(\i_MIPS/Register/register[18][28] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][29]  ( .D(\i_MIPS/Register/n561 ), 
        .CK(clk), .RN(n6271), .Q(\i_MIPS/Register/register[18][29] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][30]  ( .D(\i_MIPS/Register/n562 ), 
        .CK(clk), .RN(n6271), .Q(\i_MIPS/Register/register[18][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][31]  ( .D(\i_MIPS/Register/n563 ), 
        .CK(clk), .RN(n6271), .Q(\i_MIPS/Register/register[18][31] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][2]  ( .D(\i_MIPS/Register/n1046 ), 
        .CK(clk), .RN(n6231), .Q(\i_MIPS/Register/register[2][2] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][6]  ( .D(\i_MIPS/Register/n1050 ), 
        .CK(clk), .RN(n6231), .Q(\i_MIPS/Register/register[2][6] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][7]  ( .D(\i_MIPS/Register/n1051 ), 
        .CK(clk), .RN(n6231), .Q(\i_MIPS/Register/register[2][7] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][9]  ( .D(\i_MIPS/Register/n1053 ), 
        .CK(clk), .RN(n6230), .Q(\i_MIPS/Register/register[2][9] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][10]  ( .D(\i_MIPS/Register/n1054 ), 
        .CK(clk), .RN(n6230), .Q(\i_MIPS/Register/register[2][10] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][13]  ( .D(\i_MIPS/Register/n1057 ), 
        .CK(clk), .RN(n6230), .Q(\i_MIPS/Register/register[2][13] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][14]  ( .D(\i_MIPS/Register/n1058 ), 
        .CK(clk), .RN(n6230), .Q(\i_MIPS/Register/register[2][14] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][15]  ( .D(\i_MIPS/Register/n1059 ), 
        .CK(clk), .RN(n6230), .Q(\i_MIPS/Register/register[2][15] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][22]  ( .D(\i_MIPS/Register/n1066 ), 
        .CK(clk), .RN(n6229), .Q(\i_MIPS/Register/register[2][22] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][23]  ( .D(\i_MIPS/Register/n1067 ), 
        .CK(clk), .RN(n6229), .Q(\i_MIPS/Register/register[2][23] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][24]  ( .D(\i_MIPS/Register/n1068 ), 
        .CK(clk), .RN(n6229), .Q(\i_MIPS/Register/register[2][24] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][25]  ( .D(\i_MIPS/Register/n1069 ), 
        .CK(clk), .RN(n6229), .Q(\i_MIPS/Register/register[2][25] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][26]  ( .D(\i_MIPS/Register/n1070 ), 
        .CK(clk), .RN(n6229), .Q(\i_MIPS/Register/register[2][26] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][28]  ( .D(\i_MIPS/Register/n1072 ), 
        .CK(clk), .RN(n6229), .Q(\i_MIPS/Register/register[2][28] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][29]  ( .D(\i_MIPS/Register/n1073 ), 
        .CK(clk), .RN(n6229), .Q(\i_MIPS/Register/register[2][29] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][30]  ( .D(\i_MIPS/Register/n1074 ), 
        .CK(clk), .RN(n6229), .Q(\i_MIPS/Register/register[2][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][31]  ( .D(\i_MIPS/Register/n1075 ), 
        .CK(clk), .RN(n6229), .Q(\i_MIPS/Register/register[2][31] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][2]  ( .D(\i_MIPS/Register/n278 ), 
        .CK(clk), .RN(n6295), .Q(\i_MIPS/Register/register[26][2] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][6]  ( .D(\i_MIPS/Register/n282 ), 
        .CK(clk), .RN(n6295), .Q(\i_MIPS/Register/register[26][6] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][9]  ( .D(\i_MIPS/Register/n285 ), 
        .CK(clk), .RN(n6294), .Q(\i_MIPS/Register/register[26][9] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][13]  ( .D(\i_MIPS/Register/n289 ), 
        .CK(clk), .RN(n6294), .Q(\i_MIPS/Register/register[26][13] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][14]  ( .D(\i_MIPS/Register/n290 ), 
        .CK(clk), .RN(n6294), .Q(\i_MIPS/Register/register[26][14] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][15]  ( .D(\i_MIPS/Register/n291 ), 
        .CK(clk), .RN(n6294), .Q(\i_MIPS/Register/register[26][15] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][22]  ( .D(\i_MIPS/Register/n298 ), 
        .CK(clk), .RN(n6293), .Q(\i_MIPS/Register/register[26][22] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][23]  ( .D(\i_MIPS/Register/n299 ), 
        .CK(clk), .RN(n6293), .Q(\i_MIPS/Register/register[26][23] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][24]  ( .D(\i_MIPS/Register/n300 ), 
        .CK(clk), .RN(n6293), .Q(\i_MIPS/Register/register[26][24] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][25]  ( .D(\i_MIPS/Register/n301 ), 
        .CK(clk), .RN(n6293), .Q(\i_MIPS/Register/register[26][25] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][28]  ( .D(\i_MIPS/Register/n304 ), 
        .CK(clk), .RN(n6293), .Q(\i_MIPS/Register/register[26][28] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][29]  ( .D(\i_MIPS/Register/n305 ), 
        .CK(clk), .RN(n6293), .Q(\i_MIPS/Register/register[26][29] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][30]  ( .D(\i_MIPS/Register/n306 ), 
        .CK(clk), .RN(n6293), .Q(\i_MIPS/Register/register[26][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][31]  ( .D(\i_MIPS/Register/n307 ), 
        .CK(clk), .RN(n6293), .Q(\i_MIPS/Register/register[26][31] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][2]  ( .D(\i_MIPS/Register/n790 ), 
        .CK(clk), .RN(n6252), .Q(\i_MIPS/Register/register[10][2] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][6]  ( .D(\i_MIPS/Register/n794 ), 
        .CK(clk), .RN(n6252), .Q(\i_MIPS/Register/register[10][6] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][7]  ( .D(\i_MIPS/Register/n795 ), 
        .CK(clk), .RN(n6252), .Q(\i_MIPS/Register/register[10][7] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][9]  ( .D(\i_MIPS/Register/n797 ), 
        .CK(clk), .RN(n6252), .Q(\i_MIPS/Register/register[10][9] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][13]  ( .D(\i_MIPS/Register/n801 ), 
        .CK(clk), .RN(n6251), .Q(\i_MIPS/Register/register[10][13] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][14]  ( .D(\i_MIPS/Register/n802 ), 
        .CK(clk), .RN(n6251), .Q(\i_MIPS/Register/register[10][14] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][15]  ( .D(\i_MIPS/Register/n803 ), 
        .CK(clk), .RN(n6251), .Q(\i_MIPS/Register/register[10][15] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][22]  ( .D(\i_MIPS/Register/n810 ), 
        .CK(clk), .RN(n6251), .Q(\i_MIPS/Register/register[10][22] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][23]  ( .D(\i_MIPS/Register/n811 ), 
        .CK(clk), .RN(n6251), .Q(\i_MIPS/Register/register[10][23] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][24]  ( .D(\i_MIPS/Register/n812 ), 
        .CK(clk), .RN(n6250), .Q(\i_MIPS/Register/register[10][24] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][25]  ( .D(\i_MIPS/Register/n813 ), 
        .CK(clk), .RN(n6250), .Q(\i_MIPS/Register/register[10][25] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][28]  ( .D(\i_MIPS/Register/n816 ), 
        .CK(clk), .RN(n6250), .Q(\i_MIPS/Register/register[10][28] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][29]  ( .D(\i_MIPS/Register/n817 ), 
        .CK(clk), .RN(n6250), .Q(\i_MIPS/Register/register[10][29] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][30]  ( .D(\i_MIPS/Register/n818 ), 
        .CK(clk), .RN(n6250), .Q(\i_MIPS/Register/register[10][30] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][31]  ( .D(\i_MIPS/Register/n819 ), 
        .CK(clk), .RN(n6250), .Q(\i_MIPS/Register/register[10][31] ) );
  DFFRX1 \i_MIPS/IF_ID_reg[25]  ( .D(\i_MIPS/N42 ), .CK(clk), .RN(n6332), .Q(
        \i_MIPS/IF_ID[25] ), .QN(\i_MIPS/n178 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[23]  ( .D(\i_MIPS/N40 ), .CK(clk), .RN(n6332), .Q(
        \i_MIPS/IF_ID[23] ), .QN(\i_MIPS/n176 ) );
  DFFRX1 \i_MIPS/Register/register_reg[31][14]  ( .D(n11558), .CK(clk), .RN(
        n6307), .QN(n167) );
  DFFRX1 \i_MIPS/Register/register_reg[31][31]  ( .D(n11541), .CK(clk), .RN(
        n6306), .QN(n222) );
  DFFRX1 \i_MIPS/ID_EX_reg[70]  ( .D(\i_MIPS/n309 ), .CK(clk), .RN(n6329), .Q(
        \i_MIPS/ID_EX[70] ), .QN(\i_MIPS/n186 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[67]  ( .D(\i_MIPS/n315 ), .CK(clk), .RN(n6329), .Q(
        \i_MIPS/ID_EX[67] ), .QN(\i_MIPS/n192 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[72]  ( .D(\i_MIPS/n305 ), .CK(clk), .RN(n6330), .Q(
        n3547), .QN(\i_MIPS/n182 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[66]  ( .D(\i_MIPS/n317 ), .CK(clk), .RN(n6329), .Q(
        \i_MIPS/ID_EX[66] ), .QN(\i_MIPS/n194 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[71]  ( .D(\i_MIPS/n307 ), .CK(clk), .RN(n6329), .Q(
        \i_MIPS/ID_EX[71] ), .QN(\i_MIPS/n184 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[3]  ( .D(\i_MIPS/n455 ), .CK(clk), .RN(n6314), .Q(
        \i_MIPS/ID_EX_3 ), .QN(\i_MIPS/n265 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[0]  ( .D(\i_MIPS/n458 ), .CK(clk), .RN(n6314), .Q(
        \i_MIPS/ID_EX_0 ), .QN(\i_MIPS/n302 ) );
  DFFRX1 \I_cache/cache_reg[0][154]  ( .D(n11613), .CK(clk), .RN(n6017), .Q(
        \I_cache/cache[0][154] ), .QN(n2883) );
  DFFRX1 \I_cache/cache_reg[1][154]  ( .D(n11612), .CK(clk), .RN(n6017), .Q(
        \I_cache/cache[1][154] ), .QN(n1265) );
  DFFRX1 \I_cache/cache_reg[2][154]  ( .D(n11611), .CK(clk), .RN(n6017), .Q(
        \I_cache/cache[2][154] ), .QN(n2884) );
  DFFRX1 \I_cache/cache_reg[3][154]  ( .D(n11610), .CK(clk), .RN(n6017), .Q(
        \I_cache/cache[3][154] ), .QN(n1266) );
  DFFRX1 \I_cache/cache_reg[4][154]  ( .D(n11609), .CK(clk), .RN(n6017), .Q(
        \I_cache/cache[4][154] ), .QN(n2885) );
  DFFRX1 \I_cache/cache_reg[5][154]  ( .D(n11608), .CK(clk), .RN(n6017), .Q(
        \I_cache/cache[5][154] ), .QN(n1267) );
  DFFRX1 \I_cache/cache_reg[6][154]  ( .D(n11607), .CK(clk), .RN(n6017), .Q(
        \I_cache/cache[6][154] ), .QN(n2939) );
  DFFRX1 \I_cache/cache_reg[7][154]  ( .D(n11606), .CK(clk), .RN(n6017), .Q(
        \I_cache/cache[7][154] ), .QN(n1305) );
  DFFRX1 \i_MIPS/Register/register_reg[29][14]  ( .D(\i_MIPS/Register/n194 ), 
        .CK(clk), .RN(n6302), .Q(\i_MIPS/Register/register[29][14] ), .QN(n163) );
  DFFRX1 \i_MIPS/Register/register_reg[29][30]  ( .D(\i_MIPS/Register/n210 ), 
        .CK(clk), .RN(n6301), .Q(\i_MIPS/Register/register[29][30] ), .QN(n367) );
  DFFRX1 \i_MIPS/Register/register_reg[29][31]  ( .D(\i_MIPS/Register/n211 ), 
        .CK(clk), .RN(n6301), .Q(\i_MIPS/Register/register[29][31] ), .QN(n162) );
  DFFRX1 \i_MIPS/Register/register_reg[27][14]  ( .D(\i_MIPS/Register/n258 ), 
        .CK(clk), .RN(n6297), .Q(\i_MIPS/Register/register[27][14] ), .QN(n161) );
  DFFRX1 \i_MIPS/Register/register_reg[27][31]  ( .D(\i_MIPS/Register/n275 ), 
        .CK(clk), .RN(n6295), .Q(\i_MIPS/Register/register[27][31] ), .QN(n241) );
  DFFRX1 \i_MIPS/Register/register_reg[25][14]  ( .D(\i_MIPS/Register/n322 ), 
        .CK(clk), .RN(n6291), .Q(\i_MIPS/Register/register[25][14] ), .QN(n363) );
  DFFRX1 \i_MIPS/Register/register_reg[25][30]  ( .D(\i_MIPS/Register/n338 ), 
        .CK(clk), .RN(n6290), .Q(\i_MIPS/Register/register[25][30] ), .QN(n239) );
  DFFRX1 \i_MIPS/Register/register_reg[25][31]  ( .D(\i_MIPS/Register/n339 ), 
        .CK(clk), .RN(n6290), .Q(\i_MIPS/Register/register[25][31] ), .QN(n372) );
  DFFRX1 \i_MIPS/Register/register_reg[23][14]  ( .D(\i_MIPS/Register/n386 ), 
        .CK(clk), .RN(n6286), .Q(\i_MIPS/Register/register[23][14] ), .QN(n245) );
  DFFRX1 \i_MIPS/Register/register_reg[23][31]  ( .D(\i_MIPS/Register/n403 ), 
        .CK(clk), .RN(n6285), .Q(\i_MIPS/Register/register[23][31] ), .QN(n373) );
  DFFRX1 \i_MIPS/Register/register_reg[21][14]  ( .D(\i_MIPS/Register/n450 ), 
        .CK(clk), .RN(n6281), .Q(\i_MIPS/Register/register[21][14] ), .QN(n178) );
  DFFRX1 \i_MIPS/Register/register_reg[21][30]  ( .D(\i_MIPS/Register/n466 ), 
        .CK(clk), .RN(n6279), .Q(\i_MIPS/Register/register[21][30] ), .QN(
        n1989) );
  DFFRX1 \i_MIPS/Register/register_reg[21][31]  ( .D(\i_MIPS/Register/n467 ), 
        .CK(clk), .RN(n6279), .Q(\i_MIPS/Register/register[21][31] ), .QN(n244) );
  DFFRX1 \i_MIPS/Register/register_reg[19][14]  ( .D(\i_MIPS/Register/n514 ), 
        .CK(clk), .RN(n6275), .Q(\i_MIPS/Register/register[19][14] ), .QN(n179) );
  DFFRX1 \i_MIPS/Register/register_reg[19][30]  ( .D(\i_MIPS/Register/n530 ), 
        .CK(clk), .RN(n6274), .Q(\i_MIPS/Register/register[19][30] ), .QN(
        n2002) );
  DFFRX1 \i_MIPS/Register/register_reg[19][31]  ( .D(\i_MIPS/Register/n531 ), 
        .CK(clk), .RN(n6274), .Q(\i_MIPS/Register/register[19][31] ), .QN(n374) );
  DFFRX1 \i_MIPS/Register/register_reg[17][14]  ( .D(\i_MIPS/Register/n578 ), 
        .CK(clk), .RN(n6270), .Q(\i_MIPS/Register/register[17][14] ), .QN(
        n2001) );
  DFFRX1 \i_MIPS/Register/register_reg[17][30]  ( .D(\i_MIPS/Register/n594 ), 
        .CK(clk), .RN(n6269), .Q(\i_MIPS/Register/register[17][30] ), .QN(
        n2007) );
  DFFRX1 \i_MIPS/Register/register_reg[17][31]  ( .D(\i_MIPS/Register/n595 ), 
        .CK(clk), .RN(n6269), .Q(\i_MIPS/Register/register[17][31] ), .QN(
        n1998) );
  DFFRX1 \i_MIPS/Register/register_reg[15][14]  ( .D(\i_MIPS/Register/n642 ), 
        .CK(clk), .RN(n6265), .Q(\i_MIPS/Register/register[15][14] ), .QN(n177) );
  DFFRX1 \i_MIPS/Register/register_reg[13][14]  ( .D(\i_MIPS/Register/n706 ), 
        .CK(clk), .RN(n6259), .Q(\i_MIPS/Register/register[13][14] ), .QN(n242) );
  DFFRX1 \i_MIPS/Register/register_reg[13][30]  ( .D(\i_MIPS/Register/n722 ), 
        .CK(clk), .RN(n6258), .Q(\i_MIPS/Register/register[13][30] ), .QN(n368) );
  DFFRX1 \i_MIPS/Register/register_reg[13][31]  ( .D(\i_MIPS/Register/n723 ), 
        .CK(clk), .RN(n6258), .Q(\i_MIPS/Register/register[13][31] ), .QN(n240) );
  DFFRX1 \i_MIPS/Register/register_reg[11][14]  ( .D(\i_MIPS/Register/n770 ), 
        .CK(clk), .RN(n6254), .Q(\i_MIPS/Register/register[11][14] ), .QN(n175) );
  DFFRX1 \i_MIPS/Register/register_reg[11][31]  ( .D(\i_MIPS/Register/n787 ), 
        .CK(clk), .RN(n6253), .Q(\i_MIPS/Register/register[11][31] ), .QN(n366) );
  DFFRX1 \i_MIPS/Register/register_reg[9][14]  ( .D(\i_MIPS/Register/n834 ), 
        .CK(clk), .RN(n6249), .Q(\i_MIPS/Register/register[9][14] ), .QN(n360)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][30]  ( .D(\i_MIPS/Register/n850 ), 
        .CK(clk), .RN(n6247), .Q(\i_MIPS/Register/register[9][30] ), .QN(n174)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][31]  ( .D(\i_MIPS/Register/n851 ), 
        .CK(clk), .RN(n6247), .Q(\i_MIPS/Register/register[9][31] ), .QN(n176)
         );
  DFFRX1 \i_MIPS/Register/register_reg[7][14]  ( .D(\i_MIPS/Register/n898 ), 
        .CK(clk), .RN(n6243), .Q(\i_MIPS/Register/register[7][14] ), .QN(n246)
         );
  DFFRX1 \i_MIPS/Register/register_reg[7][31]  ( .D(\i_MIPS/Register/n915 ), 
        .CK(clk), .RN(n6242), .Q(\i_MIPS/Register/register[7][31] ), .QN(n1993) );
  DFFRX1 \i_MIPS/Register/register_reg[5][14]  ( .D(\i_MIPS/Register/n962 ), 
        .CK(clk), .RN(n6238), .Q(\i_MIPS/Register/register[5][14] ), .QN(n1994) );
  DFFRX1 \i_MIPS/Register/register_reg[5][30]  ( .D(\i_MIPS/Register/n978 ), 
        .CK(clk), .RN(n6237), .Q(\i_MIPS/Register/register[5][30] ), .QN(n1990) );
  DFFRX1 \i_MIPS/Register/register_reg[5][31]  ( .D(\i_MIPS/Register/n979 ), 
        .CK(clk), .RN(n6237), .Q(\i_MIPS/Register/register[5][31] ), .QN(n1991) );
  DFFRX1 \i_MIPS/Register/register_reg[3][14]  ( .D(\i_MIPS/Register/n1026 ), 
        .CK(clk), .RN(n6233), .Q(\i_MIPS/Register/register[3][14] ), .QN(n247)
         );
  DFFRX1 \i_MIPS/Register/register_reg[3][30]  ( .D(\i_MIPS/Register/n1042 ), 
        .CK(clk), .RN(n6231), .Q(\i_MIPS/Register/register[3][30] ), .QN(n2003) );
  DFFRX1 \i_MIPS/Register/register_reg[3][31]  ( .D(\i_MIPS/Register/n1043 ), 
        .CK(clk), .RN(n6231), .Q(\i_MIPS/Register/register[3][31] ), .QN(n2004) );
  DFFRX1 \i_MIPS/Register/register_reg[1][14]  ( .D(\i_MIPS/Register/n1090 ), 
        .CK(clk), .RN(n6227), .Q(\i_MIPS/Register/register[1][14] ), .QN(n2006) );
  DFFRX1 \i_MIPS/Register/register_reg[1][30]  ( .D(\i_MIPS/Register/n1106 ), 
        .CK(clk), .RN(n6226), .Q(\i_MIPS/Register/register[1][30] ), .QN(n375)
         );
  DFFRX1 \i_MIPS/Register/register_reg[1][31]  ( .D(\i_MIPS/Register/n1107 ), 
        .CK(clk), .RN(n6226), .Q(\i_MIPS/Register/register[1][31] ), .QN(n2005) );
  DFFRX1 \i_MIPS/Register/register_reg[31][0]  ( .D(n11572), .CK(clk), .RN(
        n6308), .Q(\i_MIPS/Register/register[31][0] ), .QN(n227) );
  DFFRX1 \i_MIPS/Register/register_reg[31][1]  ( .D(n11571), .CK(clk), .RN(
        n6308), .Q(\i_MIPS/Register/register[31][1] ), .QN(n170) );
  DFFRX1 \i_MIPS/Register/register_reg[31][2]  ( .D(n11570), .CK(clk), .RN(
        n6308), .Q(\i_MIPS/Register/register[31][2] ), .QN(n237) );
  DFFRX1 \i_MIPS/Register/register_reg[31][3]  ( .D(n11569), .CK(clk), .RN(
        n6308), .Q(\i_MIPS/Register/register[31][3] ), .QN(n228) );
  DFFRX1 \i_MIPS/Register/register_reg[31][4]  ( .D(n11568), .CK(clk), .RN(
        n6308), .Q(\i_MIPS/Register/register[31][4] ), .QN(n359) );
  DFFRX1 \i_MIPS/Register/register_reg[31][5]  ( .D(n11567), .CK(clk), .RN(
        n6308), .Q(\i_MIPS/Register/register[31][5] ), .QN(n226) );
  DFFRX1 \i_MIPS/Register/register_reg[31][6]  ( .D(n11566), .CK(clk), .RN(
        n6308), .Q(\i_MIPS/Register/register[31][6] ), .QN(n232) );
  DFFRX1 \i_MIPS/Register/register_reg[31][7]  ( .D(n11565), .CK(clk), .RN(
        n6308), .Q(\i_MIPS/Register/register[31][7] ), .QN(n231) );
  DFFRX1 \i_MIPS/Register/register_reg[31][8]  ( .D(n11564), .CK(clk), .RN(
        n6308), .Q(\i_MIPS/Register/register[31][8] ), .QN(n173) );
  DFFRX1 \i_MIPS/Register/register_reg[31][9]  ( .D(n11563), .CK(clk), .RN(
        n6308), .Q(\i_MIPS/Register/register[31][9] ), .QN(n165) );
  DFFRX1 \i_MIPS/Register/register_reg[31][10]  ( .D(n11562), .CK(clk), .RN(
        n6308), .Q(\i_MIPS/Register/register[31][10] ), .QN(n164) );
  DFFRX1 \i_MIPS/Register/register_reg[31][11]  ( .D(n11561), .CK(clk), .RN(
        n6308), .Q(\i_MIPS/Register/register[31][11] ), .QN(n172) );
  DFFRX1 \i_MIPS/Register/register_reg[31][12]  ( .D(n11560), .CK(clk), .RN(
        n6307), .Q(\i_MIPS/Register/register[31][12] ), .QN(n171) );
  DFFRX1 \i_MIPS/Register/register_reg[31][13]  ( .D(n11559), .CK(clk), .RN(
        n6307), .Q(\i_MIPS/Register/register[31][13] ), .QN(n159) );
  DFFRX1 \i_MIPS/Register/register_reg[31][15]  ( .D(n11557), .CK(clk), .RN(
        n6307), .Q(\i_MIPS/Register/register[31][15] ), .QN(n160) );
  DFFRX1 \i_MIPS/Register/register_reg[31][16]  ( .D(n11556), .CK(clk), .RN(
        n6307), .Q(\i_MIPS/Register/register[31][16] ), .QN(n229) );
  DFFRX1 \i_MIPS/Register/register_reg[31][17]  ( .D(n11555), .CK(clk), .RN(
        n6307), .Q(\i_MIPS/Register/register[31][17] ), .QN(n169) );
  DFFRX1 \i_MIPS/Register/register_reg[31][18]  ( .D(n11554), .CK(clk), .RN(
        n6307), .Q(\i_MIPS/Register/register[31][18] ), .QN(n225) );
  DFFRX1 \i_MIPS/Register/register_reg[31][19]  ( .D(n11553), .CK(clk), .RN(
        n6307), .Q(\i_MIPS/Register/register[31][19] ), .QN(n158) );
  DFFRX1 \i_MIPS/Register/register_reg[31][20]  ( .D(n11552), .CK(clk), .RN(
        n6307), .Q(\i_MIPS/Register/register[31][20] ), .QN(n356) );
  DFFRX1 \i_MIPS/Register/register_reg[31][21]  ( .D(n11551), .CK(clk), .RN(
        n6307), .Q(\i_MIPS/Register/register[31][21] ), .QN(n230) );
  DFFRX1 \i_MIPS/Register/register_reg[31][23]  ( .D(n11549), .CK(clk), .RN(
        n6307), .Q(\i_MIPS/Register/register[31][23] ), .QN(n236) );
  DFFRX1 \i_MIPS/Register/register_reg[31][24]  ( .D(n11548), .CK(clk), .RN(
        n6306), .Q(\i_MIPS/Register/register[31][24] ), .QN(n224) );
  DFFRX1 \i_MIPS/Register/register_reg[31][25]  ( .D(n11547), .CK(clk), .RN(
        n6306), .Q(\i_MIPS/Register/register[31][25] ), .QN(n238) );
  DFFRX1 \i_MIPS/Register/register_reg[31][26]  ( .D(n11546), .CK(clk), .RN(
        n6306), .Q(\i_MIPS/Register/register[31][26] ), .QN(n235) );
  DFFRX1 \i_MIPS/Register/register_reg[31][27]  ( .D(n11545), .CK(clk), .RN(
        n6306), .Q(\i_MIPS/Register/register[31][27] ), .QN(n259) );
  DFFRX1 \i_MIPS/Register/register_reg[31][28]  ( .D(n11544), .CK(clk), .RN(
        n6306), .Q(\i_MIPS/Register/register[31][28] ), .QN(n234) );
  DFFRX1 \i_MIPS/Register/register_reg[31][29]  ( .D(n11543), .CK(clk), .RN(
        n6306), .Q(\i_MIPS/Register/register[31][29] ), .QN(n233) );
  DFFRX1 \D_cache/cache_reg[0][0]  ( .D(\D_cache/n1795 ), .CK(clk), .RN(n6223), 
        .Q(\D_cache/cache[0][0] ), .QN(n1116) );
  DFFRX1 \D_cache/cache_reg[1][0]  ( .D(\D_cache/n1794 ), .CK(clk), .RN(n6223), 
        .Q(\D_cache/cache[1][0] ), .QN(n2739) );
  DFFRX1 \D_cache/cache_reg[2][0]  ( .D(\D_cache/n1793 ), .CK(clk), .RN(n6223), 
        .Q(\D_cache/cache[2][0] ), .QN(n1115) );
  DFFRX1 \D_cache/cache_reg[3][0]  ( .D(\D_cache/n1792 ), .CK(clk), .RN(n6223), 
        .Q(\D_cache/cache[3][0] ), .QN(n2738) );
  DFFRX1 \D_cache/cache_reg[4][0]  ( .D(\D_cache/n1791 ), .CK(clk), .RN(n6223), 
        .Q(\D_cache/cache[4][0] ), .QN(n606) );
  DFFRX1 \D_cache/cache_reg[5][0]  ( .D(\D_cache/n1790 ), .CK(clk), .RN(n6223), 
        .Q(\D_cache/cache[5][0] ), .QN(n2224) );
  DFFRX1 \D_cache/cache_reg[6][0]  ( .D(\D_cache/n1789 ), .CK(clk), .RN(n6223), 
        .Q(\D_cache/cache[6][0] ), .QN(n2124) );
  DFFRX1 \D_cache/cache_reg[7][0]  ( .D(\D_cache/n1796 ), .CK(clk), .RN(n6223), 
        .Q(\D_cache/cache[7][0] ), .QN(n499) );
  DFFRX1 \D_cache/cache_reg[0][1]  ( .D(\D_cache/n1788 ), .CK(clk), .RN(n6222), 
        .Q(\D_cache/cache[0][1] ), .QN(n1110) );
  DFFRX1 \D_cache/cache_reg[1][1]  ( .D(\D_cache/n1787 ), .CK(clk), .RN(n6222), 
        .Q(\D_cache/cache[1][1] ), .QN(n2733) );
  DFFRX1 \D_cache/cache_reg[2][1]  ( .D(\D_cache/n1786 ), .CK(clk), .RN(n6222), 
        .Q(\D_cache/cache[2][1] ), .QN(n2135) );
  DFFRX1 \D_cache/cache_reg[3][1]  ( .D(\D_cache/n1785 ), .CK(clk), .RN(n6222), 
        .Q(\D_cache/cache[3][1] ), .QN(n510) );
  DFFRX1 \D_cache/cache_reg[4][1]  ( .D(\D_cache/n1784 ), .CK(clk), .RN(n6222), 
        .Q(\D_cache/cache[4][1] ), .QN(n1176) );
  DFFRX1 \D_cache/cache_reg[5][1]  ( .D(\D_cache/n1783 ), .CK(clk), .RN(n6222), 
        .Q(\D_cache/cache[5][1] ), .QN(n2799) );
  DFFRX1 \D_cache/cache_reg[6][1]  ( .D(\D_cache/n1782 ), .CK(clk), .RN(n6222), 
        .Q(\D_cache/cache[6][1] ), .QN(n1109) );
  DFFRX1 \D_cache/cache_reg[7][1]  ( .D(\D_cache/n1781 ), .CK(clk), .RN(n6222), 
        .Q(\D_cache/cache[7][1] ), .QN(n2732) );
  DFFRX1 \D_cache/cache_reg[0][2]  ( .D(\D_cache/n1780 ), .CK(clk), .RN(n6222), 
        .Q(\D_cache/cache[0][2] ), .QN(n949) );
  DFFRX1 \D_cache/cache_reg[1][2]  ( .D(\D_cache/n1779 ), .CK(clk), .RN(n6222), 
        .Q(\D_cache/cache[1][2] ), .QN(n2636) );
  DFFRX1 \D_cache/cache_reg[2][2]  ( .D(\D_cache/n1778 ), .CK(clk), .RN(n6222), 
        .Q(\D_cache/cache[2][2] ), .QN(n1010) );
  DFFRX1 \D_cache/cache_reg[3][2]  ( .D(\D_cache/n1777 ), .CK(clk), .RN(n6222), 
        .Q(\D_cache/cache[3][2] ), .QN(n2635) );
  DFFRX1 \D_cache/cache_reg[4][2]  ( .D(\D_cache/n1776 ), .CK(clk), .RN(n6221), 
        .Q(\D_cache/cache[4][2] ), .QN(n1207) );
  DFFRX1 \D_cache/cache_reg[5][2]  ( .D(\D_cache/n1775 ), .CK(clk), .RN(n6221), 
        .Q(\D_cache/cache[5][2] ), .QN(n2830) );
  DFFRX1 \D_cache/cache_reg[6][2]  ( .D(\D_cache/n1774 ), .CK(clk), .RN(n6221), 
        .Q(\D_cache/cache[6][2] ), .QN(n1009) );
  DFFRX1 \D_cache/cache_reg[7][2]  ( .D(\D_cache/n1773 ), .CK(clk), .RN(n6221), 
        .Q(\D_cache/cache[7][2] ), .QN(n2634) );
  DFFRX1 \D_cache/cache_reg[0][3]  ( .D(\D_cache/n1772 ), .CK(clk), .RN(n6221), 
        .Q(\D_cache/cache[0][3] ), .QN(n663) );
  DFFRX1 \D_cache/cache_reg[1][3]  ( .D(\D_cache/n1771 ), .CK(clk), .RN(n6221), 
        .Q(\D_cache/cache[1][3] ), .QN(n2281) );
  DFFRX1 \D_cache/cache_reg[2][3]  ( .D(\D_cache/n1770 ), .CK(clk), .RN(n6221), 
        .Q(\D_cache/cache[2][3] ), .QN(n992) );
  DFFRX1 \D_cache/cache_reg[3][3]  ( .D(\D_cache/n1769 ), .CK(clk), .RN(n6221), 
        .Q(\D_cache/cache[3][3] ), .QN(n2617) );
  DFFRX1 \D_cache/cache_reg[4][3]  ( .D(\D_cache/n1768 ), .CK(clk), .RN(n6221), 
        .Q(\D_cache/cache[4][3] ), .QN(n2900) );
  DFFRX1 \D_cache/cache_reg[5][3]  ( .D(\D_cache/n1767 ), .CK(clk), .RN(n6221), 
        .Q(\D_cache/cache[5][3] ), .QN(n1079) );
  DFFRX1 \D_cache/cache_reg[6][3]  ( .D(\D_cache/n1766 ), .CK(clk), .RN(n6221), 
        .Q(\D_cache/cache[6][3] ), .QN(n565) );
  DFFRX1 \D_cache/cache_reg[7][3]  ( .D(\D_cache/n1765 ), .CK(clk), .RN(n6221), 
        .Q(\D_cache/cache[7][3] ), .QN(n2280) );
  DFFRX1 \D_cache/cache_reg[0][4]  ( .D(\D_cache/n1764 ), .CK(clk), .RN(n6220), 
        .Q(\D_cache/cache[0][4] ), .QN(n950) );
  DFFRX1 \D_cache/cache_reg[1][4]  ( .D(\D_cache/n1763 ), .CK(clk), .RN(n6220), 
        .Q(\D_cache/cache[1][4] ), .QN(n2668) );
  DFFRX1 \D_cache/cache_reg[2][4]  ( .D(\D_cache/n1762 ), .CK(clk), .RN(n6220), 
        .Q(\D_cache/cache[2][4] ), .QN(n1041) );
  DFFRX1 \D_cache/cache_reg[3][4]  ( .D(\D_cache/n1761 ), .CK(clk), .RN(n6220), 
        .Q(\D_cache/cache[3][4] ), .QN(n2667) );
  DFFRX1 \D_cache/cache_reg[5][4]  ( .D(\D_cache/n1759 ), .CK(clk), .RN(n6220), 
        .Q(\D_cache/cache[5][4] ), .QN(n2031) );
  DFFRX1 \D_cache/cache_reg[6][4]  ( .D(\D_cache/n1758 ), .CK(clk), .RN(n6220), 
        .Q(\D_cache/cache[6][4] ), .QN(n2089) );
  DFFRX1 \D_cache/cache_reg[7][4]  ( .D(\D_cache/n1757 ), .CK(clk), .RN(n6220), 
        .Q(\D_cache/cache[7][4] ), .QN(n463) );
  DFFRX1 \D_cache/cache_reg[0][5]  ( .D(\D_cache/n1756 ), .CK(clk), .RN(n6220), 
        .Q(\D_cache/cache[0][5] ), .QN(n688) );
  DFFRX1 \D_cache/cache_reg[1][5]  ( .D(\D_cache/n1755 ), .CK(clk), .RN(n6220), 
        .Q(\D_cache/cache[1][5] ), .QN(n2306) );
  DFFRX1 \D_cache/cache_reg[2][5]  ( .D(\D_cache/n1754 ), .CK(clk), .RN(n6220), 
        .Q(\D_cache/cache[2][5] ), .QN(n2074) );
  DFFRX1 \D_cache/cache_reg[3][5]  ( .D(\D_cache/n1753 ), .CK(clk), .RN(n6220), 
        .Q(\D_cache/cache[3][5] ), .QN(n449) );
  DFFRX1 \D_cache/cache_reg[4][5]  ( .D(\D_cache/n1752 ), .CK(clk), .RN(n6219), 
        .Q(\D_cache/cache[4][5] ), .QN(n1192) );
  DFFRX1 \D_cache/cache_reg[5][5]  ( .D(\D_cache/n1751 ), .CK(clk), .RN(n6219), 
        .Q(\D_cache/cache[5][5] ), .QN(n2815) );
  DFFRX1 \D_cache/cache_reg[6][5]  ( .D(\D_cache/n1750 ), .CK(clk), .RN(n6219), 
        .Q(\D_cache/cache[6][5] ), .QN(n687) );
  DFFRX1 \D_cache/cache_reg[7][5]  ( .D(\D_cache/n1749 ), .CK(clk), .RN(n6219), 
        .Q(\D_cache/cache[7][5] ), .QN(n2305) );
  DFFRX1 \D_cache/cache_reg[0][6]  ( .D(\D_cache/n1748 ), .CK(clk), .RN(n6219), 
        .Q(\D_cache/cache[0][6] ), .QN(n957) );
  DFFRX1 \D_cache/cache_reg[1][6]  ( .D(\D_cache/n1747 ), .CK(clk), .RN(n6219), 
        .Q(\D_cache/cache[1][6] ), .QN(n2689) );
  DFFRX1 \D_cache/cache_reg[2][6]  ( .D(\D_cache/n1746 ), .CK(clk), .RN(n6219), 
        .Q(\D_cache/cache[2][6] ), .QN(n2096) );
  DFFRX1 \D_cache/cache_reg[3][6]  ( .D(\D_cache/n1745 ), .CK(clk), .RN(n6219), 
        .Q(\D_cache/cache[3][6] ), .QN(n470) );
  DFFRX1 \D_cache/cache_reg[4][6]  ( .D(\D_cache/n1744 ), .CK(clk), .RN(n6219), 
        .Q(\D_cache/cache[4][6] ), .QN(n577) );
  DFFRX1 \D_cache/cache_reg[5][6]  ( .D(\D_cache/n1743 ), .CK(clk), .RN(n6219), 
        .Q(\D_cache/cache[5][6] ), .QN(n2195) );
  DFFRX1 \D_cache/cache_reg[6][6]  ( .D(\D_cache/n1742 ), .CK(clk), .RN(n6219), 
        .Q(\D_cache/cache[6][6] ), .QN(n1061) );
  DFFRX1 \D_cache/cache_reg[7][6]  ( .D(\D_cache/n1741 ), .CK(clk), .RN(n6219), 
        .Q(\D_cache/cache[7][6] ), .QN(n2688) );
  DFFRX1 \D_cache/cache_reg[0][7]  ( .D(\D_cache/n1740 ), .CK(clk), .RN(n6218), 
        .Q(\D_cache/cache[0][7] ), .QN(n620) );
  DFFRX1 \D_cache/cache_reg[1][7]  ( .D(\D_cache/n1739 ), .CK(clk), .RN(n6218), 
        .Q(\D_cache/cache[1][7] ), .QN(n2238) );
  DFFRX1 \D_cache/cache_reg[2][7]  ( .D(\D_cache/n1738 ), .CK(clk), .RN(n6218), 
        .Q(\D_cache/cache[2][7] ), .QN(n1049) );
  DFFRX1 \D_cache/cache_reg[3][7]  ( .D(\D_cache/n1737 ), .CK(clk), .RN(n6218), 
        .Q(\D_cache/cache[3][7] ), .QN(n2676) );
  DFFRX1 \D_cache/cache_reg[4][7]  ( .D(\D_cache/n1736 ), .CK(clk), .RN(n6218), 
        .Q(\D_cache/cache[4][7] ), .QN(n1218) );
  DFFRX1 \D_cache/cache_reg[5][7]  ( .D(\D_cache/n1735 ), .CK(clk), .RN(n6218), 
        .Q(\D_cache/cache[5][7] ), .QN(n2841) );
  DFFRX1 \D_cache/cache_reg[6][7]  ( .D(\D_cache/n1734 ), .CK(clk), .RN(n6218), 
        .Q(\D_cache/cache[6][7] ), .QN(n1048) );
  DFFRX1 \D_cache/cache_reg[7][7]  ( .D(\D_cache/n1733 ), .CK(clk), .RN(n6218), 
        .Q(\D_cache/cache[7][7] ), .QN(n2675) );
  DFFRX1 \D_cache/cache_reg[0][8]  ( .D(\D_cache/n1732 ), .CK(clk), .RN(n6218), 
        .Q(\D_cache/cache[0][8] ), .QN(n1131) );
  DFFRX1 \D_cache/cache_reg[1][8]  ( .D(\D_cache/n1731 ), .CK(clk), .RN(n6218), 
        .Q(\D_cache/cache[1][8] ), .QN(n2754) );
  DFFRX1 \D_cache/cache_reg[2][8]  ( .D(\D_cache/n1730 ), .CK(clk), .RN(n6218), 
        .Q(\D_cache/cache[2][8] ), .QN(n1130) );
  DFFRX1 \D_cache/cache_reg[3][8]  ( .D(\D_cache/n1729 ), .CK(clk), .RN(n6218), 
        .Q(\D_cache/cache[3][8] ), .QN(n2753) );
  DFFRX1 \D_cache/cache_reg[4][8]  ( .D(\D_cache/n1728 ), .CK(clk), .RN(n6217), 
        .Q(\D_cache/cache[4][8] ), .QN(n1237) );
  DFFRX1 \D_cache/cache_reg[5][8]  ( .D(\D_cache/n1727 ), .CK(clk), .RN(n6217), 
        .Q(\D_cache/cache[5][8] ), .QN(n2859) );
  DFFRX1 \D_cache/cache_reg[6][8]  ( .D(\D_cache/n1726 ), .CK(clk), .RN(n6217), 
        .Q(\D_cache/cache[6][8] ), .QN(n1129) );
  DFFRX1 \D_cache/cache_reg[7][8]  ( .D(\D_cache/n1725 ), .CK(clk), .RN(n6217), 
        .Q(\D_cache/cache[7][8] ), .QN(n2752) );
  DFFRX1 \D_cache/cache_reg[0][9]  ( .D(\D_cache/n1724 ), .CK(clk), .RN(n6217), 
        .Q(\D_cache/cache[0][9] ), .QN(n1045) );
  DFFRX1 \D_cache/cache_reg[1][9]  ( .D(\D_cache/n1723 ), .CK(clk), .RN(n6217), 
        .Q(\D_cache/cache[1][9] ), .QN(n2672) );
  DFFRX1 \D_cache/cache_reg[2][9]  ( .D(\D_cache/n1722 ), .CK(clk), .RN(n6217), 
        .Q(\D_cache/cache[2][9] ), .QN(n1044) );
  DFFRX1 \D_cache/cache_reg[3][9]  ( .D(\D_cache/n1721 ), .CK(clk), .RN(n6217), 
        .Q(\D_cache/cache[3][9] ), .QN(n2671) );
  DFFRX1 \D_cache/cache_reg[4][9]  ( .D(\D_cache/n1720 ), .CK(clk), .RN(n6217), 
        .Q(\D_cache/cache[4][9] ), .QN(n1205) );
  DFFRX1 \D_cache/cache_reg[5][9]  ( .D(\D_cache/n1719 ), .CK(clk), .RN(n6217), 
        .Q(\D_cache/cache[5][9] ), .QN(n2828) );
  DFFRX1 \D_cache/cache_reg[6][9]  ( .D(\D_cache/n1718 ), .CK(clk), .RN(n6217), 
        .Q(\D_cache/cache[6][9] ), .QN(n1043) );
  DFFRX1 \D_cache/cache_reg[7][9]  ( .D(\D_cache/n1717 ), .CK(clk), .RN(n6217), 
        .Q(\D_cache/cache[7][9] ), .QN(n2670) );
  DFFRX1 \D_cache/cache_reg[0][10]  ( .D(\D_cache/n1716 ), .CK(clk), .RN(n6216), .Q(\D_cache/cache[0][10] ), .QN(n1040) );
  DFFRX1 \D_cache/cache_reg[1][10]  ( .D(\D_cache/n1715 ), .CK(clk), .RN(n6216), .Q(\D_cache/cache[1][10] ), .QN(n2666) );
  DFFRX1 \D_cache/cache_reg[2][10]  ( .D(\D_cache/n1714 ), .CK(clk), .RN(n6216), .Q(\D_cache/cache[2][10] ), .QN(n1039) );
  DFFRX1 \D_cache/cache_reg[3][10]  ( .D(\D_cache/n1713 ), .CK(clk), .RN(n6216), .Q(\D_cache/cache[3][10] ), .QN(n2665) );
  DFFRX1 \D_cache/cache_reg[4][10]  ( .D(\D_cache/n1712 ), .CK(clk), .RN(n6216), .Q(\D_cache/cache[4][10] ), .QN(n1206) );
  DFFRX1 \D_cache/cache_reg[5][10]  ( .D(\D_cache/n1711 ), .CK(clk), .RN(n6216), .Q(\D_cache/cache[5][10] ), .QN(n2829) );
  DFFRX1 \D_cache/cache_reg[6][10]  ( .D(\D_cache/n1710 ), .CK(clk), .RN(n6216), .Q(\D_cache/cache[6][10] ), .QN(n1038) );
  DFFRX1 \D_cache/cache_reg[7][10]  ( .D(\D_cache/n1709 ), .CK(clk), .RN(n6216), .Q(\D_cache/cache[7][10] ), .QN(n2664) );
  DFFRX1 \D_cache/cache_reg[0][11]  ( .D(\D_cache/n1708 ), .CK(clk), .RN(n6216), .Q(\D_cache/cache[0][11] ), .QN(n1157) );
  DFFRX1 \D_cache/cache_reg[1][11]  ( .D(\D_cache/n1707 ), .CK(clk), .RN(n6216), .Q(\D_cache/cache[1][11] ), .QN(n2780) );
  DFFRX1 \D_cache/cache_reg[2][11]  ( .D(\D_cache/n1706 ), .CK(clk), .RN(n6216), .Q(\D_cache/cache[2][11] ), .QN(n2114) );
  DFFRX1 \D_cache/cache_reg[3][11]  ( .D(\D_cache/n1705 ), .CK(clk), .RN(n6216), .Q(\D_cache/cache[3][11] ), .QN(n488) );
  DFFRX1 \D_cache/cache_reg[4][11]  ( .D(\D_cache/n1704 ), .CK(clk), .RN(n6215), .Q(\D_cache/cache[4][11] ), .QN(n968) );
  DFFRX1 \D_cache/cache_reg[5][11]  ( .D(\D_cache/n1703 ), .CK(clk), .RN(n6215), .Q(\D_cache/cache[5][11] ), .QN(n2593) );
  DFFRX1 \D_cache/cache_reg[6][11]  ( .D(\D_cache/n1702 ), .CK(clk), .RN(n6215), .Q(\D_cache/cache[6][11] ), .QN(n1156) );
  DFFRX1 \D_cache/cache_reg[7][11]  ( .D(\D_cache/n1701 ), .CK(clk), .RN(n6215), .Q(\D_cache/cache[7][11] ), .QN(n2779) );
  DFFRX1 \D_cache/cache_reg[0][12]  ( .D(\D_cache/n1700 ), .CK(clk), .RN(n6215), .Q(\D_cache/cache[0][12] ), .QN(n1128) );
  DFFRX1 \D_cache/cache_reg[1][12]  ( .D(\D_cache/n1699 ), .CK(clk), .RN(n6215), .Q(\D_cache/cache[1][12] ), .QN(n2751) );
  DFFRX1 \D_cache/cache_reg[2][12]  ( .D(\D_cache/n1698 ), .CK(clk), .RN(n6215), .Q(\D_cache/cache[2][12] ), .QN(n1127) );
  DFFRX1 \D_cache/cache_reg[3][12]  ( .D(\D_cache/n1697 ), .CK(clk), .RN(n6215), .Q(\D_cache/cache[3][12] ), .QN(n2750) );
  DFFRX1 \D_cache/cache_reg[4][12]  ( .D(\D_cache/n1696 ), .CK(clk), .RN(n6215), .Q(\D_cache/cache[4][12] ), .QN(n1235) );
  DFFRX1 \D_cache/cache_reg[5][12]  ( .D(\D_cache/n1695 ), .CK(clk), .RN(n6215), .Q(\D_cache/cache[5][12] ), .QN(n2857) );
  DFFRX1 \D_cache/cache_reg[6][12]  ( .D(\D_cache/n1694 ), .CK(clk), .RN(n6215), .Q(\D_cache/cache[6][12] ), .QN(n1126) );
  DFFRX1 \D_cache/cache_reg[7][12]  ( .D(\D_cache/n1693 ), .CK(clk), .RN(n6215), .Q(\D_cache/cache[7][12] ), .QN(n2749) );
  DFFRX1 \D_cache/cache_reg[0][13]  ( .D(\D_cache/n1692 ), .CK(clk), .RN(n6214), .Q(\D_cache/cache[0][13] ), .QN(n669) );
  DFFRX1 \D_cache/cache_reg[1][13]  ( .D(\D_cache/n1691 ), .CK(clk), .RN(n6214), .Q(\D_cache/cache[1][13] ), .QN(n2287) );
  DFFRX1 \D_cache/cache_reg[2][13]  ( .D(\D_cache/n1690 ), .CK(clk), .RN(n6214), .Q(\D_cache/cache[2][13] ), .QN(n994) );
  DFFRX1 \D_cache/cache_reg[3][13]  ( .D(\D_cache/n1689 ), .CK(clk), .RN(n6214), .Q(\D_cache/cache[3][13] ), .QN(n2619) );
  DFFRX1 \D_cache/cache_reg[4][13]  ( .D(\D_cache/n1688 ), .CK(clk), .RN(n6214), .Q(\D_cache/cache[4][13] ), .QN(n583) );
  DFFRX1 \D_cache/cache_reg[5][13]  ( .D(\D_cache/n1687 ), .CK(clk), .RN(n6214), .Q(\D_cache/cache[5][13] ), .QN(n2201) );
  DFFRX1 \D_cache/cache_reg[6][13]  ( .D(\D_cache/n1686 ), .CK(clk), .RN(n6214), .Q(\D_cache/cache[6][13] ), .QN(n668) );
  DFFRX1 \D_cache/cache_reg[7][13]  ( .D(\D_cache/n1685 ), .CK(clk), .RN(n6214), .Q(\D_cache/cache[7][13] ), .QN(n2286) );
  DFFRX1 \D_cache/cache_reg[0][14]  ( .D(\D_cache/n1684 ), .CK(clk), .RN(n6214), .Q(\D_cache/cache[0][14] ), .QN(n1016) );
  DFFRX1 \D_cache/cache_reg[1][14]  ( .D(\D_cache/n1683 ), .CK(clk), .RN(n6214), .Q(\D_cache/cache[1][14] ), .QN(n2642) );
  DFFRX1 \D_cache/cache_reg[2][14]  ( .D(\D_cache/n1682 ), .CK(clk), .RN(n6214), .Q(\D_cache/cache[2][14] ), .QN(n579) );
  DFFRX1 \D_cache/cache_reg[3][14]  ( .D(\D_cache/n1681 ), .CK(clk), .RN(n6214), .Q(\D_cache/cache[3][14] ), .QN(n2197) );
  DFFRX1 \D_cache/cache_reg[4][14]  ( .D(\D_cache/n1680 ), .CK(clk), .RN(n6213), .Q(\D_cache/cache[4][14] ), .QN(n967) );
  DFFRX1 \D_cache/cache_reg[5][14]  ( .D(\D_cache/n1679 ), .CK(clk), .RN(n6213), .Q(\D_cache/cache[5][14] ), .QN(n2592) );
  DFFRX1 \D_cache/cache_reg[6][14]  ( .D(\D_cache/n1678 ), .CK(clk), .RN(n6213), .Q(\D_cache/cache[6][14] ), .QN(n1015) );
  DFFRX1 \D_cache/cache_reg[7][14]  ( .D(\D_cache/n1677 ), .CK(clk), .RN(n6213), .Q(\D_cache/cache[7][14] ), .QN(n2641) );
  DFFRX1 \D_cache/cache_reg[0][15]  ( .D(\D_cache/n1676 ), .CK(clk), .RN(n6213), .Q(\D_cache/cache[0][15] ), .QN(n1008) );
  DFFRX1 \D_cache/cache_reg[1][15]  ( .D(\D_cache/n1675 ), .CK(clk), .RN(n6213), .Q(\D_cache/cache[1][15] ), .QN(n2633) );
  DFFRX1 \D_cache/cache_reg[2][15]  ( .D(\D_cache/n1674 ), .CK(clk), .RN(n6213), .Q(\D_cache/cache[2][15] ), .QN(n1007) );
  DFFRX1 \D_cache/cache_reg[3][15]  ( .D(\D_cache/n1673 ), .CK(clk), .RN(n6213), .Q(\D_cache/cache[3][15] ), .QN(n2632) );
  DFFRX1 \D_cache/cache_reg[4][15]  ( .D(\D_cache/n1672 ), .CK(clk), .RN(n6213), .Q(\D_cache/cache[4][15] ), .QN(n1204) );
  DFFRX1 \D_cache/cache_reg[5][15]  ( .D(\D_cache/n1671 ), .CK(clk), .RN(n6213), .Q(\D_cache/cache[5][15] ), .QN(n2827) );
  DFFRX1 \D_cache/cache_reg[6][15]  ( .D(\D_cache/n1670 ), .CK(clk), .RN(n6213), .Q(\D_cache/cache[6][15] ), .QN(n1006) );
  DFFRX1 \D_cache/cache_reg[7][15]  ( .D(\D_cache/n1669 ), .CK(clk), .RN(n6213), .Q(\D_cache/cache[7][15] ), .QN(n2631) );
  DFFRX1 \D_cache/cache_reg[0][16]  ( .D(\D_cache/n1668 ), .CK(clk), .RN(n6212), .Q(\D_cache/cache[0][16] ), .QN(n1133) );
  DFFRX1 \D_cache/cache_reg[1][16]  ( .D(\D_cache/n1667 ), .CK(clk), .RN(n6212), .Q(\D_cache/cache[1][16] ), .QN(n2756) );
  DFFRX1 \D_cache/cache_reg[2][16]  ( .D(\D_cache/n1666 ), .CK(clk), .RN(n6212), .Q(\D_cache/cache[2][16] ), .QN(n1132) );
  DFFRX1 \D_cache/cache_reg[3][16]  ( .D(\D_cache/n1665 ), .CK(clk), .RN(n6212), .Q(\D_cache/cache[3][16] ), .QN(n2755) );
  DFFRX1 \D_cache/cache_reg[4][16]  ( .D(\D_cache/n1664 ), .CK(clk), .RN(n6212), .Q(\D_cache/cache[4][16] ), .QN(n608) );
  DFFRX1 \D_cache/cache_reg[5][16]  ( .D(\D_cache/n1663 ), .CK(clk), .RN(n6212), .Q(\D_cache/cache[5][16] ), .QN(n2226) );
  DFFRX1 \D_cache/cache_reg[6][16]  ( .D(\D_cache/n1662 ), .CK(clk), .RN(n6212), .Q(\D_cache/cache[6][16] ), .QN(n2127) );
  DFFRX1 \D_cache/cache_reg[7][16]  ( .D(\D_cache/n1661 ), .CK(clk), .RN(n6212), .Q(\D_cache/cache[7][16] ), .QN(n502) );
  DFFRX1 \D_cache/cache_reg[0][17]  ( .D(\D_cache/n1660 ), .CK(clk), .RN(n6212), .Q(\D_cache/cache[0][17] ), .QN(n1160) );
  DFFRX1 \D_cache/cache_reg[1][17]  ( .D(\D_cache/n1659 ), .CK(clk), .RN(n6212), .Q(\D_cache/cache[1][17] ), .QN(n2783) );
  DFFRX1 \D_cache/cache_reg[2][17]  ( .D(\D_cache/n1658 ), .CK(clk), .RN(n6212), .Q(\D_cache/cache[2][17] ), .QN(n1159) );
  DFFRX1 \D_cache/cache_reg[3][17]  ( .D(\D_cache/n1657 ), .CK(clk), .RN(n6212), .Q(\D_cache/cache[3][17] ), .QN(n2782) );
  DFFRX1 \D_cache/cache_reg[4][17]  ( .D(\D_cache/n1656 ), .CK(clk), .RN(n6211), .Q(\D_cache/cache[4][17] ), .QN(n966) );
  DFFRX1 \D_cache/cache_reg[5][17]  ( .D(\D_cache/n1655 ), .CK(clk), .RN(n6211), .Q(\D_cache/cache[5][17] ), .QN(n2591) );
  DFFRX1 \D_cache/cache_reg[6][17]  ( .D(\D_cache/n1654 ), .CK(clk), .RN(n6211), .Q(\D_cache/cache[6][17] ), .QN(n1158) );
  DFFRX1 \D_cache/cache_reg[7][17]  ( .D(\D_cache/n1653 ), .CK(clk), .RN(n6211), .Q(\D_cache/cache[7][17] ), .QN(n2781) );
  DFFRX1 \D_cache/cache_reg[0][18]  ( .D(\D_cache/n1652 ), .CK(clk), .RN(n6211), .Q(\D_cache/cache[0][18] ), .QN(n1122) );
  DFFRX1 \D_cache/cache_reg[1][18]  ( .D(\D_cache/n1651 ), .CK(clk), .RN(n6211), .Q(\D_cache/cache[1][18] ), .QN(n2745) );
  DFFRX1 \D_cache/cache_reg[2][18]  ( .D(\D_cache/n1650 ), .CK(clk), .RN(n6211), .Q(\D_cache/cache[2][18] ), .QN(n1121) );
  DFFRX1 \D_cache/cache_reg[3][18]  ( .D(\D_cache/n1649 ), .CK(clk), .RN(n6211), .Q(\D_cache/cache[3][18] ), .QN(n2744) );
  DFFRX1 \D_cache/cache_reg[5][18]  ( .D(\D_cache/n1647 ), .CK(clk), .RN(n6211), .Q(\D_cache/cache[5][18] ), .QN(n2032) );
  DFFRX1 \D_cache/cache_reg[6][18]  ( .D(\D_cache/n1646 ), .CK(clk), .RN(n6211), .Q(\D_cache/cache[6][18] ), .QN(n1120) );
  DFFRX1 \D_cache/cache_reg[7][18]  ( .D(\D_cache/n1645 ), .CK(clk), .RN(n6211), .Q(\D_cache/cache[7][18] ), .QN(n2743) );
  DFFRX1 \D_cache/cache_reg[0][19]  ( .D(\D_cache/n1644 ), .CK(clk), .RN(n6210), .Q(\D_cache/cache[0][19] ), .QN(n665) );
  DFFRX1 \D_cache/cache_reg[1][19]  ( .D(\D_cache/n1643 ), .CK(clk), .RN(n6210), .Q(\D_cache/cache[1][19] ), .QN(n2283) );
  DFFRX1 \D_cache/cache_reg[2][19]  ( .D(\D_cache/n1642 ), .CK(clk), .RN(n6210), .Q(\D_cache/cache[2][19] ), .QN(n2130) );
  DFFRX1 \D_cache/cache_reg[3][19]  ( .D(\D_cache/n1641 ), .CK(clk), .RN(n6210), .Q(\D_cache/cache[3][19] ), .QN(n505) );
  DFFRX1 \D_cache/cache_reg[4][19]  ( .D(\D_cache/n1640 ), .CK(clk), .RN(n6210), .Q(\D_cache/cache[4][19] ), .QN(n1190) );
  DFFRX1 \D_cache/cache_reg[5][19]  ( .D(\D_cache/n1639 ), .CK(clk), .RN(n6210), .Q(\D_cache/cache[5][19] ), .QN(n2813) );
  DFFRX1 \D_cache/cache_reg[6][19]  ( .D(\D_cache/n1638 ), .CK(clk), .RN(n6210), .Q(\D_cache/cache[6][19] ), .QN(n664) );
  DFFRX1 \D_cache/cache_reg[7][19]  ( .D(\D_cache/n1637 ), .CK(clk), .RN(n6210), .Q(\D_cache/cache[7][19] ), .QN(n2282) );
  DFFRX1 \D_cache/cache_reg[0][21]  ( .D(\D_cache/n1628 ), .CK(clk), .RN(n6209), .Q(\D_cache/cache[0][21] ), .QN(n1145) );
  DFFRX1 \D_cache/cache_reg[1][21]  ( .D(\D_cache/n1627 ), .CK(clk), .RN(n6209), .Q(\D_cache/cache[1][21] ), .QN(n2768) );
  DFFRX1 \D_cache/cache_reg[2][21]  ( .D(\D_cache/n1626 ), .CK(clk), .RN(n6209), .Q(\D_cache/cache[2][21] ), .QN(n1144) );
  DFFRX1 \D_cache/cache_reg[3][21]  ( .D(\D_cache/n1625 ), .CK(clk), .RN(n6209), .Q(\D_cache/cache[3][21] ), .QN(n2767) );
  DFFRX1 \D_cache/cache_reg[5][21]  ( .D(\D_cache/n1623 ), .CK(clk), .RN(n6209), .Q(\D_cache/cache[5][21] ), .QN(n2889) );
  DFFRX1 \D_cache/cache_reg[6][21]  ( .D(\D_cache/n1622 ), .CK(clk), .RN(n6209), .Q(\D_cache/cache[6][21] ), .QN(n1143) );
  DFFRX1 \D_cache/cache_reg[7][21]  ( .D(\D_cache/n1621 ), .CK(clk), .RN(n6209), .Q(\D_cache/cache[7][21] ), .QN(n2766) );
  DFFRX1 \D_cache/cache_reg[0][22]  ( .D(\D_cache/n1620 ), .CK(clk), .RN(n6208), .Q(\D_cache/cache[0][22] ), .QN(n637) );
  DFFRX1 \D_cache/cache_reg[1][22]  ( .D(\D_cache/n1619 ), .CK(clk), .RN(n6208), .Q(\D_cache/cache[1][22] ), .QN(n2254) );
  DFFRX1 \D_cache/cache_reg[2][22]  ( .D(\D_cache/n1618 ), .CK(clk), .RN(n6208), .Q(\D_cache/cache[2][22] ), .QN(n990) );
  DFFRX1 \D_cache/cache_reg[3][22]  ( .D(\D_cache/n1617 ), .CK(clk), .RN(n6208), .Q(\D_cache/cache[3][22] ), .QN(n2615) );
  DFFRX1 \D_cache/cache_reg[4][22]  ( .D(\D_cache/n1616 ), .CK(clk), .RN(n6208), .Q(\D_cache/cache[4][22] ), .QN(n626) );
  DFFRX1 \D_cache/cache_reg[5][22]  ( .D(\D_cache/n1615 ), .CK(clk), .RN(n6208), .Q(\D_cache/cache[5][22] ), .QN(n2244) );
  DFFRX1 \D_cache/cache_reg[6][22]  ( .D(\D_cache/n1614 ), .CK(clk), .RN(n6208), .Q(\D_cache/cache[6][22] ), .QN(n636) );
  DFFRX1 \D_cache/cache_reg[7][22]  ( .D(\D_cache/n1613 ), .CK(clk), .RN(n6208), .Q(\D_cache/cache[7][22] ), .QN(n2253) );
  DFFRX1 \D_cache/cache_reg[0][23]  ( .D(\D_cache/n1612 ), .CK(clk), .RN(n6208), .Q(\D_cache/cache[0][23] ), .QN(n686) );
  DFFRX1 \D_cache/cache_reg[1][23]  ( .D(\D_cache/n1611 ), .CK(clk), .RN(n6208), .Q(\D_cache/cache[1][23] ), .QN(n2304) );
  DFFRX1 \D_cache/cache_reg[2][23]  ( .D(\D_cache/n1610 ), .CK(clk), .RN(n6208), .Q(\D_cache/cache[2][23] ), .QN(n1001) );
  DFFRX1 \D_cache/cache_reg[3][23]  ( .D(\D_cache/n1609 ), .CK(clk), .RN(n6208), .Q(\D_cache/cache[3][23] ), .QN(n2626) );
  DFFRX1 \D_cache/cache_reg[4][23]  ( .D(\D_cache/n1608 ), .CK(clk), .RN(n6207), .Q(\D_cache/cache[4][23] ), .QN(n1194) );
  DFFRX1 \D_cache/cache_reg[5][23]  ( .D(\D_cache/n1607 ), .CK(clk), .RN(n6207), .Q(\D_cache/cache[5][23] ), .QN(n2817) );
  DFFRX1 \D_cache/cache_reg[6][23]  ( .D(\D_cache/n1606 ), .CK(clk), .RN(n6207), .Q(\D_cache/cache[6][23] ), .QN(n685) );
  DFFRX1 \D_cache/cache_reg[7][23]  ( .D(\D_cache/n1605 ), .CK(clk), .RN(n6207), .Q(\D_cache/cache[7][23] ), .QN(n2303) );
  DFFRX1 \D_cache/cache_reg[0][26]  ( .D(\D_cache/n1588 ), .CK(clk), .RN(n6206), .Q(\D_cache/cache[0][26] ), .QN(n658) );
  DFFRX1 \D_cache/cache_reg[1][26]  ( .D(\D_cache/n1587 ), .CK(clk), .RN(n6206), .Q(\D_cache/cache[1][26] ), .QN(n2275) );
  DFFRX1 \D_cache/cache_reg[2][26]  ( .D(\D_cache/n1586 ), .CK(clk), .RN(n6206), .Q(\D_cache/cache[2][26] ), .QN(n1082) );
  DFFRX1 \D_cache/cache_reg[3][26]  ( .D(\D_cache/n1585 ), .CK(clk), .RN(n6206), .Q(\D_cache/cache[3][26] ), .QN(n2705) );
  DFFRX1 \D_cache/cache_reg[4][26]  ( .D(\D_cache/n1584 ), .CK(clk), .RN(n6205), .Q(\D_cache/cache[4][26] ), .QN(n1177) );
  DFFRX1 \D_cache/cache_reg[5][26]  ( .D(\D_cache/n1583 ), .CK(clk), .RN(n6205), .Q(\D_cache/cache[5][26] ), .QN(n2800) );
  DFFRX1 \D_cache/cache_reg[6][26]  ( .D(\D_cache/n1582 ), .CK(clk), .RN(n6205), .Q(\D_cache/cache[6][26] ), .QN(n657) );
  DFFRX1 \D_cache/cache_reg[7][26]  ( .D(\D_cache/n1581 ), .CK(clk), .RN(n6205), .Q(\D_cache/cache[7][26] ), .QN(n2274) );
  DFFRX1 \D_cache/cache_reg[0][27]  ( .D(\D_cache/n1580 ), .CK(clk), .RN(n6205), .Q(\D_cache/cache[0][27] ), .QN(n2893) );
  DFFRX1 \D_cache/cache_reg[1][27]  ( .D(\D_cache/n1579 ), .CK(clk), .RN(n6205), .Q(\D_cache/cache[1][27] ), .QN(n1230) );
  DFFRX1 \D_cache/cache_reg[2][27]  ( .D(\D_cache/n1578 ), .CK(clk), .RN(n6205), .Q(\D_cache/cache[2][27] ), .QN(n1068) );
  DFFRX1 \D_cache/cache_reg[3][27]  ( .D(\D_cache/n1577 ), .CK(clk), .RN(n6205), .Q(\D_cache/cache[3][27] ), .QN(n2696) );
  DFFRX1 \D_cache/cache_reg[4][27]  ( .D(\D_cache/n1576 ), .CK(clk), .RN(n6205), .Q(\D_cache/cache[4][27] ), .QN(n969) );
  DFFRX1 \D_cache/cache_reg[5][27]  ( .D(\D_cache/n1575 ), .CK(clk), .RN(n6205), .Q(\D_cache/cache[5][27] ), .QN(n2594) );
  DFFRX1 \D_cache/cache_reg[6][27]  ( .D(\D_cache/n1574 ), .CK(clk), .RN(n6205), .Q(\D_cache/cache[6][27] ), .QN(n1067) );
  DFFRX1 \D_cache/cache_reg[7][27]  ( .D(\D_cache/n1573 ), .CK(clk), .RN(n6205), .Q(\D_cache/cache[7][27] ), .QN(n2695) );
  DFFRX1 \D_cache/cache_reg[0][28]  ( .D(\D_cache/n1572 ), .CK(clk), .RN(n6204), .Q(\D_cache/cache[0][28] ), .QN(n692) );
  DFFRX1 \D_cache/cache_reg[1][28]  ( .D(\D_cache/n1571 ), .CK(clk), .RN(n6204), .Q(\D_cache/cache[1][28] ), .QN(n2310) );
  DFFRX1 \D_cache/cache_reg[2][28]  ( .D(\D_cache/n1570 ), .CK(clk), .RN(n6204), .Q(\D_cache/cache[2][28] ), .QN(n1002) );
  DFFRX1 \D_cache/cache_reg[3][28]  ( .D(\D_cache/n1569 ), .CK(clk), .RN(n6204), .Q(\D_cache/cache[3][28] ), .QN(n2627) );
  DFFRX1 \D_cache/cache_reg[4][28]  ( .D(\D_cache/n1568 ), .CK(clk), .RN(n6204), .Q(\D_cache/cache[4][28] ), .QN(n587) );
  DFFRX1 \D_cache/cache_reg[5][28]  ( .D(\D_cache/n1567 ), .CK(clk), .RN(n6204), .Q(\D_cache/cache[5][28] ), .QN(n2205) );
  DFFRX1 \D_cache/cache_reg[6][28]  ( .D(\D_cache/n1566 ), .CK(clk), .RN(n6204), .Q(\D_cache/cache[6][28] ), .QN(n691) );
  DFFRX1 \D_cache/cache_reg[7][28]  ( .D(\D_cache/n1565 ), .CK(clk), .RN(n6204), .Q(\D_cache/cache[7][28] ), .QN(n2309) );
  DFFRX1 \D_cache/cache_reg[0][29]  ( .D(\D_cache/n1564 ), .CK(clk), .RN(n6204), .Q(\D_cache/cache[0][29] ), .QN(n1231) );
  DFFRX1 \D_cache/cache_reg[1][29]  ( .D(\D_cache/n1563 ), .CK(clk), .RN(n6204), .Q(\D_cache/cache[1][29] ), .QN(n2853) );
  DFFRX1 \D_cache/cache_reg[2][29]  ( .D(\D_cache/n1562 ), .CK(clk), .RN(n6204), .Q(\D_cache/cache[2][29] ), .QN(n1072) );
  DFFRX1 \D_cache/cache_reg[3][29]  ( .D(\D_cache/n1561 ), .CK(clk), .RN(n6204), .Q(\D_cache/cache[3][29] ), .QN(n2700) );
  DFFRX1 \D_cache/cache_reg[4][29]  ( .D(\D_cache/n1560 ), .CK(clk), .RN(n6203), .Q(\D_cache/cache[4][29] ), .QN(n1281) );
  DFFRX1 \D_cache/cache_reg[5][29]  ( .D(\D_cache/n1559 ), .CK(clk), .RN(n6203), .Q(\D_cache/cache[5][29] ), .QN(n2913) );
  DFFRX1 \D_cache/cache_reg[6][29]  ( .D(\D_cache/n1558 ), .CK(clk), .RN(n6203), .Q(\D_cache/cache[6][29] ), .QN(n596) );
  DFFRX1 \D_cache/cache_reg[7][29]  ( .D(\D_cache/n1557 ), .CK(clk), .RN(n6203), .Q(\D_cache/cache[7][29] ), .QN(n2214) );
  DFFRX1 \D_cache/cache_reg[0][30]  ( .D(\D_cache/n1556 ), .CK(clk), .RN(n6203), .Q(\D_cache/cache[0][30] ), .QN(n661) );
  DFFRX1 \D_cache/cache_reg[1][30]  ( .D(\D_cache/n1555 ), .CK(clk), .RN(n6203), .Q(\D_cache/cache[1][30] ), .QN(n2278) );
  DFFRX1 \D_cache/cache_reg[2][30]  ( .D(\D_cache/n1554 ), .CK(clk), .RN(n6203), .Q(\D_cache/cache[2][30] ), .QN(n660) );
  DFFRX1 \D_cache/cache_reg[3][30]  ( .D(\D_cache/n1553 ), .CK(clk), .RN(n6203), .Q(\D_cache/cache[3][30] ), .QN(n2277) );
  DFFRX1 \D_cache/cache_reg[4][30]  ( .D(\D_cache/n1552 ), .CK(clk), .RN(n6203), .Q(\D_cache/cache[4][30] ), .QN(n1221) );
  DFFRX1 \D_cache/cache_reg[5][30]  ( .D(\D_cache/n1551 ), .CK(clk), .RN(n6203), .Q(\D_cache/cache[5][30] ), .QN(n2844) );
  DFFRX1 \D_cache/cache_reg[6][30]  ( .D(\D_cache/n1550 ), .CK(clk), .RN(n6203), .Q(\D_cache/cache[6][30] ), .QN(n659) );
  DFFRX1 \D_cache/cache_reg[7][30]  ( .D(\D_cache/n1549 ), .CK(clk), .RN(n6203), .Q(\D_cache/cache[7][30] ), .QN(n2276) );
  DFFRX1 \D_cache/cache_reg[0][31]  ( .D(\D_cache/n1548 ), .CK(clk), .RN(n6202), .Q(\D_cache/cache[0][31] ), .QN(n635) );
  DFFRX1 \D_cache/cache_reg[1][31]  ( .D(\D_cache/n1547 ), .CK(clk), .RN(n6202), .Q(\D_cache/cache[1][31] ), .QN(n2252) );
  DFFRX1 \D_cache/cache_reg[2][31]  ( .D(\D_cache/n1546 ), .CK(clk), .RN(n6202), .Q(\D_cache/cache[2][31] ), .QN(n634) );
  DFFRX1 \D_cache/cache_reg[3][31]  ( .D(\D_cache/n1545 ), .CK(clk), .RN(n6202), .Q(\D_cache/cache[3][31] ), .QN(n2251) );
  DFFRX1 \D_cache/cache_reg[4][31]  ( .D(\D_cache/n1544 ), .CK(clk), .RN(n6202), .Q(\D_cache/cache[4][31] ), .QN(n1219) );
  DFFRX1 \D_cache/cache_reg[5][31]  ( .D(\D_cache/n1543 ), .CK(clk), .RN(n6202), .Q(\D_cache/cache[5][31] ), .QN(n2842) );
  DFFRX1 \D_cache/cache_reg[6][31]  ( .D(\D_cache/n1542 ), .CK(clk), .RN(n6202), .Q(\D_cache/cache[6][31] ), .QN(n633) );
  DFFRX1 \D_cache/cache_reg[7][31]  ( .D(\D_cache/n1541 ), .CK(clk), .RN(n6202), .Q(\D_cache/cache[7][31] ), .QN(n2250) );
  DFFRX1 \D_cache/cache_reg[0][33]  ( .D(\D_cache/n1532 ), .CK(clk), .RN(n6201), .Q(\D_cache/cache[0][33] ), .QN(n1104) );
  DFFRX1 \D_cache/cache_reg[1][33]  ( .D(\D_cache/n1531 ), .CK(clk), .RN(n6201), .Q(\D_cache/cache[1][33] ), .QN(n2727) );
  DFFRX1 \D_cache/cache_reg[2][33]  ( .D(\D_cache/n1530 ), .CK(clk), .RN(n6201), .Q(\D_cache/cache[2][33] ), .QN(n2136) );
  DFFRX1 \D_cache/cache_reg[3][33]  ( .D(\D_cache/n1529 ), .CK(clk), .RN(n6201), .Q(\D_cache/cache[3][33] ), .QN(n511) );
  DFFRX1 \D_cache/cache_reg[4][33]  ( .D(\D_cache/n1528 ), .CK(clk), .RN(n6201), .Q(\D_cache/cache[4][33] ), .QN(n1166) );
  DFFRX1 \D_cache/cache_reg[5][33]  ( .D(\D_cache/n1527 ), .CK(clk), .RN(n6201), .Q(\D_cache/cache[5][33] ), .QN(n2789) );
  DFFRX1 \D_cache/cache_reg[6][33]  ( .D(\D_cache/n1526 ), .CK(clk), .RN(n6201), .Q(\D_cache/cache[6][33] ), .QN(n1103) );
  DFFRX1 \D_cache/cache_reg[7][33]  ( .D(\D_cache/n1525 ), .CK(clk), .RN(n6201), .Q(\D_cache/cache[7][33] ), .QN(n2726) );
  DFFRX1 \D_cache/cache_reg[0][34]  ( .D(\D_cache/n1524 ), .CK(clk), .RN(n6200), .Q(\D_cache/cache[0][34] ), .QN(n648) );
  DFFRX1 \D_cache/cache_reg[1][34]  ( .D(\D_cache/n1523 ), .CK(clk), .RN(n6200), .Q(\D_cache/cache[1][34] ), .QN(n2265) );
  DFFRX1 \D_cache/cache_reg[2][34]  ( .D(\D_cache/n1522 ), .CK(clk), .RN(n6200), .Q(\D_cache/cache[2][34] ), .QN(n2095) );
  DFFRX1 \D_cache/cache_reg[3][34]  ( .D(\D_cache/n1521 ), .CK(clk), .RN(n6200), .Q(\D_cache/cache[3][34] ), .QN(n469) );
  DFFRX1 \D_cache/cache_reg[4][34]  ( .D(\D_cache/n1520 ), .CK(clk), .RN(n6200), .Q(\D_cache/cache[4][34] ), .QN(n1195) );
  DFFRX1 \D_cache/cache_reg[5][34]  ( .D(\D_cache/n1519 ), .CK(clk), .RN(n6200), .Q(\D_cache/cache[5][34] ), .QN(n2818) );
  DFFRX1 \D_cache/cache_reg[6][34]  ( .D(\D_cache/n1518 ), .CK(clk), .RN(n6200), .Q(\D_cache/cache[6][34] ), .QN(n647) );
  DFFRX1 \D_cache/cache_reg[7][34]  ( .D(\D_cache/n1517 ), .CK(clk), .RN(n6200), .Q(\D_cache/cache[7][34] ), .QN(n2264) );
  DFFRX1 \D_cache/cache_reg[0][35]  ( .D(\D_cache/n1516 ), .CK(clk), .RN(n6200), .Q(\D_cache/cache[0][35] ), .QN(n653) );
  DFFRX1 \D_cache/cache_reg[1][35]  ( .D(\D_cache/n1515 ), .CK(clk), .RN(n6200), .Q(\D_cache/cache[1][35] ), .QN(n2270) );
  DFFRX1 \D_cache/cache_reg[2][35]  ( .D(\D_cache/n1514 ), .CK(clk), .RN(n6200), .Q(\D_cache/cache[2][35] ), .QN(n1100) );
  DFFRX1 \D_cache/cache_reg[3][35]  ( .D(\D_cache/n1513 ), .CK(clk), .RN(n6200), .Q(\D_cache/cache[3][35] ), .QN(n2723) );
  DFFRX1 \D_cache/cache_reg[4][35]  ( .D(\D_cache/n1512 ), .CK(clk), .RN(n6199), .Q(\D_cache/cache[4][35] ), .QN(n1087) );
  DFFRX1 \D_cache/cache_reg[5][35]  ( .D(\D_cache/n1511 ), .CK(clk), .RN(n6199), .Q(\D_cache/cache[5][35] ), .QN(n2710) );
  DFFRX1 \D_cache/cache_reg[6][35]  ( .D(\D_cache/n1510 ), .CK(clk), .RN(n6199), .Q(\D_cache/cache[6][35] ), .QN(n652) );
  DFFRX1 \D_cache/cache_reg[7][35]  ( .D(\D_cache/n1509 ), .CK(clk), .RN(n6199), .Q(\D_cache/cache[7][35] ), .QN(n2269) );
  DFFRX1 \D_cache/cache_reg[7][36]  ( .D(\D_cache/n1501 ), .CK(clk), .RN(n6199), .Q(\D_cache/cache[7][36] ), .QN(n564) );
  DFFRX1 \D_cache/cache_reg[0][37]  ( .D(\D_cache/n1500 ), .CK(clk), .RN(n6198), .Q(\D_cache/cache[0][37] ), .QN(n676) );
  DFFRX1 \D_cache/cache_reg[1][37]  ( .D(\D_cache/n1499 ), .CK(clk), .RN(n6198), .Q(\D_cache/cache[1][37] ), .QN(n2294) );
  DFFRX1 \D_cache/cache_reg[2][37]  ( .D(\D_cache/n1498 ), .CK(clk), .RN(n6198), .Q(\D_cache/cache[2][37] ), .QN(n998) );
  DFFRX1 \D_cache/cache_reg[3][37]  ( .D(\D_cache/n1497 ), .CK(clk), .RN(n6198), .Q(\D_cache/cache[3][37] ), .QN(n2623) );
  DFFRX1 \D_cache/cache_reg[4][37]  ( .D(\D_cache/n1496 ), .CK(clk), .RN(n6198), .Q(\D_cache/cache[4][37] ), .QN(n1182) );
  DFFRX1 \D_cache/cache_reg[5][37]  ( .D(\D_cache/n1495 ), .CK(clk), .RN(n6198), .Q(\D_cache/cache[5][37] ), .QN(n2805) );
  DFFRX1 \D_cache/cache_reg[6][37]  ( .D(\D_cache/n1494 ), .CK(clk), .RN(n6198), .Q(\D_cache/cache[6][37] ), .QN(n675) );
  DFFRX1 \D_cache/cache_reg[7][37]  ( .D(\D_cache/n1493 ), .CK(clk), .RN(n6198), .Q(\D_cache/cache[7][37] ), .QN(n2293) );
  DFFRX1 \D_cache/cache_reg[0][38]  ( .D(\D_cache/n1492 ), .CK(clk), .RN(n6198), .Q(\D_cache/cache[0][38] ), .QN(n619) );
  DFFRX1 \D_cache/cache_reg[1][38]  ( .D(\D_cache/n1491 ), .CK(clk), .RN(n6198), .Q(\D_cache/cache[1][38] ), .QN(n2237) );
  DFFRX1 \D_cache/cache_reg[2][38]  ( .D(\D_cache/n1490 ), .CK(clk), .RN(n6198), .Q(\D_cache/cache[2][38] ), .QN(n2094) );
  DFFRX1 \D_cache/cache_reg[3][38]  ( .D(\D_cache/n1489 ), .CK(clk), .RN(n6198), .Q(\D_cache/cache[3][38] ), .QN(n468) );
  DFFRX1 \D_cache/cache_reg[4][38]  ( .D(\D_cache/n1488 ), .CK(clk), .RN(n6197), .Q(\D_cache/cache[4][38] ), .QN(n1215) );
  DFFRX1 \D_cache/cache_reg[5][38]  ( .D(\D_cache/n1487 ), .CK(clk), .RN(n6197), .Q(\D_cache/cache[5][38] ), .QN(n2838) );
  DFFRX1 \D_cache/cache_reg[6][38]  ( .D(\D_cache/n1486 ), .CK(clk), .RN(n6197), .Q(\D_cache/cache[6][38] ), .QN(n1052) );
  DFFRX1 \D_cache/cache_reg[7][38]  ( .D(\D_cache/n1485 ), .CK(clk), .RN(n6197), .Q(\D_cache/cache[7][38] ), .QN(n2679) );
  DFFRX1 \D_cache/cache_reg[0][39]  ( .D(\D_cache/n1484 ), .CK(clk), .RN(n6197), .Q(\D_cache/cache[0][39] ), .QN(n2151) );
  DFFRX1 \D_cache/cache_reg[1][39]  ( .D(\D_cache/n1483 ), .CK(clk), .RN(n6197), .Q(\D_cache/cache[1][39] ), .QN(n526) );
  DFFRX1 \D_cache/cache_reg[2][39]  ( .D(\D_cache/n1482 ), .CK(clk), .RN(n6197), .Q(\D_cache/cache[2][39] ), .QN(n2137) );
  DFFRX1 \D_cache/cache_reg[3][39]  ( .D(\D_cache/n1481 ), .CK(clk), .RN(n6197), .Q(\D_cache/cache[3][39] ), .QN(n512) );
  DFFRX1 \D_cache/cache_reg[4][39]  ( .D(\D_cache/n1480 ), .CK(clk), .RN(n6197), .Q(\D_cache/cache[4][39] ), .QN(n623) );
  DFFRX1 \D_cache/cache_reg[5][39]  ( .D(\D_cache/n1479 ), .CK(clk), .RN(n6197), .Q(\D_cache/cache[5][39] ), .QN(n2241) );
  DFFRX1 \D_cache/cache_reg[6][39]  ( .D(\D_cache/n1478 ), .CK(clk), .RN(n6197), .Q(\D_cache/cache[6][39] ), .QN(n2141) );
  DFFRX1 \D_cache/cache_reg[7][39]  ( .D(\D_cache/n1477 ), .CK(clk), .RN(n6197), .Q(\D_cache/cache[7][39] ), .QN(n516) );
  DFFRX1 \D_cache/cache_reg[0][40]  ( .D(\D_cache/n1476 ), .CK(clk), .RN(n6196), .Q(\D_cache/cache[0][40] ), .QN(n1107) );
  DFFRX1 \D_cache/cache_reg[1][40]  ( .D(\D_cache/n1475 ), .CK(clk), .RN(n6196), .Q(\D_cache/cache[1][40] ), .QN(n2730) );
  DFFRX1 \D_cache/cache_reg[2][40]  ( .D(\D_cache/n1474 ), .CK(clk), .RN(n6196), .Q(\D_cache/cache[2][40] ), .QN(n2091) );
  DFFRX1 \D_cache/cache_reg[3][40]  ( .D(\D_cache/n1473 ), .CK(clk), .RN(n6196), .Q(\D_cache/cache[3][40] ), .QN(n465) );
  DFFRX1 \D_cache/cache_reg[4][40]  ( .D(\D_cache/n1472 ), .CK(clk), .RN(n6196), .Q(\D_cache/cache[4][40] ), .QN(n584) );
  DFFRX1 \D_cache/cache_reg[5][40]  ( .D(\D_cache/n1471 ), .CK(clk), .RN(n6196), .Q(\D_cache/cache[5][40] ), .QN(n2202) );
  DFFRX1 \D_cache/cache_reg[6][40]  ( .D(\D_cache/n1470 ), .CK(clk), .RN(n6196), .Q(\D_cache/cache[6][40] ), .QN(n614) );
  DFFRX1 \D_cache/cache_reg[7][40]  ( .D(\D_cache/n1469 ), .CK(clk), .RN(n6196), .Q(\D_cache/cache[7][40] ), .QN(n2232) );
  DFFRX1 \D_cache/cache_reg[0][42]  ( .D(\D_cache/n1460 ), .CK(clk), .RN(n6195), .Q(\D_cache/cache[0][42] ), .QN(n617) );
  DFFRX1 \D_cache/cache_reg[1][42]  ( .D(\D_cache/n1459 ), .CK(clk), .RN(n6195), .Q(\D_cache/cache[1][42] ), .QN(n2235) );
  DFFRX1 \D_cache/cache_reg[2][42]  ( .D(\D_cache/n1458 ), .CK(clk), .RN(n6195), .Q(\D_cache/cache[2][42] ), .QN(n1108) );
  DFFRX1 \D_cache/cache_reg[3][42]  ( .D(\D_cache/n1457 ), .CK(clk), .RN(n6195), .Q(\D_cache/cache[3][42] ), .QN(n2731) );
  DFFRX1 \D_cache/cache_reg[4][42]  ( .D(\D_cache/n1456 ), .CK(clk), .RN(n6195), .Q(\D_cache/cache[4][42] ), .QN(n1171) );
  DFFRX1 \D_cache/cache_reg[5][42]  ( .D(\D_cache/n1455 ), .CK(clk), .RN(n6195), .Q(\D_cache/cache[5][42] ), .QN(n2794) );
  DFFRX1 \D_cache/cache_reg[6][42]  ( .D(\D_cache/n1454 ), .CK(clk), .RN(n6195), .Q(\D_cache/cache[6][42] ), .QN(n591) );
  DFFRX1 \D_cache/cache_reg[7][42]  ( .D(\D_cache/n1453 ), .CK(clk), .RN(n6195), .Q(\D_cache/cache[7][42] ), .QN(n2209) );
  DFFRX1 \D_cache/cache_reg[0][43]  ( .D(\D_cache/n1452 ), .CK(clk), .RN(n6194), .Q(\D_cache/cache[0][43] ), .QN(n983) );
  DFFRX1 \D_cache/cache_reg[1][43]  ( .D(\D_cache/n1451 ), .CK(clk), .RN(n6194), .Q(\D_cache/cache[1][43] ), .QN(n2608) );
  DFFRX1 \D_cache/cache_reg[2][43]  ( .D(\D_cache/n1450 ), .CK(clk), .RN(n6194), .Q(\D_cache/cache[2][43] ), .QN(n1150) );
  DFFRX1 \D_cache/cache_reg[3][43]  ( .D(\D_cache/n1449 ), .CK(clk), .RN(n6194), .Q(\D_cache/cache[3][43] ), .QN(n2773) );
  DFFRX1 \D_cache/cache_reg[4][43]  ( .D(\D_cache/n1448 ), .CK(clk), .RN(n6194), .Q(\D_cache/cache[4][43] ), .QN(n1168) );
  DFFRX1 \D_cache/cache_reg[5][43]  ( .D(\D_cache/n1447 ), .CK(clk), .RN(n6194), .Q(\D_cache/cache[5][43] ), .QN(n2791) );
  DFFRX1 \D_cache/cache_reg[6][43]  ( .D(\D_cache/n1446 ), .CK(clk), .RN(n6194), .Q(\D_cache/cache[6][43] ), .QN(n1149) );
  DFFRX1 \D_cache/cache_reg[7][43]  ( .D(\D_cache/n1445 ), .CK(clk), .RN(n6194), .Q(\D_cache/cache[7][43] ), .QN(n2772) );
  DFFRX1 \D_cache/cache_reg[0][44]  ( .D(\D_cache/n1444 ), .CK(clk), .RN(n6194), .Q(\D_cache/cache[0][44] ), .QN(n1102) );
  DFFRX1 \D_cache/cache_reg[1][44]  ( .D(\D_cache/n1443 ), .CK(clk), .RN(n6194), .Q(\D_cache/cache[1][44] ), .QN(n2725) );
  DFFRX1 \D_cache/cache_reg[2][44]  ( .D(\D_cache/n1442 ), .CK(clk), .RN(n6194), .Q(\D_cache/cache[2][44] ), .QN(n1101) );
  DFFRX1 \D_cache/cache_reg[3][44]  ( .D(\D_cache/n1441 ), .CK(clk), .RN(n6194), .Q(\D_cache/cache[3][44] ), .QN(n2724) );
  DFFRX1 \D_cache/cache_reg[4][44]  ( .D(\D_cache/n1440 ), .CK(clk), .RN(n6193), .Q(\D_cache/cache[4][44] ), .QN(n1167) );
  DFFRX1 \D_cache/cache_reg[5][44]  ( .D(\D_cache/n1439 ), .CK(clk), .RN(n6193), .Q(\D_cache/cache[5][44] ), .QN(n2790) );
  DFFRX1 \D_cache/cache_reg[6][44]  ( .D(\D_cache/n1438 ), .CK(clk), .RN(n6193), .Q(\D_cache/cache[6][44] ), .QN(n578) );
  DFFRX1 \D_cache/cache_reg[7][44]  ( .D(\D_cache/n1437 ), .CK(clk), .RN(n6193), .Q(\D_cache/cache[7][44] ), .QN(n2196) );
  DFFRX1 \D_cache/cache_reg[0][46]  ( .D(\D_cache/n1428 ), .CK(clk), .RN(n6192), .Q(\D_cache/cache[0][46] ), .QN(n1012) );
  DFFRX1 \D_cache/cache_reg[1][46]  ( .D(\D_cache/n1427 ), .CK(clk), .RN(n6192), .Q(\D_cache/cache[1][46] ), .QN(n2638) );
  DFFRX1 \D_cache/cache_reg[2][46]  ( .D(\D_cache/n1426 ), .CK(clk), .RN(n6192), .Q(\D_cache/cache[2][46] ), .QN(n2072) );
  DFFRX1 \D_cache/cache_reg[3][46]  ( .D(\D_cache/n1425 ), .CK(clk), .RN(n6192), .Q(\D_cache/cache[3][46] ), .QN(n447) );
  DFFRX1 \D_cache/cache_reg[4][46]  ( .D(\D_cache/n1424 ), .CK(clk), .RN(n6192), .Q(\D_cache/cache[4][46] ), .QN(n971) );
  DFFRX1 \D_cache/cache_reg[5][46]  ( .D(\D_cache/n1423 ), .CK(clk), .RN(n6192), .Q(\D_cache/cache[5][46] ), .QN(n2596) );
  DFFRX1 \D_cache/cache_reg[6][46]  ( .D(\D_cache/n1422 ), .CK(clk), .RN(n6192), .Q(\D_cache/cache[6][46] ), .QN(n1011) );
  DFFRX1 \D_cache/cache_reg[7][46]  ( .D(\D_cache/n1421 ), .CK(clk), .RN(n6192), .Q(\D_cache/cache[7][46] ), .QN(n2637) );
  DFFRX1 \D_cache/cache_reg[0][47]  ( .D(\D_cache/n1420 ), .CK(clk), .RN(n6192), .Q(\D_cache/cache[0][47] ), .QN(n1057) );
  DFFRX1 \D_cache/cache_reg[1][47]  ( .D(\D_cache/n1419 ), .CK(clk), .RN(n6192), .Q(\D_cache/cache[1][47] ), .QN(n2684) );
  DFFRX1 \D_cache/cache_reg[2][47]  ( .D(\D_cache/n1418 ), .CK(clk), .RN(n6192), .Q(\D_cache/cache[2][47] ), .QN(n1056) );
  DFFRX1 \D_cache/cache_reg[3][47]  ( .D(\D_cache/n1417 ), .CK(clk), .RN(n6192), .Q(\D_cache/cache[3][47] ), .QN(n2683) );
  DFFRX1 \D_cache/cache_reg[4][47]  ( .D(\D_cache/n1416 ), .CK(clk), .RN(n6191), .Q(\D_cache/cache[4][47] ), .QN(n1213) );
  DFFRX1 \D_cache/cache_reg[5][47]  ( .D(\D_cache/n1415 ), .CK(clk), .RN(n6191), .Q(\D_cache/cache[5][47] ), .QN(n2836) );
  DFFRX1 \D_cache/cache_reg[6][47]  ( .D(\D_cache/n1414 ), .CK(clk), .RN(n6191), .Q(\D_cache/cache[6][47] ), .QN(n1055) );
  DFFRX1 \D_cache/cache_reg[7][47]  ( .D(\D_cache/n1413 ), .CK(clk), .RN(n6191), .Q(\D_cache/cache[7][47] ), .QN(n2682) );
  DFFRX1 \D_cache/cache_reg[0][48]  ( .D(\D_cache/n1412 ), .CK(clk), .RN(n6191), .Q(\D_cache/cache[0][48] ), .QN(n965) );
  DFFRX1 \D_cache/cache_reg[1][48]  ( .D(\D_cache/n1411 ), .CK(clk), .RN(n6191), .Q(\D_cache/cache[1][48] ), .QN(n2590) );
  DFFRX1 \D_cache/cache_reg[2][48]  ( .D(\D_cache/n1410 ), .CK(clk), .RN(n6191), .Q(\D_cache/cache[2][48] ), .QN(n610) );
  DFFRX1 \D_cache/cache_reg[3][48]  ( .D(\D_cache/n1409 ), .CK(clk), .RN(n6191), .Q(\D_cache/cache[3][48] ), .QN(n2228) );
  DFFRX1 \D_cache/cache_reg[4][48]  ( .D(\D_cache/n1408 ), .CK(clk), .RN(n6191), .Q(\D_cache/cache[4][48] ), .QN(n575) );
  DFFRX1 \D_cache/cache_reg[5][48]  ( .D(\D_cache/n1407 ), .CK(clk), .RN(n6191), .Q(\D_cache/cache[5][48] ), .QN(n2193) );
  DFFRX1 \D_cache/cache_reg[6][48]  ( .D(\D_cache/n1406 ), .CK(clk), .RN(n6191), .Q(\D_cache/cache[6][48] ), .QN(n621) );
  DFFRX1 \D_cache/cache_reg[7][48]  ( .D(\D_cache/n1405 ), .CK(clk), .RN(n6191), .Q(\D_cache/cache[7][48] ), .QN(n2239) );
  DFFRX1 \D_cache/cache_reg[0][49]  ( .D(\D_cache/n1404 ), .CK(clk), .RN(n6190), .Q(\D_cache/cache[0][49] ), .QN(n1155) );
  DFFRX1 \D_cache/cache_reg[1][49]  ( .D(\D_cache/n1403 ), .CK(clk), .RN(n6190), .Q(\D_cache/cache[1][49] ), .QN(n2778) );
  DFFRX1 \D_cache/cache_reg[2][49]  ( .D(\D_cache/n1402 ), .CK(clk), .RN(n6190), .Q(\D_cache/cache[2][49] ), .QN(n1154) );
  DFFRX1 \D_cache/cache_reg[3][49]  ( .D(\D_cache/n1401 ), .CK(clk), .RN(n6190), .Q(\D_cache/cache[3][49] ), .QN(n2777) );
  DFFRX1 \D_cache/cache_reg[4][49]  ( .D(\D_cache/n1400 ), .CK(clk), .RN(n6190), .Q(\D_cache/cache[4][49] ), .QN(n1181) );
  DFFRX1 \D_cache/cache_reg[5][49]  ( .D(\D_cache/n1399 ), .CK(clk), .RN(n6190), .Q(\D_cache/cache[5][49] ), .QN(n2804) );
  DFFRX1 \D_cache/cache_reg[6][49]  ( .D(\D_cache/n1398 ), .CK(clk), .RN(n6190), .Q(\D_cache/cache[6][49] ), .QN(n1153) );
  DFFRX1 \D_cache/cache_reg[7][49]  ( .D(\D_cache/n1397 ), .CK(clk), .RN(n6190), .Q(\D_cache/cache[7][49] ), .QN(n2776) );
  DFFRX1 \D_cache/cache_reg[0][53]  ( .D(\D_cache/n1372 ), .CK(clk), .RN(n6188), .Q(\D_cache/cache[0][53] ), .QN(n2148) );
  DFFRX1 \D_cache/cache_reg[1][53]  ( .D(\D_cache/n1371 ), .CK(clk), .RN(n6188), .Q(\D_cache/cache[1][53] ), .QN(n523) );
  DFFRX1 \D_cache/cache_reg[2][53]  ( .D(\D_cache/n1370 ), .CK(clk), .RN(n6188), .Q(\D_cache/cache[2][53] ), .QN(n613) );
  DFFRX1 \D_cache/cache_reg[3][53]  ( .D(\D_cache/n1369 ), .CK(clk), .RN(n6188), .Q(\D_cache/cache[3][53] ), .QN(n2231) );
  DFFRX1 \D_cache/cache_reg[4][53]  ( .D(\D_cache/n1368 ), .CK(clk), .RN(n6187), .Q(\D_cache/cache[4][53] ), .QN(n622) );
  DFFRX1 \D_cache/cache_reg[5][53]  ( .D(\D_cache/n1367 ), .CK(clk), .RN(n6187), .Q(\D_cache/cache[5][53] ), .QN(n2240) );
  DFFRX1 \D_cache/cache_reg[6][53]  ( .D(\D_cache/n1366 ), .CK(clk), .RN(n6187), .Q(\D_cache/cache[6][53] ), .QN(n2142) );
  DFFRX1 \D_cache/cache_reg[7][53]  ( .D(\D_cache/n1365 ), .CK(clk), .RN(n6187), .Q(\D_cache/cache[7][53] ), .QN(n517) );
  DFFRX1 \D_cache/cache_reg[0][54]  ( .D(\D_cache/n1364 ), .CK(clk), .RN(n6187), .Q(\D_cache/cache[0][54] ), .QN(n1229) );
  DFFRX1 \D_cache/cache_reg[1][54]  ( .D(\D_cache/n1363 ), .CK(clk), .RN(n6187), .Q(\D_cache/cache[1][54] ), .QN(n2852) );
  DFFRX1 \D_cache/cache_reg[2][54]  ( .D(\D_cache/n1362 ), .CK(clk), .RN(n6187), .Q(\D_cache/cache[2][54] ), .QN(n972) );
  DFFRX1 \D_cache/cache_reg[3][54]  ( .D(\D_cache/n1361 ), .CK(clk), .RN(n6187), .Q(\D_cache/cache[3][54] ), .QN(n2597) );
  DFFRX1 \D_cache/cache_reg[4][54]  ( .D(\D_cache/n1360 ), .CK(clk), .RN(n6187), .Q(\D_cache/cache[4][54] ), .QN(n1211) );
  DFFRX1 \D_cache/cache_reg[5][54]  ( .D(\D_cache/n1359 ), .CK(clk), .RN(n6187), .Q(\D_cache/cache[5][54] ), .QN(n2834) );
  DFFRX1 \D_cache/cache_reg[6][54]  ( .D(\D_cache/n1358 ), .CK(clk), .RN(n6187), .Q(\D_cache/cache[6][54] ), .QN(n1228) );
  DFFRX1 \D_cache/cache_reg[7][54]  ( .D(\D_cache/n1357 ), .CK(clk), .RN(n6187), .Q(\D_cache/cache[7][54] ), .QN(n2851) );
  DFFRX1 \D_cache/cache_reg[0][55]  ( .D(\D_cache/n1356 ), .CK(clk), .RN(n6186), .Q(\D_cache/cache[0][55] ), .QN(n667) );
  DFFRX1 \D_cache/cache_reg[1][55]  ( .D(\D_cache/n1355 ), .CK(clk), .RN(n6186), .Q(\D_cache/cache[1][55] ), .QN(n2285) );
  DFFRX1 \D_cache/cache_reg[2][55]  ( .D(\D_cache/n1354 ), .CK(clk), .RN(n6186), .Q(\D_cache/cache[2][55] ), .QN(n993) );
  DFFRX1 \D_cache/cache_reg[3][55]  ( .D(\D_cache/n1353 ), .CK(clk), .RN(n6186), .Q(\D_cache/cache[3][55] ), .QN(n2618) );
  DFFRX1 \D_cache/cache_reg[4][55]  ( .D(\D_cache/n1352 ), .CK(clk), .RN(n6186), .Q(\D_cache/cache[4][55] ), .QN(n1084) );
  DFFRX1 \D_cache/cache_reg[5][55]  ( .D(\D_cache/n1351 ), .CK(clk), .RN(n6186), .Q(\D_cache/cache[5][55] ), .QN(n2707) );
  DFFRX1 \D_cache/cache_reg[6][55]  ( .D(\D_cache/n1350 ), .CK(clk), .RN(n6186), .Q(\D_cache/cache[6][55] ), .QN(n666) );
  DFFRX1 \D_cache/cache_reg[7][55]  ( .D(\D_cache/n1349 ), .CK(clk), .RN(n6186), .Q(\D_cache/cache[7][55] ), .QN(n2284) );
  DFFRX1 \D_cache/cache_reg[0][58]  ( .D(\D_cache/n1332 ), .CK(clk), .RN(n6184), .Q(\D_cache/cache[0][58] ), .QN(n618) );
  DFFRX1 \D_cache/cache_reg[1][58]  ( .D(\D_cache/n1331 ), .CK(clk), .RN(n6184), .Q(\D_cache/cache[1][58] ), .QN(n2236) );
  DFFRX1 \D_cache/cache_reg[2][58]  ( .D(\D_cache/n1330 ), .CK(clk), .RN(n6184), .Q(\D_cache/cache[2][58] ), .QN(n1086) );
  DFFRX1 \D_cache/cache_reg[3][58]  ( .D(\D_cache/n1329 ), .CK(clk), .RN(n6184), .Q(\D_cache/cache[3][58] ), .QN(n2709) );
  DFFRX1 \D_cache/cache_reg[5][58]  ( .D(\D_cache/n1327 ), .CK(clk), .RN(n6184), .Q(\D_cache/cache[5][58] ), .QN(n2033) );
  DFFRX1 \D_cache/cache_reg[6][58]  ( .D(\D_cache/n1326 ), .CK(clk), .RN(n6184), .Q(\D_cache/cache[6][58] ), .QN(n978) );
  DFFRX1 \D_cache/cache_reg[7][58]  ( .D(\D_cache/n1325 ), .CK(clk), .RN(n6184), .Q(\D_cache/cache[7][58] ), .QN(n2603) );
  DFFRX1 \D_cache/cache_reg[0][59]  ( .D(\D_cache/n1324 ), .CK(clk), .RN(n6184), .Q(\D_cache/cache[0][59] ), .QN(n682) );
  DFFRX1 \D_cache/cache_reg[1][59]  ( .D(\D_cache/n1323 ), .CK(clk), .RN(n6184), .Q(\D_cache/cache[1][59] ), .QN(n2300) );
  DFFRX1 \D_cache/cache_reg[2][59]  ( .D(\D_cache/n1322 ), .CK(clk), .RN(n6184), .Q(\D_cache/cache[2][59] ), .QN(n1000) );
  DFFRX1 \D_cache/cache_reg[3][59]  ( .D(\D_cache/n1321 ), .CK(clk), .RN(n6184), .Q(\D_cache/cache[3][59] ), .QN(n2625) );
  DFFRX1 \D_cache/cache_reg[4][59]  ( .D(\D_cache/n1320 ), .CK(clk), .RN(n6183), .Q(\D_cache/cache[4][59] ), .QN(n1193) );
  DFFRX1 \D_cache/cache_reg[5][59]  ( .D(\D_cache/n1319 ), .CK(clk), .RN(n6183), .Q(\D_cache/cache[5][59] ), .QN(n2816) );
  DFFRX1 \D_cache/cache_reg[6][59]  ( .D(\D_cache/n1318 ), .CK(clk), .RN(n6183), .Q(\D_cache/cache[6][59] ), .QN(n681) );
  DFFRX1 \D_cache/cache_reg[7][59]  ( .D(\D_cache/n1317 ), .CK(clk), .RN(n6183), .Q(\D_cache/cache[7][59] ), .QN(n2299) );
  DFFRX1 \D_cache/cache_reg[0][60]  ( .D(\D_cache/n1316 ), .CK(clk), .RN(n6183), .Q(\D_cache/cache[0][60] ), .QN(n671) );
  DFFRX1 \D_cache/cache_reg[1][60]  ( .D(\D_cache/n1315 ), .CK(clk), .RN(n6183), .Q(\D_cache/cache[1][60] ), .QN(n2289) );
  DFFRX1 \D_cache/cache_reg[2][60]  ( .D(\D_cache/n1314 ), .CK(clk), .RN(n6183), .Q(\D_cache/cache[2][60] ), .QN(n995) );
  DFFRX1 \D_cache/cache_reg[3][60]  ( .D(\D_cache/n1313 ), .CK(clk), .RN(n6183), .Q(\D_cache/cache[3][60] ), .QN(n2620) );
  DFFRX1 \D_cache/cache_reg[4][60]  ( .D(\D_cache/n1312 ), .CK(clk), .RN(n6183), .Q(\D_cache/cache[4][60] ), .QN(n2150) );
  DFFRX1 \D_cache/cache_reg[5][60]  ( .D(\D_cache/n1311 ), .CK(clk), .RN(n6183), .Q(\D_cache/cache[5][60] ), .QN(n525) );
  DFFRX1 \D_cache/cache_reg[6][60]  ( .D(\D_cache/n1310 ), .CK(clk), .RN(n6183), .Q(\D_cache/cache[6][60] ), .QN(n670) );
  DFFRX1 \D_cache/cache_reg[7][60]  ( .D(\D_cache/n1309 ), .CK(clk), .RN(n6183), .Q(\D_cache/cache[7][60] ), .QN(n2288) );
  DFFRX1 \D_cache/cache_reg[0][61]  ( .D(\D_cache/n1308 ), .CK(clk), .RN(n6182), .Q(\D_cache/cache[0][61] ), .QN(n1224) );
  DFFRX1 \D_cache/cache_reg[1][61]  ( .D(\D_cache/n1307 ), .CK(clk), .RN(n6182), .Q(\D_cache/cache[1][61] ), .QN(n2847) );
  DFFRX1 \D_cache/cache_reg[2][61]  ( .D(\D_cache/n1306 ), .CK(clk), .RN(n6182), .Q(\D_cache/cache[2][61] ), .QN(n996) );
  DFFRX1 \D_cache/cache_reg[3][61]  ( .D(\D_cache/n1305 ), .CK(clk), .RN(n6182), .Q(\D_cache/cache[3][61] ), .QN(n2621) );
  DFFRX1 \D_cache/cache_reg[4][61]  ( .D(\D_cache/n1304 ), .CK(clk), .RN(n6182), .Q(\D_cache/cache[4][61] ), .QN(n1284) );
  DFFRX1 \D_cache/cache_reg[5][61]  ( .D(\D_cache/n1303 ), .CK(clk), .RN(n6182), .Q(\D_cache/cache[5][61] ), .QN(n2916) );
  DFFRX1 \D_cache/cache_reg[6][61]  ( .D(\D_cache/n1302 ), .CK(clk), .RN(n6182), .Q(\D_cache/cache[6][61] ), .QN(n672) );
  DFFRX1 \D_cache/cache_reg[7][61]  ( .D(\D_cache/n1301 ), .CK(clk), .RN(n6182), .Q(\D_cache/cache[7][61] ), .QN(n2290) );
  DFFRX1 \D_cache/cache_reg[0][62]  ( .D(\D_cache/n1300 ), .CK(clk), .RN(n6182), .Q(\D_cache/cache[0][62] ), .QN(n656) );
  DFFRX1 \D_cache/cache_reg[1][62]  ( .D(\D_cache/n1299 ), .CK(clk), .RN(n6182), .Q(\D_cache/cache[1][62] ), .QN(n2273) );
  DFFRX1 \D_cache/cache_reg[2][62]  ( .D(\D_cache/n1298 ), .CK(clk), .RN(n6182), .Q(\D_cache/cache[2][62] ), .QN(n655) );
  DFFRX1 \D_cache/cache_reg[3][62]  ( .D(\D_cache/n1297 ), .CK(clk), .RN(n6182), .Q(\D_cache/cache[3][62] ), .QN(n2272) );
  DFFRX1 \D_cache/cache_reg[4][62]  ( .D(\D_cache/n1296 ), .CK(clk), .RN(n6181), .Q(\D_cache/cache[4][62] ), .QN(n1220) );
  DFFRX1 \D_cache/cache_reg[5][62]  ( .D(\D_cache/n1295 ), .CK(clk), .RN(n6181), .Q(\D_cache/cache[5][62] ), .QN(n2843) );
  DFFRX1 \D_cache/cache_reg[6][62]  ( .D(\D_cache/n1294 ), .CK(clk), .RN(n6181), .Q(\D_cache/cache[6][62] ), .QN(n654) );
  DFFRX1 \D_cache/cache_reg[7][62]  ( .D(\D_cache/n1293 ), .CK(clk), .RN(n6181), .Q(\D_cache/cache[7][62] ), .QN(n2271) );
  DFFRX1 \D_cache/cache_reg[0][64]  ( .D(\D_cache/n1284 ), .CK(clk), .RN(n6180), .Q(\D_cache/cache[0][64] ), .QN(n699) );
  DFFRX1 \D_cache/cache_reg[1][64]  ( .D(\D_cache/n1283 ), .CK(clk), .RN(n6180), .Q(\D_cache/cache[1][64] ), .QN(n2317) );
  DFFRX1 \D_cache/cache_reg[2][64]  ( .D(\D_cache/n1282 ), .CK(clk), .RN(n6180), .Q(\D_cache/cache[2][64] ), .QN(n1019) );
  DFFRX1 \D_cache/cache_reg[3][64]  ( .D(\D_cache/n1281 ), .CK(clk), .RN(n6180), .Q(\D_cache/cache[3][64] ), .QN(n2645) );
  DFFRX1 \D_cache/cache_reg[4][64]  ( .D(\D_cache/n1280 ), .CK(clk), .RN(n6180), .Q(\D_cache/cache[4][64] ), .QN(n1191) );
  DFFRX1 \D_cache/cache_reg[5][64]  ( .D(\D_cache/n1279 ), .CK(clk), .RN(n6180), .Q(\D_cache/cache[5][64] ), .QN(n2814) );
  DFFRX1 \D_cache/cache_reg[6][64]  ( .D(\D_cache/n1278 ), .CK(clk), .RN(n6180), .Q(\D_cache/cache[6][64] ), .QN(n698) );
  DFFRX1 \D_cache/cache_reg[7][64]  ( .D(\D_cache/n1277 ), .CK(clk), .RN(n6180), .Q(\D_cache/cache[7][64] ), .QN(n2316) );
  DFFRX1 \D_cache/cache_reg[0][65]  ( .D(\D_cache/n1276 ), .CK(clk), .RN(n6180), .Q(\D_cache/cache[0][65] ), .QN(n694) );
  DFFRX1 \D_cache/cache_reg[1][65]  ( .D(\D_cache/n1275 ), .CK(clk), .RN(n6180), .Q(\D_cache/cache[1][65] ), .QN(n2312) );
  DFFRX1 \D_cache/cache_reg[2][65]  ( .D(\D_cache/n1274 ), .CK(clk), .RN(n6180), .Q(\D_cache/cache[2][65] ), .QN(n2133) );
  DFFRX1 \D_cache/cache_reg[3][65]  ( .D(\D_cache/n1273 ), .CK(clk), .RN(n6180), .Q(\D_cache/cache[3][65] ), .QN(n508) );
  DFFRX1 \D_cache/cache_reg[4][65]  ( .D(\D_cache/n1272 ), .CK(clk), .RN(n6179), .Q(\D_cache/cache[4][65] ), .QN(n1183) );
  DFFRX1 \D_cache/cache_reg[5][65]  ( .D(\D_cache/n1271 ), .CK(clk), .RN(n6179), .Q(\D_cache/cache[5][65] ), .QN(n2806) );
  DFFRX1 \D_cache/cache_reg[6][65]  ( .D(\D_cache/n1270 ), .CK(clk), .RN(n6179), .Q(\D_cache/cache[6][65] ), .QN(n693) );
  DFFRX1 \D_cache/cache_reg[7][65]  ( .D(\D_cache/n1269 ), .CK(clk), .RN(n6179), .Q(\D_cache/cache[7][65] ), .QN(n2311) );
  DFFRX1 \D_cache/cache_reg[0][66]  ( .D(\D_cache/n1268 ), .CK(clk), .RN(n6179), .Q(\D_cache/cache[0][66] ), .QN(n1042) );
  DFFRX1 \D_cache/cache_reg[1][66]  ( .D(\D_cache/n1267 ), .CK(clk), .RN(n6179), .Q(\D_cache/cache[1][66] ), .QN(n2669) );
  DFFRX1 \D_cache/cache_reg[2][66]  ( .D(\D_cache/n1266 ), .CK(clk), .RN(n6179), .Q(\D_cache/cache[2][66] ), .QN(n2098) );
  DFFRX1 \D_cache/cache_reg[3][66]  ( .D(\D_cache/n1265 ), .CK(clk), .RN(n6179), .Q(\D_cache/cache[3][66] ), .QN(n472) );
  DFFRX1 \D_cache/cache_reg[4][66]  ( .D(\D_cache/n1264 ), .CK(clk), .RN(n6179), .Q(\D_cache/cache[4][66] ), .QN(n1209) );
  DFFRX1 \D_cache/cache_reg[5][66]  ( .D(\D_cache/n1263 ), .CK(clk), .RN(n6179), .Q(\D_cache/cache[5][66] ), .QN(n2832) );
  DFFRX1 \D_cache/cache_reg[6][66]  ( .D(\D_cache/n1262 ), .CK(clk), .RN(n6179), .Q(\D_cache/cache[6][66] ), .QN(n602) );
  DFFRX1 \D_cache/cache_reg[7][66]  ( .D(\D_cache/n1261 ), .CK(clk), .RN(n6179), .Q(\D_cache/cache[7][66] ), .QN(n2220) );
  DFFRX1 \D_cache/cache_reg[0][67]  ( .D(\D_cache/n1260 ), .CK(clk), .RN(n6178), .Q(\D_cache/cache[0][67] ), .QN(n560) );
  DFFRX1 \D_cache/cache_reg[1][67]  ( .D(\D_cache/n1259 ), .CK(clk), .RN(n6178), .Q(\D_cache/cache[1][67] ), .QN(n2181) );
  DFFRX1 \D_cache/cache_reg[2][67]  ( .D(\D_cache/n1258 ), .CK(clk), .RN(n6178), .Q(\D_cache/cache[2][67] ), .QN(n1018) );
  DFFRX1 \D_cache/cache_reg[3][67]  ( .D(\D_cache/n1257 ), .CK(clk), .RN(n6178), .Q(\D_cache/cache[3][67] ), .QN(n2644) );
  DFFRX1 \D_cache/cache_reg[4][67]  ( .D(\D_cache/n1256 ), .CK(clk), .RN(n6178), .Q(\D_cache/cache[4][67] ), .QN(n1278) );
  DFFRX1 \D_cache/cache_reg[5][67]  ( .D(\D_cache/n1255 ), .CK(clk), .RN(n6178), .Q(\D_cache/cache[5][67] ), .QN(n2910) );
  DFFRX1 \D_cache/cache_reg[6][67]  ( .D(\D_cache/n1254 ), .CK(clk), .RN(n6178), .Q(\D_cache/cache[6][67] ), .QN(n697) );
  DFFRX1 \D_cache/cache_reg[7][67]  ( .D(\D_cache/n1253 ), .CK(clk), .RN(n6178), .Q(\D_cache/cache[7][67] ), .QN(n2315) );
  DFFRX1 \D_cache/cache_reg[0][68]  ( .D(\D_cache/n1252 ), .CK(clk), .RN(n6178), .Q(\D_cache/cache[0][68] ), .QN(n567) );
  DFFRX1 \D_cache/cache_reg[1][68]  ( .D(\D_cache/n1251 ), .CK(clk), .RN(n6178), .Q(\D_cache/cache[1][68] ), .QN(n2319) );
  DFFRX1 \D_cache/cache_reg[2][68]  ( .D(\D_cache/n1250 ), .CK(clk), .RN(n6178), .Q(\D_cache/cache[2][68] ), .QN(n600) );
  DFFRX1 \D_cache/cache_reg[3][68]  ( .D(\D_cache/n1249 ), .CK(clk), .RN(n6178), .Q(\D_cache/cache[3][68] ), .QN(n2218) );
  DFFRX1 \D_cache/cache_reg[4][68]  ( .D(\D_cache/n1248 ), .CK(clk), .RN(n6177), .Q(\D_cache/cache[4][68] ), .QN(n1075) );
  DFFRX1 \D_cache/cache_reg[5][68]  ( .D(\D_cache/n1247 ), .CK(clk), .RN(n6177), .Q(\D_cache/cache[5][68] ), .QN(n2581) );
  DFFRX1 \D_cache/cache_reg[6][68]  ( .D(\D_cache/n1246 ), .CK(clk), .RN(n6177), .Q(\D_cache/cache[6][68] ), .QN(n566) );
  DFFRX1 \D_cache/cache_reg[7][68]  ( .D(\D_cache/n1245 ), .CK(clk), .RN(n6177), .Q(\D_cache/cache[7][68] ), .QN(n2318) );
  DFFRX1 \D_cache/cache_reg[0][69]  ( .D(\D_cache/n1244 ), .CK(clk), .RN(n6177), .Q(\D_cache/cache[0][69] ), .QN(n1035) );
  DFFRX1 \D_cache/cache_reg[1][69]  ( .D(\D_cache/n1243 ), .CK(clk), .RN(n6177), .Q(\D_cache/cache[1][69] ), .QN(n2661) );
  DFFRX1 \D_cache/cache_reg[2][69]  ( .D(\D_cache/n1242 ), .CK(clk), .RN(n6177), .Q(\D_cache/cache[2][69] ), .QN(n1034) );
  DFFRX1 \D_cache/cache_reg[3][69]  ( .D(\D_cache/n1241 ), .CK(clk), .RN(n6177), .Q(\D_cache/cache[3][69] ), .QN(n2660) );
  DFFRX1 \D_cache/cache_reg[4][69]  ( .D(\D_cache/n1240 ), .CK(clk), .RN(n6177), .Q(\D_cache/cache[4][69] ), .QN(n986) );
  DFFRX1 \D_cache/cache_reg[5][69]  ( .D(\D_cache/n1239 ), .CK(clk), .RN(n6177), .Q(\D_cache/cache[5][69] ), .QN(n2611) );
  DFFRX1 \D_cache/cache_reg[6][69]  ( .D(\D_cache/n1238 ), .CK(clk), .RN(n6177), .Q(\D_cache/cache[6][69] ), .QN(n2080) );
  DFFRX1 \D_cache/cache_reg[7][69]  ( .D(\D_cache/n1237 ), .CK(clk), .RN(n6177), .Q(\D_cache/cache[7][69] ), .QN(n455) );
  DFFRX1 \D_cache/cache_reg[0][70]  ( .D(\D_cache/n1236 ), .CK(clk), .RN(n6176), .Q(\D_cache/cache[0][70] ), .QN(n1047) );
  DFFRX1 \D_cache/cache_reg[1][70]  ( .D(\D_cache/n1235 ), .CK(clk), .RN(n6176), .Q(\D_cache/cache[1][70] ), .QN(n2674) );
  DFFRX1 \D_cache/cache_reg[2][70]  ( .D(\D_cache/n1234 ), .CK(clk), .RN(n6176), .Q(\D_cache/cache[2][70] ), .QN(n1046) );
  DFFRX1 \D_cache/cache_reg[3][70]  ( .D(\D_cache/n1233 ), .CK(clk), .RN(n6176), .Q(\D_cache/cache[3][70] ), .QN(n2673) );
  DFFRX1 \D_cache/cache_reg[4][70]  ( .D(\D_cache/n1232 ), .CK(clk), .RN(n6176), .Q(\D_cache/cache[4][70] ), .QN(n1212) );
  DFFRX1 \D_cache/cache_reg[5][70]  ( .D(\D_cache/n1231 ), .CK(clk), .RN(n6176), .Q(\D_cache/cache[5][70] ), .QN(n2835) );
  DFFRX1 \D_cache/cache_reg[6][70]  ( .D(\D_cache/n1230 ), .CK(clk), .RN(n6176), .Q(\D_cache/cache[6][70] ), .QN(n2107) );
  DFFRX1 \D_cache/cache_reg[7][70]  ( .D(\D_cache/n1229 ), .CK(clk), .RN(n6176), .Q(\D_cache/cache[7][70] ), .QN(n481) );
  DFFRX1 \D_cache/cache_reg[0][71]  ( .D(\D_cache/n1228 ), .CK(clk), .RN(n6176), .Q(\D_cache/cache[0][71] ), .QN(n1033) );
  DFFRX1 \D_cache/cache_reg[1][71]  ( .D(\D_cache/n1227 ), .CK(clk), .RN(n6176), .Q(\D_cache/cache[1][71] ), .QN(n2659) );
  DFFRX1 \D_cache/cache_reg[2][71]  ( .D(\D_cache/n1226 ), .CK(clk), .RN(n6176), .Q(\D_cache/cache[2][71] ), .QN(n1032) );
  DFFRX1 \D_cache/cache_reg[3][71]  ( .D(\D_cache/n1225 ), .CK(clk), .RN(n6176), .Q(\D_cache/cache[3][71] ), .QN(n2658) );
  DFFRX1 \D_cache/cache_reg[4][71]  ( .D(\D_cache/n1224 ), .CK(clk), .RN(n6175), .Q(\D_cache/cache[4][71] ), .QN(n1208) );
  DFFRX1 \D_cache/cache_reg[5][71]  ( .D(\D_cache/n1223 ), .CK(clk), .RN(n6175), .Q(\D_cache/cache[5][71] ), .QN(n2831) );
  DFFRX1 \D_cache/cache_reg[6][71]  ( .D(\D_cache/n1222 ), .CK(clk), .RN(n6175), .Q(\D_cache/cache[6][71] ), .QN(n1031) );
  DFFRX1 \D_cache/cache_reg[7][71]  ( .D(\D_cache/n1221 ), .CK(clk), .RN(n6175), .Q(\D_cache/cache[7][71] ), .QN(n2657) );
  DFFRX1 \D_cache/cache_reg[0][72]  ( .D(\D_cache/n1220 ), .CK(clk), .RN(n6175), .Q(\D_cache/cache[0][72] ), .QN(n706) );
  DFFRX1 \D_cache/cache_reg[1][72]  ( .D(\D_cache/n1219 ), .CK(clk), .RN(n6175), .Q(\D_cache/cache[1][72] ), .QN(n2326) );
  DFFRX1 \D_cache/cache_reg[2][72]  ( .D(\D_cache/n1218 ), .CK(clk), .RN(n6175), .Q(\D_cache/cache[2][72] ), .QN(n1024) );
  DFFRX1 \D_cache/cache_reg[3][72]  ( .D(\D_cache/n1217 ), .CK(clk), .RN(n6175), .Q(\D_cache/cache[3][72] ), .QN(n2650) );
  DFFRX1 \D_cache/cache_reg[4][72]  ( .D(\D_cache/n1216 ), .CK(clk), .RN(n6175), .Q(\D_cache/cache[4][72] ), .QN(n592) );
  DFFRX1 \D_cache/cache_reg[5][72]  ( .D(\D_cache/n1215 ), .CK(clk), .RN(n6175), .Q(\D_cache/cache[5][72] ), .QN(n2210) );
  DFFRX1 \D_cache/cache_reg[6][72]  ( .D(\D_cache/n1214 ), .CK(clk), .RN(n6175), .Q(\D_cache/cache[6][72] ), .QN(n705) );
  DFFRX1 \D_cache/cache_reg[7][72]  ( .D(\D_cache/n1213 ), .CK(clk), .RN(n6175), .Q(\D_cache/cache[7][72] ), .QN(n2325) );
  DFFRX1 \D_cache/cache_reg[0][73]  ( .D(\D_cache/n1212 ), .CK(clk), .RN(n6174), .Q(\D_cache/cache[0][73] ), .QN(n1027) );
  DFFRX1 \D_cache/cache_reg[1][73]  ( .D(\D_cache/n1211 ), .CK(clk), .RN(n6174), .Q(\D_cache/cache[1][73] ), .QN(n2653) );
  DFFRX1 \D_cache/cache_reg[2][73]  ( .D(\D_cache/n1210 ), .CK(clk), .RN(n6174), .Q(\D_cache/cache[2][73] ), .QN(n1026) );
  DFFRX1 \D_cache/cache_reg[3][73]  ( .D(\D_cache/n1209 ), .CK(clk), .RN(n6174), .Q(\D_cache/cache[3][73] ), .QN(n2652) );
  DFFRX1 \D_cache/cache_reg[4][73]  ( .D(\D_cache/n1208 ), .CK(clk), .RN(n6174), .Q(\D_cache/cache[4][73] ), .QN(n1197) );
  DFFRX1 \D_cache/cache_reg[5][73]  ( .D(\D_cache/n1207 ), .CK(clk), .RN(n6174), .Q(\D_cache/cache[5][73] ), .QN(n2820) );
  DFFRX1 \D_cache/cache_reg[6][73]  ( .D(\D_cache/n1206 ), .CK(clk), .RN(n6174), .Q(\D_cache/cache[6][73] ), .QN(n1025) );
  DFFRX1 \D_cache/cache_reg[7][73]  ( .D(\D_cache/n1205 ), .CK(clk), .RN(n6174), .Q(\D_cache/cache[7][73] ), .QN(n2651) );
  DFFRX1 \D_cache/cache_reg[0][74]  ( .D(\D_cache/n1204 ), .CK(clk), .RN(n6174), .Q(\D_cache/cache[0][74] ), .QN(n558) );
  DFFRX1 \D_cache/cache_reg[1][74]  ( .D(\D_cache/n1203 ), .CK(clk), .RN(n6174), .Q(\D_cache/cache[1][74] ), .QN(n2179) );
  DFFRX1 \D_cache/cache_reg[2][74]  ( .D(\D_cache/n1202 ), .CK(clk), .RN(n6174), .Q(\D_cache/cache[2][74] ), .QN(n1081) );
  DFFRX1 \D_cache/cache_reg[3][74]  ( .D(\D_cache/n1201 ), .CK(clk), .RN(n6174), .Q(\D_cache/cache[3][74] ), .QN(n2704) );
  DFFRX1 \D_cache/cache_reg[4][74]  ( .D(\D_cache/n1200 ), .CK(clk), .RN(n6173), .Q(\D_cache/cache[4][74] ), .QN(n1276) );
  DFFRX1 \D_cache/cache_reg[5][74]  ( .D(\D_cache/n1199 ), .CK(clk), .RN(n6173), .Q(\D_cache/cache[5][74] ), .QN(n2908) );
  DFFRX1 \D_cache/cache_reg[6][74]  ( .D(\D_cache/n1198 ), .CK(clk), .RN(n6173), .Q(\D_cache/cache[6][74] ), .QN(n707) );
  DFFRX1 \D_cache/cache_reg[7][74]  ( .D(\D_cache/n1197 ), .CK(clk), .RN(n6173), .Q(\D_cache/cache[7][74] ), .QN(n2327) );
  DFFRX1 \D_cache/cache_reg[0][75]  ( .D(\D_cache/n1196 ), .CK(clk), .RN(n6173), .Q(\D_cache/cache[0][75] ), .QN(n701) );
  DFFRX1 \D_cache/cache_reg[1][75]  ( .D(\D_cache/n1195 ), .CK(clk), .RN(n6173), .Q(\D_cache/cache[1][75] ), .QN(n2321) );
  DFFRX1 \D_cache/cache_reg[2][75]  ( .D(\D_cache/n1194 ), .CK(clk), .RN(n6173), .Q(\D_cache/cache[2][75] ), .QN(n1020) );
  DFFRX1 \D_cache/cache_reg[3][75]  ( .D(\D_cache/n1193 ), .CK(clk), .RN(n6173), .Q(\D_cache/cache[3][75] ), .QN(n2646) );
  DFFRX1 \D_cache/cache_reg[4][75]  ( .D(\D_cache/n1192 ), .CK(clk), .RN(n6173), .Q(\D_cache/cache[4][75] ), .QN(n1186) );
  DFFRX1 \D_cache/cache_reg[5][75]  ( .D(\D_cache/n1191 ), .CK(clk), .RN(n6173), .Q(\D_cache/cache[5][75] ), .QN(n2809) );
  DFFRX1 \D_cache/cache_reg[6][75]  ( .D(\D_cache/n1190 ), .CK(clk), .RN(n6173), .Q(\D_cache/cache[6][75] ), .QN(n700) );
  DFFRX1 \D_cache/cache_reg[7][75]  ( .D(\D_cache/n1189 ), .CK(clk), .RN(n6173), .Q(\D_cache/cache[7][75] ), .QN(n2320) );
  DFFRX1 \D_cache/cache_reg[0][76]  ( .D(\D_cache/n1188 ), .CK(clk), .RN(n6172), .Q(\D_cache/cache[0][76] ), .QN(n696) );
  DFFRX1 \D_cache/cache_reg[1][76]  ( .D(\D_cache/n1187 ), .CK(clk), .RN(n6172), .Q(\D_cache/cache[1][76] ), .QN(n2314) );
  DFFRX1 \D_cache/cache_reg[2][76]  ( .D(\D_cache/n1186 ), .CK(clk), .RN(n6172), .Q(\D_cache/cache[2][76] ), .QN(n1017) );
  DFFRX1 \D_cache/cache_reg[3][76]  ( .D(\D_cache/n1185 ), .CK(clk), .RN(n6172), .Q(\D_cache/cache[3][76] ), .QN(n2643) );
  DFFRX1 \D_cache/cache_reg[4][76]  ( .D(\D_cache/n1184 ), .CK(clk), .RN(n6172), .Q(\D_cache/cache[4][76] ), .QN(n1189) );
  DFFRX1 \D_cache/cache_reg[5][76]  ( .D(\D_cache/n1183 ), .CK(clk), .RN(n6172), .Q(\D_cache/cache[5][76] ), .QN(n2812) );
  DFFRX1 \D_cache/cache_reg[6][76]  ( .D(\D_cache/n1182 ), .CK(clk), .RN(n6172), .Q(\D_cache/cache[6][76] ), .QN(n695) );
  DFFRX1 \D_cache/cache_reg[7][76]  ( .D(\D_cache/n1181 ), .CK(clk), .RN(n6172), .Q(\D_cache/cache[7][76] ), .QN(n2313) );
  DFFRX1 \D_cache/cache_reg[0][77]  ( .D(\D_cache/n1180 ), .CK(clk), .RN(n6172), .Q(\D_cache/cache[0][77] ), .QN(n1030) );
  DFFRX1 \D_cache/cache_reg[1][77]  ( .D(\D_cache/n1179 ), .CK(clk), .RN(n6172), .Q(\D_cache/cache[1][77] ), .QN(n2656) );
  DFFRX1 \D_cache/cache_reg[2][77]  ( .D(\D_cache/n1178 ), .CK(clk), .RN(n6172), .Q(\D_cache/cache[2][77] ), .QN(n1029) );
  DFFRX1 \D_cache/cache_reg[3][77]  ( .D(\D_cache/n1177 ), .CK(clk), .RN(n6172), .Q(\D_cache/cache[3][77] ), .QN(n2655) );
  DFFRX1 \D_cache/cache_reg[4][77]  ( .D(\D_cache/n1176 ), .CK(clk), .RN(n6171), .Q(\D_cache/cache[4][77] ), .QN(n1198) );
  DFFRX1 \D_cache/cache_reg[5][77]  ( .D(\D_cache/n1175 ), .CK(clk), .RN(n6171), .Q(\D_cache/cache[5][77] ), .QN(n2821) );
  DFFRX1 \D_cache/cache_reg[6][77]  ( .D(\D_cache/n1174 ), .CK(clk), .RN(n6171), .Q(\D_cache/cache[6][77] ), .QN(n1028) );
  DFFRX1 \D_cache/cache_reg[7][77]  ( .D(\D_cache/n1173 ), .CK(clk), .RN(n6171), .Q(\D_cache/cache[7][77] ), .QN(n2654) );
  DFFRX1 \D_cache/cache_reg[0][78]  ( .D(\D_cache/n1172 ), .CK(clk), .RN(n6171), .Q(\D_cache/cache[0][78] ), .QN(n557) );
  DFFRX1 \D_cache/cache_reg[1][78]  ( .D(\D_cache/n1171 ), .CK(clk), .RN(n6171), .Q(\D_cache/cache[1][78] ), .QN(n2178) );
  DFFRX1 \D_cache/cache_reg[2][78]  ( .D(\D_cache/n1170 ), .CK(clk), .RN(n6171), .Q(\D_cache/cache[2][78] ), .QN(n1054) );
  DFFRX1 \D_cache/cache_reg[3][78]  ( .D(\D_cache/n1169 ), .CK(clk), .RN(n6171), .Q(\D_cache/cache[3][78] ), .QN(n2681) );
  DFFRX1 \D_cache/cache_reg[4][78]  ( .D(\D_cache/n1168 ), .CK(clk), .RN(n6171), .Q(\D_cache/cache[4][78] ), .QN(n1201) );
  DFFRX1 \D_cache/cache_reg[5][78]  ( .D(\D_cache/n1167 ), .CK(clk), .RN(n6171), .Q(\D_cache/cache[5][78] ), .QN(n2824) );
  DFFRX1 \D_cache/cache_reg[6][78]  ( .D(\D_cache/n1166 ), .CK(clk), .RN(n6171), .Q(\D_cache/cache[6][78] ), .QN(n1053) );
  DFFRX1 \D_cache/cache_reg[7][78]  ( .D(\D_cache/n1165 ), .CK(clk), .RN(n6171), .Q(\D_cache/cache[7][78] ), .QN(n2680) );
  DFFRX1 \D_cache/cache_reg[0][79]  ( .D(\D_cache/n1164 ), .CK(clk), .RN(n6170), .Q(\D_cache/cache[0][79] ), .QN(n1051) );
  DFFRX1 \D_cache/cache_reg[1][79]  ( .D(\D_cache/n1163 ), .CK(clk), .RN(n6170), .Q(\D_cache/cache[1][79] ), .QN(n2678) );
  DFFRX1 \D_cache/cache_reg[2][79]  ( .D(\D_cache/n1162 ), .CK(clk), .RN(n6170), .Q(\D_cache/cache[2][79] ), .QN(n1050) );
  DFFRX1 \D_cache/cache_reg[3][79]  ( .D(\D_cache/n1161 ), .CK(clk), .RN(n6170), .Q(\D_cache/cache[3][79] ), .QN(n2677) );
  DFFRX1 \D_cache/cache_reg[4][79]  ( .D(\D_cache/n1160 ), .CK(clk), .RN(n6170), .Q(\D_cache/cache[4][79] ), .QN(n1210) );
  DFFRX1 \D_cache/cache_reg[5][79]  ( .D(\D_cache/n1159 ), .CK(clk), .RN(n6170), .Q(\D_cache/cache[5][79] ), .QN(n2833) );
  DFFRX1 \D_cache/cache_reg[6][79]  ( .D(\D_cache/n1158 ), .CK(clk), .RN(n6170), .Q(\D_cache/cache[6][79] ), .QN(n594) );
  DFFRX1 \D_cache/cache_reg[7][79]  ( .D(\D_cache/n1157 ), .CK(clk), .RN(n6170), .Q(\D_cache/cache[7][79] ), .QN(n2212) );
  DFFRX1 \D_cache/cache_reg[0][80]  ( .D(\D_cache/n1156 ), .CK(clk), .RN(n6170), .Q(\D_cache/cache[0][80] ), .QN(n640) );
  DFFRX1 \D_cache/cache_reg[1][80]  ( .D(\D_cache/n1155 ), .CK(clk), .RN(n6170), .Q(\D_cache/cache[1][80] ), .QN(n2257) );
  DFFRX1 \D_cache/cache_reg[2][80]  ( .D(\D_cache/n1154 ), .CK(clk), .RN(n6170), .Q(\D_cache/cache[2][80] ), .QN(n639) );
  DFFRX1 \D_cache/cache_reg[3][80]  ( .D(\D_cache/n1153 ), .CK(clk), .RN(n6170), .Q(\D_cache/cache[3][80] ), .QN(n2256) );
  DFFRX1 \D_cache/cache_reg[4][80]  ( .D(\D_cache/n1152 ), .CK(clk), .RN(n6169), .Q(\D_cache/cache[4][80] ), .QN(n625) );
  DFFRX1 \D_cache/cache_reg[5][80]  ( .D(\D_cache/n1151 ), .CK(clk), .RN(n6169), .Q(\D_cache/cache[5][80] ), .QN(n2243) );
  DFFRX1 \D_cache/cache_reg[6][80]  ( .D(\D_cache/n1150 ), .CK(clk), .RN(n6169), .Q(\D_cache/cache[6][80] ), .QN(n638) );
  DFFRX1 \D_cache/cache_reg[7][80]  ( .D(\D_cache/n1149 ), .CK(clk), .RN(n6169), .Q(\D_cache/cache[7][80] ), .QN(n2255) );
  DFFRX1 \D_cache/cache_reg[0][81]  ( .D(\D_cache/n1148 ), .CK(clk), .RN(n6169), .Q(\D_cache/cache[0][81] ), .QN(n2152) );
  DFFRX1 \D_cache/cache_reg[1][81]  ( .D(\D_cache/n1147 ), .CK(clk), .RN(n6169), .Q(\D_cache/cache[1][81] ), .QN(n527) );
  DFFRX1 \D_cache/cache_reg[2][81]  ( .D(\D_cache/n1146 ), .CK(clk), .RN(n6169), .Q(\D_cache/cache[2][81] ), .QN(n2147) );
  DFFRX1 \D_cache/cache_reg[3][81]  ( .D(\D_cache/n1145 ), .CK(clk), .RN(n6169), .Q(\D_cache/cache[3][81] ), .QN(n522) );
  DFFRX1 \D_cache/cache_reg[4][81]  ( .D(\D_cache/n1144 ), .CK(clk), .RN(n6169), .Q(\D_cache/cache[4][81] ), .QN(n2149) );
  DFFRX1 \D_cache/cache_reg[5][81]  ( .D(\D_cache/n1143 ), .CK(clk), .RN(n6169), .Q(\D_cache/cache[5][81] ), .QN(n524) );
  DFFRX1 \D_cache/cache_reg[6][81]  ( .D(\D_cache/n1142 ), .CK(clk), .RN(n6169), .Q(\D_cache/cache[6][81] ), .QN(n574) );
  DFFRX1 \D_cache/cache_reg[7][81]  ( .D(\D_cache/n1141 ), .CK(clk), .RN(n6169), .Q(\D_cache/cache[7][81] ), .QN(n2192) );
  DFFRX1 \D_cache/cache_reg[0][82]  ( .D(\D_cache/n1140 ), .CK(clk), .RN(n6168), .Q(\D_cache/cache[0][82] ), .QN(n1091) );
  DFFRX1 \D_cache/cache_reg[1][82]  ( .D(\D_cache/n1139 ), .CK(clk), .RN(n6168), .Q(\D_cache/cache[1][82] ), .QN(n2714) );
  DFFRX1 \D_cache/cache_reg[2][82]  ( .D(\D_cache/n1138 ), .CK(clk), .RN(n6168), .Q(\D_cache/cache[2][82] ), .QN(n1090) );
  DFFRX1 \D_cache/cache_reg[3][82]  ( .D(\D_cache/n1137 ), .CK(clk), .RN(n6168), .Q(\D_cache/cache[3][82] ), .QN(n2713) );
  DFFRX1 \D_cache/cache_reg[4][82]  ( .D(\D_cache/n1136 ), .CK(clk), .RN(n6168), .Q(\D_cache/cache[4][82] ), .QN(n1165) );
  DFFRX1 \D_cache/cache_reg[5][82]  ( .D(\D_cache/n1135 ), .CK(clk), .RN(n6168), .Q(\D_cache/cache[5][82] ), .QN(n2788) );
  DFFRX1 \D_cache/cache_reg[6][82]  ( .D(\D_cache/n1134 ), .CK(clk), .RN(n6168), .Q(\D_cache/cache[6][82] ), .QN(n1089) );
  DFFRX1 \D_cache/cache_reg[7][82]  ( .D(\D_cache/n1133 ), .CK(clk), .RN(n6168), .Q(\D_cache/cache[7][82] ), .QN(n2712) );
  DFFRX1 \D_cache/cache_reg[0][83]  ( .D(\D_cache/n1132 ), .CK(clk), .RN(n6168), .Q(\D_cache/cache[0][83] ), .QN(n989) );
  DFFRX1 \D_cache/cache_reg[1][83]  ( .D(\D_cache/n1131 ), .CK(clk), .RN(n6168), .Q(\D_cache/cache[1][83] ), .QN(n2614) );
  DFFRX1 \D_cache/cache_reg[2][83]  ( .D(\D_cache/n1130 ), .CK(clk), .RN(n6168), .Q(\D_cache/cache[2][83] ), .QN(n644) );
  DFFRX1 \D_cache/cache_reg[3][83]  ( .D(\D_cache/n1129 ), .CK(clk), .RN(n6168), .Q(\D_cache/cache[3][83] ), .QN(n2261) );
  DFFRX1 \D_cache/cache_reg[4][83]  ( .D(\D_cache/n1128 ), .CK(clk), .RN(n6167), .Q(\D_cache/cache[4][83] ), .QN(n1277) );
  DFFRX1 \D_cache/cache_reg[5][83]  ( .D(\D_cache/n1127 ), .CK(clk), .RN(n6167), .Q(\D_cache/cache[5][83] ), .QN(n2909) );
  DFFRX1 \D_cache/cache_reg[6][83]  ( .D(\D_cache/n1126 ), .CK(clk), .RN(n6167), .Q(\D_cache/cache[6][83] ), .QN(n2144) );
  DFFRX1 \D_cache/cache_reg[7][83]  ( .D(\D_cache/n1125 ), .CK(clk), .RN(n6167), .Q(\D_cache/cache[7][83] ), .QN(n519) );
  DFFRX1 \D_cache/cache_reg[0][84]  ( .D(\D_cache/n1124 ), .CK(clk), .RN(n6167), .Q(\D_cache/cache[0][84] ), .QN(n643) );
  DFFRX1 \D_cache/cache_reg[1][84]  ( .D(\D_cache/n1123 ), .CK(clk), .RN(n6167), .Q(\D_cache/cache[1][84] ), .QN(n2260) );
  DFFRX1 \D_cache/cache_reg[2][84]  ( .D(\D_cache/n1122 ), .CK(clk), .RN(n6167), .Q(\D_cache/cache[2][84] ), .QN(n642) );
  DFFRX1 \D_cache/cache_reg[3][84]  ( .D(\D_cache/n1121 ), .CK(clk), .RN(n6167), .Q(\D_cache/cache[3][84] ), .QN(n2259) );
  DFFRX1 \D_cache/cache_reg[4][84]  ( .D(\D_cache/n1120 ), .CK(clk), .RN(n6167), .Q(\D_cache/cache[4][84] ), .QN(n624) );
  DFFRX1 \D_cache/cache_reg[5][84]  ( .D(\D_cache/n1119 ), .CK(clk), .RN(n6167), .Q(\D_cache/cache[5][84] ), .QN(n2242) );
  DFFRX1 \D_cache/cache_reg[6][84]  ( .D(\D_cache/n1118 ), .CK(clk), .RN(n6167), .Q(\D_cache/cache[6][84] ), .QN(n641) );
  DFFRX1 \D_cache/cache_reg[7][84]  ( .D(\D_cache/n1117 ), .CK(clk), .RN(n6167), .Q(\D_cache/cache[7][84] ), .QN(n2258) );
  DFFRX1 \D_cache/cache_reg[0][85]  ( .D(\D_cache/n1116 ), .CK(clk), .RN(n6166), .Q(\D_cache/cache[0][85] ), .QN(n1114) );
  DFFRX1 \D_cache/cache_reg[1][85]  ( .D(\D_cache/n1115 ), .CK(clk), .RN(n6166), .Q(\D_cache/cache[1][85] ), .QN(n2737) );
  DFFRX1 \D_cache/cache_reg[2][85]  ( .D(\D_cache/n1114 ), .CK(clk), .RN(n6166), .Q(\D_cache/cache[2][85] ), .QN(n2132) );
  DFFRX1 \D_cache/cache_reg[3][85]  ( .D(\D_cache/n1113 ), .CK(clk), .RN(n6166), .Q(\D_cache/cache[3][85] ), .QN(n507) );
  DFFRX1 \D_cache/cache_reg[4][85]  ( .D(\D_cache/n1112 ), .CK(clk), .RN(n6166), .Q(\D_cache/cache[4][85] ), .QN(n974) );
  DFFRX1 \D_cache/cache_reg[5][85]  ( .D(\D_cache/n1111 ), .CK(clk), .RN(n6166), .Q(\D_cache/cache[5][85] ), .QN(n2599) );
  DFFRX1 \D_cache/cache_reg[6][85]  ( .D(\D_cache/n1110 ), .CK(clk), .RN(n6166), .Q(\D_cache/cache[6][85] ), .QN(n604) );
  DFFRX1 \D_cache/cache_reg[7][85]  ( .D(\D_cache/n1109 ), .CK(clk), .RN(n6166), .Q(\D_cache/cache[7][85] ), .QN(n2222) );
  DFFRX1 \D_cache/cache_reg[0][86]  ( .D(\D_cache/n1108 ), .CK(clk), .RN(n6166), .Q(\D_cache/cache[0][86] ), .QN(n646) );
  DFFRX1 \D_cache/cache_reg[1][86]  ( .D(\D_cache/n1107 ), .CK(clk), .RN(n6166), .Q(\D_cache/cache[1][86] ), .QN(n2263) );
  DFFRX1 \D_cache/cache_reg[2][86]  ( .D(\D_cache/n1106 ), .CK(clk), .RN(n6166), .Q(\D_cache/cache[2][86] ), .QN(n609) );
  DFFRX1 \D_cache/cache_reg[3][86]  ( .D(\D_cache/n1105 ), .CK(clk), .RN(n6166), .Q(\D_cache/cache[3][86] ), .QN(n2227) );
  DFFRX1 \D_cache/cache_reg[4][86]  ( .D(\D_cache/n1104 ), .CK(clk), .RN(n6165), .Q(\D_cache/cache[4][86] ), .QN(n988) );
  DFFRX1 \D_cache/cache_reg[5][86]  ( .D(\D_cache/n1103 ), .CK(clk), .RN(n6165), .Q(\D_cache/cache[5][86] ), .QN(n2613) );
  DFFRX1 \D_cache/cache_reg[6][86]  ( .D(\D_cache/n1102 ), .CK(clk), .RN(n6165), .Q(\D_cache/cache[6][86] ), .QN(n645) );
  DFFRX1 \D_cache/cache_reg[7][86]  ( .D(\D_cache/n1101 ), .CK(clk), .RN(n6165), .Q(\D_cache/cache[7][86] ), .QN(n2262) );
  DFFRX1 \D_cache/cache_reg[0][87]  ( .D(\D_cache/n1100 ), .CK(clk), .RN(n6165), .Q(\D_cache/cache[0][87] ), .QN(n632) );
  DFFRX1 \D_cache/cache_reg[1][87]  ( .D(\D_cache/n1099 ), .CK(clk), .RN(n6165), .Q(\D_cache/cache[1][87] ), .QN(n2249) );
  DFFRX1 \D_cache/cache_reg[2][87]  ( .D(\D_cache/n1098 ), .CK(clk), .RN(n6165), .Q(\D_cache/cache[2][87] ), .QN(n631) );
  DFFRX1 \D_cache/cache_reg[3][87]  ( .D(\D_cache/n1097 ), .CK(clk), .RN(n6165), .Q(\D_cache/cache[3][87] ), .QN(n2248) );
  DFFRX1 \D_cache/cache_reg[4][87]  ( .D(\D_cache/n1096 ), .CK(clk), .RN(n6165), .Q(\D_cache/cache[4][87] ), .QN(n987) );
  DFFRX1 \D_cache/cache_reg[5][87]  ( .D(\D_cache/n1095 ), .CK(clk), .RN(n6165), .Q(\D_cache/cache[5][87] ), .QN(n2612) );
  DFFRX1 \D_cache/cache_reg[6][87]  ( .D(\D_cache/n1094 ), .CK(clk), .RN(n6165), .Q(\D_cache/cache[6][87] ), .QN(n630) );
  DFFRX1 \D_cache/cache_reg[7][87]  ( .D(\D_cache/n1093 ), .CK(clk), .RN(n6165), .Q(\D_cache/cache[7][87] ), .QN(n2247) );
  DFFRX1 \D_cache/cache_reg[0][88]  ( .D(\D_cache/n1092 ), .CK(clk), .RN(n6164), .Q(\D_cache/cache[0][88] ), .QN(n1225) );
  DFFRX1 \D_cache/cache_reg[1][88]  ( .D(\D_cache/n1091 ), .CK(clk), .RN(n6164), .Q(\D_cache/cache[1][88] ), .QN(n2848) );
  DFFRX1 \D_cache/cache_reg[2][88]  ( .D(\D_cache/n1090 ), .CK(clk), .RN(n6164), .Q(\D_cache/cache[2][88] ), .QN(n1014) );
  DFFRX1 \D_cache/cache_reg[3][88]  ( .D(\D_cache/n1089 ), .CK(clk), .RN(n6164), .Q(\D_cache/cache[3][88] ), .QN(n2640) );
  DFFRX1 \D_cache/cache_reg[4][88]  ( .D(\D_cache/n1088 ), .CK(clk), .RN(n6164), .Q(\D_cache/cache[4][88] ), .QN(n1285) );
  DFFRX1 \D_cache/cache_reg[5][88]  ( .D(\D_cache/n1087 ), .CK(clk), .RN(n6164), .Q(\D_cache/cache[5][88] ), .QN(n2917) );
  DFFRX1 \D_cache/cache_reg[6][88]  ( .D(\D_cache/n1086 ), .CK(clk), .RN(n6164), .Q(\D_cache/cache[6][88] ), .QN(n1013) );
  DFFRX1 \D_cache/cache_reg[7][88]  ( .D(\D_cache/n1085 ), .CK(clk), .RN(n6164), .Q(\D_cache/cache[7][88] ), .QN(n2639) );
  DFFRX1 \D_cache/cache_reg[0][89]  ( .D(\D_cache/n1084 ), .CK(clk), .RN(n6164), .Q(\D_cache/cache[0][89] ), .QN(n1223) );
  DFFRX1 \D_cache/cache_reg[1][89]  ( .D(\D_cache/n1083 ), .CK(clk), .RN(n6164), .Q(\D_cache/cache[1][89] ), .QN(n2846) );
  DFFRX1 \D_cache/cache_reg[2][89]  ( .D(\D_cache/n1082 ), .CK(clk), .RN(n6164), .Q(\D_cache/cache[2][89] ), .QN(n991) );
  DFFRX1 \D_cache/cache_reg[3][89]  ( .D(\D_cache/n1081 ), .CK(clk), .RN(n6164), .Q(\D_cache/cache[3][89] ), .QN(n2616) );
  DFFRX1 \D_cache/cache_reg[4][89]  ( .D(\D_cache/n1080 ), .CK(clk), .RN(n6163), .Q(\D_cache/cache[4][89] ), .QN(n2886) );
  DFFRX1 \D_cache/cache_reg[5][89]  ( .D(\D_cache/n1079 ), .CK(clk), .RN(n6163), .Q(\D_cache/cache[5][89] ), .QN(n1268) );
  DFFRX1 \D_cache/cache_reg[6][89]  ( .D(\D_cache/n1078 ), .CK(clk), .RN(n6163), .Q(\D_cache/cache[6][89] ), .QN(n649) );
  DFFRX1 \D_cache/cache_reg[7][89]  ( .D(\D_cache/n1077 ), .CK(clk), .RN(n6163), .Q(\D_cache/cache[7][89] ), .QN(n2266) );
  DFFRX1 \D_cache/cache_reg[0][90]  ( .D(\D_cache/n1076 ), .CK(clk), .RN(n6163), .Q(\D_cache/cache[0][90] ), .QN(n615) );
  DFFRX1 \D_cache/cache_reg[1][90]  ( .D(\D_cache/n1075 ), .CK(clk), .RN(n6163), .Q(\D_cache/cache[1][90] ), .QN(n2233) );
  DFFRX1 \D_cache/cache_reg[2][90]  ( .D(\D_cache/n1074 ), .CK(clk), .RN(n6163), .Q(\D_cache/cache[2][90] ), .QN(n1085) );
  DFFRX1 \D_cache/cache_reg[3][90]  ( .D(\D_cache/n1073 ), .CK(clk), .RN(n6163), .Q(\D_cache/cache[3][90] ), .QN(n2708) );
  DFFRX1 \D_cache/cache_reg[4][90]  ( .D(\D_cache/n1072 ), .CK(clk), .RN(n6163), .Q(\D_cache/cache[4][90] ), .QN(n597) );
  DFFRX1 \D_cache/cache_reg[5][90]  ( .D(\D_cache/n1071 ), .CK(clk), .RN(n6163), .Q(\D_cache/cache[5][90] ), .QN(n2215) );
  DFFRX1 \D_cache/cache_reg[6][90]  ( .D(\D_cache/n1070 ), .CK(clk), .RN(n6163), .Q(\D_cache/cache[6][90] ), .QN(n982) );
  DFFRX1 \D_cache/cache_reg[7][90]  ( .D(\D_cache/n1069 ), .CK(clk), .RN(n6163), .Q(\D_cache/cache[7][90] ), .QN(n2607) );
  DFFRX1 \D_cache/cache_reg[0][91]  ( .D(\D_cache/n1068 ), .CK(clk), .RN(n6162), .Q(\D_cache/cache[0][91] ), .QN(n662) );
  DFFRX1 \D_cache/cache_reg[1][91]  ( .D(\D_cache/n1067 ), .CK(clk), .RN(n6162), .Q(\D_cache/cache[1][91] ), .QN(n2279) );
  DFFRX1 \D_cache/cache_reg[2][91]  ( .D(\D_cache/n1066 ), .CK(clk), .RN(n6162), .Q(\D_cache/cache[2][91] ), .QN(n2102) );
  DFFRX1 \D_cache/cache_reg[3][91]  ( .D(\D_cache/n1065 ), .CK(clk), .RN(n6162), .Q(\D_cache/cache[3][91] ), .QN(n476) );
  DFFRX1 \D_cache/cache_reg[4][91]  ( .D(\D_cache/n1064 ), .CK(clk), .RN(n6162), .Q(\D_cache/cache[4][91] ), .QN(n1083) );
  DFFRX1 \D_cache/cache_reg[5][91]  ( .D(\D_cache/n1063 ), .CK(clk), .RN(n6162), .Q(\D_cache/cache[5][91] ), .QN(n2706) );
  DFFRX1 \D_cache/cache_reg[6][91]  ( .D(\D_cache/n1062 ), .CK(clk), .RN(n6162), .Q(\D_cache/cache[6][91] ), .QN(n2075) );
  DFFRX1 \D_cache/cache_reg[7][91]  ( .D(\D_cache/n1061 ), .CK(clk), .RN(n6162), .Q(\D_cache/cache[7][91] ), .QN(n450) );
  DFFRX1 \D_cache/cache_reg[0][92]  ( .D(\D_cache/n1060 ), .CK(clk), .RN(n6162), .Q(\D_cache/cache[0][92] ), .QN(n1099) );
  DFFRX1 \D_cache/cache_reg[1][92]  ( .D(\D_cache/n1059 ), .CK(clk), .RN(n6162), .Q(\D_cache/cache[1][92] ), .QN(n2722) );
  DFFRX1 \D_cache/cache_reg[2][92]  ( .D(\D_cache/n1058 ), .CK(clk), .RN(n6162), .Q(\D_cache/cache[2][92] ), .QN(n1098) );
  DFFRX1 \D_cache/cache_reg[3][92]  ( .D(\D_cache/n1057 ), .CK(clk), .RN(n6162), .Q(\D_cache/cache[3][92] ), .QN(n2721) );
  DFFRX1 \D_cache/cache_reg[4][92]  ( .D(\D_cache/n1056 ), .CK(clk), .RN(n6161), .Q(\D_cache/cache[4][92] ), .QN(n1170) );
  DFFRX1 \D_cache/cache_reg[5][92]  ( .D(\D_cache/n1055 ), .CK(clk), .RN(n6161), .Q(\D_cache/cache[5][92] ), .QN(n2793) );
  DFFRX1 \D_cache/cache_reg[6][92]  ( .D(\D_cache/n1054 ), .CK(clk), .RN(n6161), .Q(\D_cache/cache[6][92] ), .QN(n595) );
  DFFRX1 \D_cache/cache_reg[7][92]  ( .D(\D_cache/n1053 ), .CK(clk), .RN(n6161), .Q(\D_cache/cache[7][92] ), .QN(n2213) );
  DFFRX1 \D_cache/cache_reg[0][93]  ( .D(\D_cache/n1052 ), .CK(clk), .RN(n6161), .Q(\D_cache/cache[0][93] ), .QN(n1148) );
  DFFRX1 \D_cache/cache_reg[1][93]  ( .D(\D_cache/n1051 ), .CK(clk), .RN(n6161), .Q(\D_cache/cache[1][93] ), .QN(n2771) );
  DFFRX1 \D_cache/cache_reg[2][93]  ( .D(\D_cache/n1050 ), .CK(clk), .RN(n6161), .Q(\D_cache/cache[2][93] ), .QN(n1147) );
  DFFRX1 \D_cache/cache_reg[3][93]  ( .D(\D_cache/n1049 ), .CK(clk), .RN(n6161), .Q(\D_cache/cache[3][93] ), .QN(n2770) );
  DFFRX1 \D_cache/cache_reg[4][93]  ( .D(\D_cache/n1048 ), .CK(clk), .RN(n6161), .Q(\D_cache/cache[4][93] ), .QN(n1172) );
  DFFRX1 \D_cache/cache_reg[5][93]  ( .D(\D_cache/n1047 ), .CK(clk), .RN(n6161), .Q(\D_cache/cache[5][93] ), .QN(n2795) );
  DFFRX1 \D_cache/cache_reg[6][93]  ( .D(\D_cache/n1046 ), .CK(clk), .RN(n6161), .Q(\D_cache/cache[6][93] ), .QN(n599) );
  DFFRX1 \D_cache/cache_reg[7][93]  ( .D(\D_cache/n1045 ), .CK(clk), .RN(n6161), .Q(\D_cache/cache[7][93] ), .QN(n2217) );
  DFFRX1 \D_cache/cache_reg[0][94]  ( .D(\D_cache/n1044 ), .CK(clk), .RN(n6160), .Q(\D_cache/cache[0][94] ), .QN(n651) );
  DFFRX1 \D_cache/cache_reg[1][94]  ( .D(\D_cache/n1043 ), .CK(clk), .RN(n6160), .Q(\D_cache/cache[1][94] ), .QN(n2268) );
  DFFRX1 \D_cache/cache_reg[2][94]  ( .D(\D_cache/n1042 ), .CK(clk), .RN(n6160), .Q(\D_cache/cache[2][94] ), .QN(n650) );
  DFFRX1 \D_cache/cache_reg[3][94]  ( .D(\D_cache/n1041 ), .CK(clk), .RN(n6160), .Q(\D_cache/cache[3][94] ), .QN(n2267) );
  DFFRX1 \D_cache/cache_reg[4][94]  ( .D(\D_cache/n1040 ), .CK(clk), .RN(n6160), .Q(\D_cache/cache[4][94] ), .QN(n976) );
  DFFRX1 \D_cache/cache_reg[5][94]  ( .D(\D_cache/n1039 ), .CK(clk), .RN(n6160), .Q(\D_cache/cache[5][94] ), .QN(n2601) );
  DFFRX1 \D_cache/cache_reg[6][94]  ( .D(\D_cache/n1038 ), .CK(clk), .RN(n6160), .Q(\D_cache/cache[6][94] ), .QN(n2110) );
  DFFRX1 \D_cache/cache_reg[7][94]  ( .D(\D_cache/n1037 ), .CK(clk), .RN(n6160), .Q(\D_cache/cache[7][94] ), .QN(n484) );
  DFFRX1 \D_cache/cache_reg[0][95]  ( .D(\D_cache/n1036 ), .CK(clk), .RN(n6160), .Q(\D_cache/cache[0][95] ), .QN(n1164) );
  DFFRX1 \D_cache/cache_reg[1][95]  ( .D(\D_cache/n1035 ), .CK(clk), .RN(n6160), .Q(\D_cache/cache[1][95] ), .QN(n2787) );
  DFFRX1 \D_cache/cache_reg[2][95]  ( .D(\D_cache/n1034 ), .CK(clk), .RN(n6160), .Q(\D_cache/cache[2][95] ), .QN(n2090) );
  DFFRX1 \D_cache/cache_reg[3][95]  ( .D(\D_cache/n1033 ), .CK(clk), .RN(n6160), .Q(\D_cache/cache[3][95] ), .QN(n464) );
  DFFRX1 \D_cache/cache_reg[4][95]  ( .D(\D_cache/n1032 ), .CK(clk), .RN(n6159), .Q(\D_cache/cache[4][95] ), .QN(n2907) );
  DFFRX1 \D_cache/cache_reg[5][95]  ( .D(\D_cache/n1031 ), .CK(clk), .RN(n6159), .Q(\D_cache/cache[5][95] ), .QN(n1240) );
  DFFRX1 \D_cache/cache_reg[6][95]  ( .D(\D_cache/n1030 ), .CK(clk), .RN(n6159), .Q(\D_cache/cache[6][95] ), .QN(n593) );
  DFFRX1 \D_cache/cache_reg[7][95]  ( .D(\D_cache/n1029 ), .CK(clk), .RN(n6159), .Q(\D_cache/cache[7][95] ), .QN(n2211) );
  DFFRX1 \D_cache/cache_reg[0][96]  ( .D(\D_cache/n1028 ), .CK(clk), .RN(n6159), .Q(\D_cache/cache[0][96] ), .QN(n1094) );
  DFFRX1 \D_cache/cache_reg[1][96]  ( .D(\D_cache/n1027 ), .CK(clk), .RN(n6159), .Q(\D_cache/cache[1][96] ), .QN(n2717) );
  DFFRX1 \D_cache/cache_reg[2][96]  ( .D(\D_cache/n1026 ), .CK(clk), .RN(n6159), .Q(\D_cache/cache[2][96] ), .QN(n1093) );
  DFFRX1 \D_cache/cache_reg[3][96]  ( .D(\D_cache/n1025 ), .CK(clk), .RN(n6159), .Q(\D_cache/cache[3][96] ), .QN(n2716) );
  DFFRX1 \D_cache/cache_reg[4][96]  ( .D(\D_cache/n1024 ), .CK(clk), .RN(n6159), .Q(\D_cache/cache[4][96] ), .QN(n1173) );
  DFFRX1 \D_cache/cache_reg[5][96]  ( .D(\D_cache/n1023 ), .CK(clk), .RN(n6159), .Q(\D_cache/cache[5][96] ), .QN(n2796) );
  DFFRX1 \D_cache/cache_reg[6][96]  ( .D(\D_cache/n1022 ), .CK(clk), .RN(n6159), .Q(\D_cache/cache[6][96] ), .QN(n1092) );
  DFFRX1 \D_cache/cache_reg[7][96]  ( .D(\D_cache/n1021 ), .CK(clk), .RN(n6159), .Q(\D_cache/cache[7][96] ), .QN(n2715) );
  DFFRX1 \D_cache/cache_reg[1][97]  ( .D(\D_cache/n1019 ), .CK(clk), .RN(n6158), .Q(\D_cache/cache[1][97] ), .QN(n958) );
  DFFRX1 \D_cache/cache_reg[2][97]  ( .D(\D_cache/n1018 ), .CK(clk), .RN(n6158), .Q(\D_cache/cache[2][97] ), .QN(n2057) );
  DFFRX1 \D_cache/cache_reg[3][97]  ( .D(\D_cache/n1017 ), .CK(clk), .RN(n6158), .Q(\D_cache/cache[3][97] ), .QN(n432) );
  DFFRX1 \D_cache/cache_reg[4][97]  ( .D(\D_cache/n1016 ), .CK(clk), .RN(n6158), .Q(\D_cache/cache[4][97] ), .QN(n563) );
  DFFRX1 \D_cache/cache_reg[5][97]  ( .D(\D_cache/n1015 ), .CK(clk), .RN(n6158), .Q(\D_cache/cache[5][97] ), .QN(n2185) );
  DFFRX1 \D_cache/cache_reg[6][97]  ( .D(\D_cache/n1014 ), .CK(clk), .RN(n6158), .Q(\D_cache/cache[6][97] ), .QN(n2056) );
  DFFRX1 \D_cache/cache_reg[7][97]  ( .D(\D_cache/n1013 ), .CK(clk), .RN(n6158), .Q(\D_cache/cache[7][97] ), .QN(n431) );
  DFFRX1 \D_cache/cache_reg[0][98]  ( .D(\D_cache/n1012 ), .CK(clk), .RN(n6158), .Q(\D_cache/cache[0][98] ), .QN(n684) );
  DFFRX1 \D_cache/cache_reg[1][98]  ( .D(\D_cache/n1011 ), .CK(clk), .RN(n6158), .Q(\D_cache/cache[1][98] ), .QN(n2302) );
  DFFRX1 \D_cache/cache_reg[2][98]  ( .D(\D_cache/n1010 ), .CK(clk), .RN(n6158), .Q(\D_cache/cache[2][98] ), .QN(n2097) );
  DFFRX1 \D_cache/cache_reg[3][98]  ( .D(\D_cache/n1009 ), .CK(clk), .RN(n6158), .Q(\D_cache/cache[3][98] ), .QN(n471) );
  DFFRX1 \D_cache/cache_reg[4][98]  ( .D(\D_cache/n1008 ), .CK(clk), .RN(n6157), .Q(\D_cache/cache[4][98] ), .QN(n1199) );
  DFFRX1 \D_cache/cache_reg[5][98]  ( .D(\D_cache/n1007 ), .CK(clk), .RN(n6157), .Q(\D_cache/cache[5][98] ), .QN(n2822) );
  DFFRX1 \D_cache/cache_reg[6][98]  ( .D(\D_cache/n1006 ), .CK(clk), .RN(n6157), .Q(\D_cache/cache[6][98] ), .QN(n683) );
  DFFRX1 \D_cache/cache_reg[7][98]  ( .D(\D_cache/n1005 ), .CK(clk), .RN(n6157), .Q(\D_cache/cache[7][98] ), .QN(n2301) );
  DFFRX1 \D_cache/cache_reg[0][99]  ( .D(\D_cache/n1004 ), .CK(clk), .RN(n6157), .Q(\D_cache/cache[0][99] ), .QN(n1106) );
  DFFRX1 \D_cache/cache_reg[1][99]  ( .D(\D_cache/n1003 ), .CK(clk), .RN(n6157), .Q(\D_cache/cache[1][99] ), .QN(n2729) );
  DFFRX1 \D_cache/cache_reg[2][99]  ( .D(\D_cache/n1002 ), .CK(clk), .RN(n6157), .Q(\D_cache/cache[2][99] ), .QN(n1105) );
  DFFRX1 \D_cache/cache_reg[3][99]  ( .D(\D_cache/n1001 ), .CK(clk), .RN(n6157), .Q(\D_cache/cache[3][99] ), .QN(n2728) );
  DFFRX1 \D_cache/cache_reg[4][99]  ( .D(\D_cache/n1000 ), .CK(clk), .RN(n6157), .Q(\D_cache/cache[4][99] ), .QN(n975) );
  DFFRX1 \D_cache/cache_reg[5][99]  ( .D(\D_cache/n999 ), .CK(clk), .RN(n6157), 
        .Q(\D_cache/cache[5][99] ), .QN(n2600) );
  DFFRX1 \D_cache/cache_reg[6][99]  ( .D(\D_cache/n998 ), .CK(clk), .RN(n6157), 
        .Q(\D_cache/cache[6][99] ), .QN(n603) );
  DFFRX1 \D_cache/cache_reg[7][99]  ( .D(\D_cache/n997 ), .CK(clk), .RN(n6157), 
        .Q(\D_cache/cache[7][99] ), .QN(n2221) );
  DFFRX1 \D_cache/cache_reg[0][100]  ( .D(\D_cache/n996 ), .CK(clk), .RN(n6156), .Q(\D_cache/cache[0][100] ), .QN(n2906) );
  DFFRX1 \D_cache/cache_reg[1][100]  ( .D(\D_cache/n995 ), .CK(clk), .RN(n6156), .Q(\D_cache/cache[1][100] ), .QN(n1239) );
  DFFRX1 \D_cache/cache_reg[2][100]  ( .D(\D_cache/n994 ), .CK(clk), .RN(n6156), .Q(\D_cache/cache[2][100] ), .QN(n2905) );
  DFFRX1 \D_cache/cache_reg[3][100]  ( .D(\D_cache/n993 ), .CK(clk), .RN(n6156), .Q(\D_cache/cache[3][100] ), .QN(n1238) );
  DFFRX1 \D_cache/cache_reg[4][100]  ( .D(\D_cache/n992 ), .CK(clk), .RN(n6156), .Q(\D_cache/cache[4][100] ), .QN(n1185) );
  DFFRX1 \D_cache/cache_reg[5][100]  ( .D(\D_cache/n991 ), .CK(clk), .RN(n6156), .Q(\D_cache/cache[5][100] ), .QN(n2808) );
  DFFRX1 \D_cache/cache_reg[6][100]  ( .D(\D_cache/n990 ), .CK(clk), .RN(n6156), .Q(\D_cache/cache[6][100] ), .QN(n1146) );
  DFFRX1 \D_cache/cache_reg[7][100]  ( .D(\D_cache/n989 ), .CK(clk), .RN(n6156), .Q(\D_cache/cache[7][100] ), .QN(n2769) );
  DFFRX1 \D_cache/cache_reg[0][101]  ( .D(\D_cache/n988 ), .CK(clk), .RN(n6156), .Q(\D_cache/cache[0][101] ), .QN(n680) );
  DFFRX1 \D_cache/cache_reg[1][101]  ( .D(\D_cache/n987 ), .CK(clk), .RN(n6156), .Q(\D_cache/cache[1][101] ), .QN(n2298) );
  DFFRX1 \D_cache/cache_reg[2][101]  ( .D(\D_cache/n986 ), .CK(clk), .RN(n6156), .Q(\D_cache/cache[2][101] ), .QN(n2083) );
  DFFRX1 \D_cache/cache_reg[3][101]  ( .D(\D_cache/n985 ), .CK(clk), .RN(n6156), .Q(\D_cache/cache[3][101] ), .QN(n457) );
  DFFRX1 \D_cache/cache_reg[4][101]  ( .D(\D_cache/n984 ), .CK(clk), .RN(n6155), .Q(\D_cache/cache[4][101] ), .QN(n1188) );
  DFFRX1 \D_cache/cache_reg[5][101]  ( .D(\D_cache/n983 ), .CK(clk), .RN(n6155), .Q(\D_cache/cache[5][101] ), .QN(n2811) );
  DFFRX1 \D_cache/cache_reg[6][101]  ( .D(\D_cache/n982 ), .CK(clk), .RN(n6155), .Q(\D_cache/cache[6][101] ), .QN(n679) );
  DFFRX1 \D_cache/cache_reg[7][101]  ( .D(\D_cache/n981 ), .CK(clk), .RN(n6155), .Q(\D_cache/cache[7][101] ), .QN(n2297) );
  DFFRX1 \D_cache/cache_reg[0][102]  ( .D(\D_cache/n980 ), .CK(clk), .RN(n6155), .Q(\D_cache/cache[0][102] ), .QN(n690) );
  DFFRX1 \D_cache/cache_reg[1][102]  ( .D(\D_cache/n979 ), .CK(clk), .RN(n6155), .Q(\D_cache/cache[1][102] ), .QN(n2308) );
  DFFRX1 \D_cache/cache_reg[2][102]  ( .D(\D_cache/n978 ), .CK(clk), .RN(n6155), .Q(\D_cache/cache[2][102] ), .QN(n605) );
  DFFRX1 \D_cache/cache_reg[3][102]  ( .D(\D_cache/n977 ), .CK(clk), .RN(n6155), .Q(\D_cache/cache[3][102] ), .QN(n2223) );
  DFFRX1 \D_cache/cache_reg[4][102]  ( .D(\D_cache/n976 ), .CK(clk), .RN(n6155), .Q(\D_cache/cache[4][102] ), .QN(n1202) );
  DFFRX1 \D_cache/cache_reg[5][102]  ( .D(\D_cache/n975 ), .CK(clk), .RN(n6155), .Q(\D_cache/cache[5][102] ), .QN(n2825) );
  DFFRX1 \D_cache/cache_reg[6][102]  ( .D(\D_cache/n974 ), .CK(clk), .RN(n6155), .Q(\D_cache/cache[6][102] ), .QN(n689) );
  DFFRX1 \D_cache/cache_reg[7][102]  ( .D(\D_cache/n973 ), .CK(clk), .RN(n6155), .Q(\D_cache/cache[7][102] ), .QN(n2307) );
  DFFRX1 \D_cache/cache_reg[0][103]  ( .D(\D_cache/n972 ), .CK(clk), .RN(n6154), .Q(\D_cache/cache[0][103] ), .QN(n616) );
  DFFRX1 \D_cache/cache_reg[1][103]  ( .D(\D_cache/n971 ), .CK(clk), .RN(n6154), .Q(\D_cache/cache[1][103] ), .QN(n2234) );
  DFFRX1 \D_cache/cache_reg[2][103]  ( .D(\D_cache/n970 ), .CK(clk), .RN(n6154), .Q(\D_cache/cache[2][103] ), .QN(n1161) );
  DFFRX1 \D_cache/cache_reg[3][103]  ( .D(\D_cache/n969 ), .CK(clk), .RN(n6154), .Q(\D_cache/cache[3][103] ), .QN(n2784) );
  DFFRX1 \D_cache/cache_reg[4][103]  ( .D(\D_cache/n968 ), .CK(clk), .RN(n6154), .Q(\D_cache/cache[4][103] ), .QN(n1200) );
  DFFRX1 \D_cache/cache_reg[5][103]  ( .D(\D_cache/n967 ), .CK(clk), .RN(n6154), .Q(\D_cache/cache[5][103] ), .QN(n2823) );
  DFFRX1 \D_cache/cache_reg[6][103]  ( .D(\D_cache/n966 ), .CK(clk), .RN(n6154), .Q(\D_cache/cache[6][103] ), .QN(n979) );
  DFFRX1 \D_cache/cache_reg[7][103]  ( .D(\D_cache/n965 ), .CK(clk), .RN(n6154), .Q(\D_cache/cache[7][103] ), .QN(n2604) );
  DFFRX1 \D_cache/cache_reg[0][104]  ( .D(\D_cache/n964 ), .CK(clk), .RN(n6154), .Q(\D_cache/cache[0][104] ), .QN(n1119) );
  DFFRX1 \D_cache/cache_reg[1][104]  ( .D(\D_cache/n963 ), .CK(clk), .RN(n6154), .Q(\D_cache/cache[1][104] ), .QN(n2742) );
  DFFRX1 \D_cache/cache_reg[2][104]  ( .D(\D_cache/n962 ), .CK(clk), .RN(n6154), .Q(\D_cache/cache[2][104] ), .QN(n1118) );
  DFFRX1 \D_cache/cache_reg[3][104]  ( .D(\D_cache/n961 ), .CK(clk), .RN(n6154), .Q(\D_cache/cache[3][104] ), .QN(n2741) );
  DFFRX1 \D_cache/cache_reg[4][104]  ( .D(\D_cache/n960 ), .CK(clk), .RN(n6153), .Q(\D_cache/cache[4][104] ), .QN(n1236) );
  DFFRX1 \D_cache/cache_reg[5][104]  ( .D(\D_cache/n959 ), .CK(clk), .RN(n6153), .Q(\D_cache/cache[5][104] ), .QN(n2858) );
  DFFRX1 \D_cache/cache_reg[6][104]  ( .D(\D_cache/n958 ), .CK(clk), .RN(n6153), .Q(\D_cache/cache[6][104] ), .QN(n1117) );
  DFFRX1 \D_cache/cache_reg[7][104]  ( .D(\D_cache/n957 ), .CK(clk), .RN(n6153), .Q(\D_cache/cache[7][104] ), .QN(n2740) );
  DFFRX1 \D_cache/cache_reg[0][105]  ( .D(\D_cache/n956 ), .CK(clk), .RN(n6153), .Q(\D_cache/cache[0][105] ), .QN(n1142) );
  DFFRX1 \D_cache/cache_reg[1][105]  ( .D(\D_cache/n955 ), .CK(clk), .RN(n6153), .Q(\D_cache/cache[1][105] ), .QN(n2765) );
  DFFRX1 \D_cache/cache_reg[2][105]  ( .D(\D_cache/n954 ), .CK(clk), .RN(n6153), .Q(\D_cache/cache[2][105] ), .QN(n1141) );
  DFFRX1 \D_cache/cache_reg[3][105]  ( .D(\D_cache/n953 ), .CK(clk), .RN(n6153), .Q(\D_cache/cache[3][105] ), .QN(n2764) );
  DFFRX1 \D_cache/cache_reg[4][105]  ( .D(\D_cache/n952 ), .CK(clk), .RN(n6153), .Q(\D_cache/cache[4][105] ), .QN(n585) );
  DFFRX1 \D_cache/cache_reg[5][105]  ( .D(\D_cache/n951 ), .CK(clk), .RN(n6153), .Q(\D_cache/cache[5][105] ), .QN(n2203) );
  DFFRX1 \D_cache/cache_reg[6][105]  ( .D(\D_cache/n950 ), .CK(clk), .RN(n6153), .Q(\D_cache/cache[6][105] ), .QN(n1140) );
  DFFRX1 \D_cache/cache_reg[7][105]  ( .D(\D_cache/n949 ), .CK(clk), .RN(n6153), .Q(\D_cache/cache[7][105] ), .QN(n2763) );
  DFFRX1 \D_cache/cache_reg[0][106]  ( .D(\D_cache/n948 ), .CK(clk), .RN(n6152), .Q(\D_cache/cache[0][106] ), .QN(n1136) );
  DFFRX1 \D_cache/cache_reg[1][106]  ( .D(\D_cache/n947 ), .CK(clk), .RN(n6152), .Q(\D_cache/cache[1][106] ), .QN(n2759) );
  DFFRX1 \D_cache/cache_reg[2][106]  ( .D(\D_cache/n946 ), .CK(clk), .RN(n6152), .Q(\D_cache/cache[2][106] ), .QN(n1135) );
  DFFRX1 \D_cache/cache_reg[3][106]  ( .D(\D_cache/n945 ), .CK(clk), .RN(n6152), .Q(\D_cache/cache[3][106] ), .QN(n2758) );
  DFFRX1 \D_cache/cache_reg[4][106]  ( .D(\D_cache/n944 ), .CK(clk), .RN(n6152), .Q(\D_cache/cache[4][106] ), .QN(n1175) );
  DFFRX1 \D_cache/cache_reg[5][106]  ( .D(\D_cache/n943 ), .CK(clk), .RN(n6152), .Q(\D_cache/cache[5][106] ), .QN(n2798) );
  DFFRX1 \D_cache/cache_reg[6][106]  ( .D(\D_cache/n942 ), .CK(clk), .RN(n6152), .Q(\D_cache/cache[6][106] ), .QN(n1134) );
  DFFRX1 \D_cache/cache_reg[7][106]  ( .D(\D_cache/n941 ), .CK(clk), .RN(n6152), .Q(\D_cache/cache[7][106] ), .QN(n2757) );
  DFFRX1 \D_cache/cache_reg[0][107]  ( .D(\D_cache/n940 ), .CK(clk), .RN(n6152), .Q(\D_cache/cache[0][107] ), .QN(n1097) );
  DFFRX1 \D_cache/cache_reg[1][107]  ( .D(\D_cache/n939 ), .CK(clk), .RN(n6152), .Q(\D_cache/cache[1][107] ), .QN(n2720) );
  DFFRX1 \D_cache/cache_reg[2][107]  ( .D(\D_cache/n938 ), .CK(clk), .RN(n6152), .Q(\D_cache/cache[2][107] ), .QN(n1096) );
  DFFRX1 \D_cache/cache_reg[3][107]  ( .D(\D_cache/n937 ), .CK(clk), .RN(n6152), .Q(\D_cache/cache[3][107] ), .QN(n2719) );
  DFFRX1 \D_cache/cache_reg[4][107]  ( .D(\D_cache/n936 ), .CK(clk), .RN(n6151), .Q(\D_cache/cache[4][107] ), .QN(n1169) );
  DFFRX1 \D_cache/cache_reg[5][107]  ( .D(\D_cache/n935 ), .CK(clk), .RN(n6151), .Q(\D_cache/cache[5][107] ), .QN(n2792) );
  DFFRX1 \D_cache/cache_reg[6][107]  ( .D(\D_cache/n934 ), .CK(clk), .RN(n6151), .Q(\D_cache/cache[6][107] ), .QN(n1095) );
  DFFRX1 \D_cache/cache_reg[7][107]  ( .D(\D_cache/n933 ), .CK(clk), .RN(n6151), .Q(\D_cache/cache[7][107] ), .QN(n2718) );
  DFFRX1 \D_cache/cache_reg[0][108]  ( .D(\D_cache/n932 ), .CK(clk), .RN(n6151), .Q(\D_cache/cache[0][108] ), .QN(n1124) );
  DFFRX1 \D_cache/cache_reg[1][108]  ( .D(\D_cache/n931 ), .CK(clk), .RN(n6151), .Q(\D_cache/cache[1][108] ), .QN(n2747) );
  DFFRX1 \D_cache/cache_reg[2][108]  ( .D(\D_cache/n930 ), .CK(clk), .RN(n6151), .Q(\D_cache/cache[2][108] ), .QN(n1123) );
  DFFRX1 \D_cache/cache_reg[3][108]  ( .D(\D_cache/n929 ), .CK(clk), .RN(n6151), .Q(\D_cache/cache[3][108] ), .QN(n2746) );
  DFFRX1 \D_cache/cache_reg[4][108]  ( .D(\D_cache/n928 ), .CK(clk), .RN(n6151), .Q(\D_cache/cache[4][108] ), .QN(n1174) );
  DFFRX1 \D_cache/cache_reg[5][108]  ( .D(\D_cache/n927 ), .CK(clk), .RN(n6151), .Q(\D_cache/cache[5][108] ), .QN(n2797) );
  DFFRX1 \D_cache/cache_reg[6][108]  ( .D(\D_cache/n926 ), .CK(clk), .RN(n6151), .Q(\D_cache/cache[6][108] ), .QN(n2071) );
  DFFRX1 \D_cache/cache_reg[7][108]  ( .D(\D_cache/n925 ), .CK(clk), .RN(n6151), .Q(\D_cache/cache[7][108] ), .QN(n446) );
  DFFRX1 \D_cache/cache_reg[0][109]  ( .D(\D_cache/n924 ), .CK(clk), .RN(n6150), .Q(\D_cache/cache[0][109] ), .QN(n1152) );
  DFFRX1 \D_cache/cache_reg[1][109]  ( .D(\D_cache/n923 ), .CK(clk), .RN(n6150), .Q(\D_cache/cache[1][109] ), .QN(n2775) );
  DFFRX1 \D_cache/cache_reg[2][109]  ( .D(\D_cache/n922 ), .CK(clk), .RN(n6150), .Q(\D_cache/cache[2][109] ), .QN(n1151) );
  DFFRX1 \D_cache/cache_reg[3][109]  ( .D(\D_cache/n921 ), .CK(clk), .RN(n6150), .Q(\D_cache/cache[3][109] ), .QN(n2774) );
  DFFRX1 \D_cache/cache_reg[4][109]  ( .D(\D_cache/n920 ), .CK(clk), .RN(n6150), .Q(\D_cache/cache[4][109] ), .QN(n1179) );
  DFFRX1 \D_cache/cache_reg[5][109]  ( .D(\D_cache/n919 ), .CK(clk), .RN(n6150), .Q(\D_cache/cache[5][109] ), .QN(n2802) );
  DFFRX1 \D_cache/cache_reg[6][109]  ( .D(\D_cache/n918 ), .CK(clk), .RN(n6150), .Q(\D_cache/cache[6][109] ), .QN(n2116) );
  DFFRX1 \D_cache/cache_reg[7][109]  ( .D(\D_cache/n917 ), .CK(clk), .RN(n6150), .Q(\D_cache/cache[7][109] ), .QN(n490) );
  DFFRX1 \D_cache/cache_reg[0][110]  ( .D(\D_cache/n916 ), .CK(clk), .RN(n6150), .Q(\D_cache/cache[0][110] ), .QN(n1066) );
  DFFRX1 \D_cache/cache_reg[1][110]  ( .D(\D_cache/n915 ), .CK(clk), .RN(n6150), .Q(\D_cache/cache[1][110] ), .QN(n2694) );
  DFFRX1 \D_cache/cache_reg[2][110]  ( .D(\D_cache/n914 ), .CK(clk), .RN(n6150), .Q(\D_cache/cache[2][110] ), .QN(n580) );
  DFFRX1 \D_cache/cache_reg[3][110]  ( .D(\D_cache/n913 ), .CK(clk), .RN(n6150), .Q(\D_cache/cache[3][110] ), .QN(n2198) );
  DFFRX1 \D_cache/cache_reg[4][110]  ( .D(\D_cache/n912 ), .CK(clk), .RN(n6149), .Q(\D_cache/cache[4][110] ), .QN(n581) );
  DFFRX1 \D_cache/cache_reg[5][110]  ( .D(\D_cache/n911 ), .CK(clk), .RN(n6149), .Q(\D_cache/cache[5][110] ), .QN(n2199) );
  DFFRX1 \D_cache/cache_reg[6][110]  ( .D(\D_cache/n910 ), .CK(clk), .RN(n6149), .Q(\D_cache/cache[6][110] ), .QN(n1065) );
  DFFRX1 \D_cache/cache_reg[7][110]  ( .D(\D_cache/n909 ), .CK(clk), .RN(n6149), .Q(\D_cache/cache[7][110] ), .QN(n2693) );
  DFFRX1 \D_cache/cache_reg[0][111]  ( .D(\D_cache/n908 ), .CK(clk), .RN(n6149), .Q(\D_cache/cache[0][111] ), .QN(n1071) );
  DFFRX1 \D_cache/cache_reg[1][111]  ( .D(\D_cache/n907 ), .CK(clk), .RN(n6149), .Q(\D_cache/cache[1][111] ), .QN(n2699) );
  DFFRX1 \D_cache/cache_reg[2][111]  ( .D(\D_cache/n906 ), .CK(clk), .RN(n6149), .Q(\D_cache/cache[2][111] ), .QN(n1070) );
  DFFRX1 \D_cache/cache_reg[3][111]  ( .D(\D_cache/n905 ), .CK(clk), .RN(n6149), .Q(\D_cache/cache[3][111] ), .QN(n2698) );
  DFFRX1 \D_cache/cache_reg[4][111]  ( .D(\D_cache/n904 ), .CK(clk), .RN(n6149), .Q(\D_cache/cache[4][111] ), .QN(n1217) );
  DFFRX1 \D_cache/cache_reg[5][111]  ( .D(\D_cache/n903 ), .CK(clk), .RN(n6149), .Q(\D_cache/cache[5][111] ), .QN(n2840) );
  DFFRX1 \D_cache/cache_reg[6][111]  ( .D(\D_cache/n902 ), .CK(clk), .RN(n6149), .Q(\D_cache/cache[6][111] ), .QN(n1069) );
  DFFRX1 \D_cache/cache_reg[7][111]  ( .D(\D_cache/n901 ), .CK(clk), .RN(n6149), .Q(\D_cache/cache[7][111] ), .QN(n2697) );
  DFFRX1 \D_cache/cache_reg[0][112]  ( .D(\D_cache/n900 ), .CK(clk), .RN(n6148), .Q(\D_cache/cache[0][112] ), .QN(n1125) );
  DFFRX1 \D_cache/cache_reg[1][112]  ( .D(\D_cache/n899 ), .CK(clk), .RN(n6148), .Q(\D_cache/cache[1][112] ), .QN(n2748) );
  DFFRX1 \D_cache/cache_reg[2][112]  ( .D(\D_cache/n898 ), .CK(clk), .RN(n6148), .Q(\D_cache/cache[2][112] ), .QN(n2125) );
  DFFRX1 \D_cache/cache_reg[3][112]  ( .D(\D_cache/n897 ), .CK(clk), .RN(n6148), .Q(\D_cache/cache[3][112] ), .QN(n500) );
  DFFRX1 \D_cache/cache_reg[4][112]  ( .D(\D_cache/n896 ), .CK(clk), .RN(n6148), .Q(\D_cache/cache[4][112] ), .QN(n607) );
  DFFRX1 \D_cache/cache_reg[5][112]  ( .D(\D_cache/n895 ), .CK(clk), .RN(n6148), .Q(\D_cache/cache[5][112] ), .QN(n2225) );
  DFFRX1 \D_cache/cache_reg[6][112]  ( .D(\D_cache/n894 ), .CK(clk), .RN(n6148), .Q(\D_cache/cache[6][112] ), .QN(n977) );
  DFFRX1 \D_cache/cache_reg[7][112]  ( .D(\D_cache/n893 ), .CK(clk), .RN(n6148), .Q(\D_cache/cache[7][112] ), .QN(n2602) );
  DFFRX1 \D_cache/cache_reg[0][113]  ( .D(\D_cache/n892 ), .CK(clk), .RN(n6148), .Q(\D_cache/cache[0][113] ), .QN(n1163) );
  DFFRX1 \D_cache/cache_reg[1][113]  ( .D(\D_cache/n891 ), .CK(clk), .RN(n6148), .Q(\D_cache/cache[1][113] ), .QN(n2786) );
  DFFRX1 \D_cache/cache_reg[2][113]  ( .D(\D_cache/n890 ), .CK(clk), .RN(n6148), .Q(\D_cache/cache[2][113] ), .QN(n1162) );
  DFFRX1 \D_cache/cache_reg[3][113]  ( .D(\D_cache/n889 ), .CK(clk), .RN(n6148), .Q(\D_cache/cache[3][113] ), .QN(n2785) );
  DFFRX1 \D_cache/cache_reg[4][113]  ( .D(\D_cache/n888 ), .CK(clk), .RN(n6147), .Q(\D_cache/cache[4][113] ), .QN(n1196) );
  DFFRX1 \D_cache/cache_reg[5][113]  ( .D(\D_cache/n887 ), .CK(clk), .RN(n6147), .Q(\D_cache/cache[5][113] ), .QN(n2819) );
  DFFRX1 \D_cache/cache_reg[6][113]  ( .D(\D_cache/n886 ), .CK(clk), .RN(n6147), .Q(\D_cache/cache[6][113] ), .QN(n2128) );
  DFFRX1 \D_cache/cache_reg[7][113]  ( .D(\D_cache/n885 ), .CK(clk), .RN(n6147), .Q(\D_cache/cache[7][113] ), .QN(n503) );
  DFFRX1 \D_cache/cache_reg[0][114]  ( .D(\D_cache/n884 ), .CK(clk), .RN(n6147), .Q(\D_cache/cache[0][114] ), .QN(n1113) );
  DFFRX1 \D_cache/cache_reg[1][114]  ( .D(\D_cache/n883 ), .CK(clk), .RN(n6147), .Q(\D_cache/cache[1][114] ), .QN(n2736) );
  DFFRX1 \D_cache/cache_reg[2][114]  ( .D(\D_cache/n882 ), .CK(clk), .RN(n6147), .Q(\D_cache/cache[2][114] ), .QN(n1112) );
  DFFRX1 \D_cache/cache_reg[3][114]  ( .D(\D_cache/n881 ), .CK(clk), .RN(n6147), .Q(\D_cache/cache[3][114] ), .QN(n2735) );
  DFFRX1 \D_cache/cache_reg[4][114]  ( .D(\D_cache/n880 ), .CK(clk), .RN(n6147), .Q(\D_cache/cache[4][114] ), .QN(n973) );
  DFFRX1 \D_cache/cache_reg[5][114]  ( .D(\D_cache/n879 ), .CK(clk), .RN(n6147), .Q(\D_cache/cache[5][114] ), .QN(n2598) );
  DFFRX1 \D_cache/cache_reg[6][114]  ( .D(\D_cache/n878 ), .CK(clk), .RN(n6147), .Q(\D_cache/cache[6][114] ), .QN(n1111) );
  DFFRX1 \D_cache/cache_reg[7][114]  ( .D(\D_cache/n877 ), .CK(clk), .RN(n6147), .Q(\D_cache/cache[7][114] ), .QN(n2734) );
  DFFRX1 \D_cache/cache_reg[0][115]  ( .D(\D_cache/n876 ), .CK(clk), .RN(n6146), .Q(\D_cache/cache[0][115] ), .QN(n955) );
  DFFRX1 \D_cache/cache_reg[1][115]  ( .D(\D_cache/n875 ), .CK(clk), .RN(n6146), .Q(\D_cache/cache[1][115] ), .QN(n2579) );
  DFFRX1 \D_cache/cache_reg[2][115]  ( .D(\D_cache/n874 ), .CK(clk), .RN(n6146), .Q(\D_cache/cache[2][115] ), .QN(n954) );
  DFFRX1 \D_cache/cache_reg[3][115]  ( .D(\D_cache/n873 ), .CK(clk), .RN(n6146), .Q(\D_cache/cache[3][115] ), .QN(n2578) );
  DFFRX1 \D_cache/cache_reg[4][115]  ( .D(\D_cache/n872 ), .CK(clk), .RN(n6146), .Q(\D_cache/cache[4][115] ), .QN(n956) );
  DFFRX1 \D_cache/cache_reg[5][115]  ( .D(\D_cache/n871 ), .CK(clk), .RN(n6146), .Q(\D_cache/cache[5][115] ), .QN(n2580) );
  DFFRX1 \D_cache/cache_reg[6][115]  ( .D(\D_cache/n870 ), .CK(clk), .RN(n6146), .Q(\D_cache/cache[6][115] ), .QN(n2055) );
  DFFRX1 \D_cache/cache_reg[7][115]  ( .D(\D_cache/n869 ), .CK(clk), .RN(n6146), .Q(\D_cache/cache[7][115] ), .QN(n430) );
  DFFRX1 \D_cache/cache_reg[0][116]  ( .D(\D_cache/n868 ), .CK(clk), .RN(n6146), .Q(\D_cache/cache[0][116] ), .QN(n1139) );
  DFFRX1 \D_cache/cache_reg[1][116]  ( .D(\D_cache/n867 ), .CK(clk), .RN(n6146), .Q(\D_cache/cache[1][116] ), .QN(n2762) );
  DFFRX1 \D_cache/cache_reg[2][116]  ( .D(\D_cache/n866 ), .CK(clk), .RN(n6146), .Q(\D_cache/cache[2][116] ), .QN(n980) );
  DFFRX1 \D_cache/cache_reg[3][116]  ( .D(\D_cache/n865 ), .CK(clk), .RN(n6146), .Q(\D_cache/cache[3][116] ), .QN(n2605) );
  DFFRX1 \D_cache/cache_reg[4][116]  ( .D(\D_cache/n864 ), .CK(clk), .RN(n6145), .Q(\D_cache/cache[4][116] ), .QN(n1178) );
  DFFRX1 \D_cache/cache_reg[5][116]  ( .D(\D_cache/n863 ), .CK(clk), .RN(n6145), .Q(\D_cache/cache[5][116] ), .QN(n2801) );
  DFFRX1 \D_cache/cache_reg[6][116]  ( .D(\D_cache/n862 ), .CK(clk), .RN(n6145), .Q(\D_cache/cache[6][116] ), .QN(n2145) );
  DFFRX1 \D_cache/cache_reg[7][116]  ( .D(\D_cache/n861 ), .CK(clk), .RN(n6145), .Q(\D_cache/cache[7][116] ), .QN(n520) );
  DFFRX1 \D_cache/cache_reg[0][117]  ( .D(\D_cache/n860 ), .CK(clk), .RN(n6145), .Q(\D_cache/cache[0][117] ), .QN(n1138) );
  DFFRX1 \D_cache/cache_reg[1][117]  ( .D(\D_cache/n859 ), .CK(clk), .RN(n6145), .Q(\D_cache/cache[1][117] ), .QN(n2761) );
  DFFRX1 \D_cache/cache_reg[2][117]  ( .D(\D_cache/n858 ), .CK(clk), .RN(n6145), .Q(\D_cache/cache[2][117] ), .QN(n2134) );
  DFFRX1 \D_cache/cache_reg[3][117]  ( .D(\D_cache/n857 ), .CK(clk), .RN(n6145), .Q(\D_cache/cache[3][117] ), .QN(n509) );
  DFFRX1 \D_cache/cache_reg[4][117]  ( .D(\D_cache/n856 ), .CK(clk), .RN(n6145), .Q(\D_cache/cache[4][117] ), .QN(n1180) );
  DFFRX1 \D_cache/cache_reg[5][117]  ( .D(\D_cache/n855 ), .CK(clk), .RN(n6145), .Q(\D_cache/cache[5][117] ), .QN(n2803) );
  DFFRX1 \D_cache/cache_reg[6][117]  ( .D(\D_cache/n854 ), .CK(clk), .RN(n6145), .Q(\D_cache/cache[6][117] ), .QN(n1137) );
  DFFRX1 \D_cache/cache_reg[7][117]  ( .D(\D_cache/n853 ), .CK(clk), .RN(n6145), .Q(\D_cache/cache[7][117] ), .QN(n2760) );
  DFFRX1 \D_cache/cache_reg[0][118]  ( .D(\D_cache/n852 ), .CK(clk), .RN(n6144), .Q(\D_cache/cache[0][118] ), .QN(n1005) );
  DFFRX1 \D_cache/cache_reg[1][118]  ( .D(\D_cache/n851 ), .CK(clk), .RN(n6144), .Q(\D_cache/cache[1][118] ), .QN(n2630) );
  DFFRX1 \D_cache/cache_reg[2][118]  ( .D(\D_cache/n850 ), .CK(clk), .RN(n6144), .Q(\D_cache/cache[2][118] ), .QN(n1004) );
  DFFRX1 \D_cache/cache_reg[3][118]  ( .D(\D_cache/n849 ), .CK(clk), .RN(n6144), .Q(\D_cache/cache[3][118] ), .QN(n2629) );
  DFFRX1 \D_cache/cache_reg[4][118]  ( .D(\D_cache/n848 ), .CK(clk), .RN(n6144), .Q(\D_cache/cache[4][118] ), .QN(n1088) );
  DFFRX1 \D_cache/cache_reg[5][118]  ( .D(\D_cache/n847 ), .CK(clk), .RN(n6144), .Q(\D_cache/cache[5][118] ), .QN(n2711) );
  DFFRX1 \D_cache/cache_reg[6][118]  ( .D(\D_cache/n846 ), .CK(clk), .RN(n6144), .Q(\D_cache/cache[6][118] ), .QN(n1003) );
  DFFRX1 \D_cache/cache_reg[7][118]  ( .D(\D_cache/n845 ), .CK(clk), .RN(n6144), .Q(\D_cache/cache[7][118] ), .QN(n2628) );
  DFFRX1 \D_cache/cache_reg[0][119]  ( .D(\D_cache/n844 ), .CK(clk), .RN(n6144), .Q(\D_cache/cache[0][119] ), .QN(n674) );
  DFFRX1 \D_cache/cache_reg[1][119]  ( .D(\D_cache/n843 ), .CK(clk), .RN(n6144), .Q(\D_cache/cache[1][119] ), .QN(n2292) );
  DFFRX1 \D_cache/cache_reg[2][119]  ( .D(\D_cache/n842 ), .CK(clk), .RN(n6144), .Q(\D_cache/cache[2][119] ), .QN(n997) );
  DFFRX1 \D_cache/cache_reg[3][119]  ( .D(\D_cache/n841 ), .CK(clk), .RN(n6144), .Q(\D_cache/cache[3][119] ), .QN(n2622) );
  DFFRX1 \D_cache/cache_reg[4][119]  ( .D(\D_cache/n840 ), .CK(clk), .RN(n6143), .Q(\D_cache/cache[4][119] ), .QN(n1184) );
  DFFRX1 \D_cache/cache_reg[5][119]  ( .D(\D_cache/n839 ), .CK(clk), .RN(n6143), .Q(\D_cache/cache[5][119] ), .QN(n2807) );
  DFFRX1 \D_cache/cache_reg[6][119]  ( .D(\D_cache/n838 ), .CK(clk), .RN(n6143), .Q(\D_cache/cache[6][119] ), .QN(n673) );
  DFFRX1 \D_cache/cache_reg[7][119]  ( .D(\D_cache/n837 ), .CK(clk), .RN(n6143), .Q(\D_cache/cache[7][119] ), .QN(n2291) );
  DFFRX1 \D_cache/cache_reg[0][120]  ( .D(\D_cache/n836 ), .CK(clk), .RN(n6143), .Q(\D_cache/cache[0][120] ), .QN(n1234) );
  DFFRX1 \D_cache/cache_reg[1][120]  ( .D(\D_cache/n835 ), .CK(clk), .RN(n6143), .Q(\D_cache/cache[1][120] ), .QN(n2856) );
  DFFRX1 \D_cache/cache_reg[2][120]  ( .D(\D_cache/n834 ), .CK(clk), .RN(n6143), .Q(\D_cache/cache[2][120] ), .QN(n1233) );
  DFFRX1 \D_cache/cache_reg[3][120]  ( .D(\D_cache/n833 ), .CK(clk), .RN(n6143), .Q(\D_cache/cache[3][120] ), .QN(n2855) );
  DFFRX1 \D_cache/cache_reg[4][120]  ( .D(\D_cache/n832 ), .CK(clk), .RN(n6143), .Q(\D_cache/cache[4][120] ), .QN(n1283) );
  DFFRX1 \D_cache/cache_reg[5][120]  ( .D(\D_cache/n831 ), .CK(clk), .RN(n6143), .Q(\D_cache/cache[5][120] ), .QN(n2915) );
  DFFRX1 \D_cache/cache_reg[6][120]  ( .D(\D_cache/n830 ), .CK(clk), .RN(n6143), .Q(\D_cache/cache[6][120] ), .QN(n962) );
  DFFRX1 \D_cache/cache_reg[7][120]  ( .D(\D_cache/n829 ), .CK(clk), .RN(n6143), .Q(\D_cache/cache[7][120] ), .QN(n2587) );
  DFFRX1 \D_cache/cache_reg[0][121]  ( .D(\D_cache/n828 ), .CK(clk), .RN(n6142), .Q(\D_cache/cache[0][121] ), .QN(n1232) );
  DFFRX1 \D_cache/cache_reg[1][121]  ( .D(\D_cache/n827 ), .CK(clk), .RN(n6142), .Q(\D_cache/cache[1][121] ), .QN(n2854) );
  DFFRX1 \D_cache/cache_reg[2][121]  ( .D(\D_cache/n826 ), .CK(clk), .RN(n6142), .Q(\D_cache/cache[2][121] ), .QN(n1074) );
  DFFRX1 \D_cache/cache_reg[3][121]  ( .D(\D_cache/n825 ), .CK(clk), .RN(n6142), .Q(\D_cache/cache[3][121] ), .QN(n2702) );
  DFFRX1 \D_cache/cache_reg[4][121]  ( .D(\D_cache/n824 ), .CK(clk), .RN(n6142), .Q(\D_cache/cache[4][121] ), .QN(n1282) );
  DFFRX1 \D_cache/cache_reg[5][121]  ( .D(\D_cache/n823 ), .CK(clk), .RN(n6142), .Q(\D_cache/cache[5][121] ), .QN(n2914) );
  DFFRX1 \D_cache/cache_reg[6][121]  ( .D(\D_cache/n822 ), .CK(clk), .RN(n6142), .Q(\D_cache/cache[6][121] ), .QN(n1073) );
  DFFRX1 \D_cache/cache_reg[7][121]  ( .D(\D_cache/n821 ), .CK(clk), .RN(n6142), .Q(\D_cache/cache[7][121] ), .QN(n2701) );
  DFFRX1 \D_cache/cache_reg[0][122]  ( .D(\D_cache/n820 ), .CK(clk), .RN(n6142), .Q(\D_cache/cache[0][122] ), .QN(n1080) );
  DFFRX1 \D_cache/cache_reg[1][122]  ( .D(\D_cache/n819 ), .CK(clk), .RN(n6142), .Q(\D_cache/cache[1][122] ), .QN(n2703) );
  DFFRX1 \D_cache/cache_reg[2][122]  ( .D(\D_cache/n818 ), .CK(clk), .RN(n6142), .Q(\D_cache/cache[2][122] ), .QN(n1037) );
  DFFRX1 \D_cache/cache_reg[3][122]  ( .D(\D_cache/n817 ), .CK(clk), .RN(n6142), .Q(\D_cache/cache[3][122] ), .QN(n2663) );
  DFFRX1 \D_cache/cache_reg[4][122]  ( .D(\D_cache/n816 ), .CK(clk), .RN(n6141), .Q(\D_cache/cache[4][122] ), .QN(n1203) );
  DFFRX1 \D_cache/cache_reg[5][122]  ( .D(\D_cache/n815 ), .CK(clk), .RN(n6141), .Q(\D_cache/cache[5][122] ), .QN(n2826) );
  DFFRX1 \D_cache/cache_reg[6][122]  ( .D(\D_cache/n814 ), .CK(clk), .RN(n6141), .Q(\D_cache/cache[6][122] ), .QN(n1036) );
  DFFRX1 \D_cache/cache_reg[7][122]  ( .D(\D_cache/n813 ), .CK(clk), .RN(n6141), .Q(\D_cache/cache[7][122] ), .QN(n2662) );
  DFFRX1 \D_cache/cache_reg[0][123]  ( .D(\D_cache/n812 ), .CK(clk), .RN(n6141), .Q(\D_cache/cache[0][123] ), .QN(n1059) );
  DFFRX1 \D_cache/cache_reg[1][123]  ( .D(\D_cache/n811 ), .CK(clk), .RN(n6141), .Q(\D_cache/cache[1][123] ), .QN(n2686) );
  DFFRX1 \D_cache/cache_reg[2][123]  ( .D(\D_cache/n810 ), .CK(clk), .RN(n6141), .Q(\D_cache/cache[2][123] ), .QN(n1060) );
  DFFRX1 \D_cache/cache_reg[3][123]  ( .D(\D_cache/n809 ), .CK(clk), .RN(n6141), .Q(\D_cache/cache[3][123] ), .QN(n2687) );
  DFFRX1 \D_cache/cache_reg[4][123]  ( .D(\D_cache/n808 ), .CK(clk), .RN(n6141), .Q(\D_cache/cache[4][123] ), .QN(n1214) );
  DFFRX1 \D_cache/cache_reg[5][123]  ( .D(\D_cache/n807 ), .CK(clk), .RN(n6141), .Q(\D_cache/cache[5][123] ), .QN(n2837) );
  DFFRX1 \D_cache/cache_reg[6][123]  ( .D(\D_cache/n806 ), .CK(clk), .RN(n6141), .Q(\D_cache/cache[6][123] ), .QN(n1058) );
  DFFRX1 \D_cache/cache_reg[7][123]  ( .D(\D_cache/n805 ), .CK(clk), .RN(n6141), .Q(\D_cache/cache[7][123] ), .QN(n2685) );
  DFFRX1 \D_cache/cache_reg[0][124]  ( .D(\D_cache/n804 ), .CK(clk), .RN(n6140), .Q(\D_cache/cache[0][124] ), .QN(n678) );
  DFFRX1 \D_cache/cache_reg[1][124]  ( .D(\D_cache/n803 ), .CK(clk), .RN(n6140), .Q(\D_cache/cache[1][124] ), .QN(n2296) );
  DFFRX1 \D_cache/cache_reg[2][124]  ( .D(\D_cache/n802 ), .CK(clk), .RN(n6140), .Q(\D_cache/cache[2][124] ), .QN(n999) );
  DFFRX1 \D_cache/cache_reg[3][124]  ( .D(\D_cache/n801 ), .CK(clk), .RN(n6140), .Q(\D_cache/cache[3][124] ), .QN(n2624) );
  DFFRX1 \D_cache/cache_reg[4][124]  ( .D(\D_cache/n800 ), .CK(clk), .RN(n6140), .Q(\D_cache/cache[4][124] ), .QN(n1187) );
  DFFRX1 \D_cache/cache_reg[5][124]  ( .D(\D_cache/n799 ), .CK(clk), .RN(n6140), .Q(\D_cache/cache[5][124] ), .QN(n2810) );
  DFFRX1 \D_cache/cache_reg[6][124]  ( .D(\D_cache/n798 ), .CK(clk), .RN(n6140), .Q(\D_cache/cache[6][124] ), .QN(n677) );
  DFFRX1 \D_cache/cache_reg[7][124]  ( .D(\D_cache/n797 ), .CK(clk), .RN(n6140), .Q(\D_cache/cache[7][124] ), .QN(n2295) );
  DFFRX1 \D_cache/cache_reg[0][125]  ( .D(\D_cache/n796 ), .CK(clk), .RN(n6140), .Q(\D_cache/cache[0][125] ), .QN(n1064) );
  DFFRX1 \D_cache/cache_reg[1][125]  ( .D(\D_cache/n795 ), .CK(clk), .RN(n6140), .Q(\D_cache/cache[1][125] ), .QN(n2692) );
  DFFRX1 \D_cache/cache_reg[2][125]  ( .D(\D_cache/n794 ), .CK(clk), .RN(n6140), .Q(\D_cache/cache[2][125] ), .QN(n1063) );
  DFFRX1 \D_cache/cache_reg[3][125]  ( .D(\D_cache/n793 ), .CK(clk), .RN(n6140), .Q(\D_cache/cache[3][125] ), .QN(n2691) );
  DFFRX1 \D_cache/cache_reg[4][125]  ( .D(\D_cache/n792 ), .CK(clk), .RN(n6139), .Q(\D_cache/cache[4][125] ), .QN(n1216) );
  DFFRX1 \D_cache/cache_reg[5][125]  ( .D(\D_cache/n791 ), .CK(clk), .RN(n6139), .Q(\D_cache/cache[5][125] ), .QN(n2839) );
  DFFRX1 \D_cache/cache_reg[6][125]  ( .D(\D_cache/n790 ), .CK(clk), .RN(n6139), .Q(\D_cache/cache[6][125] ), .QN(n1062) );
  DFFRX1 \D_cache/cache_reg[7][125]  ( .D(\D_cache/n789 ), .CK(clk), .RN(n6139), .Q(\D_cache/cache[7][125] ), .QN(n2690) );
  DFFRX1 \D_cache/cache_reg[0][126]  ( .D(\D_cache/n788 ), .CK(clk), .RN(n6139), .Q(\D_cache/cache[0][126] ), .QN(n1022) );
  DFFRX1 \D_cache/cache_reg[1][126]  ( .D(\D_cache/n787 ), .CK(clk), .RN(n6139), .Q(\D_cache/cache[1][126] ), .QN(n2648) );
  DFFRX1 \D_cache/cache_reg[2][126]  ( .D(\D_cache/n786 ), .CK(clk), .RN(n6139), .Q(\D_cache/cache[2][126] ), .QN(n1021) );
  DFFRX1 \D_cache/cache_reg[3][126]  ( .D(\D_cache/n785 ), .CK(clk), .RN(n6139), .Q(\D_cache/cache[3][126] ), .QN(n2647) );
  DFFRX1 \D_cache/cache_reg[4][126]  ( .D(\D_cache/n784 ), .CK(clk), .RN(n6139), .Q(\D_cache/cache[4][126] ), .QN(n1222) );
  DFFRX1 \D_cache/cache_reg[5][126]  ( .D(\D_cache/n783 ), .CK(clk), .RN(n6139), .Q(\D_cache/cache[5][126] ), .QN(n2845) );
  DFFRX1 \D_cache/cache_reg[6][126]  ( .D(\D_cache/n782 ), .CK(clk), .RN(n6139), .Q(\D_cache/cache[6][126] ), .QN(n702) );
  DFFRX1 \D_cache/cache_reg[7][126]  ( .D(\D_cache/n781 ), .CK(clk), .RN(n6139), .Q(\D_cache/cache[7][126] ), .QN(n2322) );
  DFFRX1 \D_cache/cache_reg[0][127]  ( .D(\D_cache/n780 ), .CK(clk), .RN(n6138), .Q(\D_cache/cache[0][127] ), .QN(n704) );
  DFFRX1 \D_cache/cache_reg[1][127]  ( .D(\D_cache/n779 ), .CK(clk), .RN(n6138), .Q(\D_cache/cache[1][127] ), .QN(n2324) );
  DFFRX1 \D_cache/cache_reg[2][127]  ( .D(\D_cache/n778 ), .CK(clk), .RN(n6138), .Q(\D_cache/cache[2][127] ), .QN(n1023) );
  DFFRX1 \D_cache/cache_reg[3][127]  ( .D(\D_cache/n777 ), .CK(clk), .RN(n6138), .Q(\D_cache/cache[3][127] ), .QN(n2649) );
  DFFRX1 \D_cache/cache_reg[4][127]  ( .D(\D_cache/n776 ), .CK(clk), .RN(n6138), .Q(\D_cache/cache[4][127] ), .QN(n1280) );
  DFFRX1 \D_cache/cache_reg[5][127]  ( .D(\D_cache/n775 ), .CK(clk), .RN(n6138), .Q(\D_cache/cache[5][127] ), .QN(n2912) );
  DFFRX1 \D_cache/cache_reg[6][127]  ( .D(\D_cache/n774 ), .CK(clk), .RN(n6138), .Q(\D_cache/cache[6][127] ), .QN(n703) );
  DFFRX1 \D_cache/cache_reg[7][127]  ( .D(\D_cache/n773 ), .CK(clk), .RN(n6138), .Q(\D_cache/cache[7][127] ), .QN(n2323) );
  DFFRX1 \D_cache/cache_reg[0][128]  ( .D(\D_cache/n772 ), .CK(clk), .RN(n6138), .Q(\D_cache/cache[0][128] ), .QN(n1304) );
  DFFRX1 \D_cache/cache_reg[1][128]  ( .D(\D_cache/n771 ), .CK(clk), .RN(n6138), .Q(\D_cache/cache[1][128] ), .QN(n2990) );
  DFFRX1 \D_cache/cache_reg[4][128]  ( .D(\D_cache/n768 ), .CK(clk), .RN(n6137), .Q(\D_cache/cache[4][128] ), .QN(n1273) );
  DFFRX1 \D_cache/cache_reg[5][128]  ( .D(\D_cache/n767 ), .CK(clk), .RN(n6137), .Q(\D_cache/cache[5][128] ), .QN(n2902) );
  DFFRX1 \D_cache/cache_reg[0][145]  ( .D(\D_cache/n636 ), .CK(clk), .RN(n6127), .Q(\D_cache/cache[0][145] ), .QN(n2955) );
  DFFRX1 \D_cache/cache_reg[1][145]  ( .D(\D_cache/n635 ), .CK(clk), .RN(n6126), .Q(\D_cache/cache[1][145] ), .QN(n1314) );
  DFFRX1 \D_cache/cache_reg[4][145]  ( .D(\D_cache/n632 ), .CK(clk), .RN(n6126), .Q(\D_cache/cache[4][145] ), .QN(n2953) );
  DFFRX1 \D_cache/cache_reg[5][145]  ( .D(\D_cache/n631 ), .CK(clk), .RN(n6126), .Q(\D_cache/cache[5][145] ), .QN(n1312) );
  DFFRX1 \D_cache/cache_reg[0][147]  ( .D(\D_cache/n620 ), .CK(clk), .RN(n6125), .Q(\D_cache/cache[0][147] ), .QN(n1334) );
  DFFRX1 \D_cache/cache_reg[1][147]  ( .D(\D_cache/n619 ), .CK(clk), .RN(n6125), .Q(\D_cache/cache[1][147] ), .QN(n2987) );
  DFFRX1 \D_cache/cache_reg[4][147]  ( .D(\D_cache/n616 ), .CK(clk), .RN(n6125), .Q(\D_cache/cache[4][147] ), .QN(n1335) );
  DFFRX1 \D_cache/cache_reg[5][147]  ( .D(\D_cache/n615 ), .CK(clk), .RN(n6125), .Q(\D_cache/cache[5][147] ), .QN(n2988) );
  DFFRX1 \D_cache/cache_reg[4][149]  ( .D(\D_cache/n600 ), .CK(clk), .RN(n6124), .Q(\D_cache/cache[4][149] ), .QN(n1272) );
  DFFRX1 \D_cache/cache_reg[0][150]  ( .D(\D_cache/n596 ), .CK(clk), .RN(n6123), .Q(\D_cache/cache[0][150] ), .QN(n2954) );
  DFFRX1 \D_cache/cache_reg[1][150]  ( .D(\D_cache/n595 ), .CK(clk), .RN(n6123), .Q(\D_cache/cache[1][150] ), .QN(n1313) );
  DFFRX1 \D_cache/cache_reg[4][150]  ( .D(\D_cache/n592 ), .CK(clk), .RN(n6123), .Q(\D_cache/cache[4][150] ), .QN(n1333) );
  DFFRX1 \D_cache/cache_reg[5][150]  ( .D(\D_cache/n591 ), .CK(clk), .RN(n6123), .Q(\D_cache/cache[5][150] ), .QN(n2986) );
  DFFRX1 \D_cache/cache_reg[0][153]  ( .D(\D_cache/n572 ), .CK(clk), .RN(n6121), .Q(\D_cache/cache[0][153] ), .QN(n1274) );
  DFFRX1 \D_cache/cache_reg[1][153]  ( .D(\D_cache/n571 ), .CK(clk), .RN(n6121), .Q(\D_cache/cache[1][153] ), .QN(n2903) );
  DFFRX1 \D_cache/cache_reg[2][153]  ( .D(\D_cache/n570 ), .CK(clk), .RN(n6121), .Q(\D_cache/cache[2][153] ), .QN(n1279) );
  DFFRX1 \D_cache/cache_reg[3][153]  ( .D(\D_cache/n569 ), .CK(clk), .RN(n6121), .Q(\D_cache/cache[3][153] ), .QN(n2911) );
  DFFRX1 \D_cache/cache_reg[4][153]  ( .D(\D_cache/n568 ), .CK(clk), .RN(n6121), .Q(\D_cache/cache[4][153] ), .QN(n1275) );
  DFFRX1 \D_cache/cache_reg[5][153]  ( .D(\D_cache/n567 ), .CK(clk), .RN(n6121), .Q(\D_cache/cache[5][153] ), .QN(n2904) );
  DFFRX1 \D_cache/cache_reg[6][153]  ( .D(\D_cache/n566 ), .CK(clk), .RN(n6121), .Q(\D_cache/cache[6][153] ), .QN(n1271) );
  DFFRX1 \D_cache/cache_reg[7][153]  ( .D(\D_cache/n565 ), .CK(clk), .RN(n6121), .Q(\D_cache/cache[7][153] ), .QN(n2895) );
  DFFRX1 \I_cache/cache_reg[5][0]  ( .D(n12839), .CK(clk), .RN(n6119), .Q(
        \I_cache/cache[5][0] ), .QN(n3127) );
  DFFRX1 \I_cache/cache_reg[6][0]  ( .D(n12838), .CK(clk), .RN(n6119), .Q(
        \I_cache/cache[6][0] ), .QN(n1530) );
  DFFRX1 \I_cache/cache_reg[7][0]  ( .D(n12845), .CK(clk), .RN(n6119), .Q(
        \I_cache/cache[7][0] ), .QN(n3217) );
  DFFRX1 \I_cache/cache_reg[5][1]  ( .D(n12832), .CK(clk), .RN(n6119), .Q(
        \I_cache/cache[5][1] ), .QN(n3199) );
  DFFRX1 \I_cache/cache_reg[6][1]  ( .D(n12831), .CK(clk), .RN(n6119), .Q(
        \I_cache/cache[6][1] ), .QN(n1577) );
  DFFRX1 \I_cache/cache_reg[7][1]  ( .D(n12830), .CK(clk), .RN(n6119), .Q(
        \I_cache/cache[7][1] ), .QN(n3264) );
  DFFRX1 \I_cache/cache_reg[5][2]  ( .D(n12824), .CK(clk), .RN(n6118), .Q(
        \I_cache/cache[5][2] ), .QN(n3196) );
  DFFRX1 \I_cache/cache_reg[6][2]  ( .D(n12823), .CK(clk), .RN(n6118), .Q(
        \I_cache/cache[6][2] ), .QN(n1575) );
  DFFRX1 \I_cache/cache_reg[7][2]  ( .D(n12822), .CK(clk), .RN(n6118), .Q(
        \I_cache/cache[7][2] ), .QN(n3263) );
  DFFRX1 \I_cache/cache_reg[5][3]  ( .D(n12816), .CK(clk), .RN(n6117), .Q(
        \I_cache/cache[5][3] ), .QN(n3193) );
  DFFRX1 \I_cache/cache_reg[6][3]  ( .D(n12815), .CK(clk), .RN(n6117), .Q(
        \I_cache/cache[6][3] ), .QN(n1573) );
  DFFRX1 \I_cache/cache_reg[7][3]  ( .D(n12814), .CK(clk), .RN(n6117), .Q(
        \I_cache/cache[7][3] ), .QN(n3261) );
  DFFRX1 \I_cache/cache_reg[5][4]  ( .D(n12808), .CK(clk), .RN(n6117), .Q(
        \I_cache/cache[5][4] ), .QN(n3190) );
  DFFRX1 \I_cache/cache_reg[6][4]  ( .D(n12807), .CK(clk), .RN(n6117), .Q(
        \I_cache/cache[6][4] ), .QN(n1571) );
  DFFRX1 \I_cache/cache_reg[7][4]  ( .D(n12806), .CK(clk), .RN(n6117), .Q(
        \I_cache/cache[7][4] ), .QN(n3259) );
  DFFRX1 \I_cache/cache_reg[5][5]  ( .D(n12800), .CK(clk), .RN(n6116), .Q(
        \I_cache/cache[5][5] ), .QN(n3187) );
  DFFRX1 \I_cache/cache_reg[6][5]  ( .D(n12799), .CK(clk), .RN(n6116), .Q(
        \I_cache/cache[6][5] ), .QN(n1569) );
  DFFRX1 \I_cache/cache_reg[7][5]  ( .D(n12798), .CK(clk), .RN(n6116), .Q(
        \I_cache/cache[7][5] ), .QN(n3257) );
  DFFRX1 \I_cache/cache_reg[5][6]  ( .D(n12792), .CK(clk), .RN(n6115), .Q(
        \I_cache/cache[5][6] ), .QN(n3184) );
  DFFRX1 \I_cache/cache_reg[6][6]  ( .D(n12791), .CK(clk), .RN(n6115), .Q(
        \I_cache/cache[6][6] ), .QN(n1567) );
  DFFRX1 \I_cache/cache_reg[7][6]  ( .D(n12790), .CK(clk), .RN(n6115), .Q(
        \I_cache/cache[7][6] ), .QN(n3255) );
  DFFRX1 \I_cache/cache_reg[5][7]  ( .D(n12784), .CK(clk), .RN(n6115), .Q(
        \I_cache/cache[5][7] ), .QN(n3181) );
  DFFRX1 \I_cache/cache_reg[6][7]  ( .D(n12783), .CK(clk), .RN(n6115), .Q(
        \I_cache/cache[6][7] ), .QN(n1565) );
  DFFRX1 \I_cache/cache_reg[7][7]  ( .D(n12782), .CK(clk), .RN(n6115), .Q(
        \I_cache/cache[7][7] ), .QN(n3253) );
  DFFRX1 \I_cache/cache_reg[5][8]  ( .D(n12776), .CK(clk), .RN(n6114), .Q(
        \I_cache/cache[5][8] ), .QN(n3178) );
  DFFRX1 \I_cache/cache_reg[6][8]  ( .D(n12775), .CK(clk), .RN(n6114), .Q(
        \I_cache/cache[6][8] ), .QN(n1563) );
  DFFRX1 \I_cache/cache_reg[7][8]  ( .D(n12774), .CK(clk), .RN(n6114), .Q(
        \I_cache/cache[7][8] ), .QN(n3251) );
  DFFRX1 \I_cache/cache_reg[5][9]  ( .D(n12768), .CK(clk), .RN(n6113), .Q(
        \I_cache/cache[5][9] ), .QN(n3175) );
  DFFRX1 \I_cache/cache_reg[6][9]  ( .D(n12767), .CK(clk), .RN(n6113), .Q(
        \I_cache/cache[6][9] ), .QN(n1561) );
  DFFRX1 \I_cache/cache_reg[7][9]  ( .D(n12766), .CK(clk), .RN(n6113), .Q(
        \I_cache/cache[7][9] ), .QN(n3249) );
  DFFRX1 \I_cache/cache_reg[5][10]  ( .D(n12760), .CK(clk), .RN(n6113), .Q(
        \I_cache/cache[5][10] ), .QN(n3172) );
  DFFRX1 \I_cache/cache_reg[6][10]  ( .D(n12759), .CK(clk), .RN(n6113), .Q(
        \I_cache/cache[6][10] ), .QN(n1559) );
  DFFRX1 \I_cache/cache_reg[7][10]  ( .D(n12758), .CK(clk), .RN(n6113), .Q(
        \I_cache/cache[7][10] ), .QN(n3247) );
  DFFRX1 \I_cache/cache_reg[5][11]  ( .D(n12752), .CK(clk), .RN(n6112), .Q(
        \I_cache/cache[5][11] ), .QN(n3169) );
  DFFRX1 \I_cache/cache_reg[6][11]  ( .D(n12751), .CK(clk), .RN(n6112), .Q(
        \I_cache/cache[6][11] ), .QN(n1557) );
  DFFRX1 \I_cache/cache_reg[7][11]  ( .D(n12750), .CK(clk), .RN(n6112), .Q(
        \I_cache/cache[7][11] ), .QN(n3245) );
  DFFRX1 \I_cache/cache_reg[5][12]  ( .D(n12744), .CK(clk), .RN(n6111), .Q(
        \I_cache/cache[5][12] ), .QN(n3166) );
  DFFRX1 \I_cache/cache_reg[6][12]  ( .D(n12743), .CK(clk), .RN(n6111), .Q(
        \I_cache/cache[6][12] ), .QN(n1555) );
  DFFRX1 \I_cache/cache_reg[7][12]  ( .D(n12742), .CK(clk), .RN(n6111), .Q(
        \I_cache/cache[7][12] ), .QN(n3243) );
  DFFRX1 \I_cache/cache_reg[5][13]  ( .D(n12736), .CK(clk), .RN(n6111), .Q(
        \I_cache/cache[5][13] ), .QN(n3163) );
  DFFRX1 \I_cache/cache_reg[6][13]  ( .D(n12735), .CK(clk), .RN(n6111), .Q(
        \I_cache/cache[6][13] ), .QN(n1553) );
  DFFRX1 \I_cache/cache_reg[7][13]  ( .D(n12734), .CK(clk), .RN(n6111), .Q(
        \I_cache/cache[7][13] ), .QN(n3241) );
  DFFRX1 \I_cache/cache_reg[5][14]  ( .D(n12728), .CK(clk), .RN(n6110), .Q(
        \I_cache/cache[5][14] ), .QN(n3160) );
  DFFRX1 \I_cache/cache_reg[6][14]  ( .D(n12727), .CK(clk), .RN(n6110), .Q(
        \I_cache/cache[6][14] ), .QN(n1551) );
  DFFRX1 \I_cache/cache_reg[7][14]  ( .D(n12726), .CK(clk), .RN(n6110), .Q(
        \I_cache/cache[7][14] ), .QN(n3239) );
  DFFRX1 \I_cache/cache_reg[5][15]  ( .D(n12720), .CK(clk), .RN(n6109), .Q(
        \I_cache/cache[5][15] ), .QN(n3157) );
  DFFRX1 \I_cache/cache_reg[6][15]  ( .D(n12719), .CK(clk), .RN(n6109), .Q(
        \I_cache/cache[6][15] ), .QN(n1549) );
  DFFRX1 \I_cache/cache_reg[7][15]  ( .D(n12718), .CK(clk), .RN(n6109), .Q(
        \I_cache/cache[7][15] ), .QN(n3237) );
  DFFRX1 \I_cache/cache_reg[5][16]  ( .D(n12712), .CK(clk), .RN(n6109), .Q(
        \I_cache/cache[5][16] ), .QN(n3154) );
  DFFRX1 \I_cache/cache_reg[6][16]  ( .D(n12711), .CK(clk), .RN(n6109), .Q(
        \I_cache/cache[6][16] ), .QN(n1547) );
  DFFRX1 \I_cache/cache_reg[7][16]  ( .D(n12710), .CK(clk), .RN(n6109), .Q(
        \I_cache/cache[7][16] ), .QN(n3235) );
  DFFRX1 \I_cache/cache_reg[5][17]  ( .D(n12704), .CK(clk), .RN(n6108), .Q(
        \I_cache/cache[5][17] ), .QN(n3151) );
  DFFRX1 \I_cache/cache_reg[6][17]  ( .D(n12703), .CK(clk), .RN(n6108), .Q(
        \I_cache/cache[6][17] ), .QN(n1545) );
  DFFRX1 \I_cache/cache_reg[7][17]  ( .D(n12702), .CK(clk), .RN(n6108), .Q(
        \I_cache/cache[7][17] ), .QN(n3233) );
  DFFRX1 \I_cache/cache_reg[5][18]  ( .D(n12696), .CK(clk), .RN(n6107), .Q(
        \I_cache/cache[5][18] ), .QN(n3148) );
  DFFRX1 \I_cache/cache_reg[6][18]  ( .D(n12695), .CK(clk), .RN(n6107), .Q(
        \I_cache/cache[6][18] ), .QN(n1544) );
  DFFRX1 \I_cache/cache_reg[7][18]  ( .D(n12694), .CK(clk), .RN(n6107), .Q(
        \I_cache/cache[7][18] ), .QN(n3231) );
  DFFRX1 \I_cache/cache_reg[5][19]  ( .D(n12688), .CK(clk), .RN(n6107), .Q(
        \I_cache/cache[5][19] ), .QN(n3284) );
  DFFRX1 \I_cache/cache_reg[6][19]  ( .D(n12687), .CK(clk), .RN(n6107), .Q(
        \I_cache/cache[6][19] ), .QN(n1600) );
  DFFRX1 \I_cache/cache_reg[7][19]  ( .D(n12686), .CK(clk), .RN(n6107), .Q(
        \I_cache/cache[7][19] ), .QN(n3287) );
  DFFRX1 \I_cache/cache_reg[5][20]  ( .D(n12680), .CK(clk), .RN(n6106), .Q(
        \I_cache/cache[5][20] ), .QN(n3145) );
  DFFRX1 \I_cache/cache_reg[6][20]  ( .D(n12679), .CK(clk), .RN(n6106), .Q(
        \I_cache/cache[6][20] ), .QN(n1542) );
  DFFRX1 \I_cache/cache_reg[7][20]  ( .D(n12678), .CK(clk), .RN(n6106), .Q(
        \I_cache/cache[7][20] ), .QN(n3229) );
  DFFRX1 \I_cache/cache_reg[5][21]  ( .D(n12672), .CK(clk), .RN(n6105), .Q(
        \I_cache/cache[5][21] ), .QN(n3142) );
  DFFRX1 \I_cache/cache_reg[6][21]  ( .D(n12671), .CK(clk), .RN(n6105), .Q(
        \I_cache/cache[6][21] ), .QN(n1540) );
  DFFRX1 \I_cache/cache_reg[7][21]  ( .D(n12670), .CK(clk), .RN(n6105), .Q(
        \I_cache/cache[7][21] ), .QN(n3227) );
  DFFRX1 \I_cache/cache_reg[5][22]  ( .D(n12664), .CK(clk), .RN(n6105), .Q(
        \I_cache/cache[5][22] ), .QN(n3139) );
  DFFRX1 \I_cache/cache_reg[6][22]  ( .D(n12663), .CK(clk), .RN(n6105), .Q(
        \I_cache/cache[6][22] ), .QN(n1538) );
  DFFRX1 \I_cache/cache_reg[7][22]  ( .D(n12662), .CK(clk), .RN(n6105), .Q(
        \I_cache/cache[7][22] ), .QN(n3225) );
  DFFRX1 \I_cache/cache_reg[5][23]  ( .D(n12656), .CK(clk), .RN(n6104), .Q(
        \I_cache/cache[5][23] ), .QN(n3136) );
  DFFRX1 \I_cache/cache_reg[6][23]  ( .D(n12655), .CK(clk), .RN(n6104), .Q(
        \I_cache/cache[6][23] ), .QN(n1536) );
  DFFRX1 \I_cache/cache_reg[7][23]  ( .D(n12654), .CK(clk), .RN(n6104), .Q(
        \I_cache/cache[7][23] ), .QN(n3223) );
  DFFRX1 \I_cache/cache_reg[5][24]  ( .D(n12648), .CK(clk), .RN(n6103), .Q(
        \I_cache/cache[5][24] ), .QN(n3133) );
  DFFRX1 \I_cache/cache_reg[6][24]  ( .D(n12647), .CK(clk), .RN(n6103), .Q(
        \I_cache/cache[6][24] ), .QN(n1534) );
  DFFRX1 \I_cache/cache_reg[7][24]  ( .D(n12646), .CK(clk), .RN(n6103), .Q(
        \I_cache/cache[7][24] ), .QN(n3221) );
  DFFRX1 \I_cache/cache_reg[5][25]  ( .D(n12640), .CK(clk), .RN(n6103), .Q(
        \I_cache/cache[5][25] ), .QN(n3130) );
  DFFRX1 \I_cache/cache_reg[6][25]  ( .D(n12639), .CK(clk), .RN(n6103), .Q(
        \I_cache/cache[6][25] ), .QN(n1532) );
  DFFRX1 \I_cache/cache_reg[7][25]  ( .D(n12638), .CK(clk), .RN(n6103), .Q(
        \I_cache/cache[7][25] ), .QN(n3219) );
  DFFRX1 \I_cache/cache_reg[5][26]  ( .D(n12632), .CK(clk), .RN(n6102), .Q(
        \I_cache/cache[5][26] ), .QN(n3214) );
  DFFRX1 \I_cache/cache_reg[6][26]  ( .D(n12631), .CK(clk), .RN(n6102), .Q(
        \I_cache/cache[6][26] ), .QN(n1588) );
  DFFRX1 \I_cache/cache_reg[7][26]  ( .D(n12630), .CK(clk), .RN(n6102), .Q(
        \I_cache/cache[7][26] ), .QN(n3275) );
  DFFRX1 \I_cache/cache_reg[5][27]  ( .D(n12624), .CK(clk), .RN(n6101), .Q(
        \I_cache/cache[5][27] ), .QN(n3211) );
  DFFRX1 \I_cache/cache_reg[6][27]  ( .D(n12623), .CK(clk), .RN(n6101), .Q(
        \I_cache/cache[6][27] ), .QN(n1586) );
  DFFRX1 \I_cache/cache_reg[7][27]  ( .D(n12622), .CK(clk), .RN(n6101), .Q(
        \I_cache/cache[7][27] ), .QN(n3273) );
  DFFRX1 \I_cache/cache_reg[5][28]  ( .D(n12616), .CK(clk), .RN(n6101), .Q(
        \I_cache/cache[5][28] ), .QN(n3208) );
  DFFRX1 \I_cache/cache_reg[6][28]  ( .D(n12615), .CK(clk), .RN(n6101), .Q(
        \I_cache/cache[6][28] ), .QN(n1584) );
  DFFRX1 \I_cache/cache_reg[7][28]  ( .D(n12614), .CK(clk), .RN(n6101), .Q(
        \I_cache/cache[7][28] ), .QN(n3271) );
  DFFRX1 \I_cache/cache_reg[5][29]  ( .D(n12608), .CK(clk), .RN(n6100), .Q(
        \I_cache/cache[5][29] ), .QN(n3205) );
  DFFRX1 \I_cache/cache_reg[6][29]  ( .D(n12607), .CK(clk), .RN(n6100), .Q(
        \I_cache/cache[6][29] ), .QN(n1582) );
  DFFRX1 \I_cache/cache_reg[7][29]  ( .D(n12606), .CK(clk), .RN(n6100), .Q(
        \I_cache/cache[7][29] ), .QN(n3269) );
  DFFRX1 \I_cache/cache_reg[5][30]  ( .D(n12600), .CK(clk), .RN(n6099), .Q(
        \I_cache/cache[5][30] ), .QN(n3202) );
  DFFRX1 \I_cache/cache_reg[6][30]  ( .D(n12599), .CK(clk), .RN(n6099), .Q(
        \I_cache/cache[6][30] ), .QN(n1580) );
  DFFRX1 \I_cache/cache_reg[7][30]  ( .D(n12598), .CK(clk), .RN(n6099), .Q(
        \I_cache/cache[7][30] ), .QN(n3267) );
  DFFRX1 \I_cache/cache_reg[3][32]  ( .D(n12586), .CK(clk), .RN(n6098), .Q(
        \I_cache/cache[3][32] ), .QN(n3382) );
  DFFRX1 \I_cache/cache_reg[4][32]  ( .D(n12585), .CK(clk), .RN(n6098), .Q(
        \I_cache/cache[4][32] ), .QN(n1693) );
  DFFRX1 \I_cache/cache_reg[5][32]  ( .D(n12584), .CK(clk), .RN(n6098), .Q(
        \I_cache/cache[5][32] ), .QN(n3381) );
  DFFRX1 \I_cache/cache_reg[6][32]  ( .D(n12583), .CK(clk), .RN(n6098), .Q(
        \I_cache/cache[6][32] ), .QN(n1790) );
  DFFRX1 \I_cache/cache_reg[7][32]  ( .D(n12582), .CK(clk), .RN(n6098), .Q(
        \I_cache/cache[7][32] ), .QN(n3478) );
  DFFRX1 \I_cache/cache_reg[3][33]  ( .D(n12578), .CK(clk), .RN(n6098), .Q(
        \I_cache/cache[3][33] ), .QN(n3454) );
  DFFRX1 \I_cache/cache_reg[4][33]  ( .D(n12577), .CK(clk), .RN(n6097), .Q(
        \I_cache/cache[4][33] ), .QN(n1765) );
  DFFRX1 \I_cache/cache_reg[5][33]  ( .D(n12576), .CK(clk), .RN(n6097), .Q(
        \I_cache/cache[5][33] ), .QN(n3453) );
  DFFRX1 \I_cache/cache_reg[6][33]  ( .D(n12575), .CK(clk), .RN(n6097), .Q(
        \I_cache/cache[6][33] ), .QN(n1834) );
  DFFRX1 \I_cache/cache_reg[7][33]  ( .D(n12574), .CK(clk), .RN(n6097), .Q(
        \I_cache/cache[7][33] ), .QN(n3522) );
  DFFRX1 \I_cache/cache_reg[3][34]  ( .D(n12570), .CK(clk), .RN(n6097), .Q(
        \I_cache/cache[3][34] ), .QN(n3451) );
  DFFRX1 \I_cache/cache_reg[4][34]  ( .D(n12569), .CK(clk), .RN(n6097), .Q(
        \I_cache/cache[4][34] ), .QN(n1762) );
  DFFRX1 \I_cache/cache_reg[5][34]  ( .D(n12568), .CK(clk), .RN(n6097), .Q(
        \I_cache/cache[5][34] ), .QN(n3450) );
  DFFRX1 \I_cache/cache_reg[6][34]  ( .D(n12567), .CK(clk), .RN(n6097), .Q(
        \I_cache/cache[6][34] ), .QN(n1833) );
  DFFRX1 \I_cache/cache_reg[7][34]  ( .D(n12566), .CK(clk), .RN(n6097), .Q(
        \I_cache/cache[7][34] ), .QN(n3521) );
  DFFRX1 \I_cache/cache_reg[3][35]  ( .D(n12562), .CK(clk), .RN(n6096), .Q(
        \I_cache/cache[3][35] ), .QN(n3448) );
  DFFRX1 \I_cache/cache_reg[4][35]  ( .D(n12561), .CK(clk), .RN(n6096), .Q(
        \I_cache/cache[4][35] ), .QN(n1759) );
  DFFRX1 \I_cache/cache_reg[5][35]  ( .D(n12560), .CK(clk), .RN(n6096), .Q(
        \I_cache/cache[5][35] ), .QN(n3447) );
  DFFRX1 \I_cache/cache_reg[6][35]  ( .D(n12559), .CK(clk), .RN(n6096), .Q(
        \I_cache/cache[6][35] ), .QN(n1832) );
  DFFRX1 \I_cache/cache_reg[7][35]  ( .D(n12558), .CK(clk), .RN(n6096), .Q(
        \I_cache/cache[7][35] ), .QN(n3520) );
  DFFRX1 \I_cache/cache_reg[3][36]  ( .D(n12554), .CK(clk), .RN(n6096), .Q(
        \I_cache/cache[3][36] ), .QN(n3445) );
  DFFRX1 \I_cache/cache_reg[4][36]  ( .D(n12553), .CK(clk), .RN(n6095), .Q(
        \I_cache/cache[4][36] ), .QN(n1756) );
  DFFRX1 \I_cache/cache_reg[5][36]  ( .D(n12552), .CK(clk), .RN(n6095), .Q(
        \I_cache/cache[5][36] ), .QN(n3444) );
  DFFRX1 \I_cache/cache_reg[6][36]  ( .D(n12551), .CK(clk), .RN(n6095), .Q(
        \I_cache/cache[6][36] ), .QN(n1830) );
  DFFRX1 \I_cache/cache_reg[7][36]  ( .D(n12550), .CK(clk), .RN(n6095), .Q(
        \I_cache/cache[7][36] ), .QN(n3518) );
  DFFRX1 \I_cache/cache_reg[3][37]  ( .D(n12546), .CK(clk), .RN(n6095), .Q(
        \I_cache/cache[3][37] ), .QN(n3442) );
  DFFRX1 \I_cache/cache_reg[4][37]  ( .D(n12545), .CK(clk), .RN(n6095), .Q(
        \I_cache/cache[4][37] ), .QN(n1753) );
  DFFRX1 \I_cache/cache_reg[5][37]  ( .D(n12544), .CK(clk), .RN(n6095), .Q(
        \I_cache/cache[5][37] ), .QN(n3441) );
  DFFRX1 \I_cache/cache_reg[6][37]  ( .D(n12543), .CK(clk), .RN(n6095), .Q(
        \I_cache/cache[6][37] ), .QN(n1829) );
  DFFRX1 \I_cache/cache_reg[7][37]  ( .D(n12542), .CK(clk), .RN(n6095), .Q(
        \I_cache/cache[7][37] ), .QN(n3517) );
  DFFRX1 \I_cache/cache_reg[3][38]  ( .D(n12538), .CK(clk), .RN(n6094), .Q(
        \I_cache/cache[3][38] ), .QN(n3439) );
  DFFRX1 \I_cache/cache_reg[4][38]  ( .D(n12537), .CK(clk), .RN(n6094), .Q(
        \I_cache/cache[4][38] ), .QN(n1750) );
  DFFRX1 \I_cache/cache_reg[5][38]  ( .D(n12536), .CK(clk), .RN(n6094), .Q(
        \I_cache/cache[5][38] ), .QN(n3438) );
  DFFRX1 \I_cache/cache_reg[6][38]  ( .D(n12535), .CK(clk), .RN(n6094), .Q(
        \I_cache/cache[6][38] ), .QN(n1827) );
  DFFRX1 \I_cache/cache_reg[7][38]  ( .D(n12534), .CK(clk), .RN(n6094), .Q(
        \I_cache/cache[7][38] ), .QN(n3515) );
  DFFRX1 \I_cache/cache_reg[3][39]  ( .D(n12530), .CK(clk), .RN(n6094), .Q(
        \I_cache/cache[3][39] ), .QN(n3436) );
  DFFRX1 \I_cache/cache_reg[4][39]  ( .D(n12529), .CK(clk), .RN(n6093), .Q(
        \I_cache/cache[4][39] ), .QN(n1747) );
  DFFRX1 \I_cache/cache_reg[5][39]  ( .D(n12528), .CK(clk), .RN(n6093), .Q(
        \I_cache/cache[5][39] ), .QN(n3435) );
  DFFRX1 \I_cache/cache_reg[6][39]  ( .D(n12527), .CK(clk), .RN(n6093), .Q(
        \I_cache/cache[6][39] ), .QN(n1825) );
  DFFRX1 \I_cache/cache_reg[7][39]  ( .D(n12526), .CK(clk), .RN(n6093), .Q(
        \I_cache/cache[7][39] ), .QN(n3513) );
  DFFRX1 \I_cache/cache_reg[3][40]  ( .D(n12522), .CK(clk), .RN(n6093), .Q(
        \I_cache/cache[3][40] ), .QN(n3433) );
  DFFRX1 \I_cache/cache_reg[4][40]  ( .D(n12521), .CK(clk), .RN(n6093), .Q(
        \I_cache/cache[4][40] ), .QN(n1744) );
  DFFRX1 \I_cache/cache_reg[5][40]  ( .D(n12520), .CK(clk), .RN(n6093), .Q(
        \I_cache/cache[5][40] ), .QN(n3432) );
  DFFRX1 \I_cache/cache_reg[6][40]  ( .D(n12519), .CK(clk), .RN(n6093), .Q(
        \I_cache/cache[6][40] ), .QN(n1823) );
  DFFRX1 \I_cache/cache_reg[7][40]  ( .D(n12518), .CK(clk), .RN(n6093), .Q(
        \I_cache/cache[7][40] ), .QN(n3511) );
  DFFRX1 \I_cache/cache_reg[3][41]  ( .D(n12514), .CK(clk), .RN(n6092), .Q(
        \I_cache/cache[3][41] ), .QN(n3430) );
  DFFRX1 \I_cache/cache_reg[4][41]  ( .D(n12513), .CK(clk), .RN(n6092), .Q(
        \I_cache/cache[4][41] ), .QN(n1741) );
  DFFRX1 \I_cache/cache_reg[5][41]  ( .D(n12512), .CK(clk), .RN(n6092), .Q(
        \I_cache/cache[5][41] ), .QN(n3429) );
  DFFRX1 \I_cache/cache_reg[6][41]  ( .D(n12511), .CK(clk), .RN(n6092), .Q(
        \I_cache/cache[6][41] ), .QN(n1821) );
  DFFRX1 \I_cache/cache_reg[7][41]  ( .D(n12510), .CK(clk), .RN(n6092), .Q(
        \I_cache/cache[7][41] ), .QN(n3509) );
  DFFRX1 \I_cache/cache_reg[3][42]  ( .D(n12506), .CK(clk), .RN(n6092), .Q(
        \I_cache/cache[3][42] ), .QN(n3427) );
  DFFRX1 \I_cache/cache_reg[4][42]  ( .D(n12505), .CK(clk), .RN(n6091), .Q(
        \I_cache/cache[4][42] ), .QN(n1738) );
  DFFRX1 \I_cache/cache_reg[5][42]  ( .D(n12504), .CK(clk), .RN(n6091), .Q(
        \I_cache/cache[5][42] ), .QN(n3426) );
  DFFRX1 \I_cache/cache_reg[6][42]  ( .D(n12503), .CK(clk), .RN(n6091), .Q(
        \I_cache/cache[6][42] ), .QN(n1819) );
  DFFRX1 \I_cache/cache_reg[7][42]  ( .D(n12502), .CK(clk), .RN(n6091), .Q(
        \I_cache/cache[7][42] ), .QN(n3507) );
  DFFRX1 \I_cache/cache_reg[3][43]  ( .D(n12498), .CK(clk), .RN(n6091), .Q(
        \I_cache/cache[3][43] ), .QN(n3424) );
  DFFRX1 \I_cache/cache_reg[4][43]  ( .D(n12497), .CK(clk), .RN(n6091), .Q(
        \I_cache/cache[4][43] ), .QN(n1735) );
  DFFRX1 \I_cache/cache_reg[5][43]  ( .D(n12496), .CK(clk), .RN(n6091), .Q(
        \I_cache/cache[5][43] ), .QN(n3423) );
  DFFRX1 \I_cache/cache_reg[6][43]  ( .D(n12495), .CK(clk), .RN(n6091), .Q(
        \I_cache/cache[6][43] ), .QN(n1817) );
  DFFRX1 \I_cache/cache_reg[7][43]  ( .D(n12494), .CK(clk), .RN(n6091), .Q(
        \I_cache/cache[7][43] ), .QN(n3505) );
  DFFRX1 \I_cache/cache_reg[3][44]  ( .D(n12490), .CK(clk), .RN(n6090), .Q(
        \I_cache/cache[3][44] ), .QN(n3421) );
  DFFRX1 \I_cache/cache_reg[4][44]  ( .D(n12489), .CK(clk), .RN(n6090), .Q(
        \I_cache/cache[4][44] ), .QN(n1732) );
  DFFRX1 \I_cache/cache_reg[5][44]  ( .D(n12488), .CK(clk), .RN(n6090), .Q(
        \I_cache/cache[5][44] ), .QN(n3420) );
  DFFRX1 \I_cache/cache_reg[6][44]  ( .D(n12487), .CK(clk), .RN(n6090), .Q(
        \I_cache/cache[6][44] ), .QN(n1815) );
  DFFRX1 \I_cache/cache_reg[7][44]  ( .D(n12486), .CK(clk), .RN(n6090), .Q(
        \I_cache/cache[7][44] ), .QN(n3503) );
  DFFRX1 \I_cache/cache_reg[3][45]  ( .D(n12482), .CK(clk), .RN(n6090), .Q(
        \I_cache/cache[3][45] ), .QN(n3418) );
  DFFRX1 \I_cache/cache_reg[4][45]  ( .D(n12481), .CK(clk), .RN(n6089), .Q(
        \I_cache/cache[4][45] ), .QN(n1729) );
  DFFRX1 \I_cache/cache_reg[5][45]  ( .D(n12480), .CK(clk), .RN(n6089), .Q(
        \I_cache/cache[5][45] ), .QN(n3417) );
  DFFRX1 \I_cache/cache_reg[6][45]  ( .D(n12479), .CK(clk), .RN(n6089), .Q(
        \I_cache/cache[6][45] ), .QN(n1813) );
  DFFRX1 \I_cache/cache_reg[7][45]  ( .D(n12478), .CK(clk), .RN(n6089), .Q(
        \I_cache/cache[7][45] ), .QN(n3501) );
  DFFRX1 \I_cache/cache_reg[3][46]  ( .D(n12474), .CK(clk), .RN(n6089), .Q(
        \I_cache/cache[3][46] ), .QN(n3415) );
  DFFRX1 \I_cache/cache_reg[4][46]  ( .D(n12473), .CK(clk), .RN(n6089), .Q(
        \I_cache/cache[4][46] ), .QN(n1726) );
  DFFRX1 \I_cache/cache_reg[5][46]  ( .D(n12472), .CK(clk), .RN(n6089), .Q(
        \I_cache/cache[5][46] ), .QN(n3414) );
  DFFRX1 \I_cache/cache_reg[6][46]  ( .D(n12471), .CK(clk), .RN(n6089), .Q(
        \I_cache/cache[6][46] ), .QN(n1811) );
  DFFRX1 \I_cache/cache_reg[7][46]  ( .D(n12470), .CK(clk), .RN(n6089), .Q(
        \I_cache/cache[7][46] ), .QN(n3499) );
  DFFRX1 \I_cache/cache_reg[3][47]  ( .D(n12466), .CK(clk), .RN(n6088), .Q(
        \I_cache/cache[3][47] ), .QN(n3412) );
  DFFRX1 \I_cache/cache_reg[4][47]  ( .D(n12465), .CK(clk), .RN(n6088), .Q(
        \I_cache/cache[4][47] ), .QN(n1723) );
  DFFRX1 \I_cache/cache_reg[5][47]  ( .D(n12464), .CK(clk), .RN(n6088), .Q(
        \I_cache/cache[5][47] ), .QN(n3411) );
  DFFRX1 \I_cache/cache_reg[6][47]  ( .D(n12463), .CK(clk), .RN(n6088), .Q(
        \I_cache/cache[6][47] ), .QN(n1809) );
  DFFRX1 \I_cache/cache_reg[7][47]  ( .D(n12462), .CK(clk), .RN(n6088), .Q(
        \I_cache/cache[7][47] ), .QN(n3497) );
  DFFRX1 \I_cache/cache_reg[3][48]  ( .D(n12458), .CK(clk), .RN(n6088), .Q(
        \I_cache/cache[3][48] ), .QN(n3409) );
  DFFRX1 \I_cache/cache_reg[4][48]  ( .D(n12457), .CK(clk), .RN(n6087), .Q(
        \I_cache/cache[4][48] ), .QN(n1720) );
  DFFRX1 \I_cache/cache_reg[5][48]  ( .D(n12456), .CK(clk), .RN(n6087), .Q(
        \I_cache/cache[5][48] ), .QN(n3408) );
  DFFRX1 \I_cache/cache_reg[6][48]  ( .D(n12455), .CK(clk), .RN(n6087), .Q(
        \I_cache/cache[6][48] ), .QN(n1807) );
  DFFRX1 \I_cache/cache_reg[7][48]  ( .D(n12454), .CK(clk), .RN(n6087), .Q(
        \I_cache/cache[7][48] ), .QN(n3495) );
  DFFRX1 \I_cache/cache_reg[3][49]  ( .D(n12450), .CK(clk), .RN(n6087), .Q(
        \I_cache/cache[3][49] ), .QN(n3406) );
  DFFRX1 \I_cache/cache_reg[4][49]  ( .D(n12449), .CK(clk), .RN(n6087), .Q(
        \I_cache/cache[4][49] ), .QN(n1717) );
  DFFRX1 \I_cache/cache_reg[5][49]  ( .D(n12448), .CK(clk), .RN(n6087), .Q(
        \I_cache/cache[5][49] ), .QN(n3405) );
  DFFRX1 \I_cache/cache_reg[6][49]  ( .D(n12447), .CK(clk), .RN(n6087), .Q(
        \I_cache/cache[6][49] ), .QN(n1805) );
  DFFRX1 \I_cache/cache_reg[7][49]  ( .D(n12446), .CK(clk), .RN(n6087), .Q(
        \I_cache/cache[7][49] ), .QN(n3493) );
  DFFRX1 \I_cache/cache_reg[3][50]  ( .D(n12442), .CK(clk), .RN(n6086), .Q(
        \I_cache/cache[3][50] ), .QN(n3403) );
  DFFRX1 \I_cache/cache_reg[4][50]  ( .D(n12441), .CK(clk), .RN(n6086), .Q(
        \I_cache/cache[4][50] ), .QN(n1714) );
  DFFRX1 \I_cache/cache_reg[5][50]  ( .D(n12440), .CK(clk), .RN(n6086), .Q(
        \I_cache/cache[5][50] ), .QN(n3402) );
  DFFRX1 \I_cache/cache_reg[6][50]  ( .D(n12439), .CK(clk), .RN(n6086), .Q(
        \I_cache/cache[6][50] ), .QN(n1803) );
  DFFRX1 \I_cache/cache_reg[7][50]  ( .D(n12438), .CK(clk), .RN(n6086), .Q(
        \I_cache/cache[7][50] ), .QN(n3491) );
  DFFRX1 \I_cache/cache_reg[3][51]  ( .D(n12434), .CK(clk), .RN(n6086), .Q(
        \I_cache/cache[3][51] ), .QN(n3540) );
  DFFRX1 \I_cache/cache_reg[4][51]  ( .D(n12433), .CK(clk), .RN(n6085), .Q(
        \I_cache/cache[4][51] ), .QN(n1852) );
  DFFRX1 \I_cache/cache_reg[5][51]  ( .D(n12432), .CK(clk), .RN(n6085), .Q(
        \I_cache/cache[5][51] ), .QN(n3539) );
  DFFRX1 \I_cache/cache_reg[6][51]  ( .D(n12431), .CK(clk), .RN(n6085), .Q(
        \I_cache/cache[6][51] ), .QN(n1855) );
  DFFRX1 \I_cache/cache_reg[7][51]  ( .D(n12430), .CK(clk), .RN(n6085), .Q(
        \I_cache/cache[7][51] ), .QN(n3542) );
  DFFRX1 \I_cache/cache_reg[3][52]  ( .D(n12426), .CK(clk), .RN(n6085), .Q(
        \I_cache/cache[3][52] ), .QN(n3400) );
  DFFRX1 \I_cache/cache_reg[4][52]  ( .D(n12425), .CK(clk), .RN(n6085), .Q(
        \I_cache/cache[4][52] ), .QN(n1711) );
  DFFRX1 \I_cache/cache_reg[5][52]  ( .D(n12424), .CK(clk), .RN(n6085), .Q(
        \I_cache/cache[5][52] ), .QN(n3399) );
  DFFRX1 \I_cache/cache_reg[6][52]  ( .D(n12423), .CK(clk), .RN(n6085), .Q(
        \I_cache/cache[6][52] ), .QN(n1801) );
  DFFRX1 \I_cache/cache_reg[7][52]  ( .D(n12422), .CK(clk), .RN(n6085), .Q(
        \I_cache/cache[7][52] ), .QN(n3489) );
  DFFRX1 \I_cache/cache_reg[3][53]  ( .D(n12418), .CK(clk), .RN(n6084), .Q(
        \I_cache/cache[3][53] ), .QN(n3397) );
  DFFRX1 \I_cache/cache_reg[4][53]  ( .D(n12417), .CK(clk), .RN(n6084), .Q(
        \I_cache/cache[4][53] ), .QN(n1708) );
  DFFRX1 \I_cache/cache_reg[5][53]  ( .D(n12416), .CK(clk), .RN(n6084), .Q(
        \I_cache/cache[5][53] ), .QN(n3396) );
  DFFRX1 \I_cache/cache_reg[6][53]  ( .D(n12415), .CK(clk), .RN(n6084), .Q(
        \I_cache/cache[6][53] ), .QN(n1799) );
  DFFRX1 \I_cache/cache_reg[7][53]  ( .D(n12414), .CK(clk), .RN(n6084), .Q(
        \I_cache/cache[7][53] ), .QN(n3487) );
  DFFRX1 \I_cache/cache_reg[3][54]  ( .D(n12410), .CK(clk), .RN(n6084), .Q(
        \I_cache/cache[3][54] ), .QN(n3394) );
  DFFRX1 \I_cache/cache_reg[4][54]  ( .D(n12409), .CK(clk), .RN(n6083), .Q(
        \I_cache/cache[4][54] ), .QN(n1705) );
  DFFRX1 \I_cache/cache_reg[5][54]  ( .D(n12408), .CK(clk), .RN(n6083), .Q(
        \I_cache/cache[5][54] ), .QN(n3393) );
  DFFRX1 \I_cache/cache_reg[6][54]  ( .D(n12407), .CK(clk), .RN(n6083), .Q(
        \I_cache/cache[6][54] ), .QN(n1797) );
  DFFRX1 \I_cache/cache_reg[7][54]  ( .D(n12406), .CK(clk), .RN(n6083), .Q(
        \I_cache/cache[7][54] ), .QN(n3485) );
  DFFRX1 \I_cache/cache_reg[3][55]  ( .D(n12402), .CK(clk), .RN(n6083), .Q(
        \I_cache/cache[3][55] ), .QN(n3391) );
  DFFRX1 \I_cache/cache_reg[4][55]  ( .D(n12401), .CK(clk), .RN(n6083), .Q(
        \I_cache/cache[4][55] ), .QN(n1702) );
  DFFRX1 \I_cache/cache_reg[5][55]  ( .D(n12400), .CK(clk), .RN(n6083), .Q(
        \I_cache/cache[5][55] ), .QN(n3390) );
  DFFRX1 \I_cache/cache_reg[6][55]  ( .D(n12399), .CK(clk), .RN(n6083), .Q(
        \I_cache/cache[6][55] ), .QN(n1795) );
  DFFRX1 \I_cache/cache_reg[7][55]  ( .D(n12398), .CK(clk), .RN(n6083), .Q(
        \I_cache/cache[7][55] ), .QN(n3483) );
  DFFRX1 \I_cache/cache_reg[3][56]  ( .D(n12394), .CK(clk), .RN(n6082), .Q(
        \I_cache/cache[3][56] ), .QN(n3388) );
  DFFRX1 \I_cache/cache_reg[4][56]  ( .D(n12393), .CK(clk), .RN(n6082), .Q(
        \I_cache/cache[4][56] ), .QN(n1699) );
  DFFRX1 \I_cache/cache_reg[5][56]  ( .D(n12392), .CK(clk), .RN(n6082), .Q(
        \I_cache/cache[5][56] ), .QN(n3387) );
  DFFRX1 \I_cache/cache_reg[6][56]  ( .D(n12391), .CK(clk), .RN(n6082), .Q(
        \I_cache/cache[6][56] ), .QN(n1793) );
  DFFRX1 \I_cache/cache_reg[7][56]  ( .D(n12390), .CK(clk), .RN(n6082), .Q(
        \I_cache/cache[7][56] ), .QN(n3481) );
  DFFRX1 \I_cache/cache_reg[3][57]  ( .D(n12386), .CK(clk), .RN(n6082), .Q(
        \I_cache/cache[3][57] ), .QN(n3385) );
  DFFRX1 \I_cache/cache_reg[4][57]  ( .D(n12385), .CK(clk), .RN(n6081), .Q(
        \I_cache/cache[4][57] ), .QN(n1696) );
  DFFRX1 \I_cache/cache_reg[5][57]  ( .D(n12384), .CK(clk), .RN(n6081), .Q(
        \I_cache/cache[5][57] ), .QN(n3384) );
  DFFRX1 \I_cache/cache_reg[6][57]  ( .D(n12383), .CK(clk), .RN(n6081), .Q(
        \I_cache/cache[6][57] ), .QN(n1792) );
  DFFRX1 \I_cache/cache_reg[7][57]  ( .D(n12382), .CK(clk), .RN(n6081), .Q(
        \I_cache/cache[7][57] ), .QN(n3480) );
  DFFRX1 \I_cache/cache_reg[3][58]  ( .D(n12378), .CK(clk), .RN(n6081), .Q(
        \I_cache/cache[3][58] ), .QN(n3472) );
  DFFRX1 \I_cache/cache_reg[4][58]  ( .D(n12377), .CK(clk), .RN(n6081), .Q(
        \I_cache/cache[4][58] ), .QN(n1783) );
  DFFRX1 \I_cache/cache_reg[5][58]  ( .D(n12376), .CK(clk), .RN(n6081), .Q(
        \I_cache/cache[5][58] ), .QN(n3471) );
  DFFRX1 \I_cache/cache_reg[6][58]  ( .D(n12375), .CK(clk), .RN(n6081), .Q(
        \I_cache/cache[6][58] ), .QN(n1846) );
  DFFRX1 \I_cache/cache_reg[7][58]  ( .D(n12374), .CK(clk), .RN(n6081), .Q(
        \I_cache/cache[7][58] ), .QN(n3534) );
  DFFRX1 \I_cache/cache_reg[3][59]  ( .D(n12370), .CK(clk), .RN(n6080), .Q(
        \I_cache/cache[3][59] ), .QN(n3469) );
  DFFRX1 \I_cache/cache_reg[4][59]  ( .D(n12369), .CK(clk), .RN(n6080), .Q(
        \I_cache/cache[4][59] ), .QN(n1780) );
  DFFRX1 \I_cache/cache_reg[5][59]  ( .D(n12368), .CK(clk), .RN(n6080), .Q(
        \I_cache/cache[5][59] ), .QN(n3468) );
  DFFRX1 \I_cache/cache_reg[6][59]  ( .D(n12367), .CK(clk), .RN(n6080), .Q(
        \I_cache/cache[6][59] ), .QN(n1844) );
  DFFRX1 \I_cache/cache_reg[7][59]  ( .D(n12366), .CK(clk), .RN(n6080), .Q(
        \I_cache/cache[7][59] ), .QN(n3532) );
  DFFRX1 \I_cache/cache_reg[3][60]  ( .D(n12362), .CK(clk), .RN(n6080), .Q(
        \I_cache/cache[3][60] ), .QN(n3466) );
  DFFRX1 \I_cache/cache_reg[4][60]  ( .D(n12361), .CK(clk), .RN(n6079), .Q(
        \I_cache/cache[4][60] ), .QN(n1777) );
  DFFRX1 \I_cache/cache_reg[5][60]  ( .D(n12360), .CK(clk), .RN(n6079), .Q(
        \I_cache/cache[5][60] ), .QN(n3465) );
  DFFRX1 \I_cache/cache_reg[6][60]  ( .D(n12359), .CK(clk), .RN(n6079), .Q(
        \I_cache/cache[6][60] ), .QN(n1842) );
  DFFRX1 \I_cache/cache_reg[7][60]  ( .D(n12358), .CK(clk), .RN(n6079), .Q(
        \I_cache/cache[7][60] ), .QN(n3530) );
  DFFRX1 \I_cache/cache_reg[3][61]  ( .D(n12354), .CK(clk), .RN(n6079), .Q(
        \I_cache/cache[3][61] ), .QN(n3463) );
  DFFRX1 \I_cache/cache_reg[4][61]  ( .D(n12353), .CK(clk), .RN(n6079), .Q(
        \I_cache/cache[4][61] ), .QN(n1774) );
  DFFRX1 \I_cache/cache_reg[5][61]  ( .D(n12352), .CK(clk), .RN(n6079), .Q(
        \I_cache/cache[5][61] ), .QN(n3462) );
  DFFRX1 \I_cache/cache_reg[6][61]  ( .D(n12351), .CK(clk), .RN(n6079), .Q(
        \I_cache/cache[6][61] ), .QN(n1840) );
  DFFRX1 \I_cache/cache_reg[7][61]  ( .D(n12350), .CK(clk), .RN(n6079), .Q(
        \I_cache/cache[7][61] ), .QN(n3528) );
  DFFRX1 \I_cache/cache_reg[3][62]  ( .D(n12346), .CK(clk), .RN(n6078), .Q(
        \I_cache/cache[3][62] ), .QN(n3460) );
  DFFRX1 \I_cache/cache_reg[4][62]  ( .D(n12345), .CK(clk), .RN(n6078), .Q(
        \I_cache/cache[4][62] ), .QN(n1771) );
  DFFRX1 \I_cache/cache_reg[5][62]  ( .D(n12344), .CK(clk), .RN(n6078), .Q(
        \I_cache/cache[5][62] ), .QN(n3459) );
  DFFRX1 \I_cache/cache_reg[6][62]  ( .D(n12343), .CK(clk), .RN(n6078), .Q(
        \I_cache/cache[6][62] ), .QN(n1838) );
  DFFRX1 \I_cache/cache_reg[7][62]  ( .D(n12342), .CK(clk), .RN(n6078), .Q(
        \I_cache/cache[7][62] ), .QN(n3526) );
  DFFRX1 \I_cache/cache_reg[3][63]  ( .D(n12338), .CK(clk), .RN(n6078), .Q(
        \I_cache/cache[3][63] ), .QN(n3457) );
  DFFRX1 \I_cache/cache_reg[4][63]  ( .D(n12337), .CK(clk), .RN(n6077), .Q(
        \I_cache/cache[4][63] ), .QN(n1768) );
  DFFRX1 \I_cache/cache_reg[5][63]  ( .D(n12336), .CK(clk), .RN(n6077), .Q(
        \I_cache/cache[5][63] ), .QN(n3456) );
  DFFRX1 \I_cache/cache_reg[6][63]  ( .D(n12335), .CK(clk), .RN(n6077), .Q(
        \I_cache/cache[6][63] ), .QN(n1836) );
  DFFRX1 \I_cache/cache_reg[7][63]  ( .D(n12334), .CK(clk), .RN(n6077), .Q(
        \I_cache/cache[7][63] ), .QN(n3524) );
  DFFRX1 \I_cache/cache_reg[3][64]  ( .D(n12330), .CK(clk), .RN(n6077), .Q(
        \I_cache/cache[3][64] ), .QN(n3291) );
  DFFRX1 \I_cache/cache_reg[4][64]  ( .D(n12329), .CK(clk), .RN(n6077), .Q(
        \I_cache/cache[4][64] ), .QN(n1602) );
  DFFRX1 \I_cache/cache_reg[5][64]  ( .D(n12328), .CK(clk), .RN(n6077), .Q(
        \I_cache/cache[5][64] ), .QN(n3290) );
  DFFRX1 \I_cache/cache_reg[6][64]  ( .D(n12327), .CK(clk), .RN(n6077), .Q(
        \I_cache/cache[6][64] ), .QN(n1789) );
  DFFRX1 \I_cache/cache_reg[7][64]  ( .D(n12326), .CK(clk), .RN(n6077), .Q(
        \I_cache/cache[7][64] ), .QN(n3477) );
  DFFRX1 \I_cache/cache_reg[3][65]  ( .D(n12322), .CK(clk), .RN(n6076), .Q(
        \I_cache/cache[3][65] ), .QN(n349) );
  DFFRX1 \I_cache/cache_reg[4][65]  ( .D(n12321), .CK(clk), .RN(n6076), .Q(
        \I_cache/cache[4][65] ), .QN(n1672) );
  DFFRX1 \I_cache/cache_reg[5][65]  ( .D(n12320), .CK(clk), .RN(n6076), .Q(
        \I_cache/cache[5][65] ), .QN(n3361) );
  DFFRX1 \I_cache/cache_reg[6][65]  ( .D(n12319), .CK(clk), .RN(n6076), .Q(
        \I_cache/cache[6][65] ), .QN(n1788) );
  DFFRX1 \I_cache/cache_reg[7][65]  ( .D(n12318), .CK(clk), .RN(n6076), .Q(
        \I_cache/cache[7][65] ), .QN(n3476) );
  DFFRX1 \I_cache/cache_reg[3][66]  ( .D(n12314), .CK(clk), .RN(n6076), .Q(
        \I_cache/cache[3][66] ), .QN(n3360) );
  DFFRX1 \I_cache/cache_reg[4][66]  ( .D(n12313), .CK(clk), .RN(n6075), .Q(
        \I_cache/cache[4][66] ), .QN(n1670) );
  DFFRX1 \I_cache/cache_reg[5][66]  ( .D(n12312), .CK(clk), .RN(n6075), .Q(
        \I_cache/cache[5][66] ), .QN(n3359) );
  DFFRX1 \I_cache/cache_reg[6][66]  ( .D(n12311), .CK(clk), .RN(n6075), .Q(
        \I_cache/cache[6][66] ), .QN(n1787) );
  DFFRX1 \I_cache/cache_reg[7][66]  ( .D(n12310), .CK(clk), .RN(n6075), .Q(
        \I_cache/cache[7][66] ), .QN(n3475) );
  DFFRX1 \I_cache/cache_reg[3][67]  ( .D(n12306), .CK(clk), .RN(n6075), .Q(
        \I_cache/cache[3][67] ), .QN(n3357) );
  DFFRX1 \I_cache/cache_reg[4][67]  ( .D(n12305), .CK(clk), .RN(n6075), .Q(
        \I_cache/cache[4][67] ), .QN(n1667) );
  DFFRX1 \I_cache/cache_reg[5][67]  ( .D(n12304), .CK(clk), .RN(n6075), .Q(
        \I_cache/cache[5][67] ), .QN(n3356) );
  DFFRX1 \I_cache/cache_reg[6][67]  ( .D(n12303), .CK(clk), .RN(n6075), .Q(
        \I_cache/cache[6][67] ), .QN(n1831) );
  DFFRX1 \I_cache/cache_reg[7][67]  ( .D(n12302), .CK(clk), .RN(n6075), .Q(
        \I_cache/cache[7][67] ), .QN(n3519) );
  DFFRX1 \I_cache/cache_reg[3][68]  ( .D(n12298), .CK(clk), .RN(n6074), .Q(
        \I_cache/cache[3][68] ), .QN(n3354) );
  DFFRX1 \I_cache/cache_reg[4][68]  ( .D(n12297), .CK(clk), .RN(n6074), .Q(
        \I_cache/cache[4][68] ), .QN(n1664) );
  DFFRX1 \I_cache/cache_reg[5][68]  ( .D(n12296), .CK(clk), .RN(n6074), .Q(
        \I_cache/cache[5][68] ), .QN(n3353) );
  DFFRX1 \I_cache/cache_reg[6][68]  ( .D(n12295), .CK(clk), .RN(n6074), .Q(
        \I_cache/cache[6][68] ), .QN(n1786) );
  DFFRX1 \I_cache/cache_reg[7][68]  ( .D(n12294), .CK(clk), .RN(n6074), .Q(
        \I_cache/cache[7][68] ), .QN(n3474) );
  DFFRX1 \I_cache/cache_reg[3][69]  ( .D(n12290), .CK(clk), .RN(n6074), .Q(
        \I_cache/cache[3][69] ), .QN(n3351) );
  DFFRX1 \I_cache/cache_reg[4][69]  ( .D(n12289), .CK(clk), .RN(n6073), .Q(
        \I_cache/cache[4][69] ), .QN(n1661) );
  DFFRX1 \I_cache/cache_reg[5][69]  ( .D(n12288), .CK(clk), .RN(n6073), .Q(
        \I_cache/cache[5][69] ), .QN(n3350) );
  DFFRX1 \I_cache/cache_reg[6][69]  ( .D(n12287), .CK(clk), .RN(n6073), .Q(
        \I_cache/cache[6][69] ), .QN(n1828) );
  DFFRX1 \I_cache/cache_reg[7][69]  ( .D(n12286), .CK(clk), .RN(n6073), .Q(
        \I_cache/cache[7][69] ), .QN(n3516) );
  DFFRX1 \I_cache/cache_reg[3][70]  ( .D(n12282), .CK(clk), .RN(n6073), .Q(
        \I_cache/cache[3][70] ), .QN(n3348) );
  DFFRX1 \I_cache/cache_reg[4][70]  ( .D(n12281), .CK(clk), .RN(n6073), .Q(
        \I_cache/cache[4][70] ), .QN(n1658) );
  DFFRX1 \I_cache/cache_reg[5][70]  ( .D(n12280), .CK(clk), .RN(n6073), .Q(
        \I_cache/cache[5][70] ), .QN(n3347) );
  DFFRX1 \I_cache/cache_reg[6][70]  ( .D(n12279), .CK(clk), .RN(n6073), .Q(
        \I_cache/cache[6][70] ), .QN(n1826) );
  DFFRX1 \I_cache/cache_reg[7][70]  ( .D(n12278), .CK(clk), .RN(n6073), .Q(
        \I_cache/cache[7][70] ), .QN(n3514) );
  DFFRX1 \I_cache/cache_reg[3][71]  ( .D(n12274), .CK(clk), .RN(n6072), .Q(
        \I_cache/cache[3][71] ), .QN(n3345) );
  DFFRX1 \I_cache/cache_reg[4][71]  ( .D(n12273), .CK(clk), .RN(n6072), .Q(
        \I_cache/cache[4][71] ), .QN(n1655) );
  DFFRX1 \I_cache/cache_reg[5][71]  ( .D(n12272), .CK(clk), .RN(n6072), .Q(
        \I_cache/cache[5][71] ), .QN(n3344) );
  DFFRX1 \I_cache/cache_reg[6][71]  ( .D(n12271), .CK(clk), .RN(n6072), .Q(
        \I_cache/cache[6][71] ), .QN(n1824) );
  DFFRX1 \I_cache/cache_reg[7][71]  ( .D(n12270), .CK(clk), .RN(n6072), .Q(
        \I_cache/cache[7][71] ), .QN(n3512) );
  DFFRX1 \I_cache/cache_reg[3][72]  ( .D(n12266), .CK(clk), .RN(n6072), .Q(
        \I_cache/cache[3][72] ), .QN(n3342) );
  DFFRX1 \I_cache/cache_reg[5][72]  ( .D(n12264), .CK(clk), .RN(n6071), .Q(
        \I_cache/cache[5][72] ), .QN(n3341) );
  DFFRX1 \I_cache/cache_reg[6][72]  ( .D(n12263), .CK(clk), .RN(n6071), .Q(
        \I_cache/cache[6][72] ), .QN(n1822) );
  DFFRX1 \I_cache/cache_reg[7][72]  ( .D(n12262), .CK(clk), .RN(n6071), .Q(
        \I_cache/cache[7][72] ), .QN(n3510) );
  DFFRX1 \I_cache/cache_reg[3][73]  ( .D(n12258), .CK(clk), .RN(n6071), .Q(
        \I_cache/cache[3][73] ), .QN(n3339) );
  DFFRX1 \I_cache/cache_reg[4][73]  ( .D(n12257), .CK(clk), .RN(n6071), .Q(
        \I_cache/cache[4][73] ), .QN(n1649) );
  DFFRX1 \I_cache/cache_reg[5][73]  ( .D(n12256), .CK(clk), .RN(n6071), .Q(
        \I_cache/cache[5][73] ), .QN(n3338) );
  DFFRX1 \I_cache/cache_reg[6][73]  ( .D(n12255), .CK(clk), .RN(n6071), .Q(
        \I_cache/cache[6][73] ), .QN(n1820) );
  DFFRX1 \I_cache/cache_reg[7][73]  ( .D(n12254), .CK(clk), .RN(n6071), .Q(
        \I_cache/cache[7][73] ), .QN(n3508) );
  DFFRX1 \I_cache/cache_reg[3][74]  ( .D(n12250), .CK(clk), .RN(n6070), .Q(
        \I_cache/cache[3][74] ), .QN(n3336) );
  DFFRX1 \I_cache/cache_reg[4][74]  ( .D(n12249), .CK(clk), .RN(n6070), .Q(
        \I_cache/cache[4][74] ), .QN(n1646) );
  DFFRX1 \I_cache/cache_reg[5][74]  ( .D(n12248), .CK(clk), .RN(n6070), .Q(
        \I_cache/cache[5][74] ), .QN(n3335) );
  DFFRX1 \I_cache/cache_reg[6][74]  ( .D(n12247), .CK(clk), .RN(n6070), .Q(
        \I_cache/cache[6][74] ), .QN(n1818) );
  DFFRX1 \I_cache/cache_reg[7][74]  ( .D(n12246), .CK(clk), .RN(n6070), .Q(
        \I_cache/cache[7][74] ), .QN(n3506) );
  DFFRX1 \I_cache/cache_reg[3][75]  ( .D(n12242), .CK(clk), .RN(n6070), .Q(
        \I_cache/cache[3][75] ), .QN(n3333) );
  DFFRX1 \I_cache/cache_reg[4][75]  ( .D(n12241), .CK(clk), .RN(n6069), .Q(
        \I_cache/cache[4][75] ), .QN(n1643) );
  DFFRX1 \I_cache/cache_reg[5][75]  ( .D(n12240), .CK(clk), .RN(n6069), .Q(
        \I_cache/cache[5][75] ), .QN(n3332) );
  DFFRX1 \I_cache/cache_reg[6][75]  ( .D(n12239), .CK(clk), .RN(n6069), .Q(
        \I_cache/cache[6][75] ), .QN(n1816) );
  DFFRX1 \I_cache/cache_reg[7][75]  ( .D(n12238), .CK(clk), .RN(n6069), .Q(
        \I_cache/cache[7][75] ), .QN(n3504) );
  DFFRX1 \I_cache/cache_reg[3][76]  ( .D(n12234), .CK(clk), .RN(n6069), .Q(
        \I_cache/cache[3][76] ), .QN(n3330) );
  DFFRX1 \I_cache/cache_reg[4][76]  ( .D(n12233), .CK(clk), .RN(n6069), .Q(
        \I_cache/cache[4][76] ), .QN(n1640) );
  DFFRX1 \I_cache/cache_reg[5][76]  ( .D(n12232), .CK(clk), .RN(n6069), .Q(
        \I_cache/cache[5][76] ), .QN(n3329) );
  DFFRX1 \I_cache/cache_reg[6][76]  ( .D(n12231), .CK(clk), .RN(n6069), .Q(
        \I_cache/cache[6][76] ), .QN(n1814) );
  DFFRX1 \I_cache/cache_reg[7][76]  ( .D(n12230), .CK(clk), .RN(n6069), .Q(
        \I_cache/cache[7][76] ), .QN(n3502) );
  DFFRX1 \I_cache/cache_reg[3][77]  ( .D(n12226), .CK(clk), .RN(n6068), .Q(
        \I_cache/cache[3][77] ), .QN(n3327) );
  DFFRX1 \I_cache/cache_reg[4][77]  ( .D(n12225), .CK(clk), .RN(n6068), .Q(
        \I_cache/cache[4][77] ), .QN(n1637) );
  DFFRX1 \I_cache/cache_reg[5][77]  ( .D(n12224), .CK(clk), .RN(n6068), .Q(
        \I_cache/cache[5][77] ), .QN(n3326) );
  DFFRX1 \I_cache/cache_reg[6][77]  ( .D(n12223), .CK(clk), .RN(n6068), .Q(
        \I_cache/cache[6][77] ), .QN(n1812) );
  DFFRX1 \I_cache/cache_reg[7][77]  ( .D(n12222), .CK(clk), .RN(n6068), .Q(
        \I_cache/cache[7][77] ), .QN(n3500) );
  DFFRX1 \I_cache/cache_reg[3][78]  ( .D(n12218), .CK(clk), .RN(n6068), .Q(
        \I_cache/cache[3][78] ), .QN(n3324) );
  DFFRX1 \I_cache/cache_reg[4][78]  ( .D(n12217), .CK(clk), .RN(n6067), .Q(
        \I_cache/cache[4][78] ), .QN(n1634) );
  DFFRX1 \I_cache/cache_reg[5][78]  ( .D(n12216), .CK(clk), .RN(n6067), .Q(
        \I_cache/cache[5][78] ), .QN(n3323) );
  DFFRX1 \I_cache/cache_reg[6][78]  ( .D(n12215), .CK(clk), .RN(n6067), .Q(
        \I_cache/cache[6][78] ), .QN(n1810) );
  DFFRX1 \I_cache/cache_reg[7][78]  ( .D(n12214), .CK(clk), .RN(n6067), .Q(
        \I_cache/cache[7][78] ), .QN(n3498) );
  DFFRX1 \I_cache/cache_reg[3][79]  ( .D(n12210), .CK(clk), .RN(n6067), .Q(
        \I_cache/cache[3][79] ), .QN(n3321) );
  DFFRX1 \I_cache/cache_reg[4][79]  ( .D(n12209), .CK(clk), .RN(n6067), .Q(
        \I_cache/cache[4][79] ), .QN(n1631) );
  DFFRX1 \I_cache/cache_reg[5][79]  ( .D(n12208), .CK(clk), .RN(n6067), .Q(
        \I_cache/cache[5][79] ), .QN(n3320) );
  DFFRX1 \I_cache/cache_reg[6][79]  ( .D(n12207), .CK(clk), .RN(n6067), .Q(
        \I_cache/cache[6][79] ), .QN(n1808) );
  DFFRX1 \I_cache/cache_reg[7][79]  ( .D(n12206), .CK(clk), .RN(n6067), .Q(
        \I_cache/cache[7][79] ), .QN(n3496) );
  DFFRX1 \I_cache/cache_reg[3][80]  ( .D(n12202), .CK(clk), .RN(n6066), .Q(
        \I_cache/cache[3][80] ), .QN(n3318) );
  DFFRX1 \I_cache/cache_reg[4][80]  ( .D(n12201), .CK(clk), .RN(n6066), .Q(
        \I_cache/cache[4][80] ), .QN(n1628) );
  DFFRX1 \I_cache/cache_reg[5][80]  ( .D(n12200), .CK(clk), .RN(n6066), .Q(
        \I_cache/cache[5][80] ), .QN(n3317) );
  DFFRX1 \I_cache/cache_reg[6][80]  ( .D(n12199), .CK(clk), .RN(n6066), .Q(
        \I_cache/cache[6][80] ), .QN(n1806) );
  DFFRX1 \I_cache/cache_reg[7][80]  ( .D(n12198), .CK(clk), .RN(n6066), .Q(
        \I_cache/cache[7][80] ), .QN(n3494) );
  DFFRX1 \I_cache/cache_reg[3][81]  ( .D(n12194), .CK(clk), .RN(n6066), .Q(
        \I_cache/cache[3][81] ), .QN(n3315) );
  DFFRX1 \I_cache/cache_reg[4][81]  ( .D(n12193), .CK(clk), .RN(n6065), .Q(
        \I_cache/cache[4][81] ), .QN(n1626) );
  DFFRX1 \I_cache/cache_reg[5][81]  ( .D(n12192), .CK(clk), .RN(n6065), .Q(
        \I_cache/cache[5][81] ), .QN(n3314) );
  DFFRX1 \I_cache/cache_reg[6][81]  ( .D(n12191), .CK(clk), .RN(n6065), .Q(
        \I_cache/cache[6][81] ), .QN(n1804) );
  DFFRX1 \I_cache/cache_reg[7][81]  ( .D(n12190), .CK(clk), .RN(n6065), .Q(
        \I_cache/cache[7][81] ), .QN(n3492) );
  DFFRX1 \I_cache/cache_reg[3][82]  ( .D(n12186), .CK(clk), .RN(n6065), .Q(
        \I_cache/cache[3][82] ), .QN(n3312) );
  DFFRX1 \I_cache/cache_reg[4][82]  ( .D(n12185), .CK(clk), .RN(n6065), .Q(
        \I_cache/cache[4][82] ), .QN(n1623) );
  DFFRX1 \I_cache/cache_reg[5][82]  ( .D(n12184), .CK(clk), .RN(n6065), .Q(
        \I_cache/cache[5][82] ), .QN(n3311) );
  DFFRX1 \I_cache/cache_reg[6][82]  ( .D(n12183), .CK(clk), .RN(n6065), .Q(
        \I_cache/cache[6][82] ), .QN(n1802) );
  DFFRX1 \I_cache/cache_reg[7][82]  ( .D(n12182), .CK(clk), .RN(n6065), .Q(
        \I_cache/cache[7][82] ), .QN(n3490) );
  DFFRX1 \I_cache/cache_reg[3][83]  ( .D(n12178), .CK(clk), .RN(n6064), .Q(
        \I_cache/cache[3][83] ), .QN(n3537) );
  DFFRX1 \I_cache/cache_reg[4][83]  ( .D(n12177), .CK(clk), .RN(n6064), .Q(
        \I_cache/cache[4][83] ), .QN(n1848) );
  DFFRX1 \I_cache/cache_reg[5][83]  ( .D(n12176), .CK(clk), .RN(n6064), .Q(
        \I_cache/cache[5][83] ), .QN(n3536) );
  DFFRX1 \I_cache/cache_reg[6][83]  ( .D(n12175), .CK(clk), .RN(n6064), .Q(
        \I_cache/cache[6][83] ), .QN(n1854) );
  DFFRX1 \I_cache/cache_reg[7][83]  ( .D(n12174), .CK(clk), .RN(n6064), .Q(
        \I_cache/cache[7][83] ), .QN(n3541) );
  DFFRX1 \I_cache/cache_reg[3][84]  ( .D(n12170), .CK(clk), .RN(n6064), .Q(
        \I_cache/cache[3][84] ), .QN(n3309) );
  DFFRX1 \I_cache/cache_reg[4][84]  ( .D(n12169), .CK(clk), .RN(n6063), .Q(
        \I_cache/cache[4][84] ), .QN(n1620) );
  DFFRX1 \I_cache/cache_reg[5][84]  ( .D(n12168), .CK(clk), .RN(n6063), .Q(
        \I_cache/cache[5][84] ), .QN(n3308) );
  DFFRX1 \I_cache/cache_reg[6][84]  ( .D(n12167), .CK(clk), .RN(n6063), .Q(
        \I_cache/cache[6][84] ), .QN(n1800) );
  DFFRX1 \I_cache/cache_reg[7][84]  ( .D(n12166), .CK(clk), .RN(n6063), .Q(
        \I_cache/cache[7][84] ), .QN(n3488) );
  DFFRX1 \I_cache/cache_reg[3][85]  ( .D(n12162), .CK(clk), .RN(n6063), .Q(
        \I_cache/cache[3][85] ), .QN(n3306) );
  DFFRX1 \I_cache/cache_reg[4][85]  ( .D(n12161), .CK(clk), .RN(n6063), .Q(
        \I_cache/cache[4][85] ), .QN(n1617) );
  DFFRX1 \I_cache/cache_reg[5][85]  ( .D(n12160), .CK(clk), .RN(n6063), .Q(
        \I_cache/cache[5][85] ), .QN(n3305) );
  DFFRX1 \I_cache/cache_reg[6][85]  ( .D(n12159), .CK(clk), .RN(n6063), .Q(
        \I_cache/cache[6][85] ), .QN(n1798) );
  DFFRX1 \I_cache/cache_reg[7][85]  ( .D(n12158), .CK(clk), .RN(n6063), .Q(
        \I_cache/cache[7][85] ), .QN(n3486) );
  DFFRX1 \I_cache/cache_reg[3][86]  ( .D(n12154), .CK(clk), .RN(n6062), .Q(
        \I_cache/cache[3][86] ), .QN(n3303) );
  DFFRX1 \I_cache/cache_reg[4][86]  ( .D(n12153), .CK(clk), .RN(n6062), .Q(
        \I_cache/cache[4][86] ), .QN(n1614) );
  DFFRX1 \I_cache/cache_reg[5][86]  ( .D(n12152), .CK(clk), .RN(n6062), .Q(
        \I_cache/cache[5][86] ), .QN(n3302) );
  DFFRX1 \I_cache/cache_reg[6][86]  ( .D(n12151), .CK(clk), .RN(n6062), .Q(
        \I_cache/cache[6][86] ), .QN(n1796) );
  DFFRX1 \I_cache/cache_reg[7][86]  ( .D(n12150), .CK(clk), .RN(n6062), .Q(
        \I_cache/cache[7][86] ), .QN(n3484) );
  DFFRX1 \I_cache/cache_reg[3][87]  ( .D(n12146), .CK(clk), .RN(n6062), .Q(
        \I_cache/cache[3][87] ), .QN(n3300) );
  DFFRX1 \I_cache/cache_reg[4][87]  ( .D(n12145), .CK(clk), .RN(n6061), .Q(
        \I_cache/cache[4][87] ), .QN(n1611) );
  DFFRX1 \I_cache/cache_reg[5][87]  ( .D(n12144), .CK(clk), .RN(n6061), .Q(
        \I_cache/cache[5][87] ), .QN(n3299) );
  DFFRX1 \I_cache/cache_reg[6][87]  ( .D(n12143), .CK(clk), .RN(n6061), .Q(
        \I_cache/cache[6][87] ), .QN(n1794) );
  DFFRX1 \I_cache/cache_reg[7][87]  ( .D(n12142), .CK(clk), .RN(n6061), .Q(
        \I_cache/cache[7][87] ), .QN(n3482) );
  DFFRX1 \I_cache/cache_reg[3][88]  ( .D(n12138), .CK(clk), .RN(n6061), .Q(
        \I_cache/cache[3][88] ), .QN(n3297) );
  DFFRX1 \I_cache/cache_reg[4][88]  ( .D(n12137), .CK(clk), .RN(n6061), .Q(
        \I_cache/cache[4][88] ), .QN(n1608) );
  DFFRX1 \I_cache/cache_reg[5][88]  ( .D(n12136), .CK(clk), .RN(n6061), .Q(
        \I_cache/cache[5][88] ), .QN(n3296) );
  DFFRX1 \I_cache/cache_reg[6][88]  ( .D(n12135), .CK(clk), .RN(n6061), .Q(
        \I_cache/cache[6][88] ), .QN(n1785) );
  DFFRX1 \I_cache/cache_reg[7][88]  ( .D(n12134), .CK(clk), .RN(n6061), .Q(
        \I_cache/cache[7][88] ), .QN(n3473) );
  DFFRX1 \I_cache/cache_reg[3][89]  ( .D(n12130), .CK(clk), .RN(n6060), .Q(
        \I_cache/cache[3][89] ), .QN(n3294) );
  DFFRX1 \I_cache/cache_reg[4][89]  ( .D(n12129), .CK(clk), .RN(n6060), .Q(
        \I_cache/cache[4][89] ), .QN(n1605) );
  DFFRX1 \I_cache/cache_reg[5][89]  ( .D(n12128), .CK(clk), .RN(n6060), .Q(
        \I_cache/cache[5][89] ), .QN(n3293) );
  DFFRX1 \I_cache/cache_reg[6][89]  ( .D(n12127), .CK(clk), .RN(n6060), .Q(
        \I_cache/cache[6][89] ), .QN(n1791) );
  DFFRX1 \I_cache/cache_reg[7][89]  ( .D(n12126), .CK(clk), .RN(n6060), .Q(
        \I_cache/cache[7][89] ), .QN(n3479) );
  DFFRX1 \I_cache/cache_reg[3][90]  ( .D(n12122), .CK(clk), .RN(n6060), .Q(
        \I_cache/cache[3][90] ), .QN(n3379) );
  DFFRX1 \I_cache/cache_reg[4][90]  ( .D(n12121), .CK(clk), .RN(n6059), .Q(
        \I_cache/cache[4][90] ), .QN(n1690) );
  DFFRX1 \I_cache/cache_reg[5][90]  ( .D(n12120), .CK(clk), .RN(n6059), .Q(
        \I_cache/cache[5][90] ), .QN(n3378) );
  DFFRX1 \I_cache/cache_reg[6][90]  ( .D(n12119), .CK(clk), .RN(n6059), .Q(
        \I_cache/cache[6][90] ), .QN(n1845) );
  DFFRX1 \I_cache/cache_reg[7][90]  ( .D(n12118), .CK(clk), .RN(n6059), .Q(
        \I_cache/cache[7][90] ), .QN(n3533) );
  DFFRX1 \I_cache/cache_reg[3][91]  ( .D(n12114), .CK(clk), .RN(n6059), .Q(
        \I_cache/cache[3][91] ), .QN(n3376) );
  DFFRX1 \I_cache/cache_reg[4][91]  ( .D(n12113), .CK(clk), .RN(n6059), .Q(
        \I_cache/cache[4][91] ), .QN(n1687) );
  DFFRX1 \I_cache/cache_reg[5][91]  ( .D(n12112), .CK(clk), .RN(n6059), .Q(
        \I_cache/cache[5][91] ), .QN(n3375) );
  DFFRX1 \I_cache/cache_reg[6][91]  ( .D(n12111), .CK(clk), .RN(n6059), .Q(
        \I_cache/cache[6][91] ), .QN(n1843) );
  DFFRX1 \I_cache/cache_reg[7][91]  ( .D(n12110), .CK(clk), .RN(n6059), .Q(
        \I_cache/cache[7][91] ), .QN(n3531) );
  DFFRX1 \I_cache/cache_reg[3][92]  ( .D(n12106), .CK(clk), .RN(n6058), .Q(
        \I_cache/cache[3][92] ), .QN(n3373) );
  DFFRX1 \I_cache/cache_reg[4][92]  ( .D(n12105), .CK(clk), .RN(n6058), .Q(
        \I_cache/cache[4][92] ), .QN(n1684) );
  DFFRX1 \I_cache/cache_reg[5][92]  ( .D(n12104), .CK(clk), .RN(n6058), .Q(
        \I_cache/cache[5][92] ), .QN(n3372) );
  DFFRX1 \I_cache/cache_reg[6][92]  ( .D(n12103), .CK(clk), .RN(n6058), .Q(
        \I_cache/cache[6][92] ), .QN(n1841) );
  DFFRX1 \I_cache/cache_reg[7][92]  ( .D(n12102), .CK(clk), .RN(n6058), .Q(
        \I_cache/cache[7][92] ), .QN(n3529) );
  DFFRX1 \I_cache/cache_reg[3][93]  ( .D(n12098), .CK(clk), .RN(n6058), .Q(
        \I_cache/cache[3][93] ), .QN(n3370) );
  DFFRX1 \I_cache/cache_reg[4][93]  ( .D(n12097), .CK(clk), .RN(n6057), .Q(
        \I_cache/cache[4][93] ), .QN(n1681) );
  DFFRX1 \I_cache/cache_reg[5][93]  ( .D(n12096), .CK(clk), .RN(n6057), .Q(
        \I_cache/cache[5][93] ), .QN(n3369) );
  DFFRX1 \I_cache/cache_reg[6][93]  ( .D(n12095), .CK(clk), .RN(n6057), .Q(
        \I_cache/cache[6][93] ), .QN(n1839) );
  DFFRX1 \I_cache/cache_reg[7][93]  ( .D(n12094), .CK(clk), .RN(n6057), .Q(
        \I_cache/cache[7][93] ), .QN(n3527) );
  DFFRX1 \I_cache/cache_reg[3][94]  ( .D(n12090), .CK(clk), .RN(n6057), .Q(
        \I_cache/cache[3][94] ), .QN(n3367) );
  DFFRX1 \I_cache/cache_reg[4][94]  ( .D(n12089), .CK(clk), .RN(n6057), .Q(
        \I_cache/cache[4][94] ), .QN(n1678) );
  DFFRX1 \I_cache/cache_reg[5][94]  ( .D(n12088), .CK(clk), .RN(n6057), .Q(
        \I_cache/cache[5][94] ), .QN(n3366) );
  DFFRX1 \I_cache/cache_reg[6][94]  ( .D(n12087), .CK(clk), .RN(n6057), .Q(
        \I_cache/cache[6][94] ), .QN(n1837) );
  DFFRX1 \I_cache/cache_reg[7][94]  ( .D(n12086), .CK(clk), .RN(n6057), .Q(
        \I_cache/cache[7][94] ), .QN(n3525) );
  DFFRX1 \I_cache/cache_reg[3][95]  ( .D(n12082), .CK(clk), .RN(n6056), .Q(
        \I_cache/cache[3][95] ), .QN(n3364) );
  DFFRX1 \I_cache/cache_reg[4][95]  ( .D(n12081), .CK(clk), .RN(n6056), .Q(
        \I_cache/cache[4][95] ), .QN(n1675) );
  DFFRX1 \I_cache/cache_reg[5][95]  ( .D(n12080), .CK(clk), .RN(n6056), .Q(
        \I_cache/cache[5][95] ), .QN(n3363) );
  DFFRX1 \I_cache/cache_reg[6][95]  ( .D(n12079), .CK(clk), .RN(n6056), .Q(
        \I_cache/cache[6][95] ), .QN(n1835) );
  DFFRX1 \I_cache/cache_reg[7][95]  ( .D(n12078), .CK(clk), .RN(n6056), .Q(
        \I_cache/cache[7][95] ), .QN(n3523) );
  DFFRX1 \I_cache/cache_reg[3][96]  ( .D(n12074), .CK(clk), .RN(n6056), .Q(
        \I_cache/cache[3][96] ), .QN(n3036) );
  DFFRX1 \I_cache/cache_reg[4][96]  ( .D(n12073), .CK(clk), .RN(n6055), .Q(
        \I_cache/cache[4][96] ), .QN(n1348) );
  DFFRX1 \I_cache/cache_reg[5][96]  ( .D(n12072), .CK(clk), .RN(n6055), .Q(
        \I_cache/cache[5][96] ), .QN(n3035) );
  DFFRX1 \I_cache/cache_reg[6][96]  ( .D(n12071), .CK(clk), .RN(n6055), .Q(
        \I_cache/cache[6][96] ), .QN(n1529) );
  DFFRX1 \I_cache/cache_reg[7][96]  ( .D(n12070), .CK(clk), .RN(n6055), .Q(
        \I_cache/cache[7][96] ), .QN(n3216) );
  DFFRX1 \I_cache/cache_reg[3][97]  ( .D(n12066), .CK(clk), .RN(n6055), .Q(
        \I_cache/cache[3][97] ), .QN(n3107) );
  DFFRX1 \I_cache/cache_reg[4][97]  ( .D(n12065), .CK(clk), .RN(n6055), .Q(
        \I_cache/cache[4][97] ), .QN(n1419) );
  DFFRX1 \I_cache/cache_reg[5][97]  ( .D(n12064), .CK(clk), .RN(n6055), .Q(
        \I_cache/cache[5][97] ), .QN(n3106) );
  DFFRX1 \I_cache/cache_reg[6][97]  ( .D(n12063), .CK(clk), .RN(n6055), .Q(
        \I_cache/cache[6][97] ), .QN(n1576) );
  DFFRX1 \I_cache/cache_reg[7][97]  ( .D(n12062), .CK(clk), .RN(n6055), .Q(
        \I_cache/cache[7][97] ), .QN(n3288) );
  DFFRX1 \I_cache/cache_reg[3][98]  ( .D(n12058), .CK(clk), .RN(n6054), .Q(
        \I_cache/cache[3][98] ), .QN(n3104) );
  DFFRX1 \I_cache/cache_reg[4][98]  ( .D(n12057), .CK(clk), .RN(n6054), .Q(
        \I_cache/cache[4][98] ), .QN(n1416) );
  DFFRX1 \I_cache/cache_reg[5][98]  ( .D(n12056), .CK(clk), .RN(n6054), .Q(
        \I_cache/cache[5][98] ), .QN(n3103) );
  DFFRX1 \I_cache/cache_reg[6][98]  ( .D(n12055), .CK(clk), .RN(n6054), .Q(
        \I_cache/cache[6][98] ), .QN(n1574) );
  DFFRX1 \I_cache/cache_reg[7][98]  ( .D(n12054), .CK(clk), .RN(n6054), .Q(
        \I_cache/cache[7][98] ), .QN(n3262) );
  DFFRX1 \I_cache/cache_reg[3][99]  ( .D(n12050), .CK(clk), .RN(n6054), .Q(
        \I_cache/cache[3][99] ), .QN(n3101) );
  DFFRX1 \I_cache/cache_reg[4][99]  ( .D(n12049), .CK(clk), .RN(n6053), .Q(
        \I_cache/cache[4][99] ), .QN(n1413) );
  DFFRX1 \I_cache/cache_reg[5][99]  ( .D(n12048), .CK(clk), .RN(n6053), .Q(
        \I_cache/cache[5][99] ), .QN(n3100) );
  DFFRX1 \I_cache/cache_reg[6][99]  ( .D(n12047), .CK(clk), .RN(n6053), .Q(
        \I_cache/cache[6][99] ), .QN(n1572) );
  DFFRX1 \I_cache/cache_reg[7][99]  ( .D(n12046), .CK(clk), .RN(n6053), .Q(
        \I_cache/cache[7][99] ), .QN(n3260) );
  DFFRX1 \I_cache/cache_reg[3][100]  ( .D(n12042), .CK(clk), .RN(n6053), .Q(
        \I_cache/cache[3][100] ), .QN(n3098) );
  DFFRX1 \I_cache/cache_reg[4][100]  ( .D(n12041), .CK(clk), .RN(n6053), .Q(
        \I_cache/cache[4][100] ), .QN(n1410) );
  DFFRX1 \I_cache/cache_reg[5][100]  ( .D(n12040), .CK(clk), .RN(n6053), .Q(
        \I_cache/cache[5][100] ), .QN(n3097) );
  DFFRX1 \I_cache/cache_reg[6][100]  ( .D(n12039), .CK(clk), .RN(n6053), .Q(
        \I_cache/cache[6][100] ), .QN(n1570) );
  DFFRX1 \I_cache/cache_reg[7][100]  ( .D(n12038), .CK(clk), .RN(n6053), .Q(
        \I_cache/cache[7][100] ), .QN(n3258) );
  DFFRX1 \I_cache/cache_reg[3][101]  ( .D(n12034), .CK(clk), .RN(n6052), .Q(
        \I_cache/cache[3][101] ), .QN(n3095) );
  DFFRX1 \I_cache/cache_reg[4][101]  ( .D(n12033), .CK(clk), .RN(n6052), .Q(
        \I_cache/cache[4][101] ), .QN(n1407) );
  DFFRX1 \I_cache/cache_reg[5][101]  ( .D(n12032), .CK(clk), .RN(n6052), .Q(
        \I_cache/cache[5][101] ), .QN(n3094) );
  DFFRX1 \I_cache/cache_reg[6][101]  ( .D(n12031), .CK(clk), .RN(n6052), .Q(
        \I_cache/cache[6][101] ), .QN(n1568) );
  DFFRX1 \I_cache/cache_reg[7][101]  ( .D(n12030), .CK(clk), .RN(n6052), .Q(
        \I_cache/cache[7][101] ), .QN(n3256) );
  DFFRX1 \I_cache/cache_reg[3][102]  ( .D(n12026), .CK(clk), .RN(n6052), .Q(
        \I_cache/cache[3][102] ), .QN(n3092) );
  DFFRX1 \I_cache/cache_reg[4][102]  ( .D(n12025), .CK(clk), .RN(n6051), .Q(
        \I_cache/cache[4][102] ), .QN(n1404) );
  DFFRX1 \I_cache/cache_reg[5][102]  ( .D(n12024), .CK(clk), .RN(n6051), .Q(
        \I_cache/cache[5][102] ), .QN(n3091) );
  DFFRX1 \I_cache/cache_reg[6][102]  ( .D(n12023), .CK(clk), .RN(n6051), .Q(
        \I_cache/cache[6][102] ), .QN(n1566) );
  DFFRX1 \I_cache/cache_reg[7][102]  ( .D(n12022), .CK(clk), .RN(n6051), .Q(
        \I_cache/cache[7][102] ), .QN(n3254) );
  DFFRX1 \I_cache/cache_reg[3][103]  ( .D(n12018), .CK(clk), .RN(n6051), .Q(
        \I_cache/cache[3][103] ), .QN(n3089) );
  DFFRX1 \I_cache/cache_reg[4][103]  ( .D(n12017), .CK(clk), .RN(n6051), .Q(
        \I_cache/cache[4][103] ), .QN(n1401) );
  DFFRX1 \I_cache/cache_reg[5][103]  ( .D(n12016), .CK(clk), .RN(n6051), .Q(
        \I_cache/cache[5][103] ), .QN(n3088) );
  DFFRX1 \I_cache/cache_reg[6][103]  ( .D(n12015), .CK(clk), .RN(n6051), .Q(
        \I_cache/cache[6][103] ), .QN(n1564) );
  DFFRX1 \I_cache/cache_reg[7][103]  ( .D(n12014), .CK(clk), .RN(n6051), .Q(
        \I_cache/cache[7][103] ), .QN(n3252) );
  DFFRX1 \I_cache/cache_reg[3][104]  ( .D(n12010), .CK(clk), .RN(n6050), .Q(
        \I_cache/cache[3][104] ), .QN(n3086) );
  DFFRX1 \I_cache/cache_reg[4][104]  ( .D(n12009), .CK(clk), .RN(n6050), .Q(
        \I_cache/cache[4][104] ), .QN(n1398) );
  DFFRX1 \I_cache/cache_reg[5][104]  ( .D(n12008), .CK(clk), .RN(n6050), .Q(
        \I_cache/cache[5][104] ), .QN(n3085) );
  DFFRX1 \I_cache/cache_reg[6][104]  ( .D(n12007), .CK(clk), .RN(n6050), .Q(
        \I_cache/cache[6][104] ), .QN(n1562) );
  DFFRX1 \I_cache/cache_reg[7][104]  ( .D(n12006), .CK(clk), .RN(n6050), .Q(
        \I_cache/cache[7][104] ), .QN(n3250) );
  DFFRX1 \I_cache/cache_reg[3][105]  ( .D(n12002), .CK(clk), .RN(n6050), .Q(
        \I_cache/cache[3][105] ), .QN(n3083) );
  DFFRX1 \I_cache/cache_reg[4][105]  ( .D(n12001), .CK(clk), .RN(n6049), .Q(
        \I_cache/cache[4][105] ), .QN(n1395) );
  DFFRX1 \I_cache/cache_reg[5][105]  ( .D(n12000), .CK(clk), .RN(n6049), .Q(
        \I_cache/cache[5][105] ), .QN(n3082) );
  DFFRX1 \I_cache/cache_reg[6][105]  ( .D(n11999), .CK(clk), .RN(n6049), .Q(
        \I_cache/cache[6][105] ), .QN(n1560) );
  DFFRX1 \I_cache/cache_reg[7][105]  ( .D(n11998), .CK(clk), .RN(n6049), .Q(
        \I_cache/cache[7][105] ), .QN(n3248) );
  DFFRX1 \I_cache/cache_reg[3][106]  ( .D(n11994), .CK(clk), .RN(n6049), .Q(
        \I_cache/cache[3][106] ), .QN(n3080) );
  DFFRX1 \I_cache/cache_reg[4][106]  ( .D(n11993), .CK(clk), .RN(n6049), .Q(
        \I_cache/cache[4][106] ), .QN(n1392) );
  DFFRX1 \I_cache/cache_reg[5][106]  ( .D(n11992), .CK(clk), .RN(n6049), .Q(
        \I_cache/cache[5][106] ), .QN(n3079) );
  DFFRX1 \I_cache/cache_reg[6][106]  ( .D(n11991), .CK(clk), .RN(n6049), .Q(
        \I_cache/cache[6][106] ), .QN(n1558) );
  DFFRX1 \I_cache/cache_reg[7][106]  ( .D(n11990), .CK(clk), .RN(n6049), .Q(
        \I_cache/cache[7][106] ), .QN(n3246) );
  DFFRX1 \I_cache/cache_reg[3][107]  ( .D(n11986), .CK(clk), .RN(n6048), .Q(
        \I_cache/cache[3][107] ), .QN(n3077) );
  DFFRX1 \I_cache/cache_reg[4][107]  ( .D(n11985), .CK(clk), .RN(n6048), .Q(
        \I_cache/cache[4][107] ), .QN(n1389) );
  DFFRX1 \I_cache/cache_reg[5][107]  ( .D(n11984), .CK(clk), .RN(n6048), .Q(
        \I_cache/cache[5][107] ), .QN(n3076) );
  DFFRX1 \I_cache/cache_reg[6][107]  ( .D(n11983), .CK(clk), .RN(n6048), .Q(
        \I_cache/cache[6][107] ), .QN(n1556) );
  DFFRX1 \I_cache/cache_reg[7][107]  ( .D(n11982), .CK(clk), .RN(n6048), .Q(
        \I_cache/cache[7][107] ), .QN(n3244) );
  DFFRX1 \I_cache/cache_reg[3][108]  ( .D(n11978), .CK(clk), .RN(n6048), .Q(
        \I_cache/cache[3][108] ), .QN(n3074) );
  DFFRX1 \I_cache/cache_reg[4][108]  ( .D(n11977), .CK(clk), .RN(n6047), .Q(
        \I_cache/cache[4][108] ), .QN(n1386) );
  DFFRX1 \I_cache/cache_reg[5][108]  ( .D(n11976), .CK(clk), .RN(n6047), .Q(
        \I_cache/cache[5][108] ), .QN(n3073) );
  DFFRX1 \I_cache/cache_reg[6][108]  ( .D(n11975), .CK(clk), .RN(n6047), .Q(
        \I_cache/cache[6][108] ), .QN(n1554) );
  DFFRX1 \I_cache/cache_reg[7][108]  ( .D(n11974), .CK(clk), .RN(n6047), .Q(
        \I_cache/cache[7][108] ), .QN(n3242) );
  DFFRX1 \I_cache/cache_reg[3][109]  ( .D(n11970), .CK(clk), .RN(n6047), .Q(
        \I_cache/cache[3][109] ), .QN(n3071) );
  DFFRX1 \I_cache/cache_reg[4][109]  ( .D(n11969), .CK(clk), .RN(n6047), .Q(
        \I_cache/cache[4][109] ), .QN(n1383) );
  DFFRX1 \I_cache/cache_reg[5][109]  ( .D(n11968), .CK(clk), .RN(n6047), .Q(
        \I_cache/cache[5][109] ), .QN(n3070) );
  DFFRX1 \I_cache/cache_reg[6][109]  ( .D(n11967), .CK(clk), .RN(n6047), .Q(
        \I_cache/cache[6][109] ), .QN(n1552) );
  DFFRX1 \I_cache/cache_reg[7][109]  ( .D(n11966), .CK(clk), .RN(n6047), .Q(
        \I_cache/cache[7][109] ), .QN(n3240) );
  DFFRX1 \I_cache/cache_reg[3][110]  ( .D(n11962), .CK(clk), .RN(n6046), .Q(
        \I_cache/cache[3][110] ), .QN(n3068) );
  DFFRX1 \I_cache/cache_reg[4][110]  ( .D(n11961), .CK(clk), .RN(n6046), .Q(
        \I_cache/cache[4][110] ), .QN(n1380) );
  DFFRX1 \I_cache/cache_reg[5][110]  ( .D(n11960), .CK(clk), .RN(n6046), .Q(
        \I_cache/cache[5][110] ), .QN(n3067) );
  DFFRX1 \I_cache/cache_reg[6][110]  ( .D(n11959), .CK(clk), .RN(n6046), .Q(
        \I_cache/cache[6][110] ), .QN(n1550) );
  DFFRX1 \I_cache/cache_reg[7][110]  ( .D(n11958), .CK(clk), .RN(n6046), .Q(
        \I_cache/cache[7][110] ), .QN(n3238) );
  DFFRX1 \I_cache/cache_reg[3][111]  ( .D(n11954), .CK(clk), .RN(n6046), .Q(
        \I_cache/cache[3][111] ), .QN(n3065) );
  DFFRX1 \I_cache/cache_reg[4][111]  ( .D(n11953), .CK(clk), .RN(n6045), .Q(
        \I_cache/cache[4][111] ), .QN(n1377) );
  DFFRX1 \I_cache/cache_reg[5][111]  ( .D(n11952), .CK(clk), .RN(n6045), .Q(
        \I_cache/cache[5][111] ), .QN(n3064) );
  DFFRX1 \I_cache/cache_reg[6][111]  ( .D(n11951), .CK(clk), .RN(n6045), .Q(
        \I_cache/cache[6][111] ), .QN(n1548) );
  DFFRX1 \I_cache/cache_reg[7][111]  ( .D(n11950), .CK(clk), .RN(n6045), .Q(
        \I_cache/cache[7][111] ), .QN(n3236) );
  DFFRX1 \I_cache/cache_reg[3][112]  ( .D(n11946), .CK(clk), .RN(n6045), .Q(
        \I_cache/cache[3][112] ), .QN(n3062) );
  DFFRX1 \I_cache/cache_reg[4][112]  ( .D(n11945), .CK(clk), .RN(n6045), .Q(
        \I_cache/cache[4][112] ), .QN(n1374) );
  DFFRX1 \I_cache/cache_reg[5][112]  ( .D(n11944), .CK(clk), .RN(n6045), .Q(
        \I_cache/cache[5][112] ), .QN(n3061) );
  DFFRX1 \I_cache/cache_reg[6][112]  ( .D(n11943), .CK(clk), .RN(n6045), .Q(
        \I_cache/cache[6][112] ), .QN(n1546) );
  DFFRX1 \I_cache/cache_reg[7][112]  ( .D(n11942), .CK(clk), .RN(n6045), .Q(
        \I_cache/cache[7][112] ), .QN(n3234) );
  DFFRX1 \I_cache/cache_reg[3][113]  ( .D(n11938), .CK(clk), .RN(n6044), .Q(
        \I_cache/cache[3][113] ), .QN(n3059) );
  DFFRX1 \I_cache/cache_reg[4][113]  ( .D(n11937), .CK(clk), .RN(n6044), .Q(
        \I_cache/cache[4][113] ), .QN(n1371) );
  DFFRX1 \I_cache/cache_reg[5][113]  ( .D(n11936), .CK(clk), .RN(n6044), .Q(
        \I_cache/cache[5][113] ), .QN(n3058) );
  DFFRX1 \I_cache/cache_reg[6][113]  ( .D(n11935), .CK(clk), .RN(n6044), .Q(
        \I_cache/cache[6][113] ), .QN(n1344) );
  DFFRX1 \I_cache/cache_reg[7][113]  ( .D(n11934), .CK(clk), .RN(n6044), .Q(
        \I_cache/cache[7][113] ), .QN(n3232) );
  DFFRX1 \I_cache/cache_reg[3][114]  ( .D(n11930), .CK(clk), .RN(n6044), .Q(
        \I_cache/cache[3][114] ), .QN(n3057) );
  DFFRX1 \I_cache/cache_reg[4][114]  ( .D(n11929), .CK(clk), .RN(n6043), .Q(
        \I_cache/cache[4][114] ), .QN(n1369) );
  DFFRX1 \I_cache/cache_reg[5][114]  ( .D(n11928), .CK(clk), .RN(n6043), .Q(
        \I_cache/cache[5][114] ), .QN(n3056) );
  DFFRX1 \I_cache/cache_reg[6][114]  ( .D(n11927), .CK(clk), .RN(n6043), .Q(
        \I_cache/cache[6][114] ), .QN(n1543) );
  DFFRX1 \I_cache/cache_reg[7][114]  ( .D(n11926), .CK(clk), .RN(n6043), .Q(
        \I_cache/cache[7][114] ), .QN(n3230) );
  DFFRX1 \I_cache/cache_reg[3][115]  ( .D(n11922), .CK(clk), .RN(n6043), .Q(
        \I_cache/cache[3][115] ), .QN(n3282) );
  DFFRX1 \I_cache/cache_reg[4][115]  ( .D(n11921), .CK(clk), .RN(n6043), .Q(
        \I_cache/cache[4][115] ), .QN(n1594) );
  DFFRX1 \I_cache/cache_reg[5][115]  ( .D(n11920), .CK(clk), .RN(n6043), .Q(
        \I_cache/cache[5][115] ), .QN(n3281) );
  DFFRX1 \I_cache/cache_reg[6][115]  ( .D(n11919), .CK(clk), .RN(n6043), .Q(
        \I_cache/cache[6][115] ), .QN(n1599) );
  DFFRX1 \I_cache/cache_reg[7][115]  ( .D(n11918), .CK(clk), .RN(n6043), .Q(
        \I_cache/cache[7][115] ), .QN(n3286) );
  DFFRX1 \I_cache/cache_reg[3][116]  ( .D(n11914), .CK(clk), .RN(n6042), .Q(
        \I_cache/cache[3][116] ), .QN(n3054) );
  DFFRX1 \I_cache/cache_reg[4][116]  ( .D(n11913), .CK(clk), .RN(n6042), .Q(
        \I_cache/cache[4][116] ), .QN(n1366) );
  DFFRX1 \I_cache/cache_reg[5][116]  ( .D(n11912), .CK(clk), .RN(n6042), .Q(
        \I_cache/cache[5][116] ), .QN(n3053) );
  DFFRX1 \I_cache/cache_reg[6][116]  ( .D(n11911), .CK(clk), .RN(n6042), .Q(
        \I_cache/cache[6][116] ), .QN(n1541) );
  DFFRX1 \I_cache/cache_reg[7][116]  ( .D(n11910), .CK(clk), .RN(n6042), .Q(
        \I_cache/cache[7][116] ), .QN(n3228) );
  DFFRX1 \I_cache/cache_reg[3][117]  ( .D(n11906), .CK(clk), .RN(n6042), .Q(
        \I_cache/cache[3][117] ), .QN(n3051) );
  DFFRX1 \I_cache/cache_reg[4][117]  ( .D(n11905), .CK(clk), .RN(n6041), .Q(
        \I_cache/cache[4][117] ), .QN(n1363) );
  DFFRX1 \I_cache/cache_reg[5][117]  ( .D(n11904), .CK(clk), .RN(n6041), .Q(
        \I_cache/cache[5][117] ), .QN(n3050) );
  DFFRX1 \I_cache/cache_reg[6][117]  ( .D(n11903), .CK(clk), .RN(n6041), .Q(
        \I_cache/cache[6][117] ), .QN(n1539) );
  DFFRX1 \I_cache/cache_reg[7][117]  ( .D(n11902), .CK(clk), .RN(n6041), .Q(
        \I_cache/cache[7][117] ), .QN(n3226) );
  DFFRX1 \I_cache/cache_reg[3][118]  ( .D(n11898), .CK(clk), .RN(n6041), .Q(
        \I_cache/cache[3][118] ), .QN(n3048) );
  DFFRX1 \I_cache/cache_reg[4][118]  ( .D(n11897), .CK(clk), .RN(n6041), .Q(
        \I_cache/cache[4][118] ), .QN(n1360) );
  DFFRX1 \I_cache/cache_reg[5][118]  ( .D(n11896), .CK(clk), .RN(n6041), .Q(
        \I_cache/cache[5][118] ), .QN(n3047) );
  DFFRX1 \I_cache/cache_reg[6][118]  ( .D(n11895), .CK(clk), .RN(n6041), .Q(
        \I_cache/cache[6][118] ), .QN(n1537) );
  DFFRX1 \I_cache/cache_reg[7][118]  ( .D(n11894), .CK(clk), .RN(n6041), .Q(
        \I_cache/cache[7][118] ), .QN(n3224) );
  DFFRX1 \I_cache/cache_reg[3][119]  ( .D(n11890), .CK(clk), .RN(n6040), .Q(
        \I_cache/cache[3][119] ), .QN(n3045) );
  DFFRX1 \I_cache/cache_reg[4][119]  ( .D(n11889), .CK(clk), .RN(n6040), .Q(
        \I_cache/cache[4][119] ), .QN(n1357) );
  DFFRX1 \I_cache/cache_reg[5][119]  ( .D(n11888), .CK(clk), .RN(n6040), .Q(
        \I_cache/cache[5][119] ), .QN(n3044) );
  DFFRX1 \I_cache/cache_reg[6][119]  ( .D(n11887), .CK(clk), .RN(n6040), .Q(
        \I_cache/cache[6][119] ), .QN(n1535) );
  DFFRX1 \I_cache/cache_reg[7][119]  ( .D(n11886), .CK(clk), .RN(n6040), .Q(
        \I_cache/cache[7][119] ), .QN(n3222) );
  DFFRX1 \I_cache/cache_reg[3][120]  ( .D(n11882), .CK(clk), .RN(n6040), .Q(
        \I_cache/cache[3][120] ), .QN(n3042) );
  DFFRX1 \I_cache/cache_reg[4][120]  ( .D(n11881), .CK(clk), .RN(n6039), .Q(
        \I_cache/cache[4][120] ), .QN(n1354) );
  DFFRX1 \I_cache/cache_reg[5][120]  ( .D(n11880), .CK(clk), .RN(n6039), .Q(
        \I_cache/cache[5][120] ), .QN(n3041) );
  DFFRX1 \I_cache/cache_reg[6][120]  ( .D(n11879), .CK(clk), .RN(n6039), .Q(
        \I_cache/cache[6][120] ), .QN(n1533) );
  DFFRX1 \I_cache/cache_reg[7][120]  ( .D(n11878), .CK(clk), .RN(n6039), .Q(
        \I_cache/cache[7][120] ), .QN(n3220) );
  DFFRX1 \I_cache/cache_reg[3][121]  ( .D(n11874), .CK(clk), .RN(n6039), .Q(
        \I_cache/cache[3][121] ), .QN(n3039) );
  DFFRX1 \I_cache/cache_reg[4][121]  ( .D(n11873), .CK(clk), .RN(n6039), .Q(
        \I_cache/cache[4][121] ), .QN(n1351) );
  DFFRX1 \I_cache/cache_reg[5][121]  ( .D(n11872), .CK(clk), .RN(n6039), .Q(
        \I_cache/cache[5][121] ), .QN(n3038) );
  DFFRX1 \I_cache/cache_reg[6][121]  ( .D(n11871), .CK(clk), .RN(n6039), .Q(
        \I_cache/cache[6][121] ), .QN(n1531) );
  DFFRX1 \I_cache/cache_reg[7][121]  ( .D(n11870), .CK(clk), .RN(n6039), .Q(
        \I_cache/cache[7][121] ), .QN(n3218) );
  DFFRX1 \I_cache/cache_reg[3][122]  ( .D(n11866), .CK(clk), .RN(n6038), .Q(
        \I_cache/cache[3][122] ), .QN(n3125) );
  DFFRX1 \I_cache/cache_reg[4][122]  ( .D(n11865), .CK(clk), .RN(n6038), .Q(
        \I_cache/cache[4][122] ), .QN(n1437) );
  DFFRX1 \I_cache/cache_reg[5][122]  ( .D(n11864), .CK(clk), .RN(n6038), .Q(
        \I_cache/cache[5][122] ), .QN(n3124) );
  DFFRX1 \I_cache/cache_reg[6][122]  ( .D(n11863), .CK(clk), .RN(n6038), .Q(
        \I_cache/cache[6][122] ), .QN(n1587) );
  DFFRX1 \I_cache/cache_reg[7][122]  ( .D(n11862), .CK(clk), .RN(n6038), .Q(
        \I_cache/cache[7][122] ), .QN(n3274) );
  DFFRX1 \I_cache/cache_reg[3][123]  ( .D(n11858), .CK(clk), .RN(n6038), .Q(
        \I_cache/cache[3][123] ), .QN(n3122) );
  DFFRX1 \I_cache/cache_reg[4][123]  ( .D(n11857), .CK(clk), .RN(n6037), .Q(
        \I_cache/cache[4][123] ), .QN(n1434) );
  DFFRX1 \I_cache/cache_reg[5][123]  ( .D(n11856), .CK(clk), .RN(n6037), .Q(
        \I_cache/cache[5][123] ), .QN(n3121) );
  DFFRX1 \I_cache/cache_reg[6][123]  ( .D(n11855), .CK(clk), .RN(n6037), .Q(
        \I_cache/cache[6][123] ), .QN(n1585) );
  DFFRX1 \I_cache/cache_reg[7][123]  ( .D(n11854), .CK(clk), .RN(n6037), .Q(
        \I_cache/cache[7][123] ), .QN(n3272) );
  DFFRX1 \I_cache/cache_reg[3][124]  ( .D(n11850), .CK(clk), .RN(n6037), .Q(
        \I_cache/cache[3][124] ), .QN(n3119) );
  DFFRX1 \I_cache/cache_reg[4][124]  ( .D(n11849), .CK(clk), .RN(n6037), .Q(
        \I_cache/cache[4][124] ), .QN(n1431) );
  DFFRX1 \I_cache/cache_reg[5][124]  ( .D(n11848), .CK(clk), .RN(n6037), .Q(
        \I_cache/cache[5][124] ), .QN(n3118) );
  DFFRX1 \I_cache/cache_reg[6][124]  ( .D(n11847), .CK(clk), .RN(n6037), .Q(
        \I_cache/cache[6][124] ), .QN(n1583) );
  DFFRX1 \I_cache/cache_reg[7][124]  ( .D(n11846), .CK(clk), .RN(n6037), .Q(
        \I_cache/cache[7][124] ), .QN(n3270) );
  DFFRX1 \I_cache/cache_reg[3][125]  ( .D(n11842), .CK(clk), .RN(n6036), .Q(
        \I_cache/cache[3][125] ), .QN(n3116) );
  DFFRX1 \I_cache/cache_reg[4][125]  ( .D(n11841), .CK(clk), .RN(n6036), .Q(
        \I_cache/cache[4][125] ), .QN(n1428) );
  DFFRX1 \I_cache/cache_reg[5][125]  ( .D(n11840), .CK(clk), .RN(n6036), .Q(
        \I_cache/cache[5][125] ), .QN(n3115) );
  DFFRX1 \I_cache/cache_reg[6][125]  ( .D(n11839), .CK(clk), .RN(n6036), .Q(
        \I_cache/cache[6][125] ), .QN(n1581) );
  DFFRX1 \I_cache/cache_reg[7][125]  ( .D(n11838), .CK(clk), .RN(n6036), .Q(
        \I_cache/cache[7][125] ), .QN(n3268) );
  DFFRX1 \I_cache/cache_reg[3][126]  ( .D(n11834), .CK(clk), .RN(n6036), .Q(
        \I_cache/cache[3][126] ), .QN(n3113) );
  DFFRX1 \I_cache/cache_reg[4][126]  ( .D(n11833), .CK(clk), .RN(n6035), .Q(
        \I_cache/cache[4][126] ), .QN(n1425) );
  DFFRX1 \I_cache/cache_reg[5][126]  ( .D(n11832), .CK(clk), .RN(n6035), .Q(
        \I_cache/cache[5][126] ), .QN(n3112) );
  DFFRX1 \I_cache/cache_reg[6][126]  ( .D(n11831), .CK(clk), .RN(n6035), .Q(
        \I_cache/cache[6][126] ), .QN(n1579) );
  DFFRX1 \I_cache/cache_reg[7][126]  ( .D(n11830), .CK(clk), .RN(n6035), .Q(
        \I_cache/cache[7][126] ), .QN(n3266) );
  DFFRX1 \I_cache/cache_reg[3][127]  ( .D(n11826), .CK(clk), .RN(n6035), .Q(
        \I_cache/cache[3][127] ), .QN(n3110) );
  DFFRX1 \I_cache/cache_reg[4][127]  ( .D(n11825), .CK(clk), .RN(n6035), .Q(
        \I_cache/cache[4][127] ), .QN(n1422) );
  DFFRX1 \I_cache/cache_reg[5][127]  ( .D(n11824), .CK(clk), .RN(n6035), .Q(
        \I_cache/cache[5][127] ), .QN(n3109) );
  DFFRX1 \I_cache/cache_reg[6][127]  ( .D(n11823), .CK(clk), .RN(n6035), .Q(
        \I_cache/cache[6][127] ), .QN(n1578) );
  DFFRX1 \I_cache/cache_reg[7][127]  ( .D(n11822), .CK(clk), .RN(n6035), .Q(
        \I_cache/cache[7][127] ), .QN(n3265) );
  DFFRX1 \I_cache/cache_reg[0][153]  ( .D(n11621), .CK(clk), .RN(n6018), .Q(
        \I_cache/cache[0][153] ), .QN(n2582) );
  DFFRX1 \I_cache/cache_reg[1][153]  ( .D(n11620), .CK(clk), .RN(n6018), .Q(
        \I_cache/cache[1][153] ), .QN(n1076) );
  DFFRX1 \I_cache/cache_reg[2][153]  ( .D(n11619), .CK(clk), .RN(n6018), .Q(
        \I_cache/cache[2][153] ), .QN(n2583) );
  DFFRX1 \I_cache/cache_reg[3][153]  ( .D(n11618), .CK(clk), .RN(n6018), .Q(
        \I_cache/cache[3][153] ), .QN(n1077) );
  DFFRX1 \I_cache/cache_reg[4][153]  ( .D(n11617), .CK(clk), .RN(n6018), .Q(
        \I_cache/cache[4][153] ), .QN(n2584) );
  DFFRX1 \I_cache/cache_reg[5][153]  ( .D(n11616), .CK(clk), .RN(n6017), .Q(
        \I_cache/cache[5][153] ), .QN(n1078) );
  DFFRX1 \I_cache/cache_reg[6][153]  ( .D(n11615), .CK(clk), .RN(n6017), .Q(
        \I_cache/cache[6][153] ), .QN(n1286) );
  DFFRX1 \I_cache/cache_reg[7][153]  ( .D(n11614), .CK(clk), .RN(n6017), .Q(
        \I_cache/cache[7][153] ), .QN(n2935) );
  DFFRX1 \D_cache/cache_reg[6][136]  ( .D(\D_cache/n702 ), .CK(clk), .RN(n6132), .Q(\D_cache/cache[6][136] ), .QN(n2113) );
  DFFRX1 \D_cache/cache_reg[7][148]  ( .D(\D_cache/n605 ), .CK(clk), .RN(n6124), .Q(\D_cache/cache[7][148] ), .QN(n2037) );
  DFFRX1 \D_cache/cache_reg[2][137]  ( .D(\D_cache/n698 ), .CK(clk), .RN(n6132), .Q(\D_cache/cache[2][137] ), .QN(n2082) );
  DFFRX1 \D_cache/cache_reg[6][131]  ( .D(\D_cache/n742 ), .CK(clk), .RN(n6135), .Q(\D_cache/cache[6][131] ), .QN(n2069) );
  DFFRX1 \D_cache/cache_reg[7][142]  ( .D(\D_cache/n653 ), .CK(clk), .RN(n6128), .Q(\D_cache/cache[7][142] ), .QN(n489) );
  DFFRX1 \D_cache/cache_reg[3][129]  ( .D(\D_cache/n761 ), .CK(clk), .RN(n6137), .Q(\D_cache/cache[3][129] ), .QN(n501) );
  DFFRX1 \D_cache/cache_reg[6][133]  ( .D(\D_cache/n726 ), .CK(clk), .RN(n6134), .Q(\D_cache/cache[6][133] ), .QN(n2129) );
  DFFRX1 \D_cache/cache_reg[2][130]  ( .D(\D_cache/n754 ), .CK(clk), .RN(n6136), .Q(\D_cache/cache[2][130] ), .QN(n2120) );
  DFFRX1 \D_cache/cache_reg[3][138]  ( .D(\D_cache/n689 ), .CK(clk), .RN(n6131), .Q(\D_cache/cache[3][138] ), .QN(n477) );
  DFFRX1 \D_cache/cache_reg[3][139]  ( .D(\D_cache/n681 ), .CK(clk), .RN(n6130), .Q(\D_cache/cache[3][139] ), .QN(n2034) );
  DFFRX1 \D_cache/cache_reg[6][137]  ( .D(\D_cache/n694 ), .CK(clk), .RN(n6131), .Q(\D_cache/cache[6][137] ), .QN(n2070) );
  DFFRX1 \D_cache/cache_reg[7][129]  ( .D(\D_cache/n757 ), .CK(clk), .RN(n6137), .Q(\D_cache/cache[7][129] ), .QN(n443) );
  DFFRX1 \D_cache/cache_reg[6][130]  ( .D(\D_cache/n750 ), .CK(clk), .RN(n6136), .Q(\D_cache/cache[6][130] ), .QN(n2153) );
  DFFRX1 \D_cache/cache_reg[7][138]  ( .D(\D_cache/n685 ), .CK(clk), .RN(n6131), .Q(\D_cache/cache[7][138] ), .QN(n498) );
  DFFRX1 \D_cache/cache_reg[3][134]  ( .D(\D_cache/n721 ), .CK(clk), .RN(n6134), .Q(\D_cache/cache[3][134] ), .QN(n494) );
  DFFRX1 \D_cache/cache_reg[3][132]  ( .D(\D_cache/n737 ), .CK(clk), .RN(n6135), .Q(\D_cache/cache[3][132] ), .QN(n518) );
  DFFRX1 \D_cache/cache_reg[3][136]  ( .D(\D_cache/n705 ), .CK(clk), .RN(n6132), .Q(\D_cache/cache[3][136] ), .QN(n462) );
  DFFRX1 \D_cache/cache_reg[2][140]  ( .D(\D_cache/n674 ), .CK(clk), .RN(n6130), .Q(\D_cache/cache[2][140] ), .QN(n2108) );
  DFFRX1 \D_cache/cache_reg[3][133]  ( .D(\D_cache/n729 ), .CK(clk), .RN(n6134), .Q(\D_cache/cache[3][133] ), .QN(n496) );
  DFFRX1 \D_cache/cache_reg[7][134]  ( .D(\D_cache/n717 ), .CK(clk), .RN(n6133), .Q(\D_cache/cache[7][134] ), .QN(n2038) );
  DFFRX1 \D_cache/cache_reg[7][132]  ( .D(\D_cache/n733 ), .CK(clk), .RN(n6135), .Q(\D_cache/cache[7][132] ), .QN(n2039) );
  DFFRX1 \I_cache/cache_reg[0][149]  ( .D(n11653), .CK(clk), .RN(n6021), .Q(
        \I_cache/cache[0][149] ), .QN(n984) );
  DFFRX1 \D_cache/cache_reg[7][144]  ( .D(\D_cache/n637 ), .CK(clk), .RN(n6127), .Q(\D_cache/cache[7][144] ), .QN(n2035) );
  DFFRX1 \D_cache/cache_reg[7][136]  ( .D(\D_cache/n701 ), .CK(clk), .RN(n6132), .Q(\D_cache/cache[7][136] ), .QN(n487) );
  DFFRX1 \D_cache/cache_reg[3][137]  ( .D(\D_cache/n697 ), .CK(clk), .RN(n6132), .Q(\D_cache/cache[3][137] ), .QN(n456) );
  DFFRX1 \D_cache/cache_reg[7][131]  ( .D(\D_cache/n741 ), .CK(clk), .RN(n6135), .Q(\D_cache/cache[7][131] ), .QN(n444) );
  DFFRX1 \D_cache/cache_reg[7][133]  ( .D(\D_cache/n725 ), .CK(clk), .RN(n6134), .Q(\D_cache/cache[7][133] ), .QN(n504) );
  DFFRX1 \D_cache/cache_reg[3][130]  ( .D(\D_cache/n753 ), .CK(clk), .RN(n6136), .Q(\D_cache/cache[3][130] ), .QN(n495) );
  DFFRX1 \D_cache/cache_reg[6][135]  ( .D(\D_cache/n710 ), .CK(clk), .RN(n6133), .Q(\D_cache/cache[6][135] ), .QN(n2131) );
  DFFRX1 \I_cache/cache_reg[2][149]  ( .D(n11651), .CK(clk), .RN(n6020), .Q(
        \I_cache/cache[2][149] ), .QN(n1227) );
  DFFRX1 \I_cache/cache_reg[0][147]  ( .D(n11669), .CK(clk), .RN(n6022), .Q(
        \I_cache/cache[0][147] ), .QN(n2066) );
  DFFRX1 \D_cache/cache_reg[7][137]  ( .D(\D_cache/n693 ), .CK(clk), .RN(n6131), .Q(\D_cache/cache[7][137] ), .QN(n445) );
  DFFRX1 \D_cache/cache_reg[7][130]  ( .D(\D_cache/n749 ), .CK(clk), .RN(n6136), .Q(\D_cache/cache[7][130] ), .QN(n528) );
  DFFRX1 \I_cache/cache_reg[0][148]  ( .D(n11661), .CK(clk), .RN(n6021), .Q(
        \I_cache/cache[0][148] ), .QN(n572) );
  DFFRX1 \I_cache/cache_reg[4][149]  ( .D(n11649), .CK(clk), .RN(n6020), .Q(
        \I_cache/cache[4][149] ), .QN(n2100) );
  DFFRX1 \D_cache/cache_reg[7][135]  ( .D(\D_cache/n709 ), .CK(clk), .RN(n6133), .Q(\D_cache/cache[7][135] ), .QN(n506) );
  DFFRX1 \I_cache/cache_reg[0][144]  ( .D(n11693), .CK(clk), .RN(n6024), .Q(
        \I_cache/cache[0][144] ), .QN(n2086) );
  DFFRX1 \I_cache/cache_reg[2][147]  ( .D(n11667), .CK(clk), .RN(n6022), .Q(
        \I_cache/cache[2][147] ), .QN(n2099) );
  DFFRX1 \I_cache/cache_reg[6][149]  ( .D(n11647), .CK(clk), .RN(n6020), .Q(
        \I_cache/cache[6][149] ), .QN(n964) );
  DFFRX1 \I_cache/cache_reg[1][149]  ( .D(n11652), .CK(clk), .RN(n6020), .Q(
        \I_cache/cache[1][149] ), .QN(n2609) );
  DFFRX1 \I_cache/cache_reg[0][129]  ( .D(n11813), .CK(clk), .RN(n6034), .Q(
        \I_cache/cache[0][129] ), .QN(n627) );
  DFFRX1 \D_cache/cache_reg[3][140]  ( .D(\D_cache/n673 ), .CK(clk), .RN(n6130), .Q(\D_cache/cache[3][140] ), .QN(n482) );
  DFFRX1 \I_cache/cache_reg[2][148]  ( .D(n11659), .CK(clk), .RN(n6021), .Q(
        \I_cache/cache[2][148] ), .QN(n2118) );
  DFFRX1 \I_cache/cache_reg[4][147]  ( .D(n11665), .CK(clk), .RN(n6022), .Q(
        \I_cache/cache[4][147] ), .QN(n571) );
  DFFRX1 \I_cache/cache_reg[2][144]  ( .D(n11691), .CK(clk), .RN(n6024), .Q(
        \I_cache/cache[2][144] ), .QN(n570) );
  DFFRX1 \I_cache/cache_reg[4][148]  ( .D(n11657), .CK(clk), .RN(n6021), .Q(
        \I_cache/cache[4][148] ), .QN(n629) );
  DFFRX1 \I_cache/cache_reg[0][130]  ( .D(n11805), .CK(clk), .RN(n6033), .Q(
        \I_cache/cache[0][130] ), .QN(n2146) );
  DFFRX1 \I_cache/cache_reg[6][147]  ( .D(n11663), .CK(clk), .RN(n6021), .Q(
        \I_cache/cache[6][147] ), .QN(n598) );
  DFFRX1 \I_cache/cache_reg[1][147]  ( .D(n11668), .CK(clk), .RN(n6022), .Q(
        \I_cache/cache[1][147] ), .QN(n441) );
  DFFRX1 \I_cache/cache_reg[2][129]  ( .D(n11811), .CK(clk), .RN(n6034), .Q(
        \I_cache/cache[2][129] ), .QN(n589) );
  DFFRX1 \I_cache/cache_reg[3][149]  ( .D(n11650), .CK(clk), .RN(n6020), .Q(
        \I_cache/cache[3][149] ), .QN(n2850) );
  DFFRX1 \I_cache/cache_reg[4][144]  ( .D(n11689), .CK(clk), .RN(n6024), .Q(
        \I_cache/cache[4][144] ), .QN(n2064) );
  DFFRX1 \I_cache/cache_reg[6][148]  ( .D(n11655), .CK(clk), .RN(n6021), .Q(
        \I_cache/cache[6][148] ), .QN(n2081) );
  DFFRX1 \I_cache/cache_reg[1][148]  ( .D(n11660), .CK(clk), .RN(n6021), .Q(
        \I_cache/cache[1][148] ), .QN(n2190) );
  DFFRX1 \I_cache/cache_reg[4][129]  ( .D(n11809), .CK(clk), .RN(n6034), .Q(
        \I_cache/cache[4][129] ), .QN(n2076) );
  DFFRX1 \I_cache/cache_reg[6][144]  ( .D(n11687), .CK(clk), .RN(n6023), .Q(
        \I_cache/cache[6][144] ), .QN(n433) );
  DFFRX1 \I_cache/cache_reg[1][144]  ( .D(n11692), .CK(clk), .RN(n6024), .Q(
        \I_cache/cache[1][144] ), .QN(n460) );
  DFFRX1 \I_cache/cache_reg[2][130]  ( .D(n11803), .CK(clk), .RN(n6033), .Q(
        \I_cache/cache[2][130] ), .QN(n573) );
  DFFRX1 \I_cache/cache_reg[3][147]  ( .D(n11666), .CK(clk), .RN(n6022), .Q(
        \I_cache/cache[3][147] ), .QN(n473) );
  DFFRX1 \I_cache/cache_reg[5][149]  ( .D(n11648), .CK(clk), .RN(n6020), .Q(
        \I_cache/cache[5][149] ), .QN(n474) );
  DFFRX1 \I_cache/cache_reg[1][129]  ( .D(n11812), .CK(clk), .RN(n6034), .Q(
        \I_cache/cache[1][129] ), .QN(n2245) );
  DFFRX1 \I_cache/cache_reg[6][129]  ( .D(n11807), .CK(clk), .RN(n6033), .Q(
        \I_cache/cache[6][129] ), .QN(n576) );
  DFFRX1 \I_cache/cache_reg[4][130]  ( .D(n11801), .CK(clk), .RN(n6033), .Q(
        \I_cache/cache[4][130] ), .QN(n2062) );
  DFFRX1 \I_cache/cache_reg[3][148]  ( .D(n11658), .CK(clk), .RN(n6021), .Q(
        \I_cache/cache[3][148] ), .QN(n492) );
  DFFRX1 \I_cache/cache_reg[3][144]  ( .D(n11690), .CK(clk), .RN(n6024), .Q(
        \I_cache/cache[3][144] ), .QN(n2188) );
  DFFRX1 \I_cache/cache_reg[1][130]  ( .D(n11804), .CK(clk), .RN(n6033), .Q(
        \I_cache/cache[1][130] ), .QN(n521) );
  DFFRX1 \I_cache/cache_reg[5][147]  ( .D(n11664), .CK(clk), .RN(n6021), .Q(
        \I_cache/cache[5][147] ), .QN(n2189) );
  DFFRX1 \I_cache/cache_reg[7][149]  ( .D(n11646), .CK(clk), .RN(n6020), .Q(
        \I_cache/cache[7][149] ), .QN(n2589) );
  DFFRX1 \I_cache/cache_reg[6][130]  ( .D(n11799), .CK(clk), .RN(n6033), .Q(
        \I_cache/cache[6][130] ), .QN(n2078) );
  DFFRX1 \I_cache/cache_reg[3][129]  ( .D(n11810), .CK(clk), .RN(n6034), .Q(
        \I_cache/cache[3][129] ), .QN(n2207) );
  DFFRX1 \I_cache/cache_reg[5][148]  ( .D(n11656), .CK(clk), .RN(n6021), .Q(
        \I_cache/cache[5][148] ), .QN(n2246) );
  DFFRX1 \I_cache/cache_reg[5][144]  ( .D(n11688), .CK(clk), .RN(n6023), .Q(
        \I_cache/cache[5][144] ), .QN(n439) );
  DFFRX1 \I_cache/cache_reg[3][130]  ( .D(n11802), .CK(clk), .RN(n6033), .Q(
        \I_cache/cache[3][130] ), .QN(n2191) );
  DFFRX1 \I_cache/cache_reg[7][147]  ( .D(n11662), .CK(clk), .RN(n6021), .Q(
        \I_cache/cache[7][147] ), .QN(n2216) );
  DFFRX1 \I_cache/cache_reg[5][129]  ( .D(n11808), .CK(clk), .RN(n6033), .Q(
        \I_cache/cache[5][129] ), .QN(n451) );
  DFFRX1 \I_cache/cache_reg[7][148]  ( .D(n11654), .CK(clk), .RN(n6021), .Q(
        \I_cache/cache[7][148] ), .QN(n435) );
  DFFRX1 \I_cache/cache_reg[7][144]  ( .D(n11686), .CK(clk), .RN(n6023), .Q(
        \I_cache/cache[7][144] ), .QN(n2059) );
  DFFRX1 \I_cache/cache_reg[5][130]  ( .D(n11800), .CK(clk), .RN(n6033), .Q(
        \I_cache/cache[5][130] ), .QN(n437) );
  DFFRX1 \I_cache/cache_reg[7][129]  ( .D(n11806), .CK(clk), .RN(n6033), .Q(
        \I_cache/cache[7][129] ), .QN(n2194) );
  DFFRX1 \I_cache/cache_reg[7][130]  ( .D(n11798), .CK(clk), .RN(n6033), .Q(
        \I_cache/cache[7][130] ), .QN(n453) );
  DFFRX1 \I_cache/cache_reg[5][152]  ( .D(n11624), .CK(clk), .RN(n6018), .Q(
        \I_cache/cache[5][152] ) );
  DFFRX1 \D_cache/cache_reg[2][129]  ( .D(\D_cache/n762 ), .CK(clk), .RN(n6137), .Q(\D_cache/cache[2][129] ), .QN(n2126) );
  DFFRX1 \D_cache/cache_reg[6][129]  ( .D(\D_cache/n758 ), .CK(clk), .RN(n6137), .Q(\D_cache/cache[6][129] ), .QN(n2068) );
  DFFRX1 \D_cache/cache_reg[2][131]  ( .D(\D_cache/n746 ), .CK(clk), .RN(n6136), .Q(\D_cache/cache[2][131] ), .QN(n2058) );
  DFFRX1 \D_cache/cache_reg[2][132]  ( .D(\D_cache/n738 ), .CK(clk), .RN(n6135), .Q(\D_cache/cache[2][132] ), .QN(n2143) );
  DFFRX1 \D_cache/cache_reg[2][133]  ( .D(\D_cache/n730 ), .CK(clk), .RN(n6134), .Q(\D_cache/cache[2][133] ), .QN(n2121) );
  DFFRX1 \D_cache/cache_reg[2][134]  ( .D(\D_cache/n722 ), .CK(clk), .RN(n6134), .Q(\D_cache/cache[2][134] ), .QN(n2119) );
  DFFRX1 \D_cache/cache_reg[2][136]  ( .D(\D_cache/n706 ), .CK(clk), .RN(n6132), .Q(\D_cache/cache[2][136] ), .QN(n2088) );
  DFFRX1 \D_cache/cache_reg[2][138]  ( .D(\D_cache/n690 ), .CK(clk), .RN(n6131), .Q(\D_cache/cache[2][138] ), .QN(n2103) );
  DFFRX1 \D_cache/cache_reg[6][138]  ( .D(\D_cache/n686 ), .CK(clk), .RN(n6131), .Q(\D_cache/cache[6][138] ), .QN(n2123) );
  DFFRX1 \D_cache/cache_reg[0][139]  ( .D(\D_cache/n684 ), .CK(clk), .RN(n6131), .Q(\D_cache/cache[0][139] ), .QN(n1938) );
  DFFRX1 \D_cache/cache_reg[1][139]  ( .D(\D_cache/n683 ), .CK(clk), .RN(n6130), .Q(\D_cache/cache[1][139] ), .QN(n353) );
  DFFRX1 \D_cache/cache_reg[4][139]  ( .D(\D_cache/n680 ), .CK(clk), .RN(n6130), .Q(\D_cache/cache[4][139] ), .QN(n2024) );
  DFFRX1 \D_cache/cache_reg[5][139]  ( .D(\D_cache/n679 ), .CK(clk), .RN(n6130), .Q(\D_cache/cache[5][139] ), .QN(n405) );
  DFFRX1 \D_cache/cache_reg[0][140]  ( .D(\D_cache/n676 ), .CK(clk), .RN(n6130), .Q(\D_cache/cache[0][140] ), .QN(n2028) );
  DFFRX1 \D_cache/cache_reg[1][140]  ( .D(\D_cache/n675 ), .CK(clk), .RN(n6130), .Q(\D_cache/cache[1][140] ), .QN(n409) );
  DFFRX1 \D_cache/cache_reg[4][140]  ( .D(\D_cache/n672 ), .CK(clk), .RN(n6130), .Q(\D_cache/cache[4][140] ), .QN(n413) );
  DFFRX1 \D_cache/cache_reg[5][140]  ( .D(\D_cache/n671 ), .CK(clk), .RN(n6129), .Q(\D_cache/cache[5][140] ), .QN(n257) );
  DFFRX1 \D_cache/cache_reg[2][141]  ( .D(\D_cache/n666 ), .CK(clk), .RN(n6129), .Q(\D_cache/cache[2][141] ), .QN(n2105) );
  DFFRX1 \D_cache/cache_reg[3][141]  ( .D(\D_cache/n665 ), .CK(clk), .RN(n6129), .Q(\D_cache/cache[3][141] ), .QN(n479) );
  DFFRX1 \D_cache/cache_reg[6][141]  ( .D(\D_cache/n662 ), .CK(clk), .RN(n6129), .Q(\D_cache/cache[6][141] ), .QN(n2073) );
  DFFRX1 \D_cache/cache_reg[7][141]  ( .D(\D_cache/n661 ), .CK(clk), .RN(n6129), .Q(\D_cache/cache[7][141] ), .QN(n448) );
  DFFRX1 \D_cache/cache_reg[2][142]  ( .D(\D_cache/n658 ), .CK(clk), .RN(n6128), .Q(\D_cache/cache[2][142] ), .QN(n2063) );
  DFFRX1 \D_cache/cache_reg[3][142]  ( .D(\D_cache/n657 ), .CK(clk), .RN(n6128), .Q(\D_cache/cache[3][142] ), .QN(n438) );
  DFFRX1 \D_cache/cache_reg[6][142]  ( .D(\D_cache/n654 ), .CK(clk), .RN(n6128), .Q(\D_cache/cache[6][142] ), .QN(n2115) );
  DFFRX1 \D_cache/cache_reg[2][143]  ( .D(\D_cache/n650 ), .CK(clk), .RN(n6128), .Q(\D_cache/cache[2][143] ), .QN(n2101) );
  DFFRX1 \D_cache/cache_reg[3][143]  ( .D(\D_cache/n649 ), .CK(clk), .RN(n6128), .Q(\D_cache/cache[3][143] ), .QN(n475) );
  DFFRX1 \D_cache/cache_reg[6][143]  ( .D(\D_cache/n646 ), .CK(clk), .RN(n6127), .Q(\D_cache/cache[6][143] ), .QN(n582) );
  DFFRX1 \D_cache/cache_reg[7][143]  ( .D(\D_cache/n645 ), .CK(clk), .RN(n6127), .Q(\D_cache/cache[7][143] ), .QN(n2200) );
  DFFRX1 \D_cache/cache_reg[0][144]  ( .D(\D_cache/n644 ), .CK(clk), .RN(n6127), .Q(\D_cache/cache[0][144] ), .QN(n2027) );
  DFFRX1 \D_cache/cache_reg[1][144]  ( .D(\D_cache/n643 ), .CK(clk), .RN(n6127), .Q(\D_cache/cache[1][144] ), .QN(n408) );
  DFFRX1 \D_cache/cache_reg[4][144]  ( .D(\D_cache/n640 ), .CK(clk), .RN(n6127), .Q(\D_cache/cache[4][144] ), .QN(n412) );
  DFFRX1 \D_cache/cache_reg[5][144]  ( .D(\D_cache/n639 ), .CK(clk), .RN(n6127), .Q(\D_cache/cache[5][144] ), .QN(n256) );
  DFFRX1 \D_cache/cache_reg[2][146]  ( .D(\D_cache/n626 ), .CK(clk), .RN(n6126), .Q(\D_cache/cache[2][146] ), .QN(n2040) );
  DFFRX1 \D_cache/cache_reg[6][146]  ( .D(\D_cache/n622 ), .CK(clk), .RN(n6125), .Q(\D_cache/cache[6][146] ), .QN(n2106) );
  DFFRX1 \D_cache/cache_reg[7][146]  ( .D(\D_cache/n621 ), .CK(clk), .RN(n6125), .Q(\D_cache/cache[7][146] ), .QN(n480) );
  DFFRX1 \D_cache/cache_reg[3][148]  ( .D(\D_cache/n609 ), .CK(clk), .RN(n6124), .Q(\D_cache/cache[3][148] ), .QN(n2036) );
  DFFRX1 \D_cache/cache_reg[2][151]  ( .D(\D_cache/n586 ), .CK(clk), .RN(n6122), .Q(\D_cache/cache[2][151] ), .QN(n2138) );
  DFFRX1 \D_cache/cache_reg[3][151]  ( .D(\D_cache/n585 ), .CK(clk), .RN(n6122), .Q(\D_cache/cache[3][151] ), .QN(n513) );
  DFFRX1 \D_cache/cache_reg[6][151]  ( .D(\D_cache/n582 ), .CK(clk), .RN(n6122), .Q(\D_cache/cache[6][151] ), .QN(n2065) );
  DFFRX1 \D_cache/cache_reg[7][151]  ( .D(\D_cache/n581 ), .CK(clk), .RN(n6122), .Q(\D_cache/cache[7][151] ), .QN(n440) );
  DFFRX1 \D_cache/cache_reg[0][152]  ( .D(\D_cache/n580 ), .CK(clk), .RN(n6122), .Q(\D_cache/cache[0][152] ), .QN(n2017) );
  DFFRX1 \D_cache/cache_reg[1][152]  ( .D(\D_cache/n579 ), .CK(clk), .RN(n6122), .Q(\D_cache/cache[1][152] ), .QN(n398) );
  DFFRX1 \D_cache/cache_reg[2][152]  ( .D(\D_cache/n578 ), .CK(clk), .RN(n6122), .Q(\D_cache/cache[2][152] ), .QN(n2112) );
  DFFRX1 \D_cache/cache_reg[3][152]  ( .D(\D_cache/n577 ), .CK(clk), .RN(n6122), .Q(\D_cache/cache[3][152] ), .QN(n486) );
  DFFRX1 \D_cache/cache_reg[4][152]  ( .D(\D_cache/n576 ), .CK(clk), .RN(n6122), .Q(\D_cache/cache[4][152] ), .QN(n2016) );
  DFFRX1 \D_cache/cache_reg[5][152]  ( .D(\D_cache/n575 ), .CK(clk), .RN(n6121), .Q(\D_cache/cache[5][152] ), .QN(n397) );
  DFFRX1 \D_cache/cache_reg[6][152]  ( .D(\D_cache/n574 ), .CK(clk), .RN(n6121), .Q(\D_cache/cache[6][152] ), .QN(n2109) );
  DFFRX1 \D_cache/cache_reg[7][152]  ( .D(\D_cache/n573 ), .CK(clk), .RN(n6121), .Q(\D_cache/cache[7][152] ), .QN(n483) );
  DFFRX1 \D_cache/cache_reg[4][143]  ( .D(\D_cache/n648 ), .CK(clk), .RN(n6128), .Q(\D_cache/cache[4][143] ), .QN(n2918) );
  DFFRX1 \D_cache/cache_reg[0][143]  ( .D(\D_cache/n652 ), .CK(clk), .RN(n6128), .Q(\D_cache/cache[0][143] ), .QN(n2354) );
  DFFRX1 \D_cache/cache_reg[1][143]  ( .D(\D_cache/n651 ), .CK(clk), .RN(n6128), .Q(\D_cache/cache[1][143] ), .QN(n904) );
  DFFRX1 \D_cache/cache_reg[2][128]  ( .D(\D_cache/n770 ), .CK(clk), .RN(n6138), .Q(\D_cache/cache[2][128] ), .QN(n2888) );
  DFFRX1 \D_cache/cache_reg[3][128]  ( .D(\D_cache/n769 ), .CK(clk), .RN(n6138), .Q(\D_cache/cache[3][128] ), .QN(n1270) );
  DFFRX1 \D_cache/cache_reg[6][128]  ( .D(\D_cache/n766 ), .CK(clk), .RN(n6137), .Q(\D_cache/cache[6][128] ), .QN(n2887) );
  DFFRX1 \D_cache/cache_reg[7][128]  ( .D(\D_cache/n765 ), .CK(clk), .RN(n6121), .Q(\D_cache/cache[7][128] ), .QN(n1269) );
  DFFRX1 \D_cache/cache_reg[4][146]  ( .D(\D_cache/n624 ), .CK(clk), .RN(n6126), .Q(\D_cache/cache[4][146] ), .QN(n2015) );
  DFFRX1 \D_cache/cache_reg[5][146]  ( .D(\D_cache/n623 ), .CK(clk), .RN(n6125), .Q(\D_cache/cache[5][146] ), .QN(n396) );
  DFFRX1 \D_cache/cache_reg[4][141]  ( .D(\D_cache/n664 ), .CK(clk), .RN(n6129), .Q(\D_cache/cache[4][141] ), .QN(n2023) );
  DFFRX1 \D_cache/cache_reg[5][141]  ( .D(\D_cache/n663 ), .CK(clk), .RN(n6129), .Q(\D_cache/cache[5][141] ), .QN(n404) );
  DFFRX1 \D_cache/cache_reg[0][146]  ( .D(\D_cache/n628 ), .CK(clk), .RN(n6126), .Q(\D_cache/cache[0][146] ), .QN(n1336) );
  DFFRX1 \D_cache/cache_reg[1][146]  ( .D(\D_cache/n627 ), .CK(clk), .RN(n6126), .Q(\D_cache/cache[1][146] ), .QN(n2989) );
  DFFRX1 \D_cache/cache_reg[0][141]  ( .D(\D_cache/n668 ), .CK(clk), .RN(n6129), .Q(\D_cache/cache[0][141] ), .QN(n2957) );
  DFFRX1 \D_cache/cache_reg[1][141]  ( .D(\D_cache/n667 ), .CK(clk), .RN(n6129), .Q(\D_cache/cache[1][141] ), .QN(n1316) );
  DFFRX1 \D_cache/cache_reg[4][138]  ( .D(\D_cache/n688 ), .CK(clk), .RN(n6131), .Q(\D_cache/cache[4][138] ), .QN(n2021) );
  DFFRX1 \D_cache/cache_reg[5][138]  ( .D(\D_cache/n687 ), .CK(clk), .RN(n6131), .Q(\D_cache/cache[5][138] ), .QN(n402) );
  DFFRX1 \D_cache/cache_reg[4][142]  ( .D(\D_cache/n656 ), .CK(clk), .RN(n6128), .Q(\D_cache/cache[4][142] ), .QN(n2022) );
  DFFRX1 \D_cache/cache_reg[5][142]  ( .D(\D_cache/n655 ), .CK(clk), .RN(n6128), .Q(\D_cache/cache[5][142] ), .QN(n403) );
  DFFRX1 \D_cache/cache_reg[0][142]  ( .D(\D_cache/n660 ), .CK(clk), .RN(n6129), .Q(\D_cache/cache[0][142] ), .QN(n1331) );
  DFFRX1 \D_cache/cache_reg[1][142]  ( .D(\D_cache/n659 ), .CK(clk), .RN(n6128), .Q(\D_cache/cache[1][142] ), .QN(n2984) );
  DFFRX1 \D_cache/cache_reg[4][131]  ( .D(\D_cache/n744 ), .CK(clk), .RN(n6136), .Q(\D_cache/cache[4][131] ), .QN(n2029) );
  DFFRX1 \D_cache/cache_reg[5][131]  ( .D(\D_cache/n743 ), .CK(clk), .RN(n6135), .Q(\D_cache/cache[5][131] ), .QN(n410) );
  DFFRX1 \D_cache/cache_reg[4][129]  ( .D(\D_cache/n760 ), .CK(clk), .RN(n6137), .Q(\D_cache/cache[4][129] ), .QN(n2014) );
  DFFRX1 \D_cache/cache_reg[5][129]  ( .D(\D_cache/n759 ), .CK(clk), .RN(n6137), .Q(\D_cache/cache[5][129] ), .QN(n395) );
  DFFRX1 \D_cache/cache_reg[4][134]  ( .D(\D_cache/n720 ), .CK(clk), .RN(n6134), .Q(\D_cache/cache[4][134] ), .QN(n2026) );
  DFFRX1 \D_cache/cache_reg[5][134]  ( .D(\D_cache/n719 ), .CK(clk), .RN(n6133), .Q(\D_cache/cache[5][134] ), .QN(n407) );
  DFFRX1 \D_cache/cache_reg[0][138]  ( .D(\D_cache/n692 ), .CK(clk), .RN(n6131), .Q(\D_cache/cache[0][138] ), .QN(n2019) );
  DFFRX1 \D_cache/cache_reg[1][138]  ( .D(\D_cache/n691 ), .CK(clk), .RN(n6131), .Q(\D_cache/cache[1][138] ), .QN(n400) );
  DFFRX1 \D_cache/cache_reg[0][131]  ( .D(\D_cache/n748 ), .CK(clk), .RN(n6136), .Q(\D_cache/cache[0][131] ), .QN(n2952) );
  DFFRX1 \D_cache/cache_reg[1][131]  ( .D(\D_cache/n747 ), .CK(clk), .RN(n6136), .Q(\D_cache/cache[1][131] ), .QN(n1311) );
  DFFRX1 \D_cache/cache_reg[4][133]  ( .D(\D_cache/n728 ), .CK(clk), .RN(n6134), .Q(\D_cache/cache[4][133] ), .QN(n2897) );
  DFFRX1 \D_cache/cache_reg[5][133]  ( .D(\D_cache/n727 ), .CK(clk), .RN(n6134), .Q(\D_cache/cache[5][133] ), .QN(n2352) );
  DFFRX1 \D_cache/cache_reg[0][129]  ( .D(\D_cache/n764 ), .CK(clk), .RN(n6137), .Q(\D_cache/cache[0][129] ), .QN(n2956) );
  DFFRX1 \D_cache/cache_reg[1][129]  ( .D(\D_cache/n763 ), .CK(clk), .RN(n6137), .Q(\D_cache/cache[1][129] ), .QN(n1315) );
  DFFRX1 \D_cache/cache_reg[4][130]  ( .D(\D_cache/n752 ), .CK(clk), .RN(n6136), .Q(\D_cache/cache[4][130] ), .QN(n414) );
  DFFRX1 \D_cache/cache_reg[5][130]  ( .D(\D_cache/n751 ), .CK(clk), .RN(n6136), .Q(\D_cache/cache[5][130] ), .QN(n258) );
  DFFRX1 \D_cache/cache_reg[0][134]  ( .D(\D_cache/n724 ), .CK(clk), .RN(n6134), .Q(\D_cache/cache[0][134] ), .QN(n2020) );
  DFFRX1 \D_cache/cache_reg[1][134]  ( .D(\D_cache/n723 ), .CK(clk), .RN(n6134), .Q(\D_cache/cache[1][134] ), .QN(n401) );
  DFFRX1 \D_cache/cache_reg[0][130]  ( .D(\D_cache/n756 ), .CK(clk), .RN(n6137), .Q(\D_cache/cache[0][130] ), .QN(n2958) );
  DFFRX1 \D_cache/cache_reg[1][130]  ( .D(\D_cache/n755 ), .CK(clk), .RN(n6136), .Q(\D_cache/cache[1][130] ), .QN(n1317) );
  DFFRX1 \D_cache/cache_reg[0][133]  ( .D(\D_cache/n732 ), .CK(clk), .RN(n6135), .Q(\D_cache/cache[0][133] ), .QN(n1338) );
  DFFRX1 \D_cache/cache_reg[1][133]  ( .D(\D_cache/n731 ), .CK(clk), .RN(n6134), .Q(\D_cache/cache[1][133] ), .QN(n2992) );
  DFFRX1 \D_cache/cache_reg[4][151]  ( .D(\D_cache/n584 ), .CK(clk), .RN(n6122), .Q(\D_cache/cache[4][151] ), .QN(n411) );
  DFFRX1 \D_cache/cache_reg[5][151]  ( .D(\D_cache/n583 ), .CK(clk), .RN(n6122), .Q(\D_cache/cache[5][151] ), .QN(n255) );
  DFFRX1 \D_cache/cache_reg[0][151]  ( .D(\D_cache/n588 ), .CK(clk), .RN(n6123), .Q(\D_cache/cache[0][151] ), .QN(n1337) );
  DFFRX1 \D_cache/cache_reg[1][151]  ( .D(\D_cache/n587 ), .CK(clk), .RN(n6122), .Q(\D_cache/cache[1][151] ), .QN(n2991) );
  DFFRX1 \D_cache/cache_reg[4][148]  ( .D(\D_cache/n608 ), .CK(clk), .RN(n6124), .Q(\D_cache/cache[4][148] ), .QN(n2018) );
  DFFRX1 \D_cache/cache_reg[5][148]  ( .D(\D_cache/n607 ), .CK(clk), .RN(n6124), .Q(\D_cache/cache[5][148] ), .QN(n399) );
  DFFRX1 \D_cache/cache_reg[4][137]  ( .D(\D_cache/n696 ), .CK(clk), .RN(n6132), .Q(\D_cache/cache[4][137] ), .QN(n2355) );
  DFFRX1 \D_cache/cache_reg[5][137]  ( .D(\D_cache/n695 ), .CK(clk), .RN(n6131), .Q(\D_cache/cache[5][137] ), .QN(n905) );
  DFFRX1 \D_cache/cache_reg[0][148]  ( .D(\D_cache/n612 ), .CK(clk), .RN(n6125), .Q(\D_cache/cache[0][148] ), .QN(n2891) );
  DFFRX1 \D_cache/cache_reg[1][148]  ( .D(\D_cache/n611 ), .CK(clk), .RN(n6124), .Q(\D_cache/cache[1][148] ), .QN(n2951) );
  DFFRX1 \D_cache/cache_reg[0][137]  ( .D(\D_cache/n700 ), .CK(clk), .RN(n6132), .Q(\D_cache/cache[0][137] ), .QN(n2898) );
  DFFRX1 \D_cache/cache_reg[4][132]  ( .D(\D_cache/n736 ), .CK(clk), .RN(n6135), .Q(\D_cache/cache[4][132] ), .QN(n906) );
  DFFRX1 \D_cache/cache_reg[5][132]  ( .D(\D_cache/n735 ), .CK(clk), .RN(n6135), .Q(\D_cache/cache[5][132] ), .QN(n299) );
  DFFRX1 \D_cache/cache_reg[4][136]  ( .D(\D_cache/n704 ), .CK(clk), .RN(n6132), .Q(\D_cache/cache[4][136] ), .QN(n2353) );
  DFFRX1 \D_cache/cache_reg[5][136]  ( .D(\D_cache/n703 ), .CK(clk), .RN(n6132), .Q(\D_cache/cache[5][136] ), .QN(n903) );
  DFFRX1 \D_cache/cache_reg[0][135]  ( .D(\D_cache/n716 ), .CK(clk), .RN(n6133), .Q(\D_cache/cache[0][135] ), .QN(n2177) );
  DFFRX1 \D_cache/cache_reg[1][135]  ( .D(\D_cache/n715 ), .CK(clk), .RN(n6133), .Q(\D_cache/cache[1][135] ), .QN(n2890) );
  DFFRX1 \D_cache/cache_reg[0][132]  ( .D(\D_cache/n740 ), .CK(clk), .RN(n6135), .Q(\D_cache/cache[0][132] ), .QN(n2959) );
  DFFRX1 \D_cache/cache_reg[1][132]  ( .D(\D_cache/n739 ), .CK(clk), .RN(n6135), .Q(\D_cache/cache[1][132] ), .QN(n1318) );
  DFFRX1 \D_cache/cache_reg[0][136]  ( .D(\D_cache/n708 ), .CK(clk), .RN(n6133), .Q(\D_cache/cache[0][136] ), .QN(n1332) );
  DFFRX1 \D_cache/cache_reg[1][136]  ( .D(\D_cache/n707 ), .CK(clk), .RN(n6132), .Q(\D_cache/cache[1][136] ), .QN(n2985) );
  DFFRX1 \D_cache/cache_reg[4][135]  ( .D(\D_cache/n712 ), .CK(clk), .RN(n6133), .Q(\D_cache/cache[4][135] ), .QN(n2025) );
  DFFRX1 \D_cache/cache_reg[5][135]  ( .D(\D_cache/n711 ), .CK(clk), .RN(n6133), .Q(\D_cache/cache[5][135] ), .QN(n406) );
  DFFRX1 \I_cache/cache_reg[0][128]  ( .D(n11821), .CK(clk), .RN(n6034), .Q(
        \I_cache/cache[0][128] ), .QN(n2154) );
  DFFRX1 \D_cache/cache_reg[6][149]  ( .D(\D_cache/n598 ), .CK(clk), .RN(n6123), .Q(\D_cache/cache[6][149] ), .QN(n434) );
  DFFRX1 \D_cache/cache_reg[7][149]  ( .D(\D_cache/n597 ), .CK(clk), .RN(n6123), .Q(\D_cache/cache[7][149] ), .QN(n2060) );
  DFFRX1 \I_cache/cache_reg[0][133]  ( .D(n11781), .CK(clk), .RN(n6031), .Q(
        \I_cache/cache[0][133] ), .QN(n2104) );
  DFFRX1 \D_cache/cache_reg[2][149]  ( .D(\D_cache/n602 ), .CK(clk), .RN(n6124), .Q(\D_cache/cache[2][149] ), .QN(n1339) );
  DFFRX1 \D_cache/cache_reg[3][149]  ( .D(\D_cache/n601 ), .CK(clk), .RN(n6124), .Q(\D_cache/cache[3][149] ), .QN(n2994) );
  DFFRX1 \I_cache/cache_reg[4][137]  ( .D(n11745), .CK(clk), .RN(n6028), .Q(
        \I_cache/cache[4][137] ), .QN(n2977) );
  DFFRX1 \I_cache/cache_reg[0][143]  ( .D(n11701), .CK(clk), .RN(n6025), .Q(
        \I_cache/cache[0][143] ), .QN(n612) );
  DFFRX1 \D_cache/cache_reg[6][150]  ( .D(\D_cache/n590 ), .CK(clk), .RN(n6123), .Q(\D_cache/cache[6][150] ), .QN(n588) );
  DFFRX1 \D_cache/cache_reg[7][150]  ( .D(\D_cache/n589 ), .CK(clk), .RN(n6123), .Q(\D_cache/cache[7][150] ), .QN(n2206) );
  DFFRX1 \D_cache/cache_reg[6][147]  ( .D(\D_cache/n614 ), .CK(clk), .RN(n6125), .Q(\D_cache/cache[6][147] ), .QN(n586) );
  DFFRX1 \D_cache/cache_reg[7][147]  ( .D(\D_cache/n613 ), .CK(clk), .RN(n6125), .Q(\D_cache/cache[7][147] ), .QN(n2204) );
  DFFRX1 \D_cache/cache_reg[6][145]  ( .D(\D_cache/n630 ), .CK(clk), .RN(n6126), .Q(\D_cache/cache[6][145] ), .QN(n2970) );
  DFFRX1 \D_cache/cache_reg[7][145]  ( .D(\D_cache/n629 ), .CK(clk), .RN(n6126), .Q(\D_cache/cache[7][145] ), .QN(n1321) );
  DFFRX1 \D_cache/cache_reg[2][150]  ( .D(\D_cache/n594 ), .CK(clk), .RN(n6123), .Q(\D_cache/cache[2][150] ), .QN(n2092) );
  DFFRX1 \D_cache/cache_reg[3][150]  ( .D(\D_cache/n593 ), .CK(clk), .RN(n6123), .Q(\D_cache/cache[3][150] ), .QN(n466) );
  DFFRX1 \D_cache/cache_reg[2][147]  ( .D(\D_cache/n618 ), .CK(clk), .RN(n6125), .Q(\D_cache/cache[2][147] ), .QN(n2087) );
  DFFRX1 \D_cache/cache_reg[3][147]  ( .D(\D_cache/n617 ), .CK(clk), .RN(n6125), .Q(\D_cache/cache[3][147] ), .QN(n461) );
  DFFRX1 \D_cache/cache_reg[2][145]  ( .D(\D_cache/n634 ), .CK(clk), .RN(n6126), .Q(\D_cache/cache[2][145] ), .QN(n2960) );
  DFFRX1 \I_cache/cache_reg[4][139]  ( .D(n11729), .CK(clk), .RN(n6027), .Q(
        \I_cache/cache[4][139] ), .QN(n709) );
  DFFRX1 \I_cache/cache_reg[4][135]  ( .D(n11761), .CK(clk), .RN(n6030), .Q(
        \I_cache/cache[4][135] ), .QN(n2978) );
  DFFRX1 \I_cache/cache_reg[2][133]  ( .D(n11779), .CK(clk), .RN(n6031), .Q(
        \I_cache/cache[2][133] ), .QN(n2111) );
  DFFRX1 \I_cache/cache_reg[4][131]  ( .D(n11793), .CK(clk), .RN(n6032), .Q(
        \I_cache/cache[4][131] ), .QN(n2976) );
  DFFRX1 \I_cache/cache_reg[4][136]  ( .D(n11753), .CK(clk), .RN(n6029), .Q(
        \I_cache/cache[4][136] ), .QN(n2979) );
  DFFRX1 \I_cache/cache_reg[2][143]  ( .D(n11699), .CK(clk), .RN(n6024), .Q(
        \I_cache/cache[2][143] ), .QN(n2139) );
  DFFRX1 \I_cache/cache_reg[0][137]  ( .D(n11749), .CK(clk), .RN(n6029), .Q(
        \I_cache/cache[0][137] ), .QN(n985) );
  DFFRX1 \I_cache/cache_reg[4][128]  ( .D(n11817), .CK(clk), .RN(n6034), .Q(
        \I_cache/cache[4][128] ), .QN(n2924) );
  DFFRX1 \I_cache/cache_reg[4][133]  ( .D(n11777), .CK(clk), .RN(n6031), .Q(
        \I_cache/cache[4][133] ), .QN(n611) );
  DFFRX1 \I_cache/cache_reg[4][140]  ( .D(n11721), .CK(clk), .RN(n6026), .Q(
        \I_cache/cache[4][140] ), .QN(n708) );
  DFFRX1 \I_cache/cache_reg[6][143]  ( .D(n11695), .CK(clk), .RN(n6024), .Q(
        \I_cache/cache[6][143] ), .QN(n2968) );
  DFFRX1 \I_cache/cache_reg[1][143]  ( .D(n11700), .CK(clk), .RN(n6024), .Q(
        \I_cache/cache[1][143] ), .QN(n2230) );
  DFFRX1 \I_cache/cache_reg[5][137]  ( .D(n11744), .CK(clk), .RN(n6028), .Q(
        \I_cache/cache[5][137] ), .QN(n1325) );
  DFFRX1 \I_cache/cache_reg[6][133]  ( .D(n11775), .CK(clk), .RN(n6031), .Q(
        \I_cache/cache[6][133] ), .QN(n1330) );
  DFFRX1 \I_cache/cache_reg[1][133]  ( .D(n11780), .CK(clk), .RN(n6031), .Q(
        \I_cache/cache[1][133] ), .QN(n478) );
  DFFRX1 \I_cache/cache_reg[5][139]  ( .D(n11728), .CK(clk), .RN(n6027), .Q(
        \I_cache/cache[5][139] ), .QN(n2329) );
  DFFRX1 \I_cache/cache_reg[4][143]  ( .D(n11697), .CK(clk), .RN(n6024), .Q(
        \I_cache/cache[4][143] ), .QN(n2155) );
  DFFRX1 \I_cache/cache_reg[5][135]  ( .D(n11760), .CK(clk), .RN(n6029), .Q(
        \I_cache/cache[5][135] ), .QN(n1326) );
  DFFRX1 \I_cache/cache_reg[5][131]  ( .D(n11792), .CK(clk), .RN(n6032), .Q(
        \I_cache/cache[5][131] ), .QN(n1324) );
  DFFRX1 \I_cache/cache_reg[2][137]  ( .D(n11747), .CK(clk), .RN(n6028), .Q(
        \I_cache/cache[2][137] ), .QN(n1226) );
  DFFRX1 \I_cache/cache_reg[0][135]  ( .D(n11765), .CK(clk), .RN(n6030), .Q(
        \I_cache/cache[0][135] ), .QN(n981) );
  DFFRX1 \I_cache/cache_reg[0][131]  ( .D(n11797), .CK(clk), .RN(n6033), .Q(
        \I_cache/cache[0][131] ), .QN(n559) );
  DFFRX1 \I_cache/cache_reg[2][128]  ( .D(n11819), .CK(clk), .RN(n6034), .Q(
        \I_cache/cache[2][128] ), .QN(n535) );
  DFFRX1 \I_cache/cache_reg[5][136]  ( .D(n11752), .CK(clk), .RN(n6029), .Q(
        \I_cache/cache[5][136] ), .QN(n1327) );
  DFFRX1 \I_cache/cache_reg[3][143]  ( .D(n11698), .CK(clk), .RN(n6024), .Q(
        \I_cache/cache[3][143] ), .QN(n514) );
  DFFRX1 \I_cache/cache_reg[5][140]  ( .D(n11720), .CK(clk), .RN(n6026), .Q(
        \I_cache/cache[5][140] ), .QN(n2328) );
  DFFRX1 \I_cache/cache_reg[0][139]  ( .D(n11733), .CK(clk), .RN(n6027), .Q(
        \I_cache/cache[0][139] ), .QN(n2084) );
  DFFRX1 \I_cache/cache_reg[7][152]  ( .D(n11622), .CK(clk), .RN(n6018), .Q(
        \I_cache/cache[7][152] ), .QN(n530) );
  DFFRX1 \I_cache/cache_reg[4][134]  ( .D(n11769), .CK(clk), .RN(n6030), .Q(
        \I_cache/cache[4][134] ), .QN(n2975) );
  DFFRX1 \I_cache/cache_reg[0][136]  ( .D(n11757), .CK(clk), .RN(n6029), .Q(
        \I_cache/cache[0][136] ), .QN(n568) );
  DFFRX1 \I_cache/cache_reg[3][133]  ( .D(n11778), .CK(clk), .RN(n6031), .Q(
        \I_cache/cache[3][133] ), .QN(n485) );
  DFFRX1 \I_cache/cache_reg[2][135]  ( .D(n11763), .CK(clk), .RN(n6030), .Q(
        \I_cache/cache[2][135] ), .QN(n2117) );
  DFFRX1 \D_cache/cache_reg[5][149]  ( .D(\D_cache/n599 ), .CK(clk), .RN(n6123), .Q(\D_cache/cache[5][149] ), .QN(n2901) );
  DFFRX1 \I_cache/cache_reg[5][143]  ( .D(n11696), .CK(clk), .RN(n6024), .Q(
        \I_cache/cache[5][143] ), .QN(n531) );
  DFFRX1 \I_cache/cache_reg[4][132]  ( .D(n11785), .CK(clk), .RN(n6032), .Q(
        \I_cache/cache[4][132] ), .QN(n2974) );
  DFFRX1 \I_cache/cache_reg[2][131]  ( .D(n11795), .CK(clk), .RN(n6032), .Q(
        \I_cache/cache[2][131] ), .QN(n970) );
  DFFRX1 \I_cache/cache_reg[0][151]  ( .D(n11637), .CK(clk), .RN(n6019), .Q(
        \I_cache/cache[0][151] ), .QN(n534) );
  DFFRX1 \I_cache/cache_reg[2][139]  ( .D(n11731), .CK(clk), .RN(n6027), .Q(
        \I_cache/cache[2][139] ), .QN(n2067) );
  DFFRX1 \I_cache/cache_reg[6][137]  ( .D(n11743), .CK(clk), .RN(n6028), .Q(
        \I_cache/cache[6][137] ), .QN(n961) );
  DFFRX1 \I_cache/cache_reg[4][138]  ( .D(n11737), .CK(clk), .RN(n6028), .Q(
        \I_cache/cache[4][138] ), .QN(n2936) );
  DFFRX1 \I_cache/cache_reg[1][137]  ( .D(n11748), .CK(clk), .RN(n6028), .Q(
        \I_cache/cache[1][137] ), .QN(n2610) );
  DFFRX1 \I_cache/cache_reg[2][136]  ( .D(n11755), .CK(clk), .RN(n6029), .Q(
        \I_cache/cache[2][136] ), .QN(n960) );
  DFFRX1 \I_cache/cache_reg[7][133]  ( .D(n11774), .CK(clk), .RN(n6031), .Q(
        \I_cache/cache[7][133] ), .QN(n2983) );
  DFFRX1 \I_cache/cache_reg[5][133]  ( .D(n11776), .CK(clk), .RN(n6031), .Q(
        \I_cache/cache[5][133] ), .QN(n2229) );
  DFFRX1 \I_cache/cache_reg[5][134]  ( .D(n11768), .CK(clk), .RN(n6030), .Q(
        \I_cache/cache[5][134] ), .QN(n1323) );
  DFFRX1 \I_cache/cache_reg[7][143]  ( .D(n11694), .CK(clk), .RN(n6024), .Q(
        \I_cache/cache[7][143] ), .QN(n1320) );
  DFFRX1 \I_cache/cache_reg[4][151]  ( .D(n11633), .CK(clk), .RN(n6019), .Q(
        \I_cache/cache[4][151] ), .QN(n2923) );
  DFFRX1 \I_cache/cache_reg[0][140]  ( .D(n11725), .CK(clk), .RN(n6027), .Q(
        \I_cache/cache[0][140] ), .QN(n2085) );
  DFFRX1 \I_cache/cache_reg[5][132]  ( .D(n11784), .CK(clk), .RN(n6031), .Q(
        \I_cache/cache[5][132] ), .QN(n1322) );
  DFFRX1 \I_cache/cache_reg[4][142]  ( .D(n11705), .CK(clk), .RN(n6025), .Q(
        \I_cache/cache[4][142] ), .QN(n2980) );
  DFFRX1 \I_cache/cache_reg[6][135]  ( .D(n11759), .CK(clk), .RN(n6029), .Q(
        \I_cache/cache[6][135] ), .QN(n963) );
  DFFRX1 \I_cache/cache_reg[1][135]  ( .D(n11764), .CK(clk), .RN(n6030), .Q(
        \I_cache/cache[1][135] ), .QN(n2606) );
  DFFRX1 \I_cache/cache_reg[6][131]  ( .D(n11791), .CK(clk), .RN(n6032), .Q(
        \I_cache/cache[6][131] ), .QN(n2093) );
  DFFRX1 \I_cache/cache_reg[1][131]  ( .D(n11796), .CK(clk), .RN(n6032), .Q(
        \I_cache/cache[1][131] ), .QN(n2180) );
  DFFRX1 \I_cache/cache_reg[5][138]  ( .D(n11736), .CK(clk), .RN(n6027), .Q(
        \I_cache/cache[5][138] ), .QN(n4680) );
  DFFRX1 \I_cache/cache_reg[3][137]  ( .D(n11746), .CK(clk), .RN(n6028), .Q(
        \I_cache/cache[3][137] ), .QN(n2849) );
  DFFRX1 \I_cache/cache_reg[6][139]  ( .D(n11727), .CK(clk), .RN(n6027), .Q(
        \I_cache/cache[6][139] ), .QN(n2077) );
  DFFRX1 \I_cache/cache_reg[1][139]  ( .D(n11732), .CK(clk), .RN(n6027), .Q(
        \I_cache/cache[1][139] ), .QN(n458) );
  DFFRX1 \I_cache/cache_reg[2][140]  ( .D(n11723), .CK(clk), .RN(n6026), .Q(
        \I_cache/cache[2][140] ), .QN(n2061) );
  DFFRX1 \I_cache/cache_reg[6][136]  ( .D(n11751), .CK(clk), .RN(n6029), .Q(
        \I_cache/cache[6][136] ), .QN(n569) );
  DFFRX1 \I_cache/cache_reg[1][136]  ( .D(n11756), .CK(clk), .RN(n6029), .Q(
        \I_cache/cache[1][136] ), .QN(n2186) );
  DFFRX1 \I_cache/cache_reg[3][135]  ( .D(n11762), .CK(clk), .RN(n6030), .Q(
        \I_cache/cache[3][135] ), .QN(n491) );
  DFFRX1 \I_cache/cache_reg[3][131]  ( .D(n11794), .CK(clk), .RN(n6032), .Q(
        \I_cache/cache[3][131] ), .QN(n2595) );
  DFFRX1 \I_cache/cache_reg[4][145]  ( .D(n11681), .CK(clk), .RN(n6023), .Q(
        \I_cache/cache[4][145] ), .QN(n2922) );
  DFFRX1 \I_cache/cache_reg[5][128]  ( .D(n11816), .CK(clk), .RN(n6034), .Q(
        \I_cache/cache[5][128] ) );
  DFFRX1 \I_cache/cache_reg[3][139]  ( .D(n11730), .CK(clk), .RN(n6027), .Q(
        \I_cache/cache[3][139] ), .QN(n442) );
  DFFRX1 \I_cache/cache_reg[5][142]  ( .D(n11704), .CK(clk), .RN(n6025), .Q(
        \I_cache/cache[5][142] ), .QN(n1328) );
  DFFRX1 \I_cache/cache_reg[3][136]  ( .D(n11754), .CK(clk), .RN(n6029), .Q(
        \I_cache/cache[3][136] ), .QN(n2585) );
  DFFRX1 \I_cache/cache_reg[6][140]  ( .D(n11719), .CK(clk), .RN(n6026), .Q(
        \I_cache/cache[6][140] ), .QN(n2079) );
  DFFRX1 \I_cache/cache_reg[1][140]  ( .D(n11724), .CK(clk), .RN(n6026), .Q(
        \I_cache/cache[1][140] ), .QN(n459) );
  DFFRX1 \I_cache/cache_reg[7][137]  ( .D(n11742), .CK(clk), .RN(n6028), .Q(
        \I_cache/cache[7][137] ), .QN(n2586) );
  DFFRX1 \I_cache/cache_reg[0][134]  ( .D(n11773), .CK(clk), .RN(n6031), .Q(
        \I_cache/cache[0][134] ), .QN(n394) );
  DFFRX1 \I_cache/cache_reg[6][128]  ( .D(n11815), .CK(clk), .RN(n6034), .Q(
        \I_cache/cache[6][128] ), .QN(n536) );
  DFFRX1 \I_cache/cache_reg[2][151]  ( .D(n11635), .CK(clk), .RN(n6019), .Q(
        \I_cache/cache[2][151] ), .QN(n2972) );
  DFFRX1 \I_cache/cache_reg[1][128]  ( .D(n11820), .CK(clk), .RN(n6034), .Q(
        \I_cache/cache[1][128] ), .QN(n529) );
  DFFRX1 \I_cache/cache_reg[3][140]  ( .D(n11722), .CK(clk), .RN(n6026), .Q(
        \I_cache/cache[3][140] ), .QN(n436) );
  DFFRX1 \I_cache/cache_reg[0][145]  ( .D(n11685), .CK(clk), .RN(n6023), .Q(
        \I_cache/cache[0][145] ), .QN(n2971) );
  DFFRX1 \I_cache/cache_reg[7][135]  ( .D(n11758), .CK(clk), .RN(n6029), .Q(
        \I_cache/cache[7][135] ), .QN(n2588) );
  DFFRX1 \I_cache/cache_reg[7][131]  ( .D(n11790), .CK(clk), .RN(n6032), .Q(
        \I_cache/cache[7][131] ), .QN(n467) );
  DFFRX1 \I_cache/cache_reg[2][134]  ( .D(n11771), .CK(clk), .RN(n6030), .Q(
        \I_cache/cache[2][134] ), .QN(n590) );
  DFFRX1 \I_cache/cache_reg[7][139]  ( .D(n11726), .CK(clk), .RN(n6027), .Q(
        \I_cache/cache[7][139] ), .QN(n452) );
  DFFRX1 \I_cache/cache_reg[0][132]  ( .D(n11789), .CK(clk), .RN(n6032), .Q(
        \I_cache/cache[0][132] ), .QN(n2140) );
  DFFRX1 \I_cache/cache_reg[7][136]  ( .D(n11750), .CK(clk), .RN(n6029), .Q(
        \I_cache/cache[7][136] ), .QN(n2187) );
  DFFRX1 \I_cache/cache_reg[0][138]  ( .D(n11741), .CK(clk), .RN(n6028), .Q(
        \I_cache/cache[0][138] ), .QN(n376) );
  DFFRX1 \I_cache/cache_reg[1][134]  ( .D(n11772), .CK(clk), .RN(n6030), .Q(
        \I_cache/cache[1][134] ), .QN(n2030) );
  DFFRX1 \I_cache/cache_reg[2][132]  ( .D(n11787), .CK(clk), .RN(n6032), .Q(
        \I_cache/cache[2][132] ), .QN(n2122) );
  DFFRX1 \I_cache/cache_reg[6][134]  ( .D(n11767), .CK(clk), .RN(n6030), .Q(
        \I_cache/cache[6][134] ), .QN(n601) );
  DFFRX1 \I_cache/cache_reg[7][140]  ( .D(n11718), .CK(clk), .RN(n6026), .Q(
        \I_cache/cache[7][140] ), .QN(n454) );
  DFFRX1 \I_cache/cache_reg[5][151]  ( .D(n11632), .CK(clk), .RN(n6019), .Q(
        \I_cache/cache[5][151] ) );
  DFFRX1 \I_cache/cache_reg[2][138]  ( .D(n11739), .CK(clk), .RN(n6028), .Q(
        \I_cache/cache[2][138] ), .QN(n532) );
  DFFRX1 \I_cache/cache_reg[3][134]  ( .D(n11770), .CK(clk), .RN(n6030), .Q(
        \I_cache/cache[3][134] ), .QN(n2208) );
  DFFRX1 \I_cache/cache_reg[1][132]  ( .D(n11788), .CK(clk), .RN(n6032), .Q(
        \I_cache/cache[1][132] ), .QN(n515) );
  DFFRX1 \I_cache/cache_reg[6][132]  ( .D(n11783), .CK(clk), .RN(n6031), .Q(
        \I_cache/cache[6][132] ), .QN(n628) );
  DFFRX1 \I_cache/cache_reg[0][142]  ( .D(n11709), .CK(clk), .RN(n6025), .Q(
        \I_cache/cache[0][142] ), .QN(n533) );
  DFFRX1 \I_cache/cache_reg[3][128]  ( .D(n11818), .CK(clk), .RN(n6034), .Q(
        \I_cache/cache[3][128] ), .QN(n2964) );
  DFFRX1 \i_MIPS/ID_EX_reg[104]  ( .D(\i_MIPS/n417 ), .CK(clk), .RN(n6320), 
        .Q(\i_MIPS/ID_EX[104] ), .QN(n4772) );
  DFFRX1 \i_MIPS/ID_EX_reg[93]  ( .D(\i_MIPS/n428 ), .CK(clk), .RN(n6319), .Q(
        \i_MIPS/ID_EX[93] ), .QN(n4778) );
  DFFRX1 \i_MIPS/ID_EX_reg[89]  ( .D(\i_MIPS/n432 ), .CK(clk), .RN(n6318), .Q(
        \i_MIPS/ID_EX[89] ), .QN(n4781) );
  DFFRX1 \i_MIPS/ID_EX_reg[90]  ( .D(\i_MIPS/n431 ), .CK(clk), .RN(n6319), .Q(
        \i_MIPS/ID_EX[90] ), .QN(n4780) );
  DFFRX1 \i_MIPS/ID_EX_reg[92]  ( .D(\i_MIPS/n429 ), .CK(clk), .RN(n6319), .Q(
        \i_MIPS/ID_EX[92] ), .QN(n4779) );
  DFFRX1 \i_MIPS/ID_EX_reg[91]  ( .D(\i_MIPS/n430 ), .CK(clk), .RN(n6319), .Q(
        \i_MIPS/ID_EX[91] ), .QN(n4777) );
  DFFRX1 \D_cache/cache_reg[0][154]  ( .D(\D_cache/n564 ), .CK(clk), .RN(n6120), .Q(\D_cache/cache[0][154] ) );
  DFFRX1 \D_cache/cache_reg[1][154]  ( .D(\D_cache/n563 ), .CK(clk), .RN(n6120), .Q(\D_cache/cache[1][154] ) );
  DFFRX1 \D_cache/cache_reg[3][154]  ( .D(\D_cache/n561 ), .CK(clk), .RN(n6120), .Q(\D_cache/cache[3][154] ) );
  DFFRX1 \D_cache/cache_reg[4][154]  ( .D(\D_cache/n560 ), .CK(clk), .RN(n6120), .Q(\D_cache/cache[4][154] ), .QN(n3889) );
  DFFRX1 \D_cache/cache_reg[5][154]  ( .D(\D_cache/n559 ), .CK(clk), .RN(n6120), .Q(\D_cache/cache[5][154] ), .QN(n2012) );
  DFFRX1 \D_cache/cache_reg[6][154]  ( .D(\D_cache/n558 ), .CK(clk), .RN(n6120), .Q(\D_cache/cache[6][154] ) );
  DFFRX1 \D_cache/cache_reg[7][154]  ( .D(\D_cache/n557 ), .CK(clk), .RN(n6120), .Q(\D_cache/cache[7][154] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][0]  ( .D(\i_MIPS/Register/n148 ), 
        .CK(clk), .RN(n6306), .Q(\i_MIPS/Register/register[30][0] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][1]  ( .D(\i_MIPS/Register/n149 ), 
        .CK(clk), .RN(n6306), .Q(\i_MIPS/Register/register[30][1] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][2]  ( .D(\i_MIPS/Register/n150 ), 
        .CK(clk), .RN(n6306), .Q(\i_MIPS/Register/register[30][2] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][3]  ( .D(\i_MIPS/Register/n151 ), 
        .CK(clk), .RN(n6306), .Q(\i_MIPS/Register/register[30][3] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][4]  ( .D(\i_MIPS/Register/n152 ), 
        .CK(clk), .RN(n6305), .Q(\i_MIPS/Register/register[30][4] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][5]  ( .D(\i_MIPS/Register/n153 ), 
        .CK(clk), .RN(n6305), .Q(\i_MIPS/Register/register[30][5] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][6]  ( .D(\i_MIPS/Register/n154 ), 
        .CK(clk), .RN(n6305), .Q(\i_MIPS/Register/register[30][6] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][7]  ( .D(\i_MIPS/Register/n155 ), 
        .CK(clk), .RN(n6305), .Q(\i_MIPS/Register/register[30][7] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][8]  ( .D(\i_MIPS/Register/n156 ), 
        .CK(clk), .RN(n6305), .Q(\i_MIPS/Register/register[30][8] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][9]  ( .D(\i_MIPS/Register/n157 ), 
        .CK(clk), .RN(n6305), .Q(\i_MIPS/Register/register[30][9] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][10]  ( .D(\i_MIPS/Register/n158 ), 
        .CK(clk), .RN(n6305), .Q(\i_MIPS/Register/register[30][10] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][11]  ( .D(\i_MIPS/Register/n159 ), 
        .CK(clk), .RN(n6305), .Q(\i_MIPS/Register/register[30][11] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][12]  ( .D(\i_MIPS/Register/n160 ), 
        .CK(clk), .RN(n6305), .Q(\i_MIPS/Register/register[30][12] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][13]  ( .D(\i_MIPS/Register/n161 ), 
        .CK(clk), .RN(n6305), .Q(\i_MIPS/Register/register[30][13] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][15]  ( .D(\i_MIPS/Register/n163 ), 
        .CK(clk), .RN(n6305), .Q(\i_MIPS/Register/register[30][15] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][16]  ( .D(\i_MIPS/Register/n164 ), 
        .CK(clk), .RN(n6304), .Q(\i_MIPS/Register/register[30][16] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][17]  ( .D(\i_MIPS/Register/n165 ), 
        .CK(clk), .RN(n6304), .Q(\i_MIPS/Register/register[30][17] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][18]  ( .D(\i_MIPS/Register/n166 ), 
        .CK(clk), .RN(n6304), .Q(\i_MIPS/Register/register[30][18] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][19]  ( .D(\i_MIPS/Register/n167 ), 
        .CK(clk), .RN(n6304), .Q(\i_MIPS/Register/register[30][19] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][20]  ( .D(\i_MIPS/Register/n168 ), 
        .CK(clk), .RN(n6304), .Q(\i_MIPS/Register/register[30][20] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][21]  ( .D(\i_MIPS/Register/n169 ), 
        .CK(clk), .RN(n6304), .Q(\i_MIPS/Register/register[30][21] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][22]  ( .D(\i_MIPS/Register/n170 ), 
        .CK(clk), .RN(n6304), .Q(\i_MIPS/Register/register[30][22] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][23]  ( .D(\i_MIPS/Register/n171 ), 
        .CK(clk), .RN(n6304), .Q(\i_MIPS/Register/register[30][23] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][24]  ( .D(\i_MIPS/Register/n172 ), 
        .CK(clk), .RN(n6304), .Q(\i_MIPS/Register/register[30][24] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][25]  ( .D(\i_MIPS/Register/n173 ), 
        .CK(clk), .RN(n6304), .Q(\i_MIPS/Register/register[30][25] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][26]  ( .D(\i_MIPS/Register/n174 ), 
        .CK(clk), .RN(n6304), .Q(\i_MIPS/Register/register[30][26] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][27]  ( .D(\i_MIPS/Register/n175 ), 
        .CK(clk), .RN(n6304), .Q(\i_MIPS/Register/register[30][27] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][28]  ( .D(\i_MIPS/Register/n176 ), 
        .CK(clk), .RN(n6303), .Q(\i_MIPS/Register/register[30][28] ) );
  DFFRX1 \i_MIPS/Register/register_reg[30][29]  ( .D(\i_MIPS/Register/n177 ), 
        .CK(clk), .RN(n6303), .Q(\i_MIPS/Register/register[30][29] ) );
  DFFRX1 \i_MIPS/Register/register_reg[29][22]  ( .D(\i_MIPS/Register/n202 ), 
        .CK(clk), .RN(n6301), .Q(\i_MIPS/Register/register[29][22] ) );
  DFFRX1 \i_MIPS/Register/register_reg[27][22]  ( .D(\i_MIPS/Register/n266 ), 
        .CK(clk), .RN(n6296), .Q(\i_MIPS/Register/register[27][22] ) );
  DFFRX1 \i_MIPS/Register/register_reg[25][22]  ( .D(\i_MIPS/Register/n330 ), 
        .CK(clk), .RN(n6291), .Q(\i_MIPS/Register/register[25][22] ) );
  DFFRX1 \i_MIPS/Register/register_reg[15][22]  ( .D(\i_MIPS/Register/n650 ), 
        .CK(clk), .RN(n6264), .Q(\i_MIPS/Register/register[15][22] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][0]  ( .D(\i_MIPS/Register/n660 ), 
        .CK(clk), .RN(n6263), .Q(\i_MIPS/Register/register[14][0] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][1]  ( .D(\i_MIPS/Register/n661 ), 
        .CK(clk), .RN(n6263), .Q(\i_MIPS/Register/register[14][1] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][2]  ( .D(\i_MIPS/Register/n662 ), 
        .CK(clk), .RN(n6263), .Q(\i_MIPS/Register/register[14][2] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][3]  ( .D(\i_MIPS/Register/n663 ), 
        .CK(clk), .RN(n6263), .Q(\i_MIPS/Register/register[14][3] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][4]  ( .D(\i_MIPS/Register/n664 ), 
        .CK(clk), .RN(n6263), .Q(\i_MIPS/Register/register[14][4] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][5]  ( .D(\i_MIPS/Register/n665 ), 
        .CK(clk), .RN(n6263), .Q(\i_MIPS/Register/register[14][5] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][6]  ( .D(\i_MIPS/Register/n666 ), 
        .CK(clk), .RN(n6263), .Q(\i_MIPS/Register/register[14][6] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][7]  ( .D(\i_MIPS/Register/n667 ), 
        .CK(clk), .RN(n6263), .Q(\i_MIPS/Register/register[14][7] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][8]  ( .D(\i_MIPS/Register/n668 ), 
        .CK(clk), .RN(n6262), .Q(\i_MIPS/Register/register[14][8] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][9]  ( .D(\i_MIPS/Register/n669 ), 
        .CK(clk), .RN(n6262), .Q(\i_MIPS/Register/register[14][9] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][10]  ( .D(\i_MIPS/Register/n670 ), 
        .CK(clk), .RN(n6262), .Q(\i_MIPS/Register/register[14][10] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][11]  ( .D(\i_MIPS/Register/n671 ), 
        .CK(clk), .RN(n6262), .Q(\i_MIPS/Register/register[14][11] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][12]  ( .D(\i_MIPS/Register/n672 ), 
        .CK(clk), .RN(n6262), .Q(\i_MIPS/Register/register[14][12] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][13]  ( .D(\i_MIPS/Register/n673 ), 
        .CK(clk), .RN(n6262), .Q(\i_MIPS/Register/register[14][13] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][15]  ( .D(\i_MIPS/Register/n675 ), 
        .CK(clk), .RN(n6262), .Q(\i_MIPS/Register/register[14][15] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][16]  ( .D(\i_MIPS/Register/n676 ), 
        .CK(clk), .RN(n6262), .Q(\i_MIPS/Register/register[14][16] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][17]  ( .D(\i_MIPS/Register/n677 ), 
        .CK(clk), .RN(n6262), .Q(\i_MIPS/Register/register[14][17] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][18]  ( .D(\i_MIPS/Register/n678 ), 
        .CK(clk), .RN(n6262), .Q(\i_MIPS/Register/register[14][18] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][19]  ( .D(\i_MIPS/Register/n679 ), 
        .CK(clk), .RN(n6262), .Q(\i_MIPS/Register/register[14][19] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][20]  ( .D(\i_MIPS/Register/n680 ), 
        .CK(clk), .RN(n6261), .Q(\i_MIPS/Register/register[14][20] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][21]  ( .D(\i_MIPS/Register/n681 ), 
        .CK(clk), .RN(n6261), .Q(\i_MIPS/Register/register[14][21] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][22]  ( .D(\i_MIPS/Register/n682 ), 
        .CK(clk), .RN(n6261), .Q(\i_MIPS/Register/register[14][22] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][23]  ( .D(\i_MIPS/Register/n683 ), 
        .CK(clk), .RN(n6261), .Q(\i_MIPS/Register/register[14][23] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][24]  ( .D(\i_MIPS/Register/n684 ), 
        .CK(clk), .RN(n6261), .Q(\i_MIPS/Register/register[14][24] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][25]  ( .D(\i_MIPS/Register/n685 ), 
        .CK(clk), .RN(n6261), .Q(\i_MIPS/Register/register[14][25] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][26]  ( .D(\i_MIPS/Register/n686 ), 
        .CK(clk), .RN(n6261), .Q(\i_MIPS/Register/register[14][26] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][27]  ( .D(\i_MIPS/Register/n687 ), 
        .CK(clk), .RN(n6261), .Q(\i_MIPS/Register/register[14][27] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][28]  ( .D(\i_MIPS/Register/n688 ), 
        .CK(clk), .RN(n6261), .Q(\i_MIPS/Register/register[14][28] ) );
  DFFRX1 \i_MIPS/Register/register_reg[14][29]  ( .D(\i_MIPS/Register/n689 ), 
        .CK(clk), .RN(n6261), .Q(\i_MIPS/Register/register[14][29] ) );
  DFFRX1 \i_MIPS/Register/register_reg[13][22]  ( .D(\i_MIPS/Register/n714 ), 
        .CK(clk), .RN(n6259), .Q(\i_MIPS/Register/register[13][22] ) );
  DFFRX1 \i_MIPS/Register/register_reg[11][22]  ( .D(\i_MIPS/Register/n778 ), 
        .CK(clk), .RN(n6253), .Q(\i_MIPS/Register/register[11][22] ) );
  DFFRX1 \i_MIPS/Register/register_reg[9][22]  ( .D(\i_MIPS/Register/n842 ), 
        .CK(clk), .RN(n6248), .Q(\i_MIPS/Register/register[9][22] ) );
  DFFRX1 \i_MIPS/Register/register_reg[23][22]  ( .D(\i_MIPS/Register/n394 ), 
        .CK(clk), .RN(n6285), .Q(\i_MIPS/Register/register[23][22] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][0]  ( .D(\i_MIPS/Register/n404 ), 
        .CK(clk), .RN(n6284), .Q(\i_MIPS/Register/register[22][0] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][1]  ( .D(\i_MIPS/Register/n405 ), 
        .CK(clk), .RN(n6284), .Q(\i_MIPS/Register/register[22][1] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][2]  ( .D(\i_MIPS/Register/n406 ), 
        .CK(clk), .RN(n6284), .Q(\i_MIPS/Register/register[22][2] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][3]  ( .D(\i_MIPS/Register/n407 ), 
        .CK(clk), .RN(n6284), .Q(\i_MIPS/Register/register[22][3] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][4]  ( .D(\i_MIPS/Register/n408 ), 
        .CK(clk), .RN(n6284), .Q(\i_MIPS/Register/register[22][4] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][5]  ( .D(\i_MIPS/Register/n409 ), 
        .CK(clk), .RN(n6284), .Q(\i_MIPS/Register/register[22][5] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][6]  ( .D(\i_MIPS/Register/n410 ), 
        .CK(clk), .RN(n6284), .Q(\i_MIPS/Register/register[22][6] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][7]  ( .D(\i_MIPS/Register/n411 ), 
        .CK(clk), .RN(n6284), .Q(\i_MIPS/Register/register[22][7] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][8]  ( .D(\i_MIPS/Register/n412 ), 
        .CK(clk), .RN(n6284), .Q(\i_MIPS/Register/register[22][8] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][9]  ( .D(\i_MIPS/Register/n413 ), 
        .CK(clk), .RN(n6284), .Q(\i_MIPS/Register/register[22][9] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][10]  ( .D(\i_MIPS/Register/n414 ), 
        .CK(clk), .RN(n6284), .Q(\i_MIPS/Register/register[22][10] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][11]  ( .D(\i_MIPS/Register/n415 ), 
        .CK(clk), .RN(n6284), .Q(\i_MIPS/Register/register[22][11] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][12]  ( .D(\i_MIPS/Register/n416 ), 
        .CK(clk), .RN(n6283), .Q(\i_MIPS/Register/register[22][12] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][13]  ( .D(\i_MIPS/Register/n417 ), 
        .CK(clk), .RN(n6283), .Q(\i_MIPS/Register/register[22][13] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][16]  ( .D(\i_MIPS/Register/n420 ), 
        .CK(clk), .RN(n6283), .Q(\i_MIPS/Register/register[22][16] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][17]  ( .D(\i_MIPS/Register/n421 ), 
        .CK(clk), .RN(n6283), .Q(\i_MIPS/Register/register[22][17] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][18]  ( .D(\i_MIPS/Register/n422 ), 
        .CK(clk), .RN(n6283), .Q(\i_MIPS/Register/register[22][18] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][19]  ( .D(\i_MIPS/Register/n423 ), 
        .CK(clk), .RN(n6283), .Q(\i_MIPS/Register/register[22][19] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][20]  ( .D(\i_MIPS/Register/n424 ), 
        .CK(clk), .RN(n6283), .Q(\i_MIPS/Register/register[22][20] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][21]  ( .D(\i_MIPS/Register/n425 ), 
        .CK(clk), .RN(n6283), .Q(\i_MIPS/Register/register[22][21] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][22]  ( .D(\i_MIPS/Register/n426 ), 
        .CK(clk), .RN(n6283), .Q(\i_MIPS/Register/register[22][22] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][23]  ( .D(\i_MIPS/Register/n427 ), 
        .CK(clk), .RN(n6283), .Q(\i_MIPS/Register/register[22][23] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][24]  ( .D(\i_MIPS/Register/n428 ), 
        .CK(clk), .RN(n6282), .Q(\i_MIPS/Register/register[22][24] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][26]  ( .D(\i_MIPS/Register/n430 ), 
        .CK(clk), .RN(n6282), .Q(\i_MIPS/Register/register[22][26] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][27]  ( .D(\i_MIPS/Register/n431 ), 
        .CK(clk), .RN(n6282), .Q(\i_MIPS/Register/register[22][27] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][28]  ( .D(\i_MIPS/Register/n432 ), 
        .CK(clk), .RN(n6282), .Q(\i_MIPS/Register/register[22][28] ) );
  DFFRX1 \i_MIPS/Register/register_reg[22][29]  ( .D(\i_MIPS/Register/n433 ), 
        .CK(clk), .RN(n6282), .Q(\i_MIPS/Register/register[22][29] ) );
  DFFRX1 \i_MIPS/Register/register_reg[7][22]  ( .D(\i_MIPS/Register/n906 ), 
        .CK(clk), .RN(n6243), .Q(\i_MIPS/Register/register[7][22] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][0]  ( .D(\i_MIPS/Register/n916 ), 
        .CK(clk), .RN(n6242), .Q(\i_MIPS/Register/register[6][0] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][1]  ( .D(\i_MIPS/Register/n917 ), 
        .CK(clk), .RN(n6242), .Q(\i_MIPS/Register/register[6][1] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][2]  ( .D(\i_MIPS/Register/n918 ), 
        .CK(clk), .RN(n6242), .Q(\i_MIPS/Register/register[6][2] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][3]  ( .D(\i_MIPS/Register/n919 ), 
        .CK(clk), .RN(n6242), .Q(\i_MIPS/Register/register[6][3] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][4]  ( .D(\i_MIPS/Register/n920 ), 
        .CK(clk), .RN(n6241), .Q(\i_MIPS/Register/register[6][4] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][5]  ( .D(\i_MIPS/Register/n921 ), 
        .CK(clk), .RN(n6241), .Q(\i_MIPS/Register/register[6][5] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][6]  ( .D(\i_MIPS/Register/n922 ), 
        .CK(clk), .RN(n6241), .Q(\i_MIPS/Register/register[6][6] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][7]  ( .D(\i_MIPS/Register/n923 ), 
        .CK(clk), .RN(n6241), .Q(\i_MIPS/Register/register[6][7] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][8]  ( .D(\i_MIPS/Register/n924 ), 
        .CK(clk), .RN(n6241), .Q(\i_MIPS/Register/register[6][8] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][9]  ( .D(\i_MIPS/Register/n925 ), 
        .CK(clk), .RN(n6241), .Q(\i_MIPS/Register/register[6][9] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][10]  ( .D(\i_MIPS/Register/n926 ), 
        .CK(clk), .RN(n6241), .Q(\i_MIPS/Register/register[6][10] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][11]  ( .D(\i_MIPS/Register/n927 ), 
        .CK(clk), .RN(n6241), .Q(\i_MIPS/Register/register[6][11] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][12]  ( .D(\i_MIPS/Register/n928 ), 
        .CK(clk), .RN(n6241), .Q(\i_MIPS/Register/register[6][12] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][13]  ( .D(\i_MIPS/Register/n929 ), 
        .CK(clk), .RN(n6241), .Q(\i_MIPS/Register/register[6][13] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][16]  ( .D(\i_MIPS/Register/n932 ), 
        .CK(clk), .RN(n6240), .Q(\i_MIPS/Register/register[6][16] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][17]  ( .D(\i_MIPS/Register/n933 ), 
        .CK(clk), .RN(n6240), .Q(\i_MIPS/Register/register[6][17] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][18]  ( .D(\i_MIPS/Register/n934 ), 
        .CK(clk), .RN(n6240), .Q(\i_MIPS/Register/register[6][18] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][19]  ( .D(\i_MIPS/Register/n935 ), 
        .CK(clk), .RN(n6240), .Q(\i_MIPS/Register/register[6][19] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][20]  ( .D(\i_MIPS/Register/n936 ), 
        .CK(clk), .RN(n6240), .Q(\i_MIPS/Register/register[6][20] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][21]  ( .D(\i_MIPS/Register/n937 ), 
        .CK(clk), .RN(n6240), .Q(\i_MIPS/Register/register[6][21] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][22]  ( .D(\i_MIPS/Register/n938 ), 
        .CK(clk), .RN(n6240), .Q(\i_MIPS/Register/register[6][22] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][23]  ( .D(\i_MIPS/Register/n939 ), 
        .CK(clk), .RN(n6240), .Q(\i_MIPS/Register/register[6][23] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][24]  ( .D(\i_MIPS/Register/n940 ), 
        .CK(clk), .RN(n6240), .Q(\i_MIPS/Register/register[6][24] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][26]  ( .D(\i_MIPS/Register/n942 ), 
        .CK(clk), .RN(n6240), .Q(\i_MIPS/Register/register[6][26] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][27]  ( .D(\i_MIPS/Register/n943 ), 
        .CK(clk), .RN(n6240), .Q(\i_MIPS/Register/register[6][27] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][28]  ( .D(\i_MIPS/Register/n944 ), 
        .CK(clk), .RN(n6239), .Q(\i_MIPS/Register/register[6][28] ) );
  DFFRX1 \i_MIPS/Register/register_reg[6][29]  ( .D(\i_MIPS/Register/n945 ), 
        .CK(clk), .RN(n6239), .Q(\i_MIPS/Register/register[6][29] ) );
  DFFRX1 \i_MIPS/Register/register_reg[29][0]  ( .D(\i_MIPS/Register/n180 ), 
        .CK(clk), .RN(n6303), .Q(\i_MIPS/Register/register[29][0] ), .QN(n272)
         );
  DFFRX1 \i_MIPS/Register/register_reg[29][1]  ( .D(\i_MIPS/Register/n181 ), 
        .CK(clk), .RN(n6303), .Q(\i_MIPS/Register/register[29][1] ), .QN(n859)
         );
  DFFRX1 \i_MIPS/Register/register_reg[29][2]  ( .D(\i_MIPS/Register/n182 ), 
        .CK(clk), .RN(n6303), .Q(\i_MIPS/Register/register[29][2] ), .QN(n887)
         );
  DFFRX1 \i_MIPS/Register/register_reg[29][3]  ( .D(\i_MIPS/Register/n183 ), 
        .CK(clk), .RN(n6303), .Q(\i_MIPS/Register/register[29][3] ), .QN(n792)
         );
  DFFRX1 \i_MIPS/Register/register_reg[29][4]  ( .D(\i_MIPS/Register/n184 ), 
        .CK(clk), .RN(n6303), .Q(\i_MIPS/Register/register[29][4] ), .QN(n875)
         );
  DFFRX1 \i_MIPS/Register/register_reg[29][5]  ( .D(\i_MIPS/Register/n185 ), 
        .CK(clk), .RN(n6303), .Q(\i_MIPS/Register/register[29][5] ), .QN(n782)
         );
  DFFRX1 \i_MIPS/Register/register_reg[29][6]  ( .D(\i_MIPS/Register/n186 ), 
        .CK(clk), .RN(n6303), .Q(\i_MIPS/Register/register[29][6] ), .QN(n884)
         );
  DFFRX1 \i_MIPS/Register/register_reg[29][7]  ( .D(\i_MIPS/Register/n187 ), 
        .CK(clk), .RN(n6303), .Q(\i_MIPS/Register/register[29][7] ), .QN(n880)
         );
  DFFRX1 \i_MIPS/Register/register_reg[29][8]  ( .D(\i_MIPS/Register/n188 ), 
        .CK(clk), .RN(n6302), .Q(\i_MIPS/Register/register[29][8] ), .QN(n867)
         );
  DFFRX1 \i_MIPS/Register/register_reg[29][9]  ( .D(\i_MIPS/Register/n189 ), 
        .CK(clk), .RN(n6302), .Q(\i_MIPS/Register/register[29][9] ), .QN(n384)
         );
  DFFRX1 \i_MIPS/Register/register_reg[29][10]  ( .D(\i_MIPS/Register/n190 ), 
        .CK(clk), .RN(n6302), .Q(\i_MIPS/Register/register[29][10] ), .QN(n380) );
  DFFRX1 \i_MIPS/Register/register_reg[29][11]  ( .D(\i_MIPS/Register/n191 ), 
        .CK(clk), .RN(n6302), .Q(\i_MIPS/Register/register[29][11] ), .QN(n294) );
  DFFRX1 \i_MIPS/Register/register_reg[29][12]  ( .D(\i_MIPS/Register/n192 ), 
        .CK(clk), .RN(n6302), .Q(\i_MIPS/Register/register[29][12] ), .QN(n860) );
  DFFRX1 \i_MIPS/Register/register_reg[29][13]  ( .D(\i_MIPS/Register/n193 ), 
        .CK(clk), .RN(n6302), .Q(\i_MIPS/Register/register[29][13] ), .QN(n804) );
  DFFRX1 \i_MIPS/Register/register_reg[29][15]  ( .D(\i_MIPS/Register/n195 ), 
        .CK(clk), .RN(n6302), .Q(\i_MIPS/Register/register[29][15] ), .QN(n889) );
  DFFRX1 \i_MIPS/Register/register_reg[29][16]  ( .D(\i_MIPS/Register/n196 ), 
        .CK(clk), .RN(n6302), .Q(\i_MIPS/Register/register[29][16] ), .QN(n275) );
  DFFRX1 \i_MIPS/Register/register_reg[29][17]  ( .D(\i_MIPS/Register/n197 ), 
        .CK(clk), .RN(n6302), .Q(\i_MIPS/Register/register[29][17] ), .QN(n855) );
  DFFRX1 \i_MIPS/Register/register_reg[29][18]  ( .D(\i_MIPS/Register/n198 ), 
        .CK(clk), .RN(n6302), .Q(\i_MIPS/Register/register[29][18] ), .QN(n293) );
  DFFRX1 \i_MIPS/Register/register_reg[29][19]  ( .D(\i_MIPS/Register/n199 ), 
        .CK(clk), .RN(n6302), .Q(\i_MIPS/Register/register[29][19] ), .QN(n863) );
  DFFRX1 \i_MIPS/Register/register_reg[29][20]  ( .D(\i_MIPS/Register/n200 ), 
        .CK(clk), .RN(n6301), .Q(\i_MIPS/Register/register[29][20] ), .QN(n295) );
  DFFRX1 \i_MIPS/Register/register_reg[29][21]  ( .D(\i_MIPS/Register/n201 ), 
        .CK(clk), .RN(n6301), .Q(\i_MIPS/Register/register[29][21] ), .QN(n297) );
  DFFRX1 \i_MIPS/Register/register_reg[29][23]  ( .D(\i_MIPS/Register/n203 ), 
        .CK(clk), .RN(n6301), .Q(\i_MIPS/Register/register[29][23] ), .QN(n812) );
  DFFRX1 \i_MIPS/Register/register_reg[29][24]  ( .D(\i_MIPS/Register/n204 ), 
        .CK(clk), .RN(n6301), .Q(\i_MIPS/Register/register[29][24] ), .QN(n775) );
  DFFRX1 \i_MIPS/Register/register_reg[29][25]  ( .D(\i_MIPS/Register/n205 ), 
        .CK(clk), .RN(n6301), .Q(\i_MIPS/Register/register[29][25] ), .QN(n893) );
  DFFRX1 \i_MIPS/Register/register_reg[29][26]  ( .D(\i_MIPS/Register/n206 ), 
        .CK(clk), .RN(n6301), .Q(\i_MIPS/Register/register[29][26] ), .QN(n870) );
  DFFRX1 \i_MIPS/Register/register_reg[29][27]  ( .D(\i_MIPS/Register/n207 ), 
        .CK(clk), .RN(n6301), .Q(\i_MIPS/Register/register[29][27] ), .QN(n894) );
  DFFRX1 \i_MIPS/Register/register_reg[29][28]  ( .D(\i_MIPS/Register/n208 ), 
        .CK(clk), .RN(n6301), .Q(\i_MIPS/Register/register[29][28] ), .QN(n885) );
  DFFRX1 \i_MIPS/Register/register_reg[29][29]  ( .D(\i_MIPS/Register/n209 ), 
        .CK(clk), .RN(n6301), .Q(\i_MIPS/Register/register[29][29] ), .QN(n820) );
  DFFRX1 \i_MIPS/Register/register_reg[28][0]  ( .D(\i_MIPS/Register/n212 ), 
        .CK(clk), .RN(n6300), .Q(\i_MIPS/Register/register[28][0] ), .QN(n830)
         );
  DFFRX1 \i_MIPS/Register/register_reg[28][1]  ( .D(\i_MIPS/Register/n213 ), 
        .CK(clk), .RN(n6300), .Q(\i_MIPS/Register/register[28][1] ), .QN(n285)
         );
  DFFRX1 \i_MIPS/Register/register_reg[28][3]  ( .D(\i_MIPS/Register/n215 ), 
        .CK(clk), .RN(n6300), .Q(\i_MIPS/Register/register[28][3] ), .QN(n266)
         );
  DFFRX1 \i_MIPS/Register/register_reg[28][4]  ( .D(\i_MIPS/Register/n216 ), 
        .CK(clk), .RN(n6300), .Q(\i_MIPS/Register/register[28][4] ), .QN(n283)
         );
  DFFRX1 \i_MIPS/Register/register_reg[28][5]  ( .D(\i_MIPS/Register/n217 ), 
        .CK(clk), .RN(n6300), .Q(\i_MIPS/Register/register[28][5] ), .QN(n263)
         );
  DFFRX1 \i_MIPS/Register/register_reg[28][6]  ( .D(\i_MIPS/Register/n218 ), 
        .CK(clk), .RN(n6300), .Q(\i_MIPS/Register/register[28][6] ), .QN(n897)
         );
  DFFRX1 \i_MIPS/Register/register_reg[28][7]  ( .D(\i_MIPS/Register/n219 ), 
        .CK(clk), .RN(n6300), .Q(\i_MIPS/Register/register[28][7] ), .QN(n896)
         );
  DFFRX1 \i_MIPS/Register/register_reg[28][8]  ( .D(\i_MIPS/Register/n220 ), 
        .CK(clk), .RN(n6300), .Q(\i_MIPS/Register/register[28][8] ), .QN(n832)
         );
  DFFRX1 \i_MIPS/Register/register_reg[28][9]  ( .D(\i_MIPS/Register/n221 ), 
        .CK(clk), .RN(n6300), .Q(\i_MIPS/Register/register[28][9] ), .QN(n562)
         );
  DFFRX1 \i_MIPS/Register/register_reg[28][10]  ( .D(\i_MIPS/Register/n222 ), 
        .CK(clk), .RN(n6300), .Q(\i_MIPS/Register/register[28][10] ), .QN(n723) );
  DFFRX1 \i_MIPS/Register/register_reg[28][11]  ( .D(\i_MIPS/Register/n223 ), 
        .CK(clk), .RN(n6300), .Q(\i_MIPS/Register/register[28][11] ), .QN(n827) );
  DFFRX1 \i_MIPS/Register/register_reg[28][12]  ( .D(\i_MIPS/Register/n224 ), 
        .CK(clk), .RN(n6299), .Q(\i_MIPS/Register/register[28][12] ), .QN(n831) );
  DFFRX1 \i_MIPS/Register/register_reg[28][13]  ( .D(\i_MIPS/Register/n225 ), 
        .CK(clk), .RN(n6299), .Q(\i_MIPS/Register/register[28][13] ), .QN(n853) );
  DFFRX1 \i_MIPS/Register/register_reg[28][16]  ( .D(\i_MIPS/Register/n228 ), 
        .CK(clk), .RN(n6299), .Q(\i_MIPS/Register/register[28][16] ), .QN(n829) );
  DFFRX1 \i_MIPS/Register/register_reg[28][17]  ( .D(\i_MIPS/Register/n229 ), 
        .CK(clk), .RN(n6299), .Q(\i_MIPS/Register/register[28][17] ), .QN(n262) );
  DFFRX1 \i_MIPS/Register/register_reg[28][18]  ( .D(\i_MIPS/Register/n230 ), 
        .CK(clk), .RN(n6299), .Q(\i_MIPS/Register/register[28][18] ), .QN(n415) );
  DFFRX1 \i_MIPS/Register/register_reg[28][19]  ( .D(\i_MIPS/Register/n231 ), 
        .CK(clk), .RN(n6299), .Q(\i_MIPS/Register/register[28][19] ), .QN(n828) );
  DFFRX1 \i_MIPS/Register/register_reg[28][20]  ( .D(\i_MIPS/Register/n232 ), 
        .CK(clk), .RN(n6299), .Q(\i_MIPS/Register/register[28][20] ), .QN(n895) );
  DFFRX1 \i_MIPS/Register/register_reg[28][21]  ( .D(\i_MIPS/Register/n233 ), 
        .CK(clk), .RN(n6299), .Q(\i_MIPS/Register/register[28][21] ), .QN(n424) );
  DFFRX1 \i_MIPS/Register/register_reg[28][23]  ( .D(\i_MIPS/Register/n235 ), 
        .CK(clk), .RN(n6299), .Q(\i_MIPS/Register/register[28][23] ), .QN(n284) );
  DFFRX1 \i_MIPS/Register/register_reg[28][26]  ( .D(\i_MIPS/Register/n238 ), 
        .CK(clk), .RN(n6298), .Q(\i_MIPS/Register/register[28][26] ), .QN(n898) );
  DFFRX1 \i_MIPS/Register/register_reg[28][27]  ( .D(\i_MIPS/Register/n239 ), 
        .CK(clk), .RN(n6298), .Q(\i_MIPS/Register/register[28][27] ), .QN(n833) );
  DFFRX1 \i_MIPS/Register/register_reg[27][0]  ( .D(\i_MIPS/Register/n244 ), 
        .CK(clk), .RN(n6298), .Q(\i_MIPS/Register/register[27][0] ), .QN(n783)
         );
  DFFRX1 \i_MIPS/Register/register_reg[27][1]  ( .D(\i_MIPS/Register/n245 ), 
        .CK(clk), .RN(n6298), .Q(\i_MIPS/Register/register[27][1] ), .QN(n776)
         );
  DFFRX1 \i_MIPS/Register/register_reg[27][2]  ( .D(\i_MIPS/Register/n246 ), 
        .CK(clk), .RN(n6298), .Q(\i_MIPS/Register/register[27][2] ), .QN(n816)
         );
  DFFRX1 \i_MIPS/Register/register_reg[27][3]  ( .D(\i_MIPS/Register/n247 ), 
        .CK(clk), .RN(n6298), .Q(\i_MIPS/Register/register[27][3] ), .QN(n791)
         );
  DFFRX1 \i_MIPS/Register/register_reg[27][4]  ( .D(\i_MIPS/Register/n248 ), 
        .CK(clk), .RN(n6297), .Q(\i_MIPS/Register/register[27][4] ), .QN(n874)
         );
  DFFRX1 \i_MIPS/Register/register_reg[27][5]  ( .D(\i_MIPS/Register/n249 ), 
        .CK(clk), .RN(n6297), .Q(\i_MIPS/Register/register[27][5] ), .QN(n781)
         );
  DFFRX1 \i_MIPS/Register/register_reg[27][6]  ( .D(\i_MIPS/Register/n250 ), 
        .CK(clk), .RN(n6297), .Q(\i_MIPS/Register/register[27][6] ), .QN(n883)
         );
  DFFRX1 \i_MIPS/Register/register_reg[27][7]  ( .D(\i_MIPS/Register/n251 ), 
        .CK(clk), .RN(n6297), .Q(\i_MIPS/Register/register[27][7] ), .QN(n879)
         );
  DFFRX1 \i_MIPS/Register/register_reg[27][8]  ( .D(\i_MIPS/Register/n252 ), 
        .CK(clk), .RN(n6297), .Q(\i_MIPS/Register/register[27][8] ), .QN(n279)
         );
  DFFRX1 \i_MIPS/Register/register_reg[27][9]  ( .D(\i_MIPS/Register/n253 ), 
        .CK(clk), .RN(n6297), .Q(\i_MIPS/Register/register[27][9] ), .QN(n249)
         );
  DFFRX1 \i_MIPS/Register/register_reg[27][10]  ( .D(\i_MIPS/Register/n254 ), 
        .CK(clk), .RN(n6297), .Q(\i_MIPS/Register/register[27][10] ), .QN(n379) );
  DFFRX1 \i_MIPS/Register/register_reg[27][11]  ( .D(\i_MIPS/Register/n255 ), 
        .CK(clk), .RN(n6297), .Q(\i_MIPS/Register/register[27][11] ), .QN(n796) );
  DFFRX1 \i_MIPS/Register/register_reg[27][12]  ( .D(\i_MIPS/Register/n256 ), 
        .CK(clk), .RN(n6297), .Q(\i_MIPS/Register/register[27][12] ), .QN(n270) );
  DFFRX1 \i_MIPS/Register/register_reg[27][13]  ( .D(\i_MIPS/Register/n257 ), 
        .CK(clk), .RN(n6297), .Q(\i_MIPS/Register/register[27][13] ), .QN(n281) );
  DFFRX1 \i_MIPS/Register/register_reg[27][15]  ( .D(\i_MIPS/Register/n259 ), 
        .CK(clk), .RN(n6297), .Q(\i_MIPS/Register/register[27][15] ), .QN(n888) );
  DFFRX1 \i_MIPS/Register/register_reg[27][16]  ( .D(\i_MIPS/Register/n260 ), 
        .CK(clk), .RN(n6296), .Q(\i_MIPS/Register/register[27][16] ), .QN(n797) );
  DFFRX1 \i_MIPS/Register/register_reg[27][17]  ( .D(\i_MIPS/Register/n261 ), 
        .CK(clk), .RN(n6296), .Q(\i_MIPS/Register/register[27][17] ), .QN(n854) );
  DFFRX1 \i_MIPS/Register/register_reg[27][18]  ( .D(\i_MIPS/Register/n262 ), 
        .CK(clk), .RN(n6296), .Q(\i_MIPS/Register/register[27][18] ), .QN(n780) );
  DFFRX1 \i_MIPS/Register/register_reg[27][19]  ( .D(\i_MIPS/Register/n263 ), 
        .CK(clk), .RN(n6296), .Q(\i_MIPS/Register/register[27][19] ), .QN(n278) );
  DFFRX1 \i_MIPS/Register/register_reg[27][20]  ( .D(\i_MIPS/Register/n264 ), 
        .CK(clk), .RN(n6296), .Q(\i_MIPS/Register/register[27][20] ), .QN(n862) );
  DFFRX1 \i_MIPS/Register/register_reg[27][21]  ( .D(\i_MIPS/Register/n265 ), 
        .CK(clk), .RN(n6296), .Q(\i_MIPS/Register/register[27][21] ), .QN(n802) );
  DFFRX1 \i_MIPS/Register/register_reg[27][23]  ( .D(\i_MIPS/Register/n267 ), 
        .CK(clk), .RN(n6296), .Q(\i_MIPS/Register/register[27][23] ), .QN(n811) );
  DFFRX1 \i_MIPS/Register/register_reg[27][24]  ( .D(\i_MIPS/Register/n268 ), 
        .CK(clk), .RN(n6296), .Q(\i_MIPS/Register/register[27][24] ), .QN(n774) );
  DFFRX1 \i_MIPS/Register/register_reg[27][25]  ( .D(\i_MIPS/Register/n269 ), 
        .CK(clk), .RN(n6296), .Q(\i_MIPS/Register/register[27][25] ), .QN(n822) );
  DFFRX1 \i_MIPS/Register/register_reg[27][26]  ( .D(\i_MIPS/Register/n270 ), 
        .CK(clk), .RN(n6296), .Q(\i_MIPS/Register/register[27][26] ), .QN(n869) );
  DFFRX1 \i_MIPS/Register/register_reg[27][27]  ( .D(\i_MIPS/Register/n271 ), 
        .CK(clk), .RN(n6296), .Q(\i_MIPS/Register/register[27][27] ), .QN(n823) );
  DFFRX1 \i_MIPS/Register/register_reg[27][28]  ( .D(\i_MIPS/Register/n272 ), 
        .CK(clk), .RN(n6295), .Q(\i_MIPS/Register/register[27][28] ), .QN(n809) );
  DFFRX1 \i_MIPS/Register/register_reg[27][29]  ( .D(\i_MIPS/Register/n273 ), 
        .CK(clk), .RN(n6295), .Q(\i_MIPS/Register/register[27][29] ), .QN(n387) );
  DFFRX1 \i_MIPS/Register/register_reg[25][0]  ( .D(\i_MIPS/Register/n308 ), 
        .CK(clk), .RN(n6292), .Q(\i_MIPS/Register/register[25][0] ), .QN(n420)
         );
  DFFRX1 \i_MIPS/Register/register_reg[25][1]  ( .D(\i_MIPS/Register/n309 ), 
        .CK(clk), .RN(n6292), .Q(\i_MIPS/Register/register[25][1] ), .QN(n836)
         );
  DFFRX1 \i_MIPS/Register/register_reg[25][2]  ( .D(\i_MIPS/Register/n310 ), 
        .CK(clk), .RN(n6292), .Q(\i_MIPS/Register/register[25][2] ), .QN(n200)
         );
  DFFRX1 \i_MIPS/Register/register_reg[25][3]  ( .D(\i_MIPS/Register/n311 ), 
        .CK(clk), .RN(n6292), .Q(\i_MIPS/Register/register[25][3] ), .QN(n734)
         );
  DFFRX1 \i_MIPS/Register/register_reg[25][4]  ( .D(\i_MIPS/Register/n312 ), 
        .CK(clk), .RN(n6292), .Q(\i_MIPS/Register/register[25][4] ), .QN(n762)
         );
  DFFRX1 \i_MIPS/Register/register_reg[25][5]  ( .D(\i_MIPS/Register/n313 ), 
        .CK(clk), .RN(n6292), .Q(\i_MIPS/Register/register[25][5] ), .QN(n378)
         );
  DFFRX1 \i_MIPS/Register/register_reg[25][6]  ( .D(\i_MIPS/Register/n314 ), 
        .CK(clk), .RN(n6292), .Q(\i_MIPS/Register/register[25][6] ), .QN(n751)
         );
  DFFRX1 \i_MIPS/Register/register_reg[25][7]  ( .D(\i_MIPS/Register/n315 ), 
        .CK(clk), .RN(n6292), .Q(\i_MIPS/Register/register[25][7] ), .QN(n749)
         );
  DFFRX1 \i_MIPS/Register/register_reg[25][8]  ( .D(\i_MIPS/Register/n316 ), 
        .CK(clk), .RN(n6292), .Q(\i_MIPS/Register/register[25][8] ), .QN(n754)
         );
  DFFRX1 \i_MIPS/Register/register_reg[25][9]  ( .D(\i_MIPS/Register/n317 ), 
        .CK(clk), .RN(n6292), .Q(\i_MIPS/Register/register[25][9] ), .QN(n742)
         );
  DFFRX1 \i_MIPS/Register/register_reg[25][10]  ( .D(\i_MIPS/Register/n318 ), 
        .CK(clk), .RN(n6292), .Q(\i_MIPS/Register/register[25][10] ), .QN(n841) );
  DFFRX1 \i_MIPS/Register/register_reg[25][11]  ( .D(\i_MIPS/Register/n319 ), 
        .CK(clk), .RN(n6292), .Q(\i_MIPS/Register/register[25][11] ), .QN(n427) );
  DFFRX1 \i_MIPS/Register/register_reg[25][12]  ( .D(\i_MIPS/Register/n320 ), 
        .CK(clk), .RN(n6291), .Q(\i_MIPS/Register/register[25][12] ), .QN(n752) );
  DFFRX1 \i_MIPS/Register/register_reg[25][13]  ( .D(\i_MIPS/Register/n321 ), 
        .CK(clk), .RN(n6291), .Q(\i_MIPS/Register/register[25][13] ), .QN(n553) );
  DFFRX1 \i_MIPS/Register/register_reg[25][15]  ( .D(\i_MIPS/Register/n323 ), 
        .CK(clk), .RN(n6291), .Q(\i_MIPS/Register/register[25][15] ), .QN(n185) );
  DFFRX1 \i_MIPS/Register/register_reg[25][16]  ( .D(\i_MIPS/Register/n324 ), 
        .CK(clk), .RN(n6291), .Q(\i_MIPS/Register/register[25][16] ), .QN(n422) );
  DFFRX1 \i_MIPS/Register/register_reg[25][17]  ( .D(\i_MIPS/Register/n325 ), 
        .CK(clk), .RN(n6291), .Q(\i_MIPS/Register/register[25][17] ), .QN(n760) );
  DFFRX1 \i_MIPS/Register/register_reg[25][18]  ( .D(\i_MIPS/Register/n326 ), 
        .CK(clk), .RN(n6291), .Q(\i_MIPS/Register/register[25][18] ), .QN(n726) );
  DFFRX1 \i_MIPS/Register/register_reg[25][19]  ( .D(\i_MIPS/Register/n327 ), 
        .CK(clk), .RN(n6291), .Q(\i_MIPS/Register/register[25][19] ), .QN(n840) );
  DFFRX1 \i_MIPS/Register/register_reg[25][20]  ( .D(\i_MIPS/Register/n328 ), 
        .CK(clk), .RN(n6291), .Q(\i_MIPS/Register/register[25][20] ), .QN(n425) );
  DFFRX1 \i_MIPS/Register/register_reg[25][21]  ( .D(\i_MIPS/Register/n329 ), 
        .CK(clk), .RN(n6291), .Q(\i_MIPS/Register/register[25][21] ), .QN(n729) );
  DFFRX1 \i_MIPS/Register/register_reg[25][23]  ( .D(\i_MIPS/Register/n331 ), 
        .CK(clk), .RN(n6291), .Q(\i_MIPS/Register/register[25][23] ), .QN(n209) );
  DFFRX1 \i_MIPS/Register/register_reg[25][24]  ( .D(\i_MIPS/Register/n332 ), 
        .CK(clk), .RN(n6290), .Q(\i_MIPS/Register/register[25][24] ), .QN(n213) );
  DFFRX1 \i_MIPS/Register/register_reg[25][25]  ( .D(\i_MIPS/Register/n333 ), 
        .CK(clk), .RN(n6290), .Q(\i_MIPS/Register/register[25][25] ), .QN(n217) );
  DFFRX1 \i_MIPS/Register/register_reg[25][26]  ( .D(\i_MIPS/Register/n334 ), 
        .CK(clk), .RN(n6290), .Q(\i_MIPS/Register/register[25][26] ), .QN(n725) );
  DFFRX1 \i_MIPS/Register/register_reg[25][27]  ( .D(\i_MIPS/Register/n335 ), 
        .CK(clk), .RN(n6290), .Q(\i_MIPS/Register/register[25][27] ), .QN(n748) );
  DFFRX1 \i_MIPS/Register/register_reg[25][28]  ( .D(\i_MIPS/Register/n336 ), 
        .CK(clk), .RN(n6290), .Q(\i_MIPS/Register/register[25][28] ), .QN(n746) );
  DFFRX1 \i_MIPS/Register/register_reg[25][29]  ( .D(\i_MIPS/Register/n337 ), 
        .CK(clk), .RN(n6290), .Q(\i_MIPS/Register/register[25][29] ), .QN(n211) );
  DFFRX1 \i_MIPS/Register/register_reg[24][0]  ( .D(\i_MIPS/Register/n340 ), 
        .CK(clk), .RN(n6290), .Q(\i_MIPS/Register/register[24][0] ), .QN(n838)
         );
  DFFRX1 \i_MIPS/Register/register_reg[24][1]  ( .D(\i_MIPS/Register/n341 ), 
        .CK(clk), .RN(n6290), .Q(\i_MIPS/Register/register[24][1] ), .QN(n204)
         );
  DFFRX1 \i_MIPS/Register/register_reg[24][2]  ( .D(\i_MIPS/Register/n342 ), 
        .CK(clk), .RN(n6290), .Q(\i_MIPS/Register/register[24][2] ), .QN(n191)
         );
  DFFRX1 \i_MIPS/Register/register_reg[24][3]  ( .D(\i_MIPS/Register/n343 ), 
        .CK(clk), .RN(n6290), .Q(\i_MIPS/Register/register[24][3] ), .QN(n194)
         );
  DFFRX1 \i_MIPS/Register/register_reg[24][4]  ( .D(\i_MIPS/Register/n344 ), 
        .CK(clk), .RN(n6289), .Q(\i_MIPS/Register/register[24][4] ), .QN(n195)
         );
  DFFRX1 \i_MIPS/Register/register_reg[24][5]  ( .D(\i_MIPS/Register/n345 ), 
        .CK(clk), .RN(n6289), .Q(\i_MIPS/Register/register[24][5] ), .QN(n196)
         );
  DFFRX1 \i_MIPS/Register/register_reg[24][6]  ( .D(\i_MIPS/Register/n346 ), 
        .CK(clk), .RN(n6289), .Q(\i_MIPS/Register/register[24][6] ), .QN(n766)
         );
  DFFRX1 \i_MIPS/Register/register_reg[24][7]  ( .D(\i_MIPS/Register/n347 ), 
        .CK(clk), .RN(n6289), .Q(\i_MIPS/Register/register[24][7] ), .QN(n765)
         );
  DFFRX1 \i_MIPS/Register/register_reg[24][8]  ( .D(\i_MIPS/Register/n348 ), 
        .CK(clk), .RN(n6289), .Q(\i_MIPS/Register/register[24][8] ), .QN(n736)
         );
  DFFRX1 \i_MIPS/Register/register_reg[24][9]  ( .D(\i_MIPS/Register/n349 ), 
        .CK(clk), .RN(n6289), .Q(\i_MIPS/Register/register[24][9] ), .QN(n770)
         );
  DFFRX1 \i_MIPS/Register/register_reg[24][10]  ( .D(\i_MIPS/Register/n350 ), 
        .CK(clk), .RN(n6289), .Q(\i_MIPS/Register/register[24][10] ), .QN(n724) );
  DFFRX1 \i_MIPS/Register/register_reg[24][11]  ( .D(\i_MIPS/Register/n351 ), 
        .CK(clk), .RN(n6289), .Q(\i_MIPS/Register/register[24][11] ), .QN(n768) );
  DFFRX1 \i_MIPS/Register/register_reg[24][12]  ( .D(\i_MIPS/Register/n352 ), 
        .CK(clk), .RN(n6289), .Q(\i_MIPS/Register/register[24][12] ), .QN(n738) );
  DFFRX1 \i_MIPS/Register/register_reg[24][13]  ( .D(\i_MIPS/Register/n353 ), 
        .CK(clk), .RN(n6289), .Q(\i_MIPS/Register/register[24][13] ), .QN(n756) );
  DFFRX1 \i_MIPS/Register/register_reg[24][16]  ( .D(\i_MIPS/Register/n356 ), 
        .CK(clk), .RN(n6288), .Q(\i_MIPS/Register/register[24][16] ), .QN(n728) );
  DFFRX1 \i_MIPS/Register/register_reg[24][17]  ( .D(\i_MIPS/Register/n357 ), 
        .CK(clk), .RN(n6288), .Q(\i_MIPS/Register/register[24][17] ), .QN(n212) );
  DFFRX1 \i_MIPS/Register/register_reg[24][18]  ( .D(\i_MIPS/Register/n358 ), 
        .CK(clk), .RN(n6288), .Q(\i_MIPS/Register/register[24][18] ), .QN(n767) );
  DFFRX1 \i_MIPS/Register/register_reg[24][19]  ( .D(\i_MIPS/Register/n359 ), 
        .CK(clk), .RN(n6288), .Q(\i_MIPS/Register/register[24][19] ), .QN(n834) );
  DFFRX1 \i_MIPS/Register/register_reg[24][20]  ( .D(\i_MIPS/Register/n360 ), 
        .CK(clk), .RN(n6288), .Q(\i_MIPS/Register/register[24][20] ), .QN(n551) );
  DFFRX1 \i_MIPS/Register/register_reg[24][21]  ( .D(\i_MIPS/Register/n361 ), 
        .CK(clk), .RN(n6288), .Q(\i_MIPS/Register/register[24][21] ), .QN(n556) );
  DFFRX1 \i_MIPS/Register/register_reg[24][23]  ( .D(\i_MIPS/Register/n363 ), 
        .CK(clk), .RN(n6288), .Q(\i_MIPS/Register/register[24][23] ), .QN(n207) );
  DFFRX1 \i_MIPS/Register/register_reg[24][26]  ( .D(\i_MIPS/Register/n366 ), 
        .CK(clk), .RN(n6288), .Q(\i_MIPS/Register/register[24][26] ), .QN(n759) );
  DFFRX1 \i_MIPS/Register/register_reg[24][27]  ( .D(\i_MIPS/Register/n367 ), 
        .CK(clk), .RN(n6288), .Q(\i_MIPS/Register/register[24][27] ), .QN(n741) );
  DFFRX1 \i_MIPS/Register/register_reg[24][28]  ( .D(\i_MIPS/Register/n368 ), 
        .CK(clk), .RN(n6287), .Q(\i_MIPS/Register/register[24][28] ), .QN(n758) );
  DFFRX1 \i_MIPS/Register/register_reg[24][29]  ( .D(\i_MIPS/Register/n369 ), 
        .CK(clk), .RN(n6287), .Q(\i_MIPS/Register/register[24][29] ), .QN(n189) );
  DFFRX1 \i_MIPS/Register/register_reg[15][0]  ( .D(\i_MIPS/Register/n628 ), 
        .CK(clk), .RN(n6266), .Q(\i_MIPS/Register/register[15][0] ), .QN(n789)
         );
  DFFRX1 \i_MIPS/Register/register_reg[15][1]  ( .D(\i_MIPS/Register/n629 ), 
        .CK(clk), .RN(n6266), .Q(\i_MIPS/Register/register[15][1] ), .QN(n777)
         );
  DFFRX1 \i_MIPS/Register/register_reg[15][2]  ( .D(\i_MIPS/Register/n630 ), 
        .CK(clk), .RN(n6266), .Q(\i_MIPS/Register/register[15][2] ), .QN(n817)
         );
  DFFRX1 \i_MIPS/Register/register_reg[15][3]  ( .D(\i_MIPS/Register/n631 ), 
        .CK(clk), .RN(n6266), .Q(\i_MIPS/Register/register[15][3] ), .QN(n793)
         );
  DFFRX1 \i_MIPS/Register/register_reg[15][4]  ( .D(\i_MIPS/Register/n632 ), 
        .CK(clk), .RN(n6265), .Q(\i_MIPS/Register/register[15][4] ), .QN(n876)
         );
  DFFRX1 \i_MIPS/Register/register_reg[15][5]  ( .D(\i_MIPS/Register/n633 ), 
        .CK(clk), .RN(n6265), .Q(\i_MIPS/Register/register[15][5] ), .QN(n786)
         );
  DFFRX1 \i_MIPS/Register/register_reg[15][6]  ( .D(\i_MIPS/Register/n634 ), 
        .CK(clk), .RN(n6265), .Q(\i_MIPS/Register/register[15][6] ), .QN(n806)
         );
  DFFRX1 \i_MIPS/Register/register_reg[15][7]  ( .D(\i_MIPS/Register/n635 ), 
        .CK(clk), .RN(n6265), .Q(\i_MIPS/Register/register[15][7] ), .QN(n390)
         );
  DFFRX1 \i_MIPS/Register/register_reg[15][8]  ( .D(\i_MIPS/Register/n636 ), 
        .CK(clk), .RN(n6265), .Q(\i_MIPS/Register/register[15][8] ), .QN(n203)
         );
  DFFRX1 \i_MIPS/Register/register_reg[15][9]  ( .D(\i_MIPS/Register/n637 ), 
        .CK(clk), .RN(n6265), .Q(\i_MIPS/Register/register[15][9] ), .QN(n180)
         );
  DFFRX1 \i_MIPS/Register/register_reg[15][10]  ( .D(\i_MIPS/Register/n638 ), 
        .CK(clk), .RN(n6265), .Q(\i_MIPS/Register/register[15][10] ), .QN(n381) );
  DFFRX1 \i_MIPS/Register/register_reg[15][11]  ( .D(\i_MIPS/Register/n639 ), 
        .CK(clk), .RN(n6265), .Q(\i_MIPS/Register/register[15][11] ), .QN(n798) );
  DFFRX1 \i_MIPS/Register/register_reg[15][12]  ( .D(\i_MIPS/Register/n640 ), 
        .CK(clk), .RN(n6265), .Q(\i_MIPS/Register/register[15][12] ), .QN(n201) );
  DFFRX1 \i_MIPS/Register/register_reg[15][13]  ( .D(\i_MIPS/Register/n641 ), 
        .CK(clk), .RN(n6265), .Q(\i_MIPS/Register/register[15][13] ), .QN(n181) );
  DFFRX1 \i_MIPS/Register/register_reg[15][15]  ( .D(\i_MIPS/Register/n643 ), 
        .CK(clk), .RN(n6265), .Q(\i_MIPS/Register/register[15][15] ), .QN(n890) );
  DFFRX1 \i_MIPS/Register/register_reg[15][16]  ( .D(\i_MIPS/Register/n644 ), 
        .CK(clk), .RN(n6264), .Q(\i_MIPS/Register/register[15][16] ), .QN(n800) );
  DFFRX1 \i_MIPS/Register/register_reg[15][17]  ( .D(\i_MIPS/Register/n645 ), 
        .CK(clk), .RN(n6264), .Q(\i_MIPS/Register/register[15][17] ), .QN(n856) );
  DFFRX1 \i_MIPS/Register/register_reg[15][18]  ( .D(\i_MIPS/Register/n646 ), 
        .CK(clk), .RN(n6264), .Q(\i_MIPS/Register/register[15][18] ), .QN(n784) );
  DFFRX1 \i_MIPS/Register/register_reg[15][19]  ( .D(\i_MIPS/Register/n647 ), 
        .CK(clk), .RN(n6264), .Q(\i_MIPS/Register/register[15][19] ), .QN(n202) );
  DFFRX1 \i_MIPS/Register/register_reg[15][20]  ( .D(\i_MIPS/Register/n648 ), 
        .CK(clk), .RN(n6264), .Q(\i_MIPS/Register/register[15][20] ), .QN(n864) );
  DFFRX1 \i_MIPS/Register/register_reg[15][21]  ( .D(\i_MIPS/Register/n649 ), 
        .CK(clk), .RN(n6264), .Q(\i_MIPS/Register/register[15][21] ), .QN(n866) );
  DFFRX1 \i_MIPS/Register/register_reg[15][23]  ( .D(\i_MIPS/Register/n651 ), 
        .CK(clk), .RN(n6264), .Q(\i_MIPS/Register/register[15][23] ), .QN(n813) );
  DFFRX1 \i_MIPS/Register/register_reg[15][24]  ( .D(\i_MIPS/Register/n652 ), 
        .CK(clk), .RN(n6264), .Q(\i_MIPS/Register/register[15][24] ), .QN(n391) );
  DFFRX1 \i_MIPS/Register/register_reg[15][25]  ( .D(\i_MIPS/Register/n653 ), 
        .CK(clk), .RN(n6264), .Q(\i_MIPS/Register/register[15][25] ), .QN(n909) );
  DFFRX1 \i_MIPS/Register/register_reg[15][26]  ( .D(\i_MIPS/Register/n654 ), 
        .CK(clk), .RN(n6264), .Q(\i_MIPS/Register/register[15][26] ), .QN(n871) );
  DFFRX1 \i_MIPS/Register/register_reg[15][27]  ( .D(\i_MIPS/Register/n655 ), 
        .CK(clk), .RN(n6264), .Q(\i_MIPS/Register/register[15][27] ), .QN(n824) );
  DFFRX1 \i_MIPS/Register/register_reg[15][28]  ( .D(\i_MIPS/Register/n656 ), 
        .CK(clk), .RN(n6263), .Q(\i_MIPS/Register/register[15][28] ), .QN(n386) );
  DFFRX1 \i_MIPS/Register/register_reg[15][29]  ( .D(\i_MIPS/Register/n657 ), 
        .CK(clk), .RN(n6263), .Q(\i_MIPS/Register/register[15][29] ), .QN(n388) );
  DFFRX1 \i_MIPS/Register/register_reg[13][0]  ( .D(\i_MIPS/Register/n692 ), 
        .CK(clk), .RN(n6260), .Q(\i_MIPS/Register/register[13][0] ), .QN(n274)
         );
  DFFRX1 \i_MIPS/Register/register_reg[13][1]  ( .D(\i_MIPS/Register/n693 ), 
        .CK(clk), .RN(n6260), .Q(\i_MIPS/Register/register[13][1] ), .QN(n779)
         );
  DFFRX1 \i_MIPS/Register/register_reg[13][2]  ( .D(\i_MIPS/Register/n694 ), 
        .CK(clk), .RN(n6260), .Q(\i_MIPS/Register/register[13][2] ), .QN(n819)
         );
  DFFRX1 \i_MIPS/Register/register_reg[13][3]  ( .D(\i_MIPS/Register/n695 ), 
        .CK(clk), .RN(n6260), .Q(\i_MIPS/Register/register[13][3] ), .QN(n795)
         );
  DFFRX1 \i_MIPS/Register/register_reg[13][4]  ( .D(\i_MIPS/Register/n696 ), 
        .CK(clk), .RN(n6260), .Q(\i_MIPS/Register/register[13][4] ), .QN(n878)
         );
  DFFRX1 \i_MIPS/Register/register_reg[13][5]  ( .D(\i_MIPS/Register/n697 ), 
        .CK(clk), .RN(n6260), .Q(\i_MIPS/Register/register[13][5] ), .QN(n788)
         );
  DFFRX1 \i_MIPS/Register/register_reg[13][6]  ( .D(\i_MIPS/Register/n698 ), 
        .CK(clk), .RN(n6260), .Q(\i_MIPS/Register/register[13][6] ), .QN(n808)
         );
  DFFRX1 \i_MIPS/Register/register_reg[13][7]  ( .D(\i_MIPS/Register/n699 ), 
        .CK(clk), .RN(n6260), .Q(\i_MIPS/Register/register[13][7] ), .QN(n882)
         );
  DFFRX1 \i_MIPS/Register/register_reg[13][8]  ( .D(\i_MIPS/Register/n700 ), 
        .CK(clk), .RN(n6260), .Q(\i_MIPS/Register/register[13][8] ), .QN(n868)
         );
  DFFRX1 \i_MIPS/Register/register_reg[13][9]  ( .D(\i_MIPS/Register/n701 ), 
        .CK(clk), .RN(n6260), .Q(\i_MIPS/Register/register[13][9] ), .QN(n385)
         );
  DFFRX1 \i_MIPS/Register/register_reg[13][10]  ( .D(\i_MIPS/Register/n702 ), 
        .CK(clk), .RN(n6260), .Q(\i_MIPS/Register/register[13][10] ), .QN(n383) );
  DFFRX1 \i_MIPS/Register/register_reg[13][11]  ( .D(\i_MIPS/Register/n703 ), 
        .CK(clk), .RN(n6260), .Q(\i_MIPS/Register/register[13][11] ), .QN(n276) );
  DFFRX1 \i_MIPS/Register/register_reg[13][12]  ( .D(\i_MIPS/Register/n704 ), 
        .CK(clk), .RN(n6259), .Q(\i_MIPS/Register/register[13][12] ), .QN(n861) );
  DFFRX1 \i_MIPS/Register/register_reg[13][13]  ( .D(\i_MIPS/Register/n705 ), 
        .CK(clk), .RN(n6259), .Q(\i_MIPS/Register/register[13][13] ), .QN(n805) );
  DFFRX1 \i_MIPS/Register/register_reg[13][15]  ( .D(\i_MIPS/Register/n707 ), 
        .CK(clk), .RN(n6259), .Q(\i_MIPS/Register/register[13][15] ), .QN(n892) );
  DFFRX1 \i_MIPS/Register/register_reg[13][16]  ( .D(\i_MIPS/Register/n708 ), 
        .CK(clk), .RN(n6259), .Q(\i_MIPS/Register/register[13][16] ), .QN(n277) );
  DFFRX1 \i_MIPS/Register/register_reg[13][17]  ( .D(\i_MIPS/Register/n709 ), 
        .CK(clk), .RN(n6259), .Q(\i_MIPS/Register/register[13][17] ), .QN(n858) );
  DFFRX1 \i_MIPS/Register/register_reg[13][18]  ( .D(\i_MIPS/Register/n710 ), 
        .CK(clk), .RN(n6259), .Q(\i_MIPS/Register/register[13][18] ), .QN(n273) );
  DFFRX1 \i_MIPS/Register/register_reg[13][19]  ( .D(\i_MIPS/Register/n711 ), 
        .CK(clk), .RN(n6259), .Q(\i_MIPS/Register/register[13][19] ), .QN(n554) );
  DFFRX1 \i_MIPS/Register/register_reg[13][20]  ( .D(\i_MIPS/Register/n712 ), 
        .CK(clk), .RN(n6259), .Q(\i_MIPS/Register/register[13][20] ), .QN(n296) );
  DFFRX1 \i_MIPS/Register/register_reg[13][21]  ( .D(\i_MIPS/Register/n713 ), 
        .CK(clk), .RN(n6259), .Q(\i_MIPS/Register/register[13][21] ), .QN(n298) );
  DFFRX1 \i_MIPS/Register/register_reg[13][23]  ( .D(\i_MIPS/Register/n715 ), 
        .CK(clk), .RN(n6259), .Q(\i_MIPS/Register/register[13][23] ), .QN(n815) );
  DFFRX1 \i_MIPS/Register/register_reg[13][24]  ( .D(\i_MIPS/Register/n716 ), 
        .CK(clk), .RN(n6258), .Q(\i_MIPS/Register/register[13][24] ), .QN(n908) );
  DFFRX1 \i_MIPS/Register/register_reg[13][25]  ( .D(\i_MIPS/Register/n717 ), 
        .CK(clk), .RN(n6258), .Q(\i_MIPS/Register/register[13][25] ), .QN(n911) );
  DFFRX1 \i_MIPS/Register/register_reg[13][26]  ( .D(\i_MIPS/Register/n718 ), 
        .CK(clk), .RN(n6258), .Q(\i_MIPS/Register/register[13][26] ), .QN(n873) );
  DFFRX1 \i_MIPS/Register/register_reg[13][27]  ( .D(\i_MIPS/Register/n719 ), 
        .CK(clk), .RN(n6258), .Q(\i_MIPS/Register/register[13][27] ), .QN(n826) );
  DFFRX1 \i_MIPS/Register/register_reg[13][28]  ( .D(\i_MIPS/Register/n720 ), 
        .CK(clk), .RN(n6258), .Q(\i_MIPS/Register/register[13][28] ), .QN(n886) );
  DFFRX1 \i_MIPS/Register/register_reg[13][29]  ( .D(\i_MIPS/Register/n721 ), 
        .CK(clk), .RN(n6258), .Q(\i_MIPS/Register/register[13][29] ), .QN(n821) );
  DFFRX1 \i_MIPS/Register/register_reg[12][0]  ( .D(\i_MIPS/Register/n724 ), 
        .CK(clk), .RN(n6258), .Q(\i_MIPS/Register/register[12][0] ), .QN(n846)
         );
  DFFRX1 \i_MIPS/Register/register_reg[12][1]  ( .D(\i_MIPS/Register/n725 ), 
        .CK(clk), .RN(n6258), .Q(\i_MIPS/Register/register[12][1] ), .QN(n289)
         );
  DFFRX1 \i_MIPS/Register/register_reg[12][3]  ( .D(\i_MIPS/Register/n727 ), 
        .CK(clk), .RN(n6258), .Q(\i_MIPS/Register/register[12][3] ), .QN(n267)
         );
  DFFRX1 \i_MIPS/Register/register_reg[12][4]  ( .D(\i_MIPS/Register/n728 ), 
        .CK(clk), .RN(n6257), .Q(\i_MIPS/Register/register[12][4] ), .QN(n288)
         );
  DFFRX1 \i_MIPS/Register/register_reg[12][5]  ( .D(\i_MIPS/Register/n729 ), 
        .CK(clk), .RN(n6257), .Q(\i_MIPS/Register/register[12][5] ), .QN(n265)
         );
  DFFRX1 \i_MIPS/Register/register_reg[12][6]  ( .D(\i_MIPS/Register/n730 ), 
        .CK(clk), .RN(n6257), .Q(\i_MIPS/Register/register[12][6] ), .QN(n849)
         );
  DFFRX1 \i_MIPS/Register/register_reg[12][7]  ( .D(\i_MIPS/Register/n731 ), 
        .CK(clk), .RN(n6257), .Q(\i_MIPS/Register/register[12][7] ), .QN(n901)
         );
  DFFRX1 \i_MIPS/Register/register_reg[12][8]  ( .D(\i_MIPS/Register/n732 ), 
        .CK(clk), .RN(n6257), .Q(\i_MIPS/Register/register[12][8] ), .QN(n848)
         );
  DFFRX1 \i_MIPS/Register/register_reg[12][9]  ( .D(\i_MIPS/Register/n733 ), 
        .CK(clk), .RN(n6257), .Q(\i_MIPS/Register/register[12][9] ), .QN(n561)
         );
  DFFRX1 \i_MIPS/Register/register_reg[12][10]  ( .D(\i_MIPS/Register/n734 ), 
        .CK(clk), .RN(n6257), .Q(\i_MIPS/Register/register[12][10] ), .QN(n722) );
  DFFRX1 \i_MIPS/Register/register_reg[12][11]  ( .D(\i_MIPS/Register/n735 ), 
        .CK(clk), .RN(n6257), .Q(\i_MIPS/Register/register[12][11] ), .QN(n843) );
  DFFRX1 \i_MIPS/Register/register_reg[12][12]  ( .D(\i_MIPS/Register/n736 ), 
        .CK(clk), .RN(n6257), .Q(\i_MIPS/Register/register[12][12] ), .QN(n847) );
  DFFRX1 \i_MIPS/Register/register_reg[12][13]  ( .D(\i_MIPS/Register/n737 ), 
        .CK(clk), .RN(n6257), .Q(\i_MIPS/Register/register[12][13] ), .QN(n851) );
  DFFRX1 \i_MIPS/Register/register_reg[12][16]  ( .D(\i_MIPS/Register/n740 ), 
        .CK(clk), .RN(n6256), .Q(\i_MIPS/Register/register[12][16] ), .QN(n845) );
  DFFRX1 \i_MIPS/Register/register_reg[12][17]  ( .D(\i_MIPS/Register/n741 ), 
        .CK(clk), .RN(n6256), .Q(\i_MIPS/Register/register[12][17] ), .QN(n264) );
  DFFRX1 \i_MIPS/Register/register_reg[12][18]  ( .D(\i_MIPS/Register/n742 ), 
        .CK(clk), .RN(n6256), .Q(\i_MIPS/Register/register[12][18] ), .QN(n416) );
  DFFRX1 \i_MIPS/Register/register_reg[12][19]  ( .D(\i_MIPS/Register/n743 ), 
        .CK(clk), .RN(n6256), .Q(\i_MIPS/Register/register[12][19] ), .QN(n844) );
  DFFRX1 \i_MIPS/Register/register_reg[12][20]  ( .D(\i_MIPS/Register/n744 ), 
        .CK(clk), .RN(n6256), .Q(\i_MIPS/Register/register[12][20] ), .QN(n418) );
  DFFRX1 \i_MIPS/Register/register_reg[12][21]  ( .D(\i_MIPS/Register/n745 ), 
        .CK(clk), .RN(n6256), .Q(\i_MIPS/Register/register[12][21] ), .QN(n417) );
  DFFRX1 \i_MIPS/Register/register_reg[12][23]  ( .D(\i_MIPS/Register/n747 ), 
        .CK(clk), .RN(n6256), .Q(\i_MIPS/Register/register[12][23] ), .QN(n290) );
  DFFRX1 \i_MIPS/Register/register_reg[12][26]  ( .D(\i_MIPS/Register/n750 ), 
        .CK(clk), .RN(n6256), .Q(\i_MIPS/Register/register[12][26] ), .QN(n850) );
  DFFRX1 \i_MIPS/Register/register_reg[12][27]  ( .D(\i_MIPS/Register/n751 ), 
        .CK(clk), .RN(n6256), .Q(\i_MIPS/Register/register[12][27] ), .QN(n852) );
  DFFRX1 \i_MIPS/Register/register_reg[11][0]  ( .D(\i_MIPS/Register/n756 ), 
        .CK(clk), .RN(n6255), .Q(\i_MIPS/Register/register[11][0] ), .QN(n790)
         );
  DFFRX1 \i_MIPS/Register/register_reg[11][1]  ( .D(\i_MIPS/Register/n757 ), 
        .CK(clk), .RN(n6255), .Q(\i_MIPS/Register/register[11][1] ), .QN(n778)
         );
  DFFRX1 \i_MIPS/Register/register_reg[11][2]  ( .D(\i_MIPS/Register/n758 ), 
        .CK(clk), .RN(n6255), .Q(\i_MIPS/Register/register[11][2] ), .QN(n818)
         );
  DFFRX1 \i_MIPS/Register/register_reg[11][3]  ( .D(\i_MIPS/Register/n759 ), 
        .CK(clk), .RN(n6255), .Q(\i_MIPS/Register/register[11][3] ), .QN(n794)
         );
  DFFRX1 \i_MIPS/Register/register_reg[11][4]  ( .D(\i_MIPS/Register/n760 ), 
        .CK(clk), .RN(n6255), .Q(\i_MIPS/Register/register[11][4] ), .QN(n877)
         );
  DFFRX1 \i_MIPS/Register/register_reg[11][5]  ( .D(\i_MIPS/Register/n761 ), 
        .CK(clk), .RN(n6255), .Q(\i_MIPS/Register/register[11][5] ), .QN(n787)
         );
  DFFRX1 \i_MIPS/Register/register_reg[11][6]  ( .D(\i_MIPS/Register/n762 ), 
        .CK(clk), .RN(n6255), .Q(\i_MIPS/Register/register[11][6] ), .QN(n807)
         );
  DFFRX1 \i_MIPS/Register/register_reg[11][7]  ( .D(\i_MIPS/Register/n763 ), 
        .CK(clk), .RN(n6255), .Q(\i_MIPS/Register/register[11][7] ), .QN(n881)
         );
  DFFRX1 \i_MIPS/Register/register_reg[11][8]  ( .D(\i_MIPS/Register/n764 ), 
        .CK(clk), .RN(n6254), .Q(\i_MIPS/Register/register[11][8] ), .QN(n280)
         );
  DFFRX1 \i_MIPS/Register/register_reg[11][9]  ( .D(\i_MIPS/Register/n765 ), 
        .CK(clk), .RN(n6254), .Q(\i_MIPS/Register/register[11][9] ), .QN(n250)
         );
  DFFRX1 \i_MIPS/Register/register_reg[11][10]  ( .D(\i_MIPS/Register/n766 ), 
        .CK(clk), .RN(n6254), .Q(\i_MIPS/Register/register[11][10] ), .QN(n382) );
  DFFRX1 \i_MIPS/Register/register_reg[11][11]  ( .D(\i_MIPS/Register/n767 ), 
        .CK(clk), .RN(n6254), .Q(\i_MIPS/Register/register[11][11] ), .QN(n799) );
  DFFRX1 \i_MIPS/Register/register_reg[11][12]  ( .D(\i_MIPS/Register/n768 ), 
        .CK(clk), .RN(n6254), .Q(\i_MIPS/Register/register[11][12] ), .QN(n271) );
  DFFRX1 \i_MIPS/Register/register_reg[11][13]  ( .D(\i_MIPS/Register/n769 ), 
        .CK(clk), .RN(n6254), .Q(\i_MIPS/Register/register[11][13] ), .QN(n282) );
  DFFRX1 \i_MIPS/Register/register_reg[11][15]  ( .D(\i_MIPS/Register/n771 ), 
        .CK(clk), .RN(n6254), .Q(\i_MIPS/Register/register[11][15] ), .QN(n891) );
  DFFRX1 \i_MIPS/Register/register_reg[11][16]  ( .D(\i_MIPS/Register/n772 ), 
        .CK(clk), .RN(n6254), .Q(\i_MIPS/Register/register[11][16] ), .QN(n801) );
  DFFRX1 \i_MIPS/Register/register_reg[11][17]  ( .D(\i_MIPS/Register/n773 ), 
        .CK(clk), .RN(n6254), .Q(\i_MIPS/Register/register[11][17] ), .QN(n857) );
  DFFRX1 \i_MIPS/Register/register_reg[11][18]  ( .D(\i_MIPS/Register/n774 ), 
        .CK(clk), .RN(n6254), .Q(\i_MIPS/Register/register[11][18] ), .QN(n785) );
  DFFRX1 \i_MIPS/Register/register_reg[11][19]  ( .D(\i_MIPS/Register/n775 ), 
        .CK(clk), .RN(n6254), .Q(\i_MIPS/Register/register[11][19] ), .QN(n260) );
  DFFRX1 \i_MIPS/Register/register_reg[11][20]  ( .D(\i_MIPS/Register/n776 ), 
        .CK(clk), .RN(n6253), .Q(\i_MIPS/Register/register[11][20] ), .QN(n865) );
  DFFRX1 \i_MIPS/Register/register_reg[11][21]  ( .D(\i_MIPS/Register/n777 ), 
        .CK(clk), .RN(n6253), .Q(\i_MIPS/Register/register[11][21] ), .QN(n803) );
  DFFRX1 \i_MIPS/Register/register_reg[11][23]  ( .D(\i_MIPS/Register/n779 ), 
        .CK(clk), .RN(n6253), .Q(\i_MIPS/Register/register[11][23] ), .QN(n814) );
  DFFRX1 \i_MIPS/Register/register_reg[11][24]  ( .D(\i_MIPS/Register/n780 ), 
        .CK(clk), .RN(n6253), .Q(\i_MIPS/Register/register[11][24] ), .QN(n907) );
  DFFRX1 \i_MIPS/Register/register_reg[11][25]  ( .D(\i_MIPS/Register/n781 ), 
        .CK(clk), .RN(n6253), .Q(\i_MIPS/Register/register[11][25] ), .QN(n910) );
  DFFRX1 \i_MIPS/Register/register_reg[11][26]  ( .D(\i_MIPS/Register/n782 ), 
        .CK(clk), .RN(n6253), .Q(\i_MIPS/Register/register[11][26] ), .QN(n872) );
  DFFRX1 \i_MIPS/Register/register_reg[11][27]  ( .D(\i_MIPS/Register/n783 ), 
        .CK(clk), .RN(n6253), .Q(\i_MIPS/Register/register[11][27] ), .QN(n825) );
  DFFRX1 \i_MIPS/Register/register_reg[11][28]  ( .D(\i_MIPS/Register/n784 ), 
        .CK(clk), .RN(n6253), .Q(\i_MIPS/Register/register[11][28] ), .QN(n810) );
  DFFRX1 \i_MIPS/Register/register_reg[11][29]  ( .D(\i_MIPS/Register/n785 ), 
        .CK(clk), .RN(n6253), .Q(\i_MIPS/Register/register[11][29] ), .QN(n389) );
  DFFRX1 \i_MIPS/Register/register_reg[9][0]  ( .D(\i_MIPS/Register/n820 ), 
        .CK(clk), .RN(n6250), .Q(\i_MIPS/Register/register[9][0] ), .QN(n421)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][1]  ( .D(\i_MIPS/Register/n821 ), 
        .CK(clk), .RN(n6250), .Q(\i_MIPS/Register/register[9][1] ), .QN(n837)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][2]  ( .D(\i_MIPS/Register/n822 ), 
        .CK(clk), .RN(n6250), .Q(\i_MIPS/Register/register[9][2] ), .QN(n199)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][3]  ( .D(\i_MIPS/Register/n823 ), 
        .CK(clk), .RN(n6250), .Q(\i_MIPS/Register/register[9][3] ), .QN(n735)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][4]  ( .D(\i_MIPS/Register/n824 ), 
        .CK(clk), .RN(n6249), .Q(\i_MIPS/Register/register[9][4] ), .QN(n763)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][5]  ( .D(\i_MIPS/Register/n825 ), 
        .CK(clk), .RN(n6249), .Q(\i_MIPS/Register/register[9][5] ), .QN(n743)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][6]  ( .D(\i_MIPS/Register/n826 ), 
        .CK(clk), .RN(n6249), .Q(\i_MIPS/Register/register[9][6] ), .QN(n731)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][7]  ( .D(\i_MIPS/Register/n827 ), 
        .CK(clk), .RN(n6249), .Q(\i_MIPS/Register/register[9][7] ), .QN(n750)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][8]  ( .D(\i_MIPS/Register/n828 ), 
        .CK(clk), .RN(n6249), .Q(\i_MIPS/Register/register[9][8] ), .QN(n755)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][9]  ( .D(\i_MIPS/Register/n829 ), 
        .CK(clk), .RN(n6249), .Q(\i_MIPS/Register/register[9][9] ), .QN(n377)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][10]  ( .D(\i_MIPS/Register/n830 ), 
        .CK(clk), .RN(n6249), .Q(\i_MIPS/Register/register[9][10] ), .QN(n842)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][11]  ( .D(\i_MIPS/Register/n831 ), 
        .CK(clk), .RN(n6249), .Q(\i_MIPS/Register/register[9][11] ), .QN(n772)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][12]  ( .D(\i_MIPS/Register/n832 ), 
        .CK(clk), .RN(n6249), .Q(\i_MIPS/Register/register[9][12] ), .QN(n753)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][13]  ( .D(\i_MIPS/Register/n833 ), 
        .CK(clk), .RN(n6249), .Q(\i_MIPS/Register/register[9][13] ), .QN(n744)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][15]  ( .D(\i_MIPS/Register/n835 ), 
        .CK(clk), .RN(n6249), .Q(\i_MIPS/Register/register[9][15] ), .QN(n184)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][16]  ( .D(\i_MIPS/Register/n836 ), 
        .CK(clk), .RN(n6248), .Q(\i_MIPS/Register/register[9][16] ), .QN(n423)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][17]  ( .D(\i_MIPS/Register/n837 ), 
        .CK(clk), .RN(n6248), .Q(\i_MIPS/Register/register[9][17] ), .QN(n761)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][18]  ( .D(\i_MIPS/Register/n838 ), 
        .CK(clk), .RN(n6248), .Q(\i_MIPS/Register/register[9][18] ), .QN(n773)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][19]  ( .D(\i_MIPS/Register/n839 ), 
        .CK(clk), .RN(n6248), .Q(\i_MIPS/Register/register[9][19] ), .QN(n555)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][20]  ( .D(\i_MIPS/Register/n840 ), 
        .CK(clk), .RN(n6248), .Q(\i_MIPS/Register/register[9][20] ), .QN(n426)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][21]  ( .D(\i_MIPS/Register/n841 ), 
        .CK(clk), .RN(n6248), .Q(\i_MIPS/Register/register[9][21] ), .QN(n419)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][23]  ( .D(\i_MIPS/Register/n843 ), 
        .CK(clk), .RN(n6248), .Q(\i_MIPS/Register/register[9][23] ), .QN(n210)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][24]  ( .D(\i_MIPS/Register/n844 ), 
        .CK(clk), .RN(n6248), .Q(\i_MIPS/Register/register[9][24] ), .QN(n218)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][25]  ( .D(\i_MIPS/Register/n845 ), 
        .CK(clk), .RN(n6248), .Q(\i_MIPS/Register/register[9][25] ), .QN(n216)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][26]  ( .D(\i_MIPS/Register/n846 ), 
        .CK(clk), .RN(n6248), .Q(\i_MIPS/Register/register[9][26] ), .QN(n900)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][27]  ( .D(\i_MIPS/Register/n847 ), 
        .CK(clk), .RN(n6248), .Q(\i_MIPS/Register/register[9][27] ), .QN(n730)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][28]  ( .D(\i_MIPS/Register/n848 ), 
        .CK(clk), .RN(n6247), .Q(\i_MIPS/Register/register[9][28] ), .QN(n747)
         );
  DFFRX1 \i_MIPS/Register/register_reg[9][29]  ( .D(\i_MIPS/Register/n849 ), 
        .CK(clk), .RN(n6247), .Q(\i_MIPS/Register/register[9][29] ), .QN(n198)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][0]  ( .D(\i_MIPS/Register/n852 ), 
        .CK(clk), .RN(n6247), .Q(\i_MIPS/Register/register[8][0] ), .QN(n839)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][1]  ( .D(\i_MIPS/Register/n853 ), 
        .CK(clk), .RN(n6247), .Q(\i_MIPS/Register/register[8][1] ), .QN(n206)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][2]  ( .D(\i_MIPS/Register/n854 ), 
        .CK(clk), .RN(n6247), .Q(\i_MIPS/Register/register[8][2] ), .QN(n190)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][3]  ( .D(\i_MIPS/Register/n855 ), 
        .CK(clk), .RN(n6247), .Q(\i_MIPS/Register/register[8][3] ), .QN(n193)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][4]  ( .D(\i_MIPS/Register/n856 ), 
        .CK(clk), .RN(n6247), .Q(\i_MIPS/Register/register[8][4] ), .QN(n192)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][5]  ( .D(\i_MIPS/Register/n857 ), 
        .CK(clk), .RN(n6247), .Q(\i_MIPS/Register/register[8][5] ), .QN(n188)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][6]  ( .D(\i_MIPS/Register/n858 ), 
        .CK(clk), .RN(n6247), .Q(\i_MIPS/Register/register[8][6] ), .QN(n745)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][7]  ( .D(\i_MIPS/Register/n859 ), 
        .CK(clk), .RN(n6247), .Q(\i_MIPS/Register/register[8][7] ), .QN(n764)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][8]  ( .D(\i_MIPS/Register/n860 ), 
        .CK(clk), .RN(n6246), .Q(\i_MIPS/Register/register[8][8] ), .QN(n733)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][9]  ( .D(\i_MIPS/Register/n861 ), 
        .CK(clk), .RN(n6246), .Q(\i_MIPS/Register/register[8][9] ), .QN(n720)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][10]  ( .D(\i_MIPS/Register/n862 ), 
        .CK(clk), .RN(n6246), .Q(\i_MIPS/Register/register[8][10] ), .QN(n721)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][11]  ( .D(\i_MIPS/Register/n863 ), 
        .CK(clk), .RN(n6246), .Q(\i_MIPS/Register/register[8][11] ), .QN(n769)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][12]  ( .D(\i_MIPS/Register/n864 ), 
        .CK(clk), .RN(n6246), .Q(\i_MIPS/Register/register[8][12] ), .QN(n737)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][13]  ( .D(\i_MIPS/Register/n865 ), 
        .CK(clk), .RN(n6246), .Q(\i_MIPS/Register/register[8][13] ), .QN(n739)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][16]  ( .D(\i_MIPS/Register/n868 ), 
        .CK(clk), .RN(n6246), .Q(\i_MIPS/Register/register[8][16] ), .QN(n727)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][17]  ( .D(\i_MIPS/Register/n869 ), 
        .CK(clk), .RN(n6246), .Q(\i_MIPS/Register/register[8][17] ), .QN(n197)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][18]  ( .D(\i_MIPS/Register/n870 ), 
        .CK(clk), .RN(n6246), .Q(\i_MIPS/Register/register[8][18] ), .QN(n771)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][19]  ( .D(\i_MIPS/Register/n871 ), 
        .CK(clk), .RN(n6246), .Q(\i_MIPS/Register/register[8][19] ), .QN(n835)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][20]  ( .D(\i_MIPS/Register/n872 ), 
        .CK(clk), .RN(n6245), .Q(\i_MIPS/Register/register[8][20] ), .QN(n550)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][21]  ( .D(\i_MIPS/Register/n873 ), 
        .CK(clk), .RN(n6245), .Q(\i_MIPS/Register/register[8][21] ), .QN(n552)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][23]  ( .D(\i_MIPS/Register/n875 ), 
        .CK(clk), .RN(n6245), .Q(\i_MIPS/Register/register[8][23] ), .QN(n205)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][26]  ( .D(\i_MIPS/Register/n878 ), 
        .CK(clk), .RN(n6245), .Q(\i_MIPS/Register/register[8][26] ), .QN(n732)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][27]  ( .D(\i_MIPS/Register/n879 ), 
        .CK(clk), .RN(n6245), .Q(\i_MIPS/Register/register[8][27] ), .QN(n740)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][28]  ( .D(\i_MIPS/Register/n880 ), 
        .CK(clk), .RN(n6245), .Q(\i_MIPS/Register/register[8][28] ), .QN(n757)
         );
  DFFRX1 \i_MIPS/Register/register_reg[8][29]  ( .D(\i_MIPS/Register/n881 ), 
        .CK(clk), .RN(n6245), .Q(\i_MIPS/Register/register[8][29] ), .QN(n208)
         );
  DFFRX1 \i_MIPS/Register/register_reg[23][0]  ( .D(\i_MIPS/Register/n372 ), 
        .CK(clk), .RN(n6287), .Q(\i_MIPS/Register/register[23][0] ), .QN(n2380) );
  DFFRX1 \i_MIPS/Register/register_reg[23][1]  ( .D(\i_MIPS/Register/n373 ), 
        .CK(clk), .RN(n6287), .Q(\i_MIPS/Register/register[23][1] ), .QN(n2370) );
  DFFRX1 \i_MIPS/Register/register_reg[23][2]  ( .D(\i_MIPS/Register/n374 ), 
        .CK(clk), .RN(n6287), .Q(\i_MIPS/Register/register[23][2] ), .QN(n2426) );
  DFFRX1 \i_MIPS/Register/register_reg[23][3]  ( .D(\i_MIPS/Register/n375 ), 
        .CK(clk), .RN(n6287), .Q(\i_MIPS/Register/register[23][3] ), .QN(n2389) );
  DFFRX1 \i_MIPS/Register/register_reg[23][4]  ( .D(\i_MIPS/Register/n376 ), 
        .CK(clk), .RN(n6287), .Q(\i_MIPS/Register/register[23][4] ), .QN(n2498) );
  DFFRX1 \i_MIPS/Register/register_reg[23][5]  ( .D(\i_MIPS/Register/n377 ), 
        .CK(clk), .RN(n6287), .Q(\i_MIPS/Register/register[23][5] ), .QN(n2377) );
  DFFRX1 \i_MIPS/Register/register_reg[23][6]  ( .D(\i_MIPS/Register/n378 ), 
        .CK(clk), .RN(n6287), .Q(\i_MIPS/Register/register[23][6] ), .QN(n2510) );
  DFFRX1 \i_MIPS/Register/register_reg[23][7]  ( .D(\i_MIPS/Register/n379 ), 
        .CK(clk), .RN(n6287), .Q(\i_MIPS/Register/register[23][7] ), .QN(n2504) );
  DFFRX1 \i_MIPS/Register/register_reg[23][8]  ( .D(\i_MIPS/Register/n380 ), 
        .CK(clk), .RN(n6286), .Q(\i_MIPS/Register/register[23][8] ), .QN(n313)
         );
  DFFRX1 \i_MIPS/Register/register_reg[23][9]  ( .D(\i_MIPS/Register/n381 ), 
        .CK(clk), .RN(n6286), .Q(\i_MIPS/Register/register[23][9] ), .QN(n251)
         );
  DFFRX1 \i_MIPS/Register/register_reg[23][10]  ( .D(\i_MIPS/Register/n382 ), 
        .CK(clk), .RN(n6286), .Q(\i_MIPS/Register/register[23][10] ), .QN(
        n2405) );
  DFFRX1 \i_MIPS/Register/register_reg[23][11]  ( .D(\i_MIPS/Register/n383 ), 
        .CK(clk), .RN(n6286), .Q(\i_MIPS/Register/register[23][11] ), .QN(
        n2395) );
  DFFRX1 \i_MIPS/Register/register_reg[23][12]  ( .D(\i_MIPS/Register/n384 ), 
        .CK(clk), .RN(n6286), .Q(\i_MIPS/Register/register[23][12] ), .QN(n309) );
  DFFRX1 \i_MIPS/Register/register_reg[23][13]  ( .D(\i_MIPS/Register/n385 ), 
        .CK(clk), .RN(n6286), .Q(\i_MIPS/Register/register[23][13] ), .QN(n315) );
  DFFRX1 \i_MIPS/Register/register_reg[23][15]  ( .D(\i_MIPS/Register/n387 ), 
        .CK(clk), .RN(n6286), .Q(\i_MIPS/Register/register[23][15] ), .QN(
        n2516) );
  DFFRX1 \i_MIPS/Register/register_reg[23][16]  ( .D(\i_MIPS/Register/n388 ), 
        .CK(clk), .RN(n6286), .Q(\i_MIPS/Register/register[23][16] ), .QN(
        n2397) );
  DFFRX1 \i_MIPS/Register/register_reg[23][17]  ( .D(\i_MIPS/Register/n389 ), 
        .CK(clk), .RN(n6286), .Q(\i_MIPS/Register/register[23][17] ), .QN(
        n2475) );
  DFFRX1 \i_MIPS/Register/register_reg[23][18]  ( .D(\i_MIPS/Register/n390 ), 
        .CK(clk), .RN(n6286), .Q(\i_MIPS/Register/register[23][18] ), .QN(
        n2375) );
  DFFRX1 \i_MIPS/Register/register_reg[23][19]  ( .D(\i_MIPS/Register/n391 ), 
        .CK(clk), .RN(n6286), .Q(\i_MIPS/Register/register[23][19] ), .QN(n311) );
  DFFRX1 \i_MIPS/Register/register_reg[23][20]  ( .D(\i_MIPS/Register/n392 ), 
        .CK(clk), .RN(n6285), .Q(\i_MIPS/Register/register[23][20] ), .QN(
        n2176) );
  DFFRX1 \i_MIPS/Register/register_reg[23][21]  ( .D(\i_MIPS/Register/n393 ), 
        .CK(clk), .RN(n6285), .Q(\i_MIPS/Register/register[23][21] ), .QN(
        n2488) );
  DFFRX1 \i_MIPS/Register/register_reg[23][23]  ( .D(\i_MIPS/Register/n395 ), 
        .CK(clk), .RN(n6285), .Q(\i_MIPS/Register/register[23][23] ), .QN(
        n2420) );
  DFFRX1 \i_MIPS/Register/register_reg[23][24]  ( .D(\i_MIPS/Register/n396 ), 
        .CK(clk), .RN(n6285), .Q(\i_MIPS/Register/register[23][24] ), .QN(
        n2367) );
  DFFRX1 \i_MIPS/Register/register_reg[23][25]  ( .D(\i_MIPS/Register/n397 ), 
        .CK(clk), .RN(n6285), .Q(\i_MIPS/Register/register[23][25] ), .QN(
        n2437) );
  DFFRX1 \i_MIPS/Register/register_reg[23][26]  ( .D(\i_MIPS/Register/n398 ), 
        .CK(clk), .RN(n6285), .Q(\i_MIPS/Register/register[23][26] ), .QN(
        n2492) );
  DFFRX1 \i_MIPS/Register/register_reg[23][27]  ( .D(\i_MIPS/Register/n399 ), 
        .CK(clk), .RN(n6285), .Q(\i_MIPS/Register/register[23][27] ), .QN(
        n2439) );
  DFFRX1 \i_MIPS/Register/register_reg[23][28]  ( .D(\i_MIPS/Register/n400 ), 
        .CK(clk), .RN(n6285), .Q(\i_MIPS/Register/register[23][28] ), .QN(
        n2416) );
  DFFRX1 \i_MIPS/Register/register_reg[23][29]  ( .D(\i_MIPS/Register/n401 ), 
        .CK(clk), .RN(n6285), .Q(\i_MIPS/Register/register[23][29] ), .QN(
        n2431) );
  DFFRX1 \i_MIPS/Register/register_reg[21][0]  ( .D(\i_MIPS/Register/n436 ), 
        .CK(clk), .RN(n6282), .Q(\i_MIPS/Register/register[21][0] ), .QN(n917)
         );
  DFFRX1 \i_MIPS/Register/register_reg[21][1]  ( .D(\i_MIPS/Register/n437 ), 
        .CK(clk), .RN(n6282), .Q(\i_MIPS/Register/register[21][1] ), .QN(n2481) );
  DFFRX1 \i_MIPS/Register/register_reg[21][2]  ( .D(\i_MIPS/Register/n438 ), 
        .CK(clk), .RN(n6282), .Q(\i_MIPS/Register/register[21][2] ), .QN(n2515) );
  DFFRX1 \i_MIPS/Register/register_reg[21][3]  ( .D(\i_MIPS/Register/n439 ), 
        .CK(clk), .RN(n6282), .Q(\i_MIPS/Register/register[21][3] ), .QN(n2391) );
  DFFRX1 \i_MIPS/Register/register_reg[21][4]  ( .D(\i_MIPS/Register/n440 ), 
        .CK(clk), .RN(n6281), .Q(\i_MIPS/Register/register[21][4] ), .QN(n2500) );
  DFFRX1 \i_MIPS/Register/register_reg[21][5]  ( .D(\i_MIPS/Register/n441 ), 
        .CK(clk), .RN(n6281), .Q(\i_MIPS/Register/register[21][5] ), .QN(n2379) );
  DFFRX1 \i_MIPS/Register/register_reg[21][6]  ( .D(\i_MIPS/Register/n442 ), 
        .CK(clk), .RN(n6281), .Q(\i_MIPS/Register/register[21][6] ), .QN(n2512) );
  DFFRX1 \i_MIPS/Register/register_reg[21][7]  ( .D(\i_MIPS/Register/n443 ), 
        .CK(clk), .RN(n6281), .Q(\i_MIPS/Register/register[21][7] ), .QN(n2506) );
  DFFRX1 \i_MIPS/Register/register_reg[21][8]  ( .D(\i_MIPS/Register/n444 ), 
        .CK(clk), .RN(n6281), .Q(\i_MIPS/Register/register[21][8] ), .QN(n2490) );
  DFFRX1 \i_MIPS/Register/register_reg[21][9]  ( .D(\i_MIPS/Register/n445 ), 
        .CK(clk), .RN(n6281), .Q(\i_MIPS/Register/register[21][9] ), .QN(n2009) );
  DFFRX1 \i_MIPS/Register/register_reg[21][10]  ( .D(\i_MIPS/Register/n446 ), 
        .CK(clk), .RN(n6281), .Q(\i_MIPS/Register/register[21][10] ), .QN(
        n2407) );
  DFFRX1 \i_MIPS/Register/register_reg[21][11]  ( .D(\i_MIPS/Register/n447 ), 
        .CK(clk), .RN(n6281), .Q(\i_MIPS/Register/register[21][11] ), .QN(n938) );
  DFFRX1 \i_MIPS/Register/register_reg[21][12]  ( .D(\i_MIPS/Register/n448 ), 
        .CK(clk), .RN(n6281), .Q(\i_MIPS/Register/register[21][12] ), .QN(
        n2482) );
  DFFRX1 \i_MIPS/Register/register_reg[21][13]  ( .D(\i_MIPS/Register/n449 ), 
        .CK(clk), .RN(n6281), .Q(\i_MIPS/Register/register[21][13] ), .QN(
        n2411) );
  DFFRX1 \i_MIPS/Register/register_reg[21][15]  ( .D(\i_MIPS/Register/n451 ), 
        .CK(clk), .RN(n6281), .Q(\i_MIPS/Register/register[21][15] ), .QN(
        n2518) );
  DFFRX1 \i_MIPS/Register/register_reg[21][16]  ( .D(\i_MIPS/Register/n452 ), 
        .CK(clk), .RN(n6280), .Q(\i_MIPS/Register/register[21][16] ), .QN(n920) );
  DFFRX1 \i_MIPS/Register/register_reg[21][17]  ( .D(\i_MIPS/Register/n453 ), 
        .CK(clk), .RN(n6280), .Q(\i_MIPS/Register/register[21][17] ), .QN(
        n2477) );
  DFFRX1 \i_MIPS/Register/register_reg[21][18]  ( .D(\i_MIPS/Register/n454 ), 
        .CK(clk), .RN(n6280), .Q(\i_MIPS/Register/register[21][18] ), .QN(n937) );
  DFFRX1 \i_MIPS/Register/register_reg[21][19]  ( .D(\i_MIPS/Register/n455 ), 
        .CK(clk), .RN(n6280), .Q(\i_MIPS/Register/register[21][19] ), .QN(
        n2485) );
  DFFRX1 \i_MIPS/Register/register_reg[21][20]  ( .D(\i_MIPS/Register/n456 ), 
        .CK(clk), .RN(n6280), .Q(\i_MIPS/Register/register[21][20] ), .QN(n939) );
  DFFRX1 \i_MIPS/Register/register_reg[21][21]  ( .D(\i_MIPS/Register/n457 ), 
        .CK(clk), .RN(n6280), .Q(\i_MIPS/Register/register[21][21] ), .QN(n941) );
  DFFRX1 \i_MIPS/Register/register_reg[21][23]  ( .D(\i_MIPS/Register/n459 ), 
        .CK(clk), .RN(n6280), .Q(\i_MIPS/Register/register[21][23] ), .QN(
        n2422) );
  DFFRX1 \i_MIPS/Register/register_reg[21][24]  ( .D(\i_MIPS/Register/n460 ), 
        .CK(clk), .RN(n6280), .Q(\i_MIPS/Register/register[21][24] ), .QN(
        n2369) );
  DFFRX1 \i_MIPS/Register/register_reg[21][25]  ( .D(\i_MIPS/Register/n461 ), 
        .CK(clk), .RN(n6280), .Q(\i_MIPS/Register/register[21][25] ), .QN(
        n2522) );
  DFFRX1 \i_MIPS/Register/register_reg[21][26]  ( .D(\i_MIPS/Register/n462 ), 
        .CK(clk), .RN(n6280), .Q(\i_MIPS/Register/register[21][26] ), .QN(
        n2494) );
  DFFRX1 \i_MIPS/Register/register_reg[21][27]  ( .D(\i_MIPS/Register/n463 ), 
        .CK(clk), .RN(n6280), .Q(\i_MIPS/Register/register[21][27] ), .QN(
        n2523) );
  DFFRX1 \i_MIPS/Register/register_reg[21][28]  ( .D(\i_MIPS/Register/n464 ), 
        .CK(clk), .RN(n6279), .Q(\i_MIPS/Register/register[21][28] ), .QN(
        n2513) );
  DFFRX1 \i_MIPS/Register/register_reg[21][29]  ( .D(\i_MIPS/Register/n465 ), 
        .CK(clk), .RN(n6279), .Q(\i_MIPS/Register/register[21][29] ), .QN(
        n2433) );
  DFFRX1 \i_MIPS/Register/register_reg[20][0]  ( .D(\i_MIPS/Register/n468 ), 
        .CK(clk), .RN(n6279), .Q(\i_MIPS/Register/register[20][0] ), .QN(n2448) );
  DFFRX1 \i_MIPS/Register/register_reg[20][1]  ( .D(\i_MIPS/Register/n469 ), 
        .CK(clk), .RN(n6279), .Q(\i_MIPS/Register/register[20][1] ), .QN(n2450) );
  DFFRX1 \i_MIPS/Register/register_reg[20][2]  ( .D(\i_MIPS/Register/n470 ), 
        .CK(clk), .RN(n6279), .Q(\i_MIPS/Register/register[20][2] ), .QN(n930)
         );
  DFFRX1 \i_MIPS/Register/register_reg[20][3]  ( .D(\i_MIPS/Register/n471 ), 
        .CK(clk), .RN(n6279), .Q(\i_MIPS/Register/register[20][3] ), .QN(n2357) );
  DFFRX1 \i_MIPS/Register/register_reg[20][4]  ( .D(\i_MIPS/Register/n472 ), 
        .CK(clk), .RN(n6279), .Q(\i_MIPS/Register/register[20][4] ), .QN(n2444) );
  DFFRX1 \i_MIPS/Register/register_reg[20][5]  ( .D(\i_MIPS/Register/n473 ), 
        .CK(clk), .RN(n6279), .Q(\i_MIPS/Register/register[20][5] ), .QN(n2349) );
  DFFRX1 \i_MIPS/Register/register_reg[20][6]  ( .D(\i_MIPS/Register/n474 ), 
        .CK(clk), .RN(n6279), .Q(\i_MIPS/Register/register[20][6] ), .QN(n2526) );
  DFFRX1 \i_MIPS/Register/register_reg[20][7]  ( .D(\i_MIPS/Register/n475 ), 
        .CK(clk), .RN(n6279), .Q(\i_MIPS/Register/register[20][7] ), .QN(n2525) );
  DFFRX1 \i_MIPS/Register/register_reg[20][8]  ( .D(\i_MIPS/Register/n476 ), 
        .CK(clk), .RN(n6278), .Q(\i_MIPS/Register/register[20][8] ), .QN(n2451) );
  DFFRX1 \i_MIPS/Register/register_reg[20][9]  ( .D(\i_MIPS/Register/n477 ), 
        .CK(clk), .RN(n6278), .Q(\i_MIPS/Register/register[20][9] ), .QN(n2183) );
  DFFRX1 \i_MIPS/Register/register_reg[20][10]  ( .D(\i_MIPS/Register/n478 ), 
        .CK(clk), .RN(n6278), .Q(\i_MIPS/Register/register[20][10] ), .QN(
        n2345) );
  DFFRX1 \i_MIPS/Register/register_reg[20][11]  ( .D(\i_MIPS/Register/n479 ), 
        .CK(clk), .RN(n6278), .Q(\i_MIPS/Register/register[20][11] ), .QN(
        n2445) );
  DFFRX1 \i_MIPS/Register/register_reg[20][12]  ( .D(\i_MIPS/Register/n480 ), 
        .CK(clk), .RN(n6278), .Q(\i_MIPS/Register/register[20][12] ), .QN(
        n2449) );
  DFFRX1 \i_MIPS/Register/register_reg[20][13]  ( .D(\i_MIPS/Register/n481 ), 
        .CK(clk), .RN(n6278), .Q(\i_MIPS/Register/register[20][13] ), .QN(
        n2474) );
  DFFRX1 \i_MIPS/Register/register_reg[20][16]  ( .D(\i_MIPS/Register/n484 ), 
        .CK(clk), .RN(n6278), .Q(\i_MIPS/Register/register[20][16] ), .QN(
        n2447) );
  DFFRX1 \i_MIPS/Register/register_reg[20][17]  ( .D(\i_MIPS/Register/n485 ), 
        .CK(clk), .RN(n6278), .Q(\i_MIPS/Register/register[20][17] ), .QN(
        n2348) );
  DFFRX1 \i_MIPS/Register/register_reg[20][18]  ( .D(\i_MIPS/Register/n486 ), 
        .CK(clk), .RN(n6278), .Q(\i_MIPS/Register/register[20][18] ), .QN(
        n2042) );
  DFFRX1 \i_MIPS/Register/register_reg[20][19]  ( .D(\i_MIPS/Register/n487 ), 
        .CK(clk), .RN(n6278), .Q(\i_MIPS/Register/register[20][19] ), .QN(
        n2446) );
  DFFRX1 \i_MIPS/Register/register_reg[20][20]  ( .D(\i_MIPS/Register/n488 ), 
        .CK(clk), .RN(n6277), .Q(\i_MIPS/Register/register[20][20] ), .QN(
        n2524) );
  DFFRX1 \i_MIPS/Register/register_reg[20][21]  ( .D(\i_MIPS/Register/n489 ), 
        .CK(clk), .RN(n6277), .Q(\i_MIPS/Register/register[20][21] ), .QN(
        n2051) );
  DFFRX1 \i_MIPS/Register/register_reg[20][23]  ( .D(\i_MIPS/Register/n491 ), 
        .CK(clk), .RN(n6277), .Q(\i_MIPS/Register/register[20][23] ), .QN(n928) );
  DFFRX1 \i_MIPS/Register/register_reg[20][24]  ( .D(\i_MIPS/Register/n492 ), 
        .CK(clk), .RN(n6277), .Q(\i_MIPS/Register/register[20][24] ), .QN(n953) );
  DFFRX1 \i_MIPS/Register/register_reg[20][25]  ( .D(\i_MIPS/Register/n493 ), 
        .CK(clk), .RN(n6277), .Q(\i_MIPS/Register/register[20][25] ), .QN(n951) );
  DFFRX1 \i_MIPS/Register/register_reg[20][26]  ( .D(\i_MIPS/Register/n494 ), 
        .CK(clk), .RN(n6277), .Q(\i_MIPS/Register/register[20][26] ), .QN(
        n2527) );
  DFFRX1 \i_MIPS/Register/register_reg[20][27]  ( .D(\i_MIPS/Register/n495 ), 
        .CK(clk), .RN(n6277), .Q(\i_MIPS/Register/register[20][27] ), .QN(
        n2452) );
  DFFRX1 \i_MIPS/Register/register_reg[20][28]  ( .D(\i_MIPS/Register/n496 ), 
        .CK(clk), .RN(n6277), .Q(\i_MIPS/Register/register[20][28] ), .QN(
        n2528) );
  DFFRX1 \i_MIPS/Register/register_reg[20][29]  ( .D(\i_MIPS/Register/n497 ), 
        .CK(clk), .RN(n6277), .Q(\i_MIPS/Register/register[20][29] ), .QN(n929) );
  DFFRX1 \i_MIPS/Register/register_reg[19][0]  ( .D(\i_MIPS/Register/n500 ), 
        .CK(clk), .RN(n6276), .Q(\i_MIPS/Register/register[19][0] ), .QN(n2381) );
  DFFRX1 \i_MIPS/Register/register_reg[19][1]  ( .D(\i_MIPS/Register/n501 ), 
        .CK(clk), .RN(n6276), .Q(\i_MIPS/Register/register[19][1] ), .QN(n2371) );
  DFFRX1 \i_MIPS/Register/register_reg[19][2]  ( .D(\i_MIPS/Register/n502 ), 
        .CK(clk), .RN(n6276), .Q(\i_MIPS/Register/register[19][2] ), .QN(n2427) );
  DFFRX1 \i_MIPS/Register/register_reg[19][3]  ( .D(\i_MIPS/Register/n503 ), 
        .CK(clk), .RN(n6276), .Q(\i_MIPS/Register/register[19][3] ), .QN(n2390) );
  DFFRX1 \i_MIPS/Register/register_reg[19][4]  ( .D(\i_MIPS/Register/n504 ), 
        .CK(clk), .RN(n6276), .Q(\i_MIPS/Register/register[19][4] ), .QN(n2499) );
  DFFRX1 \i_MIPS/Register/register_reg[19][5]  ( .D(\i_MIPS/Register/n505 ), 
        .CK(clk), .RN(n6276), .Q(\i_MIPS/Register/register[19][5] ), .QN(n2378) );
  DFFRX1 \i_MIPS/Register/register_reg[19][6]  ( .D(\i_MIPS/Register/n506 ), 
        .CK(clk), .RN(n6276), .Q(\i_MIPS/Register/register[19][6] ), .QN(n2511) );
  DFFRX1 \i_MIPS/Register/register_reg[19][7]  ( .D(\i_MIPS/Register/n507 ), 
        .CK(clk), .RN(n6276), .Q(\i_MIPS/Register/register[19][7] ), .QN(n2505) );
  DFFRX1 \i_MIPS/Register/register_reg[19][8]  ( .D(\i_MIPS/Register/n508 ), 
        .CK(clk), .RN(n6276), .Q(\i_MIPS/Register/register[19][8] ), .QN(n924)
         );
  DFFRX1 \i_MIPS/Register/register_reg[19][9]  ( .D(\i_MIPS/Register/n509 ), 
        .CK(clk), .RN(n6276), .Q(\i_MIPS/Register/register[19][9] ), .QN(n392)
         );
  DFFRX1 \i_MIPS/Register/register_reg[19][10]  ( .D(\i_MIPS/Register/n510 ), 
        .CK(clk), .RN(n6276), .Q(\i_MIPS/Register/register[19][10] ), .QN(
        n2406) );
  DFFRX1 \i_MIPS/Register/register_reg[19][11]  ( .D(\i_MIPS/Register/n511 ), 
        .CK(clk), .RN(n6276), .Q(\i_MIPS/Register/register[19][11] ), .QN(
        n2396) );
  DFFRX1 \i_MIPS/Register/register_reg[19][12]  ( .D(\i_MIPS/Register/n512 ), 
        .CK(clk), .RN(n6275), .Q(\i_MIPS/Register/register[19][12] ), .QN(n915) );
  DFFRX1 \i_MIPS/Register/register_reg[19][13]  ( .D(\i_MIPS/Register/n513 ), 
        .CK(clk), .RN(n6275), .Q(\i_MIPS/Register/register[19][13] ), .QN(n926) );
  DFFRX1 \i_MIPS/Register/register_reg[19][15]  ( .D(\i_MIPS/Register/n515 ), 
        .CK(clk), .RN(n6275), .Q(\i_MIPS/Register/register[19][15] ), .QN(
        n2517) );
  DFFRX1 \i_MIPS/Register/register_reg[19][16]  ( .D(\i_MIPS/Register/n516 ), 
        .CK(clk), .RN(n6275), .Q(\i_MIPS/Register/register[19][16] ), .QN(
        n2398) );
  DFFRX1 \i_MIPS/Register/register_reg[19][17]  ( .D(\i_MIPS/Register/n517 ), 
        .CK(clk), .RN(n6275), .Q(\i_MIPS/Register/register[19][17] ), .QN(
        n2476) );
  DFFRX1 \i_MIPS/Register/register_reg[19][18]  ( .D(\i_MIPS/Register/n518 ), 
        .CK(clk), .RN(n6275), .Q(\i_MIPS/Register/register[19][18] ), .QN(
        n2376) );
  DFFRX1 \i_MIPS/Register/register_reg[19][19]  ( .D(\i_MIPS/Register/n519 ), 
        .CK(clk), .RN(n6275), .Q(\i_MIPS/Register/register[19][19] ), .QN(n923) );
  DFFRX1 \i_MIPS/Register/register_reg[19][20]  ( .D(\i_MIPS/Register/n520 ), 
        .CK(clk), .RN(n6275), .Q(\i_MIPS/Register/register[19][20] ), .QN(
        n2484) );
  DFFRX1 \i_MIPS/Register/register_reg[19][21]  ( .D(\i_MIPS/Register/n521 ), 
        .CK(clk), .RN(n6275), .Q(\i_MIPS/Register/register[19][21] ), .QN(
        n2403) );
  DFFRX1 \i_MIPS/Register/register_reg[19][23]  ( .D(\i_MIPS/Register/n523 ), 
        .CK(clk), .RN(n6275), .Q(\i_MIPS/Register/register[19][23] ), .QN(
        n2421) );
  DFFRX1 \i_MIPS/Register/register_reg[19][24]  ( .D(\i_MIPS/Register/n524 ), 
        .CK(clk), .RN(n6274), .Q(\i_MIPS/Register/register[19][24] ), .QN(
        n2368) );
  DFFRX1 \i_MIPS/Register/register_reg[19][25]  ( .D(\i_MIPS/Register/n525 ), 
        .CK(clk), .RN(n6274), .Q(\i_MIPS/Register/register[19][25] ), .QN(
        n2438) );
  DFFRX1 \i_MIPS/Register/register_reg[19][26]  ( .D(\i_MIPS/Register/n526 ), 
        .CK(clk), .RN(n6274), .Q(\i_MIPS/Register/register[19][26] ), .QN(
        n2493) );
  DFFRX1 \i_MIPS/Register/register_reg[19][27]  ( .D(\i_MIPS/Register/n527 ), 
        .CK(clk), .RN(n6274), .Q(\i_MIPS/Register/register[19][27] ), .QN(
        n2440) );
  DFFRX1 \i_MIPS/Register/register_reg[19][28]  ( .D(\i_MIPS/Register/n528 ), 
        .CK(clk), .RN(n6274), .Q(\i_MIPS/Register/register[19][28] ), .QN(
        n2417) );
  DFFRX1 \i_MIPS/Register/register_reg[19][29]  ( .D(\i_MIPS/Register/n529 ), 
        .CK(clk), .RN(n6274), .Q(\i_MIPS/Register/register[19][29] ), .QN(
        n2432) );
  DFFRX1 \i_MIPS/Register/register_reg[17][0]  ( .D(\i_MIPS/Register/n564 ), 
        .CK(clk), .RN(n6271), .Q(\i_MIPS/Register/register[17][0] ), .QN(n2047) );
  DFFRX1 \i_MIPS/Register/register_reg[17][1]  ( .D(\i_MIPS/Register/n565 ), 
        .CK(clk), .RN(n6271), .Q(\i_MIPS/Register/register[17][1] ), .QN(n2455) );
  DFFRX1 \i_MIPS/Register/register_reg[17][2]  ( .D(\i_MIPS/Register/n566 ), 
        .CK(clk), .RN(n6271), .Q(\i_MIPS/Register/register[17][2] ), .QN(n308)
         );
  DFFRX1 \i_MIPS/Register/register_reg[17][3]  ( .D(\i_MIPS/Register/n567 ), 
        .CK(clk), .RN(n6271), .Q(\i_MIPS/Register/register[17][3] ), .QN(n2539) );
  DFFRX1 \i_MIPS/Register/register_reg[17][4]  ( .D(\i_MIPS/Register/n568 ), 
        .CK(clk), .RN(n6271), .Q(\i_MIPS/Register/register[17][4] ), .QN(n2567) );
  DFFRX1 \i_MIPS/Register/register_reg[17][5]  ( .D(\i_MIPS/Register/n569 ), 
        .CK(clk), .RN(n6271), .Q(\i_MIPS/Register/register[17][5] ), .QN(n2366) );
  DFFRX1 \i_MIPS/Register/register_reg[17][6]  ( .D(\i_MIPS/Register/n570 ), 
        .CK(clk), .RN(n6271), .Q(\i_MIPS/Register/register[17][6] ), .QN(n2556) );
  DFFRX1 \i_MIPS/Register/register_reg[17][7]  ( .D(\i_MIPS/Register/n571 ), 
        .CK(clk), .RN(n6271), .Q(\i_MIPS/Register/register[17][7] ), .QN(n2554) );
  DFFRX1 \i_MIPS/Register/register_reg[17][8]  ( .D(\i_MIPS/Register/n572 ), 
        .CK(clk), .RN(n6270), .Q(\i_MIPS/Register/register[17][8] ), .QN(n2559) );
  DFFRX1 \i_MIPS/Register/register_reg[17][9]  ( .D(\i_MIPS/Register/n573 ), 
        .CK(clk), .RN(n6270), .Q(\i_MIPS/Register/register[17][9] ), .QN(n2547) );
  DFFRX1 \i_MIPS/Register/register_reg[17][10]  ( .D(\i_MIPS/Register/n574 ), 
        .CK(clk), .RN(n6270), .Q(\i_MIPS/Register/register[17][10] ), .QN(
        n2460) );
  DFFRX1 \i_MIPS/Register/register_reg[17][11]  ( .D(\i_MIPS/Register/n575 ), 
        .CK(clk), .RN(n6270), .Q(\i_MIPS/Register/register[17][11] ), .QN(
        n2054) );
  DFFRX1 \i_MIPS/Register/register_reg[17][12]  ( .D(\i_MIPS/Register/n576 ), 
        .CK(clk), .RN(n6270), .Q(\i_MIPS/Register/register[17][12] ), .QN(
        n2557) );
  DFFRX1 \i_MIPS/Register/register_reg[17][13]  ( .D(\i_MIPS/Register/n577 ), 
        .CK(clk), .RN(n6270), .Q(\i_MIPS/Register/register[17][13] ), .QN(
        n2172) );
  DFFRX1 \i_MIPS/Register/register_reg[17][15]  ( .D(\i_MIPS/Register/n579 ), 
        .CK(clk), .RN(n6270), .Q(\i_MIPS/Register/register[17][15] ), .QN(n305) );
  DFFRX1 \i_MIPS/Register/register_reg[17][16]  ( .D(\i_MIPS/Register/n580 ), 
        .CK(clk), .RN(n6270), .Q(\i_MIPS/Register/register[17][16] ), .QN(
        n2049) );
  DFFRX1 \i_MIPS/Register/register_reg[17][17]  ( .D(\i_MIPS/Register/n581 ), 
        .CK(clk), .RN(n6270), .Q(\i_MIPS/Register/register[17][17] ), .QN(
        n2565) );
  DFFRX1 \i_MIPS/Register/register_reg[17][18]  ( .D(\i_MIPS/Register/n582 ), 
        .CK(clk), .RN(n6270), .Q(\i_MIPS/Register/register[17][18] ), .QN(
        n2356) );
  DFFRX1 \i_MIPS/Register/register_reg[17][19]  ( .D(\i_MIPS/Register/n583 ), 
        .CK(clk), .RN(n6270), .Q(\i_MIPS/Register/register[17][19] ), .QN(
        n2459) );
  DFFRX1 \i_MIPS/Register/register_reg[17][20]  ( .D(\i_MIPS/Register/n584 ), 
        .CK(clk), .RN(n6269), .Q(\i_MIPS/Register/register[17][20] ), .QN(
        n2052) );
  DFFRX1 \i_MIPS/Register/register_reg[17][21]  ( .D(\i_MIPS/Register/n585 ), 
        .CK(clk), .RN(n6269), .Q(\i_MIPS/Register/register[17][21] ), .QN(
        n2534) );
  DFFRX1 \i_MIPS/Register/register_reg[17][23]  ( .D(\i_MIPS/Register/n587 ), 
        .CK(clk), .RN(n6269), .Q(\i_MIPS/Register/register[17][23] ), .QN(n320) );
  DFFRX1 \i_MIPS/Register/register_reg[17][24]  ( .D(\i_MIPS/Register/n588 ), 
        .CK(clk), .RN(n6269), .Q(\i_MIPS/Register/register[17][24] ), .QN(n323) );
  DFFRX1 \i_MIPS/Register/register_reg[17][25]  ( .D(\i_MIPS/Register/n589 ), 
        .CK(clk), .RN(n6269), .Q(\i_MIPS/Register/register[17][25] ), .QN(n331) );
  DFFRX1 \i_MIPS/Register/register_reg[17][26]  ( .D(\i_MIPS/Register/n590 ), 
        .CK(clk), .RN(n6269), .Q(\i_MIPS/Register/register[17][26] ), .QN(
        n2347) );
  DFFRX1 \i_MIPS/Register/register_reg[17][27]  ( .D(\i_MIPS/Register/n591 ), 
        .CK(clk), .RN(n6269), .Q(\i_MIPS/Register/register[17][27] ), .QN(
        n2553) );
  DFFRX1 \i_MIPS/Register/register_reg[17][28]  ( .D(\i_MIPS/Register/n592 ), 
        .CK(clk), .RN(n6269), .Q(\i_MIPS/Register/register[17][28] ), .QN(
        n2551) );
  DFFRX1 \i_MIPS/Register/register_reg[17][29]  ( .D(\i_MIPS/Register/n593 ), 
        .CK(clk), .RN(n6269), .Q(\i_MIPS/Register/register[17][29] ), .QN(n322) );
  DFFRX1 \i_MIPS/Register/register_reg[16][0]  ( .D(\i_MIPS/Register/n596 ), 
        .CK(clk), .RN(n6268), .Q(\i_MIPS/Register/register[16][0] ), .QN(n2457) );
  DFFRX1 \i_MIPS/Register/register_reg[16][1]  ( .D(\i_MIPS/Register/n597 ), 
        .CK(clk), .RN(n6268), .Q(\i_MIPS/Register/register[16][1] ), .QN(n931)
         );
  DFFRX1 \i_MIPS/Register/register_reg[16][2]  ( .D(\i_MIPS/Register/n598 ), 
        .CK(clk), .RN(n6268), .Q(\i_MIPS/Register/register[16][2] ), .QN(n328)
         );
  DFFRX1 \i_MIPS/Register/register_reg[16][3]  ( .D(\i_MIPS/Register/n599 ), 
        .CK(clk), .RN(n6268), .Q(\i_MIPS/Register/register[16][3] ), .QN(n946)
         );
  DFFRX1 \i_MIPS/Register/register_reg[16][4]  ( .D(\i_MIPS/Register/n600 ), 
        .CK(clk), .RN(n6268), .Q(\i_MIPS/Register/register[16][4] ), .QN(n947)
         );
  DFFRX1 \i_MIPS/Register/register_reg[16][5]  ( .D(\i_MIPS/Register/n601 ), 
        .CK(clk), .RN(n6268), .Q(\i_MIPS/Register/register[16][5] ), .QN(n948)
         );
  DFFRX1 \i_MIPS/Register/register_reg[16][6]  ( .D(\i_MIPS/Register/n602 ), 
        .CK(clk), .RN(n6268), .Q(\i_MIPS/Register/register[16][6] ), .QN(n2571) );
  DFFRX1 \i_MIPS/Register/register_reg[16][7]  ( .D(\i_MIPS/Register/n603 ), 
        .CK(clk), .RN(n6268), .Q(\i_MIPS/Register/register[16][7] ), .QN(n2570) );
  DFFRX1 \i_MIPS/Register/register_reg[16][8]  ( .D(\i_MIPS/Register/n604 ), 
        .CK(clk), .RN(n6268), .Q(\i_MIPS/Register/register[16][8] ), .QN(n2541) );
  DFFRX1 \i_MIPS/Register/register_reg[16][9]  ( .D(\i_MIPS/Register/n605 ), 
        .CK(clk), .RN(n6268), .Q(\i_MIPS/Register/register[16][9] ), .QN(n2362) );
  DFFRX1 \i_MIPS/Register/register_reg[16][10]  ( .D(\i_MIPS/Register/n606 ), 
        .CK(clk), .RN(n6268), .Q(\i_MIPS/Register/register[16][10] ), .QN(
        n2346) );
  DFFRX1 \i_MIPS/Register/register_reg[16][11]  ( .D(\i_MIPS/Register/n607 ), 
        .CK(clk), .RN(n6268), .Q(\i_MIPS/Register/register[16][11] ), .QN(
        n2360) );
  DFFRX1 \i_MIPS/Register/register_reg[16][12]  ( .D(\i_MIPS/Register/n608 ), 
        .CK(clk), .RN(n6267), .Q(\i_MIPS/Register/register[16][12] ), .QN(
        n2543) );
  DFFRX1 \i_MIPS/Register/register_reg[16][13]  ( .D(\i_MIPS/Register/n609 ), 
        .CK(clk), .RN(n6267), .Q(\i_MIPS/Register/register[16][13] ), .QN(
        n2561) );
  DFFRX1 \i_MIPS/Register/register_reg[16][15]  ( .D(\i_MIPS/Register/n611 ), 
        .CK(clk), .RN(n6267), .Q(\i_MIPS/Register/register[16][15] ), .QN(n325) );
  DFFRX1 \i_MIPS/Register/register_reg[16][16]  ( .D(\i_MIPS/Register/n612 ), 
        .CK(clk), .RN(n6267), .Q(\i_MIPS/Register/register[16][16] ), .QN(
        n2533) );
  DFFRX1 \i_MIPS/Register/register_reg[16][17]  ( .D(\i_MIPS/Register/n613 ), 
        .CK(clk), .RN(n6267), .Q(\i_MIPS/Register/register[16][17] ), .QN(n936) );
  DFFRX1 \i_MIPS/Register/register_reg[16][18]  ( .D(\i_MIPS/Register/n614 ), 
        .CK(clk), .RN(n6267), .Q(\i_MIPS/Register/register[16][18] ), .QN(
        n2359) );
  DFFRX1 \i_MIPS/Register/register_reg[16][19]  ( .D(\i_MIPS/Register/n615 ), 
        .CK(clk), .RN(n6267), .Q(\i_MIPS/Register/register[16][19] ), .QN(
        n2453) );
  DFFRX1 \i_MIPS/Register/register_reg[16][20]  ( .D(\i_MIPS/Register/n616 ), 
        .CK(clk), .RN(n6267), .Q(\i_MIPS/Register/register[16][20] ), .QN(
        n2170) );
  DFFRX1 \i_MIPS/Register/register_reg[16][21]  ( .D(\i_MIPS/Register/n617 ), 
        .CK(clk), .RN(n6267), .Q(\i_MIPS/Register/register[16][21] ), .QN(
        n2175) );
  DFFRX1 \i_MIPS/Register/register_reg[16][23]  ( .D(\i_MIPS/Register/n619 ), 
        .CK(clk), .RN(n6267), .Q(\i_MIPS/Register/register[16][23] ), .QN(n318) );
  DFFRX1 \i_MIPS/Register/register_reg[16][24]  ( .D(\i_MIPS/Register/n620 ), 
        .CK(clk), .RN(n6266), .Q(\i_MIPS/Register/register[16][24] ), .QN(n335) );
  DFFRX1 \i_MIPS/Register/register_reg[16][25]  ( .D(\i_MIPS/Register/n621 ), 
        .CK(clk), .RN(n6266), .Q(\i_MIPS/Register/register[16][25] ), .QN(n261) );
  DFFRX1 \i_MIPS/Register/register_reg[16][26]  ( .D(\i_MIPS/Register/n622 ), 
        .CK(clk), .RN(n6266), .Q(\i_MIPS/Register/register[16][26] ), .QN(
        n2564) );
  DFFRX1 \i_MIPS/Register/register_reg[16][27]  ( .D(\i_MIPS/Register/n623 ), 
        .CK(clk), .RN(n6266), .Q(\i_MIPS/Register/register[16][27] ), .QN(
        n2546) );
  DFFRX1 \i_MIPS/Register/register_reg[16][28]  ( .D(\i_MIPS/Register/n624 ), 
        .CK(clk), .RN(n6266), .Q(\i_MIPS/Register/register[16][28] ), .QN(
        n2563) );
  DFFRX1 \i_MIPS/Register/register_reg[16][29]  ( .D(\i_MIPS/Register/n625 ), 
        .CK(clk), .RN(n6266), .Q(\i_MIPS/Register/register[16][29] ), .QN(n326) );
  DFFRX1 \i_MIPS/Register/register_reg[7][0]  ( .D(\i_MIPS/Register/n884 ), 
        .CK(clk), .RN(n6244), .Q(\i_MIPS/Register/register[7][0] ), .QN(n2387)
         );
  DFFRX1 \i_MIPS/Register/register_reg[7][1]  ( .D(\i_MIPS/Register/n885 ), 
        .CK(clk), .RN(n6244), .Q(\i_MIPS/Register/register[7][1] ), .QN(n2372)
         );
  DFFRX1 \i_MIPS/Register/register_reg[7][2]  ( .D(\i_MIPS/Register/n886 ), 
        .CK(clk), .RN(n6244), .Q(\i_MIPS/Register/register[7][2] ), .QN(n2428)
         );
  DFFRX1 \i_MIPS/Register/register_reg[7][3]  ( .D(\i_MIPS/Register/n887 ), 
        .CK(clk), .RN(n6244), .Q(\i_MIPS/Register/register[7][3] ), .QN(n2392)
         );
  DFFRX1 \i_MIPS/Register/register_reg[7][4]  ( .D(\i_MIPS/Register/n888 ), 
        .CK(clk), .RN(n6244), .Q(\i_MIPS/Register/register[7][4] ), .QN(n2501)
         );
  DFFRX1 \i_MIPS/Register/register_reg[7][5]  ( .D(\i_MIPS/Register/n889 ), 
        .CK(clk), .RN(n6244), .Q(\i_MIPS/Register/register[7][5] ), .QN(n2384)
         );
  DFFRX1 \i_MIPS/Register/register_reg[7][6]  ( .D(\i_MIPS/Register/n890 ), 
        .CK(clk), .RN(n6244), .Q(\i_MIPS/Register/register[7][6] ), .QN(n2413)
         );
  DFFRX1 \i_MIPS/Register/register_reg[7][7]  ( .D(\i_MIPS/Register/n891 ), 
        .CK(clk), .RN(n6244), .Q(\i_MIPS/Register/register[7][7] ), .QN(n2507)
         );
  DFFRX1 \i_MIPS/Register/register_reg[7][8]  ( .D(\i_MIPS/Register/n892 ), 
        .CK(clk), .RN(n6244), .Q(\i_MIPS/Register/register[7][8] ), .QN(n314)
         );
  DFFRX1 \i_MIPS/Register/register_reg[7][9]  ( .D(\i_MIPS/Register/n893 ), 
        .CK(clk), .RN(n6244), .Q(\i_MIPS/Register/register[7][9] ), .QN(n252)
         );
  DFFRX1 \i_MIPS/Register/register_reg[7][10]  ( .D(\i_MIPS/Register/n894 ), 
        .CK(clk), .RN(n6244), .Q(\i_MIPS/Register/register[7][10] ), .QN(n2408) );
  DFFRX1 \i_MIPS/Register/register_reg[7][11]  ( .D(\i_MIPS/Register/n895 ), 
        .CK(clk), .RN(n6244), .Q(\i_MIPS/Register/register[7][11] ), .QN(n2399) );
  DFFRX1 \i_MIPS/Register/register_reg[7][12]  ( .D(\i_MIPS/Register/n896 ), 
        .CK(clk), .RN(n6243), .Q(\i_MIPS/Register/register[7][12] ), .QN(n310)
         );
  DFFRX1 \i_MIPS/Register/register_reg[7][13]  ( .D(\i_MIPS/Register/n897 ), 
        .CK(clk), .RN(n6243), .Q(\i_MIPS/Register/register[7][13] ), .QN(n316)
         );
  DFFRX1 \i_MIPS/Register/register_reg[7][15]  ( .D(\i_MIPS/Register/n899 ), 
        .CK(clk), .RN(n6243), .Q(\i_MIPS/Register/register[7][15] ), .QN(n2519) );
  DFFRX1 \i_MIPS/Register/register_reg[7][16]  ( .D(\i_MIPS/Register/n900 ), 
        .CK(clk), .RN(n6243), .Q(\i_MIPS/Register/register[7][16] ), .QN(n2401) );
  DFFRX1 \i_MIPS/Register/register_reg[7][17]  ( .D(\i_MIPS/Register/n901 ), 
        .CK(clk), .RN(n6243), .Q(\i_MIPS/Register/register[7][17] ), .QN(n2478) );
  DFFRX1 \i_MIPS/Register/register_reg[7][18]  ( .D(\i_MIPS/Register/n902 ), 
        .CK(clk), .RN(n6243), .Q(\i_MIPS/Register/register[7][18] ), .QN(n2382) );
  DFFRX1 \i_MIPS/Register/register_reg[7][19]  ( .D(\i_MIPS/Register/n903 ), 
        .CK(clk), .RN(n6243), .Q(\i_MIPS/Register/register[7][19] ), .QN(n312)
         );
  DFFRX1 \i_MIPS/Register/register_reg[7][20]  ( .D(\i_MIPS/Register/n904 ), 
        .CK(clk), .RN(n6243), .Q(\i_MIPS/Register/register[7][20] ), .QN(n2486) );
  DFFRX1 \i_MIPS/Register/register_reg[7][21]  ( .D(\i_MIPS/Register/n905 ), 
        .CK(clk), .RN(n6243), .Q(\i_MIPS/Register/register[7][21] ), .QN(n2489) );
  DFFRX1 \i_MIPS/Register/register_reg[7][23]  ( .D(\i_MIPS/Register/n907 ), 
        .CK(clk), .RN(n6243), .Q(\i_MIPS/Register/register[7][23] ), .QN(n2423) );
  DFFRX1 \i_MIPS/Register/register_reg[7][24]  ( .D(\i_MIPS/Register/n908 ), 
        .CK(clk), .RN(n6242), .Q(\i_MIPS/Register/register[7][24] ), .QN(n2572) );
  DFFRX1 \i_MIPS/Register/register_reg[7][25]  ( .D(\i_MIPS/Register/n909 ), 
        .CK(clk), .RN(n6242), .Q(\i_MIPS/Register/register[7][25] ), .QN(n2575) );
  DFFRX1 \i_MIPS/Register/register_reg[7][26]  ( .D(\i_MIPS/Register/n910 ), 
        .CK(clk), .RN(n6242), .Q(\i_MIPS/Register/register[7][26] ), .QN(n2495) );
  DFFRX1 \i_MIPS/Register/register_reg[7][27]  ( .D(\i_MIPS/Register/n911 ), 
        .CK(clk), .RN(n6242), .Q(\i_MIPS/Register/register[7][27] ), .QN(n2441) );
  DFFRX1 \i_MIPS/Register/register_reg[7][28]  ( .D(\i_MIPS/Register/n912 ), 
        .CK(clk), .RN(n6242), .Q(\i_MIPS/Register/register[7][28] ), .QN(n2418) );
  DFFRX1 \i_MIPS/Register/register_reg[7][29]  ( .D(\i_MIPS/Register/n913 ), 
        .CK(clk), .RN(n6242), .Q(\i_MIPS/Register/register[7][29] ), .QN(n2434) );
  DFFRX1 \i_MIPS/Register/register_reg[5][0]  ( .D(\i_MIPS/Register/n948 ), 
        .CK(clk), .RN(n6239), .Q(\i_MIPS/Register/register[5][0] ), .QN(n919)
         );
  DFFRX1 \i_MIPS/Register/register_reg[5][1]  ( .D(\i_MIPS/Register/n949 ), 
        .CK(clk), .RN(n6239), .Q(\i_MIPS/Register/register[5][1] ), .QN(n2374)
         );
  DFFRX1 \i_MIPS/Register/register_reg[5][2]  ( .D(\i_MIPS/Register/n950 ), 
        .CK(clk), .RN(n6239), .Q(\i_MIPS/Register/register[5][2] ), .QN(n2430)
         );
  DFFRX1 \i_MIPS/Register/register_reg[5][3]  ( .D(\i_MIPS/Register/n951 ), 
        .CK(clk), .RN(n6239), .Q(\i_MIPS/Register/register[5][3] ), .QN(n2394)
         );
  DFFRX1 \i_MIPS/Register/register_reg[5][4]  ( .D(\i_MIPS/Register/n952 ), 
        .CK(clk), .RN(n6239), .Q(\i_MIPS/Register/register[5][4] ), .QN(n2503)
         );
  DFFRX1 \i_MIPS/Register/register_reg[5][5]  ( .D(\i_MIPS/Register/n953 ), 
        .CK(clk), .RN(n6239), .Q(\i_MIPS/Register/register[5][5] ), .QN(n2386)
         );
  DFFRX1 \i_MIPS/Register/register_reg[5][6]  ( .D(\i_MIPS/Register/n954 ), 
        .CK(clk), .RN(n6239), .Q(\i_MIPS/Register/register[5][6] ), .QN(n2415)
         );
  DFFRX1 \i_MIPS/Register/register_reg[5][7]  ( .D(\i_MIPS/Register/n955 ), 
        .CK(clk), .RN(n6239), .Q(\i_MIPS/Register/register[5][7] ), .QN(n2509)
         );
  DFFRX1 \i_MIPS/Register/register_reg[5][8]  ( .D(\i_MIPS/Register/n956 ), 
        .CK(clk), .RN(n6238), .Q(\i_MIPS/Register/register[5][8] ), .QN(n2491)
         );
  DFFRX1 \i_MIPS/Register/register_reg[5][9]  ( .D(\i_MIPS/Register/n957 ), 
        .CK(clk), .RN(n6238), .Q(\i_MIPS/Register/register[5][9] ), .QN(n2010)
         );
  DFFRX1 \i_MIPS/Register/register_reg[5][10]  ( .D(\i_MIPS/Register/n958 ), 
        .CK(clk), .RN(n6238), .Q(\i_MIPS/Register/register[5][10] ), .QN(n2410) );
  DFFRX1 \i_MIPS/Register/register_reg[5][11]  ( .D(\i_MIPS/Register/n959 ), 
        .CK(clk), .RN(n6238), .Q(\i_MIPS/Register/register[5][11] ), .QN(n921)
         );
  DFFRX1 \i_MIPS/Register/register_reg[5][12]  ( .D(\i_MIPS/Register/n960 ), 
        .CK(clk), .RN(n6238), .Q(\i_MIPS/Register/register[5][12] ), .QN(n2483) );
  DFFRX1 \i_MIPS/Register/register_reg[5][13]  ( .D(\i_MIPS/Register/n961 ), 
        .CK(clk), .RN(n6238), .Q(\i_MIPS/Register/register[5][13] ), .QN(n2412) );
  DFFRX1 \i_MIPS/Register/register_reg[5][15]  ( .D(\i_MIPS/Register/n963 ), 
        .CK(clk), .RN(n6238), .Q(\i_MIPS/Register/register[5][15] ), .QN(n2521) );
  DFFRX1 \i_MIPS/Register/register_reg[5][16]  ( .D(\i_MIPS/Register/n964 ), 
        .CK(clk), .RN(n6238), .Q(\i_MIPS/Register/register[5][16] ), .QN(n922)
         );
  DFFRX1 \i_MIPS/Register/register_reg[5][17]  ( .D(\i_MIPS/Register/n965 ), 
        .CK(clk), .RN(n6238), .Q(\i_MIPS/Register/register[5][17] ), .QN(n2480) );
  DFFRX1 \i_MIPS/Register/register_reg[5][18]  ( .D(\i_MIPS/Register/n966 ), 
        .CK(clk), .RN(n6238), .Q(\i_MIPS/Register/register[5][18] ), .QN(n918)
         );
  DFFRX1 \i_MIPS/Register/register_reg[5][19]  ( .D(\i_MIPS/Register/n967 ), 
        .CK(clk), .RN(n6238), .Q(\i_MIPS/Register/register[5][19] ), .QN(n2173) );
  DFFRX1 \i_MIPS/Register/register_reg[5][20]  ( .D(\i_MIPS/Register/n968 ), 
        .CK(clk), .RN(n6237), .Q(\i_MIPS/Register/register[5][20] ), .QN(n940)
         );
  DFFRX1 \i_MIPS/Register/register_reg[5][21]  ( .D(\i_MIPS/Register/n969 ), 
        .CK(clk), .RN(n6237), .Q(\i_MIPS/Register/register[5][21] ), .QN(n942)
         );
  DFFRX1 \i_MIPS/Register/register_reg[5][23]  ( .D(\i_MIPS/Register/n971 ), 
        .CK(clk), .RN(n6237), .Q(\i_MIPS/Register/register[5][23] ), .QN(n2425) );
  DFFRX1 \i_MIPS/Register/register_reg[5][24]  ( .D(\i_MIPS/Register/n972 ), 
        .CK(clk), .RN(n6237), .Q(\i_MIPS/Register/register[5][24] ), .QN(n2574) );
  DFFRX1 \i_MIPS/Register/register_reg[5][25]  ( .D(\i_MIPS/Register/n973 ), 
        .CK(clk), .RN(n6237), .Q(\i_MIPS/Register/register[5][25] ), .QN(n2577) );
  DFFRX1 \i_MIPS/Register/register_reg[5][26]  ( .D(\i_MIPS/Register/n974 ), 
        .CK(clk), .RN(n6237), .Q(\i_MIPS/Register/register[5][26] ), .QN(n2497) );
  DFFRX1 \i_MIPS/Register/register_reg[5][27]  ( .D(\i_MIPS/Register/n975 ), 
        .CK(clk), .RN(n6237), .Q(\i_MIPS/Register/register[5][27] ), .QN(n2443) );
  DFFRX1 \i_MIPS/Register/register_reg[5][28]  ( .D(\i_MIPS/Register/n976 ), 
        .CK(clk), .RN(n6237), .Q(\i_MIPS/Register/register[5][28] ), .QN(n2514) );
  DFFRX1 \i_MIPS/Register/register_reg[5][29]  ( .D(\i_MIPS/Register/n977 ), 
        .CK(clk), .RN(n6237), .Q(\i_MIPS/Register/register[5][29] ), .QN(n2436) );
  DFFRX1 \i_MIPS/Register/register_reg[4][0]  ( .D(\i_MIPS/Register/n980 ), 
        .CK(clk), .RN(n6236), .Q(\i_MIPS/Register/register[4][0] ), .QN(n2466)
         );
  DFFRX1 \i_MIPS/Register/register_reg[4][1]  ( .D(\i_MIPS/Register/n981 ), 
        .CK(clk), .RN(n6236), .Q(\i_MIPS/Register/register[4][1] ), .QN(n2468)
         );
  DFFRX1 \i_MIPS/Register/register_reg[4][2]  ( .D(\i_MIPS/Register/n982 ), 
        .CK(clk), .RN(n6236), .Q(\i_MIPS/Register/register[4][2] ), .QN(n935)
         );
  DFFRX1 \i_MIPS/Register/register_reg[4][3]  ( .D(\i_MIPS/Register/n983 ), 
        .CK(clk), .RN(n6236), .Q(\i_MIPS/Register/register[4][3] ), .QN(n2358)
         );
  DFFRX1 \i_MIPS/Register/register_reg[4][4]  ( .D(\i_MIPS/Register/n984 ), 
        .CK(clk), .RN(n6236), .Q(\i_MIPS/Register/register[4][4] ), .QN(n2462)
         );
  DFFRX1 \i_MIPS/Register/register_reg[4][5]  ( .D(\i_MIPS/Register/n985 ), 
        .CK(clk), .RN(n6236), .Q(\i_MIPS/Register/register[4][5] ), .QN(n2351)
         );
  DFFRX1 \i_MIPS/Register/register_reg[4][6]  ( .D(\i_MIPS/Register/n986 ), 
        .CK(clk), .RN(n6236), .Q(\i_MIPS/Register/register[4][6] ), .QN(n2470)
         );
  DFFRX1 \i_MIPS/Register/register_reg[4][7]  ( .D(\i_MIPS/Register/n987 ), 
        .CK(clk), .RN(n6236), .Q(\i_MIPS/Register/register[4][7] ), .QN(n2530)
         );
  DFFRX1 \i_MIPS/Register/register_reg[4][8]  ( .D(\i_MIPS/Register/n988 ), 
        .CK(clk), .RN(n6236), .Q(\i_MIPS/Register/register[4][8] ), .QN(n2469)
         );
  DFFRX1 \i_MIPS/Register/register_reg[4][9]  ( .D(\i_MIPS/Register/n989 ), 
        .CK(clk), .RN(n6236), .Q(\i_MIPS/Register/register[4][9] ), .QN(n2182)
         );
  DFFRX1 \i_MIPS/Register/register_reg[4][10]  ( .D(\i_MIPS/Register/n990 ), 
        .CK(clk), .RN(n6236), .Q(\i_MIPS/Register/register[4][10] ), .QN(n2344) );
  DFFRX1 \i_MIPS/Register/register_reg[4][11]  ( .D(\i_MIPS/Register/n991 ), 
        .CK(clk), .RN(n6236), .Q(\i_MIPS/Register/register[4][11] ), .QN(n2463) );
  DFFRX1 \i_MIPS/Register/register_reg[4][12]  ( .D(\i_MIPS/Register/n992 ), 
        .CK(clk), .RN(n6235), .Q(\i_MIPS/Register/register[4][12] ), .QN(n2467) );
  DFFRX1 \i_MIPS/Register/register_reg[4][13]  ( .D(\i_MIPS/Register/n993 ), 
        .CK(clk), .RN(n6235), .Q(\i_MIPS/Register/register[4][13] ), .QN(n2472) );
  DFFRX1 \i_MIPS/Register/register_reg[4][16]  ( .D(\i_MIPS/Register/n996 ), 
        .CK(clk), .RN(n6235), .Q(\i_MIPS/Register/register[4][16] ), .QN(n2465) );
  DFFRX1 \i_MIPS/Register/register_reg[4][17]  ( .D(\i_MIPS/Register/n997 ), 
        .CK(clk), .RN(n6235), .Q(\i_MIPS/Register/register[4][17] ), .QN(n2350) );
  DFFRX1 \i_MIPS/Register/register_reg[4][18]  ( .D(\i_MIPS/Register/n998 ), 
        .CK(clk), .RN(n6235), .Q(\i_MIPS/Register/register[4][18] ), .QN(n2043) );
  DFFRX1 \i_MIPS/Register/register_reg[4][19]  ( .D(\i_MIPS/Register/n999 ), 
        .CK(clk), .RN(n6235), .Q(\i_MIPS/Register/register[4][19] ), .QN(n2464) );
  DFFRX1 \i_MIPS/Register/register_reg[4][20]  ( .D(\i_MIPS/Register/n1000 ), 
        .CK(clk), .RN(n6235), .Q(\i_MIPS/Register/register[4][20] ), .QN(n2045) );
  DFFRX1 \i_MIPS/Register/register_reg[4][21]  ( .D(\i_MIPS/Register/n1001 ), 
        .CK(clk), .RN(n6235), .Q(\i_MIPS/Register/register[4][21] ), .QN(n2044) );
  DFFRX1 \i_MIPS/Register/register_reg[4][23]  ( .D(\i_MIPS/Register/n1003 ), 
        .CK(clk), .RN(n6235), .Q(\i_MIPS/Register/register[4][23] ), .QN(n933)
         );
  DFFRX1 \i_MIPS/Register/register_reg[4][24]  ( .D(\i_MIPS/Register/n1004 ), 
        .CK(clk), .RN(n6234), .Q(\i_MIPS/Register/register[4][24] ), .QN(n329)
         );
  DFFRX1 \i_MIPS/Register/register_reg[4][25]  ( .D(\i_MIPS/Register/n1005 ), 
        .CK(clk), .RN(n6234), .Q(\i_MIPS/Register/register[4][25] ), .QN(n952)
         );
  DFFRX1 \i_MIPS/Register/register_reg[4][26]  ( .D(\i_MIPS/Register/n1006 ), 
        .CK(clk), .RN(n6234), .Q(\i_MIPS/Register/register[4][26] ), .QN(n2471) );
  DFFRX1 \i_MIPS/Register/register_reg[4][27]  ( .D(\i_MIPS/Register/n1007 ), 
        .CK(clk), .RN(n6234), .Q(\i_MIPS/Register/register[4][27] ), .QN(n2473) );
  DFFRX1 \i_MIPS/Register/register_reg[4][28]  ( .D(\i_MIPS/Register/n1008 ), 
        .CK(clk), .RN(n6234), .Q(\i_MIPS/Register/register[4][28] ), .QN(n2531) );
  DFFRX1 \i_MIPS/Register/register_reg[4][29]  ( .D(\i_MIPS/Register/n1009 ), 
        .CK(clk), .RN(n6234), .Q(\i_MIPS/Register/register[4][29] ), .QN(n934)
         );
  DFFRX1 \i_MIPS/Register/register_reg[3][0]  ( .D(\i_MIPS/Register/n1012 ), 
        .CK(clk), .RN(n6234), .Q(\i_MIPS/Register/register[3][0] ), .QN(n2388)
         );
  DFFRX1 \i_MIPS/Register/register_reg[3][1]  ( .D(\i_MIPS/Register/n1013 ), 
        .CK(clk), .RN(n6234), .Q(\i_MIPS/Register/register[3][1] ), .QN(n2373)
         );
  DFFRX1 \i_MIPS/Register/register_reg[3][2]  ( .D(\i_MIPS/Register/n1014 ), 
        .CK(clk), .RN(n6234), .Q(\i_MIPS/Register/register[3][2] ), .QN(n2429)
         );
  DFFRX1 \i_MIPS/Register/register_reg[3][3]  ( .D(\i_MIPS/Register/n1015 ), 
        .CK(clk), .RN(n6234), .Q(\i_MIPS/Register/register[3][3] ), .QN(n2393)
         );
  DFFRX1 \i_MIPS/Register/register_reg[3][4]  ( .D(\i_MIPS/Register/n1016 ), 
        .CK(clk), .RN(n6233), .Q(\i_MIPS/Register/register[3][4] ), .QN(n2502)
         );
  DFFRX1 \i_MIPS/Register/register_reg[3][5]  ( .D(\i_MIPS/Register/n1017 ), 
        .CK(clk), .RN(n6233), .Q(\i_MIPS/Register/register[3][5] ), .QN(n2385)
         );
  DFFRX1 \i_MIPS/Register/register_reg[3][6]  ( .D(\i_MIPS/Register/n1018 ), 
        .CK(clk), .RN(n6233), .Q(\i_MIPS/Register/register[3][6] ), .QN(n2414)
         );
  DFFRX1 \i_MIPS/Register/register_reg[3][7]  ( .D(\i_MIPS/Register/n1019 ), 
        .CK(clk), .RN(n6233), .Q(\i_MIPS/Register/register[3][7] ), .QN(n2508)
         );
  DFFRX1 \i_MIPS/Register/register_reg[3][8]  ( .D(\i_MIPS/Register/n1020 ), 
        .CK(clk), .RN(n6233), .Q(\i_MIPS/Register/register[3][8] ), .QN(n925)
         );
  DFFRX1 \i_MIPS/Register/register_reg[3][9]  ( .D(\i_MIPS/Register/n1021 ), 
        .CK(clk), .RN(n6233), .Q(\i_MIPS/Register/register[3][9] ), .QN(n393)
         );
  DFFRX1 \i_MIPS/Register/register_reg[3][10]  ( .D(\i_MIPS/Register/n1022 ), 
        .CK(clk), .RN(n6233), .Q(\i_MIPS/Register/register[3][10] ), .QN(n2409) );
  DFFRX1 \i_MIPS/Register/register_reg[3][11]  ( .D(\i_MIPS/Register/n1023 ), 
        .CK(clk), .RN(n6233), .Q(\i_MIPS/Register/register[3][11] ), .QN(n2400) );
  DFFRX1 \i_MIPS/Register/register_reg[3][12]  ( .D(\i_MIPS/Register/n1024 ), 
        .CK(clk), .RN(n6233), .Q(\i_MIPS/Register/register[3][12] ), .QN(n916)
         );
  DFFRX1 \i_MIPS/Register/register_reg[3][13]  ( .D(\i_MIPS/Register/n1025 ), 
        .CK(clk), .RN(n6233), .Q(\i_MIPS/Register/register[3][13] ), .QN(n927)
         );
  DFFRX1 \i_MIPS/Register/register_reg[3][15]  ( .D(\i_MIPS/Register/n1027 ), 
        .CK(clk), .RN(n6233), .Q(\i_MIPS/Register/register[3][15] ), .QN(n2520) );
  DFFRX1 \i_MIPS/Register/register_reg[3][16]  ( .D(\i_MIPS/Register/n1028 ), 
        .CK(clk), .RN(n6232), .Q(\i_MIPS/Register/register[3][16] ), .QN(n2402) );
  DFFRX1 \i_MIPS/Register/register_reg[3][17]  ( .D(\i_MIPS/Register/n1029 ), 
        .CK(clk), .RN(n6232), .Q(\i_MIPS/Register/register[3][17] ), .QN(n2479) );
  DFFRX1 \i_MIPS/Register/register_reg[3][18]  ( .D(\i_MIPS/Register/n1030 ), 
        .CK(clk), .RN(n6232), .Q(\i_MIPS/Register/register[3][18] ), .QN(n2383) );
  DFFRX1 \i_MIPS/Register/register_reg[3][19]  ( .D(\i_MIPS/Register/n1031 ), 
        .CK(clk), .RN(n6232), .Q(\i_MIPS/Register/register[3][19] ), .QN(n429)
         );
  DFFRX1 \i_MIPS/Register/register_reg[3][20]  ( .D(\i_MIPS/Register/n1032 ), 
        .CK(clk), .RN(n6232), .Q(\i_MIPS/Register/register[3][20] ), .QN(n2487) );
  DFFRX1 \i_MIPS/Register/register_reg[3][21]  ( .D(\i_MIPS/Register/n1033 ), 
        .CK(clk), .RN(n6232), .Q(\i_MIPS/Register/register[3][21] ), .QN(n2404) );
  DFFRX1 \i_MIPS/Register/register_reg[3][23]  ( .D(\i_MIPS/Register/n1035 ), 
        .CK(clk), .RN(n6232), .Q(\i_MIPS/Register/register[3][23] ), .QN(n2424) );
  DFFRX1 \i_MIPS/Register/register_reg[3][24]  ( .D(\i_MIPS/Register/n1036 ), 
        .CK(clk), .RN(n6232), .Q(\i_MIPS/Register/register[3][24] ), .QN(n2573) );
  DFFRX1 \i_MIPS/Register/register_reg[3][25]  ( .D(\i_MIPS/Register/n1037 ), 
        .CK(clk), .RN(n6232), .Q(\i_MIPS/Register/register[3][25] ), .QN(n2576) );
  DFFRX1 \i_MIPS/Register/register_reg[3][26]  ( .D(\i_MIPS/Register/n1038 ), 
        .CK(clk), .RN(n6232), .Q(\i_MIPS/Register/register[3][26] ), .QN(n2496) );
  DFFRX1 \i_MIPS/Register/register_reg[3][27]  ( .D(\i_MIPS/Register/n1039 ), 
        .CK(clk), .RN(n6232), .Q(\i_MIPS/Register/register[3][27] ), .QN(n2442) );
  DFFRX1 \i_MIPS/Register/register_reg[3][28]  ( .D(\i_MIPS/Register/n1040 ), 
        .CK(clk), .RN(n6231), .Q(\i_MIPS/Register/register[3][28] ), .QN(n2419) );
  DFFRX1 \i_MIPS/Register/register_reg[3][29]  ( .D(\i_MIPS/Register/n1041 ), 
        .CK(clk), .RN(n6231), .Q(\i_MIPS/Register/register[3][29] ), .QN(n2435) );
  DFFRX1 \i_MIPS/Register/register_reg[1][0]  ( .D(\i_MIPS/Register/n1076 ), 
        .CK(clk), .RN(n6228), .Q(\i_MIPS/Register/register[1][0] ), .QN(n2048)
         );
  DFFRX1 \i_MIPS/Register/register_reg[1][1]  ( .D(\i_MIPS/Register/n1077 ), 
        .CK(clk), .RN(n6228), .Q(\i_MIPS/Register/register[1][1] ), .QN(n2456)
         );
  DFFRX1 \i_MIPS/Register/register_reg[1][2]  ( .D(\i_MIPS/Register/n1078 ), 
        .CK(clk), .RN(n6228), .Q(\i_MIPS/Register/register[1][2] ), .QN(n307)
         );
  DFFRX1 \i_MIPS/Register/register_reg[1][3]  ( .D(\i_MIPS/Register/n1079 ), 
        .CK(clk), .RN(n6228), .Q(\i_MIPS/Register/register[1][3] ), .QN(n2540)
         );
  DFFRX1 \i_MIPS/Register/register_reg[1][4]  ( .D(\i_MIPS/Register/n1080 ), 
        .CK(clk), .RN(n6228), .Q(\i_MIPS/Register/register[1][4] ), .QN(n2568)
         );
  DFFRX1 \i_MIPS/Register/register_reg[1][5]  ( .D(\i_MIPS/Register/n1081 ), 
        .CK(clk), .RN(n6228), .Q(\i_MIPS/Register/register[1][5] ), .QN(n2548)
         );
  DFFRX1 \i_MIPS/Register/register_reg[1][6]  ( .D(\i_MIPS/Register/n1082 ), 
        .CK(clk), .RN(n6228), .Q(\i_MIPS/Register/register[1][6] ), .QN(n2536)
         );
  DFFRX1 \i_MIPS/Register/register_reg[1][7]  ( .D(\i_MIPS/Register/n1083 ), 
        .CK(clk), .RN(n6228), .Q(\i_MIPS/Register/register[1][7] ), .QN(n2555)
         );
  DFFRX1 \i_MIPS/Register/register_reg[1][8]  ( .D(\i_MIPS/Register/n1084 ), 
        .CK(clk), .RN(n6228), .Q(\i_MIPS/Register/register[1][8] ), .QN(n2560)
         );
  DFFRX1 \i_MIPS/Register/register_reg[1][9]  ( .D(\i_MIPS/Register/n1085 ), 
        .CK(clk), .RN(n6228), .Q(\i_MIPS/Register/register[1][9] ), .QN(n2011)
         );
  DFFRX1 \i_MIPS/Register/register_reg[1][10]  ( .D(\i_MIPS/Register/n1086 ), 
        .CK(clk), .RN(n6228), .Q(\i_MIPS/Register/register[1][10] ), .QN(n2461) );
  DFFRX1 \i_MIPS/Register/register_reg[1][11]  ( .D(\i_MIPS/Register/n1087 ), 
        .CK(clk), .RN(n6228), .Q(\i_MIPS/Register/register[1][11] ), .QN(n2364) );
  DFFRX1 \i_MIPS/Register/register_reg[1][12]  ( .D(\i_MIPS/Register/n1088 ), 
        .CK(clk), .RN(n6227), .Q(\i_MIPS/Register/register[1][12] ), .QN(n2558) );
  DFFRX1 \i_MIPS/Register/register_reg[1][13]  ( .D(\i_MIPS/Register/n1089 ), 
        .CK(clk), .RN(n6227), .Q(\i_MIPS/Register/register[1][13] ), .QN(n2549) );
  DFFRX1 \i_MIPS/Register/register_reg[1][15]  ( .D(\i_MIPS/Register/n1091 ), 
        .CK(clk), .RN(n6227), .Q(\i_MIPS/Register/register[1][15] ), .QN(n304)
         );
  DFFRX1 \i_MIPS/Register/register_reg[1][16]  ( .D(\i_MIPS/Register/n1092 ), 
        .CK(clk), .RN(n6227), .Q(\i_MIPS/Register/register[1][16] ), .QN(n2050) );
  DFFRX1 \i_MIPS/Register/register_reg[1][17]  ( .D(\i_MIPS/Register/n1093 ), 
        .CK(clk), .RN(n6227), .Q(\i_MIPS/Register/register[1][17] ), .QN(n2566) );
  DFFRX1 \i_MIPS/Register/register_reg[1][18]  ( .D(\i_MIPS/Register/n1094 ), 
        .CK(clk), .RN(n6227), .Q(\i_MIPS/Register/register[1][18] ), .QN(n2365) );
  DFFRX1 \i_MIPS/Register/register_reg[1][19]  ( .D(\i_MIPS/Register/n1095 ), 
        .CK(clk), .RN(n6227), .Q(\i_MIPS/Register/register[1][19] ), .QN(n2174) );
  DFFRX1 \i_MIPS/Register/register_reg[1][20]  ( .D(\i_MIPS/Register/n1096 ), 
        .CK(clk), .RN(n6227), .Q(\i_MIPS/Register/register[1][20] ), .QN(n2053) );
  DFFRX1 \i_MIPS/Register/register_reg[1][21]  ( .D(\i_MIPS/Register/n1097 ), 
        .CK(clk), .RN(n6227), .Q(\i_MIPS/Register/register[1][21] ), .QN(n2046) );
  DFFRX1 \i_MIPS/Register/register_reg[1][23]  ( .D(\i_MIPS/Register/n1099 ), 
        .CK(clk), .RN(n6227), .Q(\i_MIPS/Register/register[1][23] ), .QN(n321)
         );
  DFFRX1 \i_MIPS/Register/register_reg[1][24]  ( .D(\i_MIPS/Register/n1100 ), 
        .CK(clk), .RN(n6226), .Q(\i_MIPS/Register/register[1][24] ), .QN(n332)
         );
  DFFRX1 \i_MIPS/Register/register_reg[1][25]  ( .D(\i_MIPS/Register/n1101 ), 
        .CK(clk), .RN(n6226), .Q(\i_MIPS/Register/register[1][25] ), .QN(n330)
         );
  DFFRX1 \i_MIPS/Register/register_reg[1][26]  ( .D(\i_MIPS/Register/n1102 ), 
        .CK(clk), .RN(n6226), .Q(\i_MIPS/Register/register[1][26] ), .QN(n2529) );
  DFFRX1 \i_MIPS/Register/register_reg[1][27]  ( .D(\i_MIPS/Register/n1103 ), 
        .CK(clk), .RN(n6226), .Q(\i_MIPS/Register/register[1][27] ), .QN(n2535) );
  DFFRX1 \i_MIPS/Register/register_reg[1][28]  ( .D(\i_MIPS/Register/n1104 ), 
        .CK(clk), .RN(n6226), .Q(\i_MIPS/Register/register[1][28] ), .QN(n2552) );
  DFFRX1 \i_MIPS/Register/register_reg[1][29]  ( .D(\i_MIPS/Register/n1105 ), 
        .CK(clk), .RN(n6226), .Q(\i_MIPS/Register/register[1][29] ), .QN(n306)
         );
  DFFRX1 \i_MIPS/Register/register_reg[0][0]  ( .D(\i_MIPS/Register/n1108 ), 
        .CK(clk), .RN(n6226), .Q(\i_MIPS/Register/register[0][0] ), .QN(n2458)
         );
  DFFRX1 \i_MIPS/Register/register_reg[0][1]  ( .D(\i_MIPS/Register/n1109 ), 
        .CK(clk), .RN(n6226), .Q(\i_MIPS/Register/register[0][1] ), .QN(n932)
         );
  DFFRX1 \i_MIPS/Register/register_reg[0][2]  ( .D(\i_MIPS/Register/n1110 ), 
        .CK(clk), .RN(n6226), .Q(\i_MIPS/Register/register[0][2] ), .QN(n327)
         );
  DFFRX1 \i_MIPS/Register/register_reg[0][3]  ( .D(\i_MIPS/Register/n1111 ), 
        .CK(clk), .RN(n6226), .Q(\i_MIPS/Register/register[0][3] ), .QN(n945)
         );
  DFFRX1 \i_MIPS/Register/register_reg[0][4]  ( .D(\i_MIPS/Register/n1112 ), 
        .CK(clk), .RN(n6225), .Q(\i_MIPS/Register/register[0][4] ), .QN(n944)
         );
  DFFRX1 \i_MIPS/Register/register_reg[0][5]  ( .D(\i_MIPS/Register/n1113 ), 
        .CK(clk), .RN(n6225), .Q(\i_MIPS/Register/register[0][5] ), .QN(n943)
         );
  DFFRX1 \i_MIPS/Register/register_reg[0][6]  ( .D(\i_MIPS/Register/n1114 ), 
        .CK(clk), .RN(n6225), .Q(\i_MIPS/Register/register[0][6] ), .QN(n2550)
         );
  DFFRX1 \i_MIPS/Register/register_reg[0][7]  ( .D(\i_MIPS/Register/n1115 ), 
        .CK(clk), .RN(n6225), .Q(\i_MIPS/Register/register[0][7] ), .QN(n2569)
         );
  DFFRX1 \i_MIPS/Register/register_reg[0][8]  ( .D(\i_MIPS/Register/n1116 ), 
        .CK(clk), .RN(n6225), .Q(\i_MIPS/Register/register[0][8] ), .QN(n2538)
         );
  DFFRX1 \i_MIPS/Register/register_reg[0][9]  ( .D(\i_MIPS/Register/n1117 ), 
        .CK(clk), .RN(n6225), .Q(\i_MIPS/Register/register[0][9] ), .QN(n2342)
         );
  DFFRX1 \i_MIPS/Register/register_reg[0][10]  ( .D(\i_MIPS/Register/n1118 ), 
        .CK(clk), .RN(n6225), .Q(\i_MIPS/Register/register[0][10] ), .QN(n2343) );
  DFFRX1 \i_MIPS/Register/register_reg[0][11]  ( .D(\i_MIPS/Register/n1119 ), 
        .CK(clk), .RN(n6225), .Q(\i_MIPS/Register/register[0][11] ), .QN(n2361) );
  DFFRX1 \i_MIPS/Register/register_reg[0][12]  ( .D(\i_MIPS/Register/n1120 ), 
        .CK(clk), .RN(n6225), .Q(\i_MIPS/Register/register[0][12] ), .QN(n2542) );
  DFFRX1 \i_MIPS/Register/register_reg[0][13]  ( .D(\i_MIPS/Register/n1121 ), 
        .CK(clk), .RN(n6225), .Q(\i_MIPS/Register/register[0][13] ), .QN(n2544) );
  DFFRX1 \i_MIPS/Register/register_reg[0][15]  ( .D(\i_MIPS/Register/n1123 ), 
        .CK(clk), .RN(n6225), .Q(\i_MIPS/Register/register[0][15] ), .QN(n324)
         );
  DFFRX1 \i_MIPS/Register/register_reg[0][16]  ( .D(\i_MIPS/Register/n1124 ), 
        .CK(clk), .RN(n6224), .Q(\i_MIPS/Register/register[0][16] ), .QN(n2532) );
  DFFRX1 \i_MIPS/Register/register_reg[0][17]  ( .D(\i_MIPS/Register/n1125 ), 
        .CK(clk), .RN(n6224), .Q(\i_MIPS/Register/register[0][17] ), .QN(n912)
         );
  DFFRX1 \i_MIPS/Register/register_reg[0][18]  ( .D(\i_MIPS/Register/n1126 ), 
        .CK(clk), .RN(n6224), .Q(\i_MIPS/Register/register[0][18] ), .QN(n2363) );
  DFFRX1 \i_MIPS/Register/register_reg[0][19]  ( .D(\i_MIPS/Register/n1127 ), 
        .CK(clk), .RN(n6224), .Q(\i_MIPS/Register/register[0][19] ), .QN(n2454) );
  DFFRX1 \i_MIPS/Register/register_reg[0][20]  ( .D(\i_MIPS/Register/n1128 ), 
        .CK(clk), .RN(n6224), .Q(\i_MIPS/Register/register[0][20] ), .QN(n2169) );
  DFFRX1 \i_MIPS/Register/register_reg[0][21]  ( .D(\i_MIPS/Register/n1129 ), 
        .CK(clk), .RN(n6224), .Q(\i_MIPS/Register/register[0][21] ), .QN(n2171) );
  DFFRX1 \i_MIPS/Register/register_reg[0][23]  ( .D(\i_MIPS/Register/n1131 ), 
        .CK(clk), .RN(n6224), .Q(\i_MIPS/Register/register[0][23] ), .QN(n317)
         );
  DFFRX1 \i_MIPS/Register/register_reg[0][24]  ( .D(\i_MIPS/Register/n1132 ), 
        .CK(clk), .RN(n6224), .Q(\i_MIPS/Register/register[0][24] ), .QN(n333)
         );
  DFFRX1 \i_MIPS/Register/register_reg[0][25]  ( .D(\i_MIPS/Register/n1133 ), 
        .CK(clk), .RN(n6224), .Q(\i_MIPS/Register/register[0][25] ), .QN(n334)
         );
  DFFRX1 \i_MIPS/Register/register_reg[0][26]  ( .D(\i_MIPS/Register/n1134 ), 
        .CK(clk), .RN(n6224), .Q(\i_MIPS/Register/register[0][26] ), .QN(n2537) );
  DFFRX1 \i_MIPS/Register/register_reg[0][27]  ( .D(\i_MIPS/Register/n1135 ), 
        .CK(clk), .RN(n6224), .Q(\i_MIPS/Register/register[0][27] ), .QN(n2545) );
  DFFRX1 \i_MIPS/Register/register_reg[0][28]  ( .D(\i_MIPS/Register/n1136 ), 
        .CK(clk), .RN(n6223), .Q(\i_MIPS/Register/register[0][28] ), .QN(n2562) );
  DFFRX1 \i_MIPS/Register/register_reg[0][29]  ( .D(\i_MIPS/Register/n1137 ), 
        .CK(clk), .RN(n6223), .Q(\i_MIPS/Register/register[0][29] ), .QN(n319)
         );
  DFFRX1 \i_MIPS/Register/register_reg[31][22]  ( .D(n11550), .CK(clk), .RN(
        n6307), .Q(\i_MIPS/Register/register[31][22] ), .QN(n3546) );
  DFFRX1 \i_MIPS/IF_ID_reg[17]  ( .D(\i_MIPS/N34 ), .CK(clk), .RN(n6331), .Q(
        \i_MIPS/IF_ID[17] ), .QN(\i_MIPS/n170 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[22]  ( .D(\i_MIPS/N39 ), .CK(clk), .RN(n6332), .Q(
        \i_MIPS/IF_ID[22] ), .QN(\i_MIPS/n175 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[21]  ( .D(\i_MIPS/N38 ), .CK(clk), .RN(n6331), .Q(
        \i_MIPS/IF_ID[21] ), .QN(\i_MIPS/n174 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[19]  ( .D(\i_MIPS/N36 ), .CK(clk), .RN(n6331), .Q(
        \i_MIPS/IF_ID[19] ), .QN(\i_MIPS/n172 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[18]  ( .D(\i_MIPS/N35 ), .CK(clk), .RN(n6331), .Q(
        \i_MIPS/IF_ID[18] ), .QN(\i_MIPS/n171 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[12]  ( .D(\i_MIPS/N29 ), .CK(clk), .RN(n6331), .Q(
        \i_MIPS/IF_ID[12] ), .QN(\i_MIPS/n165 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[13]  ( .D(\i_MIPS/N30 ), .CK(clk), .RN(n6331), .Q(
        \i_MIPS/IF_ID[13] ), .QN(\i_MIPS/n166 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[15]  ( .D(\i_MIPS/N32 ), .CK(clk), .RN(n6331), .Q(
        \i_MIPS/IF_ID[15] ), .QN(\i_MIPS/n168 ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][0]  ( .D(\i_MIPS/Register/n532 ), 
        .CK(clk), .RN(n6274), .Q(\i_MIPS/Register/register[18][0] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][1]  ( .D(\i_MIPS/Register/n533 ), 
        .CK(clk), .RN(n6274), .Q(\i_MIPS/Register/register[18][1] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][3]  ( .D(\i_MIPS/Register/n535 ), 
        .CK(clk), .RN(n6274), .Q(\i_MIPS/Register/register[18][3] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][4]  ( .D(\i_MIPS/Register/n536 ), 
        .CK(clk), .RN(n6273), .Q(\i_MIPS/Register/register[18][4] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][5]  ( .D(\i_MIPS/Register/n537 ), 
        .CK(clk), .RN(n6273), .Q(\i_MIPS/Register/register[18][5] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][8]  ( .D(\i_MIPS/Register/n540 ), 
        .CK(clk), .RN(n6273), .Q(\i_MIPS/Register/register[18][8] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][10]  ( .D(\i_MIPS/Register/n542 ), 
        .CK(clk), .RN(n6273), .Q(\i_MIPS/Register/register[18][10] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][11]  ( .D(\i_MIPS/Register/n543 ), 
        .CK(clk), .RN(n6273), .Q(\i_MIPS/Register/register[18][11] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][12]  ( .D(\i_MIPS/Register/n544 ), 
        .CK(clk), .RN(n6273), .Q(\i_MIPS/Register/register[18][12] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][16]  ( .D(\i_MIPS/Register/n548 ), 
        .CK(clk), .RN(n6272), .Q(\i_MIPS/Register/register[18][16] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][17]  ( .D(\i_MIPS/Register/n549 ), 
        .CK(clk), .RN(n6272), .Q(\i_MIPS/Register/register[18][17] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][18]  ( .D(\i_MIPS/Register/n550 ), 
        .CK(clk), .RN(n6272), .Q(\i_MIPS/Register/register[18][18] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][19]  ( .D(\i_MIPS/Register/n551 ), 
        .CK(clk), .RN(n6272), .Q(\i_MIPS/Register/register[18][19] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][20]  ( .D(\i_MIPS/Register/n552 ), 
        .CK(clk), .RN(n6272), .Q(\i_MIPS/Register/register[18][20] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][21]  ( .D(\i_MIPS/Register/n553 ), 
        .CK(clk), .RN(n6272), .Q(\i_MIPS/Register/register[18][21] ) );
  DFFRX1 \i_MIPS/Register/register_reg[18][27]  ( .D(\i_MIPS/Register/n559 ), 
        .CK(clk), .RN(n6272), .Q(\i_MIPS/Register/register[18][27] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][0]  ( .D(\i_MIPS/Register/n1044 ), 
        .CK(clk), .RN(n6231), .Q(\i_MIPS/Register/register[2][0] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][1]  ( .D(\i_MIPS/Register/n1045 ), 
        .CK(clk), .RN(n6231), .Q(\i_MIPS/Register/register[2][1] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][3]  ( .D(\i_MIPS/Register/n1047 ), 
        .CK(clk), .RN(n6231), .Q(\i_MIPS/Register/register[2][3] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][4]  ( .D(\i_MIPS/Register/n1048 ), 
        .CK(clk), .RN(n6231), .Q(\i_MIPS/Register/register[2][4] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][5]  ( .D(\i_MIPS/Register/n1049 ), 
        .CK(clk), .RN(n6231), .Q(\i_MIPS/Register/register[2][5] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][8]  ( .D(\i_MIPS/Register/n1052 ), 
        .CK(clk), .RN(n6230), .Q(\i_MIPS/Register/register[2][8] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][11]  ( .D(\i_MIPS/Register/n1055 ), 
        .CK(clk), .RN(n6230), .Q(\i_MIPS/Register/register[2][11] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][12]  ( .D(\i_MIPS/Register/n1056 ), 
        .CK(clk), .RN(n6230), .Q(\i_MIPS/Register/register[2][12] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][16]  ( .D(\i_MIPS/Register/n1060 ), 
        .CK(clk), .RN(n6230), .Q(\i_MIPS/Register/register[2][16] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][17]  ( .D(\i_MIPS/Register/n1061 ), 
        .CK(clk), .RN(n6230), .Q(\i_MIPS/Register/register[2][17] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][18]  ( .D(\i_MIPS/Register/n1062 ), 
        .CK(clk), .RN(n6230), .Q(\i_MIPS/Register/register[2][18] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][19]  ( .D(\i_MIPS/Register/n1063 ), 
        .CK(clk), .RN(n6230), .Q(\i_MIPS/Register/register[2][19] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][20]  ( .D(\i_MIPS/Register/n1064 ), 
        .CK(clk), .RN(n6229), .Q(\i_MIPS/Register/register[2][20] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][21]  ( .D(\i_MIPS/Register/n1065 ), 
        .CK(clk), .RN(n6229), .Q(\i_MIPS/Register/register[2][21] ) );
  DFFRX1 \i_MIPS/Register/register_reg[2][27]  ( .D(\i_MIPS/Register/n1071 ), 
        .CK(clk), .RN(n6229), .Q(\i_MIPS/Register/register[2][27] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][0]  ( .D(\i_MIPS/Register/n276 ), 
        .CK(clk), .RN(n6295), .Q(\i_MIPS/Register/register[26][0] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][1]  ( .D(\i_MIPS/Register/n277 ), 
        .CK(clk), .RN(n6295), .Q(\i_MIPS/Register/register[26][1] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][3]  ( .D(\i_MIPS/Register/n279 ), 
        .CK(clk), .RN(n6295), .Q(\i_MIPS/Register/register[26][3] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][4]  ( .D(\i_MIPS/Register/n280 ), 
        .CK(clk), .RN(n6295), .Q(\i_MIPS/Register/register[26][4] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][5]  ( .D(\i_MIPS/Register/n281 ), 
        .CK(clk), .RN(n6295), .Q(\i_MIPS/Register/register[26][5] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][7]  ( .D(\i_MIPS/Register/n283 ), 
        .CK(clk), .RN(n6295), .Q(\i_MIPS/Register/register[26][7] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][8]  ( .D(\i_MIPS/Register/n284 ), 
        .CK(clk), .RN(n6294), .Q(\i_MIPS/Register/register[26][8] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][10]  ( .D(\i_MIPS/Register/n286 ), 
        .CK(clk), .RN(n6294), .Q(\i_MIPS/Register/register[26][10] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][11]  ( .D(\i_MIPS/Register/n287 ), 
        .CK(clk), .RN(n6294), .Q(\i_MIPS/Register/register[26][11] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][12]  ( .D(\i_MIPS/Register/n288 ), 
        .CK(clk), .RN(n6294), .Q(\i_MIPS/Register/register[26][12] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][16]  ( .D(\i_MIPS/Register/n292 ), 
        .CK(clk), .RN(n6294), .Q(\i_MIPS/Register/register[26][16] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][17]  ( .D(\i_MIPS/Register/n293 ), 
        .CK(clk), .RN(n6294), .Q(\i_MIPS/Register/register[26][17] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][18]  ( .D(\i_MIPS/Register/n294 ), 
        .CK(clk), .RN(n6294), .Q(\i_MIPS/Register/register[26][18] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][19]  ( .D(\i_MIPS/Register/n295 ), 
        .CK(clk), .RN(n6294), .Q(\i_MIPS/Register/register[26][19] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][20]  ( .D(\i_MIPS/Register/n296 ), 
        .CK(clk), .RN(n6293), .Q(\i_MIPS/Register/register[26][20] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][21]  ( .D(\i_MIPS/Register/n297 ), 
        .CK(clk), .RN(n6293), .Q(\i_MIPS/Register/register[26][21] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][26]  ( .D(\i_MIPS/Register/n302 ), 
        .CK(clk), .RN(n6293), .Q(\i_MIPS/Register/register[26][26] ) );
  DFFRX1 \i_MIPS/Register/register_reg[26][27]  ( .D(\i_MIPS/Register/n303 ), 
        .CK(clk), .RN(n6293), .Q(\i_MIPS/Register/register[26][27] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][0]  ( .D(\i_MIPS/Register/n788 ), 
        .CK(clk), .RN(n6252), .Q(\i_MIPS/Register/register[10][0] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][1]  ( .D(\i_MIPS/Register/n789 ), 
        .CK(clk), .RN(n6252), .Q(\i_MIPS/Register/register[10][1] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][3]  ( .D(\i_MIPS/Register/n791 ), 
        .CK(clk), .RN(n6252), .Q(\i_MIPS/Register/register[10][3] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][4]  ( .D(\i_MIPS/Register/n792 ), 
        .CK(clk), .RN(n6252), .Q(\i_MIPS/Register/register[10][4] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][5]  ( .D(\i_MIPS/Register/n793 ), 
        .CK(clk), .RN(n6252), .Q(\i_MIPS/Register/register[10][5] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][8]  ( .D(\i_MIPS/Register/n796 ), 
        .CK(clk), .RN(n6252), .Q(\i_MIPS/Register/register[10][8] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][10]  ( .D(\i_MIPS/Register/n798 ), 
        .CK(clk), .RN(n6252), .Q(\i_MIPS/Register/register[10][10] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][11]  ( .D(\i_MIPS/Register/n799 ), 
        .CK(clk), .RN(n6252), .Q(\i_MIPS/Register/register[10][11] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][12]  ( .D(\i_MIPS/Register/n800 ), 
        .CK(clk), .RN(n6251), .Q(\i_MIPS/Register/register[10][12] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][16]  ( .D(\i_MIPS/Register/n804 ), 
        .CK(clk), .RN(n6251), .Q(\i_MIPS/Register/register[10][16] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][17]  ( .D(\i_MIPS/Register/n805 ), 
        .CK(clk), .RN(n6251), .Q(\i_MIPS/Register/register[10][17] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][18]  ( .D(\i_MIPS/Register/n806 ), 
        .CK(clk), .RN(n6251), .Q(\i_MIPS/Register/register[10][18] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][19]  ( .D(\i_MIPS/Register/n807 ), 
        .CK(clk), .RN(n6251), .Q(\i_MIPS/Register/register[10][19] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][20]  ( .D(\i_MIPS/Register/n808 ), 
        .CK(clk), .RN(n6251), .Q(\i_MIPS/Register/register[10][20] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][21]  ( .D(\i_MIPS/Register/n809 ), 
        .CK(clk), .RN(n6251), .Q(\i_MIPS/Register/register[10][21] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][26]  ( .D(\i_MIPS/Register/n814 ), 
        .CK(clk), .RN(n6250), .Q(\i_MIPS/Register/register[10][26] ) );
  DFFRX1 \i_MIPS/Register/register_reg[10][27]  ( .D(\i_MIPS/Register/n815 ), 
        .CK(clk), .RN(n6250), .Q(\i_MIPS/Register/register[10][27] ) );
  DFFRX1 \i_MIPS/IF_ID_reg[14]  ( .D(\i_MIPS/N31 ), .CK(clk), .RN(n6331), .Q(
        \i_MIPS/IF_ID[14] ), .QN(\i_MIPS/n167 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[0]  ( .D(\i_MIPS/n493 ), .CK(clk), .RN(n6311), .Q(
        \i_MIPS/EX_MEM_0 ), .QN(\i_MIPS/n303 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[16]  ( .D(\i_MIPS/N33 ), .CK(clk), .RN(n6331), .Q(
        \i_MIPS/IF_ID[16] ), .QN(\i_MIPS/n169 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[20]  ( .D(\i_MIPS/N37 ), .CK(clk), .RN(n6331), .Q(
        \i_MIPS/IF_ID[20] ), .QN(\i_MIPS/n173 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[36]  ( .D(\i_MIPS/n368 ), .CK(clk), .RN(n6324), 
        .Q(n12954), .QN(n4983) );
  DFFRX1 \i_MIPS/EX_MEM_reg[23]  ( .D(\i_MIPS/n381 ), .CK(clk), .RN(n6323), 
        .Q(n12967), .QN(n1941) );
  DFFRX1 \i_MIPS/EX_MEM_reg[28]  ( .D(\i_MIPS/n376 ), .CK(clk), .RN(n6324), 
        .Q(n12962), .QN(n2013) );
  DFFRX1 \i_MIPS/EX_MEM_reg[14]  ( .D(\i_MIPS/n390 ), .CK(clk), .RN(n6322), 
        .Q(n12976), .QN(n4371) );
  DFFRX1 \i_MIPS/EX_MEM_reg[13]  ( .D(\i_MIPS/n391 ), .CK(clk), .RN(n6322), 
        .Q(n12977) );
  DFFRX1 \i_MIPS/EX_MEM_reg[15]  ( .D(\i_MIPS/n389 ), .CK(clk), .RN(n6323), 
        .Q(n12975), .QN(n4002) );
  DFFRX1 \i_MIPS/EX_MEM_reg[22]  ( .D(\i_MIPS/n382 ), .CK(clk), .RN(n6323), 
        .Q(n12968), .QN(n2998) );
  DFFRX1 \i_MIPS/EX_MEM_reg[18]  ( .D(\i_MIPS/n386 ), .CK(clk), .RN(n6323), 
        .Q(n12972), .QN(n3019) );
  DFFRX1 \i_MIPS/EX_MEM_reg[25]  ( .D(\i_MIPS/n379 ), .CK(clk), .RN(n6323), 
        .Q(n12965) );
  DFFRX1 \i_MIPS/EX_MEM_reg[26]  ( .D(\i_MIPS/n378 ), .CK(clk), .RN(n6323), 
        .Q(n12964), .QN(n4365) );
  DFFRX1 \i_MIPS/EX_MEM_reg[30]  ( .D(\i_MIPS/n374 ), .CK(clk), .RN(n6324), 
        .Q(n12960), .QN(n2997) );
  DFFRX1 \i_MIPS/EX_MEM_reg[32]  ( .D(\i_MIPS/n372 ), .CK(clk), .RN(n6324), 
        .Q(n12958), .QN(n3018) );
  DFFRX1 \i_MIPS/PC/PC_o_reg[30]  ( .D(\i_MIPS/PC/n64 ), .CK(clk), .RN(n6309), 
        .Q(ICACHE_addr[28]), .QN(\i_MIPS/PC/n32 ) );
  DFFRX2 \i_MIPS/EX_MEM_reg[1]  ( .D(\i_MIPS/n456 ), .CK(clk), .RN(n6314), .Q(
        \i_MIPS/EX_MEM_1 ), .QN(\i_MIPS/n266 ) );
  DFFRX2 \i_MIPS/EX_MEM_reg[3]  ( .D(\i_MIPS/n454 ), .CK(clk), .RN(n6315), .Q(
        DCACHE_ren), .QN(\i_MIPS/n264 ) );
  DFFRX2 \i_MIPS/EX_MEM_reg[72]  ( .D(\i_MIPS/n404 ), .CK(clk), .RN(n6321), 
        .Q(\i_MIPS/Reg_W[3] ), .QN(n1931) );
  DFFRX2 \i_MIPS/EX_MEM_reg[73]  ( .D(\i_MIPS/n403 ), .CK(clk), .RN(n6321), 
        .Q(\i_MIPS/Reg_W[4] ), .QN(n1932) );
  DFFRX1 \i_MIPS/EX_MEM_reg[29]  ( .D(\i_MIPS/n375 ), .CK(clk), .RN(n6324), 
        .Q(n12961), .QN(n5024) );
  DFFRX1 \i_MIPS/EX_MEM_reg[31]  ( .D(\i_MIPS/n373 ), .CK(clk), .RN(n6324), 
        .Q(n12959), .QN(n5021) );
  DFFRX1 \i_MIPS/EX_MEM_reg[34]  ( .D(\i_MIPS/n370 ), .CK(clk), .RN(n6324), 
        .Q(n12956), .QN(n5008) );
  DFFRX1 \i_MIPS/EX_MEM_reg[24]  ( .D(\i_MIPS/n380 ), .CK(clk), .RN(n6323), 
        .Q(n12966), .QN(n4920) );
  DFFRX1 \I_cache/cache_reg[2][142]  ( .D(n11707), .CK(clk), .RN(n6025), .Q(
        \I_cache/cache[2][142] ), .QN(n2933) );
  DFFRX1 \I_cache/cache_reg[3][142]  ( .D(n11706), .CK(clk), .RN(n6025), .Q(
        \I_cache/cache[3][142] ), .QN(n1296) );
  DFFRX1 \I_cache/cache_reg[6][142]  ( .D(n11703), .CK(clk), .RN(n6025), .Q(
        \I_cache/cache[6][142] ), .QN(n1297) );
  DFFRX1 \I_cache/cache_reg[1][145]  ( .D(n11684), .CK(clk), .RN(n6023), .Q(
        \I_cache/cache[1][145] ), .QN(n1288) );
  DFFRX1 \I_cache/cache_reg[2][145]  ( .D(n11683), .CK(clk), .RN(n6023), .Q(
        \I_cache/cache[2][145] ), .QN(n2973) );
  DFFRX1 \I_cache/cache_reg[5][145]  ( .D(n11680), .CK(clk), .RN(n6023), .Q(
        \I_cache/cache[5][145] ) );
  DFFRX1 \I_cache/cache_reg[6][145]  ( .D(n11679), .CK(clk), .RN(n6023), .Q(
        \I_cache/cache[6][145] ), .QN(n1301) );
  DFFRX1 \I_cache/cache_reg[1][151]  ( .D(n11636), .CK(clk), .RN(n6019), .Q(
        \I_cache/cache[1][151] ), .QN(n2931) );
  DFFRX1 \I_cache/cache_reg[3][151]  ( .D(n11634), .CK(clk), .RN(n6019), .Q(
        \I_cache/cache[3][151] ), .QN(n1294) );
  DFFRX1 \I_cache/cache_reg[6][151]  ( .D(n11631), .CK(clk), .RN(n6019), .Q(
        \I_cache/cache[6][151] ), .QN(n1300) );
  DFFRX1 \I_cache/cache_reg[7][128]  ( .D(n11814), .CK(clk), .RN(n6017), .Q(
        \I_cache/cache[7][128] ), .QN(n2965) );
  DFFRX1 \i_MIPS/PC/PC_o_reg[25]  ( .D(\i_MIPS/PC/n59 ), .CK(clk), .RN(n6309), 
        .Q(ICACHE_addr[23]), .QN(\i_MIPS/PC/n27 ) );
  DFFRX1 \I_cache/cache_reg[7][134]  ( .D(n11766), .CK(clk), .RN(n6030), .Q(
        \I_cache/cache[7][134] ), .QN(n2219) );
  DFFRX1 \I_cache/cache_reg[7][138]  ( .D(n11734), .CK(clk), .RN(n6027), .Q(
        \I_cache/cache[7][138] ), .QN(n493) );
  DFFRX1 \I_cache/cache_reg[7][142]  ( .D(n11702), .CK(clk), .RN(n6025), .Q(
        \I_cache/cache[7][142] ), .QN(n2963) );
  DFFRX1 \I_cache/cache_reg[1][138]  ( .D(n11740), .CK(clk), .RN(n6028), .Q(
        \I_cache/cache[1][138] ), .QN(n2008) );
  DFFRX1 \I_cache/cache_reg[6][138]  ( .D(n11735), .CK(clk), .RN(n6027), .Q(
        \I_cache/cache[6][138] ), .QN(n2969) );
  DFFRX1 \I_cache/cache_reg[3][138]  ( .D(n11738), .CK(clk), .RN(n6028), .Q(
        \I_cache/cache[3][138] ), .QN(n2929) );
  DFFRX1 \I_cache/cache_reg[4][141]  ( .D(n11713), .CK(clk), .RN(n6026), .Q(
        \I_cache/cache[4][141] ), .QN(n4679) );
  DFFRX1 \I_cache/cache_reg[3][145]  ( .D(n11682), .CK(clk), .RN(n6023), .Q(
        \I_cache/cache[3][145] ), .QN(n1295) );
  DFFRX1 \I_cache/cache_reg[3][146]  ( .D(n11674), .CK(clk), .RN(n6022), .Q(
        \I_cache/cache[3][146] ), .QN(n1290) );
  DFFRX1 \I_cache/cache_reg[4][146]  ( .D(n11673), .CK(clk), .RN(n6022), .Q(
        \I_cache/cache[4][146] ), .QN(n2927) );
  DFFRX1 \I_cache/cache_reg[7][146]  ( .D(n11670), .CK(clk), .RN(n6022), .Q(
        \I_cache/cache[7][146] ), .QN(n1291) );
  DFFRX1 \I_cache/cache_reg[1][150]  ( .D(n11644), .CK(clk), .RN(n6020), .Q(
        \I_cache/cache[1][150] ), .QN(n1289) );
  DFFRX1 \I_cache/cache_reg[3][150]  ( .D(n11642), .CK(clk), .RN(n6020), .Q(
        \I_cache/cache[3][150] ), .QN(n1292) );
  DFFRX1 \I_cache/cache_reg[4][150]  ( .D(n11641), .CK(clk), .RN(n6020), .Q(
        \I_cache/cache[4][150] ), .QN(n2926) );
  DFFRX1 \I_cache/cache_reg[6][150]  ( .D(n11639), .CK(clk), .RN(n6019), .Q(
        \I_cache/cache[6][150] ), .QN(n2932) );
  DFFRX1 \I_cache/cache_reg[7][150]  ( .D(n11638), .CK(clk), .RN(n6019), .Q(
        \I_cache/cache[7][150] ), .QN(n1293) );
  DFFRX1 \I_cache/cache_reg[0][152]  ( .D(n11629), .CK(clk), .RN(n6019), .Q(
        \I_cache/cache[0][152] ), .QN(n1298) );
  DFFRX1 \I_cache/cache_reg[2][152]  ( .D(n11627), .CK(clk), .RN(n6018), .Q(
        \I_cache/cache[2][152] ), .QN(n1299) );
  DFFRX1 \I_cache/cache_reg[4][152]  ( .D(n11625), .CK(clk), .RN(n6018), .Q(
        \I_cache/cache[4][152] ), .QN(n2925) );
  DFFRX1 \I_cache/cache_reg[7][145]  ( .D(n11678), .CK(clk), .RN(n6023), .Q(
        \I_cache/cache[7][145] ), .QN(n2967) );
  DFFRX1 \I_cache/cache_reg[7][151]  ( .D(n11630), .CK(clk), .RN(n6019), .Q(
        \I_cache/cache[7][151] ), .QN(n2966) );
  DFFRX1 \I_cache/cache_reg[0][146]  ( .D(n11677), .CK(clk), .RN(n6023), .Q(
        \I_cache/cache[0][146] ), .QN(n1310) );
  DFFRX1 \I_cache/cache_reg[2][146]  ( .D(n11675), .CK(clk), .RN(n6022), .Q(
        \I_cache/cache[2][146] ), .QN(n2941) );
  DFFRX1 \I_cache/cache_reg[6][146]  ( .D(n11671), .CK(clk), .RN(n6022), .Q(
        \I_cache/cache[6][146] ), .QN(n2942) );
  DFFRX1 \I_cache/cache_reg[0][150]  ( .D(n11645), .CK(clk), .RN(n6020), .Q(
        \I_cache/cache[0][150] ), .QN(n2940) );
  DFFRX1 \I_cache/cache_reg[2][150]  ( .D(n11643), .CK(clk), .RN(n6020), .Q(
        \I_cache/cache[2][150] ), .QN(n2943) );
  DFFRX1 \I_cache/cache_reg[1][146]  ( .D(n11676), .CK(clk), .RN(n6022), .Q(
        \I_cache/cache[1][146] ), .QN(n2962) );
  DFFRX1 \I_cache/cache_reg[5][146]  ( .D(n11672), .CK(clk), .RN(n6022), .Q(
        \I_cache/cache[5][146] ) );
  DFFRX1 \I_cache/cache_reg[5][150]  ( .D(n11640), .CK(clk), .RN(n6019), .Q(
        \I_cache/cache[5][150] ) );
  DFFRX1 \I_cache/cache_reg[3][132]  ( .D(n11786), .CK(clk), .RN(n6032), .Q(
        \I_cache/cache[3][132] ), .QN(n497) );
  DFFRX1 \I_cache/cache_reg[1][142]  ( .D(n11708), .CK(clk), .RN(n6025), .Q(
        \I_cache/cache[1][142] ), .QN(n2930) );
  DFFRX1 \I_cache/cache_reg[7][132]  ( .D(n11782), .CK(clk), .RN(n6031), .Q(
        \I_cache/cache[7][132] ), .QN(n2982) );
  DFFRX1 \i_MIPS/EX_MEM_reg[8]  ( .D(\i_MIPS/n396 ), .CK(clk), .RN(n6322), .Q(
        n12980), .QN(n1319) );
  DFFRX1 \i_MIPS/EX_MEM_reg[7]  ( .D(\i_MIPS/n397 ), .CK(clk), .RN(n6322), .Q(
        n12981), .QN(n3003) );
  DFFRHQX8 \i_MIPS/ID_EX_reg[8]  ( .D(\i_MIPS/n400 ), .CK(clk), .RN(n6322), 
        .Q(net143503) );
  DFFRX4 \i_MIPS/ID_EX_reg[12]  ( .D(\i_MIPS/n489 ), .CK(clk), .RN(n6312), .Q(
        \i_MIPS/ALUin1[3] ), .QN(n2928) );
  DFFRX4 \i_MIPS/ID_EX_reg[13]  ( .D(\i_MIPS/n488 ), .CK(clk), .RN(n6312), .Q(
        \i_MIPS/ALUin1[4] ), .QN(\i_MIPS/n297 ) );
  DFFRX4 \i_MIPS/ID_EX_reg[9]  ( .D(\i_MIPS/n492 ), .CK(clk), .RN(n6311), .Q(
        \i_MIPS/ALUin1[0] ), .QN(\i_MIPS/n301 ) );
  DFFRX4 \i_MIPS/PC/PC_o_reg[3]  ( .D(\i_MIPS/PC/n37 ), .CK(clk), .RN(n6311), 
        .Q(ICACHE_addr[1]), .QN(\i_MIPS/PC/n5 ) );
  DFFRX4 \i_MIPS/PC/PC_o_reg[22]  ( .D(\i_MIPS/PC/n56 ), .CK(clk), .RN(n6309), 
        .Q(ICACHE_addr[20]), .QN(\i_MIPS/PC/n24 ) );
  DFFRX4 \i_MIPS/PC/PC_o_reg[26]  ( .D(\i_MIPS/PC/n60 ), .CK(clk), .RN(n6309), 
        .Q(ICACHE_addr[24]), .QN(\i_MIPS/PC/n28 ) );
  DFFRX4 \i_MIPS/PC/PC_o_reg[24]  ( .D(\i_MIPS/PC/n58 ), .CK(clk), .RN(n6309), 
        .Q(ICACHE_addr[22]), .QN(\i_MIPS/PC/n26 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[46]  ( .D(\i_MIPS/n357 ), .CK(clk), .RN(n6325), .Q(
        n3548), .QN(\i_MIPS/n234 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[62]  ( .D(\i_MIPS/n325 ), .CK(clk), .RN(n6328), 
        .QN(\i_MIPS/n202 ) );
  DFFRX4 \i_MIPS/ID_EX_reg[16]  ( .D(\i_MIPS/n485 ), .CK(clk), .RN(n6312), .Q(
        \i_MIPS/ALUin1[7] ), .QN(n2892) );
  DFFRX4 \i_MIPS/ID_EX_reg[107]  ( .D(\i_MIPS/n413 ), .CK(clk), .RN(n6320), 
        .Q(\i_MIPS/ID_EX[107] ), .QN(\i_MIPS/n252 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[56]  ( .D(\i_MIPS/n337 ), .CK(clk), .RN(n6327), .Q(
        n3550), .QN(\i_MIPS/n214 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[58]  ( .D(\i_MIPS/n333 ), .CK(clk), .RN(n6327), .Q(
        n3545), .QN(\i_MIPS/n210 ) );
  DFFRX4 \i_MIPS/ID_EX_reg[11]  ( .D(\i_MIPS/n490 ), .CK(clk), .RN(n6311), .Q(
        \i_MIPS/ALUin1[2] ), .QN(\i_MIPS/n299 ) );
  DFFRX4 \i_MIPS/PC/PC_o_reg[2]  ( .D(\i_MIPS/PC/n36 ), .CK(clk), .RN(n6311), 
        .Q(ICACHE_addr[0]), .QN(\i_MIPS/PC/n4 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[57]  ( .D(\i_MIPS/n335 ), .CK(clk), .RN(n6327), .Q(
        n3549), .QN(\i_MIPS/n212 ) );
  DFFRX4 \i_MIPS/ID_EX_reg[55]  ( .D(\i_MIPS/n339 ), .CK(clk), .RN(n6327), .Q(
        n3747), .QN(\i_MIPS/n216 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[54]  ( .D(\i_MIPS/n341 ), .CK(clk), .RN(n6327), .Q(
        n3543), .QN(\i_MIPS/n218 ) );
  DFFRX4 \i_MIPS/ID_EX_reg[35]  ( .D(\i_MIPS/n466 ), .CK(clk), .RN(n6313), .Q(
        \i_MIPS/ALUin1[26] ), .QN(n253) );
  DFFRX4 \i_MIPS/ID_EX_reg[23]  ( .D(\i_MIPS/n478 ), .CK(clk), .RN(n6312), .Q(
        \i_MIPS/ALUin1[14] ), .QN(\i_MIPS/n287 ) );
  DFFRX4 \i_MIPS/ID_EX_reg[19]  ( .D(\i_MIPS/n482 ), .CK(clk), .RN(n6312), .Q(
        \i_MIPS/ALUin1[10] ), .QN(n300) );
  DFFRX4 \i_MIPS/ID_EX_reg[37]  ( .D(\i_MIPS/n464 ), .CK(clk), .RN(n6314), .Q(
        \i_MIPS/ALUin1[28] ), .QN(n347) );
  DFFRX4 \i_MIPS/ID_EX_reg[24]  ( .D(\i_MIPS/n477 ), .CK(clk), .RN(n6313), .Q(
        \i_MIPS/ALUin1[15] ), .QN(n3670) );
  DFFRX4 \i_MIPS/ID_EX_reg[29]  ( .D(\i_MIPS/n472 ), .CK(clk), .RN(n6313), .Q(
        \i_MIPS/ALUin1[20] ), .QN(n2919) );
  DFFRX2 \i_MIPS/ID_EX_reg[111]  ( .D(\i_MIPS/n449 ), .CK(clk), .RN(n6316), 
        .Q(\i_MIPS/ID_EX[111] ), .QN(\i_MIPS/n259 ) );
  DFFRX4 \i_MIPS/IF_ID_reg[38]  ( .D(\i_MIPS/N55 ), .CK(clk), .RN(n6317), .Q(
        n2948), .QN(\i_MIPS/n515 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[114]  ( .D(\i_MIPS/n452 ), .CK(clk), .RN(n6315), 
        .Q(\i_MIPS/ID_EX[114] ), .QN(\i_MIPS/n262 ) );
  DFFRX4 \i_MIPS/ID_EX_reg[115]  ( .D(\i_MIPS/n453 ), .CK(clk), .RN(n6315), 
        .Q(\i_MIPS/ID_EX[115] ), .QN(\i_MIPS/n263 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[103]  ( .D(\i_MIPS/n418 ), .CK(clk), .RN(n6320), 
        .Q(\i_MIPS/ID_EX[103] ) );
  DFFRX2 \i_MIPS/ID_EX_reg[53]  ( .D(\i_MIPS/n343 ), .CK(clk), .RN(n6326), .Q(
        n3551), .QN(\i_MIPS/n220 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[58]  ( .D(\i_MIPS/N75 ), .CK(clk), .RN(n6321), .Q(
        \i_MIPS/IR[26] ), .QN(\i_MIPS/n247 ) );
  DFFRX4 \i_MIPS/IF_ID_reg[33]  ( .D(\i_MIPS/N50 ), .CK(clk), .RN(n6317), .Q(
        \i_MIPS/Sign_Extend[1] ), .QN(\i_MIPS/n520 ) );
  DFFRX4 \i_MIPS/IF_ID_reg[44]  ( .D(\i_MIPS/N61 ), .CK(clk), .RN(n6316), .Q(
        \i_MIPS/Sign_Extend[12] ), .QN(\i_MIPS/n509 ) );
  DFFRX4 \i_MIPS/IF_ID_reg[43]  ( .D(\i_MIPS/N60 ), .CK(clk), .RN(n6316), .Q(
        \i_MIPS/Sign_Extend[11] ), .QN(\i_MIPS/n510 ) );
  DFFRX4 \i_MIPS/ID_EX_reg[106]  ( .D(\i_MIPS/n412 ), .CK(clk), .RN(n6321), 
        .Q(\i_MIPS/ID_EX[106] ), .QN(\i_MIPS/n250 ) );
  DFFRX4 \i_MIPS/ID_EX_reg[42]  ( .D(\i_MIPS/n365 ), .CK(clk), .RN(n6325), 
        .QN(\i_MIPS/n242 ) );
  DFFRHQX8 \i_MIPS/ID_EX_reg[80]  ( .D(\i_MIPS/n441 ), .CK(clk), .RN(n6318), 
        .Q(n3976) );
  DFFRHQX8 \i_MIPS/EX_MEM_reg[10]  ( .D(\i_MIPS/n394 ), .CK(clk), .RN(n6322), 
        .Q(n3965) );
  DFFRX2 \i_MIPS/ID_EX_reg[113]  ( .D(\i_MIPS/n451 ), .CK(clk), .RN(n6315), 
        .Q(\i_MIPS/ID_EX[113] ), .QN(\i_MIPS/n261 ) );
  DFFRX4 \D_cache/cache_reg[3][36]  ( .D(\D_cache/n1505 ), .CK(clk), .RN(n6199), .Q(\D_cache/cache[3][36] ) );
  DFFRX4 \D_cache/cache_reg[2][36]  ( .D(\D_cache/n1506 ), .CK(clk), .RN(n6199), .Q(\D_cache/cache[2][36] ) );
  DFFRX2 \i_MIPS/ID_EX_reg[109]  ( .D(\i_MIPS/n415 ), .CK(clk), .RN(n6320), 
        .QN(\i_MIPS/n256 ) );
  DFFRX4 \i_MIPS/IF_ID_reg[45]  ( .D(\i_MIPS/N62 ), .CK(clk), .RN(n6316), .Q(
        \i_MIPS/Sign_Extend[13] ), .QN(\i_MIPS/n508 ) );
  DFFRX4 \i_MIPS/PC/PC_o_reg[31]  ( .D(\i_MIPS/PC/n65 ), .CK(clk), .RN(n6309), 
        .Q(ICACHE_addr[29]), .QN(\i_MIPS/PC/n33 ) );
  DFFRX4 \i_MIPS/IF_ID_reg[52]  ( .D(\i_MIPS/N69 ), .CK(clk), .RN(n6315), .Q(
        \i_MIPS/jump_addr[22] ), .QN(\i_MIPS/n501 ) );
  DFFRX4 \i_MIPS/ID_EX_reg[87]  ( .D(\i_MIPS/n434 ), .CK(clk), .RN(n6318), .Q(
        \i_MIPS/ID_EX[87] ), .QN(n4776) );
  DFFRX4 \i_MIPS/ID_EX_reg[101]  ( .D(\i_MIPS/n420 ), .CK(clk), .RN(n6319), 
        .Q(\i_MIPS/ID_EX[101] ) );
  DFFRX2 \i_MIPS/ID_EX_reg[50]  ( .D(\i_MIPS/n349 ), .CK(clk), .RN(n6326), .Q(
        \i_MIPS/ID_EX[50] ), .QN(\i_MIPS/n226 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[110]  ( .D(\i_MIPS/n416 ), .CK(clk), .RN(n6320), 
        .QN(\i_MIPS/n258 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[108]  ( .D(\i_MIPS/n414 ), .CK(clk), .RN(n6320), 
        .Q(n4673), .QN(\i_MIPS/n254 ) );
  DFFRX4 \i_MIPS/IF_ID_reg[40]  ( .D(\i_MIPS/N57 ), .CK(clk), .RN(n6316), .Q(
        \i_MIPS/Sign_Extend[8] ), .QN(\i_MIPS/n513 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[45]  ( .D(\i_MIPS/n359 ), .CK(clk), .RN(n6325), 
        .QN(\i_MIPS/n236 ) );
  DFFRX4 \i_MIPS/ID_EX_reg[43]  ( .D(\i_MIPS/n363 ), .CK(clk), .RN(n6325), .Q(
        \i_MIPS/ID_EX[43] ), .QN(\i_MIPS/n240 ) );
  DFFRHQX8 \i_MIPS/ID_EX_reg[75]  ( .D(\i_MIPS/n446 ), .CK(clk), .RN(n6317), 
        .Q(n3873) );
  DFFRHQX8 \i_MIPS/EX_MEM_reg[11]  ( .D(\i_MIPS/n393 ), .CK(clk), .RN(n6322), 
        .Q(n3859) );
  DFFRX4 \i_MIPS/IF_ID_reg[36]  ( .D(\i_MIPS/N53 ), .CK(clk), .RN(n6317), .Q(
        n168), .QN(\i_MIPS/n517 ) );
  DFFRX4 \i_MIPS/IF_ID_reg[35]  ( .D(\i_MIPS/N52 ), .CK(clk), .RN(n6317), .Q(
        \i_MIPS/Sign_Extend[3] ), .QN(\i_MIPS/n518 ) );
  DFFRX4 \i_MIPS/IF_ID_reg[41]  ( .D(\i_MIPS/N58 ), .CK(clk), .RN(n6316), .Q(
        \i_MIPS/Sign_Extend[9] ), .QN(\i_MIPS/n512 ) );
  DFFRX4 \D_cache/cache_reg[0][57]  ( .D(\D_cache/n1340 ), .CK(clk), .RN(n6185), .Q(\D_cache/cache[0][57] ), .QN(n1260) );
  DFFRX4 \D_cache/cache_reg[1][57]  ( .D(\D_cache/n1339 ), .CK(clk), .RN(n6185), .Q(\D_cache/cache[1][57] ), .QN(n2880) );
  DFFRX4 \D_cache/cache_reg[4][57]  ( .D(\D_cache/n1336 ), .CK(clk), .RN(n6185), .Q(\D_cache/cache[4][57] ), .QN(n1306) );
  DFFRX4 \D_cache/cache_reg[5][57]  ( .D(\D_cache/n1335 ), .CK(clk), .RN(n6185), .Q(\D_cache/cache[5][57] ), .QN(n2944) );
  DFFRX4 \D_cache/cache_reg[7][57]  ( .D(\D_cache/n1333 ), .CK(clk), .RN(n6185), .Q(\D_cache/cache[7][57] ), .QN(n2867) );
  DFFRX4 \D_cache/cache_reg[6][57]  ( .D(\D_cache/n1334 ), .CK(clk), .RN(n6185), .Q(\D_cache/cache[6][57] ), .QN(n1247) );
  DFFRX4 \D_cache/cache_reg[0][36]  ( .D(\D_cache/n1508 ), .CK(clk), .RN(n6199), .Q(\D_cache/cache[0][36] ), .QN(n714) );
  DFFRX4 \D_cache/cache_reg[1][36]  ( .D(\D_cache/n1507 ), .CK(clk), .RN(n6199), .Q(\D_cache/cache[1][36] ), .QN(n2336) );
  DFFRX4 \D_cache/cache_reg[0][32]  ( .D(\D_cache/n1540 ), .CK(clk), .RN(n6202), .Q(\D_cache/cache[0][32] ), .QN(n1242) );
  DFFRX4 \D_cache/cache_reg[4][36]  ( .D(\D_cache/n1504 ), .CK(clk), .RN(n6199), .Q(\D_cache/cache[4][36] ), .QN(n713) );
  DFFRX4 \D_cache/cache_reg[5][36]  ( .D(\D_cache/n1503 ), .CK(clk), .RN(n6199), .Q(\D_cache/cache[5][36] ), .QN(n2335) );
  DFFRX4 \D_cache/cache_reg[6][36]  ( .D(\D_cache/n1502 ), .CK(clk), .RN(n6199), .Q(\D_cache/cache[6][36] ), .QN(n2331) );
  DFFRX4 \D_cache/cache_reg[1][32]  ( .D(\D_cache/n1539 ), .CK(clk), .RN(n6202), .Q(\D_cache/cache[1][32] ), .QN(n2861) );
  DFFRX4 \D_cache/cache_reg[4][32]  ( .D(\D_cache/n1536 ), .CK(clk), .RN(n6201), .Q(\D_cache/cache[4][32] ), .QN(n710) );
  DFFRX4 \D_cache/cache_reg[5][32]  ( .D(\D_cache/n1535 ), .CK(clk), .RN(n6201), .Q(\D_cache/cache[5][32] ), .QN(n2332) );
  DFFRX4 \D_cache/cache_reg[6][32]  ( .D(\D_cache/n1534 ), .CK(clk), .RN(n6201), .Q(\D_cache/cache[6][32] ), .QN(n2166) );
  DFFRX4 \D_cache/cache_reg[7][32]  ( .D(\D_cache/n1533 ), .CK(clk), .RN(n6201), .Q(\D_cache/cache[7][32] ), .QN(n547) );
  DFFRX4 \D_cache/cache_reg[4][41]  ( .D(\D_cache/n1464 ), .CK(clk), .RN(n6195), .Q(\D_cache/cache[4][41] ), .QN(n712) );
  DFFRX4 \D_cache/cache_reg[5][41]  ( .D(\D_cache/n1463 ), .CK(clk), .RN(n6195), .Q(\D_cache/cache[5][41] ), .QN(n2334) );
  DFFRX4 \D_cache/cache_reg[4][50]  ( .D(\D_cache/n1392 ), .CK(clk), .RN(n6189), .Q(\D_cache/cache[4][50] ) );
  DFFRX4 \D_cache/cache_reg[5][50]  ( .D(\D_cache/n1391 ), .CK(clk), .RN(n6189), .Q(\D_cache/cache[5][50] ), .QN(n2041) );
  DFFRX4 \D_cache/cache_reg[1][63]  ( .D(\D_cache/n1291 ), .CK(clk), .RN(n6181), .Q(\D_cache/cache[1][63] ), .QN(n2339) );
  DFFRX4 \D_cache/cache_reg[6][41]  ( .D(\D_cache/n1462 ), .CK(clk), .RN(n6195), .Q(\D_cache/cache[6][41] ), .QN(n2158) );
  DFFRX4 \D_cache/cache_reg[7][41]  ( .D(\D_cache/n1461 ), .CK(clk), .RN(n6195), .Q(\D_cache/cache[7][41] ), .QN(n539) );
  DFFRX4 \D_cache/cache_reg[6][50]  ( .D(\D_cache/n1390 ), .CK(clk), .RN(n6189), .Q(\D_cache/cache[6][50] ), .QN(n718) );
  DFFRX4 \D_cache/cache_reg[7][50]  ( .D(\D_cache/n1389 ), .CK(clk), .RN(n6189), .Q(\D_cache/cache[7][50] ), .QN(n2340) );
  DFFRX4 \D_cache/cache_reg[0][63]  ( .D(\D_cache/n1292 ), .CK(clk), .RN(n6181), .Q(\D_cache/cache[0][63] ), .QN(n717) );
  DFFRX4 \D_cache/cache_reg[4][63]  ( .D(\D_cache/n1288 ), .CK(clk), .RN(n6181), .Q(\D_cache/cache[4][63] ), .QN(n1256) );
  DFFRX4 \D_cache/cache_reg[5][63]  ( .D(\D_cache/n1287 ), .CK(clk), .RN(n6181), .Q(\D_cache/cache[5][63] ), .QN(n2876) );
  DFFRX4 \D_cache/cache_reg[6][63]  ( .D(\D_cache/n1286 ), .CK(clk), .RN(n6181), .Q(\D_cache/cache[6][63] ), .QN(n715) );
  DFFRX4 \D_cache/cache_reg[7][63]  ( .D(\D_cache/n1285 ), .CK(clk), .RN(n6181), .Q(\D_cache/cache[7][63] ), .QN(n2337) );
  DFFRX4 \D_cache/cache_reg[2][57]  ( .D(\D_cache/n1338 ), .CK(clk), .RN(n6185), .Q(\D_cache/cache[2][57] ), .QN(n1245) );
  DFFRX4 \D_cache/cache_reg[3][57]  ( .D(\D_cache/n1337 ), .CK(clk), .RN(n6185), .Q(\D_cache/cache[3][57] ), .QN(n2865) );
  DFFRX4 \D_cache/cache_reg[2][32]  ( .D(\D_cache/n1538 ), .CK(clk), .RN(n6202), .Q(\D_cache/cache[2][32] ), .QN(n2162) );
  DFFRX4 \D_cache/cache_reg[3][32]  ( .D(\D_cache/n1537 ), .CK(clk), .RN(n6202), .Q(\D_cache/cache[3][32] ), .QN(n543) );
  DFFRX4 \D_cache/cache_reg[0][41]  ( .D(\D_cache/n1468 ), .CK(clk), .RN(n6196), .Q(\D_cache/cache[0][41] ), .QN(n2168) );
  DFFRX4 \D_cache/cache_reg[1][41]  ( .D(\D_cache/n1467 ), .CK(clk), .RN(n6196), .Q(\D_cache/cache[1][41] ), .QN(n549) );
  DFFRX4 \D_cache/cache_reg[2][41]  ( .D(\D_cache/n1466 ), .CK(clk), .RN(n6196), .Q(\D_cache/cache[2][41] ), .QN(n2163) );
  DFFRX4 \D_cache/cache_reg[3][41]  ( .D(\D_cache/n1465 ), .CK(clk), .RN(n6196), .Q(\D_cache/cache[3][41] ), .QN(n544) );
  DFFRX4 \D_cache/cache_reg[0][50]  ( .D(\D_cache/n1396 ), .CK(clk), .RN(n6190), .Q(\D_cache/cache[0][50] ), .QN(n719) );
  DFFRX4 \D_cache/cache_reg[1][50]  ( .D(\D_cache/n1395 ), .CK(clk), .RN(n6190), .Q(\D_cache/cache[1][50] ), .QN(n2341) );
  DFFRX4 \D_cache/cache_reg[2][50]  ( .D(\D_cache/n1394 ), .CK(clk), .RN(n6190), .Q(\D_cache/cache[2][50] ), .QN(n711) );
  DFFRX4 \D_cache/cache_reg[3][50]  ( .D(\D_cache/n1393 ), .CK(clk), .RN(n6190), .Q(\D_cache/cache[3][50] ), .QN(n2333) );
  DFFRX4 \D_cache/cache_reg[2][63]  ( .D(\D_cache/n1290 ), .CK(clk), .RN(n6181), .Q(\D_cache/cache[2][63] ), .QN(n716) );
  DFFRX4 \D_cache/cache_reg[3][63]  ( .D(\D_cache/n1289 ), .CK(clk), .RN(n6181), .Q(\D_cache/cache[3][63] ), .QN(n2338) );
  DFFRX4 \D_cache/cache_reg[0][56]  ( .D(\D_cache/n1348 ), .CK(clk), .RN(n6186), .Q(\D_cache/cache[0][56] ), .QN(n1259) );
  DFFRX4 \D_cache/cache_reg[1][56]  ( .D(\D_cache/n1347 ), .CK(clk), .RN(n6186), .Q(\D_cache/cache[1][56] ), .QN(n2879) );
  DFFRX4 \D_cache/cache_reg[4][56]  ( .D(\D_cache/n1344 ), .CK(clk), .RN(n6185), .Q(\D_cache/cache[4][56] ), .QN(n1309) );
  DFFRX4 \D_cache/cache_reg[5][56]  ( .D(\D_cache/n1343 ), .CK(clk), .RN(n6185), .Q(\D_cache/cache[5][56] ), .QN(n2947) );
  DFFRX4 \D_cache/cache_reg[7][56]  ( .D(\D_cache/n1341 ), .CK(clk), .RN(n6185), .Q(\D_cache/cache[7][56] ), .QN(n2866) );
  DFFRX4 \D_cache/cache_reg[6][56]  ( .D(\D_cache/n1342 ), .CK(clk), .RN(n6185), .Q(\D_cache/cache[6][56] ), .QN(n1246) );
  DFFRX4 \D_cache/cache_reg[2][56]  ( .D(\D_cache/n1346 ), .CK(clk), .RN(n6186), .Q(\D_cache/cache[2][56] ), .QN(n1258) );
  DFFRX4 \D_cache/cache_reg[3][56]  ( .D(\D_cache/n1345 ), .CK(clk), .RN(n6186), .Q(\D_cache/cache[3][56] ), .QN(n2878) );
  DFFRX4 \D_cache/cache_reg[0][45]  ( .D(\D_cache/n1436 ), .CK(clk), .RN(n6193), .Q(\D_cache/cache[0][45] ), .QN(n1249) );
  DFFRX4 \D_cache/cache_reg[1][45]  ( .D(\D_cache/n1435 ), .CK(clk), .RN(n6193), .Q(\D_cache/cache[1][45] ), .QN(n2869) );
  DFFRX4 \D_cache/cache_reg[4][45]  ( .D(\D_cache/n1432 ), .CK(clk), .RN(n6193), .Q(\D_cache/cache[4][45] ), .QN(n1253) );
  DFFRX4 \D_cache/cache_reg[5][45]  ( .D(\D_cache/n1431 ), .CK(clk), .RN(n6193), .Q(\D_cache/cache[5][45] ), .QN(n2873) );
  DFFRX4 \D_cache/cache_reg[6][45]  ( .D(\D_cache/n1430 ), .CK(clk), .RN(n6193), .Q(\D_cache/cache[6][45] ), .QN(n1248) );
  DFFRX4 \D_cache/cache_reg[7][45]  ( .D(\D_cache/n1429 ), .CK(clk), .RN(n6193), .Q(\D_cache/cache[7][45] ), .QN(n2868) );
  DFFRX4 \D_cache/cache_reg[0][51]  ( .D(\D_cache/n1388 ), .CK(clk), .RN(n6189), .Q(\D_cache/cache[0][51] ), .QN(n1252) );
  DFFRX4 \D_cache/cache_reg[1][51]  ( .D(\D_cache/n1387 ), .CK(clk), .RN(n6189), .Q(\D_cache/cache[1][51] ), .QN(n2872) );
  DFFRX4 \D_cache/cache_reg[4][51]  ( .D(\D_cache/n1384 ), .CK(clk), .RN(n6189), .Q(\D_cache/cache[4][51] ), .QN(n1254) );
  DFFRX4 \D_cache/cache_reg[5][51]  ( .D(\D_cache/n1383 ), .CK(clk), .RN(n6189), .Q(\D_cache/cache[5][51] ), .QN(n2874) );
  DFFRX4 \D_cache/cache_reg[6][51]  ( .D(\D_cache/n1382 ), .CK(clk), .RN(n6189), .Q(\D_cache/cache[6][51] ), .QN(n2157) );
  DFFRX4 \D_cache/cache_reg[7][51]  ( .D(\D_cache/n1381 ), .CK(clk), .RN(n6189), .Q(\D_cache/cache[7][51] ), .QN(n538) );
  DFFRX4 \D_cache/cache_reg[2][45]  ( .D(\D_cache/n1434 ), .CK(clk), .RN(n6193), .Q(\D_cache/cache[2][45] ), .QN(n2164) );
  DFFRX4 \D_cache/cache_reg[3][45]  ( .D(\D_cache/n1433 ), .CK(clk), .RN(n6193), .Q(\D_cache/cache[3][45] ), .QN(n545) );
  DFFRX4 \D_cache/cache_reg[2][51]  ( .D(\D_cache/n1386 ), .CK(clk), .RN(n6189), .Q(\D_cache/cache[2][51] ), .QN(n1251) );
  DFFRX4 \D_cache/cache_reg[3][51]  ( .D(\D_cache/n1385 ), .CK(clk), .RN(n6189), .Q(\D_cache/cache[3][51] ), .QN(n2871) );
  DFFRX4 \i_MIPS/IF_ID_reg[37]  ( .D(\i_MIPS/N54 ), .CK(clk), .RN(n6317), .Q(
        \i_MIPS/Sign_Extend[5] ), .QN(\i_MIPS/n516 ) );
  DFFRX4 \i_MIPS/ID_EX_reg[47]  ( .D(\i_MIPS/n355 ), .CK(clk), .RN(n6325), .Q(
        \i_MIPS/ID_EX[47] ), .QN(\i_MIPS/n232 ) );
  DFFRX4 \i_MIPS/IF_ID_reg[62]  ( .D(\i_MIPS/N79 ), .CK(clk), .RN(n6320), .Q(
        \i_MIPS/IR[30] ), .QN(\i_MIPS/n255 ) );
  DFFRX4 \i_MIPS/IF_ID_reg[60]  ( .D(\i_MIPS/N77 ), .CK(clk), .RN(n6320), .Q(
        \i_MIPS/IR[28] ), .QN(\i_MIPS/n251 ) );
  DFFRX4 \i_MIPS/IF_ID_reg[59]  ( .D(\i_MIPS/N76 ), .CK(clk), .RN(n6320), .Q(
        \i_MIPS/IR[27] ), .QN(\i_MIPS/n249 ) );
  DFFRX4 \i_MIPS/IF_ID_reg[57]  ( .D(\i_MIPS/N74 ), .CK(clk), .RN(n6315), .Q(
        n3001), .QN(\i_MIPS/n496 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[68]  ( .D(\i_MIPS/n313 ), .CK(clk), .RN(n6329), .Q(
        \i_MIPS/ID_EX[68] ), .QN(\i_MIPS/n190 ) );
  DFFRX4 \i_MIPS/ID_EX_reg[100]  ( .D(\i_MIPS/n421 ), .CK(clk), .RN(n6319), 
        .Q(\i_MIPS/ID_EX[100] ) );
  DFFRHQX8 \i_MIPS/ID_EX_reg[79]  ( .D(\i_MIPS/n442 ), .CK(clk), .RN(n6318), 
        .Q(n3704) );
  DFFRHQX8 \i_MIPS/ID_EX_reg[82]  ( .D(\i_MIPS/n439 ), .CK(clk), .RN(n6318), 
        .Q(n3673) );
  DFFRX2 \i_MIPS/ID_EX_reg[48]  ( .D(\i_MIPS/n353 ), .CK(clk), .RN(n6326), .Q(
        \i_MIPS/ID_EX[48] ), .QN(\i_MIPS/n230 ) );
  DFFRX4 \i_MIPS/IF_ID_reg[32]  ( .D(\i_MIPS/N49 ), .CK(clk), .RN(n6314), .Q(
        \i_MIPS/Sign_Extend[0] ), .QN(\i_MIPS/n521 ) );
  DFFRHQX8 \i_MIPS/ID_EX_reg[6]  ( .D(\i_MIPS/n402 ), .CK(clk), .RN(n6321), 
        .Q(n3621) );
  DFFRHQX2 \i_MIPS/ID_EX_reg[51]  ( .D(\i_MIPS/n347 ), .CK(clk), .RN(n6326), 
        .Q(n3608) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[27]  ( .D(\i_MIPS/PC/n61 ), .CK(clk), .RN(n6309), 
        .Q(ICACHE_addr[25]), .QN(\i_MIPS/PC/n29 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[35]  ( .D(\i_MIPS/n369 ), .CK(clk), .RN(n6324), 
        .Q(n12955) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[21]  ( .D(\i_MIPS/PC/n55 ), .CK(clk), .RN(n6309), 
        .Q(ICACHE_addr[19]), .QN(\i_MIPS/PC/n23 ) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[9]  ( .D(\i_MIPS/PC/n43 ), .CK(clk), .RN(n6310), 
        .Q(ICACHE_addr[7]), .QN(\i_MIPS/PC/n11 ) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[18]  ( .D(\i_MIPS/PC/n52 ), .CK(clk), .RN(n6310), 
        .Q(ICACHE_addr[16]), .QN(\i_MIPS/PC/n20 ) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[23]  ( .D(\i_MIPS/PC/n57 ), .CK(clk), .RN(n6309), 
        .Q(ICACHE_addr[21]), .QN(\i_MIPS/PC/n25 ) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[20]  ( .D(\i_MIPS/PC/n54 ), .CK(clk), .RN(n6309), 
        .Q(ICACHE_addr[18]), .QN(\i_MIPS/PC/n22 ) );
  DFFRX4 \i_MIPS/IF_ID_reg[39]  ( .D(\i_MIPS/N56 ), .CK(clk), .RN(n6317), .Q(
        n1287), .QN(\i_MIPS/n514 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[42]  ( .D(\i_MIPS/N59 ), .CK(clk), .RN(n6316), .Q(
        \i_MIPS/Sign_Extend[10] ), .QN(\i_MIPS/n511 ) );
  DFFRHQX2 \i_MIPS/ID_EX_reg[41]  ( .D(\i_MIPS/n367 ), .CK(clk), .RN(n6324), 
        .Q(n3883) );
  DFFRX2 \i_MIPS/ID_EX_reg[49]  ( .D(\i_MIPS/n351 ), .CK(clk), .RN(n6326), .Q(
        n3555), .QN(\i_MIPS/n228 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[63]  ( .D(\i_MIPS/n323 ), .CK(clk), .RN(n6328), .Q(
        \i_MIPS/ID_EX[63] ), .QN(\i_MIPS/n200 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[65]  ( .D(\i_MIPS/n319 ), .CK(clk), .RN(n6328), .Q(
        \i_MIPS/ID_EX[65] ), .QN(\i_MIPS/n196 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[59]  ( .D(\i_MIPS/n331 ), .CK(clk), .RN(n6327), .Q(
        n3554), .QN(\i_MIPS/n208 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[52]  ( .D(\i_MIPS/n345 ), .CK(clk), .RN(n6326), .Q(
        n3553), .QN(\i_MIPS/n222 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[60]  ( .D(\i_MIPS/n329 ), .CK(clk), .RN(n6328), .Q(
        n3552), .QN(\i_MIPS/n206 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[2]  ( .D(\i_MIPS/N19 ), .CK(clk), .RN(n6330), .Q(
        \i_MIPS/IF_ID[2] ), .QN(\i_MIPS/n155 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[19]  ( .D(\i_MIPS/n385 ), .CK(clk), .RN(n6323), 
        .Q(n12971), .QN(n5005) );
  DFFRX1 \i_MIPS/EX_MEM_reg[33]  ( .D(\i_MIPS/n371 ), .CK(clk), .RN(n6324), 
        .Q(n12957), .QN(n4824) );
  DFFRX1 \i_MIPS/EX_MEM_reg[27]  ( .D(\i_MIPS/n377 ), .CK(clk), .RN(n6324), 
        .Q(n12963), .QN(n4825) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[16]  ( .D(\i_MIPS/PC/n50 ), .CK(clk), .RN(n6310), 
        .Q(ICACHE_addr[14]), .QN(\i_MIPS/PC/n18 ) );
  DFFRX1 \I_cache/cache_reg[5][141]  ( .D(n11712), .CK(clk), .RN(n6025), .Q(
        \I_cache/cache[5][141] ), .QN(n3017) );
  DFFRX1 \I_cache/cache_reg[2][141]  ( .D(n11715), .CK(clk), .RN(n6026), .Q(
        \I_cache/cache[2][141] ), .QN(n3013) );
  DFFRX1 \I_cache/cache_reg[6][152]  ( .D(n11623), .CK(clk), .RN(n6018), .Q(
        \I_cache/cache[6][152] ), .QN(n3012) );
  DFFRX1 \I_cache/cache_reg[0][141]  ( .D(n11717), .CK(clk), .RN(n6026), .Q(
        \I_cache/cache[0][141] ), .QN(n3011) );
  DFFRX1 \I_cache/cache_reg[6][141]  ( .D(n11711), .CK(clk), .RN(n6025), .Q(
        \I_cache/cache[6][141] ), .QN(n3010) );
  DFFRX1 \I_cache/cache_reg[3][152]  ( .D(n11626), .CK(clk), .RN(n6018), .Q(
        \I_cache/cache[3][152] ), .QN(n3009) );
  DFFRX1 \I_cache/cache_reg[1][152]  ( .D(n11628), .CK(clk), .RN(n6018), .Q(
        \I_cache/cache[1][152] ), .QN(n3008) );
  DFFRX2 \i_MIPS/IF_ID_reg[4]  ( .D(\i_MIPS/N21 ), .CK(clk), .RN(n6330), .Q(
        \i_MIPS/IF_ID[4] ), .QN(\i_MIPS/n157 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[105]  ( .D(\i_MIPS/n411 ), .CK(clk), .RN(n6321), 
        .Q(\i_MIPS/ID_EX[105] ), .QN(\i_MIPS/n248 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[38]  ( .D(\i_MIPS/n463 ), .CK(clk), .RN(n6314), .Q(
        \i_MIPS/ALUin1[29] ), .QN(n2961) );
  DFFRX2 \i_MIPS/ID_EX_reg[31]  ( .D(\i_MIPS/n470 ), .CK(clk), .RN(n6313), .Q(
        \i_MIPS/ALUin1[22] ), .QN(n2949) );
  DFFRX2 \D_cache/cache_reg[5][25]  ( .D(\D_cache/n1591 ), .CK(clk), .RN(n6206), .Q(\D_cache/cache[5][25] ), .QN(n2946) );
  DFFRX2 \D_cache/cache_reg[5][24]  ( .D(\D_cache/n1599 ), .CK(clk), .RN(n6207), .Q(\D_cache/cache[5][24] ), .QN(n2945) );
  DFFRX2 \i_MIPS/IF_ID_reg[3]  ( .D(\i_MIPS/N20 ), .CK(clk), .RN(n6330), .Q(
        \i_MIPS/IF_ID[3] ), .QN(\i_MIPS/n156 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[14]  ( .D(\i_MIPS/n487 ), .CK(clk), .RN(n6312), .Q(
        \i_MIPS/ALUin1[5] ), .QN(\i_MIPS/n296 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[26]  ( .D(\i_MIPS/n475 ), .CK(clk), .RN(n6313), .Q(
        \i_MIPS/ALUin1[17] ), .QN(n2921) );
  DFFRX2 \D_cache/cache_reg[1][24]  ( .D(\D_cache/n1603 ), .CK(clk), .RN(n6207), .Q(\D_cache/cache[1][24] ), .QN(n2882) );
  DFFRX2 \D_cache/cache_reg[3][24]  ( .D(\D_cache/n1601 ), .CK(clk), .RN(n6207), .Q(\D_cache/cache[3][24] ), .QN(n2881) );
  DFFRX2 \D_cache/cache_reg[1][25]  ( .D(\D_cache/n1595 ), .CK(clk), .RN(n6206), .Q(\D_cache/cache[1][25] ), .QN(n2877) );
  DFFRX2 \D_cache/cache_reg[5][20]  ( .D(\D_cache/n1631 ), .CK(clk), .RN(n6209), .Q(\D_cache/cache[5][20] ), .QN(n2875) );
  DFFRX2 \D_cache/cache_reg[1][20]  ( .D(\D_cache/n1635 ), .CK(clk), .RN(n6210), .Q(\D_cache/cache[1][20] ), .QN(n2870) );
  DFFRX2 \D_cache/cache_reg[3][25]  ( .D(\D_cache/n1593 ), .CK(clk), .RN(n6206), .Q(\D_cache/cache[3][25] ), .QN(n2864) );
  DFFRX2 \D_cache/cache_reg[7][25]  ( .D(\D_cache/n1589 ), .CK(clk), .RN(n6206), .Q(\D_cache/cache[7][25] ), .QN(n2863) );
  DFFRX1 \D_cache/cache_reg[1][52]  ( .D(\D_cache/n1379 ), .CK(clk), .RN(n6188), .Q(\D_cache/cache[1][52] ), .QN(n2860) );
  DFFRX2 \i_MIPS/ID_EX_reg[34]  ( .D(\i_MIPS/n467 ), .CK(clk), .RN(n6313), .Q(
        \i_MIPS/ALUin1[25] ), .QN(n2184) );
  DFFRX1 \D_cache/cache_reg[6][52]  ( .D(\D_cache/n1374 ), .CK(clk), .RN(n6188), .Q(\D_cache/cache[6][52] ), .QN(n2167) );
  DFFRX1 \D_cache/cache_reg[2][52]  ( .D(\D_cache/n1378 ), .CK(clk), .RN(n6188), .Q(\D_cache/cache[2][52] ), .QN(n2165) );
  DFFRX2 \D_cache/cache_reg[6][20]  ( .D(\D_cache/n1630 ), .CK(clk), .RN(n6209), .Q(\D_cache/cache[6][20] ), .QN(n2161) );
  DFFRX2 \D_cache/cache_reg[2][20]  ( .D(\D_cache/n1634 ), .CK(clk), .RN(n6210), .Q(\D_cache/cache[2][20] ), .QN(n2160) );
  DFFRX2 \D_cache/cache_reg[6][24]  ( .D(\D_cache/n1598 ), .CK(clk), .RN(n6207), .Q(\D_cache/cache[6][24] ), .QN(n2159) );
  DFFRX1 \D_cache/cache_reg[4][52]  ( .D(\D_cache/n1376 ), .CK(clk), .RN(n6188), .Q(\D_cache/cache[4][52] ), .QN(n2156) );
  DFFRX2 \i_MIPS/EX_MEM_reg[69]  ( .D(\i_MIPS/n407 ), .CK(clk), .RN(n6321), 
        .Q(\i_MIPS/Reg_W[0] ), .QN(n1988) );
  DFFRX2 \i_MIPS/ID_EX_reg[36]  ( .D(\i_MIPS/n465 ), .CK(clk), .RN(n6314), .Q(
        \i_MIPS/ALUin1[27] ), .QN(n3861) );
  DFFRX2 \D_cache/cache_reg[4][25]  ( .D(\D_cache/n1592 ), .CK(clk), .RN(n6206), .Q(\D_cache/cache[4][25] ), .QN(n1308) );
  DFFRX2 \D_cache/cache_reg[4][24]  ( .D(\D_cache/n1600 ), .CK(clk), .RN(n6207), .Q(\D_cache/cache[4][24] ), .QN(n1307) );
  DFFRX1 \i_MIPS/EX_MEM_reg[17]  ( .D(\i_MIPS/n387 ), .CK(clk), .RN(n6323), 
        .Q(n12973), .QN(n1303) );
  DFFRX2 \i_MIPS/ID_EX_reg[27]  ( .D(\i_MIPS/n474 ), .CK(clk), .RN(n6313), .Q(
        \i_MIPS/ALUin1[18] ), .QN(n1264) );
  DFFRX2 \D_cache/cache_reg[0][24]  ( .D(\D_cache/n1604 ), .CK(clk), .RN(n6207), .Q(\D_cache/cache[0][24] ), .QN(n1262) );
  DFFRX2 \D_cache/cache_reg[2][24]  ( .D(\D_cache/n1602 ), .CK(clk), .RN(n6207), .Q(\D_cache/cache[2][24] ), .QN(n1261) );
  DFFRX2 \D_cache/cache_reg[0][25]  ( .D(\D_cache/n1596 ), .CK(clk), .RN(n6206), .Q(\D_cache/cache[0][25] ), .QN(n1257) );
  DFFRX2 \D_cache/cache_reg[2][25]  ( .D(\D_cache/n1594 ), .CK(clk), .RN(n6206), .Q(\D_cache/cache[2][25] ), .QN(n1244) );
  DFFRX2 \D_cache/cache_reg[6][25]  ( .D(\D_cache/n1590 ), .CK(clk), .RN(n6206), .Q(\D_cache/cache[6][25] ), .QN(n1243) );
  DFFRX1 \D_cache/cache_reg[0][52]  ( .D(\D_cache/n1380 ), .CK(clk), .RN(n6188), .Q(\D_cache/cache[0][52] ), .QN(n1241) );
  DFFRX2 \i_MIPS/ID_EX_reg[25]  ( .D(\i_MIPS/n476 ), .CK(clk), .RN(n6313), .Q(
        \i_MIPS/ALUin1[16] ), .QN(n959) );
  DFFRX1 \D_cache/cache_reg[7][52]  ( .D(\D_cache/n1373 ), .CK(clk), .RN(n6188), .Q(\D_cache/cache[7][52] ), .QN(n548) );
  DFFRX1 \D_cache/cache_reg[3][52]  ( .D(\D_cache/n1377 ), .CK(clk), .RN(n6188), .Q(\D_cache/cache[3][52] ), .QN(n546) );
  DFFRX2 \D_cache/cache_reg[7][24]  ( .D(\D_cache/n1597 ), .CK(clk), .RN(n6207), .Q(\D_cache/cache[7][24] ), .QN(n540) );
  DFFRX1 \D_cache/cache_reg[5][52]  ( .D(\D_cache/n1375 ), .CK(clk), .RN(n6188), .Q(\D_cache/cache[5][52] ), .QN(n537) );
  DFFRX2 \i_MIPS/EX_MEM_reg[70]  ( .D(\i_MIPS/n406 ), .CK(clk), .RN(n6321), 
        .Q(\i_MIPS/Reg_W[1] ), .QN(n4833) );
  DFFRX1 \i_MIPS/EX_MEM_reg[12]  ( .D(\i_MIPS/n392 ), .CK(clk), .RN(n6322), 
        .Q(n12978), .QN(n355) );
  DFFRX1 \i_MIPS/EX_MEM_reg[21]  ( .D(\i_MIPS/n383 ), .CK(clk), .RN(n6323), 
        .Q(n12969), .QN(n1329) );
  DFFRX1 \i_MIPS/EX_MEM_reg[4]  ( .D(\i_MIPS/n409 ), .CK(clk), .RN(n6321), 
        .QN(\i_MIPS/n245 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[33]  ( .D(\i_MIPS/n468 ), .CK(clk), .RN(n6313), .Q(
        \i_MIPS/ALUin1[24] ), .QN(n344) );
  DFFRX2 \i_MIPS/ID_EX_reg[28]  ( .D(\i_MIPS/n473 ), .CK(clk), .RN(n6313), .Q(
        \i_MIPS/ALUin1[19] ), .QN(n336) );
  DFFRX2 \i_MIPS/ID_EX_reg[39]  ( .D(\i_MIPS/n462 ), .CK(clk), .RN(n6314), .Q(
        \i_MIPS/ALUin1[30] ), .QN(\i_MIPS/n271 ) );
  DFFRX2 \i_MIPS/EX_MEM_reg[71]  ( .D(\i_MIPS/n405 ), .CK(clk), .RN(n6321), 
        .Q(\i_MIPS/Reg_W[2] ), .QN(n223) );
  DFFRX2 \i_MIPS/ID_EX_reg[32]  ( .D(\i_MIPS/n469 ), .CK(clk), .RN(n6313), .Q(
        \i_MIPS/ALUin1[23] ), .QN(n183) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[17]  ( .D(\i_MIPS/PC/n51 ), .CK(clk), .RN(n6310), 
        .Q(ICACHE_addr[15]), .QN(\i_MIPS/PC/n19 ) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[19]  ( .D(\i_MIPS/PC/n53 ), .CK(clk), .RN(n6310), 
        .Q(ICACHE_addr[17]), .QN(\i_MIPS/PC/n21 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[16]  ( .D(\i_MIPS/n388 ), .CK(clk), .RN(n6323), 
        .Q(n12974), .QN(n5006) );
  DFFRX1 \i_MIPS/EX_MEM_reg[20]  ( .D(\i_MIPS/n384 ), .CK(clk), .RN(n6323), 
        .Q(n12970), .QN(net118925) );
  DFFRX1 \i_MIPS/EX_MEM_reg[56]  ( .D(\i_MIPS/n328 ), .CK(clk), .RN(n6328), 
        .Q(n12994), .QN(\i_MIPS/n205 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[57]  ( .D(\i_MIPS/n326 ), .CK(clk), .RN(n6328), 
        .Q(n12993), .QN(\i_MIPS/n203 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[63]  ( .D(\i_MIPS/n314 ), .CK(clk), .RN(n6329), 
        .Q(n12987), .QN(\i_MIPS/n191 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[49]  ( .D(\i_MIPS/n342 ), .CK(clk), .RN(n6326), 
        .Q(n13001), .QN(\i_MIPS/n219 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[43]  ( .D(\i_MIPS/n354 ), .CK(clk), .RN(n6325), 
        .Q(n13007), .QN(\i_MIPS/n231 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[48]  ( .D(\i_MIPS/n344 ), .CK(clk), .RN(n6326), 
        .Q(n13002), .QN(\i_MIPS/n221 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[59]  ( .D(\i_MIPS/n322 ), .CK(clk), .RN(n6328), 
        .Q(n12991), .QN(\i_MIPS/n199 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[62]  ( .D(\i_MIPS/n316 ), .CK(clk), .RN(n6329), 
        .Q(n12988), .QN(\i_MIPS/n193 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[53]  ( .D(\i_MIPS/n334 ), .CK(clk), .RN(n6327), 
        .Q(n12997), .QN(\i_MIPS/n211 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[64]  ( .D(\i_MIPS/n312 ), .CK(clk), .RN(n6329), 
        .Q(n12986), .QN(\i_MIPS/n189 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[37]  ( .D(\i_MIPS/n366 ), .CK(clk), .RN(n6324), 
        .Q(n13013), .QN(\i_MIPS/n243 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[52]  ( .D(\i_MIPS/n336 ), .CK(clk), .RN(n6327), 
        .Q(n12998), .QN(\i_MIPS/n213 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[40]  ( .D(\i_MIPS/n360 ), .CK(clk), .RN(n6325), 
        .Q(n13010), .QN(\i_MIPS/n237 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[42]  ( .D(\i_MIPS/n356 ), .CK(clk), .RN(n6325), 
        .Q(n13008), .QN(\i_MIPS/n233 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[39]  ( .D(\i_MIPS/n362 ), .CK(clk), .RN(n6325), 
        .Q(n13011), .QN(\i_MIPS/n239 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[38]  ( .D(\i_MIPS/n364 ), .CK(clk), .RN(n6325), 
        .Q(n13012), .QN(\i_MIPS/n241 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[41]  ( .D(\i_MIPS/n358 ), .CK(clk), .RN(n6325), 
        .Q(n13009), .QN(\i_MIPS/n235 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[44]  ( .D(\i_MIPS/n352 ), .CK(clk), .RN(n6326), 
        .Q(n13006), .QN(\i_MIPS/n229 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[45]  ( .D(\i_MIPS/n350 ), .CK(clk), .RN(n6326), 
        .Q(n13005), .QN(\i_MIPS/n227 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[46]  ( .D(\i_MIPS/n348 ), .CK(clk), .RN(n6326), 
        .Q(n13004), .QN(\i_MIPS/n225 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[47]  ( .D(\i_MIPS/n346 ), .CK(clk), .RN(n6326), 
        .Q(n13003), .QN(\i_MIPS/n223 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[50]  ( .D(\i_MIPS/n340 ), .CK(clk), .RN(n6327), 
        .Q(n13000), .QN(\i_MIPS/n217 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[51]  ( .D(\i_MIPS/n338 ), .CK(clk), .RN(n6327), 
        .Q(n12999), .QN(\i_MIPS/n215 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[54]  ( .D(\i_MIPS/n332 ), .CK(clk), .RN(n6327), 
        .Q(n12996), .QN(\i_MIPS/n209 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[55]  ( .D(\i_MIPS/n330 ), .CK(clk), .RN(n6327), 
        .Q(n12995), .QN(\i_MIPS/n207 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[58]  ( .D(\i_MIPS/n324 ), .CK(clk), .RN(n6328), 
        .Q(n12992), .QN(\i_MIPS/n201 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[60]  ( .D(\i_MIPS/n320 ), .CK(clk), .RN(n6328), 
        .Q(n12990), .QN(\i_MIPS/n197 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[61]  ( .D(\i_MIPS/n318 ), .CK(clk), .RN(n6328), 
        .Q(n12989), .QN(\i_MIPS/n195 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[65]  ( .D(\i_MIPS/n310 ), .CK(clk), .RN(n6329), 
        .Q(n12985), .QN(\i_MIPS/n187 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[66]  ( .D(\i_MIPS/n308 ), .CK(clk), .RN(n6329), 
        .Q(n12984), .QN(\i_MIPS/n185 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[67]  ( .D(\i_MIPS/n306 ), .CK(clk), .RN(n6329), 
        .Q(n12983), .QN(\i_MIPS/n183 ) );
  DFFRX1 \i_MIPS/EX_MEM_reg[68]  ( .D(\i_MIPS/n304 ), .CK(clk), .RN(n6330), 
        .Q(n12982), .QN(\i_MIPS/n181 ) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[28]  ( .D(\i_MIPS/PC/n62 ), .CK(clk), .RN(n6309), 
        .Q(ICACHE_addr[26]), .QN(\i_MIPS/PC/n30 ) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[14]  ( .D(\i_MIPS/PC/n48 ), .CK(clk), .RN(n6310), 
        .Q(ICACHE_addr[12]), .QN(\i_MIPS/PC/n16 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[94]  ( .D(\i_MIPS/n427 ), .CK(clk), .RN(n6319), .Q(
        \i_MIPS/ID_EX[94] ), .QN(n4782) );
  DFFRX2 \i_MIPS/ID_EX_reg[112]  ( .D(\i_MIPS/n450 ), .CK(clk), .RN(n6316), 
        .Q(\i_MIPS/ID_EX[112] ), .QN(\i_MIPS/n260 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[99]  ( .D(\i_MIPS/n422 ), .CK(clk), .RN(n6319), .Q(
        \i_MIPS/ID_EX[99] ) );
  DFFRX1 \i_MIPS/PC/PC_o_reg[8]  ( .D(\i_MIPS/PC/n42 ), .CK(clk), .RN(n6310), 
        .Q(ICACHE_addr[6]), .QN(\i_MIPS/PC/n10 ) );
  DFFRX2 \i_MIPS/ID_EX_reg[85]  ( .D(\i_MIPS/n436 ), .CK(clk), .RN(n6318), .Q(
        \i_MIPS/ID_EX[85] ), .QN(n4775) );
  DFFRX2 \i_MIPS/ID_EX_reg[98]  ( .D(\i_MIPS/n423 ), .CK(clk), .RN(n6319), .Q(
        \i_MIPS/ID_EX[98] ) );
  DFFRX2 \i_MIPS/ID_EX_reg[22]  ( .D(\i_MIPS/n479 ), .CK(clk), .RN(n6312), .Q(
        \i_MIPS/ALUin1[13] ), .QN(n2937) );
  DFFRX1 \D_cache/cache_reg[2][154]  ( .D(\D_cache/n562 ), .CK(clk), .RN(n6120), .Q(\D_cache/cache[2][154] ), .QN(n3975) );
  DFFRX1 \i_MIPS/ID_EX_reg[102]  ( .D(\i_MIPS/n419 ), .CK(clk), .RN(n6320), 
        .Q(\i_MIPS/ID_EX[102] ) );
  DFFRX1 \D_cache/cache_reg[1][149]  ( .D(\D_cache/n603 ), .CK(clk), .RN(n6124), .Q(\D_cache/cache[1][149] ) );
  DFFRX1 \D_cache/cache_reg[0][149]  ( .D(\D_cache/n604 ), .CK(clk), .RN(n6124), .Q(\D_cache/cache[0][149] ) );
  DFFRX1 \D_cache/cache_reg[3][145]  ( .D(\D_cache/n633 ), .CK(clk), .RN(n6126), .Q(\D_cache/cache[3][145] ) );
  DFFRX1 \D_cache/cache_reg[3][146]  ( .D(\D_cache/n625 ), .CK(clk), .RN(n6126), .Q(\D_cache/cache[3][146] ) );
  DFFRX2 \i_MIPS/ID_EX_reg[86]  ( .D(\i_MIPS/n435 ), .CK(clk), .RN(n6318), .Q(
        \i_MIPS/ID_EX[86] ), .QN(n4774) );
  DFFRX1 \i_MIPS/ID_EX_reg[97]  ( .D(\i_MIPS/n424 ), .CK(clk), .RN(n6319), .Q(
        \i_MIPS/ID_EX[97] ) );
  DFFRX1 \D_cache/cache_reg[1][137]  ( .D(\D_cache/n699 ), .CK(clk), .RN(n6132), .Q(\D_cache/cache[1][137] ) );
  DFFRX2 \i_MIPS/ID_EX_reg[96]  ( .D(\i_MIPS/n425 ), .CK(clk), .RN(n6319), .Q(
        \i_MIPS/ID_EX[96] ) );
  DFFRX2 \i_MIPS/ID_EX_reg[64]  ( .D(\i_MIPS/n321 ), .CK(clk), .RN(n6328), .Q(
        \i_MIPS/ID_EX[64] ), .QN(\i_MIPS/n198 ) );
  DFFRX1 \D_cache/cache_reg[3][144]  ( .D(\D_cache/n641 ), .CK(clk), .RN(n6127), .Q(\D_cache/cache[3][144] ), .QN(n3865) );
  DFFRX1 \D_cache/cache_reg[2][144]  ( .D(\D_cache/n642 ), .CK(clk), .RN(n6127), .Q(\D_cache/cache[2][144] ) );
  DFFRX1 \D_cache/cache_reg[6][132]  ( .D(\D_cache/n734 ), .CK(clk), .RN(n6135), .Q(\D_cache/cache[6][132] ) );
  DFFRX1 \D_cache/cache_reg[6][134]  ( .D(\D_cache/n718 ), .CK(clk), .RN(n6133), .Q(\D_cache/cache[6][134] ) );
  DFFRX1 \i_MIPS/ID_EX_reg[61]  ( .D(\i_MIPS/n327 ), .CK(clk), .RN(n6328), .Q(
        n3544), .QN(\i_MIPS/n204 ) );
  DFFRX1 \D_cache/cache_reg[6][148]  ( .D(\D_cache/n606 ), .CK(clk), .RN(n6124), .Q(\D_cache/cache[6][148] ) );
  DFFRX1 \D_cache/cache_reg[2][148]  ( .D(\D_cache/n610 ), .CK(clk), .RN(n6124), .Q(\D_cache/cache[2][148] ) );
  DFFRX1 \D_cache/cache_reg[6][144]  ( .D(\D_cache/n638 ), .CK(clk), .RN(n6127), .Q(\D_cache/cache[6][144] ) );
  DFFRX1 \D_cache/cache_reg[5][143]  ( .D(\D_cache/n647 ), .CK(clk), .RN(n6127), .Q(\D_cache/cache[5][143] ) );
  DFFRX2 \D_cache/cache_reg[0][20]  ( .D(\D_cache/n1636 ), .CK(clk), .RN(n6210), .Q(\D_cache/cache[0][20] ), .QN(n1250) );
  DFFRX2 \D_cache/cache_reg[4][20]  ( .D(\D_cache/n1632 ), .CK(clk), .RN(n6209), .Q(\D_cache/cache[4][20] ), .QN(n1255) );
  DFFRX2 \D_cache/cache_reg[7][20]  ( .D(\D_cache/n1629 ), .CK(clk), .RN(n6209), .Q(\D_cache/cache[7][20] ), .QN(n542) );
  DFFRX2 \D_cache/cache_reg[3][20]  ( .D(\D_cache/n1633 ), .CK(clk), .RN(n6210), .Q(\D_cache/cache[3][20] ), .QN(n541) );
  DFFRX2 \i_MIPS/ID_EX_reg[88]  ( .D(\i_MIPS/n433 ), .CK(clk), .RN(n6318), .Q(
        \i_MIPS/ID_EX[88] ), .QN(n4791) );
  DFFRX2 \i_MIPS/ID_EX_reg[69]  ( .D(\i_MIPS/n311 ), .CK(clk), .RN(n6329), .Q(
        \i_MIPS/ID_EX[69] ), .QN(\i_MIPS/n188 ) );
  DFFRX1 \D_cache/cache_reg[4][21]  ( .D(\D_cache/n1624 ), .CK(clk), .RN(n6209), .Q(\D_cache/cache[4][21] ) );
  DFFRX1 \D_cache/cache_reg[2][139]  ( .D(\D_cache/n682 ), .CK(clk), .RN(n6130), .Q(\D_cache/cache[2][139] ) );
  DFFRX1 \D_cache/cache_reg[4][58]  ( .D(\D_cache/n1328 ), .CK(clk), .RN(n6184), .Q(\D_cache/cache[4][58] ) );
  DFFRX1 \D_cache/cache_reg[6][140]  ( .D(\D_cache/n670 ), .CK(clk), .RN(n6129), .Q(\D_cache/cache[6][140] ), .QN(n3724) );
  DFFRX1 \i_MIPS/EX_MEM_reg[5]  ( .D(\i_MIPS/n399 ), .CK(clk), .RN(n6322), .Q(
        \i_MIPS/EX_MEM[5] ) );
  DFFRX1 \D_cache/cache_reg[7][139]  ( .D(\D_cache/n677 ), .CK(clk), .RN(n6130), .Q(\D_cache/cache[7][139] ) );
  DFFRX1 \D_cache/cache_reg[6][139]  ( .D(\D_cache/n678 ), .CK(clk), .RN(n6130), .Q(\D_cache/cache[6][139] ), .QN(n3756) );
  DFFRX2 \i_MIPS/ID_EX_reg[95]  ( .D(\i_MIPS/n426 ), .CK(clk), .RN(n6319), .Q(
        \i_MIPS/ID_EX[95] ) );
  DFFRX1 \D_cache/cache_reg[3][135]  ( .D(\D_cache/n713 ), .CK(clk), .RN(n6133), .Q(\D_cache/cache[3][135] ) );
  DFFRX1 \D_cache/cache_reg[2][135]  ( .D(\D_cache/n714 ), .CK(clk), .RN(n6133), .Q(\D_cache/cache[2][135] ) );
  DFFRX1 \D_cache/cache_reg[7][140]  ( .D(\D_cache/n669 ), .CK(clk), .RN(n6129), .Q(\D_cache/cache[7][140] ) );
  DFFRX1 \i_MIPS/IF_ID_reg[11]  ( .D(\i_MIPS/N28 ), .CK(clk), .RN(n6331), .Q(
        \i_MIPS/IF_ID[11] ), .QN(\i_MIPS/n164 ) );
  DFFRX1 \D_cache/cache_reg[4][18]  ( .D(\D_cache/n1648 ), .CK(clk), .RN(n6211), .Q(\D_cache/cache[4][18] ) );
  DFFRX1 \D_cache/cache_reg[4][4]  ( .D(\D_cache/n1760 ), .CK(clk), .RN(n6220), 
        .Q(\D_cache/cache[4][4] ) );
  DFFRX1 \D_cache/cache_reg[3][131]  ( .D(\D_cache/n745 ), .CK(clk), .RN(n6136), .Q(\D_cache/cache[3][131] ), .QN(n3711) );
  DFFRX1 \i_MIPS/PC/PC_o_reg[29]  ( .D(\i_MIPS/PC/n63 ), .CK(clk), .RN(n6309), 
        .Q(ICACHE_addr[27]), .QN(\i_MIPS/PC/n31 ) );
  DFFRHQX4 \i_MIPS/ID_EX_reg[77]  ( .D(\i_MIPS/n444 ), .CK(clk), .RN(n6317), 
        .Q(n3682) );
  DFFRX1 \i_MIPS/IF_ID_reg[8]  ( .D(\i_MIPS/N25 ), .CK(clk), .RN(n6330), .Q(
        \i_MIPS/IF_ID[8] ), .QN(\i_MIPS/n161 ) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[13]  ( .D(\i_MIPS/PC/n47 ), .CK(clk), .RN(n6310), 
        .Q(ICACHE_addr[11]), .QN(\i_MIPS/PC/n15 ) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[12]  ( .D(\i_MIPS/PC/n46 ), .CK(clk), .RN(n6310), 
        .Q(ICACHE_addr[10]), .QN(\i_MIPS/PC/n14 ) );
  DFFRX2 \i_MIPS/PC/PC_o_reg[10]  ( .D(\i_MIPS/PC/n44 ), .CK(clk), .RN(n6310), 
        .Q(ICACHE_addr[8]), .QN(\i_MIPS/PC/n12 ) );
  DFFRHQX4 \i_MIPS/ID_EX_reg[44]  ( .D(\i_MIPS/n361 ), .CK(clk), .RN(n6325), 
        .Q(n3558) );
  DFFRX1 \i_MIPS/IF_ID_reg[9]  ( .D(\i_MIPS/N26 ), .CK(clk), .RN(n6330), .Q(
        \i_MIPS/IF_ID[9] ), .QN(\i_MIPS/n162 ) );
  DFFRX1 \D_cache/cache_reg[0][97]  ( .D(\D_cache/n1020 ), .CK(clk), .RN(n6158), .Q(\D_cache/cache[0][97] ), .QN(n2862) );
  DFFRX1 \I_cache/cache_reg[3][141]  ( .D(n11714), .CK(clk), .RN(n6026), .Q(
        \I_cache/cache[3][141] ), .QN(n1343) );
  DFFRX1 \I_cache/cache_reg[1][141]  ( .D(n11716), .CK(clk), .RN(n6026), .Q(
        \I_cache/cache[1][141] ), .QN(n1342) );
  DFFRX1 \I_cache/cache_reg[7][141]  ( .D(n11710), .CK(clk), .RN(n6025), .Q(
        \I_cache/cache[7][141] ), .QN(n1341) );
  DFFRX1 \i_MIPS/IF_ID_reg[10]  ( .D(\i_MIPS/N27 ), .CK(clk), .RN(n6331), .Q(
        \i_MIPS/IF_ID[10] ), .QN(\i_MIPS/n163 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[7]  ( .D(\i_MIPS/N24 ), .CK(clk), .RN(n6330), .Q(
        \i_MIPS/IF_ID[7] ), .QN(\i_MIPS/n160 ) );
  DFFRX1 \i_MIPS/IF_ID_reg[5]  ( .D(\i_MIPS/N22 ), .CK(clk), .RN(n6330), .Q(
        \i_MIPS/IF_ID[5] ), .QN(\i_MIPS/n158 ) );
  DFFRX1 \i_MIPS/ID_EX_reg[84]  ( .D(\i_MIPS/n437 ), .CK(clk), .RN(n6318), .Q(
        \i_MIPS/ID_EX[84] ), .QN(n4773) );
  DFFRX4 \i_MIPS/PC/PC_o_reg[7]  ( .D(\i_MIPS/PC/n41 ), .CK(clk), .RN(n6311), 
        .Q(ICACHE_addr[5]), .QN(\i_MIPS/PC/n9 ) );
  DFFRX4 \i_MIPS/PC/PC_o_reg[15]  ( .D(\i_MIPS/PC/n49 ), .CK(clk), .RN(n6310), 
        .Q(ICACHE_addr[13]), .QN(\i_MIPS/PC/n17 ) );
  DFFRX4 \i_MIPS/PC/PC_o_reg[11]  ( .D(\i_MIPS/PC/n45 ), .CK(clk), .RN(n6310), 
        .Q(ICACHE_addr[9]), .QN(\i_MIPS/PC/n13 ) );
  DFFRX4 \i_MIPS/IF_ID_reg[46]  ( .D(\i_MIPS/N63 ), .CK(clk), .RN(n6316), .Q(
        \i_MIPS/Sign_Extend[14] ), .QN(\i_MIPS/n507 ) );
  DFFRX4 \i_MIPS/IF_ID_reg[61]  ( .D(\i_MIPS/N78 ), .CK(clk), .RN(n6320), .Q(
        \i_MIPS/IR[29] ), .QN(\i_MIPS/n253 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[47]  ( .D(\i_MIPS/N64 ), .CK(clk), .RN(n6316), .Q(
        \i_MIPS/Sign_Extend[31] ), .QN(\i_MIPS/n506 ) );
  DFFRX2 \I_cache/cache_reg[4][72]  ( .D(n12265), .CK(clk), .RN(n6071), .Q(
        \I_cache/cache[4][72] ), .QN(n1652) );
  DFFRHQX8 \i_MIPS/ID_EX_reg[73]  ( .D(\i_MIPS/n448 ), .CK(clk), .RN(n6317), 
        .Q(n11) );
  DFFRX4 \i_MIPS/IF_ID_reg[63]  ( .D(\i_MIPS/N80 ), .CK(clk), .RN(n6320), .Q(
        \i_MIPS/IR[31] ), .QN(\i_MIPS/n257 ) );
  DFFRX2 \i_MIPS/IF_ID_reg[6]  ( .D(\i_MIPS/N23 ), .CK(clk), .RN(n6330), .Q(
        \i_MIPS/IF_ID[6] ), .QN(\i_MIPS/n159 ) );
  BUFX2 U2 ( .A(net134681), .Y(net118367) );
  AND2X6 U3 ( .A(net107196), .B(n6642), .Y(n4827) );
  NAND3BX2 U4 ( .AN(n2), .B(n122), .C(n10027), .Y(\i_MIPS/N72 ) );
  NOR2X2 U5 ( .A(n10028), .B(net143858), .Y(n2) );
  NAND3BX2 U6 ( .AN(n3), .B(n123), .C(n9983), .Y(\i_MIPS/N71 ) );
  NOR2X2 U7 ( .A(n9984), .B(net143858), .Y(n3) );
  OA22X1 U8 ( .A0(n5751), .A1(n1227), .B0(n5695), .B1(n2850), .Y(n11185) );
  BUFX8 U9 ( .A(n5707), .Y(n5695) );
  INVX1 U10 ( .A(net114325), .Y(n3594) );
  NAND3X6 U11 ( .A(n3696), .B(n8399), .C(n8398), .Y(net105336) );
  AND4X4 U12 ( .A(n8392), .B(n8391), .C(n8390), .D(n8389), .Y(n3696) );
  NAND2X2 U13 ( .A(n6408), .B(n2013), .Y(n4374) );
  AOI222X1 U14 ( .A0(n5541), .A1(n11411), .B0(mem_rdata_D[35]), .B1(n131), 
        .C0(n13010), .C1(n5540), .Y(n10766) );
  NOR2X4 U15 ( .A(net143506), .B(net143507), .Y(net139864) );
  AND2X4 U16 ( .A(net118215), .B(net104964), .Y(net143506) );
  AND2X2 U17 ( .A(net118227), .B(n8595), .Y(net143507) );
  NAND2X2 U18 ( .A(net139864), .B(net105531), .Y(n4334) );
  NAND2X4 U19 ( .A(\i_MIPS/ALUin1[6] ), .B(n6707), .Y(n7301) );
  OA22X4 U20 ( .A0(n5260), .A1(n2103), .B0(n5302), .B1(n477), .Y(n6482) );
  CLKBUFX3 U21 ( .A(net104171), .Y(n3827) );
  NAND3X8 U22 ( .A(n3960), .B(n3961), .C(net109991), .Y(net104691) );
  AND4X6 U23 ( .A(n4326), .B(n4325), .C(n4323), .D(n4324), .Y(n3917) );
  NAND4X2 U24 ( .A(net115797), .B(net134815), .C(n4676), .D(n10717), .Y(n10718) );
  INVXL U25 ( .A(n6459), .Y(n3715) );
  INVX6 U26 ( .A(n10384), .Y(n10529) );
  INVX6 U27 ( .A(n10530), .Y(n10567) );
  AO22X2 U28 ( .A0(n5121), .A1(n159), .B0(n5120), .B1(n315), .Y(n8019) );
  NAND2X6 U29 ( .A(n4001), .B(n9541), .Y(n9562) );
  BUFX2 U30 ( .A(n5655), .Y(n5651) );
  BUFX8 U31 ( .A(n11091), .Y(n5573) );
  INVX16 U32 ( .A(net104168), .Y(net143857) );
  AO22X2 U33 ( .A0(n5556), .A1(n10569), .B0(n11054), .B1(n10574), .Y(n10570)
         );
  BUFX16 U34 ( .A(n11056), .Y(n5556) );
  MXI2X1 U35 ( .A(n10414), .B(n10413), .S0(n5544), .Y(n10415) );
  OR2XL U36 ( .A(n5040), .B(n10413), .Y(n3945) );
  AND2X6 U37 ( .A(net139774), .B(net106819), .Y(n3996) );
  AND2X2 U38 ( .A(net104173), .B(n11297), .Y(n3847) );
  CLKAND2X8 U39 ( .A(n9046), .B(n9045), .Y(n3701) );
  NAND3BX4 U40 ( .AN(n4), .B(n72), .C(n9682), .Y(\i_MIPS/N79 ) );
  NOR2X2 U41 ( .A(n9683), .B(net143858), .Y(n4) );
  INVX6 U42 ( .A(net110928), .Y(net112425) );
  NAND2X4 U43 ( .A(net109510), .B(n6722), .Y(n3784) );
  AND2X4 U44 ( .A(net104173), .B(net103785), .Y(n121) );
  AND2X4 U45 ( .A(net104173), .B(n11282), .Y(n4427) );
  NAND2X6 U46 ( .A(net105834), .B(net105835), .Y(n3997) );
  NAND4X2 U47 ( .A(n7323), .B(n7322), .C(n7321), .D(n7320), .Y(n7328) );
  NAND3X6 U48 ( .A(net144666), .B(net144667), .C(net107696), .Y(net104980) );
  CLKBUFX8 U49 ( .A(n9504), .Y(n5146) );
  AND3X6 U50 ( .A(n3950), .B(n7034), .C(n7029), .Y(n7054) );
  INVX4 U51 ( .A(net104868), .Y(net111763) );
  NAND2X1 U52 ( .A(n11112), .B(n3556), .Y(n5) );
  NAND2X4 U53 ( .A(n6), .B(n9439), .Y(n9540) );
  INVX3 U54 ( .A(n5), .Y(n6) );
  NAND2X2 U55 ( .A(\i_MIPS/ALUin1[29] ), .B(n134), .Y(n11112) );
  AND2X6 U56 ( .A(n9567), .B(net117743), .Y(n9570) );
  INVX3 U57 ( .A(n9432), .Y(n9438) );
  NOR4X6 U58 ( .A(n7427), .B(n7428), .C(n7426), .D(n7425), .Y(n7436) );
  AND2X4 U59 ( .A(n7406), .B(n7405), .Y(n7428) );
  NAND3X4 U60 ( .A(n3735), .B(n3736), .C(n3737), .Y(n9054) );
  NAND3X4 U61 ( .A(n11167), .B(n11166), .C(n11165), .Y(n11595) );
  CLKINVX1 U62 ( .A(net114331), .Y(n3596) );
  AND3X8 U63 ( .A(n7686), .B(n4736), .C(n7592), .Y(n7) );
  INVX20 U64 ( .A(n7), .Y(n9423) );
  NAND2X6 U65 ( .A(n3911), .B(n7431), .Y(n4007) );
  INVX6 U66 ( .A(n9542), .Y(n9441) );
  NAND2BX4 U67 ( .AN(n3670), .B(net112410), .Y(net108868) );
  NOR2X4 U68 ( .A(n3842), .B(n8), .Y(n11093) );
  OR2X8 U69 ( .A(n3765), .B(n9138), .Y(n6654) );
  AO22X2 U70 ( .A0(n5556), .A1(n10933), .B0(n11054), .B1(
        \i_MIPS/Sign_Extend[2] ), .Y(n10934) );
  NAND2X2 U71 ( .A(n10135), .B(n10903), .Y(n10156) );
  OR2X2 U72 ( .A(n10932), .B(net143858), .Y(n102) );
  AND4X6 U73 ( .A(n3635), .B(n3634), .C(n11372), .D(net118581), .Y(n3633) );
  INVX6 U74 ( .A(net104918), .Y(net108161) );
  AOI32X1 U75 ( .A0(n3669), .A1(\i_MIPS/n300 ), .A2(n3829), .B0(net108285), 
        .B1(n128), .Y(net108281) );
  AND2X2 U76 ( .A(n8715), .B(net108285), .Y(n4632) );
  INVX1 U77 ( .A(net107689), .Y(net108285) );
  NAND3X2 U78 ( .A(n13), .B(n14), .C(n9726), .Y(\i_MIPS/N54 ) );
  INVX3 U79 ( .A(n5062), .Y(n3778) );
  OAI222X2 U80 ( .A0(n7234), .A1(n9318), .B0(net107661), .B1(n7840), .C0(n9316), .C1(n7846), .Y(n7236) );
  NAND2X6 U81 ( .A(net109168), .B(net114073), .Y(n9318) );
  OAI221X1 U82 ( .A0(\i_MIPS/ALUin1[9] ), .A1(n5072), .B0(\i_MIPS/ALUin1[8] ), 
        .B1(n5068), .C0(n7144), .Y(n7234) );
  OA22X1 U83 ( .A0(\i_MIPS/ALUin1[7] ), .A1(n5064), .B0(\i_MIPS/ALUin1[6] ), 
        .B1(n3778), .Y(n7144) );
  OA22X1 U84 ( .A0(n5251), .A1(n2130), .B0(n5291), .B1(n505), .Y(n8333) );
  OR2X8 U85 ( .A(n3840), .B(n3841), .Y(n8) );
  NAND2X6 U86 ( .A(n4401), .B(n8117), .Y(n8123) );
  INVX4 U87 ( .A(net104941), .Y(net109674) );
  INVX3 U88 ( .A(n6400), .Y(n10988) );
  INVX20 U89 ( .A(n9599), .Y(n5194) );
  CLKBUFX8 U90 ( .A(n5224), .Y(n5209) );
  NOR2BX4 U91 ( .AN(n3898), .B(n3811), .Y(n4477) );
  AOI21X4 U92 ( .A0(net108297), .A1(net111570), .B0(net134145), .Y(n4273) );
  INVX6 U93 ( .A(net112219), .Y(n4276) );
  NAND2X6 U94 ( .A(net112425), .B(n7490), .Y(n6710) );
  NAND2X4 U95 ( .A(n6705), .B(\i_MIPS/ALUin1[7] ), .Y(n8117) );
  NAND2X4 U96 ( .A(n6705), .B(n2892), .Y(n8121) );
  INVX8 U97 ( .A(net104964), .Y(net108894) );
  INVX16 U98 ( .A(n5564), .Y(n5561) );
  NAND3X2 U99 ( .A(n3939), .B(n3940), .C(n10303), .Y(\i_MIPS/PC/n53 ) );
  OR2X8 U100 ( .A(n9293), .B(net117731), .Y(net144667) );
  AND2X6 U101 ( .A(n3653), .B(n9), .Y(n9608) );
  NAND2X2 U102 ( .A(n3663), .B(n11275), .Y(n9) );
  NOR2X6 U103 ( .A(n4474), .B(n4473), .Y(n3653) );
  XNOR2X4 U104 ( .A(net104691), .B(n10811), .Y(n4337) );
  NAND2X4 U105 ( .A(net139860), .B(net105195), .Y(n10811) );
  CLKMX2X2 U106 ( .A(net107656), .B(net107657), .S0(n9319), .Y(n9320) );
  OA22XL U107 ( .A0(n5919), .A1(n963), .B0(n5877), .B1(n2588), .Y(n11173) );
  NAND3X4 U108 ( .A(\i_MIPS/PC/n6 ), .B(ICACHE_addr[3]), .C(\i_MIPS/PC/n8 ), 
        .Y(n4678) );
  BUFX12 U109 ( .A(n5935), .Y(n5943) );
  CLKAND2X2 U110 ( .A(n3663), .B(n11266), .Y(n3846) );
  INVX4 U111 ( .A(net105336), .Y(net109202) );
  OR2X4 U112 ( .A(net112329), .B(net117733), .Y(n3814) );
  AND4X6 U113 ( .A(n4056), .B(n4057), .C(n4055), .D(n4054), .Y(n3999) );
  OAI21X1 U114 ( .A0(n6815), .A1(n7027), .B0(n8696), .Y(n6727) );
  NOR3X4 U115 ( .A(n4453), .B(n4452), .C(n4454), .Y(n10230) );
  CLKAND2X2 U116 ( .A(n3663), .B(n11263), .Y(n4453) );
  AND3X6 U117 ( .A(net108623), .B(n8782), .C(n9218), .Y(n3848) );
  INVX4 U118 ( .A(n10619), .Y(n9293) );
  NAND3X2 U119 ( .A(n4419), .B(n4420), .C(n10534), .Y(\i_MIPS/PC/n62 ) );
  CLKAND2X2 U120 ( .A(net104172), .B(n11265), .Y(n4435) );
  INVX6 U121 ( .A(n6818), .Y(n6819) );
  CLKAND2X2 U122 ( .A(net104173), .B(n11296), .Y(n4436) );
  AOI222X1 U123 ( .A0(net104171), .A1(n11241), .B0(net104172), .B1(n11272), 
        .C0(net104173), .C1(n11303), .Y(n10027) );
  CLKMX2X3 U124 ( .A(n3609), .B(net134375), .S0(net143514), .Y(n6703) );
  CLKINVX4 U125 ( .A(n7048), .Y(n7029) );
  CLKINVX6 U126 ( .A(n10376), .Y(n10385) );
  CLKINVX4 U127 ( .A(n10272), .Y(n10282) );
  INVX4 U128 ( .A(n9562), .Y(n9565) );
  NAND4X1 U129 ( .A(n3950), .B(n9562), .C(n9563), .D(n9543), .Y(n9574) );
  AOI222X1 U130 ( .A0(net104171), .A1(n11240), .B0(n3663), .B1(n11271), .C0(
        net104173), .C1(n11302), .Y(n9983) );
  CLKINVX6 U131 ( .A(net105234), .Y(net109528) );
  OA22X4 U132 ( .A0(n2928), .A1(n5064), .B0(\i_MIPS/n297 ), .B1(n5059), .Y(
        n6671) );
  INVX6 U133 ( .A(n4007), .Y(n7433) );
  CLKAND2X3 U134 ( .A(n6707), .B(n1302), .Y(n3753) );
  INVX6 U135 ( .A(n6707), .Y(n6711) );
  NAND3X2 U136 ( .A(n4413), .B(n4414), .C(n10494), .Y(\i_MIPS/PC/n48 ) );
  AOI2BB1X1 U137 ( .A0N(\i_MIPS/PC/n16 ), .A1N(net115799), .B0(n10493), .Y(
        n10494) );
  INVX20 U138 ( .A(n5559), .Y(n5558) );
  OA22X2 U139 ( .A0(n5331), .A1(n625), .B0(n5356), .B1(n2243), .Y(n8830) );
  INVX12 U140 ( .A(net106822), .Y(n3648) );
  INVX12 U141 ( .A(net104828), .Y(net106822) );
  NOR3X4 U142 ( .A(n4488), .B(n4487), .C(n4489), .Y(n10049) );
  CLKAND2X2 U143 ( .A(n3898), .B(n11305), .Y(n4489) );
  CLKAND2X2 U144 ( .A(net104172), .B(n11274), .Y(n4488) );
  CLKAND2X3 U145 ( .A(n3663), .B(n11268), .Y(n3841) );
  INVX16 U146 ( .A(n3921), .Y(n3663) );
  INVX1 U147 ( .A(n8961), .Y(n8965) );
  CLKAND2X2 U148 ( .A(n3898), .B(n11293), .Y(n4481) );
  OA22X4 U149 ( .A0(n1264), .A1(n5063), .B0(n2921), .B1(n5057), .Y(n7954) );
  OR2X1 U150 ( .A(n9734), .B(n5557), .Y(n4424) );
  INVX20 U151 ( .A(n5559), .Y(n5557) );
  OA22X2 U152 ( .A0(n5330), .A1(n1255), .B0(n5359), .B1(n2875), .Y(n8422) );
  NAND2X8 U153 ( .A(n8780), .B(n8779), .Y(n9224) );
  INVX6 U154 ( .A(n6483), .Y(n11029) );
  CLKBUFX6 U155 ( .A(n11050), .Y(n5551) );
  NOR3X4 U156 ( .A(n4430), .B(n4429), .C(n4428), .Y(n10866) );
  CLKAND2X2 U157 ( .A(n3898), .B(n11285), .Y(n4430) );
  INVX3 U158 ( .A(n8298), .Y(n8292) );
  OA22X4 U159 ( .A0(n2919), .A1(n5064), .B0(n336), .B1(n5058), .Y(n7105) );
  INVX4 U160 ( .A(n6768), .Y(n6770) );
  AND2X6 U161 ( .A(n6770), .B(n6776), .Y(net134685) );
  INVX12 U162 ( .A(n3788), .Y(n3789) );
  NOR2X2 U163 ( .A(n5335), .B(n3889), .Y(n3887) );
  INVX3 U164 ( .A(n3834), .Y(n6518) );
  CLKAND2X3 U165 ( .A(n3898), .B(n11294), .Y(n4454) );
  AOI2BB1X1 U166 ( .A0N(\i_MIPS/PC/n17 ), .A1N(net115789), .B0(n10266), .Y(
        n10267) );
  CLKMX2X4 U167 ( .A(n7940), .B(n7939), .S0(net114087), .Y(net110147) );
  CLKMX2X2 U168 ( .A(n7524), .B(n7523), .S0(net114087), .Y(n7525) );
  MXI2X1 U169 ( .A(n7987), .B(n7986), .S0(net114087), .Y(n3981) );
  MX2X6 U170 ( .A(n9164), .B(n9163), .S0(net114085), .Y(net107943) );
  MXI2X1 U171 ( .A(n9345), .B(n9344), .S0(net114085), .Y(n3719) );
  MXI2X1 U172 ( .A(n7184), .B(n7183), .S0(net114085), .Y(n3891) );
  AND4X4 U173 ( .A(n6767), .B(n6766), .C(n6765), .D(n6764), .Y(net134445) );
  INVX4 U174 ( .A(n7962), .Y(n7960) );
  CLKBUFX2 U175 ( .A(n8969), .Y(n10) );
  INVXL U176 ( .A(n3831), .Y(n3833) );
  BUFX8 U177 ( .A(n10590), .Y(n140) );
  NAND2X6 U178 ( .A(n3974), .B(n4278), .Y(n4277) );
  OR3X8 U179 ( .A(n3692), .B(n3693), .C(n3694), .Y(net105071) );
  INVX3 U180 ( .A(n8862), .Y(n8966) );
  NAND2X4 U181 ( .A(n4789), .B(n4786), .Y(n7888) );
  CLKBUFX3 U182 ( .A(n9502), .Y(n5132) );
  NOR4X2 U183 ( .A(n8443), .B(n8442), .C(n8441), .D(n8440), .Y(n8444) );
  NAND2X6 U184 ( .A(net139862), .B(net105756), .Y(n4341) );
  AND3X8 U185 ( .A(\i_MIPS/ID_EX[76] ), .B(\i_MIPS/ALUOp[1] ), .C(n3622), .Y(
        n6645) );
  OAI2BB2X4 U186 ( .B0(n6964), .B1(n9425), .A0N(n6931), .A1N(n4682), .Y(n6944)
         );
  NAND3X8 U187 ( .A(n9572), .B(n148), .C(n3689), .Y(n10711) );
  AND2X2 U188 ( .A(net117743), .B(n9540), .Y(n3872) );
  INVX1 U189 ( .A(net108300), .Y(net108299) );
  BUFX20 U190 ( .A(n8466), .Y(n4883) );
  INVX6 U191 ( .A(n8974), .Y(n8969) );
  CLKINVX6 U192 ( .A(n11), .Y(n12) );
  NAND4BX2 U193 ( .AN(n4645), .B(n9179), .C(n9178), .D(n9177), .Y(n11411) );
  OA22X4 U194 ( .A0(n2949), .A1(n5063), .B0(n345), .B1(n5057), .Y(n7944) );
  NAND3BX4 U195 ( .AN(n3707), .B(n3910), .C(n8209), .Y(n8214) );
  INVX3 U196 ( .A(net107661), .Y(net109661) );
  NAND2X6 U197 ( .A(net139765), .B(net105783), .Y(n4354) );
  AND2X1 U198 ( .A(n5065), .B(n3670), .Y(n4730) );
  MXI2X2 U199 ( .A(n7221), .B(n7231), .S0(net114065), .Y(n4653) );
  OAI211X1 U200 ( .A0(\i_MIPS/ALUin1[16] ), .A1(n5068), .B0(n7158), .C0(n7157), 
        .Y(n7231) );
  NOR2X8 U201 ( .A(net108641), .B(net117731), .Y(n3695) );
  INVX6 U202 ( .A(net104794), .Y(net108641) );
  NAND2X6 U203 ( .A(n3632), .B(n8779), .Y(n8566) );
  OAI2BB1X2 U204 ( .A0N(n4709), .A1N(n7028), .B0(n7862), .Y(n7048) );
  NAND2X8 U205 ( .A(n3710), .B(n4732), .Y(n7028) );
  NAND2X6 U206 ( .A(\i_MIPS/ALUin1[11] ), .B(n6695), .Y(n8464) );
  NAND2X6 U207 ( .A(\i_MIPS/ALUin1[10] ), .B(n6691), .Y(n8467) );
  CLKINVX6 U208 ( .A(n6703), .Y(n6691) );
  INVX3 U209 ( .A(n11485), .Y(n10799) );
  CLKMX2X8 U210 ( .A(n3609), .B(net134375), .S0(net143514), .Y(n3760) );
  OAI221X2 U211 ( .A0(n10824), .A1(net143858), .B0(\i_MIPS/n521 ), .B1(
        net115793), .C0(n10823), .Y(\i_MIPS/N49 ) );
  MX2X8 U212 ( .A(\i_MIPS/n214 ), .B(n4791), .S0(net143514), .Y(net112410) );
  BUFX20 U213 ( .A(n5223), .Y(n5211) );
  OAI221X1 U214 ( .A0(n5186), .A1(n1332), .B0(n5211), .B1(n2985), .C0(n6419), 
        .Y(n6420) );
  BUFX4 U215 ( .A(n10510), .Y(n4514) );
  NAND3X2 U216 ( .A(n7694), .B(n7693), .C(n3950), .Y(n3582) );
  INVX8 U217 ( .A(n7694), .Y(n7695) );
  MXI2X4 U218 ( .A(\i_MIPS/ID_EX[47] ), .B(n5050), .S0(net143514), .Y(n6707)
         );
  MX2X6 U219 ( .A(\i_MIPS/n228 ), .B(n3903), .S0(net143514), .Y(n6704) );
  AND4X6 U220 ( .A(n3581), .B(n3582), .C(n3030), .D(n3580), .Y(n7700) );
  INVX1 U221 ( .A(net107119), .Y(n4314) );
  NAND2X2 U222 ( .A(n4738), .B(net107119), .Y(n11073) );
  CLKBUFX6 U223 ( .A(n11209), .Y(n5788) );
  NAND3BX4 U224 ( .AN(\i_MIPS/PC/n6 ), .B(ICACHE_addr[4]), .C(\i_MIPS/PC/n7 ), 
        .Y(n11209) );
  MXI2X2 U225 ( .A(n10451), .B(n10450), .S0(n5545), .Y(n10452) );
  CLKINVX3 U226 ( .A(n9957), .Y(n9959) );
  NOR2X6 U227 ( .A(n3658), .B(n9957), .Y(n4737) );
  INVX12 U228 ( .A(n5194), .Y(n5026) );
  INVX8 U229 ( .A(n5194), .Y(n4626) );
  OR2X2 U230 ( .A(n9727), .B(net143858), .Y(n13) );
  OR2X1 U231 ( .A(\i_MIPS/n516 ), .B(net115789), .Y(n14) );
  INVX3 U232 ( .A(n11317), .Y(n9727) );
  OR2X2 U233 ( .A(n10074), .B(net143858), .Y(n15) );
  OR2X2 U234 ( .A(\i_MIPS/n506 ), .B(net115793), .Y(n16) );
  NAND3X4 U235 ( .A(n15), .B(n16), .C(n10073), .Y(\i_MIPS/N64 ) );
  NOR3X4 U236 ( .A(n4435), .B(n4434), .C(n4436), .Y(n10073) );
  AND2X2 U237 ( .A(mem_rdata_I[32]), .B(n5945), .Y(n17) );
  CLKAND2X4 U238 ( .A(n5566), .B(n11250), .Y(n18) );
  OR2X6 U239 ( .A(n17), .B(n18), .Y(n6552) );
  BUFX6 U240 ( .A(n5936), .Y(n5945) );
  CLKMX2X2 U241 ( .A(\I_cache/cache[0][64] ), .B(n6552), .S0(n5625), .Y(n12333) );
  MX2X1 U242 ( .A(\I_cache/cache[1][64] ), .B(n6552), .S0(n5576), .Y(n12332)
         );
  MX2X1 U243 ( .A(\I_cache/cache[2][64] ), .B(n6552), .S0(n5716), .Y(n12331)
         );
  MX2X1 U244 ( .A(\I_cache/cache[3][64] ), .B(n6552), .S0(n5671), .Y(n12330)
         );
  MX2X1 U245 ( .A(\I_cache/cache[4][64] ), .B(n6552), .S0(n5806), .Y(n12329)
         );
  MX2X1 U246 ( .A(\I_cache/cache[5][64] ), .B(n6552), .S0(n5755), .Y(n12328)
         );
  MX2X1 U247 ( .A(\I_cache/cache[6][64] ), .B(n6552), .S0(n5893), .Y(n12327)
         );
  MX2X1 U248 ( .A(\I_cache/cache[7][64] ), .B(n6552), .S0(n5848), .Y(n12326)
         );
  AND2X2 U249 ( .A(net104171), .B(n11237), .Y(n3840) );
  NAND3X4 U250 ( .A(n3838), .B(n3839), .C(n11093), .Y(\i_MIPS/N68 ) );
  AND2X2 U251 ( .A(mem_rdata_I[53]), .B(n5944), .Y(n19) );
  CLKAND2X4 U252 ( .A(n5567), .B(n11270), .Y(n20) );
  OR2X6 U253 ( .A(n19), .B(n20), .Y(n9989) );
  CLKMX2X2 U254 ( .A(\I_cache/cache[0][85] ), .B(n9989), .S0(n5622), .Y(n12165) );
  MX2X1 U255 ( .A(\I_cache/cache[1][85] ), .B(n9989), .S0(n5579), .Y(n12164)
         );
  MX2X1 U256 ( .A(\I_cache/cache[2][85] ), .B(n9989), .S0(n5713), .Y(n12163)
         );
  MX2X1 U257 ( .A(\I_cache/cache[3][85] ), .B(n9989), .S0(n5668), .Y(n12162)
         );
  MX2X1 U258 ( .A(\I_cache/cache[4][85] ), .B(n9989), .S0(n5803), .Y(n12161)
         );
  MX2X1 U259 ( .A(\I_cache/cache[5][85] ), .B(n9989), .S0(n5757), .Y(n12160)
         );
  MX2X1 U260 ( .A(\I_cache/cache[6][85] ), .B(n9989), .S0(n5890), .Y(n12159)
         );
  MX2X1 U261 ( .A(\I_cache/cache[7][85] ), .B(n9989), .S0(n5847), .Y(n12158)
         );
  CLKAND2X3 U262 ( .A(mem_rdata_I[56]), .B(n5945), .Y(n21) );
  AND2X4 U263 ( .A(n5566), .B(n11273), .Y(n22) );
  OR2X8 U264 ( .A(n21), .B(n22), .Y(n6547) );
  NAND4X4 U265 ( .A(n6546), .B(n6545), .C(n6544), .D(n6543), .Y(n11273) );
  MX2X1 U266 ( .A(\I_cache/cache[0][88] ), .B(n6547), .S0(n5620), .Y(n12141)
         );
  MX2X1 U267 ( .A(\I_cache/cache[2][88] ), .B(n6547), .S0(n5716), .Y(n12139)
         );
  MX2X1 U268 ( .A(\I_cache/cache[3][88] ), .B(n6547), .S0(n5671), .Y(n12138)
         );
  MX2X1 U269 ( .A(\I_cache/cache[4][88] ), .B(n6547), .S0(n5806), .Y(n12137)
         );
  MX2X1 U270 ( .A(\I_cache/cache[5][88] ), .B(n6547), .S0(n5754), .Y(n12136)
         );
  MX2X1 U271 ( .A(\I_cache/cache[6][88] ), .B(n6547), .S0(n5893), .Y(n12135)
         );
  MX2X1 U272 ( .A(\I_cache/cache[7][88] ), .B(n6547), .S0(n5848), .Y(n12134)
         );
  CLKAND2X3 U273 ( .A(n4505), .B(n11458), .Y(n23) );
  AND2X2 U274 ( .A(mem_rdata_D[82]), .B(n133), .Y(n24) );
  AND2X2 U275 ( .A(n12995), .B(n5536), .Y(n25) );
  NOR3X4 U276 ( .A(n23), .B(n24), .C(n25), .Y(n10638) );
  BUFX6 U277 ( .A(n4686), .Y(n5536) );
  NAND2X1 U278 ( .A(\D_cache/cache[0][41] ), .B(n26), .Y(n27) );
  NAND2X1 U279 ( .A(n4569), .B(n5164), .Y(n28) );
  NAND2X1 U280 ( .A(n27), .B(n28), .Y(\D_cache/n1468 ) );
  INVXL U281 ( .A(n5164), .Y(n26) );
  BUFX8 U282 ( .A(n10611), .Y(n4569) );
  INVX4 U283 ( .A(n5176), .Y(n5164) );
  AND2X2 U284 ( .A(mem_rdata_I[50]), .B(n5942), .Y(n29) );
  AND2X4 U285 ( .A(n5567), .B(net103817), .Y(n30) );
  OR2X8 U286 ( .A(n29), .B(n30), .Y(n9770) );
  NAND4X4 U287 ( .A(net106718), .B(net106719), .C(net106720), .D(net106721), 
        .Y(net103817) );
  MX2X1 U288 ( .A(\I_cache/cache[0][82] ), .B(n9770), .S0(n5618), .Y(n12189)
         );
  MX2X1 U289 ( .A(\I_cache/cache[1][82] ), .B(n9770), .S0(n5581), .Y(n12188)
         );
  MX2X1 U290 ( .A(\I_cache/cache[3][82] ), .B(n9770), .S0(n5664), .Y(n12186)
         );
  MX2X1 U291 ( .A(\I_cache/cache[4][82] ), .B(n9770), .S0(n5799), .Y(n12185)
         );
  MX2X1 U292 ( .A(\I_cache/cache[6][82] ), .B(n9770), .S0(n5886), .Y(n12183)
         );
  MX2X1 U293 ( .A(\I_cache/cache[7][82] ), .B(n9770), .S0(n5843), .Y(n12182)
         );
  AND2X2 U294 ( .A(mem_rdata_I[34]), .B(n5944), .Y(n31) );
  AND2X4 U295 ( .A(n5566), .B(n11252), .Y(n32) );
  OR2X8 U296 ( .A(n31), .B(n32), .Y(n10915) );
  NAND4X4 U297 ( .A(n6533), .B(n6532), .C(n6531), .D(n6530), .Y(n11252) );
  MX2X1 U298 ( .A(\I_cache/cache[0][66] ), .B(n10915), .S0(n5623), .Y(n12317)
         );
  MX2X1 U299 ( .A(\I_cache/cache[1][66] ), .B(n10915), .S0(n5576), .Y(n12316)
         );
  MX2X1 U300 ( .A(\I_cache/cache[2][66] ), .B(n10915), .S0(n5712), .Y(n12315)
         );
  MX2X1 U301 ( .A(\I_cache/cache[3][66] ), .B(n10915), .S0(n5668), .Y(n12314)
         );
  MX2X1 U302 ( .A(\I_cache/cache[4][66] ), .B(n10915), .S0(n5798), .Y(n12313)
         );
  MX2X1 U303 ( .A(\I_cache/cache[5][66] ), .B(n10915), .S0(n4831), .Y(n12312)
         );
  MX2X1 U304 ( .A(\I_cache/cache[6][66] ), .B(n10915), .S0(n5890), .Y(n12311)
         );
  CLKAND2X2 U305 ( .A(n4505), .B(n11464), .Y(n33) );
  AND2X2 U306 ( .A(mem_rdata_D[88]), .B(n129), .Y(n34) );
  CLKAND2X3 U307 ( .A(n12989), .B(n5535), .Y(n35) );
  NOR3X2 U308 ( .A(n33), .B(n34), .C(n35), .Y(n10421) );
  NAND4X8 U309 ( .A(n6742), .B(n6741), .C(n6740), .D(n6739), .Y(n11464) );
  BUFX8 U310 ( .A(n4686), .Y(n5535) );
  NAND2X2 U311 ( .A(mem_rdata_I[33]), .B(n5945), .Y(n36) );
  NAND2X2 U312 ( .A(n5566), .B(n11251), .Y(n37) );
  NAND2X8 U313 ( .A(n36), .B(n37), .Y(n10873) );
  NAND4X4 U314 ( .A(n6537), .B(n6536), .C(n6535), .D(n6534), .Y(n11251) );
  MX2X1 U315 ( .A(\I_cache/cache[0][65] ), .B(n10873), .S0(n5619), .Y(n12325)
         );
  MX2X1 U316 ( .A(\I_cache/cache[1][65] ), .B(n10873), .S0(n5580), .Y(n12324)
         );
  MX2X1 U317 ( .A(\I_cache/cache[2][65] ), .B(n10873), .S0(n5716), .Y(n12323)
         );
  MX2X1 U318 ( .A(\I_cache/cache[4][65] ), .B(n10873), .S0(n5806), .Y(n12321)
         );
  MX2X1 U319 ( .A(\I_cache/cache[5][65] ), .B(n10873), .S0(n5759), .Y(n12320)
         );
  MX2X1 U320 ( .A(\I_cache/cache[6][65] ), .B(n10873), .S0(n5893), .Y(n12319)
         );
  CLKAND2X2 U321 ( .A(n4505), .B(n11471), .Y(n38) );
  AND2X2 U322 ( .A(mem_rdata_D[95]), .B(n130), .Y(n39) );
  CLKAND2X3 U323 ( .A(n12982), .B(n5536), .Y(n40) );
  NOR3X2 U324 ( .A(n38), .B(n39), .C(n40), .Y(n10703) );
  NAND4X6 U325 ( .A(n9524), .B(n9523), .C(n9522), .D(n9521), .Y(n11471) );
  CLKAND2X2 U326 ( .A(n4505), .B(n11440), .Y(n41) );
  AND2X2 U327 ( .A(mem_rdata_D[64]), .B(n129), .Y(n42) );
  CLKAND2X3 U328 ( .A(n13013), .B(n5535), .Y(n43) );
  NOR3X2 U329 ( .A(n41), .B(n42), .C(n43), .Y(n10742) );
  NAND4X6 U330 ( .A(n8748), .B(n8747), .C(n8746), .D(n8745), .Y(n11440) );
  NAND2X1 U331 ( .A(mem_rdata_I[48]), .B(n5942), .Y(n44) );
  NAND2X2 U332 ( .A(n5567), .B(n11266), .Y(n45) );
  NAND2X8 U333 ( .A(n44), .B(n45), .Y(n9752) );
  BUFX8 U334 ( .A(n5934), .Y(n5942) );
  NAND4X4 U335 ( .A(n9751), .B(n9750), .C(n9749), .D(n9748), .Y(n11266) );
  MX2X1 U336 ( .A(\I_cache/cache[1][80] ), .B(n9752), .S0(n5577), .Y(n12204)
         );
  MX2X1 U337 ( .A(\I_cache/cache[3][80] ), .B(n9752), .S0(n5663), .Y(n12202)
         );
  MX2X1 U338 ( .A(\I_cache/cache[4][80] ), .B(n9752), .S0(n5798), .Y(n12201)
         );
  MX2X1 U339 ( .A(\I_cache/cache[5][80] ), .B(n9752), .S0(n5755), .Y(n12200)
         );
  MX2X1 U340 ( .A(\I_cache/cache[6][80] ), .B(n9752), .S0(n5885), .Y(n12199)
         );
  MX2X1 U341 ( .A(\I_cache/cache[7][80] ), .B(n9752), .S0(n5842), .Y(n12198)
         );
  MX2X1 U342 ( .A(\I_cache/cache[0][80] ), .B(n9752), .S0(n5618), .Y(n12205)
         );
  NAND2X6 U343 ( .A(net104830), .B(net106822), .Y(n46) );
  CLKINVX4 U344 ( .A(n9729), .Y(n47) );
  NAND2X8 U345 ( .A(n46), .B(n47), .Y(n11059) );
  CLKINVX6 U346 ( .A(net106828), .Y(net104830) );
  NAND2X2 U347 ( .A(n12963), .B(mem_read_D), .Y(n48) );
  NAND2X2 U348 ( .A(mem_write_D), .B(n11524), .Y(n49) );
  NAND2X1 U349 ( .A(n48), .B(n49), .Y(n5010) );
  BUFX20 U350 ( .A(n11534), .Y(mem_read_D) );
  INVX20 U351 ( .A(n5040), .Y(mem_write_D) );
  NAND2XL U352 ( .A(n9952), .B(n9951), .Y(n50) );
  INVX1 U353 ( .A(n9950), .Y(n51) );
  NAND2X2 U354 ( .A(n50), .B(n51), .Y(n9958) );
  NAND2X2 U355 ( .A(DCACHE_addr[0]), .B(DCACHE_addr[1]), .Y(n9951) );
  NAND3X4 U356 ( .A(n9956), .B(n9959), .C(n9958), .Y(n10973) );
  OR2X2 U357 ( .A(n9631), .B(net143858), .Y(n52) );
  OR2X1 U358 ( .A(\i_MIPS/n249 ), .B(net115789), .Y(n53) );
  NAND3X4 U359 ( .A(n52), .B(n53), .C(n9630), .Y(\i_MIPS/N76 ) );
  OR2X2 U360 ( .A(n10961), .B(net143858), .Y(n54) );
  OR2X1 U361 ( .A(\i_MIPS/n518 ), .B(net115789), .Y(n55) );
  NAND3X4 U362 ( .A(n54), .B(n55), .C(n10960), .Y(\i_MIPS/N52 ) );
  AND2X4 U363 ( .A(n4506), .B(n11459), .Y(n56) );
  AND2X2 U364 ( .A(mem_rdata_D[83]), .B(n133), .Y(n57) );
  AND2X2 U365 ( .A(n5535), .B(n12994), .Y(n58) );
  NOR3X2 U366 ( .A(n56), .B(n57), .C(n58), .Y(n10968) );
  INVX16 U367 ( .A(n4504), .Y(n4506) );
  OR2X2 U368 ( .A(n9653), .B(net143858), .Y(n59) );
  OR2X1 U369 ( .A(\i_MIPS/n251 ), .B(net115789), .Y(n60) );
  NAND3X4 U370 ( .A(n59), .B(n60), .C(n9652), .Y(\i_MIPS/N77 ) );
  NAND2X1 U371 ( .A(\D_cache/cache[6][45] ), .B(n61), .Y(n62) );
  NAND2X1 U372 ( .A(n4538), .B(n3574), .Y(n63) );
  NAND2X1 U373 ( .A(n62), .B(n63), .Y(\D_cache/n1430 ) );
  INVXL U374 ( .A(n3574), .Y(n61) );
  BUFX8 U375 ( .A(n10804), .Y(n4538) );
  INVX4 U376 ( .A(n5381), .Y(n3574) );
  CLKAND2X2 U377 ( .A(n4506), .B(n11465), .Y(n64) );
  AND2X2 U378 ( .A(mem_rdata_D[89]), .B(n130), .Y(n65) );
  AND2X4 U379 ( .A(n12988), .B(n5535), .Y(n66) );
  NOR3X4 U380 ( .A(n64), .B(n65), .C(n66), .Y(n10435) );
  NAND4X6 U381 ( .A(n6861), .B(n6860), .C(n6859), .D(n6858), .Y(n11465) );
  MXI2X4 U382 ( .A(n10435), .B(n10434), .S0(n5544), .Y(n10436) );
  AND2X1 U383 ( .A(net104171), .B(n11236), .Y(n67) );
  CLKAND2X2 U384 ( .A(n3663), .B(n11267), .Y(n68) );
  CLKAND2X2 U385 ( .A(net104173), .B(n11298), .Y(n69) );
  NOR3X4 U386 ( .A(n67), .B(n68), .C(n69), .Y(n9746) );
  NAND4X4 U387 ( .A(n9739), .B(n9738), .C(n9737), .D(n9736), .Y(n11236) );
  OR2X2 U388 ( .A(n10133), .B(net143858), .Y(n70) );
  OR2X1 U389 ( .A(\i_MIPS/n509 ), .B(net115793), .Y(n71) );
  NAND3X2 U390 ( .A(n70), .B(n71), .C(n10132), .Y(\i_MIPS/N61 ) );
  CLKBUFX3 U391 ( .A(net115813), .Y(net115793) );
  OR2X1 U392 ( .A(\i_MIPS/n255 ), .B(net115789), .Y(n72) );
  CLKAND2X4 U393 ( .A(n4505), .B(n11444), .Y(n73) );
  AND2X2 U394 ( .A(mem_rdata_D[68]), .B(n131), .Y(n74) );
  AND2X1 U395 ( .A(n13009), .B(n5535), .Y(n75) );
  NOR3X4 U396 ( .A(n73), .B(n74), .C(n75), .Y(n10751) );
  NAND4X4 U397 ( .A(n9087), .B(n9086), .C(n9085), .D(n9084), .Y(n11444) );
  NAND2X1 U398 ( .A(n3560), .B(n3950), .Y(n76) );
  NAND2X1 U399 ( .A(n77), .B(n4764), .Y(n8794) );
  CLKINVX1 U400 ( .A(n76), .Y(n77) );
  OR2X1 U401 ( .A(\i_MIPS/Register/register[2][0] ), .B(n5091), .Y(n78) );
  OR2X1 U402 ( .A(\i_MIPS/Register/register[10][0] ), .B(n5087), .Y(n79) );
  NAND3X1 U403 ( .A(n78), .B(n79), .C(n8759), .Y(n8767) );
  NAND4BX2 U404 ( .AN(n8767), .B(n8766), .C(n8765), .D(n8764), .Y(n8778) );
  OR2X2 U405 ( .A(n10285), .B(n5561), .Y(n80) );
  OR2X2 U406 ( .A(n5558), .B(n10286), .Y(n81) );
  NAND3X1 U407 ( .A(n80), .B(n81), .C(n10284), .Y(\i_MIPS/PC/n51 ) );
  OR2X2 U408 ( .A(n9705), .B(net143858), .Y(n82) );
  OR2X2 U409 ( .A(\i_MIPS/n253 ), .B(net115789), .Y(n83) );
  NAND3X6 U410 ( .A(n82), .B(n83), .C(n9704), .Y(\i_MIPS/N78 ) );
  INVX3 U411 ( .A(n11340), .Y(n9705) );
  NOR3X6 U412 ( .A(n4458), .B(n4459), .C(n4460), .Y(n9704) );
  OR2X2 U413 ( .A(n9912), .B(net143858), .Y(n84) );
  OR2X2 U414 ( .A(\i_MIPS/n514 ), .B(net115791), .Y(n85) );
  NAND3X6 U415 ( .A(n84), .B(n85), .C(n9911), .Y(\i_MIPS/N56 ) );
  INVX1 U416 ( .A(n11319), .Y(n9912) );
  NAND2X1 U417 ( .A(n8034), .B(net118584), .Y(n86) );
  NAND2X2 U418 ( .A(n8033), .B(n8032), .Y(n87) );
  NAND2X2 U419 ( .A(n8031), .B(n8030), .Y(n88) );
  AND3X6 U420 ( .A(n86), .B(n87), .C(n88), .Y(n8049) );
  CLKBUFX4 U421 ( .A(net107404), .Y(net118584) );
  OR3X2 U422 ( .A(n3779), .B(n3780), .C(n3781), .Y(n8032) );
  AO22X1 U423 ( .A0(n8028), .A1(net117747), .B0(n3950), .B1(n8027), .Y(n8031)
         );
  NAND2X1 U424 ( .A(n8044), .B(n8029), .Y(n8030) );
  NAND4X6 U425 ( .A(n8049), .B(n8048), .C(n8047), .D(n8046), .Y(net105010) );
  OR2X6 U426 ( .A(net110640), .B(net117711), .Y(n89) );
  OR2X4 U427 ( .A(n4090), .B(net117731), .Y(n90) );
  NAND3X6 U428 ( .A(n89), .B(n90), .C(net110642), .Y(net105093) );
  BUFX16 U429 ( .A(net105093), .Y(n3706) );
  NAND2X4 U430 ( .A(n10763), .B(n91), .Y(n92) );
  NAND2X1 U431 ( .A(n10762), .B(n5550), .Y(n93) );
  NAND2X2 U432 ( .A(n92), .B(n93), .Y(n94) );
  INVX3 U433 ( .A(n5550), .Y(n91) );
  INVX3 U434 ( .A(n94), .Y(n10764) );
  INVX3 U435 ( .A(n11379), .Y(n10762) );
  BUFX4 U436 ( .A(n10974), .Y(n5550) );
  BUFX4 U437 ( .A(n10764), .Y(n4499) );
  OR2X2 U438 ( .A(n10253), .B(net143858), .Y(n95) );
  OR2X2 U439 ( .A(\i_MIPS/n507 ), .B(net115791), .Y(n96) );
  NAND3X6 U440 ( .A(n95), .B(n96), .C(n10252), .Y(\i_MIPS/N63 ) );
  INVX3 U441 ( .A(n11326), .Y(n10253) );
  AND2X2 U442 ( .A(mem_rdata_I[47]), .B(n5940), .Y(n97) );
  AND2X2 U443 ( .A(n5568), .B(n11265), .Y(n98) );
  OR2X6 U444 ( .A(n97), .B(n98), .Y(n10057) );
  CLKBUFX6 U445 ( .A(n5565), .Y(n5568) );
  CLKMX2X2 U446 ( .A(\I_cache/cache[0][79] ), .B(n10057), .S0(n5619), .Y(
        n12213) );
  MX2X1 U447 ( .A(\I_cache/cache[1][79] ), .B(n10057), .S0(n5576), .Y(n12212)
         );
  MX2X1 U448 ( .A(\I_cache/cache[2][79] ), .B(n10057), .S0(n5710), .Y(n12211)
         );
  MX2X1 U449 ( .A(\I_cache/cache[3][79] ), .B(n10057), .S0(n5665), .Y(n12210)
         );
  MX2X1 U450 ( .A(\I_cache/cache[4][79] ), .B(n10057), .S0(n5800), .Y(n12209)
         );
  MX2X1 U451 ( .A(\I_cache/cache[5][79] ), .B(n10057), .S0(n5754), .Y(n12208)
         );
  MX2X1 U452 ( .A(\I_cache/cache[6][79] ), .B(n10057), .S0(n5888), .Y(n12207)
         );
  MX2X1 U453 ( .A(\I_cache/cache[7][79] ), .B(n10057), .S0(n5844), .Y(n12206)
         );
  CLKAND2X2 U454 ( .A(n3800), .B(n11386), .Y(n99) );
  AND2X4 U455 ( .A(mem_rdata_D[10]), .B(n130), .Y(n100) );
  AND2X2 U456 ( .A(n13003), .B(n5538), .Y(n101) );
  NOR3X4 U457 ( .A(n99), .B(n100), .C(n101), .Y(n10778) );
  NAND4X4 U458 ( .A(n7537), .B(n7536), .C(n7535), .D(n7534), .Y(n11386) );
  MXI2X4 U459 ( .A(n10778), .B(n10777), .S0(n5550), .Y(n10779) );
  OR2X1 U460 ( .A(\i_MIPS/n519 ), .B(net115791), .Y(n103) );
  NAND3X2 U461 ( .A(n102), .B(n103), .C(n10931), .Y(\i_MIPS/N51 ) );
  OR2X1 U462 ( .A(n10171), .B(n5561), .Y(n104) );
  OR2X2 U463 ( .A(n5557), .B(n10172), .Y(n105) );
  NAND3X2 U464 ( .A(n104), .B(n105), .C(n10170), .Y(\i_MIPS/PC/n44 ) );
  OR2XL U465 ( .A(n10182), .B(n5561), .Y(n106) );
  OR2XL U466 ( .A(n5558), .B(n10183), .Y(n107) );
  NAND3X2 U467 ( .A(n106), .B(n107), .C(n10181), .Y(\i_MIPS/PC/n45 ) );
  AOI2BB1X4 U468 ( .A0N(\i_MIPS/PC/n13 ), .A1N(net115789), .B0(n10180), .Y(
        n10181) );
  OR2X1 U469 ( .A(n10476), .B(n5560), .Y(n108) );
  OR2X1 U470 ( .A(n5557), .B(n10477), .Y(n109) );
  NAND3X2 U471 ( .A(n108), .B(n109), .C(n10475), .Y(\i_MIPS/PC/n46 ) );
  INVX20 U472 ( .A(n5563), .Y(n5560) );
  OR3X6 U473 ( .A(n10263), .B(n10262), .C(n10261), .Y(n110) );
  NAND2X6 U474 ( .A(n110), .B(n10260), .Y(n10487) );
  OR2XL U475 ( .A(n10268), .B(n5561), .Y(n111) );
  OR2XL U476 ( .A(n5557), .B(n10269), .Y(n112) );
  NAND3X2 U477 ( .A(n111), .B(n112), .C(n10267), .Y(\i_MIPS/PC/n49 ) );
  OR2XL U478 ( .A(n10141), .B(n5561), .Y(n113) );
  OR2XL U479 ( .A(n5557), .B(n10142), .Y(n114) );
  NAND3X2 U480 ( .A(n113), .B(n114), .C(n10140), .Y(\i_MIPS/PC/n41 ) );
  AOI2BB1X4 U481 ( .A0N(\i_MIPS/PC/n9 ), .A1N(net115789), .B0(n10139), .Y(
        n10140) );
  NAND2X2 U482 ( .A(n10466), .B(n115), .Y(n116) );
  NAND2X2 U483 ( .A(n10465), .B(n5545), .Y(n117) );
  NAND2X2 U484 ( .A(n116), .B(n117), .Y(n118) );
  INVX1 U485 ( .A(n5545), .Y(n115) );
  INVX3 U486 ( .A(n118), .Y(n10467) );
  AOI222X4 U487 ( .A0(n5541), .A1(n11420), .B0(mem_rdata_D[44]), .B1(n133), 
        .C0(n13001), .C1(n5539), .Y(n10466) );
  INVX6 U488 ( .A(n11420), .Y(n10465) );
  BUFX4 U489 ( .A(n5542), .Y(n5545) );
  BUFX4 U490 ( .A(n10467), .Y(n4516) );
  AND2X1 U491 ( .A(net104171), .B(net103849), .Y(n119) );
  AND2X2 U492 ( .A(net104172), .B(net103817), .Y(n120) );
  NOR3X4 U493 ( .A(n119), .B(n120), .C(n121), .Y(n4312) );
  NAND4X4 U494 ( .A(net106705), .B(net106706), .C(net106707), .D(net106708), 
        .Y(net103785) );
  OR2X2 U495 ( .A(\i_MIPS/n498 ), .B(net115791), .Y(n122) );
  OR2X1 U496 ( .A(\i_MIPS/n499 ), .B(net115791), .Y(n123) );
  INVX12 U497 ( .A(n5334), .Y(n3763) );
  INVX8 U498 ( .A(n9226), .Y(n9230) );
  OAI222X4 U499 ( .A0(n9297), .A1(net107688), .B0(net107217), .B1(n9309), .C0(
        net107689), .C1(n9296), .Y(n9325) );
  BUFX16 U500 ( .A(n5247), .Y(n5255) );
  OA22X2 U501 ( .A0(n5247), .A1(n639), .B0(n5287), .B1(n2256), .Y(n8831) );
  OA22X1 U502 ( .A0(n5247), .A1(n1132), .B0(n5287), .B1(n2755), .Y(n8819) );
  OA22X1 U503 ( .A0(n5247), .A1(n1144), .B0(n5287), .B1(n2767), .Y(n8922) );
  OA22XL U504 ( .A0(n5247), .A1(n610), .B0(n5287), .B1(n2228), .Y(n8823) );
  BUFX6 U505 ( .A(n5265), .Y(n5247) );
  NOR3X6 U506 ( .A(n4697), .B(n3681), .C(n7598), .Y(n7605) );
  BUFX8 U507 ( .A(n9574), .Y(n148) );
  NAND2X2 U508 ( .A(n4813), .B(net114073), .Y(n8792) );
  AND2X1 U509 ( .A(\i_MIPS/ALUin1[0] ), .B(n5062), .Y(n4813) );
  INVX3 U510 ( .A(n6915), .Y(n6925) );
  NAND4X6 U511 ( .A(n7964), .B(n7966), .C(n7965), .D(n7967), .Y(net104700) );
  AOI211X4 U512 ( .A0(n7948), .A1(n8208), .B0(n7947), .C0(n7946), .Y(n7967) );
  BUFX3 U513 ( .A(n5261), .Y(n5254) );
  BUFX8 U514 ( .A(n9806), .Y(n5261) );
  NAND2XL U515 ( .A(net108873), .B(n8637), .Y(n7961) );
  NAND2X8 U516 ( .A(n8202), .B(n8637), .Y(n7776) );
  NAND2X6 U517 ( .A(\i_MIPS/ALUin1[13] ), .B(n6693), .Y(n8637) );
  BUFX8 U518 ( .A(net108868), .Y(n124) );
  NAND2X8 U519 ( .A(n4624), .B(n6694), .Y(net111724) );
  INVX3 U520 ( .A(n11099), .Y(n125) );
  INVX3 U521 ( .A(n125), .Y(n126) );
  MXI2X4 U522 ( .A(n10739), .B(n10738), .S0(n5549), .Y(n10740) );
  NAND3X8 U523 ( .A(net107411), .B(net107210), .C(net117759), .Y(n8704) );
  INVX6 U524 ( .A(n6705), .Y(n6708) );
  NAND2X2 U525 ( .A(n7038), .B(n3674), .Y(n7313) );
  CLKMX2X12 U526 ( .A(n8039), .B(n8962), .S0(net114065), .Y(n9295) );
  MX2X1 U527 ( .A(net118597), .B(net118592), .S0(n9428), .Y(n6929) );
  INVX3 U528 ( .A(n6928), .Y(n9428) );
  NAND4X2 U529 ( .A(n7344), .B(n7343), .C(n7342), .D(n7341), .Y(n11479) );
  OA22XL U530 ( .A0(n5250), .A1(n1049), .B0(n5298), .B1(n2676), .Y(n7343) );
  NAND4X2 U531 ( .A(n8074), .B(n8073), .C(n8072), .D(n8071), .Y(n11481) );
  OA22XL U532 ( .A0(n5391), .A1(n1043), .B0(n5434), .B1(n2670), .Y(n8071) );
  OA22XL U533 ( .A0(n5253), .A1(n1044), .B0(n5293), .B1(n2671), .Y(n8073) );
  OA22X2 U534 ( .A0(n5250), .A1(n642), .B0(n5290), .B1(n2259), .Y(n8435) );
  BUFX12 U535 ( .A(n5264), .Y(n5250) );
  OA22X2 U536 ( .A0(n5333), .A1(n1083), .B0(n5360), .B1(n2706), .Y(n7714) );
  BUFX12 U537 ( .A(n5354), .Y(n5360) );
  BUFX16 U538 ( .A(n3875), .Y(n5333) );
  BUFX3 U539 ( .A(n5260), .Y(n3923) );
  NAND2X2 U540 ( .A(n7864), .B(n7863), .Y(n7867) );
  INVX16 U541 ( .A(n10962), .Y(n4533) );
  OR2X8 U542 ( .A(n3657), .B(n9943), .Y(n10962) );
  AND4X8 U543 ( .A(n6446), .B(n6447), .C(n6444), .D(n6445), .Y(n3919) );
  CLKINVX20 U544 ( .A(net143513), .Y(net143514) );
  CLKAND2X8 U545 ( .A(n8029), .B(n7770), .Y(n3006) );
  INVX4 U546 ( .A(n7766), .Y(n7770) );
  BUFX4 U547 ( .A(n9233), .Y(n127) );
  OAI221X2 U548 ( .A0(n2919), .A1(n5071), .B0(n336), .B1(n5067), .C0(n7954), 
        .Y(n8040) );
  NAND2X8 U549 ( .A(net111416), .B(\i_MIPS/n297 ), .Y(n9303) );
  INVX16 U550 ( .A(net112414), .Y(net111416) );
  AOI22X4 U551 ( .A0(net118217), .A1(net104941), .B0(net118227), .B1(net109762), .Y(net139775) );
  CLKMX2X4 U552 ( .A(n8160), .B(n8159), .S0(net114087), .Y(net109762) );
  NAND2X8 U553 ( .A(net144187), .B(n3559), .Y(n4621) );
  CLKMX2X6 U554 ( .A(\i_MIPS/n210 ), .B(n4780), .S0(n3894), .Y(n6718) );
  CLKMX2X6 U555 ( .A(\i_MIPS/n212 ), .B(n4781), .S0(n3894), .Y(n6717) );
  MX2X6 U556 ( .A(\i_MIPS/n204 ), .B(n4778), .S0(n3894), .Y(n6723) );
  MXI2X1 U557 ( .A(\i_MIPS/ID_EX[69] ), .B(\i_MIPS/ID_EX[101] ), .S0(n3894), 
        .Y(n6947) );
  NOR2X8 U558 ( .A(n3695), .B(n3783), .Y(n4329) );
  CLKINVX6 U559 ( .A(net105227), .Y(n4342) );
  CLKBUFX3 U560 ( .A(net107665), .Y(n128) );
  NAND2X2 U561 ( .A(n11590), .B(n11589), .Y(n11585) );
  NAND2X4 U562 ( .A(n5062), .B(\i_MIPS/ALUin1[13] ), .Y(n7953) );
  AOI211X2 U563 ( .A0(n3777), .A1(n9055), .B0(n9054), .C0(n9053), .Y(n9056) );
  CLKAND2X12 U564 ( .A(net112425), .B(n3022), .Y(n4278) );
  BUFX6 U565 ( .A(n5921), .Y(n5920) );
  NAND2XL U566 ( .A(n9204), .B(n9203), .Y(n9231) );
  NAND2X8 U567 ( .A(n6699), .B(n2921), .Y(n9203) );
  AOI2BB1X1 U568 ( .A0N(n3752), .A1N(net111256), .B0(n4305), .Y(n4304) );
  MX2X1 U569 ( .A(net109172), .B(net109496), .S0(net114065), .Y(net111256) );
  OA21X2 U570 ( .A0(\i_MIPS/ALUin1[19] ), .A1(n5068), .B0(n7104), .Y(n6829) );
  AOI2BB1X4 U571 ( .A0N(n2184), .A1N(n5068), .B0(n4794), .Y(n7030) );
  OAI221X2 U572 ( .A0(\i_MIPS/n299 ), .A1(n5072), .B0(n2928), .B1(n5068), .C0(
        n6834), .Y(n8865) );
  INVX20 U573 ( .A(n5069), .Y(n5068) );
  AND3X2 U574 ( .A(n3950), .B(n6729), .C(n6848), .Y(n6734) );
  INVX4 U575 ( .A(n6848), .Y(n6822) );
  NAND2X6 U576 ( .A(n4704), .B(n3636), .Y(n6848) );
  CLKMX2X6 U577 ( .A(n7599), .B(n4813), .S0(net114065), .Y(n9055) );
  AO22X4 U578 ( .A0(mem_rdata_I[103]), .A1(n5933), .B0(n5572), .B1(n11319), 
        .Y(n9910) );
  BUFX4 U579 ( .A(n11091), .Y(n5572) );
  NAND4X8 U580 ( .A(n6853), .B(n6852), .C(n6851), .D(n6850), .Y(net105290) );
  AND3X6 U581 ( .A(n4482), .B(n4483), .C(n6450), .Y(n3718) );
  NAND2BX2 U582 ( .AN(n5352), .B(\D_cache/cache[5][143] ), .Y(n4483) );
  NAND2X4 U583 ( .A(n3938), .B(n4736), .Y(n7694) );
  INVX4 U584 ( .A(net112549), .Y(n4000) );
  OR2X2 U585 ( .A(n5045), .B(n4087), .Y(n4086) );
  INVX4 U586 ( .A(net106596), .Y(net108012) );
  CLKMX2X3 U587 ( .A(\i_MIPS/n270 ), .B(\i_MIPS/n271 ), .S0(n5062), .Y(n7784)
         );
  BUFX8 U588 ( .A(n4714), .Y(n5062) );
  NAND3X8 U589 ( .A(ICACHE_addr[6]), .B(ICACHE_addr[5]), .C(n10158), .Y(n10167) );
  CLKINVX8 U590 ( .A(n10146), .Y(n10158) );
  OR2X2 U591 ( .A(n5045), .B(n4083), .Y(n4082) );
  OR2X2 U592 ( .A(n5045), .B(n4089), .Y(n4088) );
  AND2X8 U593 ( .A(n3733), .B(net105549), .Y(n4011) );
  NAND4X4 U594 ( .A(n8003), .B(n8002), .C(n8001), .D(n8000), .Y(n11421) );
  INVX4 U595 ( .A(n11408), .Y(n10747) );
  NAND4X2 U596 ( .A(n8756), .B(n8755), .C(n8754), .D(n8753), .Y(n11408) );
  NAND2X8 U597 ( .A(n4578), .B(n336), .Y(n8288) );
  BUFX12 U598 ( .A(n6720), .Y(n4578) );
  NAND4BX4 U599 ( .AN(n10732), .B(n10731), .C(n10730), .D(n10729), .Y(
        \i_MIPS/PC/n65 ) );
  NAND3X6 U600 ( .A(n7768), .B(n7769), .C(n3006), .Y(n8466) );
  NAND2X2 U601 ( .A(n4705), .B(n7767), .Y(n7769) );
  OAI221X4 U602 ( .A0(\i_MIPS/Register/register[18][3] ), .A1(net117643), .B0(
        \i_MIPS/Register/register[26][3] ), .B1(net117661), .C0(n9158), .Y(
        n9161) );
  BUFX16 U603 ( .A(net117665), .Y(net117661) );
  OR2X2 U604 ( .A(n5170), .B(n2177), .Y(n4617) );
  BUFX8 U605 ( .A(n5184), .Y(n5170) );
  MXI2X4 U606 ( .A(n10518), .B(n10517), .S0(n5546), .Y(n10519) );
  INVX4 U607 ( .A(n11461), .Y(n10517) );
  OR2X4 U608 ( .A(n5326), .B(n2918), .Y(n4482) );
  BUFX8 U609 ( .A(n5336), .Y(n5326) );
  INVX16 U610 ( .A(net143514), .Y(net144187) );
  CLKAND2X12 U611 ( .A(n9309), .B(n7302), .Y(n4727) );
  NAND2X6 U612 ( .A(\i_MIPS/ALUin1[5] ), .B(n6712), .Y(n9309) );
  INVX12 U613 ( .A(n6717), .Y(n6698) );
  OA22X4 U614 ( .A0(n6940), .A1(net117759), .B0(n9202), .B1(n7941), .Y(n6941)
         );
  CLKMX2X6 U615 ( .A(n7785), .B(n7788), .S0(net114065), .Y(n8557) );
  CLKMX2X3 U616 ( .A(n7786), .B(n7785), .S0(\i_MIPS/ID_EX[81] ), .Y(n7847) );
  OAI221X4 U617 ( .A0(n2892), .A1(n5071), .B0(n343), .B1(n5068), .C0(n7412), 
        .Y(n7785) );
  OA22X2 U618 ( .A0(\i_MIPS/Register/register[5][7] ), .A1(net118401), .B0(
        \i_MIPS/Register/register[13][7] ), .B1(net118425), .Y(n7322) );
  OA22X1 U619 ( .A0(\i_MIPS/Register/register[21][7] ), .A1(net118401), .B0(
        \i_MIPS/Register/register[29][7] ), .B1(net118425), .Y(n7331) );
  INVX4 U620 ( .A(net118415), .Y(net118401) );
  AO22X4 U621 ( .A0(mem_rdata_I[123]), .A1(n5944), .B0(n5573), .B1(n11338), 
        .Y(n9629) );
  BUFX20 U622 ( .A(n3020), .Y(n129) );
  BUFX12 U623 ( .A(n3020), .Y(n130) );
  BUFX12 U624 ( .A(n3020), .Y(n131) );
  BUFX12 U625 ( .A(n3020), .Y(n132) );
  BUFX12 U626 ( .A(n3020), .Y(n133) );
  AND2X6 U627 ( .A(n9798), .B(mem_ready_D), .Y(n3020) );
  AO21X1 U628 ( .A0(n9802), .A1(n3634), .B0(n11584), .Y(n11091) );
  NAND3X4 U629 ( .A(n11585), .B(net36572), .C(n11586), .Y(n11584) );
  NAND2X2 U630 ( .A(n5062), .B(\i_MIPS/ALUin1[30] ), .Y(n9447) );
  OR2X6 U631 ( .A(n5212), .B(n2890), .Y(n4618) );
  CLKBUFX6 U632 ( .A(n5223), .Y(n5212) );
  BUFX8 U633 ( .A(n6938), .Y(n134) );
  BUFX4 U634 ( .A(n5788), .Y(n5785) );
  NAND2X4 U635 ( .A(\i_MIPS/ALUin1[20] ), .B(n6688), .Y(n8382) );
  INVX2 U636 ( .A(n6723), .Y(n6688) );
  NAND4X2 U637 ( .A(n7808), .B(n7807), .C(n7806), .D(n7805), .Y(n11390) );
  OA22XL U638 ( .A0(n5393), .A1(n1065), .B0(n5436), .B1(n2693), .Y(n7805) );
  BUFX12 U639 ( .A(net111270), .Y(n3974) );
  OA22X2 U640 ( .A0(n5376), .A1(n638), .B0(n5429), .B1(n2255), .Y(n8829) );
  INVX8 U641 ( .A(n11422), .Y(n10107) );
  NAND4BX4 U642 ( .AN(n4647), .B(n7811), .C(n7810), .D(n7809), .Y(n11422) );
  BUFX12 U643 ( .A(n4677), .Y(n5841) );
  NAND4X4 U644 ( .A(n7716), .B(n7715), .C(n7714), .D(n7713), .Y(n11435) );
  OA22X1 U645 ( .A0(n5255), .A1(n2102), .B0(n5295), .B1(n476), .Y(n7715) );
  CLKMX2X4 U646 ( .A(n9042), .B(n8204), .S0(net114065), .Y(n8697) );
  OAI221X4 U647 ( .A0(\i_MIPS/ALUin1[11] ), .A1(n5071), .B0(
        \i_MIPS/ALUin1[10] ), .B1(n5067), .C0(n8130), .Y(n9042) );
  INVX2 U648 ( .A(net108005), .Y(n3637) );
  BUFX8 U649 ( .A(n150), .Y(n135) );
  AOI31X2 U650 ( .A0(n8696), .A1(n8695), .A2(n8694), .B0(n8693), .Y(n8713) );
  NAND2BX2 U651 ( .AN(n7688), .B(n11097), .Y(n9433) );
  OA22X4 U652 ( .A0(n5392), .A1(n636), .B0(n5435), .B1(n2253), .Y(n7903) );
  AOI33X4 U653 ( .A0(n3950), .A1(n7962), .A2(n7963), .B0(n3950), .B1(n7961), 
        .B2(n7960), .Y(n7964) );
  NAND3BX1 U654 ( .AN(n7951), .B(net117745), .C(n7950), .Y(n7966) );
  NAND4X2 U655 ( .A(n7712), .B(n7711), .C(n7710), .D(n7709), .Y(n11403) );
  OA22X2 U656 ( .A0(n5393), .A1(n1058), .B0(n5436), .B1(n2685), .Y(n7709) );
  OA22XL U657 ( .A0(n5255), .A1(n1060), .B0(n5295), .B1(n2687), .Y(n7711) );
  CLKINVX3 U658 ( .A(n4982), .Y(n5521) );
  CLKINVX3 U659 ( .A(n4982), .Y(n5520) );
  OR2X8 U660 ( .A(n4982), .B(net117623), .Y(n3987) );
  INVX4 U661 ( .A(n5742), .Y(n136) );
  INVX3 U662 ( .A(n136), .Y(n137) );
  INVX6 U663 ( .A(n136), .Y(n138) );
  INVX8 U664 ( .A(n11415), .Y(n10683) );
  NAND4X4 U665 ( .A(n7356), .B(n7355), .C(n7354), .D(n7353), .Y(n11415) );
  INVX12 U666 ( .A(n9204), .Y(n8565) );
  BUFX6 U667 ( .A(n6947), .Y(n145) );
  BUFX8 U668 ( .A(n10735), .Y(n3677) );
  AND2XL U669 ( .A(net139859), .B(net104915), .Y(n4694) );
  AND2X8 U670 ( .A(net139859), .B(net104915), .Y(n3775) );
  AOI22X4 U671 ( .A0(net118215), .A1(net104918), .B0(net118225), .B1(net108249), .Y(net139859) );
  NOR4X2 U672 ( .A(n11), .B(\i_MIPS/ID_EX[76] ), .C(n3682), .D(n3621), .Y(
        n6651) );
  AND2X8 U673 ( .A(n6711), .B(n1302), .Y(n3854) );
  AND3X8 U674 ( .A(n4634), .B(n4635), .C(n6436), .Y(n3972) );
  NAND2X4 U675 ( .A(n5205), .B(\D_cache/cache[1][137] ), .Y(n4635) );
  MXI2X4 U676 ( .A(n10454), .B(n10453), .S0(n5545), .Y(n10455) );
  AOI222X4 U677 ( .A0(n5541), .A1(n11423), .B0(mem_rdata_D[47]), .B1(n131), 
        .C0(n12998), .C1(n5539), .Y(n10454) );
  NAND3BX2 U678 ( .AN(n7696), .B(n3950), .C(n7695), .Y(n7697) );
  AOI222X2 U679 ( .A0(n4505), .A1(n11469), .B0(mem_rdata_D[93]), .B1(n130), 
        .C0(n12984), .C1(n5536), .Y(n10559) );
  AOI222X2 U680 ( .A0(n4505), .A1(n11454), .B0(mem_rdata_D[78]), .B1(n129), 
        .C0(n12999), .C1(n5535), .Y(n10102) );
  MXI2X4 U681 ( .A(n10690), .B(n10689), .S0(n5549), .Y(n10691) );
  INVX8 U682 ( .A(n11425), .Y(n10628) );
  NAND4X4 U683 ( .A(n9270), .B(n9269), .C(n9268), .D(n9267), .Y(n11425) );
  NAND4X6 U684 ( .A(n9361), .B(n9360), .C(n9359), .D(n9358), .Y(n11413) );
  OA22XL U685 ( .A0(n5333), .A1(n986), .B0(n5358), .B1(n2611), .Y(n9359) );
  AOI222X2 U686 ( .A0(n4506), .A1(n11470), .B0(mem_rdata_D[94]), .B1(n133), 
        .C0(n12983), .C1(n5536), .Y(n10596) );
  BUFX12 U687 ( .A(n10776), .Y(n4539) );
  BUFX12 U688 ( .A(n10547), .Y(n4565) );
  AOI222X2 U689 ( .A0(n4506), .A1(n11452), .B0(mem_rdata_D[76]), .B1(n131), 
        .C0(n13001), .C1(n5535), .Y(n10460) );
  BUFX12 U690 ( .A(n10396), .Y(n4553) );
  BUFX12 U691 ( .A(n10312), .Y(n4554) );
  BUFX12 U692 ( .A(n10624), .Y(n4568) );
  AOI222X2 U693 ( .A0(n4506), .A1(n11448), .B0(mem_rdata_D[72]), .B1(n130), 
        .C0(n13005), .C1(n5536), .Y(n10651) );
  NOR4X4 U694 ( .A(n9558), .B(n9560), .C(n9559), .D(n9561), .Y(n9573) );
  OAI222X4 U695 ( .A0(n9552), .A1(net107230), .B0(n9551), .B1(n9550), .C0(
        \i_MIPS/n270 ), .C1(n9549), .Y(n9560) );
  NAND2X4 U696 ( .A(\i_MIPS/ALUin1[3] ), .B(n3698), .Y(n9126) );
  NAND2X8 U697 ( .A(n3698), .B(n2928), .Y(n9121) );
  BUFX8 U698 ( .A(n8650), .Y(n3698) );
  NAND2X4 U699 ( .A(\i_MIPS/ALUin1[1] ), .B(n3606), .Y(net111572) );
  NOR2X6 U700 ( .A(n3606), .B(\i_MIPS/n300 ), .Y(net134145) );
  NAND2X4 U701 ( .A(n3606), .B(\i_MIPS/n300 ), .Y(net111570) );
  MXI2X8 U702 ( .A(n4021), .B(\i_MIPS/n242 ), .S0(net143504), .Y(n3606) );
  OA22X4 U703 ( .A0(n10692), .A1(n3879), .B0(n10695), .B1(n4495), .Y(n7077) );
  MX2X6 U704 ( .A(n10695), .B(n10696), .S0(n4410), .Y(n3825) );
  OR2XL U705 ( .A(n5040), .B(n10695), .Y(n3946) );
  INVX3 U706 ( .A(n11431), .Y(n10695) );
  AOI222X1 U707 ( .A0(n3800), .A1(n11395), .B0(mem_rdata_D[19]), .B1(n133), 
        .C0(n5538), .C1(n12994), .Y(n10972) );
  BUFX20 U708 ( .A(n4684), .Y(n5538) );
  NOR4X4 U709 ( .A(n7606), .B(n7605), .C(n7604), .D(n7603), .Y(n7607) );
  MXI2X4 U710 ( .A(n10405), .B(n10404), .S0(n5544), .Y(n10406) );
  AOI222X4 U711 ( .A0(n4535), .A1(n11492), .B0(mem_rdata_D[116]), .B1(n133), 
        .C0(n12993), .C1(n5533), .Y(n10405) );
  BUFX8 U712 ( .A(n10419), .Y(n4556) );
  BUFX8 U713 ( .A(n10433), .Y(n4555) );
  OA22X2 U714 ( .A0(n9453), .A1(n9452), .B0(n9552), .B1(n9451), .Y(n9454) );
  OAI222X2 U715 ( .A0(n8863), .A1(n7788), .B0(net108781), .B1(n7787), .C0(
        n3673), .C1(n7847), .Y(n9451) );
  BUFX6 U716 ( .A(n9232), .Y(n139) );
  NOR4X6 U717 ( .A(n6943), .B(n6944), .C(n6945), .D(n6942), .Y(n6959) );
  OAI221X2 U718 ( .A0(n8855), .A1(n9550), .B0(net107217), .B1(n9424), .C0(
        n6941), .Y(n6942) );
  NOR2BX4 U719 ( .AN(n3762), .B(\i_MIPS/n270 ), .Y(net134069) );
  AOI32X2 U720 ( .A0(n8970), .A1(\i_MIPS/ALUin1[1] ), .A2(n3762), .B0(
        net108306), .B1(\i_MIPS/ALUin1[1] ), .Y(n8971) );
  INVX1 U721 ( .A(n5059), .Y(n3762) );
  NAND2X2 U722 ( .A(net117747), .B(n8281), .Y(n8285) );
  INVX6 U723 ( .A(n8281), .Y(n8309) );
  NAND2X2 U724 ( .A(n3665), .B(n8683), .Y(n8281) );
  NAND4X8 U725 ( .A(n139), .B(n3742), .C(n127), .D(n9234), .Y(n10619) );
  NAND2X2 U726 ( .A(n6696), .B(\i_MIPS/n287 ), .Y(net108869) );
  NOR2X8 U727 ( .A(n6696), .B(\i_MIPS/ALUin1[14] ), .Y(n3764) );
  INVX4 U728 ( .A(n6715), .Y(n6696) );
  INVX3 U729 ( .A(net111572), .Y(net112512) );
  CLKBUFX3 U730 ( .A(n5884), .Y(n5851) );
  CLKBUFX3 U731 ( .A(n5884), .Y(n5879) );
  AO21X4 U732 ( .A0(n9218), .A1(n3628), .B0(n8280), .Y(n3967) );
  OAI221X2 U733 ( .A0(n344), .A1(n5071), .B0(n183), .B1(n5067), .C0(n7944), 
        .Y(n8039) );
  INVX8 U734 ( .A(n11416), .Y(n10656) );
  NAND4X4 U735 ( .A(n8176), .B(n8175), .C(n8174), .D(n8173), .Y(n11416) );
  BUFX20 U736 ( .A(n4757), .Y(n5554) );
  CLKBUFX6 U737 ( .A(n4757), .Y(n5553) );
  AO22X4 U738 ( .A0(n4757), .A1(DCACHE_addr[18]), .B0(n5552), .B1(n11522), .Y(
        n11038) );
  AO22X4 U739 ( .A0(n4757), .A1(DCACHE_addr[11]), .B0(n5552), .B1(n11515), .Y(
        n11025) );
  AO22X4 U740 ( .A0(n4757), .A1(DCACHE_addr[23]), .B0(n5552), .B1(n11527), .Y(
        n11033) );
  AO22X4 U741 ( .A0(n4757), .A1(DCACHE_addr[15]), .B0(n5552), .B1(n11519), .Y(
        n11030) );
  CLKAND2X4 U742 ( .A(n129), .B(n10979), .Y(n4757) );
  AOI211X2 U743 ( .A0(net109168), .A1(n9322), .B0(n7958), .C0(n7957), .Y(n7965) );
  NAND3BX4 U744 ( .AN(n4817), .B(n4802), .C(n10279), .Y(n10290) );
  NAND3X6 U745 ( .A(n10487), .B(n10264), .C(n10254), .Y(n10279) );
  NAND4X2 U746 ( .A(n8436), .B(n8435), .C(n8434), .D(n8433), .Y(n11428) );
  OA22X2 U747 ( .A0(n5395), .A1(n641), .B0(n5431), .B1(n2258), .Y(n8433) );
  NAND2X6 U748 ( .A(n4737), .B(n9956), .Y(n9943) );
  INVX6 U749 ( .A(n6718), .Y(n6699) );
  MXI2X4 U750 ( .A(n10648), .B(n10647), .S0(n5548), .Y(n10649) );
  AOI222X4 U751 ( .A0(n4534), .A1(n11480), .B0(mem_rdata_D[104]), .B1(n129), 
        .C0(n13005), .C1(n5534), .Y(n10648) );
  CLKINVX8 U752 ( .A(n10711), .Y(n9597) );
  INVX16 U753 ( .A(n4533), .Y(n4535) );
  MXI2X4 U754 ( .A(n10099), .B(n10098), .S0(n5542), .Y(n10100) );
  AOI222X4 U755 ( .A0(n4535), .A1(n11486), .B0(mem_rdata_D[110]), .B1(n129), 
        .C0(n12999), .C1(n5533), .Y(n10099) );
  AOI222X1 U756 ( .A0(n4535), .A1(n11476), .B0(mem_rdata_D[100]), .B1(n130), 
        .C0(n13009), .C1(n5533), .Y(n9805) );
  OAI2BB1X4 U757 ( .A0N(n3967), .A1N(n8550), .B0(n8556), .Y(n8310) );
  INVX3 U758 ( .A(n8683), .Y(n8680) );
  CLKINVX8 U759 ( .A(n10481), .Y(n10491) );
  NAND3X8 U760 ( .A(ICACHE_addr[10]), .B(ICACHE_addr[9]), .C(n10471), .Y(
        n10481) );
  OAI221X1 U761 ( .A0(n10150), .A1(n5562), .B0(n5558), .B1(n10151), .C0(n10149), .Y(\i_MIPS/PC/n42 ) );
  XOR2X4 U762 ( .A(n11347), .B(ICACHE_addr[5]), .Y(n6384) );
  NAND4X4 U763 ( .A(n4670), .B(n6375), .C(n6374), .D(n6373), .Y(n11347) );
  INVX12 U764 ( .A(n5563), .Y(n5562) );
  OAI221X2 U765 ( .A0(n8863), .A1(n8862), .B0(n3673), .B1(n9295), .C0(n8861), 
        .Y(n9315) );
  XNOR2X4 U766 ( .A(n10716), .B(ICACHE_addr[29]), .Y(n4676) );
  CLKINVX8 U767 ( .A(n9437), .Y(n7689) );
  NAND2X4 U768 ( .A(n4739), .B(n11103), .Y(n9437) );
  MXI2X4 U769 ( .A(\i_MIPS/ID_EX[95] ), .B(\i_MIPS/ID_EX[63] ), .S0(net144187), 
        .Y(n6725) );
  AOI2BB1X1 U770 ( .A0N(\i_MIPS/PC/n10 ), .A1N(net115789), .B0(n10148), .Y(
        n10149) );
  NAND2X6 U771 ( .A(n4708), .B(n8859), .Y(n6814) );
  CLKAND2X12 U772 ( .A(n8397), .B(n8688), .Y(n4708) );
  OAI221X2 U773 ( .A0(\i_MIPS/n300 ), .A1(n5073), .B0(\i_MIPS/n299 ), .B1(
        n5067), .C0(n6671), .Y(n7599) );
  OAI222X1 U774 ( .A0(n9202), .A1(n7846), .B0(n5049), .B1(n9444), .C0(n9453), 
        .C1(n8856), .Y(n7853) );
  OAI221X2 U775 ( .A0(n7420), .A1(n8863), .B0(n3673), .B1(n7789), .C0(n8861), 
        .Y(n7846) );
  CLKMX2X4 U776 ( .A(n8040), .B(n8039), .S0(net114065), .Y(n8961) );
  NAND3BX4 U777 ( .AN(n4822), .B(n4803), .C(n10319), .Y(n10331) );
  NAND3X4 U778 ( .A(n10288), .B(n10291), .C(n10290), .Y(n10319) );
  NAND3X8 U779 ( .A(ICACHE_addr[22]), .B(ICACHE_addr[21]), .C(n10371), .Y(
        n10376) );
  CLKINVX8 U780 ( .A(n10364), .Y(n10371) );
  OAI221X4 U781 ( .A0(n10572), .A1(n5560), .B0(n5558), .B1(n10573), .C0(n10571), .Y(\i_MIPS/PC/n63 ) );
  INVX8 U782 ( .A(n10573), .Y(n10575) );
  XOR2X4 U783 ( .A(n10576), .B(ICACHE_addr[27]), .Y(n10573) );
  OAI221X2 U784 ( .A0(n10720), .A1(n10719), .B0(n3027), .B1(n10736), .C0(
        n10718), .Y(n10732) );
  NAND2X8 U785 ( .A(n6688), .B(n2919), .Y(n8688) );
  CLKINVX8 U786 ( .A(net108781), .Y(net108310) );
  BUFX16 U787 ( .A(n5197), .Y(n5225) );
  XNOR2X2 U788 ( .A(n11350), .B(ICACHE_addr[8]), .Y(n11165) );
  XNOR2X2 U789 ( .A(ICACHE_addr[7]), .B(n11349), .Y(n11166) );
  XNOR2X2 U790 ( .A(ICACHE_addr[6]), .B(n11348), .Y(n11167) );
  NAND2X4 U791 ( .A(n11046), .B(n11045), .Y(n6467) );
  NAND2X4 U792 ( .A(n11007), .B(n3007), .Y(n6443) );
  BUFX4 U793 ( .A(net134685), .Y(net118481) );
  NAND2X4 U794 ( .A(n11034), .B(n3718), .Y(n4671) );
  BUFX6 U795 ( .A(n5132), .Y(n5135) );
  CLKINVX12 U796 ( .A(net143503), .Y(net143513) );
  NAND2X2 U797 ( .A(n6939), .B(n2961), .Y(n11110) );
  AOI2BB1X1 U798 ( .A0N(\i_MIPS/ALUin1[16] ), .A1N(n5059), .B0(n4730), .Y(
        n6657) );
  AOI2BB1X1 U799 ( .A0N(\i_MIPS/ALUin1[17] ), .A1N(n5059), .B0(n4731), .Y(
        n6839) );
  INVX6 U800 ( .A(n6608), .Y(n6610) );
  NAND2X4 U801 ( .A(n248), .B(\i_MIPS/n505 ), .Y(n6608) );
  AND2X4 U802 ( .A(net108631), .B(n3674), .Y(net134907) );
  BUFX4 U803 ( .A(net118281), .Y(net118267) );
  BUFX4 U804 ( .A(net117641), .Y(net117635) );
  CLKINVX8 U805 ( .A(net118369), .Y(net118351) );
  CLKINVX4 U806 ( .A(n9556), .Y(n9555) );
  CLKINVX1 U807 ( .A(n9543), .Y(n9557) );
  CLKMX2X2 U808 ( .A(n8703), .B(n8701), .S0(net114065), .Y(n8373) );
  BUFX6 U809 ( .A(n11210), .Y(n5921) );
  CLKBUFX8 U810 ( .A(n135), .Y(n5655) );
  CLKINVX6 U811 ( .A(n5447), .Y(n3755) );
  INVX6 U812 ( .A(n5263), .Y(n3856) );
  CLKAND2X8 U813 ( .A(n8699), .B(\i_MIPS/n270 ), .Y(n4724) );
  INVX8 U814 ( .A(n8699), .Y(n8291) );
  INVX8 U815 ( .A(n5075), .Y(n5071) );
  NAND4X2 U816 ( .A(n7415), .B(n7414), .C(net107389), .D(n7413), .Y(n7427) );
  NAND4X2 U817 ( .A(n6837), .B(n6836), .C(net107389), .D(n6835), .Y(n6846) );
  OAI222X1 U818 ( .A0(n8863), .A1(n7422), .B0(net118601), .B1(n7480), .C0(
        n7478), .C1(n8699), .Y(n7159) );
  OAI222X1 U819 ( .A0(n8863), .A1(n7422), .B0(net118601), .B1(n7480), .C0(
        n7478), .C1(n8699), .Y(n3631) );
  BUFX16 U820 ( .A(n5312), .Y(n5305) );
  INVX2 U821 ( .A(n5097), .Y(n5096) );
  INVX12 U822 ( .A(net107138), .Y(net107607) );
  CLKBUFX8 U823 ( .A(net118223), .Y(net118215) );
  CLKBUFX4 U824 ( .A(n5788), .Y(n5786) );
  BUFX8 U825 ( .A(n5655), .Y(n5652) );
  BUFX2 U826 ( .A(n5788), .Y(n5787) );
  BUFX4 U827 ( .A(n5655), .Y(n5654) );
  BUFX4 U828 ( .A(n5840), .Y(n5832) );
  BUFX12 U829 ( .A(n5921), .Y(n5919) );
  BUFX4 U830 ( .A(n5404), .Y(n5385) );
  BUFX12 U831 ( .A(n5449), .Y(n5438) );
  BUFX16 U832 ( .A(n5264), .Y(n5248) );
  BUFX6 U833 ( .A(n5264), .Y(n5249) );
  BUFX16 U834 ( .A(n5185), .Y(n5175) );
  XOR2XL U835 ( .A(\i_MIPS/n497 ), .B(\i_MIPS/Reg_W[3] ), .Y(n6767) );
  CLKINVX1 U836 ( .A(n11244), .Y(n3798) );
  CLKINVX1 U837 ( .A(n11306), .Y(n3805) );
  OA22XL U838 ( .A0(n9211), .A1(n8878), .B0(n9316), .B1(n8035), .Y(n8048) );
  NAND3X4 U839 ( .A(ICACHE_addr[18]), .B(ICACHE_addr[17]), .C(n10333), .Y(
        n10341) );
  NAND4X4 U840 ( .A(n6561), .B(n6560), .C(n6559), .D(n6558), .Y(n11373) );
  INVX3 U841 ( .A(n11386), .Y(n10777) );
  CLKAND2X3 U842 ( .A(n4505), .B(n11442), .Y(n4386) );
  CLKINVX4 U843 ( .A(n11490), .Y(n10634) );
  INVX3 U844 ( .A(n11487), .Y(n10444) );
  BUFX4 U845 ( .A(\i_MIPS/jump_addr[22] ), .Y(net114079) );
  NAND3X4 U846 ( .A(ICACHE_addr[20]), .B(ICACHE_addr[19]), .C(n10354), .Y(
        n10364) );
  NAND4X1 U847 ( .A(n10882), .B(n10881), .C(n10880), .D(n10879), .Y(n11220) );
  NAND4X1 U848 ( .A(n9926), .B(n9925), .C(n9924), .D(n9923), .Y(n11225) );
  NAND4X1 U849 ( .A(n9921), .B(n9920), .C(n9919), .D(n9918), .Y(n11287) );
  INVX6 U850 ( .A(n11361), .Y(n11202) );
  NAND2X6 U851 ( .A(n11024), .B(n11023), .Y(n6495) );
  AND2X4 U852 ( .A(n10985), .B(n12962), .Y(n3782) );
  NAND2X2 U853 ( .A(n10984), .B(n10985), .Y(n6408) );
  NAND2X4 U854 ( .A(n10991), .B(n10990), .Y(n6398) );
  NAND2X4 U855 ( .A(n11032), .B(n11031), .Y(n6481) );
  NAND2X4 U856 ( .A(n11029), .B(n11028), .Y(n6486) );
  NAND2X4 U857 ( .A(n11049), .B(n11048), .Y(n6462) );
  NOR2X4 U858 ( .A(n6476), .B(n6474), .Y(n4370) );
  MX2X6 U859 ( .A(\i_MIPS/ID_EX[50] ), .B(n3673), .S0(n3894), .Y(n3583) );
  INVX3 U860 ( .A(n8026), .Y(n8028) );
  CLKINVX6 U861 ( .A(n3583), .Y(n6702) );
  BUFX4 U862 ( .A(net107615), .Y(net118243) );
  OA21X2 U863 ( .A0(\i_MIPS/ALUin1[15] ), .A1(n5073), .B0(n8131), .Y(n8132) );
  INVX4 U864 ( .A(n6724), .Y(n6689) );
  AND2X4 U865 ( .A(n11018), .B(n11017), .Y(n4099) );
  NOR2X6 U866 ( .A(n6503), .B(n6502), .Y(n6515) );
  CLKAND2X8 U867 ( .A(n11003), .B(n11002), .Y(n3882) );
  OA22XL U868 ( .A0(\i_MIPS/Register/register[6][18] ), .A1(net117685), .B0(
        \i_MIPS/Register/register[14][18] ), .B1(net117697), .Y(n8579) );
  AND4X6 U869 ( .A(n4673), .B(\i_MIPS/n258 ), .C(\i_MIPS/n256 ), .D(n3621), 
        .Y(n4672) );
  AND2X6 U870 ( .A(n9539), .B(n11108), .Y(n4728) );
  CLKINVX1 U871 ( .A(n7594), .Y(n7598) );
  NAND2XL U872 ( .A(n7585), .B(n9429), .Y(n7594) );
  NOR2BX2 U873 ( .AN(n5065), .B(\i_MIPS/n271 ), .Y(n4810) );
  BUFX4 U874 ( .A(n5132), .Y(n5136) );
  INVX3 U875 ( .A(net118409), .Y(net118407) );
  NAND2X1 U876 ( .A(n5074), .B(n2921), .Y(n7158) );
  NAND2X2 U877 ( .A(n7434), .B(net117745), .Y(n7401) );
  BUFX8 U878 ( .A(n6726), .Y(n4546) );
  AOI2BB1XL U879 ( .A0N(\i_MIPS/ALUin1[16] ), .A1N(n5073), .B0(n4746), .Y(
        n7033) );
  NAND2X1 U880 ( .A(\i_MIPS/ALUin1[27] ), .B(n6951), .Y(n11099) );
  INVX1 U881 ( .A(n6832), .Y(n6931) );
  INVX6 U882 ( .A(n3862), .Y(n4755) );
  AOI2BB1X2 U883 ( .A0N(n2928), .A1N(n5073), .B0(n4795), .Y(n7232) );
  NAND2X6 U884 ( .A(n7864), .B(n8695), .Y(n6817) );
  MX2X2 U885 ( .A(n7671), .B(n7682), .S0(net114065), .Y(n9551) );
  INVX6 U886 ( .A(net109512), .Y(net110429) );
  NAND2X6 U887 ( .A(\i_MIPS/ALUin1[17] ), .B(n6718), .Y(n9204) );
  BUFX16 U888 ( .A(n9503), .Y(n5142) );
  CLKBUFX6 U889 ( .A(n5078), .Y(n5077) );
  NAND2X6 U890 ( .A(n3995), .B(\D_cache/cache[0][154] ), .Y(n6522) );
  OR2X6 U891 ( .A(n5263), .B(n3975), .Y(n6520) );
  NOR2X2 U892 ( .A(n5353), .B(n2012), .Y(n3834) );
  AND2X2 U893 ( .A(n1319), .B(n3003), .Y(n4689) );
  CLKAND2X3 U894 ( .A(n5065), .B(n959), .Y(n4731) );
  AND2X2 U895 ( .A(n5070), .B(n2921), .Y(n4746) );
  BUFX6 U896 ( .A(net118241), .Y(net118233) );
  BUFX4 U897 ( .A(net118281), .Y(net118269) );
  NAND2X1 U898 ( .A(n3673), .B(\i_MIPS/n270 ), .Y(n7419) );
  OA22XL U899 ( .A0(\i_MIPS/Register/register[22][9] ), .A1(net139810), .B0(
        \i_MIPS/Register/register[30][9] ), .B1(net117695), .Y(n8063) );
  INVX6 U900 ( .A(net118483), .Y(net118477) );
  OA22X1 U901 ( .A0(\i_MIPS/Register/register[6][21] ), .A1(net117681), .B0(
        \i_MIPS/Register/register[14][21] ), .B1(net117697), .Y(n8903) );
  BUFX4 U902 ( .A(net118281), .Y(net118273) );
  AO21XL U903 ( .A0(n9553), .A1(n5049), .B0(net107228), .Y(n9554) );
  NAND4X2 U904 ( .A(n6634), .B(n6754), .C(n6633), .D(n10848), .Y(n6635) );
  INVX12 U905 ( .A(n5406), .Y(n3863) );
  OA22XL U906 ( .A0(\i_MIPS/Register/register[17][24] ), .A1(net118455), .B0(
        \i_MIPS/Register/register[25][24] ), .B1(net118479), .Y(n6784) );
  NAND4X1 U907 ( .A(n6774), .B(n6773), .C(n6772), .D(n6771), .Y(n6780) );
  OR2XL U908 ( .A(n9043), .B(net107987), .Y(n3910) );
  OAI221XL U909 ( .A0(\i_MIPS/Register/register[18][25] ), .A1(net117635), 
        .B0(\i_MIPS/Register/register[26][25] ), .B1(net117653), .C0(n6885), 
        .Y(n6888) );
  AO22XL U910 ( .A0(net118235), .A1(n182), .B0(net118259), .B1(n261), .Y(n6886) );
  OA22XL U911 ( .A0(\i_MIPS/Register/register[22][17] ), .A1(net117681), .B0(
        \i_MIPS/Register/register[30][17] ), .B1(net117703), .Y(n9248) );
  BUFX4 U912 ( .A(net118281), .Y(net118275) );
  CLKBUFX8 U913 ( .A(net118241), .Y(net118239) );
  NOR4X1 U914 ( .A(\i_MIPS/forward_unit/n10 ), .B(n6763), .C(n6762), .D(n6761), 
        .Y(n6764) );
  AO22XL U915 ( .A0(n5157), .A1(n555), .B0(n5153), .B1(n2174), .Y(n8350) );
  AO22XL U916 ( .A0(n5148), .A1(n554), .B0(n5144), .B1(n2173), .Y(n8351) );
  OAI221XL U917 ( .A0(\i_MIPS/Register/register[2][19] ), .A1(n5090), .B0(
        \i_MIPS/Register/register[10][19] ), .B1(n4669), .C0(n8349), .Y(n8357)
         );
  CLKINVX1 U918 ( .A(n9434), .Y(n9435) );
  CLKINVX4 U919 ( .A(n3748), .Y(n9552) );
  NAND2BX2 U920 ( .AN(n2948), .B(\i_MIPS/n161 ), .Y(n10154) );
  CLKBUFX3 U921 ( .A(n4713), .Y(n5111) );
  NAND2X4 U922 ( .A(net108310), .B(\i_MIPS/n270 ), .Y(n8861) );
  CLKINVX6 U923 ( .A(n5097), .Y(n5094) );
  NAND2BX1 U924 ( .AN(n10153), .B(n10154), .Y(n10261) );
  INVXL U925 ( .A(n8280), .Y(n3676) );
  AND3X4 U926 ( .A(n6946), .B(net117745), .C(n7585), .Y(n4733) );
  NAND2X1 U927 ( .A(n11112), .B(n11110), .Y(n6960) );
  NAND2XL U928 ( .A(n6928), .B(n9424), .Y(n6946) );
  CLKINVX1 U929 ( .A(n8137), .Y(n8790) );
  CLKMX2X4 U930 ( .A(n7583), .B(n6659), .S0(\i_MIPS/ID_EX[81] ), .Y(n8789) );
  NAND2X2 U931 ( .A(n11096), .B(n7400), .Y(n7688) );
  INVX6 U932 ( .A(n6921), .Y(n3983) );
  OA22X1 U933 ( .A0(net117757), .A1(n3613), .B0(n7431), .B1(net107217), .Y(
        n3612) );
  CLKINVX1 U934 ( .A(n6838), .Y(n3613) );
  NOR3X4 U935 ( .A(n8871), .B(n2993), .C(n8870), .Y(n8877) );
  AOI2BB1X1 U936 ( .A0N(n8875), .A1N(n8874), .B0(net107841), .Y(n8876) );
  CLKINVX2 U937 ( .A(n6932), .Y(n8879) );
  INVX4 U938 ( .A(n9049), .Y(n8372) );
  NAND2X2 U939 ( .A(n9445), .B(net114065), .Y(n8874) );
  NAND2X6 U940 ( .A(n8283), .B(n8566), .Y(n8394) );
  NAND2X1 U941 ( .A(n8370), .B(n8688), .Y(n8385) );
  INVX3 U942 ( .A(n8477), .Y(n7493) );
  NAND2X6 U943 ( .A(n9445), .B(net114073), .Y(n8878) );
  INVXL U944 ( .A(n7787), .Y(n8553) );
  NAND3BX2 U945 ( .AN(n9796), .B(DCACHE_ren), .C(n5193), .Y(n9797) );
  CLKAND2X8 U946 ( .A(n4719), .B(n4725), .Y(n4683) );
  INVX3 U947 ( .A(n5098), .Y(n5092) );
  INVX3 U948 ( .A(n5098), .Y(n5093) );
  CLKAND2X4 U949 ( .A(n3673), .B(net108631), .Y(n4718) );
  BUFX8 U950 ( .A(net108779), .Y(net118601) );
  BUFX16 U951 ( .A(n3770), .Y(n5049) );
  INVXL U952 ( .A(n8293), .Y(n7683) );
  CLKMX2X2 U953 ( .A(n8386), .B(n7599), .S0(net114065), .Y(n8137) );
  BUFX4 U954 ( .A(net118281), .Y(net118271) );
  NAND2X4 U955 ( .A(n2938), .B(net105396), .Y(n4362) );
  INVX2 U956 ( .A(n8373), .Y(n9043) );
  OA22XL U957 ( .A0(n5395), .A1(n2107), .B0(n5439), .B1(n481), .Y(n7273) );
  INVX12 U958 ( .A(n5306), .Y(n3924) );
  OA22XL U959 ( .A0(n5393), .A1(n2142), .B0(n5429), .B1(n517), .Y(n8924) );
  BUFX12 U960 ( .A(n5186), .Y(n5173) );
  CLKINVX6 U961 ( .A(n11372), .Y(n11375) );
  INVX4 U962 ( .A(n6466), .Y(n11045) );
  INVX4 U963 ( .A(n6402), .Y(n10987) );
  INVX3 U964 ( .A(n6454), .Y(n11036) );
  INVX8 U965 ( .A(n11535), .Y(n5041) );
  NAND2X6 U966 ( .A(n3748), .B(n3674), .Y(n8793) );
  OA22XL U967 ( .A0(n5400), .A1(n2159), .B0(n5440), .B1(n540), .Y(n6735) );
  OA22XL U968 ( .A0(\i_MIPS/Register/register[22][24] ), .A1(n5081), .B0(
        \i_MIPS/Register/register[30][24] ), .B1(n5076), .Y(n6620) );
  OA22XL U969 ( .A0(\i_MIPS/Register/register[6][24] ), .A1(n5081), .B0(
        \i_MIPS/Register/register[14][24] ), .B1(n5076), .Y(n6611) );
  OA22XL U970 ( .A0(\i_MIPS/Register/register[6][22] ), .A1(n5082), .B0(
        \i_MIPS/Register/register[14][22] ), .B1(n5078), .Y(n7879) );
  OA22X1 U971 ( .A0(\i_MIPS/Register/register[20][3] ), .A1(n5099), .B0(
        \i_MIPS/Register/register[28][3] ), .B1(n5096), .Y(n9198) );
  OA22X1 U972 ( .A0(\i_MIPS/Register/register[4][3] ), .A1(n5099), .B0(
        \i_MIPS/Register/register[12][3] ), .B1(n5096), .Y(n9189) );
  CLKINVX1 U973 ( .A(n10289), .Y(n10291) );
  INVX16 U974 ( .A(net107217), .Y(net107404) );
  INVX12 U975 ( .A(n3866), .Y(net107389) );
  NOR2X6 U976 ( .A(net108631), .B(n3758), .Y(n3866) );
  OA22XL U977 ( .A0(n5175), .A1(n719), .B0(n5214), .B1(n2341), .Y(n8603) );
  AOI2BB2XL U978 ( .B0(n3763), .B1(\D_cache/cache[4][50] ), .A0N(n5356), .A1N(
        n2041), .Y(n8601) );
  NAND4BX2 U979 ( .AN(n9115), .B(n9114), .C(n9113), .D(n9112), .Y(n9116) );
  OAI221XL U980 ( .A0(\i_MIPS/Register/register[18][4] ), .A1(n5088), .B0(
        \i_MIPS/Register/register[26][4] ), .B1(n5086), .C0(n9107), .Y(n9115)
         );
  NAND2X6 U981 ( .A(net109168), .B(net114065), .Y(net107689) );
  CLKMX2X3 U982 ( .A(n9041), .B(n9040), .S0(net114079), .Y(net108160) );
  CLKAND2X6 U983 ( .A(net118227), .B(n7525), .Y(net143525) );
  AND2X4 U984 ( .A(net118217), .B(net105121), .Y(net143524) );
  INVX3 U985 ( .A(net111509), .Y(net105731) );
  OAI221XL U986 ( .A0(\i_MIPS/Register/register[2][17] ), .A1(n5091), .B0(
        \i_MIPS/Register/register[10][17] ), .B1(n5086), .C0(n9273), .Y(n9281)
         );
  OA22XL U987 ( .A0(\i_MIPS/Register/register[4][5] ), .A1(n5101), .B0(
        \i_MIPS/Register/register[12][5] ), .B1(n5096), .Y(n9371) );
  AO21X1 U988 ( .A0(\i_MIPS/n510 ), .A1(\i_MIPS/n166 ), .B0(n10479), .Y(n10488) );
  AOI2BB1X1 U989 ( .A0N(\i_MIPS/IF_ID[25] ), .A1N(\i_MIPS/Sign_Extend[31] ), 
        .B0(n4769), .Y(n10375) );
  INVXL U990 ( .A(n9123), .Y(n7161) );
  OR2X4 U991 ( .A(n5462), .B(net117623), .Y(n3993) );
  INVX1 U992 ( .A(n7687), .Y(n3580) );
  CLKINVX1 U993 ( .A(n6920), .Y(n6849) );
  OAI221XL U994 ( .A0(n345), .A1(n5072), .B0(n2919), .B1(n5068), .C0(n7154), 
        .Y(n3714) );
  OAI221X1 U995 ( .A0(net107210), .A1(n7495), .B0(n7493), .B1(n3774), .C0(
        net117757), .Y(n7499) );
  NAND4X1 U996 ( .A(n6865), .B(n6864), .C(n6863), .D(n6862), .Y(n11401) );
  INVX4 U997 ( .A(n11398), .Y(n10313) );
  INVX3 U998 ( .A(n11397), .Y(n10520) );
  INVX4 U999 ( .A(n11393), .Y(n10625) );
  INVX4 U1000 ( .A(n11384), .Y(n10653) );
  INVX4 U1001 ( .A(n11378), .Y(n10192) );
  CLKINVX6 U1002 ( .A(n11376), .Y(n10744) );
  INVX4 U1003 ( .A(n11433), .Y(n10440) );
  CLKINVX1 U1004 ( .A(n11424), .Y(n10508) );
  OA22XL U1005 ( .A0(n5174), .A1(n696), .B0(n5213), .B1(n2314), .Y(n8256) );
  NAND4X2 U1006 ( .A(n9095), .B(n9094), .C(n9093), .D(n9092), .Y(n11412) );
  OA22XL U1007 ( .A0(n5245), .A1(n600), .B0(n5286), .B1(n2218), .Y(n9094) );
  OA22XL U1008 ( .A0(n5176), .A1(n567), .B0(n5215), .B1(n2319), .Y(n9095) );
  OA22XL U1009 ( .A0(n5396), .A1(n602), .B0(n5440), .B1(n2220), .Y(n7197) );
  INVX4 U1010 ( .A(n11443), .Y(n10759) );
  INVX4 U1011 ( .A(n11495), .Y(n10687) );
  CLKINVX1 U1012 ( .A(n11494), .Y(n10307) );
  BUFX16 U1013 ( .A(n5187), .Y(n5172) );
  OA22XL U1014 ( .A0(n5180), .A1(n620), .B0(n5218), .B1(n2238), .Y(n7344) );
  OA22XL U1015 ( .A0(n5334), .A1(n577), .B0(n5361), .B1(n2195), .Y(n7262) );
  OA22X2 U1016 ( .A0(n5386), .A1(n2089), .B0(n5427), .B1(n463), .Y(n9080) );
  AOI2BB2X1 U1017 ( .B0(n3763), .B1(\D_cache/cache[4][4] ), .A0N(n5357), .A1N(
        n2031), .Y(n9081) );
  INVX3 U1018 ( .A(n11474), .Y(n10186) );
  NAND3X6 U1019 ( .A(ICACHE_addr[26]), .B(ICACHE_addr[25]), .C(n10568), .Y(
        n10576) );
  NAND3X6 U1020 ( .A(ICACHE_addr[14]), .B(ICACHE_addr[13]), .C(n10282), .Y(
        n10292) );
  CLKINVX1 U1021 ( .A(n10488), .Y(n10264) );
  NAND3X2 U1022 ( .A(ICACHE_addr[12]), .B(ICACHE_addr[11]), .C(n10491), .Y(
        n10272) );
  NAND3X6 U1023 ( .A(ICACHE_addr[8]), .B(ICACHE_addr[7]), .C(n10179), .Y(
        n10265) );
  CLKAND2X3 U1024 ( .A(net118217), .B(net105010), .Y(net143547) );
  CLKAND2X8 U1025 ( .A(n9575), .B(n9573), .Y(n3689) );
  NAND4BX1 U1026 ( .AN(n9594), .B(n9593), .C(n9592), .D(n9591), .Y(n9595) );
  NAND4X1 U1027 ( .A(n10953), .B(n10952), .C(n10951), .D(n10950), .Y(n11222)
         );
  NAND4X1 U1028 ( .A(n10859), .B(n10858), .C(n10857), .D(n10856), .Y(n11223)
         );
  NAND4X1 U1029 ( .A(n9904), .B(n9903), .C(n9902), .D(n9901), .Y(n11226) );
  NAND4X1 U1030 ( .A(n9860), .B(n9859), .C(n9858), .D(n9857), .Y(n11227) );
  NAND4X1 U1031 ( .A(n9882), .B(n9881), .C(n9880), .D(n9879), .Y(n11228) );
  NAND4X1 U1032 ( .A(n9838), .B(n9837), .C(n9836), .D(n9835), .Y(n11229) );
  NAND4X1 U1033 ( .A(n10089), .B(n10088), .C(n10087), .D(n10086), .Y(n11230)
         );
  NAND4X1 U1034 ( .A(n10066), .B(n10065), .C(n10064), .D(n10063), .Y(n11234)
         );
  NAND4X1 U1035 ( .A(n9787), .B(n9786), .C(n9785), .D(n9784), .Y(n11238) );
  NAND4X2 U1036 ( .A(n6601), .B(n6600), .C(n6599), .D(n6598), .Y(n11244) );
  NAND4X1 U1037 ( .A(n9623), .B(n9622), .C(n9621), .D(n9620), .Y(n11245) );
  NAND4X1 U1038 ( .A(n9645), .B(n9644), .C(n9643), .D(n9642), .Y(n11246) );
  NAND4X1 U1039 ( .A(n9697), .B(n9696), .C(n9695), .D(n9694), .Y(n11247) );
  NAND4X1 U1040 ( .A(n9675), .B(n9674), .C(n9673), .D(n9672), .Y(n11248) );
  NAND4X1 U1041 ( .A(n6551), .B(n6550), .C(n6549), .D(n6548), .Y(n11250) );
  NAND4X2 U1042 ( .A(n9894), .B(n9893), .C(n9892), .D(n9891), .Y(n11257) );
  NAND4X2 U1043 ( .A(n10115), .B(n10114), .C(n10113), .D(n10112), .Y(n11262)
         );
  NAND4X1 U1044 ( .A(n9777), .B(n9776), .C(n9775), .D(n9774), .Y(n11269) );
  NAND4X1 U1045 ( .A(n10032), .B(n10031), .C(n10030), .D(n10029), .Y(n11274)
         );
  NAND4X1 U1046 ( .A(n9613), .B(n9612), .C(n9611), .D(n9610), .Y(n11276) );
  NAND4X1 U1047 ( .A(n9635), .B(n9634), .C(n9633), .D(n9632), .Y(n11277) );
  NAND4X1 U1048 ( .A(n9687), .B(n9686), .C(n9685), .D(n9684), .Y(n11278) );
  NAND4X1 U1049 ( .A(n6576), .B(n6575), .C(n6574), .D(n6573), .Y(n11280) );
  NAND4X1 U1050 ( .A(n6556), .B(n6555), .C(n6554), .D(n6553), .Y(n11281) );
  NAND4X1 U1051 ( .A(n10877), .B(n10876), .C(n10875), .D(n10874), .Y(n11282)
         );
  NAND4X1 U1052 ( .A(n10948), .B(n10947), .C(n10946), .D(n10945), .Y(n11284)
         );
  NAND4X1 U1053 ( .A(n10854), .B(n10853), .C(n10852), .D(n10851), .Y(n11285)
         );
  NAND4X1 U1054 ( .A(n9714), .B(n9713), .C(n9712), .D(n9711), .Y(n11286) );
  NAND4X1 U1055 ( .A(n9899), .B(n9898), .C(n9897), .D(n9896), .Y(n11288) );
  NAND4X1 U1056 ( .A(n9855), .B(n9854), .C(n9853), .D(n9852), .Y(n11289) );
  NAND4X1 U1057 ( .A(n9877), .B(n9876), .C(n9875), .D(n9874), .Y(n11290) );
  NAND4X1 U1058 ( .A(n9833), .B(n9832), .C(n9831), .D(n9830), .Y(n11291) );
  NAND4X1 U1059 ( .A(n10084), .B(n10083), .C(n10082), .D(n10081), .Y(n11292)
         );
  NAND4X1 U1060 ( .A(n10120), .B(n10119), .C(n10118), .D(n10117), .Y(n11293)
         );
  NAND4X1 U1061 ( .A(n10218), .B(n10217), .C(n10216), .D(n10215), .Y(n11294)
         );
  NAND4X1 U1062 ( .A(n10240), .B(n10239), .C(n10238), .D(n10237), .Y(n11295)
         );
  NAND4X1 U1063 ( .A(n10061), .B(n10060), .C(n10059), .D(n10058), .Y(n11296)
         );
  NAND4X1 U1064 ( .A(n9782), .B(n9781), .C(n9780), .D(n9779), .Y(n11300) );
  NAND4X1 U1065 ( .A(n10037), .B(n10036), .C(n10035), .D(n10034), .Y(n11305)
         );
  NAND4X2 U1066 ( .A(n6596), .B(n6595), .C(n6594), .D(n6593), .Y(n11306) );
  NAND4X1 U1067 ( .A(n9618), .B(n9617), .C(n9616), .D(n9615), .Y(n11307) );
  NAND4X1 U1068 ( .A(n9640), .B(n9639), .C(n9638), .D(n9637), .Y(n11308) );
  NAND4X1 U1069 ( .A(n9692), .B(n9691), .C(n9690), .D(n9689), .Y(n11309) );
  NAND4X1 U1070 ( .A(n9670), .B(n9669), .C(n9668), .D(n9667), .Y(n11310) );
  NAND4X1 U1071 ( .A(n6581), .B(n6580), .C(n6579), .D(n6578), .Y(n11311) );
  OA22X2 U1072 ( .A0(n5918), .A1(n2078), .B0(n5876), .B1(n453), .Y(n11151) );
  OA22X2 U1073 ( .A0(n5831), .A1(n2062), .B0(n5786), .B1(n437), .Y(n11152) );
  OA22X2 U1074 ( .A0(n5919), .A1(n2093), .B0(n5877), .B1(n467), .Y(n11156) );
  OA22X2 U1075 ( .A0(n5918), .A1(n2077), .B0(n5876), .B1(n452), .Y(n11136) );
  NAND4X4 U1076 ( .A(n11149), .B(n11148), .C(n11147), .D(n11146), .Y(n11359)
         );
  OA22X2 U1077 ( .A0(n5918), .A1(n2079), .B0(n5876), .B1(n454), .Y(n11146) );
  OA22X2 U1078 ( .A0(n5652), .A1(n2085), .B0(n5608), .B1(n459), .Y(n11149) );
  NAND4X6 U1079 ( .A(n4664), .B(n6381), .C(n6380), .D(n6379), .Y(n11364) );
  AOI2BB2X2 U1080 ( .B0(n4832), .B1(\I_cache/cache[5][146] ), .A0N(n5807), 
        .A1N(n2927), .Y(n6363) );
  OA22X2 U1081 ( .A0(n5654), .A1(n2066), .B0(n5608), .B1(n441), .Y(n11191) );
  AOI2BB2X2 U1082 ( .B0(n4832), .B1(\I_cache/cache[5][150] ), .A0N(n5807), 
        .A1N(n2926), .Y(n6367) );
  NAND4X6 U1083 ( .A(n4665), .B(n6378), .C(n6377), .D(n6376), .Y(n11370) );
  OA22X2 U1084 ( .A0(n5718), .A1(n2972), .B0(n5703), .B1(n1294), .Y(n6378) );
  AOI2BB2X2 U1085 ( .B0(n4829), .B1(\I_cache/cache[5][151] ), .A0N(n5838), 
        .A1N(n2923), .Y(n6377) );
  OA22X2 U1086 ( .A0(n5929), .A1(n3012), .B0(n5878), .B1(n530), .Y(n6370) );
  AOI2BB2X2 U1087 ( .B0(n4831), .B1(\I_cache/cache[5][152] ), .A0N(n5833), 
        .A1N(n2925), .Y(n6371) );
  NAND4X2 U1088 ( .A(n9176), .B(n9175), .C(n9174), .D(n9173), .Y(n11379) );
  OA22XL U1089 ( .A0(n5180), .A1(n616), .B0(n5218), .B1(n2234), .Y(n7352) );
  OA22XL U1090 ( .A0(n5391), .A1(n2116), .B0(n5434), .B1(n490), .Y(n7996) );
  NAND4X2 U1091 ( .A(n8607), .B(n8606), .C(n8605), .D(n8604), .Y(n11394) );
  NAND4X2 U1092 ( .A(n8342), .B(n8341), .C(n8340), .D(n8339), .Y(n11395) );
  OA22XL U1093 ( .A0(n5181), .A1(n674), .B0(n5218), .B1(n2292), .Y(n7072) );
  OA22XL U1094 ( .A0(n5398), .A1(n673), .B0(n5442), .B1(n2291), .Y(n7069) );
  INVX3 U1095 ( .A(n11401), .Y(n10437) );
  NAND4X2 U1096 ( .A(n8832), .B(n8831), .C(n8830), .D(n8829), .Y(n11424) );
  OA22XL U1097 ( .A0(n5175), .A1(n640), .B0(n5214), .B1(n2257), .Y(n8832) );
  NAND4X2 U1098 ( .A(n8611), .B(n8610), .C(n8609), .D(n8608), .Y(n11426) );
  OA22XL U1099 ( .A0(n5387), .A1(n604), .B0(n5428), .B1(n2222), .Y(n8932) );
  OA22X2 U1100 ( .A0(n5246), .A1(n2132), .B0(n5296), .B1(n507), .Y(n8934) );
  OA22XL U1101 ( .A0(n5177), .A1(n651), .B0(n5216), .B1(n2268), .Y(n9419) );
  OA22X2 U1102 ( .A0(n5377), .A1(n2110), .B0(n5422), .B1(n484), .Y(n9416) );
  OA22X1 U1103 ( .A0(n5248), .A1(n2162), .B0(n5288), .B1(n543), .Y(n8747) );
  OA22X2 U1104 ( .A0(n5388), .A1(n2166), .B0(n5430), .B1(n547), .Y(n8745) );
  OA22XL U1105 ( .A0(n5181), .A1(n648), .B0(n5218), .B1(n2265), .Y(n7192) );
  OA22XL U1106 ( .A0(n5396), .A1(n647), .B0(n5440), .B1(n2264), .Y(n7189) );
  OA22XL U1107 ( .A0(n5177), .A1(n676), .B0(n5216), .B1(n2294), .Y(n9353) );
  OA22X2 U1108 ( .A0(n5180), .A1(n2151), .B0(n5218), .B1(n526), .Y(n7348) );
  OA22XL U1109 ( .A0(n5252), .A1(n2091), .B0(n5292), .B1(n465), .Y(n8167) );
  OA22XL U1110 ( .A0(n5329), .A1(n584), .B0(n5354), .B1(n2202), .Y(n8166) );
  OA22X1 U1111 ( .A0(n5375), .A1(n614), .B0(n5433), .B1(n2232), .Y(n8165) );
  OA22X2 U1112 ( .A0(n5178), .A1(n2168), .B0(n5217), .B1(n549), .Y(n8078) );
  OA22X2 U1113 ( .A0(n5253), .A1(n2163), .B0(n5293), .B1(n544), .Y(n8077) );
  OA22XL U1114 ( .A0(n5253), .A1(n2164), .B0(n5293), .B1(n545), .Y(n7994) );
  OA22XL U1115 ( .A0(n5255), .A1(n2072), .B0(n5295), .B1(n447), .Y(n7803) );
  OA22X2 U1116 ( .A0(n5390), .A1(n2157), .B0(n5432), .B1(n538), .Y(n8335) );
  OA22X2 U1117 ( .A0(n5330), .A1(n2156), .B0(n5354), .B1(n537), .Y(n8426) );
  NAND4X4 U1118 ( .A(n8927), .B(n8926), .C(n8925), .D(n8924), .Y(n11461) );
  OA22XL U1119 ( .A0(n5176), .A1(n2148), .B0(n5215), .B1(n523), .Y(n8927) );
  OA22XL U1120 ( .A0(n5247), .A1(n613), .B0(n5287), .B1(n2231), .Y(n8926) );
  OA22X1 U1121 ( .A0(n5332), .A1(n622), .B0(n5357), .B1(n2240), .Y(n8925) );
  OA22XL U1122 ( .A0(n5181), .A1(n667), .B0(n5218), .B1(n2285), .Y(n7068) );
  OA22X1 U1123 ( .A0(n5398), .A1(n666), .B0(n5442), .B1(n2284), .Y(n7065) );
  OA22XL U1124 ( .A0(n5179), .A1(n682), .B0(n5213), .B1(n2300), .Y(n7708) );
  OA22XL U1125 ( .A0(n5398), .A1(n672), .B0(n5442), .B1(n2290), .Y(n6969) );
  OA22XL U1126 ( .A0(n5177), .A1(n656), .B0(n5216), .B1(n2273), .Y(n9411) );
  OA22X1 U1127 ( .A0(n5379), .A1(n654), .B0(n5422), .B1(n2271), .Y(n9408) );
  OA22XL U1128 ( .A0(n5178), .A1(n717), .B0(n5217), .B1(n2339), .Y(n9524) );
  OA22XL U1129 ( .A0(n5388), .A1(n2124), .B0(n5430), .B1(n499), .Y(n8741) );
  NAND4X2 U1130 ( .A(n9007), .B(n9006), .C(n9005), .D(n9004), .Y(n11473) );
  OA22X2 U1131 ( .A0(n5246), .A1(n2135), .B0(n5298), .B1(n510), .Y(n9006) );
  NAND4X2 U1132 ( .A(n9168), .B(n9167), .C(n9166), .D(n9165), .Y(n11475) );
  OA22XL U1133 ( .A0(n5176), .A1(n663), .B0(n5215), .B1(n2281), .Y(n9168) );
  INVX6 U1134 ( .A(n11479), .Y(n10674) );
  INVX3 U1135 ( .A(n11481), .Y(n10606) );
  NAND4X2 U1136 ( .A(n7109), .B(n7108), .C(n7107), .D(n7106), .Y(n11487) );
  AOI2BB2XL U1137 ( .B0(n3763), .B1(\D_cache/cache[4][18] ), .A0N(n5356), 
        .A1N(n2032), .Y(n8597) );
  OA22X2 U1138 ( .A0(n5250), .A1(n2160), .B0(n5290), .B1(n541), .Y(n8423) );
  NAND4X2 U1139 ( .A(n7906), .B(n7905), .C(n7904), .D(n7903), .Y(n11494) );
  OA22XL U1140 ( .A0(n5178), .A1(n637), .B0(n5217), .B1(n2254), .Y(n7906) );
  OA22XL U1141 ( .A0(n5331), .A1(n626), .B0(n5359), .B1(n2244), .Y(n7904) );
  INVX1 U1142 ( .A(n11496), .Y(n10417) );
  OA22XL U1143 ( .A0(n5180), .A1(n658), .B0(n5218), .B1(n2275), .Y(n7443) );
  OA22X1 U1144 ( .A0(n5395), .A1(n657), .B0(n5439), .B1(n2274), .Y(n7440) );
  OA22XL U1145 ( .A0(n5178), .A1(n635), .B0(n5217), .B1(n2252), .Y(n9520) );
  OA22XL U1146 ( .A0(n5376), .A1(n633), .B0(n5421), .B1(n2250), .Y(n9517) );
  INVX8 U1147 ( .A(n5041), .Y(n5043) );
  INVX8 U1148 ( .A(n11508), .Y(n11534) );
  OR2X6 U1149 ( .A(net108640), .B(net117709), .Y(n3835) );
  NAND2XL U1150 ( .A(net139864), .B(net105531), .Y(n10646) );
  NAND4X1 U1151 ( .A(n10042), .B(n10041), .C(n10040), .D(n10039), .Y(n11243)
         );
  NAND4X1 U1152 ( .A(n9665), .B(n9664), .C(n9663), .D(n9662), .Y(n11279) );
  NAND4X1 U1153 ( .A(n9719), .B(n9718), .C(n9717), .D(n9716), .Y(n11224) );
  NAND4X1 U1154 ( .A(n10223), .B(n10222), .C(n10221), .D(n10220), .Y(n11232)
         );
  NAND4X1 U1155 ( .A(n10125), .B(n10124), .C(n10123), .D(n10122), .Y(n11231)
         );
  CLKINVX1 U1156 ( .A(n11220), .Y(n3806) );
  NAND4X1 U1157 ( .A(n6586), .B(n6585), .C(n6584), .D(n6583), .Y(n11249) );
  NAND4X1 U1158 ( .A(n6591), .B(n6590), .C(n6589), .D(n6588), .Y(n11275) );
  NAND4X1 U1159 ( .A(n10245), .B(n10244), .C(n10243), .D(n10242), .Y(n11233)
         );
  NAND2XL U1160 ( .A(n3004), .B(net105479), .Y(n10416) );
  AO21X1 U1161 ( .A0(\i_MIPS/n516 ), .A1(\i_MIPS/n160 ), .B0(n4747), .Y(n10153) );
  NAND2XL U1162 ( .A(net139765), .B(net105783), .Y(n10528) );
  XOR2X1 U1163 ( .A(n10492), .B(ICACHE_addr[12]), .Y(n10496) );
  XOR2X1 U1164 ( .A(n10342), .B(ICACHE_addr[20]), .Y(n10346) );
  XOR2X1 U1165 ( .A(n10365), .B(ICACHE_addr[22]), .Y(n10369) );
  AO21X1 U1166 ( .A0(\i_MIPS/n169 ), .A1(\i_MIPS/n507 ), .B0(n4816), .Y(n10289) );
  BUFX20 U1167 ( .A(net115811), .Y(net115799) );
  NOR2BX2 U1168 ( .AN(\i_MIPS/IF_ID[10] ), .B(\i_MIPS/n513 ), .Y(n4807) );
  BUFX16 U1169 ( .A(n12977), .Y(DCACHE_addr[6]) );
  BUFX16 U1170 ( .A(n12965), .Y(DCACHE_addr[18]) );
  OAI221X1 U1171 ( .A0(n9934), .A1(net143858), .B0(\i_MIPS/n515 ), .B1(
        net115791), .C0(n9933), .Y(\i_MIPS/N55 ) );
  AND2X2 U1172 ( .A(net104172), .B(n11256), .Y(n4447) );
  INVX6 U1173 ( .A(n11362), .Y(n11216) );
  CLKAND2X8 U1174 ( .A(n4378), .B(n4379), .Y(n4367) );
  CLKINVX1 U1175 ( .A(net108004), .Y(net108847) );
  INVX8 U1176 ( .A(net108874), .Y(net112449) );
  AND2X6 U1177 ( .A(n7314), .B(n8134), .Y(n4690) );
  CLKAND2X6 U1178 ( .A(n9302), .B(n9308), .Y(n4692) );
  INVX1 U1179 ( .A(n4776), .Y(n3746) );
  OR2X6 U1180 ( .A(n6495), .B(n3019), .Y(n4403) );
  NAND2X2 U1181 ( .A(n6495), .B(n3019), .Y(n4402) );
  NAND2X6 U1182 ( .A(n11026), .B(n3005), .Y(n6490) );
  NAND2X4 U1183 ( .A(n11037), .B(n11036), .Y(n6455) );
  CLKBUFX3 U1184 ( .A(net134680), .Y(net118315) );
  CLKINVX1 U1185 ( .A(net108151), .Y(net108005) );
  INVX6 U1186 ( .A(n3704), .Y(n3705) );
  CLKINVX6 U1187 ( .A(n3682), .Y(n6646) );
  INVX6 U1188 ( .A(n3621), .Y(n3622) );
  NAND2X2 U1189 ( .A(n4727), .B(n7487), .Y(n7767) );
  INVX3 U1190 ( .A(n3850), .Y(n3851) );
  INVXL U1191 ( .A(n8120), .Y(n8660) );
  NAND2XL U1192 ( .A(n4675), .B(n6776), .Y(net139718) );
  NAND2X1 U1193 ( .A(\i_MIPS/ALU/N303 ), .B(n9556), .Y(n11106) );
  NAND2X1 U1194 ( .A(n9555), .B(\i_MIPS/n270 ), .Y(n11108) );
  CLKAND2X6 U1195 ( .A(n4814), .B(n4785), .Y(net134679) );
  AND2X4 U1196 ( .A(n254), .B(\i_MIPS/n500 ), .Y(n4675) );
  NAND2X2 U1197 ( .A(n6724), .B(n345), .Y(n8886) );
  NAND2X2 U1198 ( .A(net109965), .B(n8291), .Y(n8210) );
  CLKINVX1 U1199 ( .A(n3764), .Y(net110423) );
  CLKINVX1 U1200 ( .A(n7765), .Y(n3708) );
  AND2X1 U1201 ( .A(n4787), .B(n4722), .Y(n4759) );
  NAND4X4 U1202 ( .A(n4003), .B(n4004), .C(n4005), .D(n4006), .Y(n3793) );
  OA22X1 U1203 ( .A0(\i_MIPS/Register/register[17][18] ), .A1(net118453), .B0(
        \i_MIPS/Register/register[25][18] ), .B1(net118477), .Y(n8587) );
  OA22X1 U1204 ( .A0(\i_MIPS/Register/register[22][18] ), .A1(net117681), .B0(
        \i_MIPS/Register/register[30][18] ), .B1(net117697), .Y(n8588) );
  CLKINVX1 U1205 ( .A(n8666), .Y(n8647) );
  INVX3 U1206 ( .A(n7224), .Y(n7225) );
  NAND2X6 U1207 ( .A(n4395), .B(n4396), .Y(n7222) );
  CLKINVX4 U1208 ( .A(net118487), .Y(net118473) );
  INVX4 U1209 ( .A(net118367), .Y(net118353) );
  INVX4 U1210 ( .A(net118439), .Y(net118425) );
  AND2X2 U1211 ( .A(n5074), .B(n2937), .Y(n4745) );
  INVX3 U1212 ( .A(net108003), .Y(net108148) );
  NAND2X1 U1213 ( .A(n134), .B(n2961), .Y(n6928) );
  CLKBUFX3 U1214 ( .A(net134686), .Y(net118415) );
  CLKBUFX3 U1215 ( .A(net134686), .Y(net118413) );
  CLKINVX1 U1216 ( .A(n7424), .Y(n6913) );
  NAND2X2 U1217 ( .A(n6948), .B(n253), .Y(n11096) );
  NAND2X4 U1218 ( .A(n6668), .B(n344), .Y(n11101) );
  BUFX4 U1219 ( .A(n6823), .Y(n144) );
  CLKINVX1 U1220 ( .A(n6937), .Y(n6830) );
  AO21X1 U1221 ( .A0(n8966), .A1(n8291), .B0(n4724), .Y(n7941) );
  NAND3BX1 U1222 ( .AN(n8639), .B(net110129), .C(n7949), .Y(n7955) );
  INVX6 U1223 ( .A(n6716), .Y(n8780) );
  CLKINVX1 U1224 ( .A(n7784), .Y(n7420) );
  CLKMX2X2 U1225 ( .A(n8873), .B(n8865), .S0(net114065), .Y(n8043) );
  NOR2X2 U1226 ( .A(n8028), .B(n3774), .Y(n3780) );
  CLKINVX4 U1227 ( .A(n6725), .Y(n6685) );
  OA22X2 U1228 ( .A0(n3861), .A1(n5064), .B0(n253), .B1(n5058), .Y(n7152) );
  NAND2BX2 U1229 ( .AN(\i_MIPS/PC/n8 ), .B(n4801), .Y(n4681) );
  BUFX6 U1230 ( .A(n9809), .Y(n5454) );
  AND2X2 U1231 ( .A(\i_MIPS/n504 ), .B(\i_MIPS/n505 ), .Y(n4722) );
  CLKMX2X4 U1232 ( .A(net108284), .B(net107404), .S0(n3669), .Y(net108306) );
  MXI2X1 U1233 ( .A(n3873), .B(net134414), .S0(\i_MIPS/ID_EX[74] ), .Y(n6650)
         );
  NAND2X1 U1234 ( .A(n5075), .B(\i_MIPS/ALUin1[8] ), .Y(n8979) );
  AND2X2 U1235 ( .A(n5075), .B(\i_MIPS/ALUin1[26] ), .Y(n4794) );
  NAND2X1 U1236 ( .A(net108869), .B(net108873), .Y(net109513) );
  NOR2BX2 U1237 ( .AN(n5066), .B(\i_MIPS/n299 ), .Y(n4799) );
  OA22X1 U1238 ( .A0(\i_MIPS/Register/register[1][15] ), .A1(net118453), .B0(
        \i_MIPS/Register/register[9][15] ), .B1(net118479), .Y(n4297) );
  OR3X6 U1239 ( .A(n149), .B(n8119), .C(n8118), .Y(n4401) );
  INVX3 U1240 ( .A(n8116), .Y(n8118) );
  AND2X4 U1241 ( .A(n5065), .B(\i_MIPS/ALUin1[17] ), .Y(n4818) );
  AND2X4 U1242 ( .A(\i_MIPS/n497 ), .B(n7739), .Y(n4720) );
  AND2X4 U1243 ( .A(\i_MIPS/n499 ), .B(\i_MIPS/n500 ), .Y(n4723) );
  NAND2X4 U1244 ( .A(n3004), .B(net105479), .Y(n3828) );
  NAND2X4 U1245 ( .A(net139777), .B(net105764), .Y(n4336) );
  AND2X2 U1246 ( .A(net49779), .B(net118581), .Y(n3773) );
  NAND2X4 U1247 ( .A(net112414), .B(\i_MIPS/n297 ), .Y(n9302) );
  NOR4X4 U1248 ( .A(n6385), .B(n6384), .C(n6383), .D(n6382), .Y(n6386) );
  INVX6 U1249 ( .A(n3965), .Y(n3966) );
  BUFX3 U1250 ( .A(n5267), .Y(n5262) );
  OAI221XL U1251 ( .A0(\i_MIPS/Register/register[18][23] ), .A1(net117635), 
        .B0(\i_MIPS/Register/register[26][23] ), .B1(net117653), .C0(n7092), 
        .Y(n7095) );
  OAI221XL U1252 ( .A0(\i_MIPS/Register/register[18][19] ), .A1(net117639), 
        .B0(\i_MIPS/Register/register[26][19] ), .B1(net117659), .C0(n8324), 
        .Y(n8327) );
  OA22X1 U1253 ( .A0(\i_MIPS/Register/register[22][19] ), .A1(net117681), .B0(
        \i_MIPS/Register/register[30][19] ), .B1(net117695), .Y(n8324) );
  CLKMX2X2 U1254 ( .A(n7675), .B(net107992), .S0(net114065), .Y(n7038) );
  OAI221XL U1255 ( .A0(\i_MIPS/Register/register[18][16] ), .A1(net117641), 
        .B0(\i_MIPS/Register/register[26][16] ), .B1(net117659), .C0(n8810), 
        .Y(n8813) );
  OAI221XL U1256 ( .A0(\i_MIPS/Register/register[18][22] ), .A1(net117639), 
        .B0(\i_MIPS/Register/register[26][22] ), .B1(net117657), .C0(n7934), 
        .Y(n7937) );
  CLKINVX6 U1257 ( .A(n7025), .Y(n7864) );
  INVX4 U1258 ( .A(n8880), .Y(n7856) );
  NAND2X1 U1259 ( .A(\i_MIPS/ALUin1[21] ), .B(n6689), .Y(n8885) );
  NAND2X2 U1260 ( .A(n6725), .B(n2949), .Y(n7861) );
  CLKMX2X2 U1261 ( .A(n7788), .B(n7787), .S0(net114065), .Y(n7233) );
  CLKMX2X2 U1262 ( .A(n7480), .B(n7422), .S0(net114065), .Y(n7789) );
  INVX1 U1263 ( .A(n7949), .Y(n7777) );
  AO22X1 U1264 ( .A0(n5156), .A1(n427), .B0(n5153), .B1(n2054), .Y(n8540) );
  OA22X1 U1265 ( .A0(\i_MIPS/Register/register[6][18] ), .A1(n5083), .B0(
        \i_MIPS/Register/register[14][18] ), .B1(n5079), .Y(n8612) );
  OA22X1 U1266 ( .A0(\i_MIPS/Register/register[22][18] ), .A1(n5083), .B0(
        \i_MIPS/Register/register[30][18] ), .B1(n5079), .Y(n8621) );
  NAND2X6 U1267 ( .A(n4788), .B(n4784), .Y(n7887) );
  NOR4X1 U1268 ( .A(n8763), .B(n8762), .C(n8761), .D(n8760), .Y(n8764) );
  AO22X1 U1269 ( .A0(n5154), .A1(n421), .B0(n5153), .B1(n2048), .Y(n8760) );
  OA22XL U1270 ( .A0(\i_MIPS/Register/register[6][0] ), .A1(n5083), .B0(
        \i_MIPS/Register/register[14][0] ), .B1(n5079), .Y(n8759) );
  AO22X1 U1271 ( .A0(n5158), .A1(n420), .B0(n5153), .B1(n2047), .Y(n8769) );
  OAI221XL U1272 ( .A0(\i_MIPS/Register/register[18][0] ), .A1(n5091), .B0(
        \i_MIPS/Register/register[26][0] ), .B1(n4669), .C0(n8768), .Y(n8776)
         );
  NOR4X1 U1273 ( .A(n8583), .B(n8582), .C(n8581), .D(n8580), .Y(n8594) );
  OAI221XL U1274 ( .A0(\i_MIPS/Register/register[2][18] ), .A1(net117641), 
        .B0(\i_MIPS/Register/register[10][18] ), .B1(net117659), .C0(n8579), 
        .Y(n8582) );
  AO22X1 U1275 ( .A0(net118273), .A1(n416), .B0(net118291), .B1(n2043), .Y(
        n8581) );
  NOR4X1 U1276 ( .A(n8592), .B(n8591), .C(n8590), .D(n8589), .Y(n8593) );
  OAI221XL U1277 ( .A0(\i_MIPS/Register/register[18][18] ), .A1(net117641), 
        .B0(\i_MIPS/Register/register[26][18] ), .B1(net117659), .C0(n8588), 
        .Y(n8591) );
  AO22X1 U1278 ( .A0(net118273), .A1(n415), .B0(net118291), .B1(n2042), .Y(
        n8590) );
  NAND4X1 U1279 ( .A(n8587), .B(n8586), .C(n8585), .D(n8584), .Y(n8592) );
  INVX6 U1280 ( .A(n8632), .Y(n6674) );
  OA21XL U1281 ( .A0(n9428), .A1(n9425), .B0(n9424), .Y(n9426) );
  CLKINVX1 U1282 ( .A(n7790), .Y(n9453) );
  OAI221XL U1283 ( .A0(\i_MIPS/ALUin1[23] ), .A1(n5071), .B0(
        \i_MIPS/ALUin1[24] ), .B1(n5067), .C0(n7410), .Y(n7411) );
  OAI221XL U1284 ( .A0(\i_MIPS/Register/register[18][29] ), .A1(net117635), 
        .B0(\i_MIPS/Register/register[26][29] ), .B1(net117653), .C0(n6996), 
        .Y(n6999) );
  NAND4X2 U1285 ( .A(n11583), .B(n3726), .C(net108787), .D(n4741), .Y(n8707)
         );
  AOI31X1 U1286 ( .A0(n9204), .A1(n8687), .A2(n8686), .B0(n8685), .Y(n8691) );
  AOI21XL U1287 ( .A0(n9203), .A1(n9223), .B0(n8680), .Y(n8686) );
  NAND2X2 U1288 ( .A(\i_MIPS/ALUin1[22] ), .B(n6725), .Y(n8695) );
  AOI211X1 U1289 ( .A0(n8642), .A1(n8641), .B0(n8640), .C0(n8690), .Y(n8677)
         );
  BUFX4 U1290 ( .A(n5113), .Y(n5118) );
  OAI2BB1X2 U1291 ( .A0N(n5065), .A1N(\i_MIPS/ALU/N303 ), .B0(n9447), .Y(n7790) );
  CLKINVX1 U1292 ( .A(n7789), .Y(n7850) );
  OAI221XL U1293 ( .A0(\i_MIPS/Register/register[18][2] ), .A1(n5089), .B0(
        \i_MIPS/Register/register[26][2] ), .B1(n5084), .C0(n7210), .Y(n7218)
         );
  OAI221XL U1294 ( .A0(\i_MIPS/Register/register[2][2] ), .A1(n5089), .B0(
        \i_MIPS/Register/register[10][2] ), .B1(n5084), .C0(n7201), .Y(n7209)
         );
  NAND2X2 U1295 ( .A(n8866), .B(n3674), .Y(n9317) );
  AO22X1 U1296 ( .A0(net118237), .A1(n551), .B0(net118255), .B1(n2170), .Y(
        n8414) );
  OAI221XL U1297 ( .A0(\i_MIPS/Register/register[18][20] ), .A1(net117641), 
        .B0(\i_MIPS/Register/register[26][20] ), .B1(net117659), .C0(n8413), 
        .Y(n8416) );
  OA22X1 U1298 ( .A0(\i_MIPS/Register/register[22][20] ), .A1(net117681), .B0(
        \i_MIPS/Register/register[30][20] ), .B1(net117697), .Y(n8413) );
  NAND4X1 U1299 ( .A(n8403), .B(n8402), .C(n8401), .D(n8400), .Y(n8408) );
  AO22X1 U1300 ( .A0(net118237), .A1(n550), .B0(net118255), .B1(n2169), .Y(
        n8405) );
  OAI221XL U1301 ( .A0(\i_MIPS/Register/register[2][20] ), .A1(net117639), 
        .B0(\i_MIPS/Register/register[10][20] ), .B1(net117659), .C0(n8404), 
        .Y(n8407) );
  AO22X1 U1302 ( .A0(net118273), .A1(n418), .B0(net118291), .B1(n2045), .Y(
        n8406) );
  OAI221XL U1303 ( .A0(\i_MIPS/Register/register[18][10] ), .A1(net117637), 
        .B0(\i_MIPS/Register/register[26][10] ), .B1(net117655), .C0(n7518), 
        .Y(n7521) );
  NOR4X1 U1304 ( .A(n8010), .B(n8009), .C(n8008), .D(n8007), .Y(n8011) );
  NOR4X1 U1305 ( .A(n8019), .B(n8018), .C(n8017), .D(n8016), .Y(n8020) );
  AO22X1 U1306 ( .A0(n5157), .A1(n553), .B0(n5153), .B1(n2172), .Y(n8016) );
  AND4X1 U1307 ( .A(n1988), .B(n4833), .C(\i_MIPS/forward_unit/n25 ), .D(n223), 
        .Y(\i_MIPS/forward_unit/n10 ) );
  INVX3 U1308 ( .A(n5097), .Y(n5095) );
  OA22X1 U1309 ( .A0(\i_MIPS/Register/register[20][17] ), .A1(n5099), .B0(
        \i_MIPS/Register/register[28][17] ), .B1(n5096), .Y(n9289) );
  NOR4X2 U1310 ( .A(n9277), .B(n9276), .C(n9275), .D(n9274), .Y(n9278) );
  OA22X1 U1311 ( .A0(\i_MIPS/Register/register[4][17] ), .A1(n5101), .B0(
        \i_MIPS/Register/register[12][17] ), .B1(n5096), .Y(n9280) );
  NOR4X1 U1312 ( .A(n8951), .B(n8950), .C(n8949), .D(n8948), .Y(n8952) );
  AO22X1 U1313 ( .A0(n5155), .A1(n419), .B0(n5153), .B1(n2046), .Y(n8939) );
  OA22X1 U1314 ( .A0(\i_MIPS/Register/register[20][5] ), .A1(n5099), .B0(
        \i_MIPS/Register/register[28][5] ), .B1(n5096), .Y(n9380) );
  NAND4X1 U1315 ( .A(n9157), .B(n9156), .C(n9155), .D(n9154), .Y(n9162) );
  NAND4X1 U1316 ( .A(n9148), .B(n9147), .C(n9146), .D(n9145), .Y(n9153) );
  OAI221XL U1317 ( .A0(\i_MIPS/Register/register[2][3] ), .A1(net117643), .B0(
        \i_MIPS/Register/register[10][3] ), .B1(net117661), .C0(n9149), .Y(
        n9152) );
  NOR2BX2 U1318 ( .AN(n5069), .B(\i_MIPS/n297 ), .Y(n4795) );
  NOR2BX2 U1319 ( .AN(n5074), .B(\i_MIPS/n296 ), .Y(n4792) );
  NAND2X1 U1320 ( .A(\i_MIPS/ALUin1[2] ), .B(net112418), .Y(n7145) );
  INVX12 U1321 ( .A(net112393), .Y(net108787) );
  INVX12 U1322 ( .A(n8793), .Y(n7676) );
  CLKAND2X3 U1323 ( .A(n8963), .B(n3748), .Y(n4688) );
  NAND2X1 U1324 ( .A(n144), .B(n2184), .Y(n6919) );
  CLKAND2X8 U1325 ( .A(n8550), .B(n8288), .Y(n4706) );
  NAND2X2 U1326 ( .A(n6687), .B(n336), .Y(n8397) );
  CLKINVX1 U1327 ( .A(n7955), .Y(n7950) );
  CLKINVX1 U1328 ( .A(n9314), .Y(n8968) );
  CLKINVX1 U1329 ( .A(n8043), .Y(n9200) );
  CLKINVX1 U1330 ( .A(n8037), .Y(n8038) );
  AOI32X1 U1331 ( .A0(net111262), .A1(n7102), .A2(n4718), .B0(n7039), .B1(
        net107404), .Y(n7046) );
  NAND2BX2 U1332 ( .AN(n8874), .B(net110602), .Y(n7043) );
  OAI222X1 U1333 ( .A0(net135772), .A1(n9553), .B0(n9551), .B1(n5049), .C0(
        n7035), .C1(net117757), .Y(n7052) );
  INVX4 U1334 ( .A(n6814), .Y(n7026) );
  CLKINVX1 U1335 ( .A(n8557), .Y(n8561) );
  CLKINVX1 U1336 ( .A(n8558), .Y(n8559) );
  NAND2X4 U1337 ( .A(n8291), .B(n3748), .Y(n9210) );
  NAND3X2 U1338 ( .A(n8573), .B(n8569), .C(n3950), .Y(n3790) );
  OA22X2 U1339 ( .A0(n5626), .A1(n2582), .B0(n5612), .B1(n1076), .Y(n4663) );
  NAND2X1 U1340 ( .A(n4796), .B(n10980), .Y(n11050) );
  CLKAND2X3 U1341 ( .A(n9945), .B(n4725), .Y(n3658) );
  OA22X2 U1342 ( .A0(n5256), .A1(n2096), .B0(n5299), .B1(n470), .Y(n7263) );
  OA22X2 U1343 ( .A0(n5929), .A1(n2939), .B0(n5879), .B1(n1305), .Y(n6359) );
  BUFX4 U1344 ( .A(n5133), .Y(n5137) );
  BUFX4 U1345 ( .A(n5121), .Y(n5124) );
  XOR2XL U1346 ( .A(n6754), .B(net105477), .Y(n6641) );
  XOR2XL U1347 ( .A(n6753), .B(\i_MIPS/jump_addr[18] ), .Y(n6640) );
  CLKBUFX8 U1348 ( .A(n5113), .Y(n5117) );
  BUFX4 U1349 ( .A(n5078), .Y(n5076) );
  BUFX4 U1350 ( .A(n5121), .Y(n5122) );
  BUFX4 U1351 ( .A(n4660), .Y(n5079) );
  CLKBUFX3 U1352 ( .A(n11073), .Y(n5565) );
  BUFX6 U1353 ( .A(n5661), .Y(n5660) );
  OAI211XL U1354 ( .A0(n5051), .A1(n9136), .B0(n8980), .C0(n8979), .Y(
        net107665) );
  NAND4BX2 U1355 ( .AN(n3887), .B(n6518), .C(n6517), .D(n6516), .Y(n6524) );
  NAND2BX1 U1356 ( .AN(n5447), .B(\D_cache/cache[7][154] ), .Y(n6516) );
  OAI221XL U1357 ( .A0(\i_MIPS/Register/register[2][0] ), .A1(net117641), .B0(
        \i_MIPS/Register/register[10][0] ), .B1(net117659), .C0(n8725), .Y(
        n8728) );
  OAI221XL U1358 ( .A0(\i_MIPS/Register/register[18][0] ), .A1(net117641), 
        .B0(\i_MIPS/Register/register[26][0] ), .B1(net117659), .C0(n8734), 
        .Y(n8737) );
  NAND3BX1 U1359 ( .AN(n4746), .B(n7104), .C(n7103), .Y(net109172) );
  CLKMX2X2 U1360 ( .A(n8480), .B(net109172), .S0(net114065), .Y(n9134) );
  NAND2X4 U1361 ( .A(n6695), .B(n3744), .Y(net109176) );
  OA22X1 U1362 ( .A0(\i_MIPS/Register/register[17][15] ), .A1(net118453), .B0(
        \i_MIPS/Register/register[25][15] ), .B1(net118479), .Y(n4288) );
  OAI221XL U1363 ( .A0(\i_MIPS/Register/register[18][15] ), .A1(net117635), 
        .B0(\i_MIPS/Register/register[26][15] ), .B1(net117653), .C0(n4287), 
        .Y(n4284) );
  NOR4X2 U1364 ( .A(n9067), .B(n9066), .C(n9065), .D(n9064), .Y(n9078) );
  OAI221XL U1365 ( .A0(\i_MIPS/Register/register[2][4] ), .A1(net117643), .B0(
        \i_MIPS/Register/register[10][4] ), .B1(net117661), .C0(n9063), .Y(
        n9066) );
  NOR4X2 U1366 ( .A(n8058), .B(n8057), .C(n8056), .D(n8055), .Y(n8069) );
  AO22X1 U1367 ( .A0(net118271), .A1(n561), .B0(net118289), .B1(n2182), .Y(
        n8056) );
  OAI221XL U1368 ( .A0(\i_MIPS/Register/register[2][9] ), .A1(net117639), .B0(
        \i_MIPS/Register/register[10][9] ), .B1(net117657), .C0(n8054), .Y(
        n8057) );
  NOR4X2 U1369 ( .A(n8067), .B(n8066), .C(n8065), .D(n8064), .Y(n8068) );
  AO22X1 U1370 ( .A0(net118271), .A1(n562), .B0(net118289), .B1(n2183), .Y(
        n8065) );
  OAI221XL U1371 ( .A0(\i_MIPS/Register/register[18][9] ), .A1(net117639), 
        .B0(\i_MIPS/Register/register[26][9] ), .B1(net117657), .C0(n8063), 
        .Y(n8066) );
  OAI221XL U1372 ( .A0(\i_MIPS/Register/register[18][12] ), .A1(net117639), 
        .B0(\i_MIPS/Register/register[26][12] ), .B1(net117657), .C0(n8234), 
        .Y(n8237) );
  AO22X2 U1373 ( .A0(net118273), .A1(n424), .B0(net118291), .B1(n2051), .Y(
        n8914) );
  OA22X1 U1374 ( .A0(\i_MIPS/Register/register[22][21] ), .A1(net117681), .B0(
        \i_MIPS/Register/register[30][21] ), .B1(net117697), .Y(n8912) );
  AO22X2 U1375 ( .A0(net118273), .A1(n417), .B0(net118291), .B1(n2044), .Y(
        n8905) );
  NAND3BX1 U1376 ( .AN(net36572), .B(ICACHE_addr[1]), .C(\i_MIPS/PC/n4 ), .Y(
        net107119) );
  NAND3BX1 U1377 ( .AN(net36572), .B(ICACHE_addr[0]), .C(\i_MIPS/PC/n5 ), .Y(
        n9606) );
  NAND2X2 U1378 ( .A(n3023), .B(net105430), .Y(n4361) );
  NAND2X2 U1379 ( .A(net105581), .B(net105582), .Y(n4279) );
  NAND3BX1 U1380 ( .AN(\i_MIPS/IR[30] ), .B(n9816), .C(n9811), .Y(n9603) );
  AND2X2 U1381 ( .A(n9048), .B(n9047), .Y(n3700) );
  OR2X2 U1382 ( .A(n3627), .B(n3752), .Y(n3736) );
  OA22X1 U1383 ( .A0(n5894), .A1(n536), .B0(n5852), .B1(n2965), .Y(n6373) );
  CLKBUFX2 U1384 ( .A(n5841), .Y(n5830) );
  OA22X1 U1385 ( .A0(n5385), .A1(n574), .B0(n5426), .B1(n2192), .Y(n9267) );
  OA22X2 U1386 ( .A0(n5256), .A1(n2095), .B0(n5299), .B1(n469), .Y(n7191) );
  OA22X2 U1387 ( .A0(n5395), .A1(n2141), .B0(n5439), .B1(n516), .Y(n7345) );
  BUFX12 U1388 ( .A(n5444), .Y(n5433) );
  BUFX4 U1389 ( .A(n5404), .Y(n5386) );
  CLKBUFX3 U1390 ( .A(n5265), .Y(n5245) );
  BUFX12 U1391 ( .A(n5264), .Y(n5252) );
  CLKBUFX8 U1392 ( .A(n5307), .Y(n5292) );
  OA22X2 U1393 ( .A0(n5260), .A1(n2888), .B0(n5294), .B1(n1270), .Y(n6392) );
  INVX3 U1394 ( .A(n6469), .Y(n11043) );
  OA22X2 U1395 ( .A0(n5406), .A1(n2069), .B0(n5445), .B1(n444), .Y(n6470) );
  INVX3 U1396 ( .A(n6427), .Y(n11015) );
  INVX4 U1397 ( .A(n6492), .Y(n11024) );
  INVX4 U1398 ( .A(n6442), .Y(n11007) );
  AND3X4 U1399 ( .A(n4617), .B(n4618), .C(n6440), .Y(n3007) );
  INVX3 U1400 ( .A(n6422), .Y(n10996) );
  INVX3 U1401 ( .A(n6438), .Y(n11009) );
  OR2X1 U1402 ( .A(n5170), .B(n2898), .Y(n4634) );
  OA22X2 U1403 ( .A0(n5263), .A1(n2082), .B0(n5307), .B1(n456), .Y(n6436) );
  INVX3 U1404 ( .A(n6485), .Y(n11028) );
  OAI221X1 U1405 ( .A0(n5329), .A1(n2021), .B0(n5354), .B1(n402), .C0(n6484), 
        .Y(n6485) );
  INVX3 U1406 ( .A(n6412), .Y(n10981) );
  INVX3 U1407 ( .A(n6449), .Y(n11034) );
  INVX6 U1408 ( .A(n6405), .Y(n10985) );
  INVX3 U1409 ( .A(n5261), .Y(n3864) );
  INVX3 U1410 ( .A(n6407), .Y(n10984) );
  AOI2BB2X2 U1411 ( .B0(n3863), .B1(\D_cache/cache[6][144] ), .A0N(n5447), 
        .A1N(n2035), .Y(n6406) );
  INVX3 U1412 ( .A(n6511), .Y(n11017) );
  CLKINVX1 U1413 ( .A(n6509), .Y(n11018) );
  INVX3 U1414 ( .A(n6478), .Y(n11032) );
  OAI221X1 U1415 ( .A0(n5172), .A1(n1336), .B0(n5222), .B1(n2989), .C0(n6477), 
        .Y(n6478) );
  AOI2BB2X2 U1416 ( .B0(n3924), .B1(\D_cache/cache[3][146] ), .A0N(n5259), 
        .A1N(n2040), .Y(n6477) );
  INVX3 U1417 ( .A(n6480), .Y(n11031) );
  OAI221X1 U1418 ( .A0(n5187), .A1(n1334), .B0(n5222), .B1(n2987), .C0(n6498), 
        .Y(n6499) );
  INVX3 U1419 ( .A(n6501), .Y(n11002) );
  OAI221X1 U1420 ( .A0(n5329), .A1(n1335), .B0(n5354), .B1(n2988), .C0(n6500), 
        .Y(n6501) );
  CLKINVX3 U1421 ( .A(n6432), .Y(n11012) );
  NAND3X4 U1422 ( .A(n3738), .B(n3739), .C(n6431), .Y(n6432) );
  OR2X2 U1423 ( .A(n5185), .B(n2891), .Y(n3738) );
  INVX3 U1424 ( .A(n6417), .Y(n10999) );
  OA22X2 U1425 ( .A0(n5259), .A1(n2112), .B0(n5306), .B1(n486), .Y(n6394) );
  INVX3 U1426 ( .A(n6397), .Y(n10990) );
  OA22X2 U1427 ( .A0(n5407), .A1(n2109), .B0(n5446), .B1(n483), .Y(n6396) );
  NOR4X1 U1428 ( .A(n6780), .B(n6779), .C(n6778), .D(n6777), .Y(n6791) );
  OR2X4 U1429 ( .A(n8218), .B(n8217), .Y(n3688) );
  CLKMX2X2 U1430 ( .A(n6891), .B(n6890), .S0(n3001), .Y(n6892) );
  NOR4X1 U1431 ( .A(n6889), .B(n6888), .C(n6887), .D(n6886), .Y(n6890) );
  NOR4X1 U1432 ( .A(n6880), .B(n6879), .C(n6878), .D(n6877), .Y(n6891) );
  NOR4X2 U1433 ( .A(n9252), .B(n9251), .C(n9250), .D(n9249), .Y(n9253) );
  NOR4X2 U1434 ( .A(n9243), .B(n9242), .C(n9241), .D(n9240), .Y(n9254) );
  NAND4X1 U1435 ( .A(n9329), .B(n9328), .C(n9327), .D(n9326), .Y(n9334) );
  NOR4X2 U1436 ( .A(n9343), .B(n9342), .C(n9341), .D(n9340), .Y(n9344) );
  CLKINVX1 U1437 ( .A(n3713), .Y(n7230) );
  CLKMX2X2 U1438 ( .A(n8368), .B(n8367), .S0(net114081), .Y(n8369) );
  NAND4BX1 U1439 ( .AN(n8366), .B(n8365), .C(n8364), .D(n8363), .Y(n8367) );
  OAI221XL U1440 ( .A0(\i_MIPS/Register/register[18][19] ), .A1(n5090), .B0(
        \i_MIPS/Register/register[26][19] ), .B1(n4669), .C0(n8358), .Y(n8366)
         );
  NAND2X1 U1441 ( .A(\i_MIPS/ALUin1[30] ), .B(n3977), .Y(n9539) );
  CLKINVX1 U1442 ( .A(n9440), .Y(n3556) );
  AOI2BB1X1 U1443 ( .A0N(n9431), .A1N(n9430), .B0(n9434), .Y(n9440) );
  INVX3 U1444 ( .A(n10167), .Y(n10179) );
  AND2X6 U1445 ( .A(n7608), .B(n7610), .Y(n3832) );
  AO22X2 U1446 ( .A0(n5157), .A1(n426), .B0(n5153), .B1(n2053), .Y(n8440) );
  NOR4X2 U1447 ( .A(n8452), .B(n8451), .C(n8450), .D(n8449), .Y(n8453) );
  AO22X2 U1448 ( .A0(n5156), .A1(n425), .B0(n5153), .B1(n2052), .Y(n8449) );
  AO22XL U1449 ( .A0(n5123), .A1(n356), .B0(n5119), .B1(n2176), .Y(n8452) );
  INVX3 U1450 ( .A(n9729), .Y(n10713) );
  AO21X2 U1451 ( .A0(net105334), .A1(net105335), .B0(net117623), .Y(net105479)
         );
  OAI2BB1X1 U1452 ( .A0N(net105110), .A1N(net105111), .B0(net117631), .Y(
        net105105) );
  AOI32X1 U1453 ( .A0(net117631), .A1(n3970), .A2(n7836), .B0(n7813), .B1(
        net117631), .Y(n7814) );
  INVX3 U1454 ( .A(n4758), .Y(n5104) );
  AO22X1 U1455 ( .A0(n5155), .A1(n422), .B0(n5153), .B1(n2049), .Y(n8845) );
  AO22X1 U1456 ( .A0(n5155), .A1(n423), .B0(n5153), .B1(n2050), .Y(n8836) );
  CLKMX2X2 U1457 ( .A(n7339), .B(n7338), .S0(net114087), .Y(n7340) );
  INVX3 U1458 ( .A(n10256), .Y(n10263) );
  AND2X2 U1459 ( .A(\i_MIPS/IF_ID[13] ), .B(\i_MIPS/Sign_Extend[11] ), .Y(
        n4806) );
  CLKINVX1 U1460 ( .A(\i_MIPS/IR[31] ), .Y(n9816) );
  AND3X2 U1461 ( .A(n8573), .B(n8550), .C(n8287), .Y(n8306) );
  NAND3X4 U1462 ( .A(n3646), .B(n3647), .C(n8284), .Y(n8307) );
  AND4X4 U1463 ( .A(n6959), .B(n6958), .C(n6957), .D(n6956), .Y(n6962) );
  CLKAND2X8 U1464 ( .A(n7437), .B(n7438), .Y(n3028) );
  NOR4X4 U1465 ( .A(n6680), .B(net107841), .C(n6679), .D(n6678), .Y(n6681) );
  CLKMX2X2 U1466 ( .A(net107656), .B(net107657), .S0(n6849), .Y(n6678) );
  AOI32X1 U1467 ( .A0(n6661), .A1(n3673), .A2(n3748), .B0(n6660), .B1(n9445), 
        .Y(n6684) );
  CLKINVX1 U1468 ( .A(n8789), .Y(n6660) );
  NAND2XL U1469 ( .A(n6920), .B(n6918), .Y(n6729) );
  MXI2X6 U1470 ( .A(\i_MIPS/ID_EX[87] ), .B(\i_MIPS/ID_EX[114] ), .S0(n4790), 
        .Y(n6634) );
  OR2X6 U1471 ( .A(n9487), .B(net107141), .Y(n3994) );
  NAND4BX1 U1472 ( .AN(n9475), .B(n9474), .C(n9473), .D(n9472), .Y(n9486) );
  NAND2X1 U1473 ( .A(n6919), .B(n7431), .Y(n6826) );
  INVXL U1474 ( .A(n6918), .Y(n6825) );
  NOR4X4 U1475 ( .A(n6847), .B(n6846), .C(n6845), .D(n6844), .Y(n6851) );
  CLKINVX1 U1476 ( .A(n3612), .Y(n6845) );
  AND2X2 U1477 ( .A(n6849), .B(n6827), .Y(n6847) );
  NAND3BX1 U1478 ( .AN(n8888), .B(n8887), .C(n3950), .Y(n8896) );
  OAI222X1 U1479 ( .A0(net107217), .A1(n8382), .B0(n8372), .B1(n8856), .C0(
        n8371), .C1(net117757), .Y(n8376) );
  OA22X2 U1480 ( .A0(n8388), .A1(n8793), .B0(n8387), .B1(n8874), .Y(n8389) );
  CLKAND2X4 U1481 ( .A(net117747), .B(n8385), .Y(n4693) );
  INVX3 U1482 ( .A(n8397), .Y(n8682) );
  CLKINVX1 U1483 ( .A(n8682), .Y(n3665) );
  CLKINVX1 U1484 ( .A(n8396), .Y(n8395) );
  AND2X2 U1485 ( .A(net117745), .B(n8393), .Y(n4698) );
  INVXL U1486 ( .A(n9216), .Y(n9209) );
  NAND2XL U1487 ( .A(n8687), .B(n8681), .Y(n8567) );
  INVX3 U1488 ( .A(n10323), .Y(n10333) );
  NOR3X1 U1489 ( .A(\i_MIPS/Reg_W[0] ), .B(\i_MIPS/Reg_W[2] ), .C(n4833), .Y(
        \i_MIPS/Register/n115 ) );
  INVX3 U1490 ( .A(n10265), .Y(n10471) );
  INVX3 U1491 ( .A(n10292), .Y(n10301) );
  INVX3 U1492 ( .A(n10341), .Y(n10354) );
  NOR3X1 U1493 ( .A(\i_MIPS/Reg_W[1] ), .B(\i_MIPS/Reg_W[2] ), .C(
        \i_MIPS/Reg_W[0] ), .Y(\i_MIPS/Register/n119 ) );
  NOR3X1 U1494 ( .A(\i_MIPS/Reg_W[1] ), .B(\i_MIPS/Reg_W[2] ), .C(n1988), .Y(
        \i_MIPS/Register/n117 ) );
  NOR3X1 U1495 ( .A(n1988), .B(\i_MIPS/Reg_W[2] ), .C(n4833), .Y(
        \i_MIPS/Register/n113 ) );
  NOR3X1 U1496 ( .A(n1988), .B(\i_MIPS/Reg_W[1] ), .C(n223), .Y(
        \i_MIPS/Register/n109 ) );
  NOR3BX2 U1497 ( .AN(\i_MIPS/Register/n120 ), .B(\i_MIPS/Reg_W[3] ), .C(
        \i_MIPS/Reg_W[4] ), .Y(\i_MIPS/Register/n140 ) );
  NOR3BX2 U1498 ( .AN(\i_MIPS/Register/n120 ), .B(\i_MIPS/Reg_W[3] ), .C(n1932), .Y(\i_MIPS/Register/n122 ) );
  NOR3BX2 U1499 ( .AN(\i_MIPS/Register/n120 ), .B(\i_MIPS/Reg_W[4] ), .C(n1931), .Y(\i_MIPS/Register/n131 ) );
  NOR3X1 U1500 ( .A(n4833), .B(\i_MIPS/Reg_W[0] ), .C(n223), .Y(
        \i_MIPS/Register/n107 ) );
  NAND4X2 U1501 ( .A(n9528), .B(n9527), .C(n9526), .D(n9525), .Y(n11407) );
  OA22X1 U1502 ( .A0(n5177), .A1(n704), .B0(n5218), .B1(n2324), .Y(n9528) );
  OA22X1 U1503 ( .A0(n5374), .A1(n703), .B0(n5420), .B1(n2323), .Y(n9525) );
  OA22XL U1504 ( .A0(n5333), .A1(n581), .B0(n5360), .B1(n2199), .Y(n7806) );
  OA22XL U1505 ( .A0(n5255), .A1(n580), .B0(n5295), .B1(n2198), .Y(n7807) );
  INVX4 U1506 ( .A(n11381), .Y(n10897) );
  CLKINVX1 U1507 ( .A(n11377), .Y(n10667) );
  CLKINVX1 U1508 ( .A(n11435), .Y(n10400) );
  NAND4X1 U1509 ( .A(n7076), .B(n7075), .C(n7074), .D(n7073), .Y(n11431) );
  OA22XL U1510 ( .A0(n5397), .A1(n630), .B0(n5441), .B1(n2247), .Y(n7073) );
  OA22X1 U1511 ( .A0(n5181), .A1(n632), .B0(n5218), .B1(n2249), .Y(n7076) );
  OA22X1 U1512 ( .A0(n5241), .A1(n631), .B0(n5300), .B1(n2248), .Y(n7075) );
  OA22XL U1513 ( .A0(n5174), .A1(n643), .B0(n5213), .B1(n2260), .Y(n8436) );
  OA22XL U1514 ( .A0(n5330), .A1(n624), .B0(n5355), .B1(n2242), .Y(n8434) );
  INVX3 U1515 ( .A(n11426), .Y(n10643) );
  OAI22XL U1516 ( .A0(n5179), .A1(n557), .B0(n5218), .B1(n2178), .Y(n4647) );
  NAND4X2 U1517 ( .A(n8527), .B(n8526), .C(n8525), .D(n8524), .Y(n11419) );
  OA22X1 U1518 ( .A0(n5175), .A1(n701), .B0(n5214), .B1(n2321), .Y(n8527) );
  OA22X1 U1519 ( .A0(n5389), .A1(n700), .B0(n5439), .B1(n2320), .Y(n8524) );
  OAI22XL U1520 ( .A0(n5179), .A1(n558), .B0(n5213), .B1(n2179), .Y(n4646) );
  OA22XL U1521 ( .A0(n5394), .A1(n707), .B0(n5437), .B1(n2327), .Y(n7538) );
  OA22X1 U1522 ( .A0(n5329), .A1(n592), .B0(n5354), .B1(n2210), .Y(n8174) );
  OA22X1 U1523 ( .A0(n5374), .A1(n705), .B0(n5433), .B1(n2325), .Y(n8173) );
  OA22X1 U1524 ( .A0(n5173), .A1(n706), .B0(n5218), .B1(n2326), .Y(n8176) );
  AND2X2 U1525 ( .A(n5541), .B(n11414), .Y(n4392) );
  AND2X2 U1526 ( .A(mem_rdata_D[38]), .B(n129), .Y(n4393) );
  OAI22XL U1527 ( .A0(n5177), .A1(n560), .B0(n5216), .B1(n2181), .Y(n4645) );
  OA22X1 U1528 ( .A0(n5385), .A1(n697), .B0(n5426), .B1(n2315), .Y(n9177) );
  OA22XL U1529 ( .A0(n5176), .A1(n694), .B0(n5215), .B1(n2312), .Y(n9019) );
  OA22X1 U1530 ( .A0(n5387), .A1(n693), .B0(n5428), .B1(n2311), .Y(n9016) );
  OA22X2 U1531 ( .A0(n5246), .A1(n2133), .B0(n5296), .B1(n508), .Y(n9018) );
  OA22X1 U1532 ( .A0(n5175), .A1(n699), .B0(n5214), .B1(n2317), .Y(n8756) );
  OA22X1 U1533 ( .A0(n5388), .A1(n698), .B0(n5430), .B1(n2316), .Y(n8753) );
  BUFX20 U1534 ( .A(n10973), .Y(n5541) );
  OA22X1 U1535 ( .A0(n5180), .A1(n619), .B0(n5218), .B1(n2237), .Y(n7268) );
  NAND4X2 U1536 ( .A(n6968), .B(n6967), .C(n6966), .D(n6965), .Y(n11501) );
  OA22X1 U1537 ( .A0(n5399), .A1(n596), .B0(n5443), .B1(n2214), .Y(n6965) );
  BUFX6 U1538 ( .A(n5336), .Y(n5325) );
  BUFX4 U1539 ( .A(n5187), .Y(n5171) );
  BUFX6 U1540 ( .A(n5261), .Y(n5260) );
  INVX3 U1541 ( .A(n11477), .Y(n10891) );
  BUFX16 U1542 ( .A(n5363), .Y(n5352) );
  BUFX16 U1543 ( .A(n5335), .Y(n5327) );
  BUFX8 U1544 ( .A(n5187), .Y(n5169) );
  OAI21X2 U1545 ( .A0(n3880), .A1(n3881), .B0(n3970), .Y(net105752) );
  OA22X2 U1546 ( .A0(n10744), .A1(n3879), .B0(n10747), .B1(n4495), .Y(n8757)
         );
  INVX12 U1547 ( .A(n5193), .Y(n3969) );
  INVX4 U1548 ( .A(n3970), .Y(n5192) );
  OA22X2 U1549 ( .A0(n10437), .A1(n3877), .B0(n10440), .B1(n4495), .Y(n6870)
         );
  NAND4BX1 U1550 ( .AN(n7475), .B(n7474), .C(n7473), .D(n7472), .Y(n7476) );
  INVX8 U1551 ( .A(n3876), .Y(n3878) );
  CLKINVX1 U1552 ( .A(n11439), .Y(n10708) );
  NOR3X1 U1553 ( .A(\i_MIPS/Reg_W[0] ), .B(\i_MIPS/Reg_W[1] ), .C(n223), .Y(
        \i_MIPS/Register/n111 ) );
  CLKBUFX8 U1554 ( .A(n11085), .Y(n5571) );
  BUFX6 U1555 ( .A(n11085), .Y(n5570) );
  CLKBUFX8 U1556 ( .A(n5565), .Y(n5567) );
  CLKBUFX8 U1557 ( .A(n5565), .Y(n5566) );
  INVX3 U1558 ( .A(n10531), .Y(n10568) );
  OR2X1 U1559 ( .A(n3789), .B(n5542), .Y(n3635) );
  BUFX4 U1560 ( .A(net107977), .Y(n3752) );
  NAND2X4 U1561 ( .A(net134876), .B(net108631), .Y(net107661) );
  OA22X1 U1562 ( .A0(n8863), .A1(n7675), .B0(n7680), .B1(n8699), .Y(net111710)
         );
  CLKINVX1 U1563 ( .A(n8648), .Y(n8476) );
  OAI222X1 U1564 ( .A0(n9316), .A1(n8460), .B0(n8459), .B1(n5049), .C0(
        net107217), .C1(n8464), .Y(n8475) );
  INVX3 U1565 ( .A(n10051), .Y(n10138) );
  NOR4X1 U1566 ( .A(n9001), .B(n9000), .C(n8999), .D(n8998), .Y(n9002) );
  OAI221XL U1567 ( .A0(\i_MIPS/Register/register[2][8] ), .A1(net117639), .B0(
        \i_MIPS/Register/register[10][8] ), .B1(net117657), .C0(n8145), .Y(
        n8148) );
  NAND4X1 U1568 ( .A(n8144), .B(n8143), .C(n8142), .D(n8141), .Y(n8149) );
  INVX3 U1569 ( .A(n9802), .Y(n9935) );
  XOR2XL U1570 ( .A(\i_MIPS/ID_EX[112] ), .B(n248), .Y(
        \i_MIPS/Hazard_detection/n12 ) );
  INVX4 U1571 ( .A(n3859), .Y(n3860) );
  NAND4X1 U1572 ( .A(n6541), .B(n6540), .C(n6539), .D(n6538), .Y(n11254) );
  NAND4X1 U1573 ( .A(n9709), .B(n9708), .C(n9707), .D(n9706), .Y(n11255) );
  NAND4X1 U1574 ( .A(n9872), .B(n9871), .C(n9870), .D(n9869), .Y(n11259) );
  NAND4X1 U1575 ( .A(n9828), .B(n9827), .C(n9826), .D(n9825), .Y(n11260) );
  NAND4X1 U1576 ( .A(n10079), .B(n10078), .C(n10077), .D(n10076), .Y(n11261)
         );
  NAND4X1 U1577 ( .A(n10213), .B(n10212), .C(n10211), .D(n10210), .Y(n11263)
         );
  NAND4X1 U1578 ( .A(n10235), .B(n10234), .C(n10233), .D(n10232), .Y(n11264)
         );
  NAND4X1 U1579 ( .A(n10056), .B(n10055), .C(n10054), .D(n10053), .Y(n11265)
         );
  BUFX8 U1580 ( .A(n11537), .Y(n5951) );
  NAND2X1 U1581 ( .A(n11344), .B(n11346), .Y(n11345) );
  OA22X1 U1582 ( .A0(n5662), .A1(n2154), .B0(n5615), .B1(n529), .Y(n4670) );
  OA22X1 U1583 ( .A0(n5717), .A1(n535), .B0(n5703), .B1(n2964), .Y(n6375) );
  AOI2BB2X1 U1584 ( .B0(n4830), .B1(\I_cache/cache[5][128] ), .A0N(n5808), 
        .A1N(n2924), .Y(n6374) );
  NAND4X4 U1585 ( .A(n11163), .B(n11162), .C(n11161), .D(n11160), .Y(n11348)
         );
  OA22X1 U1586 ( .A0(n5653), .A1(n627), .B0(n5616), .B1(n2245), .Y(n11163) );
  OA22X1 U1587 ( .A0(n5919), .A1(n576), .B0(n5877), .B1(n2194), .Y(n11160) );
  NAND4X2 U1588 ( .A(n11176), .B(n11175), .C(n11174), .D(n11173), .Y(n11354)
         );
  OA22X2 U1589 ( .A0(n5748), .A1(n2117), .B0(n5695), .B1(n491), .Y(n11175) );
  OA22X1 U1590 ( .A0(n5918), .A1(n2969), .B0(n5876), .B1(n493), .Y(n11128) );
  OAI22X1 U1591 ( .A0(n5652), .A1(n376), .B0(n5608), .B1(n2008), .Y(n4644) );
  OA22X2 U1592 ( .A0(n5654), .A1(n3011), .B0(n5608), .B1(n1342), .Y(n4654) );
  OA22X2 U1593 ( .A0(n5654), .A1(n533), .B0(n5608), .B1(n2930), .Y(n4655) );
  NAND4X2 U1594 ( .A(n11186), .B(n11185), .C(n11184), .D(n11183), .Y(n11368)
         );
  NAND4X2 U1595 ( .A(n7196), .B(n7195), .C(n7194), .D(n7193), .Y(n11378) );
  OA22X1 U1596 ( .A0(n5181), .A1(n684), .B0(n5218), .B1(n2302), .Y(n7196) );
  OA22X1 U1597 ( .A0(n5396), .A1(n683), .B0(n5440), .B1(n2301), .Y(n7193) );
  OA22X1 U1598 ( .A0(n5180), .A1(n690), .B0(n5218), .B1(n2308), .Y(n7272) );
  OA22X1 U1599 ( .A0(n5396), .A1(n689), .B0(n5440), .B1(n2307), .Y(n7269) );
  OA22X2 U1600 ( .A0(n5390), .A1(n2071), .B0(n5432), .B1(n446), .Y(n8249) );
  OA22XL U1601 ( .A0(n5247), .A1(n2125), .B0(n5287), .B1(n500), .Y(n8827) );
  OA22XL U1602 ( .A0(n5331), .A1(n607), .B0(n5356), .B1(n2225), .Y(n8826) );
  NAND4X2 U1603 ( .A(n9266), .B(n9265), .C(n9264), .D(n9263), .Y(n11393) );
  OA22X1 U1604 ( .A0(n5385), .A1(n2128), .B0(n5426), .B1(n503), .Y(n9263) );
  OA22X2 U1605 ( .A0(n5394), .A1(n2145), .B0(n5431), .B1(n520), .Y(n8429) );
  NAND4X2 U1606 ( .A(n7914), .B(n7913), .C(n7912), .D(n7911), .Y(n11398) );
  INVX3 U1607 ( .A(n11403), .Y(n10397) );
  INVX3 U1608 ( .A(n11411), .Y(n10765) );
  INVX4 U1609 ( .A(n11413), .Y(n10900) );
  INVX3 U1610 ( .A(n11421), .Y(n10808) );
  OA22X1 U1611 ( .A0(n5177), .A1(n2152), .B0(n5216), .B1(n527), .Y(n9270) );
  OA22XL U1612 ( .A0(n5244), .A1(n2147), .B0(n5285), .B1(n522), .Y(n9269) );
  OA22XL U1613 ( .A0(n5333), .A1(n2149), .B0(n5358), .B1(n524), .Y(n9268) );
  OA22X2 U1614 ( .A0(n5395), .A1(n2144), .B0(n5431), .B1(n519), .Y(n8343) );
  INVX3 U1615 ( .A(n11428), .Y(n10413) );
  NAND4X2 U1616 ( .A(n6869), .B(n6868), .C(n6867), .D(n6866), .Y(n11433) );
  OA22XL U1617 ( .A0(n5335), .A1(n2886), .B0(n5360), .B1(n1268), .Y(n6867) );
  OA22X1 U1618 ( .A0(n5399), .A1(n649), .B0(n5443), .B1(n2266), .Y(n6866) );
  OA22XL U1619 ( .A0(n5334), .A1(n597), .B0(n5361), .B1(n2215), .Y(n7453) );
  OA22X1 U1620 ( .A0(n5180), .A1(n615), .B0(n5218), .B1(n2233), .Y(n7455) );
  OA22XL U1621 ( .A0(n5179), .A1(n662), .B0(n5213), .B1(n2279), .Y(n7716) );
  OA22X2 U1622 ( .A0(n5393), .A1(n2075), .B0(n5436), .B1(n450), .Y(n7713) );
  NAND4X2 U1623 ( .A(n7188), .B(n7187), .C(n7186), .D(n7185), .Y(n11474) );
  NAND4X2 U1624 ( .A(n7991), .B(n7990), .C(n7989), .D(n7988), .Y(n11485) );
  OA22XL U1625 ( .A0(n5178), .A1(n669), .B0(n5217), .B1(n2287), .Y(n7991) );
  OA22XL U1626 ( .A0(n5333), .A1(n583), .B0(n5359), .B1(n2201), .Y(n7989) );
  OA22X1 U1627 ( .A0(n5391), .A1(n668), .B0(n5434), .B1(n2286), .Y(n7988) );
  NAND4X2 U1628 ( .A(n7800), .B(n7799), .C(n7798), .D(n7797), .Y(n11486) );
  OA22XL U1629 ( .A0(n5255), .A1(n579), .B0(n5295), .B1(n2197), .Y(n7799) );
  OA22XL U1630 ( .A0(n5331), .A1(n608), .B0(n5356), .B1(n2226), .Y(n8818) );
  OA22X2 U1631 ( .A0(n5395), .A1(n2127), .B0(n5429), .B1(n502), .Y(n8817) );
  NAND4X2 U1632 ( .A(n8334), .B(n8333), .C(n8332), .D(n8331), .Y(n11491) );
  OA22XL U1633 ( .A0(n5174), .A1(n665), .B0(n5213), .B1(n2283), .Y(n8334) );
  NAND4X2 U1634 ( .A(n7064), .B(n7063), .C(n7062), .D(n7061), .Y(n11495) );
  OA22X1 U1635 ( .A0(n5181), .A1(n686), .B0(n5218), .B1(n2304), .Y(n7064) );
  OA22X1 U1636 ( .A0(n5398), .A1(n685), .B0(n5442), .B1(n2303), .Y(n7061) );
  NAND4X2 U1637 ( .A(n7614), .B(n7613), .C(n7612), .D(n7611), .Y(n11500) );
  OA22XL U1638 ( .A0(n5179), .A1(n692), .B0(n5213), .B1(n2310), .Y(n7614) );
  OA22XL U1639 ( .A0(n5333), .A1(n587), .B0(n5360), .B1(n2205), .Y(n7612) );
  NAND2X1 U1640 ( .A(n11506), .B(n4996), .Y(n11507) );
  CLKINVX1 U1641 ( .A(n6474), .Y(n11040) );
  MXI2X4 U1642 ( .A(\i_MIPS/ID_EX[85] ), .B(\i_MIPS/ID_EX[112] ), .S0(n4790), 
        .Y(n10848) );
  BUFX4 U1643 ( .A(n10409), .Y(n4549) );
  MXI2X1 U1644 ( .A(n10418), .B(n10417), .S0(n5544), .Y(n10419) );
  MXI2X1 U1645 ( .A(n10432), .B(n10431), .S0(n5544), .Y(n10433) );
  CLKMX2X2 U1646 ( .A(net112585), .B(net112586), .S0(net114079), .Y(net112328)
         );
  NAND4BX1 U1647 ( .AN(n6619), .B(n6618), .C(n6617), .D(n6616), .Y(net112585)
         );
  NAND4BX1 U1648 ( .AN(n6628), .B(n6627), .C(n6626), .D(n6625), .Y(net112586)
         );
  NAND2X1 U1649 ( .A(net117715), .B(net110227), .Y(net105435) );
  CLKINVX1 U1650 ( .A(n11226), .Y(n3799) );
  OR2X6 U1651 ( .A(n4450), .B(n4451), .Y(n3661) );
  CLKINVX1 U1652 ( .A(n11288), .Y(n3802) );
  CLKMX2X2 U1653 ( .A(net107857), .B(net107858), .S0(net114079), .Y(net107854)
         );
  CLKINVX1 U1654 ( .A(n10255), .Y(n10479) );
  AND2X2 U1655 ( .A(\i_MIPS/IF_ID[12] ), .B(\i_MIPS/Sign_Extend[10] ), .Y(
        n4797) );
  NAND4X1 U1656 ( .A(n10816), .B(n10815), .C(n10814), .D(n10813), .Y(n11219)
         );
  CLKINVX1 U1657 ( .A(n11307), .Y(n3803) );
  CLKINVX1 U1658 ( .A(n11245), .Y(n3795) );
  CLKINVX1 U1659 ( .A(n11308), .Y(n3804) );
  CLKINVX1 U1660 ( .A(n11246), .Y(n3796) );
  CLKINVX1 U1661 ( .A(n11248), .Y(n3797) );
  NAND2X6 U1662 ( .A(n3623), .B(n4629), .Y(n4630) );
  CLKMX2X2 U1663 ( .A(n7298), .B(n7297), .S0(net114081), .Y(net111276) );
  BUFX4 U1664 ( .A(n10406), .Y(n4557) );
  BUFX4 U1665 ( .A(n10969), .Y(n4536) );
  BUFX4 U1666 ( .A(n10422), .Y(n4548) );
  BUFX4 U1667 ( .A(n10704), .Y(n4562) );
  BUFX4 U1668 ( .A(n10639), .Y(n4567) );
  BUFX4 U1669 ( .A(n10743), .Y(n4541) );
  BUFX4 U1670 ( .A(n10436), .Y(n4547) );
  CLKINVX1 U1671 ( .A(n11228), .Y(n3810) );
  CLKINVX1 U1672 ( .A(n11290), .Y(n3811) );
  NAND4X1 U1673 ( .A(n10943), .B(n10942), .C(n10941), .D(n10940), .Y(n11253)
         );
  CLKINVX1 U1674 ( .A(n11222), .Y(n3807) );
  CLKINVX1 U1675 ( .A(n11223), .Y(n3808) );
  CLKMX2X2 U1676 ( .A(n7023), .B(n7022), .S0(\i_MIPS/jump_addr[22] ), .Y(
        net111762) );
  CLKMX2X4 U1677 ( .A(n9117), .B(n9116), .S0(net114079), .Y(n9120) );
  NAND4X1 U1678 ( .A(n9850), .B(n9849), .C(n9848), .D(n9847), .Y(n11258) );
  INVX3 U1679 ( .A(net105003), .Y(n4345) );
  CLKINVX1 U1680 ( .A(n11238), .Y(n3809) );
  OR2X4 U1681 ( .A(net108160), .B(net117709), .Y(n3990) );
  CLKINVX1 U1682 ( .A(n11234), .Y(n3812) );
  CLKINVX1 U1683 ( .A(n11278), .Y(n3728) );
  CLKINVX1 U1684 ( .A(n11311), .Y(n3801) );
  NAND4X1 U1685 ( .A(n9916), .B(n9915), .C(n9914), .D(n9913), .Y(n11256) );
  OR2X2 U1686 ( .A(net109989), .B(net117711), .Y(n3960) );
  AO21X2 U1687 ( .A0(n10111), .A1(n10110), .B0(net107195), .Y(n7837) );
  OR2X2 U1688 ( .A(n7839), .B(net117711), .Y(n3962) );
  INVX4 U1689 ( .A(net105167), .Y(net108491) );
  OAI2BB1X2 U1690 ( .A0N(net106037), .A1N(net106038), .B0(n3989), .Y(net107519) );
  XOR2X1 U1691 ( .A(\i_MIPS/PC/n4 ), .B(ICACHE_addr[1]), .Y(n9734) );
  INVX3 U1692 ( .A(n3558), .Y(n3559) );
  INVX3 U1693 ( .A(n3883), .Y(n6713) );
  MX2XL U1694 ( .A(net118597), .B(net118592), .S0(n7161), .Y(n7162) );
  AND2X2 U1695 ( .A(n7155), .B(net109965), .Y(n3893) );
  INVX6 U1696 ( .A(n6633), .Y(n10846) );
  CLKAND2X3 U1697 ( .A(n7503), .B(n7502), .Y(n2981) );
  INVX3 U1698 ( .A(net105010), .Y(net109840) );
  AO22X1 U1699 ( .A0(n5554), .A1(DCACHE_addr[28]), .B0(n5551), .B1(n11532), 
        .Y(n11001) );
  AO22X1 U1700 ( .A0(n5554), .A1(DCACHE_addr[28]), .B0(n5551), .B1(n11532), 
        .Y(n3794) );
  AO22X2 U1701 ( .A0(n5554), .A1(DCACHE_addr[25]), .B0(n5551), .B1(n11529), 
        .Y(n11013) );
  AO22X2 U1702 ( .A0(n5554), .A1(n12957), .B0(n5551), .B1(n11530), .Y(n11006)
         );
  AOI222X1 U1703 ( .A0(n3800), .A1(n11406), .B0(mem_rdata_D[30]), .B1(n133), 
        .C0(n12983), .C1(n5538), .Y(n10599) );
  MXI2X2 U1704 ( .A(n10562), .B(n10561), .S0(n5546), .Y(n10563) );
  MXI2X2 U1705 ( .A(n10549), .B(n10548), .S0(n5546), .Y(n10550) );
  AOI222X1 U1706 ( .A0(n3800), .A1(n11401), .B0(mem_rdata_D[25]), .B1(n131), 
        .C0(n12988), .C1(n5537), .Y(n10438) );
  AOI222X1 U1707 ( .A0(n3800), .A1(n11399), .B0(mem_rdata_D[23]), .B1(n132), 
        .C0(n12990), .C1(n5538), .Y(n10693) );
  MXI2X2 U1708 ( .A(n10521), .B(n10520), .S0(n5546), .Y(n10522) );
  AND2X2 U1709 ( .A(n4411), .B(n4412), .Y(n346) );
  NAND2XL U1710 ( .A(n10971), .B(n5549), .Y(n4412) );
  NAND2X1 U1711 ( .A(n10972), .B(n4410), .Y(n4411) );
  AOI222X1 U1712 ( .A0(n3800), .A1(n11394), .B0(mem_rdata_D[18]), .B1(n129), 
        .C0(n12995), .C1(n5538), .Y(n10641) );
  MXI2X2 U1713 ( .A(n10626), .B(n10625), .S0(n5547), .Y(n10627) );
  AOI222X1 U1714 ( .A0(n3800), .A1(n11393), .B0(mem_rdata_D[17]), .B1(n130), 
        .C0(n12996), .C1(n5538), .Y(n10626) );
  CLKBUFX3 U1715 ( .A(n10452), .Y(n4520) );
  AOI222X1 U1716 ( .A0(n3800), .A1(n11391), .B0(mem_rdata_D[15]), .B1(n129), 
        .C0(n12998), .C1(n5537), .Y(n10451) );
  AOI222X1 U1717 ( .A0(n3800), .A1(n11389), .B0(mem_rdata_D[13]), .B1(n133), 
        .C0(n13000), .C1(n5538), .Y(n10806) );
  CLKBUFX3 U1718 ( .A(n10792), .Y(n4497) );
  CLKBUFX3 U1719 ( .A(n10779), .Y(n4498) );
  AOI222X1 U1720 ( .A0(n3800), .A1(n11384), .B0(mem_rdata_D[8]), .B1(n131), 
        .C0(n13005), .C1(n5538), .Y(n10654) );
  AOI222X1 U1721 ( .A0(n3800), .A1(n11383), .B0(mem_rdata_D[7]), .B1(n131), 
        .C0(n13006), .C1(n5538), .Y(n10681) );
  MXI2X2 U1722 ( .A(n10753), .B(n3979), .S0(n5550), .Y(n10754) );
  AOI222X1 U1723 ( .A0(n3800), .A1(n11376), .B0(mem_rdata_D[0]), .B1(n133), 
        .C0(n13013), .C1(n5538), .Y(n10745) );
  MXI2X2 U1724 ( .A(n10709), .B(n10708), .S0(n5549), .Y(n10710) );
  AOI222X1 U1725 ( .A0(n5541), .A1(n11439), .B0(mem_rdata_D[63]), .B1(n129), 
        .C0(n12982), .C1(n5539), .Y(n10709) );
  MXI2X2 U1726 ( .A(n10565), .B(n10564), .S0(n5546), .Y(n10566) );
  AOI222X1 U1727 ( .A0(n5541), .A1(n11436), .B0(mem_rdata_D[60]), .B1(n129), 
        .C0(n12985), .C1(n5539), .Y(n10552) );
  AOI222X1 U1728 ( .A0(n5541), .A1(n11430), .B0(mem_rdata_D[54]), .B1(n130), 
        .C0(n12991), .C1(n5539), .Y(n10317) );
  AOI222X1 U1729 ( .A0(n5541), .A1(n11429), .B0(mem_rdata_D[53]), .B1(n132), 
        .C0(n12992), .C1(n5539), .Y(n10524) );
  BUFX4 U1730 ( .A(n10455), .Y(n4515) );
  AOI222X1 U1731 ( .A0(n5541), .A1(n11417), .B0(mem_rdata_D[41]), .B1(n130), 
        .C0(n13004), .C1(n5539), .Y(n10616) );
  INVX4 U1732 ( .A(n3578), .Y(n10757) );
  CLKMX2X2 U1733 ( .A(n10755), .B(n10756), .S0(n4410), .Y(n3578) );
  INVX4 U1734 ( .A(n3579), .Y(n10197) );
  CLKMX2X2 U1735 ( .A(n10195), .B(n10196), .S0(n4410), .Y(n3579) );
  CLKBUFX3 U1736 ( .A(n10597), .Y(n4563) );
  CLKBUFX3 U1737 ( .A(n10560), .Y(n4564) );
  BUFX4 U1738 ( .A(n10519), .Y(n4566) );
  CLKBUFX3 U1739 ( .A(n10103), .Y(n4560) );
  CLKBUFX3 U1740 ( .A(n10461), .Y(n4552) );
  CLKBUFX3 U1741 ( .A(n10652), .Y(n4570) );
  AND3X2 U1742 ( .A(n4380), .B(n4381), .C(n4382), .Y(n10678) );
  AOI222X1 U1743 ( .A0(n4505), .A1(n11445), .B0(mem_rdata_D[69]), .B1(n131), 
        .C0(n13008), .C1(n4686), .Y(n10895) );
  BUFX4 U1744 ( .A(n10752), .Y(n4540) );
  MXI2X2 U1745 ( .A(n10760), .B(n10759), .S0(n5550), .Y(n10761) );
  NOR3X1 U1746 ( .A(n4386), .B(n4387), .C(n4388), .Y(n10190) );
  AND2X2 U1747 ( .A(n13011), .B(n5535), .Y(n4388) );
  AOI222X1 U1748 ( .A0(n4506), .A1(n11441), .B0(mem_rdata_D[65]), .B1(n131), 
        .C0(n13012), .C1(n5536), .Y(n10665) );
  AOI222X1 U1749 ( .A0(n4535), .A1(n11503), .B0(mem_rdata_D[127]), .B1(n132), 
        .C0(n12982), .C1(n5534), .Y(n10700) );
  AOI222X1 U1750 ( .A0(n4534), .A1(n11499), .B0(mem_rdata_D[123]), .B1(n129), 
        .C0(n12986), .C1(n5533), .Y(n10392) );
  MXI2X2 U1751 ( .A(n10199), .B(n10198), .S0(n5543), .Y(n10200) );
  BUFX4 U1752 ( .A(n10309), .Y(n4559) );
  BUFX4 U1753 ( .A(n10636), .Y(n4574) );
  AOI222X1 U1754 ( .A0(n4535), .A1(n11489), .B0(mem_rdata_D[113]), .B1(n130), 
        .C0(n12996), .C1(n5534), .Y(n10621) );
  BUFX4 U1755 ( .A(n10446), .Y(n4558) );
  BUFX4 U1756 ( .A(n10773), .Y(n4543) );
  MXI2X1 U1757 ( .A(n10772), .B(n10771), .S0(n5550), .Y(n10773) );
  INVX12 U1758 ( .A(n5211), .Y(n5205) );
  BUFX4 U1759 ( .A(n10608), .Y(n4576) );
  BUFX4 U1760 ( .A(n10676), .Y(n4577) );
  INVX3 U1761 ( .A(n5260), .Y(n5236) );
  INVX4 U1762 ( .A(n3820), .Y(n9810) );
  CLKMX2X2 U1763 ( .A(n9804), .B(n9805), .S0(n4410), .Y(n3820) );
  BUFX6 U1764 ( .A(n10758), .Y(n4561) );
  AND2X2 U1765 ( .A(n4534), .B(n11473), .Y(n4383) );
  INVX6 U1766 ( .A(net117741), .Y(net117733) );
  INVX4 U1767 ( .A(net117715), .Y(net117713) );
  AO22X2 U1768 ( .A0(mem_rdata_I[21]), .A1(n5944), .B0(n5571), .B1(n11239), 
        .Y(n9999) );
  AO22X2 U1769 ( .A0(mem_rdata_I[17]), .A1(n5942), .B0(n5570), .B1(n11236), 
        .Y(n9740) );
  AO22X2 U1770 ( .A0(mem_rdata_I[15]), .A1(n5940), .B0(n5571), .B1(n11234), 
        .Y(n10067) );
  AO22X2 U1771 ( .A0(mem_rdata_I[5]), .A1(n5942), .B0(n5570), .B1(n11224), .Y(
        n9720) );
  AO22X2 U1772 ( .A0(mem_rdata_I[94]), .A1(n5943), .B0(n5569), .B1(n11310), 
        .Y(n9671) );
  AO22X2 U1773 ( .A0(mem_rdata_I[88]), .A1(n5939), .B0(n5569), .B1(n11304), 
        .Y(n10833) );
  AO22X2 U1774 ( .A0(mem_rdata_I[87]), .A1(n5933), .B0(n5569), .B1(n11303), 
        .Y(n10016) );
  AO22X2 U1775 ( .A0(mem_rdata_I[78]), .A1(n5943), .B0(n5569), .B1(n11295), 
        .Y(n10241) );
  AO22X2 U1776 ( .A0(mem_rdata_I[77]), .A1(n5932), .B0(n5569), .B1(n11294), 
        .Y(n10219) );
  AO22X2 U1777 ( .A0(mem_rdata_I[76]), .A1(n5943), .B0(n5569), .B1(n11293), 
        .Y(n10121) );
  AO22X2 U1778 ( .A0(mem_rdata_I[68]), .A1(n5939), .B0(n5569), .B1(n11285), 
        .Y(n10855) );
  AO22X2 U1779 ( .A0(mem_rdata_I[99]), .A1(n5941), .B0(n5573), .B1(n11315), 
        .Y(n10959) );
  INVX4 U1780 ( .A(n10075), .Y(n5462) );
  XOR2X1 U1781 ( .A(n10714), .B(\i_MIPS/PC/n32 ), .Y(n4783) );
  INVX1 U1782 ( .A(n3633), .Y(net104801) );
  INVX6 U1783 ( .A(n3592), .Y(n3591) );
  OR2XL U1784 ( .A(n9598), .B(net107138), .Y(n3986) );
  CLKBUFX3 U1785 ( .A(net115797), .Y(net115791) );
  INVX6 U1786 ( .A(n3592), .Y(n3590) );
  INVX3 U1787 ( .A(n3594), .Y(n3595) );
  INVX4 U1788 ( .A(n3602), .Y(n3603) );
  INVX1 U1789 ( .A(net114331), .Y(n3602) );
  INVX16 U1790 ( .A(n3562), .Y(DCACHE_addr[2]) );
  BUFX16 U1791 ( .A(n12954), .Y(DCACHE_addr[29]) );
  INVX12 U1792 ( .A(n1950), .Y(mem_wdata_I[1]) );
  INVX12 U1793 ( .A(n1951), .Y(mem_wdata_I[2]) );
  INVX12 U1794 ( .A(n1952), .Y(mem_wdata_I[3]) );
  INVX12 U1795 ( .A(n1953), .Y(mem_wdata_I[4]) );
  INVX12 U1796 ( .A(n1954), .Y(mem_wdata_I[5]) );
  INVX12 U1797 ( .A(n1955), .Y(mem_wdata_I[6]) );
  INVX12 U1798 ( .A(n1956), .Y(mem_wdata_I[7]) );
  INVX12 U1799 ( .A(n1957), .Y(mem_wdata_I[8]) );
  INVX12 U1800 ( .A(n1958), .Y(mem_wdata_I[9]) );
  INVX12 U1801 ( .A(n1959), .Y(mem_wdata_I[10]) );
  INVX12 U1802 ( .A(n1960), .Y(mem_wdata_I[11]) );
  INVX12 U1803 ( .A(n1961), .Y(mem_wdata_I[12]) );
  INVX12 U1804 ( .A(n1962), .Y(mem_wdata_I[13]) );
  INVX12 U1805 ( .A(n1963), .Y(mem_wdata_I[14]) );
  INVX12 U1806 ( .A(n1964), .Y(mem_wdata_I[15]) );
  INVX12 U1807 ( .A(n1965), .Y(mem_wdata_I[16]) );
  INVX12 U1808 ( .A(n1966), .Y(mem_wdata_I[17]) );
  INVX12 U1809 ( .A(n1967), .Y(mem_wdata_I[18]) );
  INVX12 U1810 ( .A(n1968), .Y(mem_wdata_I[19]) );
  INVX12 U1811 ( .A(n1969), .Y(mem_wdata_I[20]) );
  INVX12 U1812 ( .A(n1970), .Y(mem_wdata_I[21]) );
  INVX12 U1813 ( .A(n1971), .Y(mem_wdata_I[22]) );
  INVX12 U1814 ( .A(n1972), .Y(mem_wdata_I[23]) );
  INVX12 U1815 ( .A(n1973), .Y(mem_wdata_I[24]) );
  INVX12 U1816 ( .A(n1974), .Y(mem_wdata_I[25]) );
  INVX12 U1817 ( .A(n1975), .Y(mem_wdata_I[26]) );
  INVX12 U1818 ( .A(n1976), .Y(mem_wdata_I[27]) );
  INVX12 U1819 ( .A(n1977), .Y(mem_wdata_I[28]) );
  INVX12 U1820 ( .A(n1978), .Y(mem_wdata_I[29]) );
  INVX12 U1821 ( .A(n1979), .Y(mem_wdata_I[30]) );
  INVX12 U1822 ( .A(n1980), .Y(mem_wdata_I[31]) );
  INVX12 U1823 ( .A(n1981), .Y(mem_wdata_I[32]) );
  INVX12 U1824 ( .A(n1982), .Y(mem_wdata_I[33]) );
  INVX12 U1825 ( .A(n1983), .Y(mem_wdata_I[34]) );
  INVX12 U1826 ( .A(n4064), .Y(mem_wdata_I[35]) );
  NAND2BXL U1827 ( .AN(n5045), .B(n11253), .Y(n4064) );
  INVX12 U1828 ( .A(n4065), .Y(mem_wdata_I[36]) );
  OR2XL U1829 ( .A(n5045), .B(n4066), .Y(n4065) );
  CLKINVX1 U1830 ( .A(n11254), .Y(n4066) );
  INVX12 U1831 ( .A(n4067), .Y(mem_wdata_I[37]) );
  OR2XL U1832 ( .A(n5045), .B(n4068), .Y(n4067) );
  CLKINVX1 U1833 ( .A(n11255), .Y(n4068) );
  INVX12 U1834 ( .A(n4069), .Y(mem_wdata_I[38]) );
  OR2XL U1835 ( .A(n5045), .B(n4070), .Y(n4069) );
  CLKINVX1 U1836 ( .A(n11256), .Y(n4070) );
  INVX12 U1837 ( .A(n4072), .Y(mem_wdata_I[39]) );
  OR2XL U1838 ( .A(n5045), .B(n4073), .Y(n4072) );
  CLKINVX1 U1839 ( .A(n11257), .Y(n4073) );
  INVX12 U1840 ( .A(n4074), .Y(mem_wdata_I[40]) );
  OR2XL U1841 ( .A(n5045), .B(n4075), .Y(n4074) );
  CLKINVX1 U1842 ( .A(n11258), .Y(n4075) );
  INVX12 U1843 ( .A(n4076), .Y(mem_wdata_I[41]) );
  OR2XL U1844 ( .A(n5045), .B(n4077), .Y(n4076) );
  CLKINVX1 U1845 ( .A(n11259), .Y(n4077) );
  INVX12 U1846 ( .A(n4079), .Y(mem_wdata_I[42]) );
  OR2XL U1847 ( .A(n5045), .B(n4080), .Y(n4079) );
  CLKINVX1 U1848 ( .A(n11260), .Y(n4080) );
  INVX12 U1849 ( .A(n4082), .Y(mem_wdata_I[43]) );
  CLKINVX1 U1850 ( .A(n11261), .Y(n4083) );
  INVX12 U1851 ( .A(n4084), .Y(mem_wdata_I[44]) );
  OR2XL U1852 ( .A(n5045), .B(n4085), .Y(n4084) );
  CLKINVX1 U1853 ( .A(n11262), .Y(n4085) );
  INVX12 U1854 ( .A(n4086), .Y(mem_wdata_I[45]) );
  CLKINVX1 U1855 ( .A(n11263), .Y(n4087) );
  INVX12 U1856 ( .A(n4088), .Y(mem_wdata_I[46]) );
  CLKINVX1 U1857 ( .A(n11264), .Y(n4089) );
  CLKINVX12 U1858 ( .A(n4139), .Y(mem_wdata_I[49]) );
  INVX3 U1859 ( .A(n12953), .Y(n4139) );
  CLKINVX12 U1860 ( .A(n4145), .Y(mem_wdata_I[52]) );
  INVX3 U1861 ( .A(n12951), .Y(n4145) );
  CLKINVX12 U1862 ( .A(n4103), .Y(mem_wdata_I[53]) );
  INVX3 U1863 ( .A(n12950), .Y(n4103) );
  INVX16 U1864 ( .A(n4141), .Y(mem_wdata_I[54]) );
  INVX3 U1865 ( .A(n12949), .Y(n4141) );
  CLKINVX12 U1866 ( .A(n4151), .Y(mem_wdata_I[55]) );
  INVX3 U1867 ( .A(n12948), .Y(n4151) );
  CLKINVX12 U1868 ( .A(n4117), .Y(mem_wdata_I[56]) );
  INVX3 U1869 ( .A(n12947), .Y(n4117) );
  INVX16 U1870 ( .A(n4147), .Y(mem_wdata_I[57]) );
  INVX3 U1871 ( .A(n12946), .Y(n4147) );
  CLKINVX12 U1872 ( .A(n4157), .Y(mem_wdata_I[58]) );
  INVX3 U1873 ( .A(n12945), .Y(n4157) );
  CLKINVX12 U1874 ( .A(n4121), .Y(mem_wdata_I[59]) );
  INVX3 U1875 ( .A(n12944), .Y(n4121) );
  INVX16 U1876 ( .A(n4153), .Y(mem_wdata_I[60]) );
  INVX3 U1877 ( .A(n12943), .Y(n4153) );
  CLKINVX12 U1878 ( .A(n4163), .Y(mem_wdata_I[61]) );
  INVX3 U1879 ( .A(n12942), .Y(n4163) );
  CLKINVX12 U1880 ( .A(n4127), .Y(mem_wdata_I[62]) );
  INVX3 U1881 ( .A(n12941), .Y(n4127) );
  INVX16 U1882 ( .A(n4159), .Y(mem_wdata_I[63]) );
  INVX3 U1883 ( .A(n12940), .Y(n4159) );
  CLKINVX12 U1884 ( .A(n4169), .Y(mem_wdata_I[64]) );
  INVX3 U1885 ( .A(n12939), .Y(n4169) );
  CLKINVX12 U1886 ( .A(n4131), .Y(mem_wdata_I[65]) );
  INVX3 U1887 ( .A(n12938), .Y(n4131) );
  INVX16 U1888 ( .A(n4165), .Y(mem_wdata_I[66]) );
  INVX3 U1889 ( .A(n12937), .Y(n4165) );
  CLKINVX12 U1890 ( .A(n4175), .Y(mem_wdata_I[67]) );
  INVX3 U1891 ( .A(n12936), .Y(n4175) );
  CLKINVX12 U1892 ( .A(n4137), .Y(mem_wdata_I[68]) );
  INVX3 U1893 ( .A(n12935), .Y(n4137) );
  INVX16 U1894 ( .A(n4171), .Y(mem_wdata_I[69]) );
  INVX3 U1895 ( .A(n12934), .Y(n4171) );
  CLKINVX12 U1896 ( .A(n4181), .Y(mem_wdata_I[70]) );
  INVX3 U1897 ( .A(n12933), .Y(n4181) );
  CLKINVX12 U1898 ( .A(n4143), .Y(mem_wdata_I[71]) );
  INVX3 U1899 ( .A(n12932), .Y(n4143) );
  INVX16 U1900 ( .A(n4177), .Y(mem_wdata_I[72]) );
  INVX3 U1901 ( .A(n12931), .Y(n4177) );
  CLKINVX12 U1902 ( .A(n4187), .Y(mem_wdata_I[73]) );
  INVX3 U1903 ( .A(n12930), .Y(n4187) );
  CLKINVX12 U1904 ( .A(n4149), .Y(mem_wdata_I[74]) );
  INVX3 U1905 ( .A(n12929), .Y(n4149) );
  INVX16 U1906 ( .A(n4183), .Y(mem_wdata_I[75]) );
  INVX3 U1907 ( .A(n12928), .Y(n4183) );
  CLKINVX12 U1908 ( .A(n4193), .Y(mem_wdata_I[76]) );
  INVX3 U1909 ( .A(n12927), .Y(n4193) );
  CLKINVX12 U1910 ( .A(n4155), .Y(mem_wdata_I[77]) );
  INVX3 U1911 ( .A(n12926), .Y(n4155) );
  INVX16 U1912 ( .A(n4189), .Y(mem_wdata_I[78]) );
  INVX3 U1913 ( .A(n12925), .Y(n4189) );
  CLKINVX12 U1914 ( .A(n4199), .Y(mem_wdata_I[79]) );
  INVX3 U1915 ( .A(n12924), .Y(n4199) );
  CLKINVX12 U1916 ( .A(n4161), .Y(mem_wdata_I[80]) );
  INVX3 U1917 ( .A(n12923), .Y(n4161) );
  INVX16 U1918 ( .A(n4195), .Y(mem_wdata_I[81]) );
  INVX3 U1919 ( .A(n12922), .Y(n4195) );
  CLKINVX12 U1920 ( .A(n4205), .Y(mem_wdata_I[82]) );
  INVX3 U1921 ( .A(n12921), .Y(n4205) );
  CLKINVX12 U1922 ( .A(n4167), .Y(mem_wdata_I[83]) );
  INVX3 U1923 ( .A(n12920), .Y(n4167) );
  INVX16 U1924 ( .A(n4201), .Y(mem_wdata_I[84]) );
  INVX3 U1925 ( .A(n12919), .Y(n4201) );
  CLKINVX12 U1926 ( .A(n4211), .Y(mem_wdata_I[85]) );
  INVX3 U1927 ( .A(n12918), .Y(n4211) );
  CLKINVX12 U1928 ( .A(n4173), .Y(mem_wdata_I[86]) );
  INVX3 U1929 ( .A(n12917), .Y(n4173) );
  INVX16 U1930 ( .A(n4207), .Y(mem_wdata_I[87]) );
  INVX3 U1931 ( .A(n12916), .Y(n4207) );
  CLKINVX12 U1932 ( .A(n4217), .Y(mem_wdata_I[88]) );
  INVX3 U1933 ( .A(n12915), .Y(n4217) );
  CLKINVX12 U1934 ( .A(n4179), .Y(mem_wdata_I[89]) );
  INVX3 U1935 ( .A(n12914), .Y(n4179) );
  INVX16 U1936 ( .A(n4213), .Y(mem_wdata_I[90]) );
  INVX3 U1937 ( .A(n12913), .Y(n4213) );
  CLKINVX12 U1938 ( .A(n4223), .Y(mem_wdata_I[91]) );
  INVX3 U1939 ( .A(n12912), .Y(n4223) );
  CLKINVX12 U1940 ( .A(n4185), .Y(mem_wdata_I[92]) );
  INVX3 U1941 ( .A(n12911), .Y(n4185) );
  INVX16 U1942 ( .A(n4219), .Y(mem_wdata_I[93]) );
  INVX3 U1943 ( .A(n12910), .Y(n4219) );
  CLKINVX12 U1944 ( .A(n4229), .Y(mem_wdata_I[94]) );
  INVX3 U1945 ( .A(n12909), .Y(n4229) );
  CLKINVX12 U1946 ( .A(n4191), .Y(mem_wdata_I[95]) );
  INVX3 U1947 ( .A(n12908), .Y(n4191) );
  INVX16 U1948 ( .A(n4225), .Y(mem_wdata_I[96]) );
  INVX3 U1949 ( .A(n12907), .Y(n4225) );
  CLKINVX12 U1950 ( .A(n4235), .Y(mem_wdata_I[97]) );
  INVX3 U1951 ( .A(n12906), .Y(n4235) );
  CLKINVX12 U1952 ( .A(n4197), .Y(mem_wdata_I[98]) );
  INVX3 U1953 ( .A(n12905), .Y(n4197) );
  INVX16 U1954 ( .A(n4231), .Y(mem_wdata_I[99]) );
  INVX3 U1955 ( .A(n12904), .Y(n4231) );
  CLKINVX12 U1956 ( .A(n4241), .Y(mem_wdata_I[100]) );
  INVX3 U1957 ( .A(n12903), .Y(n4241) );
  CLKINVX12 U1958 ( .A(n4203), .Y(mem_wdata_I[101]) );
  INVX3 U1959 ( .A(n12902), .Y(n4203) );
  INVX16 U1960 ( .A(n4237), .Y(mem_wdata_I[102]) );
  INVX3 U1961 ( .A(n12901), .Y(n4237) );
  CLKINVX12 U1962 ( .A(n4247), .Y(mem_wdata_I[103]) );
  INVX3 U1963 ( .A(n12900), .Y(n4247) );
  CLKINVX12 U1964 ( .A(n4209), .Y(mem_wdata_I[104]) );
  INVX3 U1965 ( .A(n12899), .Y(n4209) );
  INVX16 U1966 ( .A(n4243), .Y(mem_wdata_I[105]) );
  INVX3 U1967 ( .A(n12898), .Y(n4243) );
  CLKINVX12 U1968 ( .A(n4251), .Y(mem_wdata_I[106]) );
  INVX3 U1969 ( .A(n12897), .Y(n4251) );
  CLKINVX12 U1970 ( .A(n4215), .Y(mem_wdata_I[107]) );
  INVX3 U1971 ( .A(n12896), .Y(n4215) );
  INVX16 U1972 ( .A(n4249), .Y(mem_wdata_I[108]) );
  INVX3 U1973 ( .A(n12895), .Y(n4249) );
  CLKINVX12 U1974 ( .A(n4255), .Y(mem_wdata_I[109]) );
  INVX3 U1975 ( .A(n12894), .Y(n4255) );
  CLKINVX12 U1976 ( .A(n4221), .Y(mem_wdata_I[110]) );
  INVX3 U1977 ( .A(n12893), .Y(n4221) );
  INVX16 U1978 ( .A(n4253), .Y(mem_wdata_I[111]) );
  INVX3 U1979 ( .A(n12892), .Y(n4253) );
  CLKINVX12 U1980 ( .A(n4259), .Y(mem_wdata_I[112]) );
  INVX3 U1981 ( .A(n12891), .Y(n4259) );
  CLKINVX12 U1982 ( .A(n4227), .Y(mem_wdata_I[113]) );
  INVX3 U1983 ( .A(n12890), .Y(n4227) );
  INVX16 U1984 ( .A(n4257), .Y(mem_wdata_I[114]) );
  INVX3 U1985 ( .A(n12889), .Y(n4257) );
  CLKINVX12 U1986 ( .A(n4263), .Y(mem_wdata_I[115]) );
  INVX3 U1987 ( .A(n12888), .Y(n4263) );
  CLKINVX12 U1988 ( .A(n4233), .Y(mem_wdata_I[116]) );
  INVX3 U1989 ( .A(n12887), .Y(n4233) );
  INVX16 U1990 ( .A(n4261), .Y(mem_wdata_I[117]) );
  INVX3 U1991 ( .A(n12886), .Y(n4261) );
  CLKINVX12 U1992 ( .A(n4267), .Y(mem_wdata_I[118]) );
  INVX3 U1993 ( .A(n12885), .Y(n4267) );
  CLKINVX12 U1994 ( .A(n4239), .Y(mem_wdata_I[119]) );
  INVX3 U1995 ( .A(n12884), .Y(n4239) );
  INVX16 U1996 ( .A(n4265), .Y(mem_wdata_I[120]) );
  INVX3 U1997 ( .A(n12883), .Y(n4265) );
  CLKINVX12 U1998 ( .A(n4269), .Y(mem_wdata_I[121]) );
  INVX3 U1999 ( .A(n12882), .Y(n4269) );
  CLKINVX12 U2000 ( .A(n4245), .Y(mem_wdata_I[122]) );
  INVX3 U2001 ( .A(n12881), .Y(n4245) );
  CLKINVX12 U2002 ( .A(n4271), .Y(mem_wdata_I[124]) );
  INVX3 U2003 ( .A(n12880), .Y(n4271) );
  INVX12 U2004 ( .A(n4105), .Y(mem_addr_I[8]) );
  AOI2BB2X2 U2005 ( .B0(n5047), .B1(n11348), .A0N(\i_MIPS/PC/n10 ), .A1N(n4106), .Y(n4105) );
  CLKINVX1 U2006 ( .A(mem_read_I), .Y(n4106) );
  INVX3 U2007 ( .A(n12877), .Y(n4107) );
  INVX3 U2008 ( .A(n12876), .Y(n4109) );
  INVX3 U2009 ( .A(n12874), .Y(n4113) );
  INVX3 U2010 ( .A(n12873), .Y(n4115) );
  INVX3 U2011 ( .A(n12871), .Y(n4123) );
  INVX3 U2012 ( .A(n12870), .Y(n4125) );
  INVX12 U2013 ( .A(n4579), .Y(mem_addr_I[17]) );
  INVX3 U2014 ( .A(n12869), .Y(n4579) );
  AO22X2 U2015 ( .A0(ICACHE_addr[15]), .A1(mem_read_I), .B0(n5047), .B1(n11357), .Y(n12869) );
  INVX16 U2016 ( .A(n4129), .Y(mem_addr_I[18]) );
  INVX3 U2017 ( .A(n12868), .Y(n4129) );
  INVX16 U2018 ( .A(n4133), .Y(mem_addr_I[19]) );
  INVX3 U2019 ( .A(n12867), .Y(n4133) );
  INVX16 U2020 ( .A(n4840), .Y(mem_addr_I[22]) );
  INVX3 U2021 ( .A(n12864), .Y(n4840) );
  INVX16 U2022 ( .A(n4844), .Y(mem_addr_I[24]) );
  INVX3 U2023 ( .A(n12862), .Y(n4844) );
  INVX16 U2024 ( .A(n4846), .Y(mem_addr_I[25]) );
  INVX3 U2025 ( .A(n12861), .Y(n4846) );
  INVX16 U2026 ( .A(n4848), .Y(mem_addr_I[26]) );
  INVX3 U2027 ( .A(n12860), .Y(n4848) );
  INVX16 U2028 ( .A(n4850), .Y(mem_addr_I[27]) );
  INVX3 U2029 ( .A(n12859), .Y(n4850) );
  INVX16 U2030 ( .A(n4854), .Y(mem_addr_I[29]) );
  INVX3 U2031 ( .A(n12857), .Y(n4854) );
  INVX16 U2032 ( .A(n4856), .Y(mem_addr_I[30]) );
  INVX3 U2033 ( .A(n12856), .Y(n4856) );
  INVX16 U2034 ( .A(n4858), .Y(mem_addr_I[31]) );
  INVX3 U2035 ( .A(n12855), .Y(n4858) );
  INVX3 U2036 ( .A(n11346), .Y(n11536) );
  OR2X1 U2037 ( .A(n5040), .B(n9960), .Y(n4994) );
  BUFX12 U2038 ( .A(n12854), .Y(mem_wdata_D[48]) );
  INVX12 U2039 ( .A(n1984), .Y(mem_wdata_D[50]) );
  INVX12 U2040 ( .A(n3945), .Y(mem_wdata_D[52]) );
  INVX12 U2041 ( .A(n3946), .Y(mem_wdata_D[55]) );
  INVX12 U2042 ( .A(n4932), .Y(mem_wdata_D[102]) );
  INVX16 U2043 ( .A(n3900), .Y(mem_wdata_D[123]) );
  CLKINVX1 U2044 ( .A(n1930), .Y(n3900) );
  INVX12 U2045 ( .A(n358), .Y(mem_addr_D[7]) );
  AOI22X1 U2046 ( .A0(DCACHE_addr[5]), .A1(n11534), .B0(n5042), .B1(n11509), 
        .Y(n358) );
  AND2X2 U2047 ( .A(n5043), .B(n11510), .Y(n4405) );
  AND2X2 U2048 ( .A(DCACHE_addr[6]), .B(n11534), .Y(n4404) );
  INVX12 U2049 ( .A(n1942), .Y(mem_addr_D[10]) );
  AOI22X1 U2050 ( .A0(DCACHE_addr[8]), .A1(n11534), .B0(n5042), .B1(n11512), 
        .Y(n1942) );
  INVX12 U2051 ( .A(n1943), .Y(mem_addr_D[11]) );
  AOI22X1 U2052 ( .A0(n12974), .A1(n11534), .B0(n5043), .B1(n11513), .Y(n1943)
         );
  INVX12 U2053 ( .A(n1944), .Y(mem_addr_D[12]) );
  AOI22X1 U2054 ( .A0(n12973), .A1(n11534), .B0(n5044), .B1(n11514), .Y(n1944)
         );
  INVX12 U2055 ( .A(n1945), .Y(mem_addr_D[13]) );
  AOI22X1 U2056 ( .A0(DCACHE_addr[11]), .A1(n11534), .B0(n5042), .B1(n11515), 
        .Y(n1945) );
  INVX12 U2057 ( .A(n1946), .Y(mem_addr_D[14]) );
  AOI22X1 U2058 ( .A0(n12971), .A1(n11534), .B0(n5043), .B1(n11516), .Y(n1946)
         );
  INVX12 U2059 ( .A(n1947), .Y(mem_addr_D[15]) );
  AOI22X1 U2060 ( .A0(n12970), .A1(n11534), .B0(n5044), .B1(n11517), .Y(n1947)
         );
  INVX12 U2061 ( .A(n1948), .Y(mem_addr_D[16]) );
  AOI22X1 U2062 ( .A0(n12969), .A1(n11534), .B0(n5042), .B1(n11518), .Y(n1948)
         );
  INVX12 U2063 ( .A(n1949), .Y(mem_addr_D[17]) );
  AOI22X1 U2064 ( .A0(DCACHE_addr[15]), .A1(n11534), .B0(n5043), .B1(n11519), 
        .Y(n1949) );
  INVX12 U2065 ( .A(n4929), .Y(mem_addr_D[18]) );
  CLKINVX1 U2066 ( .A(n12848), .Y(n4929) );
  INVX12 U2067 ( .A(n4941), .Y(mem_addr_D[20]) );
  CLKINVX1 U2068 ( .A(n12847), .Y(n4941) );
  CLKINVX12 U2069 ( .A(n5023), .Y(mem_addr_D[22]) );
  INVX3 U2070 ( .A(n5010), .Y(n5023) );
  AOI2BB1X1 U2071 ( .A0N(\i_MIPS/PC/n22 ), .A1N(net115799), .B0(n10325), .Y(
        n10326) );
  AOI2BB1X1 U2072 ( .A0N(\i_MIPS/PC/n25 ), .A1N(net115799), .B0(n10356), .Y(
        n10357) );
  AOI2BB1X1 U2073 ( .A0N(\i_MIPS/PC/n20 ), .A1N(net115799), .B0(n10295), .Y(
        n10296) );
  AOI2BB1X1 U2074 ( .A0N(\i_MIPS/PC/n11 ), .A1N(net115789), .B0(n10159), .Y(
        n10160) );
  AOI2BB1X1 U2075 ( .A0N(\i_MIPS/PC/n23 ), .A1N(net115789), .B0(n10335), .Y(
        n10336) );
  OAI221X1 U2076 ( .A0(n10388), .A1(n5560), .B0(n5558), .B1(n10389), .C0(
        n10387), .Y(\i_MIPS/PC/n61 ) );
  AOI2BB1X1 U2077 ( .A0N(\i_MIPS/PC/n29 ), .A1N(net115789), .B0(n10386), .Y(
        n10387) );
  OR2X1 U2078 ( .A(\i_MIPS/n510 ), .B(net115793), .Y(n3655) );
  OR2X2 U2079 ( .A(n10097), .B(net143858), .Y(n3654) );
  NAND2X1 U2080 ( .A(net104171), .B(n11231), .Y(n3662) );
  AND2X2 U2081 ( .A(n3663), .B(n11251), .Y(n4426) );
  AOI2BB1X1 U2082 ( .A0N(\i_MIPS/PC/n4 ), .A1N(net115789), .B0(n10826), .Y(
        n10827) );
  INVXL U2083 ( .A(net105137), .Y(net108323) );
  OR2XL U2084 ( .A(n5558), .B(n10496), .Y(n4414) );
  OR2X1 U2085 ( .A(n10368), .B(n4641), .Y(n4415) );
  OR2X1 U2086 ( .A(n10381), .B(n4641), .Y(n4417) );
  OR2XL U2087 ( .A(n5558), .B(n10536), .Y(n4420) );
  OR2X1 U2088 ( .A(n10345), .B(n5561), .Y(n4421) );
  CLKMX2X2 U2089 ( .A(\D_cache/cache[6][149] ), .B(n11006), .S0(n5372), .Y(
        \D_cache/n598 ) );
  CLKMX2X2 U2090 ( .A(\I_cache/cache[6][144] ), .B(n11145), .S0(n5890), .Y(
        n11687) );
  CLKMX2X2 U2091 ( .A(\I_cache/cache[6][113] ), .B(n9740), .S0(n5885), .Y(
        n11935) );
  MX2X1 U2092 ( .A(\I_cache/cache[3][65] ), .B(n10873), .S0(n5671), .Y(n12322)
         );
  CLKMX2X2 U2093 ( .A(\D_cache/cache[7][115] ), .B(n346), .S0(n5418), .Y(
        \D_cache/n869 ) );
  CLKMX2X2 U2094 ( .A(\D_cache/cache[6][115] ), .B(n346), .S0(n3574), .Y(
        \D_cache/n870 ) );
  CLKMX2X2 U2095 ( .A(\D_cache/cache[5][115] ), .B(n346), .S0(n5349), .Y(
        \D_cache/n871 ) );
  CLKMX2X2 U2096 ( .A(\D_cache/cache[4][115] ), .B(n346), .S0(n3763), .Y(
        \D_cache/n872 ) );
  CLKMX2X2 U2097 ( .A(\D_cache/cache[3][115] ), .B(n346), .S0(n5275), .Y(
        \D_cache/n873 ) );
  CLKMX2X2 U2098 ( .A(\D_cache/cache[2][115] ), .B(n346), .S0(n5235), .Y(
        \D_cache/n874 ) );
  CLKMX2X2 U2099 ( .A(\D_cache/cache[1][115] ), .B(n346), .S0(n5207), .Y(
        \D_cache/n875 ) );
  CLKMX2X2 U2100 ( .A(\D_cache/cache[0][115] ), .B(n346), .S0(n5167), .Y(
        \D_cache/n876 ) );
  CLKMX2X2 U2101 ( .A(\D_cache/cache[7][36] ), .B(n4540), .S0(n5418), .Y(
        \D_cache/n1501 ) );
  CLKMX2X2 U2102 ( .A(\D_cache/cache[0][27] ), .B(n10393), .S0(n3565), .Y(
        \D_cache/n1580 ) );
  CLKMX2X2 U2103 ( .A(\D_cache/cache[0][4] ), .B(n9810), .S0(n3564), .Y(
        \D_cache/n1764 ) );
  CLKMX2X2 U2104 ( .A(\D_cache/cache[0][2] ), .B(n10188), .S0(n5167), .Y(
        \D_cache/n1780 ) );
  CLKMX2X2 U2105 ( .A(\I_cache/cache[1][113] ), .B(n9740), .S0(n5574), .Y(
        n11940) );
  OAI221X1 U2106 ( .A0(n5562), .A1(\i_MIPS/n153 ), .B0(n5558), .B1(
        \i_MIPS/PC/n2 ), .C0(n10737), .Y(\i_MIPS/PC/n34 ) );
  OAI221X1 U2107 ( .A0(n10872), .A1(n5561), .B0(n5557), .B1(n10871), .C0(
        n10870), .Y(\i_MIPS/PC/n40 ) );
  AOI2BB1X1 U2108 ( .A0N(\i_MIPS/PC/n8 ), .A1N(net115789), .B0(n10869), .Y(
        n10870) );
  AOI2BB1X1 U2109 ( .A0N(\i_MIPS/PC/n7 ), .A1N(net115789), .B0(n10911), .Y(
        n10912) );
  OAI221X1 U2110 ( .A0(n10937), .A1(n5560), .B0(n5558), .B1(n10936), .C0(
        n10935), .Y(\i_MIPS/PC/n38 ) );
  AOI2BB1XL U2111 ( .A0N(\i_MIPS/PC/n6 ), .A1N(net115789), .B0(n10934), .Y(
        n10935) );
  XNOR2X4 U2112 ( .A(n140), .B(n141), .Y(net107134) );
  NAND3X8 U2113 ( .A(n3992), .B(n3993), .C(n3994), .Y(n141) );
  OAI211X4 U2114 ( .A0(n8303), .A1(n8556), .B0(n8302), .C0(n8301), .Y(n8304)
         );
  AND2X2 U2115 ( .A(n8664), .B(n8663), .Y(n8665) );
  OAI31X2 U2116 ( .A0(n8668), .A1(n3671), .A2(n4750), .B0(n8663), .Y(n8026) );
  NAND2X4 U2117 ( .A(\i_MIPS/ALUin1[8] ), .B(n6704), .Y(n8663) );
  NAND2X2 U2118 ( .A(n7026), .B(n8890), .Y(n7863) );
  BUFX8 U2119 ( .A(n4678), .Y(n5751) );
  CLKINVX4 U2120 ( .A(net104700), .Y(net109990) );
  AOI2BB1X1 U2121 ( .A0N(n8793), .A1N(n8792), .B0(n8791), .Y(n8795) );
  AO21XL U2122 ( .A0(net107977), .A1(n5049), .B0(n8792), .Y(n8712) );
  NAND2X2 U2123 ( .A(net107652), .B(net114073), .Y(n8112) );
  NAND2X2 U2124 ( .A(net134069), .B(net114073), .Y(net107228) );
  AND2X2 U2125 ( .A(n3898), .B(n11289), .Y(n4442) );
  AND2X8 U2126 ( .A(net139849), .B(net105105), .Y(n4363) );
  NAND2XL U2127 ( .A(n3002), .B(net105412), .Y(n10698) );
  MX2X8 U2128 ( .A(\i_MIPS/n236 ), .B(n6646), .S0(n3894), .Y(net112414) );
  AND3XL U2129 ( .A(n7026), .B(n8673), .C(n8890), .Y(n7059) );
  CLKBUFX3 U2130 ( .A(net109512), .Y(n142) );
  CLKINVX1 U2131 ( .A(n9952), .Y(n9946) );
  NAND2X2 U2132 ( .A(DCACHE_addr[1]), .B(n3003), .Y(n9952) );
  AND3X6 U2133 ( .A(net108869), .B(net108854), .C(net108873), .Y(n6701) );
  BUFX8 U2134 ( .A(n6667), .Y(n143) );
  NAND2X8 U2135 ( .A(net144187), .B(\i_MIPS/ID_EX[43] ), .Y(n3785) );
  NAND2X4 U2136 ( .A(\i_MIPS/n234 ), .B(net144187), .Y(n4395) );
  NAND2X4 U2137 ( .A(n3894), .B(n3908), .Y(n4622) );
  BUFX4 U2138 ( .A(n5450), .Y(n5430) );
  OA22X1 U2139 ( .A0(n5256), .A1(n1098), .B0(n5296), .B1(n2721), .Y(n7625) );
  BUFX3 U2140 ( .A(n5305), .Y(n5296) );
  CLKBUFX3 U2141 ( .A(n11208), .Y(n5609) );
  BUFX4 U2142 ( .A(n5609), .Y(n5607) );
  OAI31X4 U2143 ( .A0(n8691), .A1(n8690), .A2(n8889), .B0(n8689), .Y(n8694) );
  AOI222X2 U2144 ( .A0(n4535), .A1(n11491), .B0(mem_rdata_D[115]), .B1(n129), 
        .C0(n5534), .C1(n12994), .Y(n10964) );
  NAND4X4 U2145 ( .A(n11191), .B(n11190), .C(n11189), .D(n11188), .Y(n11366)
         );
  CLKBUFX8 U2146 ( .A(net118223), .Y(net118217) );
  INVX6 U2147 ( .A(n9227), .Y(n9229) );
  OR2X4 U2148 ( .A(n4632), .B(n4631), .Y(n2934) );
  AND2X4 U2149 ( .A(n8970), .B(n8716), .Y(n4631) );
  BUFX4 U2150 ( .A(n10501), .Y(n146) );
  MXI2X1 U2151 ( .A(n10500), .B(n10499), .S0(n5545), .Y(n10501) );
  MXI2X4 U2152 ( .A(n10515), .B(n10514), .S0(n5545), .Y(n10516) );
  AOI222X4 U2153 ( .A0(n4535), .A1(n11493), .B0(mem_rdata_D[117]), .B1(n132), 
        .C0(n12992), .C1(n5534), .Y(n10515) );
  BUFX4 U2154 ( .A(n10801), .Y(n147) );
  MXI2X1 U2155 ( .A(n10800), .B(n10799), .S0(n5549), .Y(n10801) );
  OAI211X2 U2156 ( .A0(\i_MIPS/ALUin1[6] ), .A1(n6707), .B0(\i_MIPS/ALUin1[5] ), .C0(n7222), .Y(n6709) );
  AND2X8 U2157 ( .A(net117723), .B(net117733), .Y(net135423) );
  INVX4 U2158 ( .A(net117723), .Y(n3989) );
  BUFX12 U2159 ( .A(net107195), .Y(net117723) );
  INVX16 U2160 ( .A(net117719), .Y(net117709) );
  OR2X6 U2161 ( .A(n9463), .B(n9462), .Y(n3870) );
  NOR3X6 U2162 ( .A(n3871), .B(n3872), .C(net134673), .Y(n9462) );
  NAND2X2 U2163 ( .A(n10711), .B(net118217), .Y(n3988) );
  INVX4 U2164 ( .A(n3854), .Y(n3727) );
  BUFX12 U2165 ( .A(n3753), .Y(n149) );
  CLKBUFX2 U2166 ( .A(n5261), .Y(n3984) );
  BUFX3 U2167 ( .A(n9809), .Y(n5453) );
  BUFX4 U2168 ( .A(n5449), .Y(n5440) );
  BUFX6 U2169 ( .A(n5402), .Y(n5395) );
  INVX1 U2170 ( .A(n3585), .Y(n3600) );
  INVX3 U2171 ( .A(net114341), .Y(n3589) );
  NAND3X1 U2172 ( .A(\i_MIPS/PC/n7 ), .B(\i_MIPS/PC/n6 ), .C(\i_MIPS/PC/n8 ), 
        .Y(n150) );
  BUFX4 U2173 ( .A(n5449), .Y(n5439) );
  CLKBUFX8 U2174 ( .A(n5307), .Y(n5287) );
  CLKBUFX4 U2175 ( .A(n5751), .Y(n5742) );
  BUFX4 U2176 ( .A(n5884), .Y(n5878) );
  CLKBUFX4 U2177 ( .A(n5261), .Y(n5256) );
  BUFX2 U2178 ( .A(n5841), .Y(n5831) );
  BUFX4 U2179 ( .A(n5921), .Y(n5917) );
  CLKBUFX3 U2180 ( .A(n11209), .Y(n5796) );
  BUFX2 U2181 ( .A(n5307), .Y(n5308) );
  CLKBUFX4 U2182 ( .A(n5307), .Y(n5285) );
  BUFX8 U2183 ( .A(n5406), .Y(n5400) );
  CLKBUFX8 U2184 ( .A(n5450), .Y(n5429) );
  BUFX2 U2185 ( .A(n5453), .Y(n5432) );
  CLKBUFX2 U2186 ( .A(n5306), .Y(n5310) );
  CLKBUFX4 U2187 ( .A(n5306), .Y(n5289) );
  CLKBUFX2 U2188 ( .A(n5265), .Y(n5266) );
  CLKINVX3 U2189 ( .A(n5357), .Y(n3575) );
  BUFX6 U2190 ( .A(n5363), .Y(n5358) );
  CLKBUFX3 U2191 ( .A(n11208), .Y(n5615) );
  CLKBUFX3 U2192 ( .A(n5705), .Y(n5704) );
  CLKINVX1 U2193 ( .A(n5796), .Y(n4832) );
  CLKBUFX4 U2194 ( .A(n5306), .Y(n5291) );
  BUFX16 U2195 ( .A(n5407), .Y(n5403) );
  BUFX4 U2196 ( .A(n5402), .Y(n5396) );
  BUFX3 U2197 ( .A(n5402), .Y(n5394) );
  BUFX8 U2198 ( .A(n5353), .Y(n5357) );
  CLKBUFX3 U2199 ( .A(n5751), .Y(n5741) );
  BUFX4 U2200 ( .A(n5264), .Y(n5251) );
  CLKBUFX3 U2201 ( .A(n5307), .Y(n5309) );
  CLKBUFX4 U2202 ( .A(n5306), .Y(n5290) );
  BUFX4 U2203 ( .A(n5407), .Y(n5404) );
  CLKBUFX3 U2204 ( .A(n135), .Y(n5661) );
  BUFX16 U2205 ( .A(n5220), .Y(n5213) );
  INVX1 U2206 ( .A(net140147), .Y(net114331) );
  INVX4 U2207 ( .A(n3600), .Y(n3601) );
  BUFX3 U2208 ( .A(n5188), .Y(n5186) );
  BUFX4 U2209 ( .A(n5185), .Y(n5176) );
  BUFX8 U2210 ( .A(n5353), .Y(n5356) );
  CLKBUFX3 U2211 ( .A(n5305), .Y(n5298) );
  BUFX16 U2212 ( .A(n5335), .Y(n5330) );
  BUFX12 U2213 ( .A(n5335), .Y(n5331) );
  BUFX8 U2214 ( .A(n3875), .Y(n5332) );
  CLKBUFX3 U2215 ( .A(n10974), .Y(n5542) );
  BUFX8 U2216 ( .A(n5188), .Y(n5184) );
  BUFX8 U2217 ( .A(n5184), .Y(n5179) );
  INVX3 U2218 ( .A(n3604), .Y(n3605) );
  CLKBUFX2 U2219 ( .A(n5453), .Y(n5421) );
  CLKBUFX2 U2220 ( .A(n5453), .Y(n5420) );
  BUFX4 U2221 ( .A(n5609), .Y(n5608) );
  CLKBUFX8 U2222 ( .A(n5267), .Y(n5264) );
  BUFX4 U2223 ( .A(n5884), .Y(n5875) );
  CLKINVX12 U2224 ( .A(n5052), .Y(n3562) );
  BUFX12 U2225 ( .A(n5932), .Y(n5940) );
  CLKBUFX3 U2226 ( .A(net140147), .Y(net114341) );
  BUFX4 U2227 ( .A(n5265), .Y(n5244) );
  BUFX2 U2228 ( .A(n5261), .Y(n5253) );
  BUFX12 U2229 ( .A(n9529), .Y(n5188) );
  BUFX6 U2230 ( .A(n5188), .Y(n5187) );
  BUFX6 U2231 ( .A(n5406), .Y(n5397) );
  BUFX4 U2232 ( .A(n5406), .Y(n5392) );
  BUFX8 U2233 ( .A(n3651), .Y(n5312) );
  BUFX12 U2234 ( .A(n3651), .Y(n5311) );
  INVX4 U2235 ( .A(net134682), .Y(net118379) );
  AND2X2 U2236 ( .A(net105255), .B(net105256), .Y(n151) );
  AND2X2 U2237 ( .A(net104698), .B(net104699), .Y(n152) );
  BUFX4 U2238 ( .A(n4658), .Y(n5707) );
  BUFX4 U2239 ( .A(n5707), .Y(n5696) );
  BUFX12 U2240 ( .A(n5338), .Y(n3875) );
  INVX4 U2241 ( .A(n4836), .Y(n11208) );
  BUFX12 U2242 ( .A(n3965), .Y(DCACHE_addr[3]) );
  BUFX12 U2243 ( .A(n3652), .Y(n5407) );
  CLKBUFX4 U2244 ( .A(n5406), .Y(n5399) );
  BUFX2 U2245 ( .A(n5406), .Y(n5398) );
  BUFX4 U2246 ( .A(n5188), .Y(n5185) );
  BUFX4 U2247 ( .A(n5184), .Y(n5177) );
  CLKBUFX8 U2248 ( .A(n5311), .Y(n5301) );
  CLKBUFX4 U2249 ( .A(n5311), .Y(n5300) );
  INVX3 U2250 ( .A(net118457), .Y(net118455) );
  BUFX16 U2251 ( .A(n5225), .Y(n5221) );
  BUFX20 U2252 ( .A(n5339), .Y(n5354) );
  INVX12 U2253 ( .A(n4018), .Y(n9806) );
  BUFX8 U2254 ( .A(n5336), .Y(n5329) );
  BUFX16 U2255 ( .A(n9809), .Y(n5448) );
  BUFX8 U2256 ( .A(n5448), .Y(n5445) );
  BUFX6 U2257 ( .A(n5448), .Y(n5444) );
  BUFX12 U2258 ( .A(n5311), .Y(n5307) );
  BUFX16 U2259 ( .A(n3652), .Y(n5408) );
  AND2X2 U2260 ( .A(net105075), .B(net105076), .Y(n153) );
  AND2X2 U2261 ( .A(net104939), .B(n3942), .Y(n154) );
  AND2X2 U2262 ( .A(net104889), .B(net104890), .Y(n155) );
  AND2X2 U2263 ( .A(net105264), .B(n3769), .Y(n156) );
  BUFX4 U2264 ( .A(net107617), .Y(net118259) );
  AND2X2 U2265 ( .A(net106602), .B(n3958), .Y(n157) );
  BUFX8 U2266 ( .A(n9505), .Y(n5153) );
  CLKBUFX6 U2267 ( .A(n5087), .Y(n5084) );
  CLKBUFX8 U2268 ( .A(n5087), .Y(n5086) );
  INVX4 U2269 ( .A(net134683), .Y(net118429) );
  INVX4 U2270 ( .A(net118441), .Y(net118423) );
  BUFX4 U2271 ( .A(n5146), .Y(n5150) );
  BUFX6 U2272 ( .A(n5146), .Y(n5149) );
  BUFX16 U2273 ( .A(net115811), .Y(net115797) );
  BUFX8 U2274 ( .A(n5221), .Y(n5215) );
  BUFX8 U2275 ( .A(n9806), .Y(n5263) );
  CLKBUFX3 U2276 ( .A(n5263), .Y(n5257) );
  BUFX2 U2277 ( .A(n5448), .Y(n5452) );
  CLKBUFX3 U2278 ( .A(n5445), .Y(n5436) );
  NAND2X2 U2279 ( .A(n4800), .B(\i_MIPS/PC/n6 ), .Y(n11210) );
  CLKBUFX2 U2280 ( .A(n5763), .Y(n5797) );
  BUFX8 U2281 ( .A(n3965), .Y(n4625) );
  CLKINVX2 U2282 ( .A(n4760), .Y(n5100) );
  NAND2X1 U2283 ( .A(net105110), .B(net105111), .Y(n10539) );
  AND2XL U2284 ( .A(net104916), .B(net104917), .Y(n357) );
  BUFX4 U2285 ( .A(n5080), .Y(n5083) );
  CLKBUFX6 U2286 ( .A(n5080), .Y(n5082) );
  CLKBUFX8 U2287 ( .A(n5080), .Y(n5081) );
  NAND2X6 U2288 ( .A(n6610), .B(n4784), .Y(n4661) );
  BUFX4 U2289 ( .A(net139810), .Y(net117681) );
  AND2X1 U2290 ( .A(net105311), .B(net105312), .Y(n166) );
  BUFX4 U2291 ( .A(n11213), .Y(n5930) );
  BUFX4 U2292 ( .A(n5115), .Y(n5120) );
  AND2X1 U2293 ( .A(net106037), .B(net106038), .Y(n341) );
  INVX6 U2294 ( .A(net134684), .Y(net118453) );
  BUFX8 U2295 ( .A(n5125), .Y(n5127) );
  BUFX6 U2296 ( .A(n5125), .Y(n5128) );
  CLKAND2X4 U2297 ( .A(n4814), .B(n6776), .Y(net134682) );
  BUFX2 U2298 ( .A(n4669), .Y(n5087) );
  BUFX6 U2299 ( .A(n5088), .Y(n5089) );
  BUFX4 U2300 ( .A(n5146), .Y(n5148) );
  BUFX8 U2301 ( .A(n5934), .Y(n5941) );
  INVX16 U2302 ( .A(net36572), .Y(n3634) );
  CLKBUFX8 U2303 ( .A(net115813), .Y(net115789) );
  CLKINVX1 U2304 ( .A(net107169), .Y(net107621) );
  BUFX12 U2305 ( .A(n5363), .Y(n5359) );
  BUFX4 U2306 ( .A(n5197), .Y(n5222) );
  BUFX8 U2307 ( .A(n5221), .Y(n5216) );
  INVX6 U2308 ( .A(n3929), .Y(n9809) );
  CLKBUFX3 U2309 ( .A(n5265), .Y(n5246) );
  CLKBUFX2 U2310 ( .A(n5305), .Y(n5299) );
  CLKINVX1 U2311 ( .A(n5762), .Y(n4829) );
  CLKINVX1 U2312 ( .A(n5788), .Y(n4828) );
  CLKINVX1 U2313 ( .A(n5761), .Y(n4830) );
  INVX3 U2314 ( .A(n5760), .Y(n4831) );
  INVX3 U2315 ( .A(n5184), .Y(n3995) );
  CLKBUFX6 U2316 ( .A(n11535), .Y(n5947) );
  INVX6 U2317 ( .A(n5041), .Y(n5042) );
  AND2XL U2318 ( .A(net105751), .B(net105752), .Y(n1934) );
  INVX4 U2319 ( .A(n5102), .Y(n5099) );
  INVX3 U2320 ( .A(n5102), .Y(n5101) );
  BUFX12 U2321 ( .A(net117703), .Y(net117697) );
  CLKBUFX8 U2322 ( .A(n9502), .Y(n5131) );
  BUFX4 U2323 ( .A(n5131), .Y(n5134) );
  BUFX12 U2324 ( .A(n5139), .Y(n5143) );
  INVX2 U2325 ( .A(net107196), .Y(net117741) );
  BUFX4 U2326 ( .A(net118261), .Y(net118253) );
  CLKBUFX3 U2327 ( .A(net107617), .Y(net118261) );
  AND2XL U2328 ( .A(net105662), .B(net105663), .Y(n337) );
  AND2X2 U2329 ( .A(net105142), .B(net105143), .Y(n338) );
  AND2XL U2330 ( .A(net104985), .B(net119263), .Y(n339) );
  AND2XL U2331 ( .A(net105232), .B(net105233), .Y(n340) );
  BUFX4 U2332 ( .A(n9506), .Y(n5158) );
  AND2X2 U2333 ( .A(net104792), .B(net104793), .Y(n342) );
  CLKBUFX6 U2334 ( .A(n4669), .Y(n5085) );
  INVX3 U2335 ( .A(n6452), .Y(n11037) );
  INVX3 U2336 ( .A(n6459), .Y(n11049) );
  OAI221X2 U2337 ( .A0(n5171), .A1(n1331), .B0(n5222), .B1(n2984), .C0(n6458), 
        .Y(n6459) );
  BUFX12 U2338 ( .A(n5936), .Y(n5939) );
  BUFX4 U2339 ( .A(n5126), .Y(n5129) );
  BUFX4 U2340 ( .A(n5146), .Y(n5147) );
  CLKINVX1 U2341 ( .A(net107168), .Y(net107615) );
  AND2X4 U2342 ( .A(n11053), .B(\i_MIPS/n497 ), .Y(n348) );
  INVX12 U2343 ( .A(n10721), .Y(n11054) );
  INVX8 U2344 ( .A(n4016), .Y(n9807) );
  BUFX6 U2345 ( .A(n5408), .Y(n5402) );
  INVX6 U2346 ( .A(\i_MIPS/n506 ), .Y(n6016) );
  NAND2X1 U2347 ( .A(DCACHE_addr[2]), .B(n11507), .Y(n350) );
  NAND2X4 U2348 ( .A(n3703), .B(\i_MIPS/n301 ), .Y(net108297) );
  AND2X1 U2349 ( .A(net108876), .B(net108869), .Y(n351) );
  AND2X2 U2350 ( .A(n10111), .B(n10110), .Y(n354) );
  NAND2X6 U2351 ( .A(n4675), .B(n348), .Y(net139810) );
  BUFX6 U2352 ( .A(net117683), .Y(net117673) );
  CLKBUFX8 U2353 ( .A(net117683), .Y(net117675) );
  CLKBUFX3 U2354 ( .A(net139810), .Y(net117683) );
  NAND3X6 U2355 ( .A(n3740), .B(n3741), .C(net107519), .Y(net106031) );
  INVX4 U2356 ( .A(n4758), .Y(n5105) );
  INVX4 U2357 ( .A(n4758), .Y(n5103) );
  INVX6 U2358 ( .A(n3903), .Y(net114065) );
  AND2X2 U2359 ( .A(n11538), .B(net118581), .Y(n428) );
  INVX16 U2360 ( .A(n5041), .Y(n5044) );
  CLKBUFX3 U2361 ( .A(net134686), .Y(net118417) );
  BUFX4 U2362 ( .A(n5141), .Y(n5145) );
  INVX3 U2363 ( .A(net107167), .Y(net107617) );
  MXI2X2 U2364 ( .A(n10976), .B(n10975), .S0(n5549), .Y(n10977) );
  NAND2X4 U2365 ( .A(n3903), .B(n3674), .Y(n8699) );
  CLKBUFX3 U2366 ( .A(net134680), .Y(net118313) );
  CLKBUFX3 U2367 ( .A(net134680), .Y(net118321) );
  INVX20 U2368 ( .A(n5065), .Y(n5064) );
  BUFX4 U2369 ( .A(net135423), .Y(net117719) );
  CLKBUFX3 U2370 ( .A(net135423), .Y(net117715) );
  BUFX4 U2371 ( .A(n4661), .Y(n5080) );
  BUFX20 U2372 ( .A(n12980), .Y(DCACHE_addr[1]) );
  BUFX4 U2373 ( .A(n11214), .Y(n5937) );
  BUFX2 U2374 ( .A(n5937), .Y(n5933) );
  BUFX4 U2375 ( .A(net118243), .Y(net118235) );
  INVX12 U2376 ( .A(n1329), .Y(DCACHE_addr[14]) );
  BUFX8 U2377 ( .A(n4660), .Y(n5078) );
  BUFX12 U2378 ( .A(n4755), .Y(n5069) );
  BUFX8 U2379 ( .A(n9500), .Y(n5121) );
  BUFX4 U2380 ( .A(n5121), .Y(n5123) );
  NAND4X4 U2381 ( .A(n4826), .B(n4827), .C(\i_MIPS/EX_MEM_0 ), .D(n6643), .Y(
        net107195) );
  BUFX4 U2382 ( .A(n9505), .Y(n5151) );
  BUFX6 U2383 ( .A(n9536), .Y(n5189) );
  AND4X8 U2384 ( .A(\i_MIPS/ALUOp[1] ), .B(n3622), .C(n3908), .D(n6646), .Y(
        n1340) );
  BUFX16 U2385 ( .A(n4756), .Y(n5074) );
  INVX2 U2386 ( .A(net112446), .Y(n3902) );
  INVX3 U2387 ( .A(n7889), .Y(n9501) );
  CLKINVX1 U2388 ( .A(net107170), .Y(net107619) );
  BUFX4 U2389 ( .A(net118297), .Y(net118291) );
  INVX4 U2390 ( .A(n11344), .Y(n11537) );
  CLKBUFX4 U2391 ( .A(n5197), .Y(n5220) );
  INVX8 U2392 ( .A(n10736), .Y(n11056) );
  BUFX12 U2393 ( .A(n9808), .Y(n5339) );
  CLKBUFX2 U2394 ( .A(n5399), .Y(n5381) );
  NAND2XL U2395 ( .A(ICACHE_addr[4]), .B(n11345), .Y(n1856) );
  NAND2X1 U2396 ( .A(n5947), .B(n11378), .Y(n1857) );
  NAND2X1 U2397 ( .A(n5947), .B(n11379), .Y(n1858) );
  NAND2X1 U2398 ( .A(n5947), .B(n11380), .Y(n1859) );
  NAND2X1 U2399 ( .A(n5947), .B(n11381), .Y(n1860) );
  NAND2X1 U2400 ( .A(n5947), .B(n11382), .Y(n1861) );
  NAND2X1 U2401 ( .A(n5947), .B(n11383), .Y(n1862) );
  NAND2X1 U2402 ( .A(n5947), .B(n11384), .Y(n1863) );
  NAND2X1 U2403 ( .A(n5947), .B(n11385), .Y(n1864) );
  NAND2X1 U2404 ( .A(n5947), .B(n11386), .Y(n1865) );
  NAND2X1 U2405 ( .A(n5947), .B(n11388), .Y(n1866) );
  NAND2X1 U2406 ( .A(n5947), .B(n11389), .Y(n1867) );
  NAND2X1 U2407 ( .A(n5947), .B(n11392), .Y(n1868) );
  NAND2X1 U2408 ( .A(n5947), .B(n11393), .Y(n1869) );
  NAND2X1 U2409 ( .A(n5947), .B(n11394), .Y(n1870) );
  NAND2X1 U2410 ( .A(n5947), .B(n11395), .Y(n1871) );
  NAND2X1 U2411 ( .A(n5947), .B(n11396), .Y(n1872) );
  NAND2X1 U2412 ( .A(n5947), .B(n11397), .Y(n1873) );
  NAND2X1 U2413 ( .A(n5947), .B(n11398), .Y(n1874) );
  NAND2X1 U2414 ( .A(n5947), .B(n11399), .Y(n1875) );
  NAND2X1 U2415 ( .A(n5947), .B(n11404), .Y(n1876) );
  NAND2X1 U2416 ( .A(n5042), .B(n11429), .Y(n1877) );
  NAND2X1 U2417 ( .A(n5042), .B(n11432), .Y(n1878) );
  NAND2X1 U2418 ( .A(n5044), .B(n11434), .Y(n1879) );
  NAND2X1 U2419 ( .A(n5042), .B(n11435), .Y(n1880) );
  NAND2XL U2420 ( .A(n5044), .B(n11437), .Y(n1881) );
  NAND2X1 U2421 ( .A(n5042), .B(n11438), .Y(n1882) );
  NAND2X1 U2422 ( .A(n5044), .B(n11440), .Y(n1883) );
  NAND2X1 U2423 ( .A(n5042), .B(n11441), .Y(n1884) );
  NAND2X1 U2424 ( .A(n5043), .B(n11445), .Y(n1885) );
  NAND2X1 U2425 ( .A(n5042), .B(n11447), .Y(n1886) );
  NAND2X1 U2426 ( .A(n5043), .B(n11448), .Y(n1887) );
  NAND2X1 U2427 ( .A(n5044), .B(n11449), .Y(n1888) );
  NAND2XL U2428 ( .A(n5042), .B(n11450), .Y(n1889) );
  NAND2X1 U2429 ( .A(n5043), .B(n11451), .Y(n1890) );
  NAND2X1 U2430 ( .A(n5044), .B(n11452), .Y(n1891) );
  NAND2XL U2431 ( .A(n5042), .B(n11453), .Y(n1892) );
  NAND2X1 U2432 ( .A(n5043), .B(n11454), .Y(n1893) );
  NAND2X1 U2433 ( .A(n5042), .B(n11456), .Y(n1894) );
  NAND2X1 U2434 ( .A(n5043), .B(n11457), .Y(n1895) );
  NAND2X1 U2435 ( .A(n5042), .B(n11459), .Y(n1896) );
  NAND2X1 U2436 ( .A(n5043), .B(n11460), .Y(n1897) );
  NAND2X1 U2437 ( .A(n5044), .B(n11461), .Y(n1898) );
  NAND2X1 U2438 ( .A(n5043), .B(n11463), .Y(n1899) );
  NAND2X1 U2439 ( .A(n5044), .B(n11464), .Y(n1900) );
  NAND2X1 U2440 ( .A(n5044), .B(n11467), .Y(n1901) );
  NAND2X1 U2441 ( .A(n5042), .B(n11468), .Y(n1902) );
  NAND2X1 U2442 ( .A(n5043), .B(n11469), .Y(n1903) );
  NAND2X1 U2443 ( .A(n5044), .B(n11470), .Y(n1904) );
  NAND2X1 U2444 ( .A(n5042), .B(n11471), .Y(n1905) );
  NAND2X1 U2445 ( .A(n5043), .B(n11472), .Y(n1906) );
  NAND2X1 U2446 ( .A(n5044), .B(n11473), .Y(n1907) );
  NAND2X1 U2447 ( .A(n5042), .B(n11474), .Y(n1908) );
  NAND2X1 U2448 ( .A(n5043), .B(n11475), .Y(n1909) );
  NAND2X1 U2449 ( .A(n5042), .B(n11477), .Y(n1910) );
  NAND2X1 U2450 ( .A(n5042), .B(n11480), .Y(n1911) );
  NAND2X1 U2451 ( .A(n5042), .B(n11483), .Y(n1912) );
  NAND2XL U2452 ( .A(n5043), .B(n11484), .Y(n1913) );
  NAND2X1 U2453 ( .A(n5044), .B(n11485), .Y(n1914) );
  NAND2X1 U2454 ( .A(n5042), .B(n11486), .Y(n1915) );
  NAND2X1 U2455 ( .A(n5043), .B(n11487), .Y(n1916) );
  NAND2X1 U2456 ( .A(n5044), .B(n11488), .Y(n1917) );
  NAND2X1 U2457 ( .A(n5042), .B(n11489), .Y(n1918) );
  NAND2X1 U2458 ( .A(n5043), .B(n11490), .Y(n1919) );
  NAND2X1 U2459 ( .A(n5044), .B(n11491), .Y(n1920) );
  NAND2X1 U2460 ( .A(n5042), .B(n11492), .Y(n1921) );
  NAND2X1 U2461 ( .A(n5042), .B(n11495), .Y(n1922) );
  NAND2X1 U2462 ( .A(n5044), .B(n11497), .Y(n1923) );
  NAND2X1 U2463 ( .A(n5042), .B(n11498), .Y(n1924) );
  NAND2X1 U2464 ( .A(n5947), .B(n11500), .Y(n1925) );
  NAND2X1 U2465 ( .A(n5043), .B(n11502), .Y(n1926) );
  NAND2XL U2466 ( .A(n5055), .B(n11507), .Y(n1927) );
  NOR2X1 U2467 ( .A(n4404), .B(n4405), .Y(n1928) );
  NOR2X1 U2468 ( .A(n4408), .B(n4409), .Y(n1929) );
  OR2X1 U2469 ( .A(n5040), .B(n9940), .Y(n4932) );
  NOR2XL U2470 ( .A(n5040), .B(n10391), .Y(n1930) );
  AND2X2 U2471 ( .A(net104866), .B(net104867), .Y(n1933) );
  AND2X2 U2472 ( .A(net105490), .B(net105491), .Y(n1935) );
  AND2XL U2473 ( .A(net105008), .B(net105009), .Y(n1936) );
  AND2X2 U2474 ( .A(net105423), .B(n3955), .Y(n1937) );
  AND2X2 U2475 ( .A(n8633), .B(n11101), .Y(n1939) );
  AND2XL U2476 ( .A(n9223), .B(n9222), .Y(n1940) );
  BUFX16 U2477 ( .A(n4683), .Y(n5539) );
  NAND2X1 U2478 ( .A(n5951), .B(n11220), .Y(n1950) );
  NAND2X1 U2479 ( .A(n5951), .B(n11221), .Y(n1951) );
  NAND2X1 U2480 ( .A(n5951), .B(n11222), .Y(n1952) );
  NAND2X1 U2481 ( .A(n5951), .B(n11223), .Y(n1953) );
  NAND2X1 U2482 ( .A(n5951), .B(n11224), .Y(n1954) );
  NAND2X1 U2483 ( .A(n5951), .B(n11225), .Y(n1955) );
  NAND2X1 U2484 ( .A(n5951), .B(n11226), .Y(n1956) );
  NAND2X1 U2485 ( .A(n5951), .B(n11227), .Y(n1957) );
  NAND2X1 U2486 ( .A(n5951), .B(n11228), .Y(n1958) );
  NAND2X1 U2487 ( .A(n5951), .B(n11229), .Y(n1959) );
  NAND2X1 U2488 ( .A(n5951), .B(n11230), .Y(n1960) );
  NAND2X1 U2489 ( .A(n5951), .B(n11231), .Y(n1961) );
  NAND2X1 U2490 ( .A(n5951), .B(n11232), .Y(n1962) );
  NAND2X1 U2491 ( .A(n5951), .B(n11233), .Y(n1963) );
  NAND2X1 U2492 ( .A(n5951), .B(n11234), .Y(n1964) );
  NAND2X1 U2493 ( .A(n5951), .B(n11235), .Y(n1965) );
  NAND2X1 U2494 ( .A(n5951), .B(n11236), .Y(n1966) );
  NAND2X1 U2495 ( .A(n5951), .B(net103849), .Y(n1967) );
  NAND2X1 U2496 ( .A(n5951), .B(n11237), .Y(n1968) );
  NAND2X1 U2497 ( .A(n5951), .B(n11238), .Y(n1969) );
  NAND2X1 U2498 ( .A(n5951), .B(n11239), .Y(n1970) );
  NAND2X1 U2499 ( .A(n5951), .B(n11240), .Y(n1971) );
  NAND2X1 U2500 ( .A(n5951), .B(n11241), .Y(n1972) );
  NAND2X1 U2501 ( .A(n5951), .B(n11242), .Y(n1973) );
  NAND2X1 U2502 ( .A(n5951), .B(n11243), .Y(n1974) );
  NAND2X1 U2503 ( .A(n5951), .B(n11244), .Y(n1975) );
  NAND2X1 U2504 ( .A(n5951), .B(n11245), .Y(n1976) );
  NAND2X1 U2505 ( .A(n5951), .B(n11246), .Y(n1977) );
  NAND2X1 U2506 ( .A(n5951), .B(n11247), .Y(n1978) );
  NAND2X1 U2507 ( .A(n5951), .B(n11248), .Y(n1979) );
  NAND2X1 U2508 ( .A(n5951), .B(n11249), .Y(n1980) );
  NAND2X1 U2509 ( .A(n5951), .B(n11250), .Y(n1981) );
  NAND2X1 U2510 ( .A(n5951), .B(n11251), .Y(n1982) );
  NAND2X1 U2511 ( .A(n5951), .B(n11252), .Y(n1983) );
  NAND2X1 U2512 ( .A(n5042), .B(n11426), .Y(n1984) );
  AOI22X2 U2513 ( .A0(n12966), .A1(n11534), .B0(n5947), .B1(n11521), .Y(n1985)
         );
  AND2X2 U2514 ( .A(net106674), .B(n4013), .Y(n1986) );
  AND2XL U2515 ( .A(net105334), .B(net105335), .Y(n1987) );
  CLKINVX1 U2516 ( .A(n128), .Y(net107659) );
  INVX1 U2517 ( .A(n10), .Y(n3896) );
  BUFX16 U2518 ( .A(n12962), .Y(DCACHE_addr[21]) );
  INVX3 U2519 ( .A(net118481), .Y(net118479) );
  INVX4 U2520 ( .A(net118345), .Y(net118327) );
  INVX6 U2521 ( .A(net118341), .Y(net118331) );
  INVX4 U2522 ( .A(net118343), .Y(net118329) );
  AND3XL U2523 ( .A(n9425), .B(n3950), .C(n6960), .Y(n2330) );
  AND2X4 U2524 ( .A(n6770), .B(n4720), .Y(net134684) );
  CLKBUFX3 U2525 ( .A(net134684), .Y(net118457) );
  AND2X2 U2526 ( .A(\i_MIPS/control_out[6] ), .B(net118581), .Y(n2894) );
  AND2X2 U2527 ( .A(net105288), .B(n3953), .Y(n2896) );
  AND2X2 U2528 ( .A(\i_MIPS/control_out[0] ), .B(net118581), .Y(n2899) );
  INVX3 U2529 ( .A(n6429), .Y(n11014) );
  MXI2X2 U2530 ( .A(n10208), .B(n10207), .S0(n5543), .Y(n10209) );
  AND2X2 U2531 ( .A(n4786), .B(n4722), .Y(n4758) );
  CLKBUFX3 U2532 ( .A(n4759), .Y(n5097) );
  NAND2X4 U2533 ( .A(n6610), .B(n4786), .Y(n4669) );
  CLKBUFX3 U2534 ( .A(net107615), .Y(net118241) );
  CLKBUFX3 U2535 ( .A(n4662), .Y(n5090) );
  NAND2X4 U2536 ( .A(n6610), .B(n4721), .Y(n4662) );
  CLKBUFX4 U2537 ( .A(n4662), .Y(n5091) );
  OAI221X4 U2538 ( .A0(\i_MIPS/n270 ), .A1(n5073), .B0(\i_MIPS/n271 ), .B1(
        n5068), .C0(n6663), .Y(n9049) );
  AOI22X4 U2539 ( .A0(net118215), .A1(net105313), .B0(net118225), .B1(n6792), 
        .Y(n2938) );
  OAI22X2 U2540 ( .A0(n10634), .A1(n3766), .B0(n9536), .B1(n10637), .Y(n2950)
         );
  CLKBUFX3 U2541 ( .A(net139810), .Y(net117685) );
  INVX8 U2542 ( .A(net117741), .Y(net117731) );
  NAND2X1 U2543 ( .A(n6951), .B(n3861), .Y(n7669) );
  BUFX12 U2544 ( .A(net139756), .Y(net117703) );
  BUFX4 U2545 ( .A(net117703), .Y(net117695) );
  BUFX16 U2546 ( .A(n5114), .Y(n5119) );
  BUFX3 U2547 ( .A(n9506), .Y(n5154) );
  BUFX12 U2548 ( .A(n5155), .Y(n5157) );
  BUFX4 U2549 ( .A(n9506), .Y(n5155) );
  OR2X6 U2550 ( .A(n8869), .B(n8872), .Y(n2993) );
  AND2X2 U2551 ( .A(n4814), .B(n348), .Y(net134680) );
  CLKBUFX3 U2552 ( .A(net134680), .Y(net118319) );
  CLKBUFX3 U2553 ( .A(n9501), .Y(n5126) );
  BUFX4 U2554 ( .A(n9501), .Y(n5125) );
  AND2X2 U2555 ( .A(n4814), .B(n4720), .Y(net134681) );
  CLKBUFX3 U2556 ( .A(net134681), .Y(net118369) );
  BUFX4 U2557 ( .A(n5142), .Y(n5140) );
  BUFX4 U2558 ( .A(net107621), .Y(net118295) );
  BUFX4 U2559 ( .A(net134686), .Y(net118409) );
  INVX3 U2560 ( .A(n7885), .Y(n9505) );
  MXI2X4 U2561 ( .A(n10620), .B(n10621), .S0(n4410), .Y(n2995) );
  AND2X6 U2562 ( .A(n4700), .B(n7100), .Y(n2996) );
  BUFX16 U2563 ( .A(n12960), .Y(DCACHE_addr[23]) );
  BUFX16 U2564 ( .A(n12968), .Y(DCACHE_addr[15]) );
  CLKAND2X8 U2565 ( .A(n6388), .B(n6389), .Y(n2999) );
  CLKAND2X8 U2566 ( .A(n4704), .B(n6918), .Y(n3776) );
  OR2X8 U2567 ( .A(n4444), .B(n4443), .Y(n3000) );
  BUFX4 U2568 ( .A(n5937), .Y(n5936) );
  CLKAND2X8 U2569 ( .A(n4719), .B(n9944), .Y(n4685) );
  CLKBUFX8 U2570 ( .A(n4685), .Y(n5534) );
  AOI22X4 U2571 ( .A0(n3625), .A1(net118217), .B0(net118225), .B1(n7099), .Y(
        n3002) );
  BUFX16 U2572 ( .A(n12981), .Y(DCACHE_addr[0]) );
  AOI22X4 U2573 ( .A0(net118215), .A1(net105336), .B0(net118227), .B1(n8420), 
        .Y(n3004) );
  NAND2X2 U2574 ( .A(n4675), .B(n4720), .Y(net139719) );
  BUFX4 U2575 ( .A(net117647), .Y(net117641) );
  BUFX4 U2576 ( .A(n11050), .Y(n5552) );
  CLKAND2X8 U2577 ( .A(n4719), .B(n4689), .Y(n4684) );
  CLKINVX1 U2578 ( .A(net108297), .Y(net108308) );
  AND3X4 U2579 ( .A(n4627), .B(n4628), .C(n6489), .Y(n3005) );
  BUFX8 U2580 ( .A(n4756), .Y(n5075) );
  AND2X2 U2581 ( .A(n4784), .B(n4722), .Y(n4760) );
  AND2X4 U2582 ( .A(n6770), .B(n4785), .Y(net134683) );
  MXI2X2 U2583 ( .A(n10687), .B(n10688), .S0(n4410), .Y(n3014) );
  MXI2X4 U2584 ( .A(n10700), .B(n10699), .S0(n5549), .Y(n10701) );
  MXI2X4 U2585 ( .A(n10895), .B(n10894), .S0(n5545), .Y(n10896) );
  NAND3X4 U2586 ( .A(n3716), .B(n3717), .C(n7152), .Y(n7422) );
  AOI22X4 U2587 ( .A0(net118225), .A1(n6892), .B0(net118217), .B1(net105290), 
        .Y(n3015) );
  NAND2X6 U2588 ( .A(net135522), .B(n10717), .Y(n3016) );
  CLKBUFX8 U2589 ( .A(n4755), .Y(n5070) );
  BUFX16 U2590 ( .A(n12958), .Y(DCACHE_addr[25]) );
  BUFX16 U2591 ( .A(n12972), .Y(DCACHE_addr[11]) );
  AND3X8 U2592 ( .A(n3643), .B(n3644), .C(net109042), .Y(n3021) );
  AND3X8 U2593 ( .A(n3727), .B(n9298), .C(n9303), .Y(n3022) );
  AOI22X4 U2594 ( .A0(n3683), .A1(net118217), .B0(net118227), .B1(n7003), .Y(
        n3023) );
  AND3X6 U2595 ( .A(n3729), .B(n3730), .C(n8702), .Y(n3024) );
  AND3X8 U2596 ( .A(n3962), .B(n3963), .C(n7837), .Y(n3025) );
  AND3X2 U2597 ( .A(n4690), .B(n4692), .C(n7486), .Y(n3026) );
  AND3X8 U2598 ( .A(n3986), .B(n3987), .C(n3988), .Y(n3027) );
  BUFX8 U2599 ( .A(net117751), .Y(net117743) );
  AOI222XL U2600 ( .A0(n5541), .A1(n11419), .B0(mem_rdata_D[43]), .B1(n131), 
        .C0(n13002), .C1(n5540), .Y(n10794) );
  NAND2X1 U2601 ( .A(n3964), .B(n3621), .Y(n3029) );
  CLKINVX1 U2602 ( .A(n10979), .Y(n10974) );
  INVX3 U2603 ( .A(n7886), .Y(n9504) );
  CLKBUFX8 U2604 ( .A(n3633), .Y(net115811) );
  INVX6 U2605 ( .A(n11374), .Y(n3788) );
  AOI22X1 U2606 ( .A0(n7685), .A1(n9445), .B0(n7684), .B1(n9442), .Y(n3030) );
  NAND2X6 U2607 ( .A(n12), .B(n3874), .Y(net112549) );
  NAND3X4 U2608 ( .A(n3687), .B(n3688), .C(n8216), .Y(net105234) );
  INVX12 U2609 ( .A(net118227), .Y(n3890) );
  INVX12 U2610 ( .A(net118592), .Y(net107657) );
  CLKINVX3 U2611 ( .A(n5211), .Y(n5204) );
  INVX16 U2612 ( .A(n355), .Y(DCACHE_addr[5]) );
  CLKBUFX2 U2613 ( .A(n5615), .Y(n5583) );
  INVX3 U2614 ( .A(n5420), .Y(n5418) );
  INVX4 U2615 ( .A(n11380), .Y(n3979) );
  BUFX4 U2616 ( .A(n5184), .Y(n5180) );
  AND2X2 U2617 ( .A(n10979), .B(mem_ready_D), .Y(n3031) );
  CLKBUFX2 U2618 ( .A(n5406), .Y(n5374) );
  BUFX8 U2619 ( .A(n5337), .Y(n5324) );
  AND2X2 U2620 ( .A(\i_MIPS/control_out[7] ), .B(net118581), .Y(n3032) );
  INVX16 U2621 ( .A(n4825), .Y(DCACHE_addr[20]) );
  INVX16 U2622 ( .A(n4824), .Y(DCACHE_addr[26]) );
  INVX16 U2623 ( .A(n5005), .Y(DCACHE_addr[12]) );
  INVX16 U2624 ( .A(n1303), .Y(DCACHE_addr[10]) );
  NAND2X4 U2625 ( .A(net104791), .B(net139850), .Y(n4328) );
  CLKINVX6 U2626 ( .A(net104343), .Y(net109359) );
  NOR3X4 U2627 ( .A(n4484), .B(n4485), .C(n4486), .Y(n9794) );
  NOR2BX2 U2628 ( .AN(net104171), .B(n3809), .Y(n4484) );
  NOR2BX2 U2629 ( .AN(net104171), .B(n3810), .Y(n4475) );
  NOR3X4 U2630 ( .A(n4475), .B(n4476), .C(n4477), .Y(n9889) );
  AOI222X2 U2631 ( .A0(net104171), .A1(n11239), .B0(n3663), .B1(n11270), .C0(
        net104173), .C1(n11301), .Y(n10005) );
  OAI221X1 U2632 ( .A0(n10006), .A1(net143858), .B0(\i_MIPS/n500 ), .B1(
        net115793), .C0(n10005), .Y(\i_MIPS/N70 ) );
  INVX4 U2633 ( .A(n12872), .Y(n4119) );
  INVX4 U2634 ( .A(n12866), .Y(n4135) );
  INVX4 U2635 ( .A(n12863), .Y(n4842) );
  CLKAND2X2 U2636 ( .A(net104171), .B(n11243), .Y(n4487) );
  CLKAND2X2 U2637 ( .A(net104172), .B(n11253), .Y(n4465) );
  CLKAND2X2 U2638 ( .A(n3663), .B(n11276), .Y(n4462) );
  CLKAND2X2 U2639 ( .A(net104172), .B(n11279), .Y(n4468) );
  CLKAND2X2 U2640 ( .A(n3663), .B(n11277), .Y(n4491) );
  CLKAND2X2 U2641 ( .A(n3663), .B(n11254), .Y(n4429) );
  CLKAND2X2 U2642 ( .A(net104172), .B(n11262), .Y(n4480) );
  CLKAND2X2 U2643 ( .A(net104172), .B(n11259), .Y(n4476) );
  CLKAND2X2 U2644 ( .A(net104172), .B(n11269), .Y(n4485) );
  NOR2BX2 U2645 ( .AN(net104171), .B(n3799), .Y(n4449) );
  CLKAND2X2 U2646 ( .A(n3898), .B(n11286), .Y(n4479) );
  AO22X4 U2647 ( .A0(mem_rdata_I[51]), .A1(n5941), .B0(n5568), .B1(n11268), 
        .Y(n11074) );
  NAND2X6 U2648 ( .A(n4372), .B(n4373), .Y(n6724) );
  NAND2X2 U2649 ( .A(n4782), .B(n3894), .Y(n4373) );
  INVX8 U2650 ( .A(net105121), .Y(net110799) );
  CLKINVX1 U2651 ( .A(n8668), .Y(n3557) );
  INVX1 U2652 ( .A(n8121), .Y(n8668) );
  INVX1 U2653 ( .A(n7404), .Y(n7406) );
  INVX4 U2654 ( .A(n9316), .Y(n8208) );
  INVXL U2655 ( .A(n8202), .Y(n8639) );
  CLKINVX1 U2656 ( .A(net144236), .Y(n3584) );
  CLKAND2X3 U2657 ( .A(n4690), .B(n7486), .Y(n4705) );
  NAND2X4 U2658 ( .A(n6819), .B(n3784), .Y(n8890) );
  NAND2X6 U2659 ( .A(n7028), .B(n3983), .Y(n7429) );
  INVX12 U2660 ( .A(n7775), .Y(n6695) );
  INVX12 U2661 ( .A(n5194), .Y(n5191) );
  MXI2X2 U2662 ( .A(n10408), .B(n10407), .S0(n5544), .Y(n10409) );
  AOI222X4 U2663 ( .A0(n4505), .A1(n11460), .B0(mem_rdata_D[84]), .B1(n133), 
        .C0(n12993), .C1(n5535), .Y(n10408) );
  OR2X6 U2664 ( .A(n6954), .B(n6953), .Y(n9432) );
  NAND2X1 U2665 ( .A(net106297), .B(net106298), .Y(n9938) );
  NAND2X1 U2666 ( .A(DCACHE_addr[4]), .B(n5190), .Y(net106297) );
  NAND3X1 U2667 ( .A(n7868), .B(n3950), .C(n7860), .Y(n7873) );
  AO22XL U2668 ( .A0(net134673), .A1(n7868), .B0(n7841), .B1(net107404), .Y(
        n7854) );
  AOI33X2 U2669 ( .A0(n7870), .A1(n7869), .A2(n3950), .B0(net117743), .B1(
        n7868), .B2(n7867), .Y(n7871) );
  CLKINVX1 U2670 ( .A(n1940), .Y(n3560) );
  INVX1 U2671 ( .A(n8044), .Y(n8468) );
  NAND2X8 U2672 ( .A(n6702), .B(n2920), .Y(n8044) );
  INVX3 U2673 ( .A(n5209), .Y(n5207) );
  MX2X1 U2674 ( .A(\D_cache/cache[0][68] ), .B(n10757), .S0(n5167), .Y(
        \D_cache/n1252 ) );
  INVX3 U2675 ( .A(n5169), .Y(n5167) );
  INVX3 U2676 ( .A(n5376), .Y(n5372) );
  CLKBUFX2 U2677 ( .A(n5406), .Y(n5376) );
  MX2X1 U2678 ( .A(\D_cache/cache[6][3] ), .B(n4561), .S0(n3574), .Y(
        \D_cache/n1766 ) );
  MX2X1 U2679 ( .A(\D_cache/cache[6][68] ), .B(n10757), .S0(n3574), .Y(
        \D_cache/n1246 ) );
  MX2X1 U2680 ( .A(\D_cache/cache[5][3] ), .B(n4561), .S0(n5349), .Y(
        \D_cache/n1767 ) );
  MX2X1 U2681 ( .A(\D_cache/cache[5][68] ), .B(n10757), .S0(n5349), .Y(
        \D_cache/n1247 ) );
  INVX3 U2682 ( .A(n5351), .Y(n5349) );
  MX2X1 U2683 ( .A(\D_cache/cache[4][3] ), .B(n4561), .S0(n3763), .Y(
        \D_cache/n1768 ) );
  MX2X1 U2684 ( .A(\D_cache/cache[4][68] ), .B(n10757), .S0(n3763), .Y(
        \D_cache/n1248 ) );
  MX2X1 U2685 ( .A(\I_cache/cache[7][97] ), .B(n10883), .S0(n5849), .Y(n12062)
         );
  INVX1 U2686 ( .A(net108623), .Y(net107828) );
  NAND3BX2 U2687 ( .AN(n9731), .B(net115797), .C(n9730), .Y(n9729) );
  NAND4X1 U2688 ( .A(\i_MIPS/n517 ), .B(\i_MIPS/n519 ), .C(\i_MIPS/n520 ), .D(
        n9602), .Y(n9730) );
  NAND2X1 U2689 ( .A(n3977), .B(\i_MIPS/n271 ), .Y(n9541) );
  NAND3X2 U2690 ( .A(n10155), .B(n10157), .C(n10156), .Y(n10256) );
  NAND2X1 U2691 ( .A(\i_MIPS/IF_ID[6] ), .B(n168), .Y(n10157) );
  INVX1 U2692 ( .A(n5439), .Y(n3561) );
  AO22X1 U2693 ( .A0(ICACHE_addr[16]), .A1(mem_read_I), .B0(mem_write_I), .B1(
        n11358), .Y(n12868) );
  NAND3X4 U2694 ( .A(ICACHE_addr[16]), .B(ICACHE_addr[15]), .C(n10301), .Y(
        n10323) );
  XOR2X1 U2695 ( .A(n11358), .B(ICACHE_addr[16]), .Y(n11592) );
  AO22X2 U2696 ( .A0(n5939), .A1(ICACHE_addr[16]), .B0(n5931), .B1(n11358), 
        .Y(n11140) );
  MXI2X2 U2697 ( .A(n10524), .B(n10523), .S0(n5546), .Y(n10525) );
  MXI2X2 U2698 ( .A(n10552), .B(n10551), .S0(n5546), .Y(n10553) );
  OAI221X4 U2699 ( .A0(n10161), .A1(n5562), .B0(n5557), .B1(n10162), .C0(
        n10160), .Y(\i_MIPS/PC/n43 ) );
  OAI221X4 U2700 ( .A0(n10337), .A1(n5561), .B0(n5557), .B1(n10338), .C0(
        n10336), .Y(\i_MIPS/PC/n55 ) );
  MXI2X2 U2701 ( .A(n10503), .B(n10502), .S0(n5545), .Y(n10504) );
  MXI2X2 U2702 ( .A(n10448), .B(n10447), .S0(n5545), .Y(n10449) );
  MXI2X1 U2703 ( .A(n10463), .B(n10462), .S0(n5545), .Y(n10464) );
  MXI2X1 U2704 ( .A(n10509), .B(n10508), .S0(n5545), .Y(n10510) );
  BUFX16 U2705 ( .A(n12964), .Y(DCACHE_addr[19]) );
  BUFX16 U2706 ( .A(n12975), .Y(DCACHE_addr[8]) );
  AND2X2 U2707 ( .A(DCACHE_addr[7]), .B(n11534), .Y(n4408) );
  BUFX16 U2708 ( .A(n12976), .Y(DCACHE_addr[7]) );
  CLKMX2X2 U2709 ( .A(n10643), .B(n10644), .S0(n4410), .Y(n3822) );
  CLKMX2X4 U2710 ( .A(n10656), .B(n10657), .S0(n4410), .Y(n3823) );
  CLKMX2X4 U2711 ( .A(n10601), .B(n10602), .S0(n4410), .Y(n3824) );
  CLKMX2X4 U2712 ( .A(n10186), .B(n10187), .S0(n4410), .Y(n3821) );
  INVX3 U2713 ( .A(n5548), .Y(n4410) );
  AO22X2 U2714 ( .A0(n5554), .A1(n12959), .B0(n5551), .B1(n11528), .Y(n11004)
         );
  INVX1 U2715 ( .A(n5180), .Y(n3564) );
  CLKINVX1 U2716 ( .A(n5180), .Y(n3565) );
  BUFX16 U2717 ( .A(n12955), .Y(DCACHE_addr[28]) );
  INVX12 U2718 ( .A(n1927), .Y(mem_addr_D[6]) );
  CLKINVX1 U2719 ( .A(n12879), .Y(n3567) );
  INVX12 U2720 ( .A(n3567), .Y(mem_addr_I[5]) );
  AND2X1 U2721 ( .A(ICACHE_addr[3]), .B(n11345), .Y(n12879) );
  CLKAND2X12 U2722 ( .A(n5043), .B(n11430), .Y(mem_wdata_D[54]) );
  CLKAND2X12 U2723 ( .A(n5043), .B(n11439), .Y(mem_wdata_D[63]) );
  CLKAND2X12 U2724 ( .A(n5043), .B(n11433), .Y(mem_wdata_D[57]) );
  CLKAND2X12 U2725 ( .A(n5046), .B(net103817), .Y(mem_wdata_I[50]) );
  INVX6 U2726 ( .A(n5045), .Y(n5046) );
  CLKAND2X12 U2727 ( .A(n5048), .B(n11266), .Y(mem_wdata_I[48]) );
  INVX6 U2728 ( .A(n5045), .Y(n5048) );
  INVX3 U2729 ( .A(n12952), .Y(n3569) );
  INVX12 U2730 ( .A(n3569), .Y(mem_wdata_I[51]) );
  CLKAND2X4 U2731 ( .A(n5047), .B(n11268), .Y(n12952) );
  INVX12 U2732 ( .A(n1856), .Y(mem_addr_I[6]) );
  CLKAND2X12 U2733 ( .A(n5046), .B(n11340), .Y(mem_wdata_I[125]) );
  INVX12 U2734 ( .A(n1928), .Y(mem_addr_D[8]) );
  INVX12 U2735 ( .A(n1929), .Y(mem_addr_D[9]) );
  BUFX16 U2736 ( .A(n12967), .Y(DCACHE_addr[16]) );
  INVXL U2737 ( .A(n5362), .Y(n5345) );
  AO22X1 U2738 ( .A0(ICACHE_addr[25]), .A1(mem_read_I), .B0(mem_write_I), .B1(
        n11367), .Y(n12859) );
  AO22XL U2739 ( .A0(ICACHE_addr[18]), .A1(mem_read_I), .B0(mem_write_I), .B1(
        n11360), .Y(n12866) );
  AO22XL U2740 ( .A0(ICACHE_addr[21]), .A1(mem_read_I), .B0(mem_write_I), .B1(
        n11363), .Y(n12863) );
  BUFX20 U2741 ( .A(n11537), .Y(mem_write_I) );
  OAI211X2 U2742 ( .A0(net112214), .A1(n6820), .B0(n6819), .C0(n7027), .Y(
        n3576) );
  INVX4 U2743 ( .A(n3576), .Y(n6954) );
  INVX4 U2744 ( .A(n6817), .Y(n7027) );
  NAND2X6 U2745 ( .A(n4624), .B(n6694), .Y(n3577) );
  AND2X8 U2746 ( .A(n8652), .B(net108003), .Y(n8654) );
  NAND3X2 U2747 ( .A(n9845), .B(n3732), .C(n3731), .Y(\i_MIPS/N59 ) );
  CLKAND2X2 U2748 ( .A(net104173), .B(n11287), .Y(n4448) );
  AO21X2 U2749 ( .A0(n7689), .A1(n9432), .B0(n7688), .Y(n7692) );
  AOI222X4 U2750 ( .A0(n5541), .A1(n11438), .B0(mem_rdata_D[62]), .B1(n132), 
        .C0(n12983), .C1(n5539), .Y(n10602) );
  AOI222X4 U2751 ( .A0(n5541), .A1(n11426), .B0(mem_rdata_D[50]), .B1(n133), 
        .C0(n12995), .C1(n5539), .Y(n10644) );
  AOI222X4 U2752 ( .A0(n5541), .A1(n11416), .B0(mem_rdata_D[40]), .B1(n131), 
        .C0(n13005), .C1(n5539), .Y(n10657) );
  CLKMX2X8 U2753 ( .A(n10670), .B(n10671), .S0(n4410), .Y(n3826) );
  AOI222X4 U2754 ( .A0(n5541), .A1(n11409), .B0(mem_rdata_D[33]), .B1(n129), 
        .C0(n13012), .C1(n5539), .Y(n10671) );
  AOI222X4 U2755 ( .A0(n3800), .A1(n11402), .B0(mem_rdata_D[26]), .B1(n131), 
        .C0(n12987), .C1(n5537), .Y(n10205) );
  CLKAND2X2 U2756 ( .A(n3898), .B(n11281), .Y(n4433) );
  OAI221X4 U2757 ( .A0(n10484), .A1(n5560), .B0(n5558), .B1(n10485), .C0(
        n10483), .Y(\i_MIPS/PC/n47 ) );
  INVX4 U2758 ( .A(n3894), .Y(net144236) );
  AOI222X4 U2759 ( .A0(n3800), .A1(n11392), .B0(mem_rdata_D[16]), .B1(n130), 
        .C0(n12997), .C1(n5537), .Y(n10506) );
  AND4X4 U2760 ( .A(n7677), .B(n7678), .C(net107389), .D(n7679), .Y(n3581) );
  AOI222X4 U2761 ( .A0(n5541), .A1(n11431), .B0(mem_rdata_D[55]), .B1(n130), 
        .C0(n12990), .C1(n5539), .Y(n10696) );
  NOR2BX2 U2762 ( .AN(net104171), .B(n3808), .Y(n4428) );
  CLKBUFX12 U2763 ( .A(net117751), .Y(net117745) );
  OAI222X4 U2764 ( .A0(net135772), .A1(net107688), .B0(net107217), .B1(n8117), 
        .C0(net107689), .C1(n8480), .Y(n7319) );
  INVXL U2765 ( .A(n7314), .Y(n8119) );
  NAND3X2 U2766 ( .A(n8134), .B(n7314), .C(n7486), .Y(n6653) );
  CLKINVX1 U2767 ( .A(net140147), .Y(n3585) );
  INVX4 U2768 ( .A(n3585), .Y(n3586) );
  INVX3 U2769 ( .A(net114331), .Y(n3587) );
  INVX8 U2770 ( .A(n3587), .Y(n3588) );
  INVX3 U2771 ( .A(net114319), .Y(n3592) );
  INVX6 U2772 ( .A(n3592), .Y(n3593) );
  INVX6 U2773 ( .A(n3596), .Y(n3597) );
  INVX3 U2774 ( .A(net114319), .Y(n3598) );
  INVX6 U2775 ( .A(n3598), .Y(n3599) );
  INVX3 U2776 ( .A(net114325), .Y(n3604) );
  CLKINVX1 U2777 ( .A(net114341), .Y(net114319) );
  CLKINVX1 U2778 ( .A(net140147), .Y(net114325) );
  INVX20 U2779 ( .A(net143514), .Y(net143504) );
  BUFX8 U2780 ( .A(n9715), .Y(n3607) );
  AO22X1 U2781 ( .A0(mem_rdata_I[69]), .A1(n5942), .B0(n5569), .B1(n11286), 
        .Y(n9715) );
  INVX6 U2782 ( .A(n3608), .Y(n3609) );
  BUFX8 U2783 ( .A(n9693), .Y(n3610) );
  AO22X1 U2784 ( .A0(mem_rdata_I[93]), .A1(n5943), .B0(n5569), .B1(n11309), 
        .Y(n9693) );
  BUFX8 U2785 ( .A(n9757), .Y(n3611) );
  AO22X1 U2786 ( .A0(mem_rdata_I[80]), .A1(n5942), .B0(n5569), .B1(n11297), 
        .Y(n9757) );
  INVX16 U2787 ( .A(n3638), .Y(net134673) );
  INVX16 U2788 ( .A(net134673), .Y(net117757) );
  NAND2X2 U2789 ( .A(\i_MIPS/ALUin1[25] ), .B(n6824), .Y(n7431) );
  BUFX8 U2790 ( .A(n11080), .Y(n3614) );
  AO22X1 U2791 ( .A0(mem_rdata_I[83]), .A1(n5939), .B0(n5569), .B1(n11299), 
        .Y(n11080) );
  OAI2BB2XL U2792 ( .B0(\i_MIPS/n161 ), .B1(net115793), .A0N(n10152), .A1N(
        n4544), .Y(\i_MIPS/N25 ) );
  BUFX8 U2793 ( .A(n9771), .Y(n3615) );
  AO22X1 U2794 ( .A0(mem_rdata_I[82]), .A1(n5942), .B0(n5569), .B1(net103785), 
        .Y(n9771) );
  OAI31X2 U2795 ( .A0(n8310), .A1(n8309), .A2(net107210), .B0(n8308), .Y(n3616) );
  NOR4X6 U2796 ( .A(n8307), .B(n8304), .C(n8305), .D(n8306), .Y(n8308) );
  CLKINVX3 U2797 ( .A(n8976), .Y(n3617) );
  NAND4BX2 U2798 ( .AN(n9372), .B(n9371), .C(n9370), .D(n9369), .Y(n9383) );
  BUFX8 U2799 ( .A(n10949), .Y(n3618) );
  AO22X1 U2800 ( .A0(mem_rdata_I[67]), .A1(n5942), .B0(n5569), .B1(n11284), 
        .Y(n10949) );
  XOR2X2 U2801 ( .A(n6609), .B(n6634), .Y(n6636) );
  INVX6 U2802 ( .A(n10334), .Y(n6609) );
  BUFX8 U2803 ( .A(n10920), .Y(n3619) );
  AO22X1 U2804 ( .A0(mem_rdata_I[66]), .A1(n5939), .B0(n5569), .B1(n11283), 
        .Y(n10920) );
  OAI221X1 U2805 ( .A0(n8863), .A1(n8862), .B0(n3673), .B1(n9295), .C0(n8861), 
        .Y(n3620) );
  NAND4BX2 U2806 ( .AN(n9381), .B(n9380), .C(n9379), .D(n9378), .Y(n9382) );
  OR2X1 U2807 ( .A(n8699), .B(n7422), .Y(n4494) );
  NOR2X1 U2808 ( .A(n8719), .B(n8720), .Y(n3623) );
  NAND2X2 U2809 ( .A(n4751), .B(n4752), .Y(n8720) );
  INVXL U2810 ( .A(net107141), .Y(net107606) );
  NAND2X8 U2811 ( .A(net117623), .B(net107141), .Y(net107138) );
  INVX1 U2812 ( .A(n7493), .Y(n3624) );
  OAI221X2 U2813 ( .A0(net107210), .A1(n3656), .B0(n9044), .B1(net107411), 
        .C0(net117759), .Y(n9047) );
  INVX1 U2814 ( .A(n9304), .Y(n9044) );
  OAI31X2 U2815 ( .A0(n7060), .A1(n7059), .A2(n7058), .B0(n7057), .Y(n3625) );
  NOR2X8 U2816 ( .A(n3912), .B(n7053), .Y(n7057) );
  INVXL U2817 ( .A(net109840), .Y(n3626) );
  OR2X1 U2818 ( .A(n9051), .B(\i_MIPS/ID_EX[81] ), .Y(n3627) );
  AND3X8 U2819 ( .A(n9216), .B(n8782), .C(net108623), .Y(n3628) );
  NAND2X4 U2820 ( .A(n6718), .B(n2921), .Y(n9216) );
  NAND2X4 U2821 ( .A(n3851), .B(n3974), .Y(net110932) );
  OR4X6 U2822 ( .A(net112393), .B(n6674), .C(n8634), .D(n6673), .Y(n3638) );
  OAI211XL U2823 ( .A0(n8471), .A1(n8467), .B0(n8199), .C0(n8464), .Y(n3629)
         );
  NAND4BX2 U2824 ( .AN(n9281), .B(n9280), .C(n9279), .D(n9278), .Y(n9292) );
  AND2X2 U2825 ( .A(net109965), .B(n8963), .Y(n4707) );
  CLKINVX12 U2826 ( .A(net107988), .Y(net109965) );
  AO22X2 U2827 ( .A0(net118237), .A1(n556), .B0(net118255), .B1(n2175), .Y(
        n8913) );
  AO22XL U2828 ( .A0(net118237), .A1(n727), .B0(net118255), .B1(n2532), .Y(
        n8802) );
  AO22XL U2829 ( .A0(net118237), .A1(n728), .B0(net118255), .B1(n2533), .Y(
        n8811) );
  BUFX4 U2830 ( .A(net118261), .Y(net118255) );
  INVXL U2831 ( .A(n4335), .Y(n3630) );
  AO22X1 U2832 ( .A0(net115799), .A1(n9824), .B0(n3584), .B1(n3586), .Y(
        \i_MIPS/n400 ) );
  CLKMX2X2 U2833 ( .A(\i_MIPS/n206 ), .B(n4779), .S0(n3894), .Y(n6720) );
  NAND2X2 U2834 ( .A(net134414), .B(n3894), .Y(n4396) );
  NAND2X4 U2835 ( .A(n3873), .B(net143514), .Y(n3786) );
  NAND3X6 U2836 ( .A(n7501), .B(n7504), .C(n2981), .Y(net105121) );
  OA22XL U2837 ( .A0(n8553), .A1(n8878), .B0(n9316), .B1(n7481), .Y(n7503) );
  CLKBUFX2 U2838 ( .A(n4729), .Y(n3632) );
  NAND2X2 U2839 ( .A(n7028), .B(n3983), .Y(n3636) );
  NAND3BX4 U2840 ( .AN(n7434), .B(net117745), .C(n11103), .Y(n7404) );
  INVX3 U2841 ( .A(n4090), .Y(net105112) );
  NOR2BX2 U2842 ( .AN(net104171), .B(n3806), .Y(n4425) );
  MX2XL U2843 ( .A(n3552), .B(net105506), .S0(n3588), .Y(\i_MIPS/n329 ) );
  OR4X6 U2844 ( .A(n6734), .B(n6733), .C(n6732), .D(n6731), .Y(net105313) );
  BUFX2 U2845 ( .A(n5450), .Y(n5441) );
  INVX8 U2846 ( .A(net112417), .Y(net108150) );
  NOR2X4 U2847 ( .A(n6704), .B(\i_MIPS/ALUin1[8] ), .Y(n4740) );
  INVX8 U2848 ( .A(n6704), .Y(n8115) );
  AOI2BB1X1 U2849 ( .A0N(\i_MIPS/PC/n21 ), .A1N(net115799), .B0(n10302), .Y(
        n10303) );
  AO22X1 U2850 ( .A0(n5555), .A1(n10978), .B0(n11054), .B1(n248), .Y(n10302)
         );
  OAI211X2 U2851 ( .A0(n8553), .A1(n9210), .B0(n8552), .C0(net107389), .Y(
        n8564) );
  INVX1 U2852 ( .A(n8467), .Y(n7479) );
  AND4X8 U2853 ( .A(n3628), .B(n7100), .C(n4700), .D(n8882), .Y(n3951) );
  INVX2 U2854 ( .A(n3577), .Y(net109511) );
  NAND2X2 U2855 ( .A(n8115), .B(\i_MIPS/ALUin1[8] ), .Y(n8124) );
  INVXL U2856 ( .A(net109674), .Y(n3639) );
  AND2X2 U2857 ( .A(n8129), .B(net118584), .Y(n3640) );
  AND2X4 U2858 ( .A(n8128), .B(n8127), .Y(n3641) );
  AND2X6 U2859 ( .A(n8126), .B(n8125), .Y(n3642) );
  NOR3X4 U2860 ( .A(n3640), .B(n3641), .C(n3642), .Y(n8139) );
  OR2X4 U2861 ( .A(net109040), .B(net117709), .Y(n3643) );
  OR2X4 U2862 ( .A(n3702), .B(net117731), .Y(n3644) );
  OAI31X1 U2863 ( .A0(n8470), .A1(n8469), .A2(n8468), .B0(n8467), .Y(n3645) );
  CLKMX2X2 U2864 ( .A(n8549), .B(n8548), .S0(net114079), .Y(net109040) );
  CLKINVX6 U2865 ( .A(n4883), .Y(n8470) );
  NAND2X4 U2866 ( .A(net108004), .B(net112417), .Y(net108149) );
  NOR3X6 U2867 ( .A(n3699), .B(n3700), .C(n3701), .Y(n9057) );
  INVX8 U2868 ( .A(net139838), .Y(net107411) );
  OAI221X2 U2869 ( .A0(net107210), .A1(n9124), .B0(net108148), .B1(n3774), 
        .C0(net117759), .Y(n7148) );
  MX2XL U2870 ( .A(DCACHE_addr[7]), .B(n3626), .S0(n3603), .Y(\i_MIPS/n390 )
         );
  INVX1 U2871 ( .A(n9298), .Y(n8659) );
  AO21X4 U2872 ( .A0(n9124), .A1(n9123), .B0(n9122), .Y(n9125) );
  BUFX4 U2873 ( .A(net117647), .Y(net117639) );
  BUFX4 U2874 ( .A(net139719), .Y(net117647) );
  OAI222X1 U2875 ( .A0(net107659), .A1(n9318), .B0(net107661), .B1(n9317), 
        .C0(n9316), .C1(n3620), .Y(n9321) );
  INVX2 U2876 ( .A(n9318), .Y(n8970) );
  CLKINVX1 U2877 ( .A(net108010), .Y(net108846) );
  INVX6 U2878 ( .A(n9549), .Y(n6675) );
  OR2X4 U2879 ( .A(n4687), .B(n8285), .Y(n3646) );
  OR2X4 U2880 ( .A(n8285), .B(n8394), .Y(n3647) );
  NAND4X2 U2881 ( .A(n4687), .B(n8286), .C(net117745), .D(n8394), .Y(n8284) );
  OAI2BB1X2 U2882 ( .A0N(net104963), .A1N(net104962), .B0(n3989), .Y(net108895) );
  NAND2X4 U2883 ( .A(n7102), .B(net108631), .Y(n9206) );
  INVXL U2884 ( .A(n9597), .Y(n3649) );
  XNOR2X4 U2885 ( .A(net105283), .B(n3650), .Y(n4055) );
  NAND2X6 U2886 ( .A(n3015), .B(net105269), .Y(n3650) );
  BUFX20 U2887 ( .A(net107607), .Y(net118225) );
  INVX20 U2888 ( .A(net117631), .Y(net117623) );
  NAND3X6 U2889 ( .A(n6391), .B(n5052), .C(n4625), .Y(n3651) );
  OA22X2 U2890 ( .A0(net107210), .A1(n3896), .B0(n3774), .B1(net108297), .Y(
        n8978) );
  NAND2X2 U2891 ( .A(n9299), .B(net107680), .Y(n8656) );
  NAND2X2 U2892 ( .A(\i_MIPS/ALUin1[5] ), .B(n7222), .Y(n9299) );
  OAI32X2 U2893 ( .A0(n8656), .A1(n8655), .A2(n8654), .B0(n8653), .B1(n9303), 
        .Y(n8658) );
  CLKINVX1 U2894 ( .A(n9299), .Y(n8653) );
  AOI211X4 U2895 ( .A0(net111249), .A1(net107652), .B0(n7316), .C0(n7315), .Y(
        n7317) );
  OAI222X2 U2896 ( .A0(n9137), .A1(n9318), .B0(net107661), .B1(n7313), .C0(
        n9316), .C1(n7312), .Y(n7316) );
  NAND3X8 U2897 ( .A(n3562), .B(n5053), .C(n5055), .Y(n3652) );
  OA22X4 U2898 ( .A0(n10404), .A1(n3766), .B0(n10407), .B1(n9536), .Y(n8438)
         );
  AND4X6 U2899 ( .A(n3815), .B(n3816), .C(n3818), .D(n3817), .Y(n4315) );
  OA22X2 U2900 ( .A0(n10674), .A1(n3766), .B0(n10677), .B1(n9536), .Y(n7358)
         );
  NAND3BX4 U2901 ( .AN(n4625), .B(n6391), .C(n5052), .Y(n9801) );
  BUFX16 U2902 ( .A(n9801), .Y(n5197) );
  CLKINVX8 U2903 ( .A(n5026), .Y(n4637) );
  ACHCINX4 U2904 ( .CIN(n4808), .A(\i_MIPS/IF_ID[26] ), .B(n6016), .CO(n10384)
         );
  AND2X2 U2905 ( .A(n3663), .B(n11280), .Y(n4471) );
  NOR2BX4 U2906 ( .AN(net104171), .B(n3798), .Y(n4473) );
  NOR2BX4 U2907 ( .AN(n3898), .B(n3805), .Y(n4474) );
  NAND3X4 U2908 ( .A(n3654), .B(n3655), .C(n10096), .Y(\i_MIPS/N60 ) );
  CLKBUFX2 U2909 ( .A(n9301), .Y(n3656) );
  INVX8 U2910 ( .A(\i_MIPS/n498 ), .Y(n11053) );
  AND2X1 U2911 ( .A(n3898), .B(n11299), .Y(n3842) );
  AND2XL U2912 ( .A(n9945), .B(n9946), .Y(n3657) );
  INVX12 U2913 ( .A(n9950), .Y(n9945) );
  AND2X2 U2914 ( .A(DCACHE_addr[0]), .B(n1319), .Y(n4725) );
  INVX20 U2915 ( .A(n3921), .Y(net104172) );
  CLKAND2X2 U2916 ( .A(n3898), .B(n11310), .Y(n4469) );
  NOR3BX2 U2917 ( .AN(n3659), .B(n4478), .C(n4479), .Y(n9726) );
  NAND2X2 U2918 ( .A(net104171), .B(n11224), .Y(n3659) );
  AND3X6 U2919 ( .A(net104830), .B(n10713), .C(net106822), .Y(n3660) );
  CLKAND2X2 U2920 ( .A(net104172), .B(n11264), .Y(n4438) );
  AOI222X2 U2921 ( .A0(net104171), .A1(n11242), .B0(net104172), .B1(n11273), 
        .C0(n3898), .C1(n11304), .Y(n10844) );
  NOR3BX2 U2922 ( .AN(n3662), .B(n4481), .C(n4480), .Y(n10132) );
  AOI222X2 U2923 ( .A0(n3827), .A1(n11221), .B0(n3663), .B1(n11252), .C0(n3898), .C1(n11283), .Y(n10931) );
  BUFX4 U2924 ( .A(n10767), .Y(n4502) );
  MXI2X2 U2925 ( .A(n10506), .B(n10505), .S0(n5545), .Y(n10507) );
  OAI221X1 U2926 ( .A0(n11061), .A1(n5560), .B0(n11060), .B1(n5557), .C0(
        n11058), .Y(\i_MIPS/PC/n59 ) );
  AND2X4 U2927 ( .A(ICACHE_addr[4]), .B(ICACHE_addr[3]), .Y(n4800) );
  NAND2X4 U2928 ( .A(net104830), .B(net106822), .Y(n10717) );
  OA22X4 U2929 ( .A0(n5744), .A1(n2061), .B0(n5694), .B1(n436), .Y(n11148) );
  CLKBUFX6 U2930 ( .A(n5707), .Y(n5694) );
  INVX12 U2931 ( .A(n3922), .Y(net104173) );
  INVX20 U2932 ( .A(n3922), .Y(n3898) );
  CLKAND2X2 U2933 ( .A(n3898), .B(n11295), .Y(n4439) );
  BUFX12 U2934 ( .A(net107120), .Y(n3921) );
  AND2X2 U2935 ( .A(n3898), .B(n11291), .Y(n4457) );
  CLKAND2X2 U2936 ( .A(n3898), .B(n11284), .Y(n4466) );
  CLKAND2X2 U2937 ( .A(n3898), .B(n11300), .Y(n4486) );
  AND2X1 U2938 ( .A(n3898), .B(n11292), .Y(n4445) );
  NOR2BX2 U2939 ( .AN(n3898), .B(n3801), .Y(n4472) );
  NOR2X6 U2940 ( .A(n4445), .B(n3000), .Y(n10096) );
  AND2X1 U2941 ( .A(n5044), .B(n11511), .Y(n4409) );
  NOR3X4 U2942 ( .A(n4425), .B(n4426), .C(n4427), .Y(n10889) );
  NAND2X6 U2943 ( .A(n3691), .B(\i_MIPS/ALUin1[2] ), .Y(net108151) );
  AND2X8 U2944 ( .A(n3785), .B(n3786), .Y(n3691) );
  OAI221X2 U2945 ( .A0(n9747), .A1(net143858), .B0(\i_MIPS/n504 ), .B1(
        net115789), .C0(n9746), .Y(\i_MIPS/N66 ) );
  CLKAND2X2 U2946 ( .A(net104172), .B(n11258), .Y(n4441) );
  INVX8 U2947 ( .A(n10604), .Y(n9487) );
  NAND4X8 U2948 ( .A(n7697), .B(n7700), .C(n7698), .D(n7699), .Y(net105425) );
  OAI211X4 U2949 ( .A0(n7691), .A1(n3749), .B0(net117745), .C0(n7690), .Y(
        n7699) );
  NAND4X2 U2950 ( .A(n7693), .B(n8635), .C(net117745), .D(n7692), .Y(n7698) );
  AOI21X2 U2951 ( .A0(net105423), .A1(net105424), .B0(net117723), .Y(net119021) );
  CLKINVX20 U2952 ( .A(net143857), .Y(net143858) );
  OA21X4 U2953 ( .A0(net106828), .A1(net104828), .B0(n9605), .Y(n3664) );
  NAND2X8 U2954 ( .A(n3664), .B(net135522), .Y(net107123) );
  CLKINVX20 U2955 ( .A(net107123), .Y(net104171) );
  AO21X2 U2956 ( .A0(n8882), .A1(n8881), .B0(n8880), .Y(n8887) );
  BUFX20 U2957 ( .A(n5408), .Y(n5401) );
  NAND2X2 U2958 ( .A(n2330), .B(n6963), .Y(n6961) );
  BUFX6 U2959 ( .A(net119018), .Y(n3947) );
  NAND3X6 U2960 ( .A(net143555), .B(net143556), .C(net109360), .Y(net105506)
         );
  CLKBUFX2 U2961 ( .A(net108874), .Y(n3666) );
  MX2X1 U2962 ( .A(DCACHE_addr[18]), .B(net105336), .S0(n3588), .Y(
        \i_MIPS/n379 ) );
  OAI21X2 U2963 ( .A0(n2950), .A1(n3855), .B0(n5193), .Y(n3667) );
  OAI21X2 U2964 ( .A0(n2950), .A1(n3855), .B0(n5193), .Y(net104963) );
  OAI22X4 U2965 ( .A0(n10640), .A1(n3877), .B0(n10643), .B1(n4495), .Y(n3855)
         );
  INVX16 U2966 ( .A(n3770), .Y(n3777) );
  INVX16 U2967 ( .A(n9547), .Y(n8976) );
  OAI2BB1X4 U2968 ( .A0N(n8027), .A1N(n8044), .B0(n8029), .Y(n7495) );
  NAND2X2 U2969 ( .A(\i_MIPS/ALUin1[9] ), .B(n3583), .Y(n8029) );
  NAND3BX2 U2970 ( .AN(n4625), .B(n5052), .C(n5055), .Y(n9808) );
  INVXL U2971 ( .A(n3606), .Y(n3668) );
  CLKINVX1 U2972 ( .A(n3668), .Y(n3669) );
  NAND2X4 U2973 ( .A(net104754), .B(net104755), .Y(n4322) );
  INVX4 U2974 ( .A(net108101), .Y(net104754) );
  INVX12 U2975 ( .A(n6669), .Y(n8634) );
  OA22X2 U2976 ( .A0(n10198), .A1(n3766), .B0(n10201), .B1(n9536), .Y(n7457)
         );
  OA22X2 U2977 ( .A0(n10738), .A1(n3766), .B0(n10741), .B1(n9536), .Y(n8758)
         );
  OA22X1 U2978 ( .A0(n10771), .A1(n3766), .B0(n10774), .B1(n9536), .Y(n7542)
         );
  OA22X2 U2979 ( .A0(n9799), .A1(n3767), .B0(n10759), .B1(n9536), .Y(n9181) );
  NAND2X4 U2980 ( .A(n4789), .B(n4721), .Y(n7889) );
  NAND2X4 U2981 ( .A(n4789), .B(n4784), .Y(n7891) );
  NAND2X4 U2982 ( .A(n4789), .B(n4787), .Y(n7890) );
  NOR4X4 U2983 ( .A(n9102), .B(n9101), .C(n9100), .D(n9099), .Y(n9103) );
  INVX2 U2984 ( .A(n7495), .Y(n7496) );
  CLKINVX3 U2985 ( .A(n6917), .Y(n4638) );
  NAND2X2 U2986 ( .A(\i_MIPS/ALUin1[16] ), .B(n6717), .Y(n9222) );
  OAI33X2 U2987 ( .A0(n3774), .A1(n1939), .A2(n6730), .B0(n1939), .B1(
        net107210), .B2(n6848), .Y(n6731) );
  NAND2BX2 U2988 ( .AN(n3861), .B(n6949), .Y(n7686) );
  NOR2X8 U2989 ( .A(net143524), .B(net143525), .Y(net139765) );
  CLKINVX1 U2990 ( .A(n8646), .Y(n3671) );
  OAI2BB1X2 U2991 ( .A0N(net104985), .A1N(net119263), .B0(net117631), .Y(
        net105549) );
  OAI21X4 U2992 ( .A0(n11373), .A1(n4637), .B0(n3789), .Y(n9798) );
  AOI32X4 U2993 ( .A0(net117743), .A1(n6838), .A2(n7402), .B0(n6827), .B1(
        n6822), .Y(n6853) );
  NAND4X8 U2994 ( .A(n4689), .B(\i_MIPS/EX_MEM_1 ), .C(DCACHE_ren), .D(n3789), 
        .Y(n9534) );
  NAND2X6 U2995 ( .A(net139775), .B(net105820), .Y(n10659) );
  MX2XL U2996 ( .A(DCACHE_addr[8]), .B(net105121), .S0(n3603), .Y(
        \i_MIPS/n389 ) );
  INVXL U2997 ( .A(n9121), .Y(n3672) );
  INVX4 U2998 ( .A(n7862), .Y(n7841) );
  NAND2X6 U2999 ( .A(\i_MIPS/ALUin1[22] ), .B(n6685), .Y(n7862) );
  NAND2X2 U3000 ( .A(n4687), .B(n8394), .Y(n8396) );
  CLKBUFX2 U3001 ( .A(net108854), .Y(n3857) );
  INVXL U3002 ( .A(n3974), .Y(net111413) );
  NAND2X2 U3003 ( .A(n6692), .B(n1263), .Y(n8211) );
  INVX12 U3004 ( .A(n6692), .Y(n6690) );
  AO21X2 U3005 ( .A0(net106602), .A1(net106603), .B0(net117623), .Y(net104755)
         );
  INVX6 U3006 ( .A(n3673), .Y(n3674) );
  NAND2X6 U3007 ( .A(n6704), .B(n343), .Y(n8134) );
  NAND2X1 U3008 ( .A(n343), .B(n8115), .Y(n8646) );
  CLKINVX8 U3009 ( .A(net105266), .Y(net110954) );
  NAND2X4 U3010 ( .A(n3673), .B(\i_MIPS/ID_EX[81] ), .Y(net108781) );
  NAND2X4 U3011 ( .A(n3673), .B(n3903), .Y(n8863) );
  CLKINVX16 U3012 ( .A(n4882), .Y(n6673) );
  CLKBUFX20 U3013 ( .A(net135551), .Y(n3950) );
  AND3XL U3014 ( .A(n3992), .B(n3993), .C(n3994), .Y(n3675) );
  NAND4BX2 U3015 ( .AN(n9290), .B(n9289), .C(n9288), .D(n9287), .Y(n9291) );
  OA22XL U3016 ( .A0(\i_MIPS/Register/register[6][17] ), .A1(n4661), .B0(
        \i_MIPS/Register/register[14][17] ), .B1(n5079), .Y(n9273) );
  OA22XL U3017 ( .A0(\i_MIPS/Register/register[22][4] ), .A1(n4661), .B0(
        \i_MIPS/Register/register[30][4] ), .B1(n5079), .Y(n9107) );
  OA22XL U3018 ( .A0(\i_MIPS/Register/register[6][4] ), .A1(n5083), .B0(
        \i_MIPS/Register/register[14][4] ), .B1(n5079), .Y(n9098) );
  CLKAND2X8 U3019 ( .A(\i_MIPS/jump_addr[18] ), .B(\i_MIPS/n504 ), .Y(n4788)
         );
  AOI22X4 U3020 ( .A0(net118225), .A1(net110569), .B0(net118217), .B1(
        net105425), .Y(net139863) );
  CLKAND2X12 U3021 ( .A(n4374), .B(n4375), .Y(n4368) );
  OA21X4 U3022 ( .A0(net108150), .A1(net108151), .B0(net108010), .Y(net112413)
         );
  NAND2X4 U3023 ( .A(\i_MIPS/ALUin1[3] ), .B(n6714), .Y(net108010) );
  NOR4X4 U3024 ( .A(n9111), .B(n9110), .C(n9109), .D(n9108), .Y(n9112) );
  OAI2BB1X4 U3025 ( .A0N(n3628), .A1N(n9218), .B0(n3676), .Y(n8573) );
  NAND2BX4 U3026 ( .AN(n7765), .B(n4883), .Y(n3906) );
  NAND2X6 U3027 ( .A(n3708), .B(n4883), .Y(n7959) );
  MX2X1 U3028 ( .A(net107656), .B(net107657), .S0(net107828), .Y(n4305) );
  AO22X4 U3029 ( .A0(n7304), .A1(net117747), .B0(n3950), .B1(n7305), .Y(n7310)
         );
  INVX4 U3030 ( .A(net104503), .Y(net111277) );
  NAND2X6 U3031 ( .A(net106040), .B(net106041), .Y(n4358) );
  CLKINVX8 U3032 ( .A(net111364), .Y(net106040) );
  MXI2X1 U3033 ( .A(\i_MIPS/ID_EX[71] ), .B(\i_MIPS/ID_EX[103] ), .S0(n3894), 
        .Y(n9422) );
  INVX6 U3034 ( .A(n4274), .Y(net111716) );
  AOI2BB1X1 U3035 ( .A0N(net109511), .A1N(net109513), .B0(net111723), .Y(n4275) );
  NAND2X6 U3036 ( .A(n348), .B(n4723), .Y(net107169) );
  NOR4X2 U3037 ( .A(n8149), .B(n8148), .C(n8147), .D(n8146), .Y(n8160) );
  BUFX4 U3038 ( .A(net118297), .Y(net118289) );
  BUFX8 U3039 ( .A(net107621), .Y(net118297) );
  NOR2X1 U3040 ( .A(n6815), .B(n6814), .Y(n6728) );
  INVX6 U3041 ( .A(net104752), .Y(net107518) );
  NAND3X8 U3042 ( .A(n6387), .B(n6386), .C(n2999), .Y(n11590) );
  XOR2X2 U3043 ( .A(ICACHE_addr[23]), .B(n6365), .Y(n6389) );
  XOR2X1 U3044 ( .A(ICACHE_addr[27]), .B(n6369), .Y(n6388) );
  MXI2X4 U3045 ( .A(n6713), .B(n12), .S0(n3894), .Y(n3703) );
  NAND4X6 U3046 ( .A(n4352), .B(n4350), .C(n4353), .D(n4351), .Y(n4346) );
  XOR2X4 U3047 ( .A(n4363), .B(n3706), .Y(n4352) );
  NAND3X6 U3048 ( .A(n7435), .B(n7436), .C(n3028), .Y(net105266) );
  AO22X4 U3049 ( .A0(net111716), .A1(net117747), .B0(n3950), .B1(net108622), 
        .Y(n4306) );
  INVX6 U3050 ( .A(net104166), .Y(n4357) );
  NAND2X2 U3051 ( .A(n4697), .B(n4711), .Y(n7608) );
  AND3X8 U3052 ( .A(n6655), .B(n3678), .C(n3679), .Y(n7101) );
  NAND4XL U3053 ( .A(net117745), .B(n6960), .C(n9429), .D(n7597), .Y(n6956) );
  INVX12 U3054 ( .A(n6721), .Y(n8283) );
  AO22X4 U3055 ( .A0(n7945), .A1(n9314), .B0(net107652), .B1(n9295), .Y(n7946)
         );
  INVXL U3056 ( .A(n9295), .Y(n9297) );
  INVX2 U3057 ( .A(n11392), .Y(n10505) );
  BUFX8 U3058 ( .A(n5404), .Y(n5387) );
  XOR3X1 U3059 ( .A(\i_MIPS/jump_addr[29] ), .B(\i_MIPS/Sign_Extend[31] ), .C(
        n10583), .Y(n10572) );
  NAND2X1 U3060 ( .A(\i_MIPS/ID_EX[74] ), .B(\i_MIPS/ID_EX[78] ), .Y(n6647) );
  CLKAND2X3 U3061 ( .A(net104171), .B(n11219), .Y(n4431) );
  INVX6 U3062 ( .A(net118313), .Y(net118307) );
  OR2X8 U3063 ( .A(n9465), .B(n9464), .Y(n3869) );
  AO21X4 U3064 ( .A0(n4727), .A1(n7487), .B0(n6653), .Y(n3678) );
  AND3X4 U3065 ( .A(n8029), .B(n7489), .C(n8124), .Y(n3679) );
  OA22X2 U3066 ( .A0(n5653), .A1(n568), .B0(n5607), .B1(n2186), .Y(n11181) );
  OA22X2 U3067 ( .A0(n5919), .A1(n569), .B0(n5877), .B1(n2187), .Y(n11178) );
  OA22X1 U3068 ( .A0(n5750), .A1(n960), .B0(n5695), .B1(n2585), .Y(n11180) );
  INVX16 U3069 ( .A(n8465), .Y(n8471) );
  NOR2X1 U3070 ( .A(net107210), .B(n7602), .Y(n3680) );
  CLKINVX1 U3071 ( .A(n3680), .Y(n3681) );
  OA22X1 U3072 ( .A0(n5919), .A1(n961), .B0(n5877), .B1(n2586), .Y(n11168) );
  NOR3X4 U3073 ( .A(n4440), .B(n4441), .C(n4442), .Y(n9867) );
  AND3X2 U3074 ( .A(n7781), .B(n7780), .C(net117747), .Y(n7783) );
  AND3X1 U3075 ( .A(net117747), .B(n7961), .C(n7955), .Y(n7958) );
  OAI31X2 U3076 ( .A0(n7223), .A1(net111413), .A2(n8659), .B0(n9299), .Y(n7224) );
  NOR4X2 U3077 ( .A(n7985), .B(n7984), .C(n7983), .D(n7982), .Y(n7986) );
  NOR4X2 U3078 ( .A(n7976), .B(n7975), .C(n7974), .D(n7973), .Y(n7987) );
  XOR2X4 U3079 ( .A(n11356), .B(ICACHE_addr[14]), .Y(n11596) );
  OAI211X2 U3080 ( .A0(n6964), .A1(n6963), .B0(n6962), .C0(n6961), .Y(n3683)
         );
  OA22X2 U3081 ( .A0(n138), .A1(n570), .B0(n5694), .B1(n2188), .Y(n11143) );
  NAND3BX2 U3082 ( .AN(n10588), .B(n10587), .C(n10586), .Y(\i_MIPS/PC/n64 ) );
  NAND2X8 U3083 ( .A(net112418), .B(\i_MIPS/n299 ), .Y(net108004) );
  NAND2X6 U3084 ( .A(n3785), .B(n3786), .Y(net112418) );
  OA22X2 U3085 ( .A0(n5833), .A1(n571), .B0(n5787), .B1(n2189), .Y(n11189) );
  XNOR2X4 U3086 ( .A(ICACHE_addr[10]), .B(n11352), .Y(n11132) );
  NAND4X4 U3087 ( .A(n11126), .B(n11125), .C(n11124), .D(n11123), .Y(n11352)
         );
  CLKMX2X2 U3088 ( .A(net118597), .B(net118592), .S0(n8551), .Y(n8552) );
  AO22X1 U3089 ( .A0(n10575), .A1(n4545), .B0(net104801), .B1(n10574), .Y(
        \i_MIPS/N46 ) );
  NOR2BX4 U3090 ( .AN(n3898), .B(n3802), .Y(n4451) );
  OR2XL U3091 ( .A(net107217), .B(n8885), .Y(n3684) );
  OR2X4 U3092 ( .A(n8884), .B(net117757), .Y(n3685) );
  OR2X2 U3093 ( .A(n9202), .B(n9315), .Y(n3686) );
  NAND3X2 U3094 ( .A(n3684), .B(n3685), .C(n3686), .Y(n8871) );
  INVX4 U3095 ( .A(n3754), .Y(n6401) );
  OR2X8 U3096 ( .A(n8220), .B(n8219), .Y(n3687) );
  OA22X2 U3097 ( .A0(n5654), .A1(n572), .B0(n5608), .B1(n2190), .Y(n11196) );
  OAI2BB1X1 U3098 ( .A0N(n9302), .A1N(n9301), .B0(n9300), .Y(n9306) );
  INVX4 U3099 ( .A(n8718), .Y(n4629) );
  NAND4X6 U3100 ( .A(n11154), .B(n11153), .C(n11152), .D(n11151), .Y(n11349)
         );
  OA22X2 U3101 ( .A0(n137), .A1(n573), .B0(n5694), .B1(n2191), .Y(n11153) );
  CLKMX2X3 U3102 ( .A(n8918), .B(n8917), .S0(net114087), .Y(n8919) );
  AO22X1 U3103 ( .A0(net118237), .A1(n767), .B0(net118255), .B1(n2359), .Y(
        n8589) );
  AO22X1 U3104 ( .A0(net118237), .A1(n768), .B0(net118255), .B1(n2360), .Y(
        n8506) );
  AO22X1 U3105 ( .A0(net118237), .A1(n769), .B0(net118255), .B1(n2361), .Y(
        n8497) );
  AO22X2 U3106 ( .A0(net118237), .A1(n552), .B0(net118255), .B1(n2171), .Y(
        n8904) );
  XOR2X1 U3107 ( .A(\i_MIPS/ID_EX[112] ), .B(n254), .Y(
        \i_MIPS/Hazard_detection/n9 ) );
  XOR2X1 U3108 ( .A(n10848), .B(n254), .Y(n6760) );
  NAND3X1 U3109 ( .A(n8637), .B(net108876), .C(n124), .Y(n8638) );
  NAND2X4 U3110 ( .A(n8673), .B(n8692), .Y(n6815) );
  NAND2X4 U3111 ( .A(n6685), .B(n2949), .Y(n8673) );
  CLKINVX6 U3112 ( .A(n9566), .Y(n9567) );
  NAND2X8 U3113 ( .A(n8650), .B(n2928), .Y(net112417) );
  INVX12 U3114 ( .A(n6714), .Y(n8650) );
  NAND2X1 U3115 ( .A(n3583), .B(n2920), .Y(n8645) );
  NAND2X6 U3116 ( .A(n6697), .B(n2937), .Y(net108873) );
  INVX6 U3117 ( .A(n6634), .Y(n10847) );
  OAI221X4 U3118 ( .A0(n10327), .A1(n5561), .B0(n5558), .B1(n10328), .C0(
        n10326), .Y(\i_MIPS/PC/n54 ) );
  OAI221X4 U3119 ( .A0(n10297), .A1(n5561), .B0(n5558), .B1(n10298), .C0(
        n10296), .Y(\i_MIPS/PC/n52 ) );
  NAND2X6 U3120 ( .A(\i_MIPS/ALUin1[20] ), .B(n6723), .Y(n8370) );
  INVX8 U3121 ( .A(n8370), .Y(n8889) );
  NAND2X2 U3122 ( .A(n6723), .B(n2919), .Y(n8381) );
  CLKINVX1 U3123 ( .A(n4071), .Y(n3690) );
  INVX4 U3124 ( .A(net105179), .Y(net105753) );
  OA22X1 U3125 ( .A0(n5400), .A1(n962), .B0(n5430), .B1(n2587), .Y(n6743) );
  OA22XL U3126 ( .A0(n5400), .A1(n1246), .B0(n5430), .B1(n2866), .Y(n6739) );
  NAND2XL U3127 ( .A(n9121), .B(net108010), .Y(n9131) );
  NAND2X2 U3128 ( .A(net135551), .B(n8286), .Y(n8303) );
  INVX20 U3129 ( .A(n3998), .Y(net135551) );
  NAND2X1 U3130 ( .A(n4755), .B(\i_MIPS/n287 ), .Y(n8131) );
  INVX20 U3131 ( .A(net107977), .Y(net109168) );
  NOR2X1 U3132 ( .A(net111930), .B(net117713), .Y(n3692) );
  NOR2X4 U3133 ( .A(net111931), .B(net117731), .Y(n3693) );
  CLKINVX1 U3134 ( .A(net111932), .Y(n3694) );
  CLKINVX4 U3135 ( .A(net105077), .Y(net111931) );
  CLKMX2X2 U3136 ( .A(\i_MIPS/ID_EX[70] ), .B(net105071), .S0(n3590), .Y(
        \i_MIPS/n309 ) );
  NAND2X6 U3137 ( .A(net108642), .B(n3835), .Y(n3783) );
  INVX1 U3138 ( .A(n8782), .Y(n9220) );
  NAND2X2 U3139 ( .A(n6717), .B(n959), .Y(n8782) );
  AND3X8 U3140 ( .A(n4672), .B(\i_MIPS/n248 ), .C(\i_MIPS/ALU_Control/n18 ), 
        .Y(n4674) );
  NAND4BBX2 U3141 ( .AN(\i_MIPS/ID_EX[105] ), .BN(n3964), .C(n4672), .D(
        \i_MIPS/ID_EX[106] ), .Y(n4835) );
  NAND2X8 U3142 ( .A(net134876), .B(net134907), .Y(n3770) );
  CLKAND2X3 U3143 ( .A(net104172), .B(n11257), .Y(n4450) );
  NAND2X2 U3144 ( .A(\i_MIPS/n222 ), .B(net144187), .Y(n4639) );
  MX2X2 U3145 ( .A(n8419), .B(n8418), .S0(net114085), .Y(n8420) );
  NOR4X2 U3146 ( .A(n9334), .B(n9333), .C(n9332), .D(n9331), .Y(n9345) );
  CLKBUFX2 U3147 ( .A(net107617), .Y(net118263) );
  OAI221X2 U3148 ( .A0(n4311), .A1(net143858), .B0(\i_MIPS/n503 ), .B1(
        net115791), .C0(n4312), .Y(\i_MIPS/N67 ) );
  NAND3X2 U3149 ( .A(\i_MIPS/PC/n6 ), .B(ICACHE_addr[4]), .C(\i_MIPS/PC/n7 ), 
        .Y(n4677) );
  INVXL U3150 ( .A(n8471), .Y(n3697) );
  NAND2X8 U3151 ( .A(n7775), .B(n3744), .Y(n8465) );
  AND2X2 U3152 ( .A(net104171), .B(n11225), .Y(n4446) );
  CLKBUFX8 U3153 ( .A(n5301), .Y(n5295) );
  CLKINVX8 U3154 ( .A(n8383), .Y(n8384) );
  INVX8 U3155 ( .A(net112410), .Y(net112446) );
  NAND2X8 U3156 ( .A(net112446), .B(n3670), .Y(net108854) );
  AND2X1 U3157 ( .A(net135551), .B(n7593), .Y(n4711) );
  INVX4 U3158 ( .A(net104934), .Y(n4343) );
  CLKMX2X8 U3159 ( .A(\i_MIPS/n218 ), .B(n4774), .S0(n3894), .Y(n6693) );
  NAND2X2 U3160 ( .A(n8290), .B(net107992), .Y(n8296) );
  INVX12 U3161 ( .A(n7845), .Y(n7102) );
  CLKINVX6 U3162 ( .A(n8200), .Y(n8201) );
  NAND4BX2 U3163 ( .AN(n8776), .B(n8775), .C(n8774), .D(n8773), .Y(n8777) );
  NOR4X1 U3164 ( .A(n8772), .B(n8771), .C(n8770), .D(n8769), .Y(n8773) );
  OA22XL U3165 ( .A0(\i_MIPS/Register/register[22][0] ), .A1(n5083), .B0(
        \i_MIPS/Register/register[30][0] ), .B1(n5079), .Y(n8768) );
  MX2XL U3166 ( .A(DCACHE_addr[29]), .B(n3649), .S0(n3591), .Y(\i_MIPS/n368 )
         );
  OAI221X1 U3167 ( .A0(n10276), .A1(n5561), .B0(n5557), .B1(n10277), .C0(
        n10275), .Y(\i_MIPS/PC/n50 ) );
  OAI221X1 U3168 ( .A0(n5562), .A1(\i_MIPS/n154 ), .B0(n5557), .B1(
        \i_MIPS/PC/n3 ), .C0(n10660), .Y(\i_MIPS/PC/n35 ) );
  OAI2BB1X4 U3169 ( .A0N(n4705), .A1N(n8116), .B0(n7770), .Y(n8027) );
  NAND2X2 U3170 ( .A(n8124), .B(n7489), .Y(n7766) );
  BUFX2 U3171 ( .A(n11209), .Y(n5795) );
  OAI221X4 U3172 ( .A0(n10358), .A1(n5561), .B0(n5558), .B1(n10359), .C0(
        n10357), .Y(\i_MIPS/PC/n57 ) );
  AOI21X1 U3173 ( .A0(net108003), .A1(n3867), .B0(net108005), .Y(n4703) );
  CLKAND2X2 U3174 ( .A(n4707), .B(n9049), .Y(n3699) );
  AO22X2 U3175 ( .A0(n9044), .A1(net117747), .B0(n3950), .B1(n3656), .Y(n9046)
         );
  NAND2XL U3176 ( .A(n9300), .B(n9302), .Y(n9045) );
  AND4X8 U3177 ( .A(n8489), .B(n8491), .C(n8490), .D(n8488), .Y(n3702) );
  OA22X1 U3178 ( .A0(n5919), .A1(n964), .B0(n5877), .B1(n2589), .Y(n11183) );
  NAND2X6 U3179 ( .A(n5075), .B(\i_MIPS/ALUin1[25] ), .Y(n7587) );
  OA22XL U3180 ( .A0(\i_MIPS/ALUin1[24] ), .A1(n5064), .B0(\i_MIPS/ALUin1[25] ), .B1(n5059), .Y(n6831) );
  OA22XL U3181 ( .A0(\i_MIPS/ALUin1[25] ), .A1(n5063), .B0(\i_MIPS/ALUin1[26] ), .B1(n5057), .Y(n7410) );
  AND2X2 U3182 ( .A(net104171), .B(n11229), .Y(n4455) );
  OR4X8 U3183 ( .A(n7052), .B(n7049), .C(n7050), .D(n7051), .Y(n7053) );
  NAND4X2 U3184 ( .A(n7046), .B(n7045), .C(n7044), .D(n7043), .Y(n7050) );
  NAND2X6 U3185 ( .A(n4639), .B(n4640), .Y(n7775) );
  NAND2X8 U3186 ( .A(net112392), .B(net108787), .Y(n3998) );
  INVX8 U3187 ( .A(n7887), .Y(n9503) );
  INVX8 U3188 ( .A(n10769), .Y(n9119) );
  XOR2X4 U3189 ( .A(n4310), .B(n3996), .Y(n4319) );
  NAND4BX1 U3190 ( .AN(n9199), .B(n9198), .C(n9197), .D(n9196), .Y(net107858)
         );
  NOR4X4 U3191 ( .A(n9195), .B(n9194), .C(n9193), .D(n9192), .Y(n9196) );
  AO22X2 U3192 ( .A0(n6935), .A1(n3748), .B0(n6934), .B1(n9314), .Y(n6943) );
  INVXL U3193 ( .A(n9452), .Y(n6934) );
  BUFX12 U3194 ( .A(n3704), .Y(n5050) );
  AND2X8 U3195 ( .A(n5050), .B(n9544), .Y(n4754) );
  MX2X1 U3196 ( .A(n3545), .B(net104980), .S0(n3597), .Y(\i_MIPS/n333 ) );
  INVX3 U3197 ( .A(n3702), .Y(n3971) );
  OA22X2 U3198 ( .A0(\i_MIPS/Register/register[22][20] ), .A1(n5083), .B0(
        \i_MIPS/Register/register[30][20] ), .B1(n5079), .Y(n8448) );
  OAI221X2 U3199 ( .A0(n9552), .A1(n7313), .B0(n9202), .B1(n7312), .C0(
        net107389), .Y(n7051) );
  AND4X6 U3200 ( .A(n4332), .B(n4333), .C(n4331), .D(n4330), .Y(n3916) );
  INVXL U3201 ( .A(n9055), .Y(n8388) );
  NOR2X2 U3202 ( .A(n8372), .B(n8210), .Y(n3707) );
  BUFX20 U3203 ( .A(n12979), .Y(n5052) );
  OA22X4 U3204 ( .A0(n5260), .A1(n2063), .B0(n5302), .B1(n438), .Y(n6458) );
  XNOR2X4 U3205 ( .A(net106031), .B(n10910), .Y(n4321) );
  OAI2BB1X2 U3206 ( .A0N(net105110), .A1N(net105111), .B0(n3989), .Y(net110642) );
  NAND2X4 U3207 ( .A(n4546), .B(n183), .Y(n7041) );
  NAND2X2 U3208 ( .A(n6920), .B(n6919), .Y(n7430) );
  INVXL U3209 ( .A(n4357), .Y(n3709) );
  OA21X4 U3210 ( .A0(n4712), .A1(n7858), .B0(n6915), .Y(n3710) );
  AND2X8 U3211 ( .A(n6652), .B(n6916), .Y(n4712) );
  NAND2X8 U3212 ( .A(n4706), .B(n8381), .Y(n7858) );
  AND2X8 U3213 ( .A(n7856), .B(n8885), .Y(n4732) );
  INVXL U3214 ( .A(n6476), .Y(n11039) );
  OA22X4 U3215 ( .A0(n5307), .A1(n3711), .B0(n5259), .B1(n2058), .Y(n6468) );
  XNOR2X4 U3216 ( .A(n3712), .B(n4362), .Y(n4054) );
  NAND3X6 U3217 ( .A(n3813), .B(n3814), .C(net112330), .Y(n3712) );
  OAI221X4 U3218 ( .A0(n345), .A1(n5072), .B0(n2919), .B1(n5068), .C0(n7154), 
        .Y(n3713) );
  OAI221X2 U3219 ( .A0(n345), .A1(n5072), .B0(n2919), .B1(n5068), .C0(n7154), 
        .Y(n7478) );
  OAI211X2 U3220 ( .A0(n4750), .A1(net110928), .B0(n8666), .C0(n7492), .Y(
        n8477) );
  AOI32X2 U3221 ( .A0(n4693), .A1(n3665), .A2(n8396), .B0(n8682), .B1(n4698), 
        .Y(n8398) );
  OR2X1 U3222 ( .A(n2961), .B(n5072), .Y(n3716) );
  OR2X1 U3223 ( .A(n5067), .B(n347), .Y(n3717) );
  INVX20 U3224 ( .A(n5074), .Y(n5072) );
  CLKAND2X2 U3225 ( .A(net104171), .B(n11249), .Y(n4470) );
  NAND2X2 U3226 ( .A(\i_MIPS/ALUin1[18] ), .B(n6700), .Y(n8556) );
  XOR2X4 U3227 ( .A(n6439), .B(n1329), .Y(n3925) );
  AOI2BB2X4 U3228 ( .B0(net118217), .B1(net104752), .A0N(n3890), .A1N(n3719), 
        .Y(net139776) );
  AND4X6 U3229 ( .A(n4338), .B(n4340), .C(n4337), .D(n4339), .Y(n3915) );
  NAND2X2 U3230 ( .A(n8293), .B(\i_MIPS/ID_EX[81] ), .Y(n4377) );
  BUFX20 U3231 ( .A(n5353), .Y(n5355) );
  OA22X2 U3232 ( .A0(n5331), .A1(n575), .B0(n5356), .B1(n2193), .Y(n8822) );
  OA22X1 U3233 ( .A0(n5175), .A1(n965), .B0(n5214), .B1(n2590), .Y(n8824) );
  CLKAND2X3 U3234 ( .A(net104171), .B(n11230), .Y(n4443) );
  OAI221X2 U3235 ( .A0(n5169), .A1(n1938), .B0(n5209), .B1(n353), .C0(n6399), 
        .Y(n3720) );
  XOR2X4 U3236 ( .A(n4671), .B(DCACHE_addr[20]), .Y(n6457) );
  NAND3BX4 U3237 ( .AN(net108787), .B(n3726), .C(n4741), .Y(net107218) );
  MX2X1 U3238 ( .A(net107657), .B(net107656), .S0(n7956), .Y(n7957) );
  XOR2X4 U3239 ( .A(n3723), .B(DCACHE_addr[26]), .Y(n6503) );
  NAND2X6 U3240 ( .A(n3931), .B(n11005), .Y(n3723) );
  NOR4X4 U3241 ( .A(n6637), .B(n6636), .C(\i_MIPS/n302 ), .D(n6756), .Y(n6638)
         );
  OAI221X2 U3242 ( .A0(net107210), .A1(n8123), .B0(n4702), .B1(n3774), .C0(
        net117759), .Y(n8127) );
  NAND2X6 U3243 ( .A(net139776), .B(net106301), .Y(n10910) );
  INVX2 U3244 ( .A(n8962), .Y(n8964) );
  INVX4 U3245 ( .A(net109196), .Y(net109496) );
  BUFX20 U3246 ( .A(n9537), .Y(n3767) );
  OA22X2 U3247 ( .A0(n9804), .A1(n3767), .B0(n10750), .B1(n9536), .Y(n9097) );
  NAND2XL U3248 ( .A(n11021), .B(n11020), .Y(n11531) );
  NAND2X8 U3249 ( .A(n11021), .B(n11020), .Y(n3725) );
  INVX8 U3250 ( .A(n6507), .Y(n11020) );
  AOI2BB2X4 U3251 ( .B0(n3755), .B1(\D_cache/cache[7][140] ), .A0N(n5407), 
        .A1N(n3724), .Y(n6411) );
  BUFX16 U3252 ( .A(n5339), .Y(n5363) );
  NAND4X4 U3253 ( .A(n8424), .B(n8423), .C(n8422), .D(n8421), .Y(n11492) );
  NAND4X4 U3254 ( .A(n7264), .B(n7263), .C(n7262), .D(n7261), .Y(n11478) );
  INVX6 U3255 ( .A(n6410), .Y(n10982) );
  CLKMX2X2 U3256 ( .A(n8962), .B(n9314), .S0(\i_MIPS/ID_EX[81] ), .Y(n6843) );
  BUFX4 U3257 ( .A(n5116), .Y(n5114) );
  OAI221X2 U3258 ( .A0(n2949), .A1(n5072), .B0(n345), .B1(n5068), .C0(n7105), 
        .Y(net109196) );
  BUFX16 U3259 ( .A(n5448), .Y(n5447) );
  OAI221X2 U3260 ( .A0(net107210), .A1(n7305), .B0(n7304), .B1(n3774), .C0(
        net117757), .Y(n7307) );
  NAND2X4 U3261 ( .A(n4788), .B(n4721), .Y(n7885) );
  NOR4X4 U3262 ( .A(n9186), .B(n9185), .C(n9184), .D(n9183), .Y(n9187) );
  XOR2X4 U3263 ( .A(n3725), .B(n12956), .Y(n6513) );
  AND2X8 U3264 ( .A(net139866), .B(net105567), .Y(n4364) );
  INVX2 U3265 ( .A(n9224), .Y(n8781) );
  MX2XL U3266 ( .A(n5053), .B(net104752), .S0(n3591), .Y(\i_MIPS/n394 ) );
  AO22XL U3267 ( .A0(n5556), .A1(n10526), .B0(n11054), .B1(n10334), .Y(n10335)
         );
  NAND2XL U3268 ( .A(n11003), .B(n11002), .Y(n11528) );
  BUFX12 U3269 ( .A(n5354), .Y(n5362) );
  INVX4 U3270 ( .A(n6673), .Y(n3726) );
  BUFX12 U3271 ( .A(n8698), .Y(n4882) );
  CLKAND2X2 U3272 ( .A(net104171), .B(n11247), .Y(n4458) );
  INVX8 U3273 ( .A(n5026), .Y(n4407) );
  CLKBUFX4 U3274 ( .A(n5353), .Y(n5351) );
  INVX3 U3275 ( .A(n10512), .Y(n8959) );
  XNOR2X4 U3276 ( .A(net105137), .B(n4327), .Y(n4325) );
  AND4X6 U3277 ( .A(n4319), .B(n4321), .C(n4318), .D(n4320), .Y(n3918) );
  NOR2BX2 U3278 ( .AN(net104172), .B(n3728), .Y(n4459) );
  OA22X1 U3279 ( .A0(net107217), .A1(n6918), .B0(n1939), .B1(net117759), .Y(
        n6682) );
  OAI221X1 U3280 ( .A0(n3897), .A1(net107210), .B0(net108308), .B1(n3774), 
        .C0(net117759), .Y(n3829) );
  AND3X4 U3281 ( .A(\i_MIPS/PC/n7 ), .B(ICACHE_addr[2]), .C(\i_MIPS/PC/n8 ), 
        .Y(n4836) );
  OA22X4 U3282 ( .A0(n5831), .A1(n2064), .B0(n5786), .B1(n439), .Y(n11142) );
  OR2X8 U3283 ( .A(net118601), .B(n3858), .Y(n3729) );
  OR2X4 U3284 ( .A(net108781), .B(n9049), .Y(n3730) );
  NAND4BX2 U3285 ( .AN(n9106), .B(n9105), .C(n9104), .D(n9103), .Y(n9117) );
  OR2X4 U3286 ( .A(n9846), .B(net143858), .Y(n3731) );
  OR2X2 U3287 ( .A(\i_MIPS/n511 ), .B(net115791), .Y(n3732) );
  NAND2X4 U3288 ( .A(n4801), .B(\i_MIPS/PC/n8 ), .Y(n4658) );
  INVX12 U3289 ( .A(n3821), .Y(n10188) );
  NAND2X6 U3290 ( .A(n11373), .B(n3789), .Y(n11504) );
  OA22X1 U3291 ( .A0(n5182), .A1(n1274), .B0(n5219), .B1(n2903), .Y(n6561) );
  OAI221X2 U3292 ( .A0(n10231), .A1(net143858), .B0(\i_MIPS/n508 ), .B1(
        net115793), .C0(n10230), .Y(\i_MIPS/N62 ) );
  NOR3X4 U3293 ( .A(n4431), .B(n4432), .C(n4433), .Y(n10823) );
  CLKAND2X2 U3294 ( .A(net104172), .B(n11250), .Y(n4432) );
  NAND4X6 U3295 ( .A(n4096), .B(n4095), .C(n4097), .D(n4098), .Y(n3791) );
  AOI2BB2X4 U3296 ( .B0(net118215), .B1(n10619), .A0N(n3890), .A1N(n3948), .Y(
        n3733) );
  INVX4 U3297 ( .A(n8205), .Y(n8206) );
  NAND3X4 U3298 ( .A(n4643), .B(n3628), .C(n2996), .Y(n4620) );
  INVXL U3299 ( .A(n9119), .Y(n3734) );
  OR2X2 U3300 ( .A(n9316), .B(n9052), .Y(n3735) );
  OR2X2 U3301 ( .A(net107987), .B(n9050), .Y(n3737) );
  OAI221X4 U3302 ( .A0(\i_MIPS/ALUin1[7] ), .A1(n5072), .B0(\i_MIPS/ALUin1[6] ), .B1(n5068), .C0(n8679), .Y(n9051) );
  CLKMX2X2 U3303 ( .A(n8204), .B(n8203), .S0(\i_MIPS/ID_EX[81] ), .Y(n9050) );
  NAND4X4 U3304 ( .A(n11171), .B(n11170), .C(n11169), .D(n11168), .Y(n11356)
         );
  NOR2BX2 U3305 ( .AN(net104173), .B(n3803), .Y(n4463) );
  NOR2BX2 U3306 ( .AN(n3898), .B(n3804), .Y(n4492) );
  CLKBUFX2 U3307 ( .A(n4658), .Y(n5706) );
  NAND2X6 U3308 ( .A(n11000), .B(n10999), .Y(n6418) );
  OA22X4 U3309 ( .A0(n5401), .A1(n2065), .B0(n5447), .B1(n440), .Y(n6416) );
  OR2X6 U3310 ( .A(n5211), .B(n2951), .Y(n3739) );
  OR2X4 U3311 ( .A(net107517), .B(net117709), .Y(n3740) );
  OR2X6 U3312 ( .A(net107518), .B(net117731), .Y(n3741) );
  CLKMX2X4 U3313 ( .A(n9383), .B(n9382), .S0(net114079), .Y(net107517) );
  OAI2BB1X4 U3314 ( .A0N(n10581), .A1N(n10578), .B0(n10579), .Y(n10722) );
  MXI2X4 U3315 ( .A(n10662), .B(n10661), .S0(n5548), .Y(n10663) );
  NOR3X2 U3316 ( .A(n4383), .B(n4384), .C(n4385), .Y(n10662) );
  AND4X8 U3317 ( .A(n4366), .B(n4367), .C(n4368), .D(n4369), .Y(n6446) );
  NOR2BX2 U3318 ( .AN(net104171), .B(n3812), .Y(n4434) );
  NAND4X4 U3319 ( .A(n8824), .B(n8823), .C(n8822), .D(n8821), .Y(n11456) );
  AND4X6 U3320 ( .A(n9214), .B(n9215), .C(n9213), .D(n9212), .Y(n3742) );
  NAND2X6 U3321 ( .A(n10987), .B(n10988), .Y(n6403) );
  MX2XL U3322 ( .A(n12957), .B(net105112), .S0(n3597), .Y(\i_MIPS/n371 ) );
  AND3X6 U3323 ( .A(n4725), .B(DCACHE_ren), .C(\i_MIPS/EX_MEM_1 ), .Y(n3743)
         );
  AND2X6 U3324 ( .A(n11374), .B(n3743), .Y(n4059) );
  NAND2X1 U3325 ( .A(n8300), .B(n8288), .Y(n8286) );
  INVX2 U3326 ( .A(n3022), .Y(n3850) );
  INVX3 U3327 ( .A(n11434), .Y(n10207) );
  OAI221X4 U3328 ( .A0(n2184), .A1(n5064), .B0(n344), .B1(n5056), .C0(n6662), 
        .Y(n3745) );
  INVX8 U3329 ( .A(n5061), .Y(n5056) );
  MXI2X4 U3330 ( .A(n3747), .B(n3746), .S0(net143514), .Y(n6715) );
  AOI22X4 U3331 ( .A0(n3856), .A1(\D_cache/cache[2][135] ), .B0(n3924), .B1(
        \D_cache/cache[3][135] ), .Y(n6440) );
  AND3X1 U3332 ( .A(net117743), .B(n7034), .C(n8673), .Y(n7056) );
  NOR2BX4 U3333 ( .AN(DCACHE_addr[16]), .B(n3720), .Y(n3787) );
  MX2XL U3334 ( .A(DCACHE_addr[15]), .B(n10619), .S0(n3595), .Y(\i_MIPS/n382 )
         );
  MX2X1 U3335 ( .A(net107656), .B(net107657), .S0(n8469), .Y(n7484) );
  AND2X8 U3336 ( .A(net134876), .B(\i_MIPS/ID_EX[83] ), .Y(n3748) );
  NAND3BX2 U3337 ( .AN(n9557), .B(n9566), .C(net117745), .Y(n9575) );
  NAND2X4 U3338 ( .A(\i_MIPS/ALUin1[21] ), .B(n6724), .Y(n8860) );
  AOI21X1 U3339 ( .A0(n7689), .A1(n9432), .B0(n7688), .Y(n3749) );
  OA22X2 U3340 ( .A0(n10777), .A1(n3878), .B0(n10780), .B1(n4495), .Y(n7541)
         );
  NOR4X4 U3341 ( .A(n8473), .B(n8474), .C(n8475), .D(n8472), .Y(n8491) );
  AOI2BB1X2 U3342 ( .A0N(n5059), .A1N(n347), .B0(n4798), .Y(n6663) );
  CLKAND2X8 U3343 ( .A(n5065), .B(\i_MIPS/ALUin1[29] ), .Y(n4798) );
  INVXL U3344 ( .A(n11012), .Y(n3750) );
  CLKINVX1 U3345 ( .A(n3750), .Y(n3751) );
  BUFX20 U3346 ( .A(n3652), .Y(n5406) );
  INVX20 U3347 ( .A(n5060), .Y(n5059) );
  OA22X4 U3348 ( .A0(\i_MIPS/n297 ), .A1(n5064), .B0(\i_MIPS/n296 ), .B1(n5059), .Y(n6834) );
  OA22X2 U3349 ( .A0(n3744), .A1(n5063), .B0(n1263), .B1(n5059), .Y(n6658) );
  AO22X4 U3350 ( .A0(n8868), .A1(n3748), .B0(n8867), .B1(n9295), .Y(n8869) );
  INVX8 U3351 ( .A(n11489), .Y(n10620) );
  NAND4X4 U3352 ( .A(n9258), .B(n9257), .C(n9256), .D(n9255), .Y(n11489) );
  OA22X1 U3353 ( .A0(n5333), .A1(n966), .B0(n5358), .B1(n2591), .Y(n9256) );
  CLKMX2X3 U3354 ( .A(n7648), .B(n7647), .S0(net114081), .Y(net110640) );
  NAND4BX2 U3355 ( .AN(n7646), .B(n7645), .C(n7644), .D(n7643), .Y(n7647) );
  NAND2X2 U3356 ( .A(n4788), .B(n4787), .Y(n7886) );
  NAND2X2 U3357 ( .A(n4788), .B(n4786), .Y(n7884) );
  CLKBUFX6 U3358 ( .A(n5311), .Y(n5294) );
  NAND2X8 U3359 ( .A(n4633), .B(n8571), .Y(net104964) );
  AOI33X4 U3360 ( .A0(n8570), .A1(n8569), .A2(net117743), .B0(n8568), .B1(
        n8567), .B2(net117743), .Y(n8571) );
  NAND2X4 U3361 ( .A(n8462), .B(net144224), .Y(n4376) );
  INVX20 U3362 ( .A(n149), .Y(n7486) );
  NAND2X8 U3363 ( .A(n11012), .B(n11011), .Y(n6435) );
  OAI2BB2X4 U3364 ( .B0(n5407), .B1(n3756), .A0N(n3755), .A1N(
        \D_cache/cache[7][139] ), .Y(n3754) );
  AO21X4 U3365 ( .A0(n8937), .A1(n8936), .B0(n5191), .Y(net105143) );
  AND2XL U3366 ( .A(\i_MIPS/EX_MEM[5] ), .B(n5190), .Y(n3757) );
  CLKMX2X8 U3367 ( .A(\i_MIPS/n182 ), .B(n4772), .S0(n3894), .Y(n9556) );
  MXI2X2 U3368 ( .A(\i_MIPS/ID_EX[68] ), .B(\i_MIPS/ID_EX[100] ), .S0(n3894), 
        .Y(n6951) );
  MXI2X2 U3369 ( .A(\i_MIPS/ID_EX[66] ), .B(\i_MIPS/ID_EX[98] ), .S0(n3894), 
        .Y(n6823) );
  MXI2X2 U3370 ( .A(\i_MIPS/ID_EX[65] ), .B(\i_MIPS/ID_EX[97] ), .S0(n3894), 
        .Y(n6667) );
  MXI2X2 U3371 ( .A(\i_MIPS/ID_EX[67] ), .B(\i_MIPS/ID_EX[99] ), .S0(n3894), 
        .Y(n6950) );
  MXI2X2 U3372 ( .A(\i_MIPS/ID_EX[64] ), .B(\i_MIPS/ID_EX[96] ), .S0(n3894), 
        .Y(n6726) );
  MX2X2 U3373 ( .A(\i_MIPS/n208 ), .B(n4777), .S0(n3894), .Y(n6719) );
  MXI2X2 U3374 ( .A(\i_MIPS/ID_EX[70] ), .B(\i_MIPS/ID_EX[102] ), .S0(n3894), 
        .Y(n6938) );
  MX2X8 U3375 ( .A(\i_MIPS/n220 ), .B(n4775), .S0(net143514), .Y(n6692) );
  OAI221X2 U3376 ( .A0(n10098), .A1(n3766), .B0(n10101), .B1(n5189), .C0(n7812), .Y(n7836) );
  AOI2BB2X2 U3377 ( .B0(n8203), .B1(n8291), .A0N(n8863), .A1N(n3745), .Y(n8702) );
  INVX3 U3378 ( .A(n8700), .Y(n8203) );
  NAND2X2 U3379 ( .A(\i_MIPS/ALUin1[29] ), .B(n6939), .Y(n9424) );
  AO22X2 U3380 ( .A0(n7225), .A1(net117747), .B0(n3950), .B1(n3909), .Y(n7227)
         );
  NAND2X6 U3381 ( .A(net105462), .B(net105463), .Y(n4327) );
  CLKINVX8 U3382 ( .A(net108412), .Y(net105462) );
  NAND2X2 U3383 ( .A(\i_MIPS/ALUin1[11] ), .B(n7775), .Y(net108851) );
  NAND2XL U3384 ( .A(n9219), .B(n8782), .Y(n8788) );
  NAND2X6 U3385 ( .A(\i_MIPS/ALUin1[16] ), .B(n6698), .Y(n9219) );
  AO21X4 U3386 ( .A0(net105255), .A1(net105256), .B0(net117625), .Y(net105582)
         );
  INVX8 U3387 ( .A(n7597), .Y(n7595) );
  NAND2X4 U3388 ( .A(\i_MIPS/ALUin1[14] ), .B(n6715), .Y(net108876) );
  NAND2X4 U3389 ( .A(n6675), .B(\i_MIPS/ALU/N303 ), .Y(n3758) );
  INVX3 U3390 ( .A(\i_MIPS/ID_EX[83] ), .Y(net108631) );
  NAND3X6 U3391 ( .A(n3990), .B(n3991), .C(net108162), .Y(net104906) );
  INVXL U3392 ( .A(net107855), .Y(n3759) );
  NAND2XL U3393 ( .A(n10982), .B(n10981), .Y(n11521) );
  CLKAND2X12 U3394 ( .A(n4400), .B(n4399), .Y(n3926) );
  INVX1 U3395 ( .A(n8481), .Y(n8478) );
  OAI21X4 U3396 ( .A0(n11582), .A1(n11581), .B0(n11580), .Y(n11583) );
  NAND3BX4 U3397 ( .AN(n9431), .B(n4728), .C(n11112), .Y(n11582) );
  NAND2X4 U3398 ( .A(n9443), .B(\i_MIPS/n271 ), .Y(n11105) );
  NAND2X2 U3399 ( .A(n10984), .B(n3782), .Y(n4375) );
  INVXL U3400 ( .A(net109359), .Y(n3761) );
  OAI31X2 U3401 ( .A0(n8310), .A1(n8309), .A2(net107210), .B0(n8308), .Y(
        net104343) );
  CLKMX2X12 U3402 ( .A(net107656), .B(net107657), .S0(n8864), .Y(n8870) );
  NAND3BX1 U3403 ( .AN(n9225), .B(n9227), .C(net117745), .Y(n9233) );
  NAND2XL U3404 ( .A(net139862), .B(net105756), .Y(n10473) );
  OA22X2 U3405 ( .A0(n5390), .A1(n578), .B0(n5432), .B1(n2196), .Y(n8245) );
  CLKMX2X3 U3406 ( .A(n7477), .B(n7476), .S0(net114081), .Y(net110953) );
  OAI221X2 U3407 ( .A0(n5329), .A1(n411), .B0(n5355), .B1(n255), .C0(n6416), 
        .Y(n6417) );
  AOI2BB2X4 U3408 ( .B0(n3763), .B1(\D_cache/cache[4][58] ), .A0N(n5361), 
        .A1N(n2033), .Y(n7445) );
  INVX16 U3409 ( .A(n3876), .Y(n3879) );
  CLKINVX12 U3410 ( .A(n9534), .Y(n3876) );
  BUFX20 U3411 ( .A(n5224), .Y(n5210) );
  MXI2X2 U3412 ( .A(n7738), .B(n7737), .S0(net114081), .Y(net119020) );
  OAI21X4 U3413 ( .A0(n3831), .A1(net112512), .B0(n9123), .Y(n3765) );
  AOI211X2 U3414 ( .A0(n3777), .A1(n8557), .B0(n7485), .C0(n7484), .Y(n7502)
         );
  OA22X2 U3415 ( .A0(n7496), .A1(net107210), .B0(n3774), .B1(n3624), .Y(n7497)
         );
  AO22X1 U3416 ( .A0(net118239), .A1(n197), .B0(net118253), .B1(n912), .Y(
        n9240) );
  NAND4X2 U3417 ( .A(n9238), .B(n9237), .C(n9236), .D(n9235), .Y(n9243) );
  MXI2X2 U3418 ( .A(net107656), .B(net107657), .S0(n8289), .Y(n8297) );
  BUFX20 U3419 ( .A(n9537), .Y(n3766) );
  XOR2X4 U3420 ( .A(n6418), .B(n12955), .Y(n6425) );
  OA22X4 U3421 ( .A0(n138), .A1(n2067), .B0(n5694), .B1(n442), .Y(n11138) );
  NAND2X6 U3422 ( .A(n6403), .B(n1941), .Y(n4378) );
  INVXL U3423 ( .A(net105265), .Y(n3768) );
  INVX1 U3424 ( .A(n3768), .Y(n3769) );
  CLKINVX1 U3425 ( .A(n8199), .Y(n8207) );
  NAND2X6 U3426 ( .A(\i_MIPS/ALUin1[12] ), .B(n6690), .Y(n8199) );
  NOR2X6 U3427 ( .A(n6424), .B(n6425), .Y(n6445) );
  AND4X8 U3428 ( .A(n9946), .B(\i_MIPS/EX_MEM_1 ), .C(DCACHE_ren), .D(n11374), 
        .Y(n3892) );
  INVX20 U3429 ( .A(n3892), .Y(n9536) );
  NAND2XL U3430 ( .A(net105375), .B(net105376), .Y(n10443) );
  OA22X1 U3431 ( .A0(n5333), .A1(n967), .B0(n5360), .B1(n2592), .Y(n7798) );
  AOI2BB2X4 U3432 ( .B0(n3856), .B1(\D_cache/cache[2][139] ), .A0N(n5303), 
        .A1N(n2034), .Y(n6399) );
  OR2X4 U3433 ( .A(net112328), .B(net117713), .Y(n3813) );
  AOI2BB2XL U3434 ( .B0(n4016), .B1(\D_cache/cache[4][21] ), .A0N(n5357), 
        .A1N(n2889), .Y(n8921) );
  AND3X4 U3435 ( .A(n3966), .B(n3930), .C(n5055), .Y(n4016) );
  NAND2X6 U3436 ( .A(n3772), .B(n3773), .Y(n3771) );
  XNOR2X4 U3437 ( .A(n4348), .B(n4349), .Y(n3772) );
  NAND2X6 U3438 ( .A(n6955), .B(n347), .Y(n9429) );
  NAND2X1 U3439 ( .A(n9429), .B(n11110), .Y(n9434) );
  INVX4 U3440 ( .A(n145), .Y(n6955) );
  INVX12 U3441 ( .A(net139838), .Y(n3774) );
  AND2X8 U3442 ( .A(net112392), .B(net112393), .Y(net139838) );
  AOI211X2 U3443 ( .A0(n8485), .A1(n8379), .B0(net107841), .C0(n8378), .Y(
        n8391) );
  NAND2X8 U3444 ( .A(\i_MIPS/ALUin1[13] ), .B(n6697), .Y(net110131) );
  MX2X1 U3445 ( .A(net107657), .B(net107656), .S0(n7591), .Y(n7589) );
  XOR2X4 U3446 ( .A(n3775), .B(net104906), .Y(n4326) );
  NAND2X2 U3447 ( .A(n6435), .B(n3018), .Y(n4399) );
  INVX12 U3448 ( .A(n5060), .Y(n5058) );
  AOI211X2 U3449 ( .A0(net107652), .A1(n9322), .B0(n9321), .C0(n9320), .Y(
        n9323) );
  AOI2BB1X4 U3450 ( .A0N(n5049), .A1N(n9208), .B0(n9207), .Y(n9214) );
  INVX1 U3451 ( .A(n9210), .Y(n8290) );
  AO22X1 U3452 ( .A0(net118239), .A1(n212), .B0(net118261), .B1(n936), .Y(
        n9249) );
  NAND4X2 U3453 ( .A(n9247), .B(n9246), .C(n9245), .D(n9244), .Y(n9252) );
  INVX4 U3454 ( .A(net104725), .Y(n4355) );
  NAND2X1 U3455 ( .A(n8485), .B(n7680), .Y(n7045) );
  OAI2BB1X4 U3456 ( .A0N(net104721), .A1N(n10783), .B0(n3989), .Y(net109042)
         );
  OR2X6 U3457 ( .A(n8959), .B(net117731), .Y(n3936) );
  NAND2X6 U3458 ( .A(n10981), .B(n10982), .Y(n6413) );
  MX2X1 U3459 ( .A(\I_cache/cache[7][148] ), .B(n11197), .S0(n5849), .Y(n11654) );
  INVX4 U3460 ( .A(net117631), .Y(net117625) );
  OA22X2 U3461 ( .A0(n10805), .A1(n3878), .B0(n10808), .B1(n4495), .Y(n8004)
         );
  INVX8 U3462 ( .A(n11396), .Y(n10410) );
  OAI2BB1X4 U3463 ( .A0N(net105232), .A1N(net105233), .B0(n3989), .Y(net109529) );
  XOR2X1 U3464 ( .A(n3001), .B(n10846), .Y(n6757) );
  NOR4X4 U3465 ( .A(n6758), .B(n6757), .C(n6756), .D(n6755), .Y(n6759) );
  OA22X2 U3466 ( .A0(n10705), .A1(n3878), .B0(n10708), .B1(n4495), .Y(n9535)
         );
  NAND4X2 U3467 ( .A(n9520), .B(n9519), .C(n9518), .D(n9517), .Y(n11503) );
  XOR2X2 U3468 ( .A(\i_MIPS/jump_addr[26] ), .B(n10847), .Y(n6755) );
  AOI21X2 U3469 ( .A0(n8477), .A1(net109179), .B0(n8476), .Y(n4753) );
  OAI2BB1X4 U3470 ( .A0N(n8758), .A1N(n8757), .B0(n3970), .Y(n4015) );
  INVX1 U3471 ( .A(n11483), .Y(n10784) );
  NAND4X2 U3472 ( .A(n8515), .B(n8514), .C(n8513), .D(n8512), .Y(n11483) );
  OA22X1 U3473 ( .A0(n5330), .A1(n968), .B0(n5357), .B1(n2593), .Y(n8513) );
  NOR2X1 U3474 ( .A(net107210), .B(n8027), .Y(n3779) );
  INVX1 U3475 ( .A(net117757), .Y(n3781) );
  AO22X4 U3476 ( .A0(n9307), .A1(net117747), .B0(n3950), .B1(n9306), .Y(n9311)
         );
  NOR2X8 U3477 ( .A(n3705), .B(n9544), .Y(n4756) );
  INVX20 U3478 ( .A(n5051), .Y(n9544) );
  CLKINVX3 U3479 ( .A(net104891), .Y(net111129) );
  OAI221X1 U3480 ( .A0(n8790), .A1(n9550), .B0(n5049), .B1(n8789), .C0(
        net107389), .Y(n8791) );
  INVX12 U3481 ( .A(net118597), .Y(net107656) );
  MX2X2 U3482 ( .A(net107656), .B(net107657), .S0(n8377), .Y(n8378) );
  OA22X4 U3483 ( .A0(n138), .A1(n532), .B0(n5694), .B1(n2929), .Y(n11130) );
  AOI21X4 U3484 ( .A0(n9734), .A1(n3634), .B0(n11584), .Y(n4738) );
  AO22X4 U3485 ( .A0(mem_rdata_I[35]), .A1(n5944), .B0(n5568), .B1(n11253), 
        .Y(n10944) );
  NAND2X4 U3486 ( .A(n5051), .B(n3705), .Y(n3862) );
  AOI222X4 U3487 ( .A0(n4735), .A1(net109168), .B0(net107652), .B1(n8961), 
        .C0(n8042), .C1(net109965), .Y(n8047) );
  MX2XL U3488 ( .A(DCACHE_addr[16]), .B(net104964), .S0(n3595), .Y(
        \i_MIPS/n381 ) );
  NAND2X8 U3489 ( .A(n3837), .B(n6952), .Y(n7597) );
  AOI21X4 U3490 ( .A0(n8372), .A1(n8291), .B0(n4724), .Y(n4715) );
  OAI221X2 U3491 ( .A0(n2892), .A1(n5064), .B0(n343), .B1(n5056), .C0(n6670), 
        .Y(n8386) );
  INVX8 U3492 ( .A(net112534), .Y(net112392) );
  AOI2BB1X1 U3493 ( .A0N(\i_MIPS/PC/n27 ), .A1N(net115789), .B0(n11057), .Y(
        n11058) );
  OA22X4 U3494 ( .A0(n345), .A1(n5063), .B0(n2919), .B1(n5057), .Y(n8109) );
  OA22X2 U3495 ( .A0(n5407), .A1(n582), .B0(n5446), .B1(n2200), .Y(n6450) );
  NAND4X2 U3496 ( .A(n8669), .B(n8671), .C(n8670), .D(n8672), .Y(n8675) );
  NAND2X1 U3497 ( .A(net108851), .B(n8648), .Y(n8662) );
  AND4X2 U3498 ( .A(n3726), .B(n8636), .C(n4726), .D(net108787), .Y(n4752) );
  AOI222X2 U3499 ( .A0(n4535), .A1(n11495), .B0(mem_rdata_D[119]), .B1(n130), 
        .C0(n12990), .C1(n5534), .Y(n10688) );
  OA22X1 U3500 ( .A0(\i_MIPS/Register/register[6][13] ), .A1(n5082), .B0(
        \i_MIPS/Register/register[14][13] ), .B1(n5078), .Y(n8006) );
  AOI2BB1X2 U3501 ( .A0N(n7773), .A1N(n3629), .B0(n7771), .Y(n7774) );
  OA22X4 U3502 ( .A0(n10397), .A1(n3877), .B0(n10400), .B1(n4495), .Y(n7717)
         );
  NAND2X6 U3503 ( .A(n4619), .B(net111416), .Y(n7487) );
  INVX12 U3504 ( .A(n7222), .Y(n6712) );
  OA22X4 U3505 ( .A0(net107210), .A1(n8201), .B0(n3774), .B1(net109666), .Y(
        n8219) );
  INVX3 U3506 ( .A(n7858), .Y(n8882) );
  AOI21X4 U3507 ( .A0(n6916), .A1(n4638), .B0(n7858), .Y(n6924) );
  AND4X6 U3508 ( .A(n3926), .B(n3925), .C(n3927), .D(n3928), .Y(n6444) );
  MX2X1 U3509 ( .A(n7422), .B(n7790), .S0(net114065), .Y(n7423) );
  NAND2X1 U3510 ( .A(net111572), .B(n3833), .Y(n9124) );
  AND4X4 U3511 ( .A(n8787), .B(n8786), .C(n8785), .D(n8784), .Y(n3959) );
  NAND4X6 U3512 ( .A(n3959), .B(n8796), .C(n8795), .D(n8794), .Y(net105167) );
  AOI33X2 U3513 ( .A0(net117743), .A1(n3560), .A2(n9224), .B0(net117743), .B1(
        n8788), .B2(n8781), .Y(n8787) );
  OA22X1 U3514 ( .A0(n5333), .A1(n969), .B0(n5360), .B1(n2594), .Y(n7702) );
  NAND4X4 U3515 ( .A(n7704), .B(n7703), .C(n7702), .D(n7701), .Y(n11499) );
  CLKINVX1 U3516 ( .A(n7430), .Y(n3905) );
  OA22X2 U3517 ( .A0(n9202), .A1(n9201), .B0(n9200), .B1(n9550), .Y(n9215) );
  INVX8 U3518 ( .A(n7402), .Y(n7405) );
  NAND2X4 U3519 ( .A(n4739), .B(n9432), .Y(n7402) );
  AO22X1 U3520 ( .A0(n10538), .A1(n4544), .B0(net104801), .B1(n10537), .Y(
        \i_MIPS/N45 ) );
  OA22XL U3521 ( .A0(n4695), .A1(n10736), .B0(\i_MIPS/PC/n2 ), .B1(net115799), 
        .Y(n10737) );
  NAND2X2 U3522 ( .A(n3787), .B(n10987), .Y(n4379) );
  CLKMX2X2 U3523 ( .A(n8594), .B(n8593), .S0(net114085), .Y(n8595) );
  OA22X4 U3524 ( .A0(n5049), .A1(n8299), .B0(n9206), .B1(n9133), .Y(n8302) );
  INVX6 U3525 ( .A(n7772), .Y(n6655) );
  CLKAND2X12 U3526 ( .A(n8780), .B(n9222), .Y(n4729) );
  NAND2X6 U3527 ( .A(n4276), .B(n4277), .Y(net110430) );
  NOR4BX2 U3528 ( .AN(n3790), .B(n8564), .C(n8563), .D(n8562), .Y(n8572) );
  INVX8 U3529 ( .A(n11448), .Y(n10650) );
  NAND4X4 U3530 ( .A(n8168), .B(n8167), .C(n8166), .D(n8165), .Y(n11448) );
  BUFX20 U3531 ( .A(n5194), .Y(n5193) );
  AND2X2 U3532 ( .A(n6677), .B(n4682), .Y(n6679) );
  NAND2X2 U3533 ( .A(n4755), .B(\i_MIPS/ALUin1[26] ), .Y(n7588) );
  XNOR2X4 U3534 ( .A(ICACHE_addr[9]), .B(n11351), .Y(n11134) );
  NAND4X4 U3535 ( .A(n11117), .B(n11116), .C(n11115), .D(n11114), .Y(n11351)
         );
  NAND3X6 U3536 ( .A(n7301), .B(n6709), .C(n8120), .Y(n7490) );
  INVX4 U3537 ( .A(net104957), .Y(n4335) );
  AO21X4 U3538 ( .A0(n7683), .A1(n8291), .B0(n4724), .Y(n8460) );
  INVX1 U3539 ( .A(n8460), .Y(n7684) );
  NOR3X8 U3540 ( .A(n3791), .B(n3792), .C(n3793), .Y(n3920) );
  OR2X8 U3541 ( .A(n6457), .B(n6456), .Y(n3792) );
  NOR2X4 U3542 ( .A(n4449), .B(n3661), .Y(n9911) );
  NAND2X8 U3543 ( .A(n6654), .B(n3895), .Y(n9301) );
  MX2X1 U3544 ( .A(\D_cache/cache[0][6] ), .B(n9942), .S0(n3565), .Y(
        \D_cache/n1748 ) );
  INVX8 U3545 ( .A(n3819), .Y(n9942) );
  NOR3X4 U3546 ( .A(n4470), .B(n4471), .C(n4472), .Y(n9660) );
  CLKINVX20 U3547 ( .A(n1985), .Y(mem_addr_D[19]) );
  NOR3X4 U3548 ( .A(n4446), .B(n4447), .C(n4448), .Y(n9933) );
  NOR2BX1 U3549 ( .AN(net104171), .B(n3795), .Y(n4461) );
  NOR2BX1 U3550 ( .AN(net104171), .B(n3796), .Y(n4490) );
  NOR2BX1 U3551 ( .AN(net104171), .B(n3797), .Y(n4467) );
  BUFX20 U3552 ( .A(n10970), .Y(n3800) );
  NAND2X6 U3553 ( .A(n9731), .B(net115797), .Y(n10721) );
  OA22X1 U3554 ( .A0(n5751), .A1(n970), .B0(n5695), .B1(n2595), .Y(n11158) );
  NOR2BX1 U3555 ( .AN(net104171), .B(n3807), .Y(n4464) );
  NOR3X4 U3556 ( .A(n4455), .B(n4456), .C(n4457), .Y(n9845) );
  CLKAND2X2 U3557 ( .A(n3663), .B(n11260), .Y(n4456) );
  AOI2BB1X1 U3558 ( .A0N(\i_MIPS/PC/n26 ), .A1N(net115799), .B0(n10366), .Y(
        n10367) );
  INVX3 U3559 ( .A(n5564), .Y(n4641) );
  NAND3BX2 U3560 ( .AN(n10728), .B(n5564), .C(n10727), .Y(n10729) );
  CLKINVX4 U3561 ( .A(n10726), .Y(n10727) );
  OA22X1 U3562 ( .A0(n5335), .A1(n1275), .B0(n5356), .B1(n2904), .Y(n6559) );
  CLKAND2X2 U3563 ( .A(net104172), .B(n11261), .Y(n4444) );
  XNOR2X4 U3564 ( .A(n4279), .B(net105250), .Y(n3815) );
  XNOR2X4 U3565 ( .A(n4359), .B(net105746), .Y(n3816) );
  XNOR2X4 U3566 ( .A(net104884), .B(n3997), .Y(n3817) );
  XNOR2X4 U3567 ( .A(n4358), .B(net106290), .Y(n3818) );
  OR2X6 U3568 ( .A(n3937), .B(n5026), .Y(net104940) );
  AOI222X1 U3569 ( .A0(n4535), .A1(n11485), .B0(mem_rdata_D[109]), .B1(n130), 
        .C0(n13000), .C1(n5534), .Y(n10800) );
  MX2X4 U3570 ( .A(n9941), .B(n9940), .S0(n5542), .Y(n3819) );
  AOI222X1 U3571 ( .A0(n5541), .A1(n11424), .B0(mem_rdata_D[48]), .B1(n133), 
        .C0(n12997), .C1(n5539), .Y(n10509) );
  CLKAND2X2 U3572 ( .A(n3898), .B(n11309), .Y(n4460) );
  NAND2XL U3573 ( .A(DCACHE_addr[2]), .B(\i_MIPS/n266 ), .Y(net106602) );
  INVX6 U3574 ( .A(n8878), .Y(n8485) );
  CLKINVX20 U3575 ( .A(n3822), .Y(n10645) );
  OAI211X2 U3576 ( .A0(n8879), .A1(n8878), .B0(n8877), .C0(n8876), .Y(n8898)
         );
  OAI221X2 U3577 ( .A0(n10050), .A1(net143858), .B0(\i_MIPS/n496 ), .B1(
        net115793), .C0(n10049), .Y(\i_MIPS/N74 ) );
  AOI222X1 U3578 ( .A0(n4535), .A1(n11488), .B0(mem_rdata_D[112]), .B1(n131), 
        .C0(n12997), .C1(n5534), .Y(n10500) );
  AOI222X1 U3579 ( .A0(n4535), .A1(n11482), .B0(mem_rdata_D[106]), .B1(n132), 
        .C0(n13003), .C1(n5534), .Y(n10772) );
  CLKINVX20 U3580 ( .A(n3823), .Y(n10658) );
  INVX12 U3581 ( .A(n4533), .Y(n4534) );
  CLKINVX20 U3582 ( .A(n3824), .Y(n10603) );
  CLKINVX20 U3583 ( .A(n3825), .Y(n10697) );
  AOI222X4 U3584 ( .A0(n3800), .A1(n11379), .B0(mem_rdata_D[3]), .B1(n129), 
        .C0(n13010), .C1(n5538), .Y(n10763) );
  CLKINVX20 U3585 ( .A(n3826), .Y(n10672) );
  MXI2X4 U3586 ( .A(n9948), .B(n9947), .S0(n5542), .Y(n9949) );
  AOI222X4 U3587 ( .A0(n4506), .A1(n11446), .B0(mem_rdata_D[70]), .B1(n133), 
        .C0(n13007), .C1(n5535), .Y(n9948) );
  OAI221X2 U3588 ( .A0(n9795), .A1(net143858), .B0(\i_MIPS/n501 ), .B1(
        net115791), .C0(n9794), .Y(\i_MIPS/N69 ) );
  BUFX20 U3589 ( .A(n10504), .Y(n4550) );
  AOI222X4 U3590 ( .A0(n4506), .A1(n11456), .B0(mem_rdata_D[80]), .B1(n131), 
        .C0(n12997), .C1(n5535), .Y(n10503) );
  AOI222X1 U3591 ( .A0(n4534), .A1(n11483), .B0(mem_rdata_D[107]), .B1(n131), 
        .C0(n13002), .C1(n5534), .Y(n10785) );
  CLKAND2X2 U3592 ( .A(net104171), .B(n11232), .Y(n4452) );
  AOI222X1 U3593 ( .A0(n4506), .A1(n11461), .B0(mem_rdata_D[85]), .B1(n132), 
        .C0(n12992), .C1(n5536), .Y(n10518) );
  AOI222X1 U3594 ( .A0(n4506), .A1(n11468), .B0(mem_rdata_D[92]), .B1(n133), 
        .C0(n12985), .C1(n5536), .Y(n10546) );
  AOI222X1 U3595 ( .A0(n4506), .A1(n11467), .B0(mem_rdata_D[91]), .B1(n132), 
        .C0(n12986), .C1(n5535), .Y(n10395) );
  AOI222X1 U3596 ( .A0(n4506), .A1(n11462), .B0(mem_rdata_D[86]), .B1(n131), 
        .C0(n12991), .C1(n5535), .Y(n10311) );
  AOI222X1 U3597 ( .A0(n4506), .A1(n11450), .B0(mem_rdata_D[74]), .B1(n133), 
        .C0(n13003), .C1(n5535), .Y(n10775) );
  OAI211X4 U3598 ( .A0(n3648), .A1(net106828), .B0(n9935), .C0(net135522), .Y(
        net104168) );
  AO22X2 U3599 ( .A0(n5939), .A1(ICACHE_addr[12]), .B0(n5930), .B1(n11354), 
        .Y(n11177) );
  AO22X2 U3600 ( .A0(n5933), .A1(ICACHE_addr[19]), .B0(n5930), .B1(n11361), 
        .Y(n11201) );
  AO22X2 U3601 ( .A0(n5939), .A1(ICACHE_addr[7]), .B0(n5930), .B1(n11349), .Y(
        n11155) );
  AO22X2 U3602 ( .A0(n5939), .A1(ICACHE_addr[14]), .B0(n5930), .B1(n11356), 
        .Y(n11172) );
  AO22X2 U3603 ( .A0(n5939), .A1(ICACHE_addr[8]), .B0(n5930), .B1(n11350), .Y(
        n11159) );
  AO22X2 U3604 ( .A0(n5939), .A1(ICACHE_addr[6]), .B0(n5930), .B1(n11348), .Y(
        n11164) );
  AO22X2 U3605 ( .A0(n5939), .A1(ICACHE_addr[17]), .B0(n5930), .B1(n11359), 
        .Y(n11150) );
  AO22X2 U3606 ( .A0(n5937), .A1(ICACHE_addr[26]), .B0(n5930), .B1(n11368), 
        .Y(n11187) );
  AO22X2 U3607 ( .A0(n5937), .A1(ICACHE_addr[24]), .B0(n5930), .B1(n11366), 
        .Y(n11192) );
  AO22XL U3608 ( .A0(ICACHE_addr[12]), .A1(mem_read_I), .B0(n5047), .B1(n11354), .Y(n12872) );
  XOR2X4 U3609 ( .A(n11354), .B(ICACHE_addr[12]), .Y(n11597) );
  OAI221X2 U3610 ( .A0(n10867), .A1(net143858), .B0(\i_MIPS/n517 ), .B1(
        net115789), .C0(n10866), .Y(\i_MIPS/N53 ) );
  AOI222X2 U3611 ( .A0(n4506), .A1(n11443), .B0(mem_rdata_D[67]), .B1(n132), 
        .C0(n13010), .C1(n5536), .Y(n10760) );
  BUFX16 U3612 ( .A(n3660), .Y(n5564) );
  BUFX12 U3613 ( .A(n3660), .Y(n5563) );
  AO21X4 U3614 ( .A0(n10585), .A1(n10584), .B0(n5562), .Y(n10586) );
  INVX6 U3615 ( .A(n10578), .Y(n10583) );
  INVXL U3616 ( .A(n10487), .Y(n10489) );
  NAND2X1 U3617 ( .A(\i_MIPS/IF_ID[5] ), .B(\i_MIPS/Sign_Extend[3] ), .Y(
        n10155) );
  AOI222X4 U3618 ( .A0(n8463), .A1(n7480), .B0(n7479), .B1(net118584), .C0(
        n8461), .C1(n3714), .Y(n7504) );
  XNOR2X4 U3619 ( .A(n3828), .B(net105329), .Y(n4331) );
  OAI221X2 U3620 ( .A0(\i_MIPS/n297 ), .A1(n5072), .B0(\i_MIPS/n296 ), .B1(
        n5068), .C0(n7036), .Y(n7675) );
  NOR2X6 U3621 ( .A(n3964), .B(n4674), .Y(n6649) );
  MX2X1 U3622 ( .A(net107657), .B(net107656), .S0(n8134), .Y(n8135) );
  INVX20 U3623 ( .A(n4504), .Y(n4505) );
  CLKINVX12 U3624 ( .A(n10966), .Y(n4504) );
  NAND4X4 U3625 ( .A(n9015), .B(n9014), .C(n9013), .D(n9012), .Y(n11377) );
  OA22X2 U3626 ( .A0(n5332), .A1(n563), .B0(n5357), .B1(n2185), .Y(n9013) );
  MX2X1 U3627 ( .A(net107656), .B(net107657), .S0(n8212), .Y(n8213) );
  OAI221X2 U3628 ( .A0(n9890), .A1(net143858), .B0(\i_MIPS/n512 ), .B1(
        net115791), .C0(n9889), .Y(\i_MIPS/N58 ) );
  OAI221X2 U3629 ( .A0(net108148), .A1(net108149), .B0(n3672), .B1(n3637), 
        .C0(net108010), .Y(n9304) );
  MXI2X4 U3630 ( .A(n10392), .B(n10391), .S0(n5543), .Y(n10393) );
  OR2X8 U3631 ( .A(n10576), .B(\i_MIPS/PC/n31 ), .Y(n10714) );
  OA22X4 U3632 ( .A0(n10505), .A1(n3878), .B0(n10508), .B1(n4495), .Y(n8833)
         );
  NAND4X4 U3633 ( .A(n11375), .B(n3789), .C(n11373), .D(n11539), .Y(n11506) );
  AOI222X2 U3634 ( .A0(n4534), .A1(n11472), .B0(mem_rdata_D[96]), .B1(n133), 
        .C0(n13013), .C1(n5534), .Y(n10739) );
  NAND4X1 U3635 ( .A(n5564), .B(n10726), .C(n10725), .D(n10728), .Y(n10730) );
  OAI2BB1X2 U3636 ( .A0N(\i_MIPS/n506 ), .A1N(n10723), .B0(n10722), .Y(n10726)
         );
  NOR3X4 U3637 ( .A(n4437), .B(n4438), .C(n4439), .Y(n10252) );
  OAI211XL U3638 ( .A0(n3764), .A1(net110131), .B0(net110406), .C0(net108625), 
        .Y(n3830) );
  CLKAND2X12 U3639 ( .A(n8969), .B(net108300), .Y(n3831) );
  AND4X8 U3640 ( .A(n8632), .B(n4882), .C(n6669), .D(net112393), .Y(net134876)
         );
  OA22X2 U3641 ( .A0(n5330), .A1(n585), .B0(n5359), .B1(n2203), .Y(n8080) );
  NAND4X4 U3642 ( .A(n8082), .B(n8081), .C(n8080), .D(n8079), .Y(n11385) );
  AND3X8 U3643 ( .A(n7607), .B(n3832), .C(n7609), .Y(n4090) );
  AOI222X4 U3644 ( .A0(n3800), .A1(n11377), .B0(mem_rdata_D[1]), .B1(n129), 
        .C0(n13012), .C1(n5538), .Y(n10668) );
  INVXL U3645 ( .A(net105424), .Y(n3954) );
  OAI2BB1X4 U3646 ( .A0N(net104940), .A1N(net104939), .B0(n3989), .Y(net109675) );
  OAI221X2 U3647 ( .A0(n9661), .A1(net143858), .B0(\i_MIPS/n257 ), .B1(
        net115789), .C0(n9660), .Y(\i_MIPS/N80 ) );
  INVX3 U3648 ( .A(n11451), .Y(n10787) );
  NAND4X2 U3649 ( .A(n8519), .B(n8518), .C(n8517), .D(n8516), .Y(n11451) );
  OAI221X4 U3650 ( .A0(\i_MIPS/Register/register[18][1] ), .A1(net117641), 
        .B0(\i_MIPS/Register/register[26][1] ), .B1(net117661), .C0(n8997), 
        .Y(n9000) );
  BUFX16 U3651 ( .A(net117639), .Y(net117643) );
  OA22X1 U3652 ( .A0(\i_MIPS/Register/register[6][4] ), .A1(net117681), .B0(
        \i_MIPS/Register/register[14][4] ), .B1(net117695), .Y(n9063) );
  OAI21X4 U3653 ( .A0(n3757), .A1(n3952), .B0(n3989), .Y(net108642) );
  OAI221X2 U3654 ( .A0(n9609), .A1(net143858), .B0(\i_MIPS/n247 ), .B1(
        net115789), .C0(n9608), .Y(\i_MIPS/N75 ) );
  INVXL U3655 ( .A(n8959), .Y(n3836) );
  AO22X4 U3656 ( .A0(n3777), .A1(n8858), .B0(n8857), .B1(n9314), .Y(n8872) );
  AO21X4 U3657 ( .A0(net104940), .A1(net104939), .B0(net117625), .Y(net105820)
         );
  INVXL U3658 ( .A(net104940), .Y(n3941) );
  OR3X6 U3659 ( .A(n6954), .B(n6953), .C(n9433), .Y(n3837) );
  OR2X2 U3660 ( .A(n11094), .B(net143858), .Y(n3838) );
  OR2XL U3661 ( .A(\i_MIPS/n502 ), .B(net115789), .Y(n3839) );
  OR2X2 U3662 ( .A(n9769), .B(net143858), .Y(n3843) );
  OR2XL U3663 ( .A(\i_MIPS/n505 ), .B(net115791), .Y(n3844) );
  NAND3X2 U3664 ( .A(n3843), .B(n3844), .C(n9768), .Y(\i_MIPS/N65 ) );
  AND2X1 U3665 ( .A(net104171), .B(n11235), .Y(n3845) );
  NOR3X2 U3666 ( .A(n3845), .B(n3846), .C(n3847), .Y(n9768) );
  CLKMX2X3 U3667 ( .A(n9078), .B(n9077), .S0(net114085), .Y(n9079) );
  NOR4X2 U3668 ( .A(n9076), .B(n9075), .C(n9074), .D(n9073), .Y(n9077) );
  INVXL U3669 ( .A(n9219), .Y(n3849) );
  OR2X8 U3670 ( .A(n3848), .B(n3849), .Y(n9226) );
  NAND3BX2 U3671 ( .AN(n9221), .B(n3950), .C(n9226), .Y(n9234) );
  OA21X2 U3672 ( .A0(\i_MIPS/ALUin1[13] ), .A1(n5068), .B0(n7299), .Y(n7300)
         );
  OAI22X4 U3673 ( .A0(n11578), .A1(n11577), .B0(n4726), .B1(n11578), .Y(n11581) );
  AO21X4 U3674 ( .A0(n11100), .A1(n126), .B0(n11098), .Y(n11578) );
  NAND4X2 U3675 ( .A(n8297), .B(n8296), .C(net107389), .D(n8295), .Y(n8305) );
  OA22X2 U3676 ( .A0(n9202), .A1(n9132), .B0(n8459), .B1(n9550), .Y(n8295) );
  INVX8 U3677 ( .A(n11399), .Y(n10692) );
  NAND4X4 U3678 ( .A(n7072), .B(n7071), .C(n7070), .D(n7069), .Y(n11399) );
  MX2XL U3679 ( .A(n6713), .B(n12), .S0(n3584), .Y(n3852) );
  CLKINVX1 U3680 ( .A(net108625), .Y(net108624) );
  OA22X4 U3681 ( .A0(net107217), .A1(net108625), .B0(net107228), .B1(net107688), .Y(n4302) );
  NAND2X2 U3682 ( .A(\i_MIPS/ALUin1[15] ), .B(net112446), .Y(net108625) );
  OAI221X4 U3683 ( .A0(n183), .A1(n5064), .B0(n2949), .B1(n5057), .C0(n7153), 
        .Y(n7480) );
  OAI221X4 U3684 ( .A0(n4021), .A1(net143504), .B0(net143514), .B1(
        \i_MIPS/n242 ), .C0(\i_MIPS/n300 ), .Y(net108300) );
  CLKINVX8 U3685 ( .A(n9219), .Y(n8783) );
  OAI211X2 U3686 ( .A0(net110429), .A1(net111724), .B0(n6701), .C0(n8283), .Y(
        n3853) );
  NAND2X6 U3687 ( .A(n6689), .B(n345), .Y(n8859) );
  CLKINVX6 U3688 ( .A(n6693), .Y(n6697) );
  NOR4X4 U3689 ( .A(n9153), .B(n9152), .C(n9151), .D(n9150), .Y(n9164) );
  OA22XL U3690 ( .A0(\i_MIPS/Register/register[6][3] ), .A1(net117681), .B0(
        \i_MIPS/Register/register[14][3] ), .B1(net117703), .Y(n9149) );
  AOI2BB2X4 U3691 ( .B0(n3856), .B1(\D_cache/cache[2][148] ), .A0N(n5306), 
        .A1N(n2036), .Y(n6431) );
  AOI2BB2X4 U3692 ( .B0(n3863), .B1(\D_cache/cache[6][148] ), .A0N(n5446), 
        .A1N(n2037), .Y(n6433) );
  OR2X8 U3693 ( .A(net108161), .B(net117731), .Y(n3991) );
  OA22X4 U3694 ( .A0(n5406), .A1(n2068), .B0(n5445), .B1(n443), .Y(n6465) );
  MXI2X1 U3695 ( .A(\i_MIPS/n203 ), .B(\i_MIPS/n204 ), .S0(n3595), .Y(
        \i_MIPS/n326 ) );
  NOR4X4 U3696 ( .A(n9162), .B(n9161), .C(n9160), .D(n9159), .Y(n9163) );
  OA22XL U3697 ( .A0(\i_MIPS/Register/register[22][3] ), .A1(net117681), .B0(
        \i_MIPS/Register/register[30][3] ), .B1(net117703), .Y(n9158) );
  OA22X4 U3698 ( .A0(n5407), .A1(n2070), .B0(n5446), .B1(n445), .Y(n6437) );
  NAND2X4 U3699 ( .A(n5062), .B(\i_MIPS/ALUin1[18] ), .Y(n7417) );
  INVX4 U3700 ( .A(n8114), .Y(n3858) );
  INVX8 U3701 ( .A(n8687), .Y(n8644) );
  NAND2X6 U3702 ( .A(\i_MIPS/ALUin1[18] ), .B(n4503), .Y(n8687) );
  OA22X1 U3703 ( .A0(n2920), .A1(n5063), .B0(n300), .B1(n5057), .Y(n7412) );
  OA22X1 U3704 ( .A0(n2937), .A1(n5063), .B0(\i_MIPS/n287 ), .B1(n5057), .Y(
        n7418) );
  OA22X1 U3705 ( .A0(\i_MIPS/ALUin1[21] ), .A1(n5063), .B0(\i_MIPS/ALUin1[22] ), .B1(n5057), .Y(n7408) );
  OA22X1 U3706 ( .A0(\i_MIPS/ALUin1[8] ), .A1(n5064), .B0(\i_MIPS/ALUin1[7] ), 
        .B1(n5057), .Y(n7311) );
  OA22X1 U3707 ( .A0(\i_MIPS/ALUin1[10] ), .A1(n5063), .B0(\i_MIPS/ALUin1[9] ), 
        .B1(n5057), .Y(n8036) );
  OA22X1 U3708 ( .A0(\i_MIPS/ALUin1[26] ), .A1(n5063), .B0(\i_MIPS/ALUin1[27] ), .B1(n5057), .Y(n7673) );
  CLKAND2X12 U3709 ( .A(n8634), .B(n6673), .Y(n4691) );
  NAND2X1 U3710 ( .A(n4682), .B(n7409), .Y(n7414) );
  AOI222X2 U3711 ( .A0(n4688), .A1(n7787), .B0(n8976), .B1(n9450), .C0(n7676), 
        .C1(n8557), .Y(n7413) );
  NAND2X4 U3712 ( .A(\i_MIPS/n299 ), .B(n3691), .Y(n9123) );
  BUFX20 U3713 ( .A(n5311), .Y(n5306) );
  AOI2BB2X4 U3714 ( .B0(n3863), .B1(\D_cache/cache[6][134] ), .A0N(n5444), 
        .A1N(n2038), .Y(n6493) );
  OAI222X1 U3715 ( .A0(net107217), .A1(net110131), .B0(net107661), .B1(n7943), 
        .C0(n7942), .C1(net117757), .Y(n7947) );
  INVX3 U3716 ( .A(n7943), .Y(n6935) );
  AOI2BB2X4 U3717 ( .B0(n3863), .B1(\D_cache/cache[6][132] ), .A0N(n5445), 
        .A1N(n2039), .Y(n6428) );
  BUFX2 U3718 ( .A(n5403), .Y(n5390) );
  OA22X1 U3719 ( .A0(\i_MIPS/ALUin1[23] ), .A1(n5064), .B0(\i_MIPS/ALUin1[24] ), .B1(n5058), .Y(n6672) );
  NAND2X6 U3720 ( .A(\i_MIPS/ALUin1[24] ), .B(n6668), .Y(n6918) );
  NAND2X8 U3721 ( .A(n4621), .B(n4622), .Y(n6714) );
  NAND2X8 U3722 ( .A(n4718), .B(net108632), .Y(net107987) );
  INVX20 U3723 ( .A(net107987), .Y(net107652) );
  OA22X4 U3724 ( .A0(n9134), .A1(net107987), .B0(net107988), .B1(n9133), .Y(
        n9142) );
  NAND4X4 U3725 ( .A(n7804), .B(n7803), .C(n7802), .D(n7801), .Y(n11454) );
  OA22X1 U3726 ( .A0(n5333), .A1(n971), .B0(n5360), .B1(n2596), .Y(n7802) );
  NAND2X6 U3727 ( .A(n6655), .B(n7765), .Y(n7100) );
  INVX8 U3728 ( .A(n9429), .Y(n11113) );
  INVX2 U3729 ( .A(n11472), .Y(n10738) );
  AOI2BB2X4 U3730 ( .B0(n3864), .B1(\D_cache/cache[2][144] ), .A0N(n5305), 
        .A1N(n3865), .Y(n6404) );
  OA22X4 U3731 ( .A0(n5406), .A1(n2073), .B0(n5445), .B1(n448), .Y(n6453) );
  OAI2BB1X4 U3732 ( .A0N(n8380), .A1N(n8381), .B0(n8382), .Y(n8880) );
  NAND2X6 U3733 ( .A(\i_MIPS/ALUin1[19] ), .B(n6687), .Y(n8300) );
  CLKINVX6 U3734 ( .A(n4578), .Y(n6687) );
  CLKBUFX2 U3735 ( .A(net108004), .Y(n3867) );
  CLKBUFX2 U3736 ( .A(n7302), .Y(n3868) );
  NAND3X8 U3737 ( .A(n3869), .B(n3870), .C(n9461), .Y(n10604) );
  AND2X4 U3738 ( .A(n9441), .B(n3950), .Y(n3871) );
  AND2XL U3739 ( .A(n9563), .B(n9541), .Y(n9465) );
  AND4X8 U3740 ( .A(n9460), .B(n9459), .C(n9458), .D(n9457), .Y(n9461) );
  OAI221XL U3741 ( .A0(n9465), .A1(n9464), .B0(n9463), .B1(n9462), .C0(n9461), 
        .Y(n4020) );
  OA22X1 U3742 ( .A0(n5254), .A1(n972), .B0(n5294), .B1(n2597), .Y(n7909) );
  NAND3X4 U3743 ( .A(n3966), .B(n6391), .C(n3930), .Y(n9529) );
  OA22X2 U3744 ( .A0(n5401), .A1(n586), .B0(n5444), .B1(n2204), .Y(n6500) );
  MX2XL U3745 ( .A(n3547), .B(n3677), .S0(n3589), .Y(\i_MIPS/n305 ) );
  OA22X4 U3746 ( .A0(n5243), .A1(n2074), .B0(n5284), .B1(n449), .Y(n9348) );
  CLKINVX12 U3747 ( .A(n5055), .Y(n6391) );
  INVX8 U3748 ( .A(n3873), .Y(n3874) );
  OA22X1 U3749 ( .A0(n5331), .A1(n973), .B0(n5356), .B1(n2598), .Y(n8605) );
  INVX6 U3750 ( .A(n7585), .Y(n9431) );
  BUFX20 U3751 ( .A(n9807), .Y(n5338) );
  NAND4BX2 U3752 ( .AN(n9039), .B(n9038), .C(n9037), .D(n9036), .Y(n9040) );
  AO22X4 U3753 ( .A0(net118217), .A1(net105257), .B0(net118227), .B1(n4280), 
        .Y(net111668) );
  OAI211X2 U3754 ( .A0(n8471), .A1(n8467), .B0(n8199), .C0(n8464), .Y(n7772)
         );
  AOI222X1 U3755 ( .A0(n5541), .A1(n11408), .B0(mem_rdata_D[32]), .B1(n132), 
        .C0(n13013), .C1(n5540), .Y(n10748) );
  OA22X1 U3756 ( .A0(\i_MIPS/ALUin1[9] ), .A1(n5063), .B0(\i_MIPS/ALUin1[8] ), 
        .B1(n5057), .Y(n8130) );
  NAND4X2 U3757 ( .A(n7117), .B(n7116), .C(n7115), .D(n7114), .Y(n11391) );
  CLKMX2X2 U3758 ( .A(n10185), .B(net105746), .S0(n3597), .Y(\i_MIPS/n363 ) );
  BUFX4 U3759 ( .A(n5397), .Y(n5393) );
  INVX3 U3760 ( .A(net108876), .Y(net111723) );
  AOI211X2 U3761 ( .A0(n3776), .A1(n6921), .B0(n7430), .C0(n7407), .Y(n6922)
         );
  NAND2X4 U3762 ( .A(n4709), .B(n7041), .Y(n6921) );
  OA22X2 U3763 ( .A0(n10520), .A1(n3878), .B0(n10523), .B1(n4495), .Y(n8936)
         );
  INVX3 U3764 ( .A(n11429), .Y(n10523) );
  NAND4X4 U3765 ( .A(n8935), .B(n8934), .C(n8933), .D(n8932), .Y(n11429) );
  OA22X1 U3766 ( .A0(n5332), .A1(n974), .B0(n5357), .B1(n2599), .Y(n8933) );
  NAND3X8 U3767 ( .A(n6644), .B(n3029), .C(\i_MIPS/ALU_Control/n20 ), .Y(
        net112393) );
  NAND4X4 U3768 ( .A(\i_MIPS/ID_EX[74] ), .B(n1340), .C(net134414), .D(n3874), 
        .Y(n8632) );
  AO22X4 U3769 ( .A0(n9445), .A1(n8558), .B0(n9442), .B1(n7421), .Y(n7426) );
  INVX16 U3770 ( .A(n3876), .Y(n3877) );
  INVX8 U3771 ( .A(n11480), .Y(n10647) );
  NAND4X4 U3772 ( .A(n8164), .B(n8163), .C(n8162), .D(n8161), .Y(n11480) );
  INVX8 U3773 ( .A(n11053), .Y(n7739) );
  CLKINVX20 U3774 ( .A(n5074), .Y(n5073) );
  INVX1 U3775 ( .A(n3857), .Y(net108853) );
  OAI22X1 U3776 ( .A0(n10186), .A1(n3766), .B0(n10189), .B1(n5189), .Y(n3880)
         );
  OAI22X1 U3777 ( .A0(n10192), .A1(n3877), .B0(n10195), .B1(n4495), .Y(n3881)
         );
  CLKINVX20 U3778 ( .A(n3969), .Y(n3970) );
  XOR2X4 U3779 ( .A(n3882), .B(n5021), .Y(n6502) );
  BUFX16 U3780 ( .A(net117667), .Y(net117657) );
  OA22X1 U3781 ( .A0(\i_MIPS/Register/register[22][12] ), .A1(net117683), .B0(
        \i_MIPS/Register/register[30][12] ), .B1(net117695), .Y(n8234) );
  MX2X1 U3782 ( .A(n8037), .B(n8040), .S0(\i_MIPS/ID_EX[81] ), .Y(n9322) );
  MX2X2 U3783 ( .A(n7682), .B(n7681), .S0(\i_MIPS/ID_EX[81] ), .Y(n8299) );
  INVXL U3784 ( .A(n11011), .Y(n3884) );
  CLKINVX1 U3785 ( .A(n3884), .Y(n3885) );
  CLKINVX4 U3786 ( .A(net111668), .Y(net105581) );
  OA22X2 U3787 ( .A0(n10971), .A1(n3879), .B0(n10975), .B1(n4495), .Y(n8347)
         );
  INVXL U3788 ( .A(net111277), .Y(n3886) );
  INVX4 U3789 ( .A(n143), .Y(n6668) );
  NAND2X8 U3790 ( .A(n3902), .B(n3670), .Y(net108623) );
  INVX8 U3791 ( .A(net118369), .Y(net118359) );
  AND2X2 U3792 ( .A(mem_ready_D), .B(n11504), .Y(n4796) );
  BUFX20 U3793 ( .A(n4714), .Y(n5060) );
  OA22X4 U3794 ( .A0(n1302), .A1(n5064), .B0(n2892), .B1(n5059), .Y(n7036) );
  OA22X2 U3795 ( .A0(n5401), .A1(n588), .B0(n5444), .B1(n2206), .Y(n6506) );
  INVX3 U3796 ( .A(n6497), .Y(n11005) );
  NAND4X2 U3797 ( .A(n7268), .B(n7267), .C(n7266), .D(n7265), .Y(n11446) );
  INVX6 U3798 ( .A(n6434), .Y(n11011) );
  NAND2X6 U3799 ( .A(n7768), .B(n7101), .Y(n4643) );
  OAI221X2 U3800 ( .A0(n3897), .A1(net107210), .B0(net108308), .B1(net107411), 
        .C0(net117759), .Y(net108284) );
  OA22X2 U3801 ( .A0(n137), .A1(n589), .B0(n5695), .B1(n2207), .Y(n11162) );
  OA22X4 U3802 ( .A0(n5832), .A1(n2076), .B0(n5796), .B1(n451), .Y(n11161) );
  BUFX20 U3803 ( .A(n5884), .Y(n5876) );
  OA22X4 U3804 ( .A0(n5918), .A1(n433), .B0(n5876), .B1(n2059), .Y(n11141) );
  BUFX8 U3805 ( .A(n4681), .Y(n5884) );
  CLKINVX8 U3806 ( .A(n7024), .Y(n7039) );
  NAND2X4 U3807 ( .A(\i_MIPS/ALUin1[23] ), .B(n6686), .Y(n7024) );
  AOI2BB1X4 U3808 ( .A0N(n1302), .A1N(n5067), .B0(n4792), .Y(n6670) );
  INVX8 U3809 ( .A(n9127), .Y(n9138) );
  OAI221X4 U3810 ( .A0(n3908), .A1(net144236), .B0(n3894), .B1(n3559), .C0(
        n2928), .Y(n9127) );
  OAI221X2 U3811 ( .A0(n5327), .A1(n2014), .B0(n5352), .B1(n395), .C0(n6465), 
        .Y(n6466) );
  BUFX4 U3812 ( .A(n4658), .Y(n5705) );
  CLKAND2X8 U3813 ( .A(\i_MIPS/EX_MEM_0 ), .B(net107141), .Y(n6765) );
  BUFX20 U3814 ( .A(net139838), .Y(net117751) );
  OAI221X2 U3815 ( .A0(n5172), .A1(n2952), .B0(n5222), .B1(n1311), .C0(n6468), 
        .Y(n6469) );
  NAND2X6 U3816 ( .A(n11014), .B(n11015), .Y(n6430) );
  CLKBUFX2 U3817 ( .A(n10403), .Y(n3888) );
  NAND2X4 U3818 ( .A(net139863), .B(net105364), .Y(n10403) );
  OA22X2 U3819 ( .A0(n5741), .A1(n590), .B0(n5706), .B1(n2208), .Y(n11121) );
  NOR2X8 U3820 ( .A(n7695), .B(n7670), .Y(n4697) );
  OAI221X4 U3821 ( .A0(net107210), .A1(n9306), .B0(n9307), .B1(net107411), 
        .C0(net117759), .Y(n9312) );
  OA22X4 U3822 ( .A0(n10431), .A1(n3766), .B0(n10434), .B1(n9536), .Y(n6871)
         );
  INVX4 U3823 ( .A(n11497), .Y(n10431) );
  OA22XL U3824 ( .A0(n5399), .A1(n1247), .B0(n5443), .B1(n2867), .Y(n6858) );
  CLKINVX12 U3825 ( .A(n6769), .Y(n6776) );
  NAND2X2 U3826 ( .A(\i_MIPS/jump_addr[23] ), .B(\i_MIPS/n499 ), .Y(n6768) );
  OA22X4 U3827 ( .A0(n5381), .A1(n2080), .B0(n5421), .B1(n455), .Y(n9358) );
  OA22X4 U3828 ( .A0(n5920), .A1(n2968), .B0(n5878), .B1(n1320), .Y(n11211) );
  OA22X4 U3829 ( .A0(n5920), .A1(n2081), .B0(n5878), .B1(n435), .Y(n11193) );
  NAND2X6 U3830 ( .A(\i_MIPS/ALUin1[4] ), .B(net112414), .Y(net107680) );
  OAI221X2 U3831 ( .A0(net107210), .A1(net108622), .B0(net111716), .B1(n3774), 
        .C0(net117759), .Y(n4309) );
  BUFX20 U3832 ( .A(n5921), .Y(n5918) );
  NAND3BX4 U3833 ( .AN(net108787), .B(n8632), .C(n4691), .Y(net107224) );
  BUFX20 U3834 ( .A(net107224), .Y(net118597) );
  BUFX20 U3835 ( .A(n5267), .Y(n5265) );
  BUFX20 U3836 ( .A(n9806), .Y(n5267) );
  NAND4X4 U3837 ( .A(n8931), .B(n8930), .C(n8929), .D(n8928), .Y(n11397) );
  OR2X8 U3838 ( .A(n6435), .B(n3018), .Y(n4400) );
  OR2X2 U3839 ( .A(n5329), .B(n2897), .Y(n4627) );
  AO21X2 U3840 ( .A0(net106297), .A1(net106298), .B0(net117625), .Y(net106041)
         );
  AO21X2 U3841 ( .A0(net104889), .A1(net104890), .B0(net117625), .Y(net105835)
         );
  ACHCINX4 U3842 ( .CIN(n10529), .A(\i_MIPS/IF_ID[27] ), .B(n6016), .CO(n10530) );
  OAI2BB2X4 U3843 ( .B0(n3890), .B1(n3891), .A0N(net118217), .A1N(net104765), 
        .Y(net111509) );
  BUFX20 U3844 ( .A(n5338), .Y(n5337) );
  NAND4X2 U3845 ( .A(n11590), .B(n11218), .C(n11217), .D(n11540), .Y(n11344)
         );
  XOR2X4 U3846 ( .A(n11366), .B(ICACHE_addr[24]), .Y(n11601) );
  NAND4X4 U3847 ( .A(n8752), .B(n8751), .C(n8750), .D(n8749), .Y(n11376) );
  OA22X4 U3848 ( .A0(n5063), .A1(n347), .B0(n3861), .B1(n5059), .Y(n7031) );
  BUFX16 U3849 ( .A(n9807), .Y(n5336) );
  NAND4BBX4 U3850 ( .AN(n7164), .BN(n3893), .C(n7163), .D(n7162), .Y(net104765) );
  CLKMX2X4 U3851 ( .A(n3745), .B(n9049), .S0(\i_MIPS/ID_EX[81] ), .Y(n6664) );
  OAI221X4 U3852 ( .A0(n2184), .A1(n5064), .B0(n344), .B1(n5056), .C0(n6662), 
        .Y(n8701) );
  INVX6 U3853 ( .A(n6494), .Y(n11023) );
  AOI21X4 U3854 ( .A0(n7841), .A1(n7041), .B0(n7039), .Y(n4704) );
  AO21X2 U3855 ( .A0(net105423), .A1(net105424), .B0(net117625), .Y(net105364)
         );
  NAND2XL U3856 ( .A(net36572), .B(n11062), .Y(n11213) );
  OA22X4 U3857 ( .A0(n10499), .A1(n3767), .B0(n10502), .B1(n5189), .Y(n8834)
         );
  NAND2XL U3858 ( .A(n3751), .B(n3885), .Y(n11529) );
  CLKINVX20 U3859 ( .A(net143513), .Y(n3894) );
  OA21X4 U3860 ( .A0(n9138), .A1(n7145), .B0(n9126), .Y(n3895) );
  OAI222X2 U3861 ( .A0(net107217), .A1(n8556), .B0(n9206), .B1(n8555), .C0(
        n8554), .C1(net117757), .Y(n8563) );
  AOI221X4 U3862 ( .A0(n3995), .A1(\D_cache/cache[0][149] ), .B0(n5205), .B1(
        \D_cache/cache[1][149] ), .C0(n3932), .Y(n3931) );
  NAND2X8 U3863 ( .A(n6675), .B(net108631), .Y(n9202) );
  MX2X1 U3864 ( .A(net107656), .B(net107657), .S0(n8471), .Y(n8472) );
  CLKINVX1 U3865 ( .A(n6815), .Y(n6816) );
  OA22X4 U3866 ( .A0(n5241), .A1(n2083), .B0(n5282), .B1(n457), .Y(n9356) );
  INVX1 U3867 ( .A(n3896), .Y(n3897) );
  NOR2BX4 U3868 ( .AN(n4719), .B(n9952), .Y(n4686) );
  INVX20 U3869 ( .A(n4875), .Y(mem_addr_D[21]) );
  CLKINVX8 U3870 ( .A(n12846), .Y(n4875) );
  OAI221X4 U3871 ( .A0(\i_MIPS/ALUin1[12] ), .A1(n5064), .B0(
        \i_MIPS/ALUin1[11] ), .B1(n5056), .C0(n7300), .Y(n8480) );
  OAI221X4 U3872 ( .A0(\i_MIPS/ALUin1[20] ), .A1(n5064), .B0(
        \i_MIPS/ALUin1[21] ), .B1(n5056), .C0(n6829), .Y(n6937) );
  OAI221X4 U3873 ( .A0(n300), .A1(n5064), .B0(n3744), .B1(n5056), .C0(n7042), 
        .Y(net110602) );
  OAI221X4 U3874 ( .A0(\i_MIPS/ALUin1[13] ), .A1(n5064), .B0(
        \i_MIPS/ALUin1[12] ), .B1(n5056), .C0(n8132), .Y(n8204) );
  MXI2X4 U3875 ( .A(n10202), .B(n10201), .S0(n5543), .Y(n10203) );
  AOI222X1 U3876 ( .A0(n4505), .A1(n11466), .B0(mem_rdata_D[90]), .B1(n132), 
        .C0(n12987), .C1(n5535), .Y(n10202) );
  CLKINVX6 U3877 ( .A(n11506), .Y(n11535) );
  OAI222X2 U3878 ( .A0(net107217), .A1(n9217), .B0(n9225), .B1(net117757), 
        .C0(n9206), .C1(n9205), .Y(n9207) );
  BUFX12 U3879 ( .A(n4313), .Y(n3922) );
  INVX12 U3880 ( .A(\i_MIPS/n502 ), .Y(n10334) );
  XNOR2X4 U3881 ( .A(n11367), .B(\i_MIPS/PC/n29 ), .Y(n11602) );
  AO21X4 U3882 ( .A0(n11109), .A1(n11108), .B0(n11107), .Y(n11579) );
  NAND2X1 U3883 ( .A(n11106), .B(n11108), .Y(n9543) );
  OAI22XL U3884 ( .A0(n5261), .A1(n1339), .B0(n5302), .B1(n2994), .Y(n3932) );
  INVX12 U3885 ( .A(n4755), .Y(n5067) );
  CLKINVX6 U3886 ( .A(n8651), .Y(n8652) );
  AO22X1 U3887 ( .A0(net118235), .A1(n770), .B0(net118253), .B1(n2362), .Y(
        n8064) );
  OAI2BB1X4 U3888 ( .A0N(n9181), .A1N(n9180), .B0(n5193), .Y(net106675) );
  NAND2X2 U3889 ( .A(\i_MIPS/ALUin1[12] ), .B(n6692), .Y(n8202) );
  OAI2BB1X2 U3890 ( .A0N(net104698), .A1N(net104699), .B0(n3989), .Y(net109991) );
  OAI2BB1X4 U3891 ( .A0N(net105264), .A1N(net105265), .B0(n3989), .Y(net110955) );
  BUFX16 U3892 ( .A(net117661), .Y(net117653) );
  OA22X2 U3893 ( .A0(n10680), .A1(n3879), .B0(n10683), .B1(n4495), .Y(n7357)
         );
  NAND2X6 U3894 ( .A(n3583), .B(n2920), .Y(n6706) );
  AO21X4 U3895 ( .A0(n6982), .A1(n6981), .B0(n5191), .Y(net105076) );
  OA22X2 U3896 ( .A0(n10963), .A1(n3767), .B0(n10967), .B1(n9536), .Y(n8348)
         );
  MXI2X1 U3897 ( .A(n9296), .B(n8038), .S0(\i_MIPS/ID_EX[81] ), .Y(n4735) );
  INVX8 U3898 ( .A(n11389), .Y(n10805) );
  NAND4X4 U3899 ( .A(n7999), .B(n7998), .C(n7997), .D(n7996), .Y(n11389) );
  OA22X4 U3900 ( .A0(n10653), .A1(n3877), .B0(n10656), .B1(n4495), .Y(n8177)
         );
  OA22X4 U3901 ( .A0(n5652), .A1(n2084), .B0(n5608), .B1(n458), .Y(n11139) );
  OA22X4 U3902 ( .A0(n5652), .A1(n2086), .B0(n5583), .B1(n460), .Y(n11144) );
  AOI2BB1X4 U3903 ( .A0N(n9565), .A1N(n9564), .B0(net107210), .Y(n9571) );
  OAI221XL U3904 ( .A0(net111762), .A1(net117713), .B0(net111763), .B1(
        net117731), .C0(net111764), .Y(n3904) );
  OA22X2 U3905 ( .A0(n10444), .A1(n3767), .B0(n10447), .B1(n9536), .Y(n7123)
         );
  OA22X4 U3906 ( .A0(n5263), .A1(n2087), .B0(n5302), .B1(n461), .Y(n6498) );
  OAI2BB1X4 U3907 ( .A0N(n3776), .A1N(n7429), .B0(n3905), .Y(n3911) );
  OA22X2 U3908 ( .A0(n10462), .A1(n3877), .B0(n10465), .B1(n4495), .Y(n8257)
         );
  INVX8 U3909 ( .A(n11450), .Y(n10774) );
  NAND4X4 U3910 ( .A(n7533), .B(n7532), .C(n7531), .D(n7530), .Y(n11450) );
  OA22X2 U3911 ( .A0(n5395), .A1(n591), .B0(n5438), .B1(n2209), .Y(n7530) );
  OAI221XL U3912 ( .A0(net112118), .A1(net117713), .B0(net112119), .B1(
        net117733), .C0(net112120), .Y(n3907) );
  INVX2 U3913 ( .A(net105290), .Y(net112119) );
  INVX3 U3914 ( .A(n6917), .Y(n6652) );
  NAND2BX4 U3915 ( .AN(n8280), .B(n8556), .Y(n6917) );
  NAND4X4 U3916 ( .A(n9407), .B(n9406), .C(n9405), .D(n9404), .Y(n11502) );
  AOI32X2 U3917 ( .A0(n3024), .A1(\i_MIPS/ID_EX[83] ), .A2(net108632), .B0(
        n8704), .B1(n8705), .Y(n8706) );
  NAND2X2 U3918 ( .A(n5191), .B(n10979), .Y(n11372) );
  OA22X4 U3919 ( .A0(n5259), .A1(n2088), .B0(n5306), .B1(n462), .Y(n6419) );
  INVX6 U3920 ( .A(n6420), .Y(n10997) );
  NAND2XL U3921 ( .A(n10984), .B(n10985), .Y(n11525) );
  MX2X1 U3922 ( .A(n7844), .B(n7843), .S0(\i_MIPS/ID_EX[81] ), .Y(n9444) );
  NAND2BX4 U3923 ( .AN(n8117), .B(n8134), .Y(n7489) );
  INVX4 U3924 ( .A(n9951), .Y(n9944) );
  OAI221X1 U3925 ( .A0(\i_MIPS/Register/register[18][17] ), .A1(net117643), 
        .B0(\i_MIPS/Register/register[26][17] ), .B1(net117661), .C0(n9248), 
        .Y(n9251) );
  OA22X2 U3926 ( .A0(n10204), .A1(n3878), .B0(n10207), .B1(n4495), .Y(n7456)
         );
  OA22X1 U3927 ( .A0(n5333), .A1(n975), .B0(n5358), .B1(n2600), .Y(n9174) );
  OA21X4 U3928 ( .A0(n344), .A1(n5067), .B0(n7587), .Y(n7153) );
  INVX1 U3929 ( .A(n7490), .Y(n7491) );
  OA22X4 U3930 ( .A0(n10580), .A1(n10579), .B0(n10582), .B1(n10722), .Y(n10585) );
  NAND3X8 U3931 ( .A(n3913), .B(n3914), .C(net111423), .Y(net105746) );
  AO21X4 U3932 ( .A0(net105751), .A1(net105752), .B0(net117723), .Y(net111423)
         );
  OR2X6 U3933 ( .A(net111422), .B(net117731), .Y(n3914) );
  NAND2X4 U3934 ( .A(\i_MIPS/ALUin1[17] ), .B(n6699), .Y(n9217) );
  NAND2X2 U3935 ( .A(net109511), .B(n142), .Y(n8282) );
  NAND3BX4 U3936 ( .AN(net112449), .B(net109176), .C(net109179), .Y(net109512)
         );
  AO21X4 U3937 ( .A0(net108310), .A1(n7784), .B0(n7159), .Y(n8560) );
  BUFX8 U3938 ( .A(n7303), .Y(n3909) );
  NAND4X4 U3939 ( .A(n7529), .B(n7528), .C(n7527), .D(n7526), .Y(n11482) );
  NAND2X6 U3940 ( .A(n10997), .B(n10996), .Y(n6423) );
  CLKAND2X2 U3941 ( .A(net104171), .B(n11233), .Y(n4437) );
  OAI221X4 U3942 ( .A0(n7851), .A1(n9550), .B0(n7850), .B1(n9553), .C0(n7849), 
        .Y(n7852) );
  AOI2BB1X1 U3943 ( .A0N(n9552), .A1N(n7840), .B0(net107841), .Y(n7855) );
  INVX12 U3944 ( .A(net107389), .Y(net107841) );
  NAND4X4 U3945 ( .A(n8172), .B(n8171), .C(n8170), .D(n8169), .Y(n11384) );
  OA22X2 U3946 ( .A0(n10456), .A1(n3766), .B0(n10459), .B1(n9536), .Y(n8258)
         );
  OA22X2 U3947 ( .A0(n10799), .A1(n3766), .B0(n10802), .B1(n9536), .Y(n8005)
         );
  OA22X4 U3948 ( .A0(n10647), .A1(n3766), .B0(n10650), .B1(n9536), .Y(n8178)
         );
  CLKBUFX20 U3949 ( .A(net107607), .Y(net118227) );
  OA22X4 U3950 ( .A0(n5254), .A1(n2090), .B0(n5294), .B1(n464), .Y(n9532) );
  NAND4X4 U3951 ( .A(n9533), .B(n9532), .C(n9531), .D(n9530), .Y(n11439) );
  OA22X2 U3952 ( .A0(n5392), .A1(n593), .B0(n5435), .B1(n2211), .Y(n9530) );
  OAI211X2 U3953 ( .A0(n9319), .A1(n9300), .B0(n7488), .C0(n9309), .Y(n7303)
         );
  OA22X4 U3954 ( .A0(n7401), .A1(n11103), .B0(n7400), .B1(n7404), .Y(n7438) );
  NAND2X2 U3955 ( .A(n6664), .B(n3674), .Y(n8133) );
  AOI222X2 U3956 ( .A0(n4534), .A1(n11498), .B0(mem_rdata_D[122]), .B1(n130), 
        .C0(n12987), .C1(n5533), .Y(n10199) );
  BUFX20 U3957 ( .A(n4685), .Y(n5533) );
  AO22X4 U3958 ( .A0(net109168), .A1(n4653), .B0(net109965), .B1(n7483), .Y(
        n7485) );
  OAI222X1 U3959 ( .A0(n7850), .A1(net107688), .B0(net107217), .B1(n3868), 
        .C0(net107689), .C1(n7221), .Y(n7239) );
  OAI221X4 U3960 ( .A0(\i_MIPS/ALUin1[11] ), .A1(n5064), .B0(
        \i_MIPS/ALUin1[10] ), .B1(n5057), .C0(n7156), .Y(n7221) );
  NOR4BX4 U3961 ( .AN(n7855), .B(n7854), .C(n7853), .D(n7852), .Y(n7874) );
  OAI221X2 U3962 ( .A0(net118601), .A1(n8873), .B0(net108781), .B1(n8975), 
        .C0(n6933), .Y(n7943) );
  AO21X4 U3963 ( .A0(n7056), .A1(n7055), .B0(n7054), .Y(n3912) );
  NAND2XL U3964 ( .A(n7027), .B(n7863), .Y(n7055) );
  OR2X2 U3965 ( .A(net111421), .B(net117711), .Y(n3913) );
  MX2X1 U3966 ( .A(n7220), .B(n7219), .S0(\i_MIPS/jump_addr[22] ), .Y(
        net111421) );
  INVX12 U3967 ( .A(net117719), .Y(net117711) );
  OR3X6 U3968 ( .A(n6695), .B(net112449), .C(n3744), .Y(n4624) );
  CLKINVX4 U3969 ( .A(n7301), .Y(n8657) );
  NAND2X4 U3970 ( .A(net105731), .B(net105732), .Y(n4359) );
  INVX3 U3971 ( .A(n134), .Y(n6939) );
  NAND2XL U3972 ( .A(net139849), .B(net105105), .Y(n10554) );
  AOI211X4 U3973 ( .A0(n3777), .A1(n8137), .B0(n8136), .C0(n8135), .Y(n8138)
         );
  NAND4X4 U3974 ( .A(n7121), .B(n7120), .C(n7119), .D(n7118), .Y(n11423) );
  OA22X2 U3975 ( .A0(n5397), .A1(n594), .B0(n5441), .B1(n2212), .Y(n7118) );
  OAI221X4 U3976 ( .A0(net111580), .A1(net117713), .B0(net111581), .B1(
        net117731), .C0(net111582), .Y(net105250) );
  MX2X1 U3977 ( .A(n7143), .B(n7142), .S0(net114081), .Y(net111580) );
  OA22X2 U3978 ( .A0(n10612), .A1(n3879), .B0(n10615), .B1(n4495), .Y(n8087)
         );
  OA22X2 U3979 ( .A0(n10606), .A1(n3767), .B0(n10609), .B1(n9536), .Y(n8088)
         );
  INVX2 U3980 ( .A(net105313), .Y(net112329) );
  NAND2X8 U3981 ( .A(n3026), .B(n9301), .Y(n7768) );
  AND4X8 U3982 ( .A(n3915), .B(n3916), .C(n3917), .D(n3918), .Y(n4317) );
  NAND4X8 U3983 ( .A(n3919), .B(n3920), .C(n6515), .D(n6514), .Y(n9599) );
  AOI222X1 U3984 ( .A0(n4534), .A1(n11502), .B0(mem_rdata_D[126]), .B1(n132), 
        .C0(n12983), .C1(n5534), .Y(n10593) );
  OAI2BB1X2 U3985 ( .A0N(net106037), .A1N(net106038), .B0(net117631), .Y(
        net106301) );
  NAND2X2 U3986 ( .A(n9950), .B(n10979), .Y(n11505) );
  OR2X8 U3987 ( .A(n5191), .B(n9796), .Y(n9950) );
  CLKINVX12 U3988 ( .A(n11590), .Y(n6528) );
  NAND4X4 U3989 ( .A(n11135), .B(n11134), .C(n11133), .D(n11132), .Y(n11591)
         );
  XNOR2X4 U3990 ( .A(ICACHE_addr[15]), .B(n11357), .Y(n11133) );
  CLKBUFX3 U3991 ( .A(n5408), .Y(n5405) );
  NAND4X4 U3992 ( .A(n9411), .B(n9410), .C(n9409), .D(n9408), .Y(n11470) );
  AO21XL U3993 ( .A0(\i_MIPS/ALUin1[0] ), .A1(n3852), .B0(net108308), .Y(n8705) );
  OAI221X2 U3994 ( .A0(n5329), .A1(n2953), .B0(n5354), .B1(n1312), .C0(n6510), 
        .Y(n6511) );
  OA22X4 U3995 ( .A0(n5262), .A1(n2092), .B0(n5302), .B1(n466), .Y(n6504) );
  OA22X2 U3996 ( .A0(n10555), .A1(n3767), .B0(n10558), .B1(n9536), .Y(n6982)
         );
  BUFX20 U3997 ( .A(net107218), .Y(net118592) );
  OAI221X2 U3998 ( .A0(net118601), .A1(n9049), .B0(n8699), .B1(n3745), .C0(
        n7419), .Y(n8111) );
  OA22X2 U3999 ( .A0(n9953), .A1(n3878), .B0(n9960), .B1(n4495), .Y(n7277) );
  INVX8 U4000 ( .A(n11414), .Y(n9960) );
  NAND4X4 U4001 ( .A(n7276), .B(n7275), .C(n7274), .D(n7273), .Y(n11414) );
  XOR2X4 U4002 ( .A(n6462), .B(n4365), .Y(n4003) );
  XOR2X4 U4003 ( .A(n6481), .B(n2997), .Y(n4095) );
  AOI22X4 U4004 ( .A0(n5236), .A1(\D_cache/cache[2][36] ), .B0(n3924), .B1(
        \D_cache/cache[3][36] ), .Y(n9086) );
  BUFX3 U4005 ( .A(n5307), .Y(n5286) );
  AO22X4 U4006 ( .A0(n4703), .A1(net117747), .B0(net135551), .B1(n9125), .Y(
        n9129) );
  NAND2X4 U4007 ( .A(n3628), .B(n8279), .Y(n6916) );
  AOI2BB2X4 U4008 ( .B0(n3924), .B1(\D_cache/cache[3][145] ), .A0N(n5258), 
        .A1N(n2960), .Y(n6508) );
  NAND3BX2 U4009 ( .AN(n11102), .B(n7403), .C(n7402), .Y(n7437) );
  NAND4X4 U4010 ( .A(n7622), .B(n7621), .C(n7620), .D(n7619), .Y(n11404) );
  XNOR2X4 U4011 ( .A(n6430), .B(n12974), .Y(n3927) );
  XNOR2X4 U4012 ( .A(n6443), .B(DCACHE_addr[12]), .Y(n3928) );
  NAND2X2 U4013 ( .A(n4773), .B(n3894), .Y(n4640) );
  AND2X8 U4014 ( .A(net115799), .B(net134815), .Y(net135522) );
  OA22X2 U4015 ( .A0(n5786), .A1(n4680), .B0(n5831), .B1(n2936), .Y(n11129) );
  AOI22X4 U4016 ( .A0(\i_MIPS/IF_ID[25] ), .A1(n6016), .B0(n10375), .B1(n10374), .Y(n4808) );
  NAND3BX4 U4017 ( .AN(n4820), .B(n4805), .C(n10373), .Y(n10374) );
  OA22X4 U4018 ( .A0(n9441), .A1(net107210), .B0(n3774), .B1(n9540), .Y(n9464)
         );
  NAND4X8 U4019 ( .A(n6674), .B(n6673), .C(net108787), .D(n8634), .Y(n9549) );
  NOR3X8 U4020 ( .A(n3930), .B(n3966), .C(n3860), .Y(n3929) );
  BUFX4 U4021 ( .A(n3965), .Y(n5053) );
  BUFX20 U4022 ( .A(n5884), .Y(n5877) );
  AOI2BB1X4 U4023 ( .A0N(n2928), .A1N(n5059), .B0(n4799), .Y(n7037) );
  OAI221X1 U4024 ( .A0(net118601), .A1(net110602), .B0(net107992), .B1(
        net108781), .C0(net111710), .Y(net107230) );
  OAI211X4 U4025 ( .A0(n3854), .A1(n9299), .B0(net110932), .C0(n7301), .Y(
        n8122) );
  OR2X6 U4026 ( .A(n5354), .B(n2352), .Y(n4628) );
  NAND4X2 U4027 ( .A(n1340), .B(n4000), .C(net134414), .D(n4021), .Y(net112544) );
  AOI222X2 U4028 ( .A0(n4707), .A1(n7790), .B0(n7229), .B1(n7228), .C0(n7227), 
        .C1(n7226), .Y(n7238) );
  OA22X4 U4029 ( .A0(n5256), .A1(n2094), .B0(n5299), .B1(n468), .Y(n7267) );
  OA22X4 U4030 ( .A0(n5239), .A1(n2097), .B0(n5299), .B1(n471), .Y(n7195) );
  OA22X4 U4031 ( .A0(n5239), .A1(n2098), .B0(n5299), .B1(n472), .Y(n7199) );
  AOI2BB1X4 U4032 ( .A0N(n3854), .A1N(n8661), .B0(n8660), .Y(n8667) );
  OA22X4 U4033 ( .A0(n138), .A1(n2099), .B0(n5696), .B1(n473), .Y(n11190) );
  NAND2X8 U4034 ( .A(n7845), .B(n9549), .Y(net108632) );
  INVX3 U4035 ( .A(n8210), .Y(n7945) );
  OAI2BB1X4 U4036 ( .A0N(net104917), .A1N(net104916), .B0(n3989), .Y(net108162) );
  OAI222X2 U4037 ( .A0(n8379), .A1(n8699), .B0(net118601), .B1(n8386), .C0(
        n3674), .C1(n9055), .Y(n8205) );
  AND2XL U4038 ( .A(net139850), .B(net104791), .Y(n4695) );
  OR2X4 U4039 ( .A(net108490), .B(net117709), .Y(n3933) );
  OR2X6 U4040 ( .A(net108491), .B(net117731), .Y(n3934) );
  NAND3X6 U4041 ( .A(n3933), .B(n3934), .C(net108492), .Y(net105160) );
  XOR2X4 U4042 ( .A(n4364), .B(net105160), .Y(n4324) );
  OA22X4 U4043 ( .A0(n5832), .A1(n2100), .B0(n5785), .B1(n474), .Y(n11184) );
  OR2X4 U4044 ( .A(n8960), .B(net117709), .Y(n3935) );
  NAND3X6 U4045 ( .A(n3935), .B(n3936), .C(n8958), .Y(net105137) );
  OA22X4 U4046 ( .A0(n5920), .A1(n1297), .B0(n5878), .B1(n2963), .Y(n11198) );
  AO22X4 U4047 ( .A0(mem_rdata_I[37]), .A1(n5943), .B0(n5567), .B1(n11255), 
        .Y(n9710) );
  OAI21X2 U4048 ( .A0(n11217), .A1(n6528), .B0(n11218), .Y(n6529) );
  AND2X8 U4049 ( .A(net139865), .B(net105517), .Y(n4060) );
  NAND2XL U4050 ( .A(net139865), .B(net105517), .Y(n10978) );
  AO21X4 U4051 ( .A0(net105662), .A1(net105663), .B0(net117625), .Y(net105517)
         );
  CLKINVX12 U4052 ( .A(n11059), .Y(n5559) );
  OA22X4 U4053 ( .A0(n5259), .A1(n2101), .B0(n5301), .B1(n475), .Y(n6448) );
  INVX20 U4054 ( .A(net134710), .Y(net107217) );
  OAI222X1 U4055 ( .A0(n9043), .A1(net107688), .B0(net107217), .B1(n9300), 
        .C0(net107689), .C1(n9042), .Y(n9058) );
  CLKAND2X12 U4056 ( .A(n8634), .B(n8632), .Y(n4741) );
  AND2X4 U4057 ( .A(n8178), .B(n8177), .Y(n3937) );
  OAI31X2 U4058 ( .A0(n6925), .A1(n6924), .A2(n6923), .B0(n6922), .Y(n3938) );
  OR2X1 U4059 ( .A(n10304), .B(n5561), .Y(n3939) );
  OR2X1 U4060 ( .A(n5558), .B(n10305), .Y(n3940) );
  NAND2X6 U4061 ( .A(\i_MIPS/ALUin1[28] ), .B(n6955), .Y(n9425) );
  NAND2X8 U4062 ( .A(ICACHE_addr[1]), .B(ICACHE_addr[0]), .Y(n9802) );
  NAND2X2 U4063 ( .A(n10715), .B(ICACHE_addr[28]), .Y(n10716) );
  OAI211X2 U4064 ( .A0(net106828), .A1(net104828), .B0(net135522), .C0(n9607), 
        .Y(net107120) );
  INVX1 U4065 ( .A(n3941), .Y(n3942) );
  AND2XL U4066 ( .A(n5044), .B(n11424), .Y(n12854) );
  NAND4X2 U4067 ( .A(n7451), .B(n7450), .C(n7449), .D(n7448), .Y(n11402) );
  OA22XL U4068 ( .A0(n5180), .A1(n1080), .B0(n5218), .B1(n2703), .Y(n7451) );
  OAI221XL U4069 ( .A0(net109201), .A1(net117709), .B0(net109202), .B1(
        net117731), .C0(net109203), .Y(n3944) );
  OAI221X2 U4070 ( .A0(net109201), .A1(net117709), .B0(net109202), .B1(
        net117731), .C0(net109203), .Y(net105329) );
  OAI2BB1X2 U4071 ( .A0N(net105490), .A1N(net105491), .B0(n3989), .Y(net105434) );
  INVX1 U4072 ( .A(n8881), .Y(n7859) );
  NAND2X6 U4073 ( .A(n4620), .B(n4712), .Y(n8881) );
  NAND4X4 U4074 ( .A(DCACHE_ren), .B(\i_MIPS/EX_MEM_1 ), .C(n9944), .D(n11374), 
        .Y(n9537) );
  NAND4X4 U4075 ( .A(n7626), .B(n7625), .C(n7624), .D(n7623), .Y(n11436) );
  OA22X2 U4076 ( .A0(n5394), .A1(n595), .B0(n5437), .B1(n2213), .Y(n7623) );
  CLKBUFX4 U4077 ( .A(n5449), .Y(n5437) );
  MXI2X2 U4078 ( .A(n9254), .B(n9253), .S0(net114085), .Y(n3948) );
  NAND2X2 U4079 ( .A(n3950), .B(n6946), .Y(n6964) );
  OAI211X2 U4080 ( .A0(n4729), .A1(n6721), .B0(n4687), .C0(n8683), .Y(n6818)
         );
  NAND2X8 U4081 ( .A(n4710), .B(n8681), .Y(n6721) );
  NAND2X8 U4082 ( .A(n6700), .B(n1264), .Y(n8681) );
  INVX12 U4083 ( .A(n4503), .Y(n6700) );
  OAI2BB1X2 U4084 ( .A0N(net105232), .A1N(net105233), .B0(net117631), .Y(
        net105756) );
  AO22X4 U4085 ( .A0(n4702), .A1(net117747), .B0(n3950), .B1(n8123), .Y(n8126)
         );
  NAND4X8 U4086 ( .A(n6710), .B(n8648), .C(n7492), .D(n8666), .Y(net112219) );
  NAND2X2 U4087 ( .A(\i_MIPS/ALUin1[10] ), .B(n3760), .Y(n8648) );
  INVX8 U4088 ( .A(n11406), .Y(n10598) );
  NAND4X4 U4089 ( .A(n9415), .B(n9414), .C(n9413), .D(n9412), .Y(n11406) );
  OAI2BB1XL U4090 ( .A0N(net106675), .A1N(net106674), .B0(n3989), .Y(n3949) );
  OAI2BB1X4 U4091 ( .A0N(n7101), .A1N(n7768), .B0(n3951), .Y(n6915) );
  OAI22X4 U4092 ( .A0(n11579), .A1(n11573), .B0(n4728), .B1(n11579), .Y(n11580) );
  OAI2BB1X4 U4093 ( .A0N(n7542), .A1N(n7541), .B0(n4407), .Y(net105120) );
  AOI21X2 U4094 ( .A0(n8758), .A1(n8757), .B0(n4626), .Y(n3952) );
  OAI2BB1X4 U4095 ( .A0N(n4706), .A1N(n8881), .B0(n8300), .Y(n8383) );
  INVX2 U4096 ( .A(n8300), .Y(n8380) );
  OAI31X2 U4097 ( .A0(n7859), .A1(n8864), .A2(n7858), .B0(n7857), .Y(n7869) );
  AO21X4 U4098 ( .A0(n8889), .A1(n8859), .B0(n8690), .Y(n7025) );
  INVX4 U4099 ( .A(n8860), .Y(n8690) );
  AO21X4 U4100 ( .A0(n6871), .A1(n6870), .B0(n5192), .Y(n3953) );
  BUFX2 U4101 ( .A(n5453), .Y(n5442) );
  NAND4X4 U4102 ( .A(n6976), .B(n6975), .C(n6974), .D(n6973), .Y(n11405) );
  OAI211X4 U4103 ( .A0(n6930), .A1(n3617), .B0(n6929), .C0(net107389), .Y(
        n6945) );
  OA21X4 U4104 ( .A0(n1263), .A1(n5064), .B0(n7953), .Y(n6840) );
  OAI2BB1X2 U4105 ( .A0N(net105662), .A1N(net105663), .B0(n3989), .Y(net109360) );
  NAND2X6 U4106 ( .A(n4636), .B(n4637), .Y(net105335) );
  NAND2XL U4107 ( .A(net139866), .B(net105567), .Y(n10511) );
  INVX1 U4108 ( .A(n10498), .Y(n5491) );
  NAND3BX2 U4109 ( .AN(n11505), .B(n11539), .C(n11504), .Y(n11508) );
  INVX1 U4110 ( .A(n11505), .Y(n10980) );
  NAND2X2 U4111 ( .A(n11505), .B(n3634), .Y(net140147) );
  AOI221X2 U4112 ( .A0(net119020), .A1(net117715), .B0(net105425), .B1(
        net117741), .C0(net119021), .Y(net119018) );
  INVX1 U4113 ( .A(n3954), .Y(n3955) );
  AOI222X2 U4114 ( .A0(n4688), .A1(n8975), .B0(n6931), .B1(n8976), .C0(n7676), 
        .C1(n8043), .Y(n6835) );
  INVXL U4115 ( .A(n7838), .Y(n3956) );
  NAND4X4 U4116 ( .A(n7455), .B(n7454), .C(n7453), .D(n7452), .Y(n11434) );
  AOI221X2 U4117 ( .A0(net117743), .A1(net109666), .B0(n8201), .B1(n3950), 
        .C0(net134673), .Y(n8218) );
  OAI2BB1X4 U4118 ( .A0N(net106603), .A1N(net106602), .B0(n3989), .Y(n9118) );
  INVXL U4119 ( .A(net106603), .Y(n3957) );
  INVX1 U4120 ( .A(n3957), .Y(n3958) );
  AOI2BB1X4 U4121 ( .A0N(n959), .A1N(n5059), .B0(n4818), .Y(n8110) );
  OR2X8 U4122 ( .A(net109359), .B(net117731), .Y(net143556) );
  CLKMX2X2 U4123 ( .A(n12966), .B(n3761), .S0(n3593), .Y(\i_MIPS/n380 ) );
  AOI211X2 U4124 ( .A0(n8680), .A1(n4693), .B0(n8376), .C0(n8375), .Y(n8392)
         );
  OAI221X2 U4125 ( .A0(net107210), .A1(n9125), .B0(n4703), .B1(n3774), .C0(
        net117759), .Y(n9130) );
  OR2X6 U4126 ( .A(net109990), .B(net117731), .Y(n3961) );
  CLKMX2X2 U4127 ( .A(n3543), .B(net104691), .S0(n3591), .Y(\i_MIPS/n341 ) );
  AO21X4 U4128 ( .A0(net105311), .A1(net105312), .B0(net117623), .Y(net105396)
         );
  AO21X4 U4129 ( .A0(net105490), .A1(net105491), .B0(net117625), .Y(net105449)
         );
  OR2X6 U4130 ( .A(n7838), .B(net117731), .Y(n3963) );
  OAI32X2 U4131 ( .A0(n8479), .A1(n8478), .A2(net107210), .B0(n4762), .B1(
        net107688), .Y(n8484) );
  AND3X2 U4132 ( .A(n3950), .B(n8486), .C(n3645), .Y(n8473) );
  AOI222X1 U4133 ( .A0(n4534), .A1(n11481), .B0(mem_rdata_D[105]), .B1(n132), 
        .C0(n13004), .C1(n5534), .Y(n10607) );
  OAI221X4 U4134 ( .A0(\i_MIPS/ALUin1[20] ), .A1(n5072), .B0(
        \i_MIPS/ALUin1[21] ), .B1(n5068), .C0(n7032), .Y(n7671) );
  AO21X4 U4135 ( .A0(n9945), .A1(n9944), .B0(n9943), .Y(n10966) );
  AO22X4 U4136 ( .A0(n5945), .A1(ICACHE_addr[21]), .B0(n5931), .B1(n11363), 
        .Y(n11145) );
  OA22X4 U4137 ( .A0(n5652), .A1(n2104), .B0(n5608), .B1(n478), .Y(n11126) );
  BUFX20 U4138 ( .A(n5930), .Y(n5931) );
  OAI211X2 U4139 ( .A0(net106828), .A1(net104828), .B0(n4314), .C0(net135522), 
        .Y(n4313) );
  OAI222X2 U4140 ( .A0(n9576), .A1(net117709), .B0(n4982), .B1(net117723), 
        .C0(n9597), .C1(net117731), .Y(n10735) );
  AND3X4 U4141 ( .A(n3950), .B(n7048), .C(n7047), .Y(n7049) );
  OA22X4 U4142 ( .A0(n5259), .A1(n2105), .B0(n5307), .B1(n479), .Y(n6451) );
  INVX12 U4143 ( .A(\i_MIPS/n503 ), .Y(net105477) );
  OAI221X4 U4144 ( .A0(\i_MIPS/ALUin1[12] ), .A1(n5071), .B0(
        \i_MIPS/ALUin1[11] ), .B1(n5068), .C0(n8036), .Y(n9296) );
  AOI222X2 U4145 ( .A0(n9122), .A1(net118584), .B0(n7149), .B1(n7148), .C0(
        n7147), .C1(n7146), .Y(n7150) );
  OAI221X2 U4146 ( .A0(n5328), .A1(n2015), .B0(n5353), .B1(n396), .C0(n6479), 
        .Y(n6480) );
  OA22X4 U4147 ( .A0(n5402), .A1(n2106), .B0(n5445), .B1(n480), .Y(n6479) );
  CLKINVX20 U4148 ( .A(net135551), .Y(net107210) );
  OAI222X2 U4149 ( .A0(n9202), .A1(n9052), .B0(n9043), .B1(n9553), .C0(n8374), 
        .C1(n5049), .Y(n8375) );
  OAI2BB1X4 U4150 ( .A0N(n3985), .A1N(n8211), .B0(n8199), .Y(n7962) );
  AOI2BB1X1 U4151 ( .A0N(n9200), .A1N(n5049), .B0(n8045), .Y(n8046) );
  NOR2X6 U4152 ( .A(n4398), .B(n8483), .Y(n8489) );
  NAND4X8 U4153 ( .A(n6673), .B(n6674), .C(n8634), .D(net112393), .Y(n7845) );
  NAND2X1 U4154 ( .A(\i_MIPS/IF_ID[3] ), .B(\i_MIPS/Sign_Extend[1] ), .Y(
        n10905) );
  AOI32X2 U4155 ( .A0(n10906), .A1(n10904), .A2(n10905), .B0(\i_MIPS/n518 ), 
        .B1(\i_MIPS/n158 ), .Y(n10135) );
  AND2X8 U4156 ( .A(n9223), .B(n9203), .Y(n4710) );
  NAND2X8 U4157 ( .A(n6698), .B(n959), .Y(n9223) );
  AND2XL U4158 ( .A(n6691), .B(n300), .Y(n3968) );
  OA22X4 U4159 ( .A0(n5920), .A1(n3010), .B0(n5878), .B1(n1341), .Y(n11203) );
  BUFX20 U4160 ( .A(net134445), .Y(net117631) );
  AOI222X2 U4161 ( .A0(n4715), .A1(n8208), .B0(n8207), .B1(net107404), .C0(
        n8206), .C1(net109661), .Y(n8209) );
  CLKINVX12 U4162 ( .A(n3016), .Y(n4545) );
  CLKINVX12 U4163 ( .A(n3016), .Y(n4544) );
  OAI222X4 U4164 ( .A0(n8790), .A1(n8793), .B0(n9547), .B1(n7600), .C0(n9202), 
        .C1(n8111), .Y(n6680) );
  AO22X1 U4165 ( .A0(n5555), .A1(net105236), .B0(n11054), .B1(
        \i_MIPS/Sign_Extend[13] ), .Y(n10266) );
  XOR2X4 U4166 ( .A(n11363), .B(ICACHE_addr[21]), .Y(n11593) );
  NAND4X4 U4167 ( .A(n11144), .B(n11143), .C(n11142), .D(n11141), .Y(n11363)
         );
  BUFX20 U4168 ( .A(n4684), .Y(n5537) );
  AOI222X4 U4169 ( .A0(n5541), .A1(n11434), .B0(mem_rdata_D[58]), .B1(n133), 
        .C0(n12987), .C1(n5539), .Y(n10208) );
  AO21X4 U4170 ( .A0(net104792), .A1(n4015), .B0(net117623), .Y(net104791) );
  OAI211X4 U4171 ( .A0(n3764), .A1(net110131), .B0(net110406), .C0(net109519), 
        .Y(net108622) );
  NAND3BX2 U4172 ( .AN(n4764), .B(n8788), .C(n3950), .Y(n8796) );
  BUFX6 U4173 ( .A(n6950), .Y(n3973) );
  AOI222X1 U4174 ( .A0(n4534), .A1(n11487), .B0(mem_rdata_D[111]), .B1(n133), 
        .C0(n12998), .C1(n5533), .Y(n10445) );
  MXI2XL U4175 ( .A(\i_MIPS/n190 ), .B(n3947), .S0(n3591), .Y(\i_MIPS/n313 )
         );
  NAND2XL U4176 ( .A(net139774), .B(net106819), .Y(n10768) );
  AO21X4 U4177 ( .A0(net106675), .A1(net106674), .B0(net117623), .Y(net106819)
         );
  NAND4X4 U4178 ( .A(n11139), .B(n11138), .C(n11137), .D(n11136), .Y(n11358)
         );
  AO21X4 U4179 ( .A0(n9604), .A1(n3634), .B0(n11584), .Y(n11085) );
  OAI211X2 U4180 ( .A0(n7026), .A1(n6817), .B0(n11101), .C0(n6816), .Y(n6953)
         );
  OAI211X2 U4181 ( .A0(n4273), .A1(net108149), .B0(net112413), .C0(net107680), 
        .Y(net111270) );
  NAND3BX2 U4182 ( .AN(n6849), .B(n6848), .C(n4701), .Y(n6850) );
  OAI222X2 U4183 ( .A0(n8561), .A1(n9550), .B0(n9202), .B1(n8560), .C0(n8559), 
        .C1(n5049), .Y(n8562) );
  OAI2BB1X4 U4184 ( .A0N(n9097), .A1N(n9096), .B0(n5193), .Y(net106603) );
  AOI222X1 U4185 ( .A0(n4534), .A1(n11501), .B0(mem_rdata_D[125]), .B1(n129), 
        .C0(n12984), .C1(n5534), .Y(n10556) );
  BUFX6 U4186 ( .A(n9422), .Y(n3977) );
  NAND3BX4 U4187 ( .AN(n8680), .B(n4698), .C(n8395), .Y(n8399) );
  OAI221X2 U4188 ( .A0(n9868), .A1(net143858), .B0(\i_MIPS/n513 ), .B1(
        net115791), .C0(n9867), .Y(\i_MIPS/N57 ) );
  OA22X2 U4189 ( .A0(n5920), .A1(n598), .B0(n5878), .B1(n2216), .Y(n11188) );
  INVXL U4190 ( .A(n3702), .Y(n3978) );
  NOR2BX4 U4191 ( .AN(\i_MIPS/jump_addr[23] ), .B(\i_MIPS/n499 ), .Y(n4814) );
  OA22X4 U4192 ( .A0(n5261), .A1(n2108), .B0(n5303), .B1(n482), .Y(n6409) );
  NAND4X4 U4193 ( .A(n9091), .B(n9090), .C(n9089), .D(n9088), .Y(n11380) );
  CLKINVX2 U4194 ( .A(net104765), .Y(net111422) );
  OAI221X2 U4195 ( .A0(n5324), .A1(n2016), .B0(n5363), .B1(n397), .C0(n6396), 
        .Y(n6397) );
  INVXL U4196 ( .A(net109528), .Y(n3980) );
  AOI2BB2X4 U4197 ( .B0(net104700), .B1(net118217), .A0N(n3890), .A1N(n3981), 
        .Y(net139860) );
  XOR2X4 U4198 ( .A(n11364), .B(ICACHE_addr[22]), .Y(n6382) );
  XOR2X4 U4199 ( .A(n11370), .B(ICACHE_addr[28]), .Y(n6383) );
  NAND4X4 U4200 ( .A(n9144), .B(n9143), .C(n9142), .D(n9141), .Y(net104367) );
  AOI222X2 U4201 ( .A0(n4623), .A1(net118584), .B0(n9131), .B1(n9130), .C0(
        n9129), .C1(n9128), .Y(n9144) );
  AOI222X4 U4202 ( .A0(n5541), .A1(n11433), .B0(mem_rdata_D[57]), .B1(n132), 
        .C0(n12988), .C1(n5539), .Y(n10441) );
  NAND4X4 U4203 ( .A(n9419), .B(n9418), .C(n9417), .D(n9416), .Y(n11438) );
  OA22X1 U4204 ( .A0(n5333), .A1(n976), .B0(n5358), .B1(n2601), .Y(n9417) );
  CLKAND2X8 U4205 ( .A(n5070), .B(\i_MIPS/ALUin1[27] ), .Y(n4793) );
  AO22X4 U4206 ( .A0(net118215), .A1(n10512), .B0(net118225), .B1(n8919), .Y(
        net108412) );
  CLKMX2X2 U4207 ( .A(DCACHE_addr[5]), .B(net104891), .S0(n3603), .Y(
        \i_MIPS/n392 ) );
  AO22X4 U4208 ( .A0(net118217), .A1(net104891), .B0(net118227), .B1(n7340), 
        .Y(net111216) );
  NAND3BX4 U4209 ( .AN(n7319), .B(n7318), .C(n7317), .Y(net104891) );
  AND2X2 U4210 ( .A(n6770), .B(n348), .Y(net134686) );
  OA22X4 U4211 ( .A0(n9316), .A1(n9132), .B0(net107991), .B1(n3617), .Y(n9143)
         );
  INVXL U4212 ( .A(net109990), .Y(n3982) );
  AOI33X2 U4213 ( .A0(n3950), .A1(n9231), .A2(n9230), .B0(n9229), .B1(n9228), 
        .B2(net117743), .Y(n9232) );
  OAI2BB1X4 U4214 ( .A0N(n8783), .A1N(n9216), .B0(n9217), .Y(n8280) );
  NAND2X8 U4215 ( .A(n2996), .B(n4643), .Y(net109519) );
  MX2X1 U4216 ( .A(n12974), .B(n3978), .S0(n3605), .Y(\i_MIPS/n388 ) );
  MX2X1 U4217 ( .A(DCACHE_addr[11]), .B(n3982), .S0(n3588), .Y(\i_MIPS/n386 )
         );
  AOI222X1 U4218 ( .A0(n3800), .A1(n11397), .B0(mem_rdata_D[21]), .B1(n130), 
        .C0(n12992), .C1(n5538), .Y(n10521) );
  NAND4X2 U4219 ( .A(n7113), .B(n7112), .C(n7111), .D(n7110), .Y(n11455) );
  OAI33X2 U4220 ( .A0(n7778), .A1(n351), .A2(net107210), .B0(n3774), .B1(n351), 
        .B2(n7780), .Y(n7796) );
  AOI211X4 U4221 ( .A0(n4696), .A1(n8208), .B0(n7792), .C0(n7791), .Y(n7793)
         );
  AOI33X2 U4222 ( .A0(n3950), .A1(n8385), .A2(n8384), .B0(n3950), .B1(n8393), 
        .B2(n8383), .Y(n8390) );
  OA22X4 U4223 ( .A0(net107217), .A1(n8300), .B0(n8309), .B1(net117759), .Y(
        n8301) );
  INVX20 U4224 ( .A(net134673), .Y(net117759) );
  AND3X2 U4225 ( .A(\i_MIPS/ID_EX[78] ), .B(n11), .C(n3873), .Y(n4834) );
  AOI222X2 U4226 ( .A0(n4707), .A1(n9314), .B0(n9313), .B1(n9312), .C0(n9311), 
        .C1(n9310), .Y(n9324) );
  INVX1 U4227 ( .A(n8041), .Y(n8042) );
  OA22X4 U4228 ( .A0(n138), .A1(n2111), .B0(n5694), .B1(n485), .Y(n11125) );
  NAND3BX1 U4229 ( .AN(n8487), .B(n4753), .C(net117745), .Y(n8488) );
  NAND2X8 U4230 ( .A(n6690), .B(n1263), .Y(net108874) );
  OAI221X2 U4231 ( .A0(n5169), .A1(n2017), .B0(n5209), .B1(n398), .C0(n6394), 
        .Y(n6395) );
  CLKMX2X4 U4232 ( .A(n7842), .B(n7786), .S0(net114065), .Y(n8558) );
  OAI221X4 U4233 ( .A0(n3744), .A1(n5071), .B0(n1263), .B1(n5068), .C0(n7418), 
        .Y(n7786) );
  NAND2BX4 U4234 ( .AN(n8663), .B(n6706), .Y(n7492) );
  NAND4BX2 U4235 ( .AN(n4646), .B(n7540), .C(n7539), .D(n7538), .Y(n11418) );
  OA22XL U4236 ( .A0(n5256), .A1(n1081), .B0(n5296), .B1(n2704), .Y(n7540) );
  MX2XL U4237 ( .A(n12963), .B(net105492), .S0(n3605), .Y(\i_MIPS/n377 ) );
  AO21X4 U4238 ( .A0(n8485), .A1(net107992), .B0(n8484), .Y(n4398) );
  OAI2BB1X4 U4239 ( .A0N(n7486), .A1N(n7303), .B0(n3868), .Y(n7305) );
  INVX8 U4240 ( .A(n11437), .Y(n10564) );
  AOI222X4 U4241 ( .A0(n5541), .A1(n11437), .B0(mem_rdata_D[61]), .B1(n129), 
        .C0(n12984), .C1(n5539), .Y(n10565) );
  NAND4X4 U4242 ( .A(n6980), .B(n6979), .C(n6978), .D(n6977), .Y(n11437) );
  OA22X2 U4243 ( .A0(n5398), .A1(n599), .B0(n5442), .B1(n2217), .Y(n6977) );
  NOR3X8 U4244 ( .A(n4346), .B(n4347), .C(n3771), .Y(n4316) );
  AO21X4 U4245 ( .A0(net105311), .A1(net105312), .B0(net117723), .Y(net112330)
         );
  NAND4X4 U4246 ( .A(n6750), .B(n6749), .C(n6748), .D(n6747), .Y(n11432) );
  MX2XL U4247 ( .A(n3873), .B(\i_MIPS/Sign_Extend[2] ), .S0(n3593), .Y(
        \i_MIPS/n446 ) );
  BUFX16 U4248 ( .A(n4754), .Y(n5066) );
  CLKINVX8 U4249 ( .A(n5055), .Y(n4019) );
  OA22X4 U4250 ( .A0(n5403), .A1(n2113), .B0(n5446), .B1(n487), .Y(n6421) );
  OAI221X2 U4251 ( .A0(n5325), .A1(n2353), .B0(n5363), .B1(n903), .C0(n6421), 
        .Y(n6422) );
  XNOR2X4 U4252 ( .A(\i_MIPS/ID_EX[106] ), .B(\i_MIPS/ID_EX[107] ), .Y(
        \i_MIPS/ALU_Control/n18 ) );
  OAI211X2 U4253 ( .A0(n8471), .A1(n8467), .B0(n3906), .C0(n8464), .Y(n3985)
         );
  XOR2X4 U4254 ( .A(net105753), .B(n3025), .Y(n4347) );
  AO21X4 U4255 ( .A0(n7358), .A1(n7357), .B0(n5026), .Y(net104890) );
  CLKMX2X2 U4256 ( .A(n9596), .B(n9595), .S0(net114085), .Y(n9598) );
  OA22X4 U4257 ( .A0(n5249), .A1(n2114), .B0(n5289), .B1(n488), .Y(n8514) );
  BUFX20 U4258 ( .A(n5403), .Y(n5389) );
  OAI2BB1X4 U4259 ( .A0N(net106675), .A1N(net106674), .B0(n3989), .Y(net107856) );
  OA22X4 U4260 ( .A0(n5401), .A1(n2115), .B0(n5444), .B1(n489), .Y(n6460) );
  OAI221X4 U4261 ( .A0(n5329), .A1(n1272), .B0(n5354), .B1(n2901), .C0(n6496), 
        .Y(n6497) );
  BUFX16 U4262 ( .A(n5454), .Y(n5450) );
  OAI221X1 U4263 ( .A0(\i_MIPS/Register/register[2][22] ), .A1(n5090), .B0(
        \i_MIPS/Register/register[10][22] ), .B1(n5085), .C0(n7879), .Y(n7882)
         );
  NAND2X8 U4264 ( .A(n4718), .B(net134876), .Y(n9550) );
  INVX16 U4265 ( .A(n9550), .Y(n9445) );
  OAI221X2 U4266 ( .A0(n5325), .A1(n2018), .B0(n5354), .B1(n399), .C0(n6433), 
        .Y(n6434) );
  NOR2X6 U4267 ( .A(n8714), .B(n2934), .Y(n8717) );
  NAND2X1 U4268 ( .A(n5066), .B(\i_MIPS/ALUin1[1] ), .Y(n8678) );
  OAI221X4 U4269 ( .A0(n5067), .A1(\i_MIPS/n301 ), .B0(\i_MIPS/n299 ), .B1(
        n5056), .C0(n8678), .Y(n7787) );
  NAND2BX4 U4270 ( .AN(n7767), .B(n7488), .Y(n8116) );
  OR2X1 U4271 ( .A(n9488), .B(net107138), .Y(n3992) );
  CLKMX2X2 U4272 ( .A(n9486), .B(n9485), .S0(net114085), .Y(n9488) );
  NAND2X8 U4273 ( .A(n4723), .B(n4720), .Y(net107167) );
  OR2X4 U4274 ( .A(n8369), .B(net117711), .Y(net143555) );
  CLKINVX3 U4275 ( .A(n7401), .Y(n7403) );
  NAND2X8 U4276 ( .A(n3777), .B(net114073), .Y(n9547) );
  INVX6 U4277 ( .A(n6505), .Y(n11021) );
  OAI221X2 U4278 ( .A0(n5173), .A1(n2954), .B0(n5217), .B1(n1313), .C0(n6504), 
        .Y(n6505) );
  OR2X8 U4279 ( .A(n9294), .B(net117709), .Y(net144666) );
  INVX3 U4280 ( .A(n11418), .Y(n10780) );
  NAND4X4 U4281 ( .A(n6522), .B(n6520), .C(n6521), .D(n6519), .Y(n6523) );
  AND2X1 U4282 ( .A(net104171), .B(n11227), .Y(n4440) );
  OA22X2 U4283 ( .A0(n5917), .A1(n601), .B0(n5875), .B1(n2219), .Y(n11119) );
  OAI221X2 U4284 ( .A0(n10890), .A1(net143858), .B0(\i_MIPS/n520 ), .B1(
        net115789), .C0(n10889), .Y(\i_MIPS/N50 ) );
  OA22X4 U4285 ( .A0(n138), .A1(n2118), .B0(n5696), .B1(n492), .Y(n11195) );
  NAND2BX1 U4286 ( .AN(n10261), .B(n10256), .Y(n10175) );
  OAI22X2 U4287 ( .A0(n5651), .A1(n394), .B0(n5607), .B1(n2030), .Y(n4651) );
  INVX6 U4288 ( .A(n9202), .Y(n9442) );
  OAI31X2 U4289 ( .A0(n7), .A1(n9428), .A2(n9427), .B0(n9426), .Y(n4001) );
  XOR2X4 U4290 ( .A(n6472), .B(n4002), .Y(n4004) );
  XNOR2X4 U4291 ( .A(n6467), .B(DCACHE_addr[6]), .Y(n4005) );
  XNOR2X4 U4292 ( .A(n4370), .B(n4371), .Y(n4006) );
  OA22X1 U4293 ( .A0(\i_MIPS/Register/register[17][25] ), .A1(net118453), .B0(
        \i_MIPS/Register/register[25][25] ), .B1(net118479), .Y(n6884) );
  OA22X1 U4294 ( .A0(\i_MIPS/Register/register[17][2] ), .A1(net118453), .B0(
        \i_MIPS/Register/register[25][2] ), .B1(net118479), .Y(n7177) );
  OA22XL U4295 ( .A0(\i_MIPS/Register/register[1][24] ), .A1(net118455), .B0(
        \i_MIPS/Register/register[9][24] ), .B1(net118479), .Y(n6774) );
  MX2X2 U4296 ( .A(net107657), .B(net107656), .S0(n9302), .Y(n9053) );
  OA22X4 U4297 ( .A0(n5263), .A1(n2119), .B0(n5302), .B1(n494), .Y(n6491) );
  NAND4X2 U4298 ( .A(n7443), .B(n7442), .C(n7441), .D(n7440), .Y(n11498) );
  OA22XL U4299 ( .A0(n5251), .A1(n1082), .B0(n5298), .B1(n2705), .Y(n7442) );
  AOI2BB1X4 U4300 ( .A0N(net108005), .A1N(net108846), .B0(n8651), .Y(n8655) );
  OA22X4 U4301 ( .A0(n5259), .A1(n2120), .B0(n5307), .B1(n495), .Y(n6473) );
  XOR2X4 U4302 ( .A(n11368), .B(ICACHE_addr[26]), .Y(n11600) );
  AO22X4 U4303 ( .A0(ICACHE_addr[26]), .A1(mem_read_I), .B0(mem_write_I), .B1(
        n11368), .Y(n12858) );
  OAI2BB1X4 U4304 ( .A0N(net111723), .A1N(net108854), .B0(n124), .Y(n6716) );
  NAND2X2 U4305 ( .A(\i_MIPS/ALUin1[28] ), .B(n145), .Y(n7585) );
  NAND2X2 U4306 ( .A(n145), .B(n347), .Y(n7591) );
  OA22X4 U4307 ( .A0(n5258), .A1(n2121), .B0(n5307), .B1(n496), .Y(n6487) );
  INVXL U4308 ( .A(net110954), .Y(n4008) );
  AO21XL U4309 ( .A0(n8758), .A1(n8757), .B0(n3969), .Y(net104793) );
  OA21X4 U4310 ( .A0(n336), .A1(n5064), .B0(n7417), .Y(n7154) );
  NAND3BX2 U4311 ( .AN(n4818), .B(n7417), .C(n7416), .Y(n7842) );
  AOI2BB1X2 U4312 ( .A0N(n7689), .A1N(n9433), .B0(n9430), .Y(n6952) );
  AO21X4 U4313 ( .A0(net119263), .A1(net104985), .B0(net117723), .Y(net107696)
         );
  OA22X4 U4314 ( .A0(n5741), .A1(n2122), .B0(n5696), .B1(n497), .Y(n11116) );
  OAI221X2 U4315 ( .A0(n5173), .A1(n2955), .B0(n5217), .B1(n1314), .C0(n6508), 
        .Y(n6509) );
  AO21X4 U4316 ( .A0(net104916), .A1(net104917), .B0(net117623), .Y(net104915)
         );
  NAND2X2 U4317 ( .A(n11103), .B(n7400), .Y(n6838) );
  INVX3 U4318 ( .A(n6821), .Y(n6827) );
  XOR2X4 U4319 ( .A(n6393), .B(DCACHE_addr[5]), .Y(n6447) );
  BUFX8 U4320 ( .A(n5186), .Y(n5183) );
  NAND2X2 U4321 ( .A(n6711), .B(\i_MIPS/ALUin1[6] ), .Y(n7302) );
  NOR2BX4 U4322 ( .AN(n11053), .B(\i_MIPS/n497 ), .Y(n4785) );
  NAND2X8 U4323 ( .A(n4785), .B(n4723), .Y(net107170) );
  NAND2X6 U4324 ( .A(n4675), .B(n4785), .Y(net139756) );
  OAI2BB1X4 U4325 ( .A0N(n9540), .A1N(n11105), .B0(n9539), .Y(n9566) );
  XOR2X4 U4326 ( .A(n4011), .B(net104980), .Y(n4320) );
  MXI2X1 U4327 ( .A(\i_MIPS/n219 ), .B(\i_MIPS/n220 ), .S0(n3589), .Y(
        \i_MIPS/n342 ) );
  INVX3 U4328 ( .A(n3853), .Y(n6722) );
  AO22XL U4329 ( .A0(n2894), .A1(n3603), .B0(n3586), .B1(n3621), .Y(
        \i_MIPS/n402 ) );
  CLKINVX20 U4330 ( .A(n5066), .Y(n5063) );
  OAI221X4 U4331 ( .A0(n5329), .A1(n1333), .B0(n5354), .B1(n2986), .C0(n6506), 
        .Y(n6507) );
  INVXL U4332 ( .A(net106675), .Y(n4012) );
  INVX1 U4333 ( .A(n4012), .Y(n4013) );
  NAND2X6 U4334 ( .A(n11043), .B(n11042), .Y(n6472) );
  INVX8 U4335 ( .A(n9553), .Y(n8867) );
  OAI222X4 U4336 ( .A0(net107217), .A1(n7686), .B0(n4762), .B1(n9553), .C0(
        n7696), .C1(net117757), .Y(n7687) );
  NAND2X8 U4337 ( .A(n7102), .B(net134907), .Y(n9553) );
  BUFX20 U4338 ( .A(n5304), .Y(n5302) );
  OAI221X2 U4339 ( .A0(n5173), .A1(n2019), .B0(n5217), .B1(n400), .C0(n6482), 
        .Y(n6483) );
  OAI221X2 U4340 ( .A0(n8863), .A1(n9049), .B0(n8373), .B1(n3673), .C0(n8861), 
        .Y(n9052) );
  OAI221X4 U4341 ( .A0(n11), .A1(net143504), .B0(n3883), .B1(net143514), .C0(
        \i_MIPS/ALUin1[0] ), .Y(n8974) );
  NOR2X4 U4342 ( .A(n10850), .B(n6635), .Y(n6756) );
  AOI222X1 U4343 ( .A0(n3800), .A1(n11398), .B0(mem_rdata_D[22]), .B1(n131), 
        .C0(n12991), .C1(n5537), .Y(n10314) );
  OAI221X2 U4344 ( .A0(n5187), .A1(n2020), .B0(n5221), .B1(n401), .C0(n6491), 
        .Y(n6492) );
  AOI222X1 U4345 ( .A0(n3800), .A1(n11378), .B0(mem_rdata_D[2]), .B1(n132), 
        .C0(n13011), .C1(n5537), .Y(n10193) );
  INVX3 U4346 ( .A(n7869), .Y(n7860) );
  AND3X8 U4347 ( .A(net105448), .B(net105447), .C(net105449), .Y(n4349) );
  OA22X4 U4348 ( .A0(n5380), .A1(n2055), .B0(n5431), .B1(n430), .Y(n8339) );
  CLKBUFX2 U4349 ( .A(net108492), .Y(n4014) );
  AOI22X4 U4350 ( .A0(net118225), .A1(net110729), .B0(net105112), .B1(
        net118217), .Y(net139849) );
  BUFX8 U4351 ( .A(n4683), .Y(n5540) );
  MXI2X1 U4352 ( .A(n10766), .B(n10765), .S0(n5550), .Y(n10767) );
  AOI222X1 U4353 ( .A0(n3800), .A1(n11405), .B0(mem_rdata_D[29]), .B1(n129), 
        .C0(n12984), .C1(n5538), .Y(n10562) );
  AOI222X1 U4354 ( .A0(n3800), .A1(n11404), .B0(mem_rdata_D[28]), .B1(n131), 
        .C0(n12985), .C1(n5538), .Y(n10549) );
  AOI222X1 U4355 ( .A0(n3800), .A1(n11407), .B0(mem_rdata_D[31]), .B1(n132), 
        .C0(n12982), .C1(n5538), .Y(n10706) );
  AOI222X1 U4356 ( .A0(n3800), .A1(n11385), .B0(mem_rdata_D[9]), .B1(n131), 
        .C0(n13004), .C1(n5538), .Y(n10613) );
  CLKMX2X2 U4357 ( .A(\D_cache/cache[0][97] ), .B(n10669), .S0(n5162), .Y(
        \D_cache/n1020 ) );
  CLKMX2X2 U4358 ( .A(\D_cache/cache[1][97] ), .B(n10669), .S0(n5202), .Y(
        \D_cache/n1019 ) );
  CLKMX2X2 U4359 ( .A(\D_cache/cache[2][97] ), .B(n10669), .S0(n5230), .Y(
        \D_cache/n1018 ) );
  CLKMX2X2 U4360 ( .A(\D_cache/cache[3][97] ), .B(n10669), .S0(n5272), .Y(
        \D_cache/n1017 ) );
  CLKMX2X2 U4361 ( .A(\D_cache/cache[4][97] ), .B(n10669), .S0(n5317), .Y(
        \D_cache/n1016 ) );
  CLKMX2X2 U4362 ( .A(\D_cache/cache[5][97] ), .B(n10669), .S0(n5344), .Y(
        \D_cache/n1015 ) );
  CLKMX2X2 U4363 ( .A(\D_cache/cache[6][97] ), .B(n10669), .S0(n5368), .Y(
        \D_cache/n1014 ) );
  CLKMX2X2 U4364 ( .A(\D_cache/cache[7][97] ), .B(n10669), .S0(n3561), .Y(
        \D_cache/n1013 ) );
  CLKINVX20 U4365 ( .A(n5950), .Y(n5045) );
  BUFX20 U4366 ( .A(n11537), .Y(n5950) );
  NAND2XL U4367 ( .A(n3931), .B(n11005), .Y(n11530) );
  INVXL U4368 ( .A(net108161), .Y(n4017) );
  NAND4X4 U4369 ( .A(n7200), .B(n7199), .C(n7198), .D(n7197), .Y(n11410) );
  MX2XL U4370 ( .A(\i_MIPS/EX_MEM[6] ), .B(n4017), .S0(n3593), .Y(
        \i_MIPS/n398 ) );
  MX2X1 U4371 ( .A(net107656), .B(net107657), .S0(n8468), .Y(n8045) );
  NOR2X8 U4372 ( .A(net143547), .B(net143548), .Y(net139778) );
  AND2X2 U4373 ( .A(net118227), .B(n8070), .Y(net143548) );
  OAI221X4 U4374 ( .A0(\i_MIPS/ALUin1[18] ), .A1(n5064), .B0(
        \i_MIPS/ALUin1[19] ), .B1(n5056), .C0(n7033), .Y(n7682) );
  NAND4X4 U4375 ( .A(n8244), .B(n8243), .C(n8242), .D(n8241), .Y(n11484) );
  INVX8 U4376 ( .A(n11484), .Y(n10456) );
  AOI222X1 U4377 ( .A0(n4534), .A1(n11484), .B0(mem_rdata_D[108]), .B1(n129), 
        .C0(n13001), .C1(n5534), .Y(n10457) );
  OA22X2 U4378 ( .A0(n5385), .A1(n603), .B0(n5426), .B1(n2221), .Y(n9173) );
  CLKAND2X12 U4379 ( .A(n7491), .B(net110932), .Y(n4750) );
  AND3X8 U4380 ( .A(n4019), .B(n3930), .C(n5053), .Y(n4018) );
  MX2XL U4381 ( .A(\i_MIPS/EX_MEM[5] ), .B(net104794), .S0(n3599), .Y(
        \i_MIPS/n399 ) );
  NAND2X8 U4382 ( .A(n4630), .B(n8717), .Y(net104794) );
  BUFX12 U4383 ( .A(n6719), .Y(n4503) );
  XOR2X1 U4384 ( .A(\i_MIPS/ID_EX[114] ), .B(n10334), .Y(
        \i_MIPS/Hazard_detection/n11 ) );
  AOI222X4 U4385 ( .A0(n3800), .A1(n11380), .B0(mem_rdata_D[4]), .B1(n131), 
        .C0(n13009), .C1(n5538), .Y(n10753) );
  OA22X4 U4386 ( .A0(n5387), .A1(n2056), .B0(n5428), .B1(n431), .Y(n9012) );
  NAND2X4 U4387 ( .A(net118225), .B(net110147), .Y(net105448) );
  CLKBUFX6 U4388 ( .A(n5454), .Y(n5449) );
  AOI211X2 U4389 ( .A0(n10470), .A1(n10259), .B0(n4797), .C0(n10468), .Y(
        n10260) );
  INVX4 U4390 ( .A(n10262), .Y(n10470) );
  NAND4X4 U4391 ( .A(n9262), .B(n9261), .C(n9260), .D(n9259), .Y(n11457) );
  INVX8 U4392 ( .A(n11457), .Y(n10622) );
  AOI222X1 U4393 ( .A0(n4506), .A1(n11457), .B0(mem_rdata_D[81]), .B1(n129), 
        .C0(n12996), .C1(n5536), .Y(n10623) );
  MXI2X4 U4394 ( .A(n10190), .B(n10189), .S0(n5542), .Y(n10191) );
  MX2XL U4395 ( .A(\i_MIPS/ID_EX[74] ), .B(\i_MIPS/Sign_Extend[1] ), .S0(n3589), .Y(\i_MIPS/n447 ) );
  AOI222X1 U4396 ( .A0(n5541), .A1(n11421), .B0(mem_rdata_D[45]), .B1(n130), 
        .C0(n13000), .C1(n5540), .Y(n10809) );
  AO21X4 U4397 ( .A0(n8529), .A1(n8528), .B0(n5026), .Y(n10783) );
  INVX3 U4398 ( .A(n11388), .Y(n10462) );
  NAND4X4 U4399 ( .A(n8523), .B(n8522), .C(n8521), .D(n8520), .Y(n11387) );
  INVX8 U4400 ( .A(n11387), .Y(n10790) );
  AOI222X4 U4401 ( .A0(n3800), .A1(n11387), .B0(mem_rdata_D[11]), .B1(n130), 
        .C0(n13002), .C1(n5538), .Y(n10791) );
  CLKAND2X12 U4402 ( .A(n5044), .B(n11387), .Y(mem_wdata_D[11]) );
  CLKAND2X12 U4403 ( .A(n5951), .B(n11219), .Y(mem_wdata_I[0]) );
  AOI222X4 U4404 ( .A0(n3800), .A1(n11403), .B0(mem_rdata_D[27]), .B1(n130), 
        .C0(n12986), .C1(n5537), .Y(n10398) );
  OA22X4 U4405 ( .A0(n10891), .A1(n3767), .B0(n10894), .B1(n9536), .Y(n9363)
         );
  OA22X4 U4406 ( .A0(n10514), .A1(n3767), .B0(n10517), .B1(n9536), .Y(n8937)
         );
  OA22X4 U4407 ( .A0(n10417), .A1(n3767), .B0(n10420), .B1(n9536), .Y(n6752)
         );
  OAI222X4 U4408 ( .A0(n9552), .A1(n8205), .B0(n8372), .B1(n9452), .C0(
        net107217), .C1(n9425), .Y(n7604) );
  NAND2X4 U4409 ( .A(n8867), .B(net144224), .Y(n9452) );
  NAND4BX4 U4410 ( .AN(n8898), .B(n8897), .C(n8896), .D(n8895), .Y(n10512) );
  AOI33X4 U4411 ( .A0(n8894), .A1(n8893), .A2(net117743), .B0(n8892), .B1(
        n8891), .B2(net117743), .Y(n8895) );
  CLKBUFX4 U4412 ( .A(n5450), .Y(n5428) );
  OA22X4 U4413 ( .A0(n5401), .A1(n2123), .B0(n5444), .B1(n498), .Y(n6484) );
  OAI221X2 U4414 ( .A0(n9120), .A1(net117709), .B0(n9119), .B1(net117731), 
        .C0(n9118), .Y(net106596) );
  CLKMX2X3 U4415 ( .A(n8069), .B(n8068), .S0(net114087), .Y(n8070) );
  NAND2X4 U4416 ( .A(n8437), .B(n8438), .Y(n4636) );
  AO22X4 U4417 ( .A0(n5945), .A1(ICACHE_addr[27]), .B0(n5931), .B1(n11369), 
        .Y(n11064) );
  AO22X4 U4418 ( .A0(n5945), .A1(ICACHE_addr[11]), .B0(n5931), .B1(n11353), 
        .Y(n11122) );
  AO22X4 U4419 ( .A0(n5945), .A1(ICACHE_addr[10]), .B0(n5931), .B1(n11352), 
        .Y(n11127) );
  AO22X4 U4420 ( .A0(n5945), .A1(ICACHE_addr[15]), .B0(n5931), .B1(n11357), 
        .Y(n11131) );
  INVX6 U4421 ( .A(n6461), .Y(n11048) );
  INVXL U4422 ( .A(net111931), .Y(n4053) );
  XNOR2X4 U4423 ( .A(net105071), .B(n4361), .Y(n4056) );
  XNOR2X4 U4424 ( .A(net104861), .B(n4360), .Y(n4057) );
  XOR2X4 U4425 ( .A(n4060), .B(net105506), .Y(n4330) );
  AOI222X4 U4426 ( .A0(n4505), .A1(n11451), .B0(mem_rdata_D[75]), .B1(n133), 
        .C0(n13002), .C1(n5536), .Y(n10788) );
  MXI2X4 U4427 ( .A(n10788), .B(n10787), .S0(n5550), .Y(n10789) );
  AO21X4 U4428 ( .A0(net105142), .A1(net105143), .B0(net117623), .Y(net105463)
         );
  BUFX12 U4429 ( .A(n5403), .Y(n5388) );
  CLKAND2X8 U4430 ( .A(n6609), .B(net110470), .Y(n4721) );
  NAND3BX4 U4431 ( .AN(n9058), .B(n9057), .C(n9056), .Y(n10769) );
  AO22X4 U4432 ( .A0(mem_rdata_I[52]), .A1(n5941), .B0(n5567), .B1(n11269), 
        .Y(n9778) );
  AO22X4 U4433 ( .A0(mem_rdata_I[42]), .A1(n5941), .B0(n5567), .B1(n11260), 
        .Y(n9829) );
  AO22X4 U4434 ( .A0(mem_rdata_I[40]), .A1(n5941), .B0(n5567), .B1(n11258), 
        .Y(n9851) );
  AO22X4 U4435 ( .A0(mem_rdata_I[84]), .A1(n5941), .B0(n5569), .B1(n11300), 
        .Y(n9783) );
  AO22X4 U4436 ( .A0(mem_rdata_I[74]), .A1(n5941), .B0(n5569), .B1(n11291), 
        .Y(n9834) );
  AO22X4 U4437 ( .A0(mem_rdata_I[72]), .A1(n5941), .B0(n5569), .B1(n11289), 
        .Y(n9856) );
  AO22X4 U4438 ( .A0(mem_rdata_I[59]), .A1(n5944), .B0(n5566), .B1(n11276), 
        .Y(n9614) );
  AO22X4 U4439 ( .A0(mem_rdata_I[58]), .A1(n5944), .B0(n5566), .B1(n11275), 
        .Y(n6592) );
  AO22X4 U4440 ( .A0(mem_rdata_I[95]), .A1(n5944), .B0(n5569), .B1(n11311), 
        .Y(n6582) );
  AO22X4 U4441 ( .A0(mem_rdata_I[92]), .A1(n5944), .B0(n5569), .B1(n11308), 
        .Y(n9641) );
  AO22X4 U4442 ( .A0(mem_rdata_I[91]), .A1(n5944), .B0(n5569), .B1(n11307), 
        .Y(n9619) );
  AO22X4 U4443 ( .A0(mem_rdata_I[90]), .A1(n5944), .B0(n5569), .B1(n11306), 
        .Y(n6597) );
  BUFX12 U4444 ( .A(n5935), .Y(n5944) );
  NAND4X4 U4445 ( .A(n7874), .B(n7873), .C(n7872), .D(n7871), .Y(net105492) );
  NAND2X4 U4446 ( .A(net118215), .B(net105492), .Y(net105447) );
  AO22X4 U4447 ( .A0(mem_rdata_I[55]), .A1(n5944), .B0(n5567), .B1(n11272), 
        .Y(n10011) );
  AO22X4 U4448 ( .A0(mem_rdata_I[54]), .A1(n5944), .B0(n5567), .B1(n11271), 
        .Y(n9967) );
  AO22X4 U4449 ( .A0(mem_rdata_I[86]), .A1(n5941), .B0(n5569), .B1(n11302), 
        .Y(n9972) );
  AO22X4 U4450 ( .A0(mem_rdata_I[85]), .A1(n5944), .B0(n5569), .B1(n11301), 
        .Y(n9994) );
  AO22X4 U4451 ( .A0(mem_rdata_I[46]), .A1(n5940), .B0(n5568), .B1(n11264), 
        .Y(n10236) );
  AO22X4 U4452 ( .A0(mem_rdata_I[45]), .A1(n5940), .B0(n5568), .B1(n11263), 
        .Y(n10214) );
  AO22X4 U4453 ( .A0(mem_rdata_I[44]), .A1(n5940), .B0(n5568), .B1(n11262), 
        .Y(n10116) );
  AO22X4 U4454 ( .A0(mem_rdata_I[89]), .A1(n5940), .B0(n5569), .B1(n11305), 
        .Y(n10038) );
  AO22X4 U4455 ( .A0(mem_rdata_I[79]), .A1(n5940), .B0(n5569), .B1(n11296), 
        .Y(n10062) );
  AO22X4 U4456 ( .A0(mem_rdata_I[75]), .A1(n5940), .B0(n5569), .B1(n11292), 
        .Y(n10085) );
  AO22X4 U4457 ( .A0(mem_rdata_I[57]), .A1(n5940), .B0(n5568), .B1(n11274), 
        .Y(n10033) );
  AO22X4 U4458 ( .A0(mem_rdata_I[43]), .A1(n5940), .B0(n5568), .B1(n11261), 
        .Y(n10080) );
  AO22X4 U4459 ( .A0(mem_rdata_I[41]), .A1(n5940), .B0(n5567), .B1(n11259), 
        .Y(n9873) );
  AO22X4 U4460 ( .A0(mem_rdata_I[39]), .A1(n5944), .B0(n5567), .B1(n11257), 
        .Y(n9895) );
  AO22X4 U4461 ( .A0(mem_rdata_I[38]), .A1(n5941), .B0(n5567), .B1(n11256), 
        .Y(n9917) );
  AO22X4 U4462 ( .A0(mem_rdata_I[73]), .A1(n5944), .B0(n5569), .B1(n11290), 
        .Y(n9878) );
  AO22X4 U4463 ( .A0(mem_rdata_I[71]), .A1(n5940), .B0(n5569), .B1(n11288), 
        .Y(n9900) );
  AO22X4 U4464 ( .A0(mem_rdata_I[70]), .A1(n5942), .B0(n5569), .B1(n11287), 
        .Y(n9922) );
  AO22X4 U4465 ( .A0(mem_rdata_I[65]), .A1(n5940), .B0(n5569), .B1(n11282), 
        .Y(n10878) );
  OA22X2 U4466 ( .A0(n10410), .A1(n3879), .B0(n10413), .B1(n4495), .Y(n8437)
         );
  BUFX2 U4467 ( .A(n5938), .Y(n5934) );
  AOI222X1 U4468 ( .A0(n4534), .A1(n11500), .B0(mem_rdata_D[124]), .B1(n130), 
        .C0(n12985), .C1(n5534), .Y(n10543) );
  OA22X2 U4469 ( .A0(n10542), .A1(n3767), .B0(n10545), .B1(n9536), .Y(n7628)
         );
  OAI211X2 U4470 ( .A0(n8973), .A1(n9318), .B0(n8971), .C0(n8972), .Y(n8983)
         );
  INVXL U4471 ( .A(net105753), .Y(n4071) );
  NAND3BX1 U4472 ( .AN(n7779), .B(n3950), .C(n7778), .Y(n7795) );
  CLKBUFX2 U4473 ( .A(n4662), .Y(n5088) );
  OA22X1 U4474 ( .A0(\i_MIPS/Register/register[6][2] ), .A1(n5081), .B0(
        \i_MIPS/Register/register[14][2] ), .B1(n5076), .Y(n7201) );
  AOI22X4 U4475 ( .A0(net118215), .A1(net104794), .B0(net118225), .B1(
        net108729), .Y(net139850) );
  NAND4X4 U4476 ( .A(n7272), .B(n7271), .C(n7270), .D(n7269), .Y(n11382) );
  OA22X2 U4477 ( .A0(n5256), .A1(n605), .B0(n5299), .B1(n2223), .Y(n7271) );
  AO21X4 U4478 ( .A0(net106297), .A1(net106298), .B0(net117723), .Y(net111278)
         );
  BUFX8 U4479 ( .A(n5306), .Y(n5288) );
  OAI221X2 U4480 ( .A0(n5171), .A1(n2956), .B0(n5222), .B1(n1315), .C0(n6463), 
        .Y(n6464) );
  OA22X4 U4481 ( .A0(n5259), .A1(n2126), .B0(n5307), .B1(n501), .Y(n6463) );
  AOI222X1 U4482 ( .A0(n4534), .A1(n11479), .B0(mem_rdata_D[103]), .B1(n131), 
        .C0(n13006), .C1(n5534), .Y(n10675) );
  AOI33X2 U4483 ( .A0(n3950), .A1(n7433), .A2(n7434), .B0(n4007), .B1(n7432), 
        .B2(n3950), .Y(n7435) );
  OAI221X1 U4484 ( .A0(net118601), .A1(n8862), .B0(n8699), .B1(n8962), .C0(
        n7419), .Y(n8035) );
  OAI221X4 U4485 ( .A0(n253), .A1(n5064), .B0(n2184), .B1(n5056), .C0(n6841), 
        .Y(n8962) );
  INVX4 U4486 ( .A(n8112), .Y(n8461) );
  INVXL U4487 ( .A(n4342), .Y(n4078) );
  BUFX2 U4488 ( .A(n5938), .Y(n5935) );
  INVX8 U4489 ( .A(n10812), .Y(n7838) );
  INVXL U4490 ( .A(n4329), .Y(n4081) );
  NAND2X6 U4491 ( .A(\i_MIPS/ALUin1[7] ), .B(n6708), .Y(n8120) );
  OA22X2 U4492 ( .A0(n5331), .A1(n710), .B0(n5356), .B1(n2332), .Y(n8746) );
  OA22X2 U4493 ( .A0(n5331), .A1(n606), .B0(n5356), .B1(n2224), .Y(n8742) );
  OAI221X4 U4494 ( .A0(net107210), .A1(n3909), .B0(n7225), .B1(n3774), .C0(
        net117759), .Y(n7228) );
  OA22X1 U4495 ( .A0(n5374), .A1(n977), .B0(n5429), .B1(n2602), .Y(n8825) );
  XOR2X4 U4496 ( .A(n6423), .B(n12970), .Y(n6424) );
  AOI22X2 U4497 ( .A0(n4815), .A1(n10154), .B0(\i_MIPS/IF_ID[8] ), .B1(n2948), 
        .Y(n4809) );
  NAND2X2 U4498 ( .A(n4809), .B(n10174), .Y(n10259) );
  AO22XL U4499 ( .A0(n5157), .A1(n729), .B0(n5153), .B1(n2534), .Y(n8948) );
  OA22X4 U4500 ( .A0(n10625), .A1(n3877), .B0(n10628), .B1(n4495), .Y(n9271)
         );
  OA22X4 U4501 ( .A0(n10762), .A1(n3878), .B0(n10765), .B1(n4495), .Y(n9180)
         );
  OA22X4 U4502 ( .A0(n10897), .A1(n3878), .B0(n10900), .B1(n4495), .Y(n9362)
         );
  OAI221X4 U4503 ( .A0(n5324), .A1(n1273), .B0(n5351), .B1(n2902), .C0(n6390), 
        .Y(n10994) );
  OA22X4 U4504 ( .A0(n5400), .A1(n2887), .B0(n5429), .B1(n1269), .Y(n6390) );
  NOR2X6 U4505 ( .A(n10994), .B(n10993), .Y(n6393) );
  MXI2X4 U4506 ( .A(\i_MIPS/ID_EX[111] ), .B(\i_MIPS/ID_EX[84] ), .S0(
        \i_MIPS/ID_EX_5 ), .Y(n6753) );
  INVXL U4507 ( .A(n4345), .Y(n4091) );
  OAI2BB2X4 U4508 ( .B0(n9571), .B1(n9570), .A0N(n9569), .A1N(n9568), .Y(n9572) );
  INVX8 U4509 ( .A(n11469), .Y(n10558) );
  NAND4X4 U4510 ( .A(n6972), .B(n6971), .C(n6970), .D(n6969), .Y(n11469) );
  NAND2X2 U4511 ( .A(\i_MIPS/ALUin1[24] ), .B(n143), .Y(n8633) );
  NAND3BX4 U4512 ( .AN(n4740), .B(n6706), .C(n8121), .Y(net110928) );
  AOI2BB1X1 U4513 ( .A0N(n9211), .A1N(n9210), .B0(net107841), .Y(n9212) );
  NAND4BX4 U4514 ( .AN(n7796), .B(n7795), .C(n7794), .D(n7793), .Y(n10812) );
  AO22X4 U4515 ( .A0(mem_rdata_I[81]), .A1(n5945), .B0(n5569), .B1(n11298), 
        .Y(n6572) );
  AO22X4 U4516 ( .A0(mem_rdata_I[64]), .A1(n5945), .B0(n5569), .B1(n11281), 
        .Y(n6557) );
  AO22X4 U4517 ( .A0(n5945), .A1(ICACHE_addr[23]), .B0(n5931), .B1(n11365), 
        .Y(n11063) );
  AO22X4 U4518 ( .A0(n5945), .A1(ICACHE_addr[29]), .B0(n5931), .B1(n11371), 
        .Y(n11068) );
  AO22X4 U4519 ( .A0(n5945), .A1(ICACHE_addr[28]), .B0(n5931), .B1(n11370), 
        .Y(n11066) );
  AO22X4 U4520 ( .A0(n5945), .A1(ICACHE_addr[22]), .B0(n5931), .B1(n11364), 
        .Y(n11065) );
  AO22X4 U4521 ( .A0(n5945), .A1(ICACHE_addr[20]), .B0(n5930), .B1(n11362), 
        .Y(n11215) );
  NAND4X6 U4522 ( .A(n7918), .B(n7917), .C(n7916), .D(n7915), .Y(n11430) );
  OA22X2 U4523 ( .A0(n5254), .A1(n609), .B0(n5294), .B1(n2227), .Y(n7917) );
  AND3X4 U4524 ( .A(net105436), .B(net105435), .C(net105434), .Y(n4348) );
  OAI221X4 U4525 ( .A0(\i_MIPS/ALUin1[19] ), .A1(n5064), .B0(
        \i_MIPS/ALUin1[20] ), .B1(n5056), .C0(n6676), .Y(n7584) );
  OAI221X4 U4526 ( .A0(\i_MIPS/ALUin1[19] ), .A1(n5071), .B0(
        \i_MIPS/ALUin1[20] ), .B1(n5068), .C0(n7408), .Y(n7844) );
  NAND4X4 U4527 ( .A(n8599), .B(n8598), .C(n8597), .D(n8596), .Y(n11490) );
  AOI222X1 U4528 ( .A0(n4534), .A1(n11490), .B0(mem_rdata_D[114]), .B1(n133), 
        .C0(n12995), .C1(n5534), .Y(n10635) );
  INVXL U4529 ( .A(n4343), .Y(n4092) );
  NAND2X6 U4530 ( .A(n3972), .B(n11009), .Y(n6439) );
  OAI221XL U4531 ( .A0(net108490), .A1(net117709), .B0(net108491), .B1(
        net117731), .C0(n4014), .Y(n4093) );
  CLKAND2X12 U4532 ( .A(net105477), .B(n6609), .Y(n4784) );
  OAI221X1 U4533 ( .A0(\i_MIPS/Register/register[18][22] ), .A1(n5090), .B0(
        \i_MIPS/Register/register[26][22] ), .B1(n5085), .C0(n7896), .Y(n7899)
         );
  OA22X1 U4534 ( .A0(\i_MIPS/Register/register[22][22] ), .A1(n5082), .B0(
        \i_MIPS/Register/register[30][22] ), .B1(n5078), .Y(n7896) );
  INVXL U4535 ( .A(n3021), .Y(n4094) );
  NAND2X4 U4536 ( .A(\i_MIPS/IF_ID[2] ), .B(\i_MIPS/Sign_Extend[0] ), .Y(
        n10134) );
  NOR4X1 U4537 ( .A(\i_MIPS/Sign_Extend[5] ), .B(\i_MIPS/Sign_Extend[0] ), .C(
        n11576), .D(\i_MIPS/n518 ), .Y(n9602) );
  AOI2BB1X4 U4538 ( .A0N(n5073), .A1N(n347), .B0(n4793), .Y(n6841) );
  OA22X4 U4539 ( .A0(n5391), .A1(n2158), .B0(n5434), .B1(n539), .Y(n8075) );
  BUFX8 U4540 ( .A(n5397), .Y(n5391) );
  AO21X4 U4541 ( .A0(net105008), .A1(net105009), .B0(net117625), .Y(net105798)
         );
  OA22X4 U4542 ( .A0(n5400), .A1(n2970), .B0(n5453), .B1(n1321), .Y(n6510) );
  OA22X4 U4543 ( .A0(n5400), .A1(n2129), .B0(n5453), .B1(n504), .Y(n6489) );
  OA22X2 U4544 ( .A0(n5400), .A1(n1271), .B0(n5440), .B1(n2895), .Y(n6558) );
  NAND2X2 U4545 ( .A(n143), .B(n344), .Y(n6920) );
  AO22X4 U4546 ( .A0(mem_rdata_I[63]), .A1(n5945), .B0(n5566), .B1(n11280), 
        .Y(n6577) );
  AO22X4 U4547 ( .A0(mem_rdata_I[49]), .A1(n5945), .B0(n5566), .B1(n11267), 
        .Y(n6567) );
  AO22X4 U4548 ( .A0(mem_rdata_I[36]), .A1(n5945), .B0(n5566), .B1(n11254), 
        .Y(n6542) );
  AO22X4 U4549 ( .A0(mem_rdata_I[62]), .A1(n5943), .B0(n5566), .B1(n11279), 
        .Y(n9666) );
  AO22X4 U4550 ( .A0(mem_rdata_I[61]), .A1(n5943), .B0(n5566), .B1(n11278), 
        .Y(n9688) );
  AO22X4 U4551 ( .A0(mem_rdata_I[60]), .A1(n5944), .B0(n5566), .B1(n11277), 
        .Y(n9636) );
  BUFX20 U4552 ( .A(n11079), .Y(n5569) );
  XNOR2X4 U4553 ( .A(n6490), .B(DCACHE_addr[10]), .Y(n4096) );
  XOR2X4 U4554 ( .A(n6486), .B(n2998), .Y(n4097) );
  AND2X8 U4555 ( .A(n4403), .B(n4402), .Y(n4098) );
  MX2XL U4556 ( .A(n3555), .B(n4092), .S0(n3605), .Y(\i_MIPS/n351 ) );
  OA22X1 U4557 ( .A0(n5392), .A1(n978), .B0(n5438), .B1(n2603), .Y(n7444) );
  NAND4X4 U4558 ( .A(n7447), .B(n7446), .C(n7445), .D(n7444), .Y(n11466) );
  OA22X2 U4559 ( .A0(n9940), .A1(n3766), .B0(n9947), .B1(n9536), .Y(n7278) );
  XOR2X4 U4560 ( .A(n4099), .B(n5024), .Y(n6512) );
  MX2XL U4561 ( .A(n3553), .B(n4094), .S0(n3605), .Y(\i_MIPS/n345 ) );
  MX2XL U4562 ( .A(n11095), .B(n3709), .S0(n3601), .Y(\i_MIPS/n315 ) );
  OAI221X1 U4563 ( .A0(n10914), .A1(n5560), .B0(n5557), .B1(n10913), .C0(
        n10912), .Y(\i_MIPS/PC/n39 ) );
  NAND2X6 U4564 ( .A(net105375), .B(net105376), .Y(n4356) );
  NAND4X4 U4565 ( .A(n7352), .B(n7351), .C(n7350), .D(n7349), .Y(n11383) );
  OA22X1 U4566 ( .A0(n5395), .A1(n979), .B0(n5439), .B1(n2604), .Y(n7349) );
  INVX8 U4567 ( .A(n11383), .Y(n10680) );
  OAI221X4 U4568 ( .A0(net111128), .A1(net117711), .B0(net111129), .B1(
        net117731), .C0(net111130), .Y(net104884) );
  NOR2BX4 U4569 ( .AN(\i_MIPS/jump_addr[18] ), .B(\i_MIPS/n504 ), .Y(n4789) );
  INVXL U4570 ( .A(n4355), .Y(n4100) );
  INVXL U4571 ( .A(net111763), .Y(n4101) );
  NAND2X2 U4572 ( .A(net110429), .B(net110430), .Y(net110129) );
  NAND2X1 U4573 ( .A(\i_MIPS/ID_EX[81] ), .B(n3674), .Y(net108779) );
  AOI22X4 U4574 ( .A0(net118217), .A1(net105234), .B0(net118227), .B1(
        net109616), .Y(net139862) );
  OAI221X2 U4575 ( .A0(n5327), .A1(n2022), .B0(n5352), .B1(n403), .C0(n6460), 
        .Y(n6461) );
  OAI221X2 U4576 ( .A0(n5327), .A1(n2023), .B0(n5352), .B1(n404), .C0(n6453), 
        .Y(n6454) );
  INVX3 U4577 ( .A(n8703), .Y(n8114) );
  OAI221X4 U4578 ( .A0(n183), .A1(n5071), .B0(n2949), .B1(n5067), .C0(n8109), 
        .Y(n8703) );
  AOI222X4 U4579 ( .A0(net107652), .A1(n4653), .B0(n7160), .B1(n8208), .C0(
        n8976), .C1(n7787), .Y(n7163) );
  NAND4X2 U4580 ( .A(n8603), .B(n8602), .C(n8601), .D(n8600), .Y(n11458) );
  OA22X2 U4581 ( .A0(n5249), .A1(n711), .B0(n5289), .B1(n2333), .Y(n8602) );
  AO21X4 U4582 ( .A0(n8890), .A1(n4708), .B0(n8889), .Y(n8892) );
  INVX3 U4583 ( .A(n8892), .Y(n8894) );
  OA22X4 U4584 ( .A0(n5393), .A1(n2161), .B0(n5431), .B1(n542), .Y(n8421) );
  AOI222X1 U4585 ( .A0(n4534), .A1(n11477), .B0(mem_rdata_D[101]), .B1(n130), 
        .C0(n13008), .C1(n5534), .Y(n10892) );
  NAND4X6 U4586 ( .A(n9349), .B(n9348), .C(n9347), .D(n9346), .Y(n11477) );
  NOR2X8 U4587 ( .A(n6513), .B(n6512), .Y(n6514) );
  AND2XL U4588 ( .A(n5046), .B(n11270), .Y(n12950) );
  INVX20 U4589 ( .A(n4107), .Y(mem_addr_I[9]) );
  AO22X1 U4590 ( .A0(ICACHE_addr[7]), .A1(mem_read_I), .B0(n5048), .B1(n11349), 
        .Y(n12877) );
  INVX20 U4591 ( .A(n4109), .Y(mem_addr_I[10]) );
  AO22X1 U4592 ( .A0(ICACHE_addr[8]), .A1(mem_read_I), .B0(n5046), .B1(n11350), 
        .Y(n12876) );
  CLKINVX6 U4593 ( .A(n12875), .Y(n4111) );
  INVX20 U4594 ( .A(n4111), .Y(mem_addr_I[11]) );
  AO22X1 U4595 ( .A0(ICACHE_addr[9]), .A1(mem_read_I), .B0(n5047), .B1(n11351), 
        .Y(n12875) );
  INVX20 U4596 ( .A(n4113), .Y(mem_addr_I[12]) );
  AO22X1 U4597 ( .A0(ICACHE_addr[10]), .A1(mem_read_I), .B0(n5048), .B1(n11352), .Y(n12874) );
  INVX20 U4598 ( .A(n4115), .Y(mem_addr_I[13]) );
  AO22X1 U4599 ( .A0(ICACHE_addr[11]), .A1(mem_read_I), .B0(n5046), .B1(n11353), .Y(n12873) );
  AND2XL U4600 ( .A(n5046), .B(n11273), .Y(n12947) );
  INVX20 U4601 ( .A(n4119), .Y(mem_addr_I[14]) );
  AND2XL U4602 ( .A(n5046), .B(n11276), .Y(n12944) );
  INVX20 U4603 ( .A(n4123), .Y(mem_addr_I[15]) );
  AO22X1 U4604 ( .A0(ICACHE_addr[13]), .A1(mem_read_I), .B0(n5048), .B1(n11355), .Y(n12871) );
  INVX20 U4605 ( .A(n4125), .Y(mem_addr_I[16]) );
  AO22X1 U4606 ( .A0(ICACHE_addr[14]), .A1(mem_read_I), .B0(n5046), .B1(n11356), .Y(n12870) );
  AND2XL U4607 ( .A(n5046), .B(n11279), .Y(n12941) );
  AND2XL U4608 ( .A(n5046), .B(n11282), .Y(n12938) );
  AO22X1 U4609 ( .A0(ICACHE_addr[17]), .A1(mem_read_I), .B0(mem_write_I), .B1(
        n11359), .Y(n12867) );
  INVX20 U4610 ( .A(n4135), .Y(mem_addr_I[20]) );
  AOI222X1 U4611 ( .A0(n3800), .A1(n11381), .B0(mem_rdata_D[5]), .B1(n129), 
        .C0(n13008), .C1(n5538), .Y(n10898) );
  NAND4X6 U4612 ( .A(n9357), .B(n9356), .C(n9355), .D(n9354), .Y(n11381) );
  OAI211X2 U4613 ( .A0(net107217), .A1(n3896), .B0(n8706), .C0(n8707), .Y(
        n8709) );
  NAND2BX4 U4614 ( .AN(n7774), .B(net110131), .Y(n7778) );
  NAND2XL U4615 ( .A(net105462), .B(net105463), .Y(n10526) );
  NAND2X4 U4616 ( .A(\i_MIPS/ALUin1[26] ), .B(n6948), .Y(n7424) );
  INVX4 U4617 ( .A(n3973), .Y(n6948) );
  OAI31X4 U4618 ( .A0(net109668), .A1(n142), .A2(net109513), .B0(n4275), .Y(
        n4274) );
  INVX4 U4619 ( .A(net110430), .Y(net109668) );
  AOI222X4 U4620 ( .A0(n4505), .A1(n11455), .B0(mem_rdata_D[79]), .B1(n132), 
        .C0(n12998), .C1(n5535), .Y(n10448) );
  CLKINVX8 U4621 ( .A(n5045), .Y(n5047) );
  AND2XL U4622 ( .A(n5046), .B(n11285), .Y(n12935) );
  AND2XL U4623 ( .A(n5048), .B(n11267), .Y(n12953) );
  AND2XL U4624 ( .A(n5047), .B(n11271), .Y(n12949) );
  AND2XL U4625 ( .A(n5046), .B(n11288), .Y(n12932) );
  AND2XL U4626 ( .A(n5048), .B(n11269), .Y(n12951) );
  AND2XL U4627 ( .A(n5047), .B(n11274), .Y(n12946) );
  AND2XL U4628 ( .A(n5046), .B(n11291), .Y(n12929) );
  AND2XL U4629 ( .A(n5048), .B(n11272), .Y(n12948) );
  AND2XL U4630 ( .A(n5047), .B(n11277), .Y(n12943) );
  AND2XL U4631 ( .A(n5046), .B(n11294), .Y(n12926) );
  AND2XL U4632 ( .A(n5048), .B(n11275), .Y(n12945) );
  AND2XL U4633 ( .A(n5047), .B(n11280), .Y(n12940) );
  AND2XL U4634 ( .A(n5046), .B(n11297), .Y(n12923) );
  AND2XL U4635 ( .A(n5048), .B(n11278), .Y(n12942) );
  AND2XL U4636 ( .A(n5047), .B(n11283), .Y(n12937) );
  AND2XL U4637 ( .A(n5046), .B(n11299), .Y(n12920) );
  AND2XL U4638 ( .A(n5048), .B(n11281), .Y(n12939) );
  AND2XL U4639 ( .A(n5047), .B(n11286), .Y(n12934) );
  AND2XL U4640 ( .A(n5046), .B(n11302), .Y(n12917) );
  AND2XL U4641 ( .A(n5048), .B(n11284), .Y(n12936) );
  AND2XL U4642 ( .A(n5047), .B(n11289), .Y(n12931) );
  AND2XL U4643 ( .A(n5046), .B(n11305), .Y(n12914) );
  AND2XL U4644 ( .A(n5048), .B(n11287), .Y(n12933) );
  AND2XL U4645 ( .A(n5047), .B(n11292), .Y(n12928) );
  AND2XL U4646 ( .A(n5046), .B(n11308), .Y(n12911) );
  AND2XL U4647 ( .A(n5048), .B(n11290), .Y(n12930) );
  AND2XL U4648 ( .A(n5047), .B(n11295), .Y(n12925) );
  AND2XL U4649 ( .A(n5046), .B(n11311), .Y(n12908) );
  AND2XL U4650 ( .A(n5048), .B(n11293), .Y(n12927) );
  AND2XL U4651 ( .A(n5047), .B(n11298), .Y(n12922) );
  AND2XL U4652 ( .A(n5046), .B(n11314), .Y(n12905) );
  AND2XL U4653 ( .A(n5048), .B(n11296), .Y(n12924) );
  AND2XL U4654 ( .A(n5047), .B(n11300), .Y(n12919) );
  AND2XL U4655 ( .A(n5046), .B(n11317), .Y(n12902) );
  AND2XL U4656 ( .A(n5048), .B(net103785), .Y(n12921) );
  AND2XL U4657 ( .A(n5047), .B(n11303), .Y(n12916) );
  AND2XL U4658 ( .A(n5046), .B(n11320), .Y(n12899) );
  AND2XL U4659 ( .A(n5048), .B(n11301), .Y(n12918) );
  AND2XL U4660 ( .A(n5047), .B(n11306), .Y(n12913) );
  AND2XL U4661 ( .A(n5046), .B(n11323), .Y(n12896) );
  AND2XL U4662 ( .A(n5048), .B(n11304), .Y(n12915) );
  AND2XL U4663 ( .A(n5047), .B(n11309), .Y(n12910) );
  AND2XL U4664 ( .A(n5046), .B(n11326), .Y(n12893) );
  AND2XL U4665 ( .A(n5048), .B(n11307), .Y(n12912) );
  AND2XL U4666 ( .A(n5047), .B(n11312), .Y(n12907) );
  AND2XL U4667 ( .A(n5046), .B(n11329), .Y(n12890) );
  AND2XL U4668 ( .A(n5048), .B(n11310), .Y(n12909) );
  AND2XL U4669 ( .A(n5047), .B(n11315), .Y(n12904) );
  AND2XL U4670 ( .A(n5046), .B(n11331), .Y(n12887) );
  AND2XL U4671 ( .A(n5048), .B(n11313), .Y(n12906) );
  AND2XL U4672 ( .A(n5047), .B(n11318), .Y(n12901) );
  AND2XL U4673 ( .A(n5046), .B(n11334), .Y(n12884) );
  AND2XL U4674 ( .A(n5048), .B(n11316), .Y(n12903) );
  AND2XL U4675 ( .A(n5047), .B(n11321), .Y(n12898) );
  AND2XL U4676 ( .A(n5046), .B(n11337), .Y(n12881) );
  AND2XL U4677 ( .A(n5048), .B(n11319), .Y(n12900) );
  AND2XL U4678 ( .A(n5047), .B(n11324), .Y(n12895) );
  AND2XL U4679 ( .A(n5048), .B(n11322), .Y(n12897) );
  AND2XL U4680 ( .A(n5047), .B(n11327), .Y(n12892) );
  AND2XL U4681 ( .A(n5048), .B(n11325), .Y(n12894) );
  AND2XL U4682 ( .A(n5047), .B(net103753), .Y(n12889) );
  AND2XL U4683 ( .A(n5048), .B(n11328), .Y(n12891) );
  AND2XL U4684 ( .A(n5047), .B(n11332), .Y(n12886) );
  AND2XL U4685 ( .A(n5048), .B(n11330), .Y(n12888) );
  AND2XL U4686 ( .A(n5047), .B(n11335), .Y(n12883) );
  AND2XL U4687 ( .A(n5048), .B(n11333), .Y(n12885) );
  CLKAND2X12 U4688 ( .A(n9945), .B(\i_MIPS/n264 ), .Y(n4719) );
  AND2XL U4689 ( .A(n5048), .B(n11336), .Y(n12882) );
  AND2XL U4690 ( .A(n5048), .B(n11339), .Y(n12880) );
  OAI221X1 U4691 ( .A0(n10845), .A1(net143858), .B0(\i_MIPS/n497 ), .B1(
        net115791), .C0(n10844), .Y(\i_MIPS/N73 ) );
  AO21X4 U4692 ( .A0(net111570), .A1(net108297), .B0(net134145), .Y(net108003)
         );
  AOI2BB1XL U4693 ( .A0N(n3668), .A1N(\i_MIPS/n300 ), .B0(net108299), .Y(
        net108290) );
  AOI21X2 U4694 ( .A0(\i_MIPS/ID_EX[78] ), .A1(n4021), .B0(net112549), .Y(
        net112555) );
  OAI31X2 U4695 ( .A0(n3968), .A1(net108852), .A2(net109668), .B0(net108851), 
        .Y(net109666) );
  NAND3BX4 U4696 ( .AN(n3577), .B(n4276), .C(n4277), .Y(net109510) );
  AOI211X2 U4697 ( .A0(n3974), .A1(n4278), .B0(net112219), .C0(n3577), .Y(
        net112214) );
  NAND4X4 U4698 ( .A(n4301), .B(n4302), .C(n4303), .D(n4304), .Y(net105257) );
  CLKMX2X2 U4699 ( .A(n4281), .B(n4282), .S0(net114087), .Y(n4280) );
  NOR4X1 U4700 ( .A(n4292), .B(n4293), .C(n4294), .D(n4295), .Y(n4281) );
  NAND4X1 U4701 ( .A(n4297), .B(n4298), .C(n4299), .D(n4300), .Y(n4292) );
  OA22XL U4702 ( .A0(\i_MIPS/Register/register[5][15] ), .A1(net118399), .B0(
        \i_MIPS/Register/register[13][15] ), .B1(net118423), .Y(n4298) );
  INVX8 U4703 ( .A(net118417), .Y(net118399) );
  OA22XL U4704 ( .A0(\i_MIPS/Register/register[3][15] ), .A1(net118351), .B0(
        \i_MIPS/Register/register[11][15] ), .B1(net118375), .Y(n4299) );
  INVX3 U4705 ( .A(net134682), .Y(net118375) );
  OA22XL U4706 ( .A0(\i_MIPS/Register/register[7][15] ), .A1(net118303), .B0(
        \i_MIPS/Register/register[15][15] ), .B1(net118327), .Y(n4300) );
  INVX6 U4707 ( .A(net118321), .Y(net118303) );
  OAI221XL U4708 ( .A0(\i_MIPS/Register/register[2][15] ), .A1(net117635), 
        .B0(\i_MIPS/Register/register[10][15] ), .B1(net117653), .C0(n4296), 
        .Y(n4293) );
  OA22XL U4709 ( .A0(\i_MIPS/Register/register[6][15] ), .A1(net117673), .B0(
        \i_MIPS/Register/register[14][15] ), .B1(net117691), .Y(n4296) );
  BUFX16 U4710 ( .A(net117697), .Y(net117691) );
  AO22X1 U4711 ( .A0(net118267), .A1(n268), .B0(net118295), .B1(n913), .Y(
        n4294) );
  AO22XL U4712 ( .A0(net118235), .A1(n186), .B0(net118259), .B1(n324), .Y(
        n4295) );
  NOR4X1 U4713 ( .A(n4283), .B(n4284), .C(n4285), .D(n4286), .Y(n4282) );
  NAND4X1 U4714 ( .A(n4288), .B(n4289), .C(n4290), .D(n4291), .Y(n4283) );
  OA22XL U4715 ( .A0(\i_MIPS/Register/register[21][15] ), .A1(net118399), .B0(
        \i_MIPS/Register/register[29][15] ), .B1(net118423), .Y(n4289) );
  OA22XL U4716 ( .A0(\i_MIPS/Register/register[19][15] ), .A1(net118351), .B0(
        \i_MIPS/Register/register[27][15] ), .B1(net118375), .Y(n4290) );
  OA22XL U4717 ( .A0(\i_MIPS/Register/register[23][15] ), .A1(net118303), .B0(
        \i_MIPS/Register/register[31][15] ), .B1(net118327), .Y(n4291) );
  OA22XL U4718 ( .A0(\i_MIPS/Register/register[22][15] ), .A1(net117673), .B0(
        \i_MIPS/Register/register[30][15] ), .B1(net117691), .Y(n4287) );
  AO22X1 U4719 ( .A0(net118267), .A1(n269), .B0(net118295), .B1(n914), .Y(
        n4285) );
  AO22XL U4720 ( .A0(net118235), .A1(n187), .B0(net118259), .B1(n325), .Y(
        n4286) );
  NAND2XL U4721 ( .A(net105581), .B(net105582), .Y(net105236) );
  AOI221X2 U4722 ( .A0(n4306), .A1(n4307), .B0(n4308), .B1(n4309), .C0(
        net107841), .Y(n4301) );
  BUFX20 U4723 ( .A(net117751), .Y(net117747) );
  NAND2XL U4724 ( .A(net108625), .B(net108623), .Y(n4307) );
  NAND2XL U4725 ( .A(n124), .B(n3857), .Y(n4308) );
  NAND2X4 U4726 ( .A(net109965), .B(n3674), .Y(net107688) );
  OA22X2 U4727 ( .A0(net107230), .A1(net107661), .B0(net135772), .B1(net107987), .Y(n4303) );
  INVX8 U4728 ( .A(net144227), .Y(net135772) );
  NAND2X8 U4729 ( .A(net134907), .B(net108632), .Y(net107977) );
  INVX3 U4730 ( .A(net105257), .Y(net111581) );
  MX2XL U4731 ( .A(n12970), .B(net105257), .S0(n3599), .Y(\i_MIPS/n384 ) );
  INVXL U4732 ( .A(net103753), .Y(n4311) );
  NAND4X1 U4733 ( .A(net106679), .B(net106680), .C(net106681), .D(net106682), 
        .Y(net103753) );
  NAND4X1 U4734 ( .A(net106692), .B(net106693), .C(net106694), .D(net106695), 
        .Y(net103849) );
  NAND4X8 U4735 ( .A(n3999), .B(n4316), .C(n4317), .D(n4315), .Y(net106828) );
  NAND2X8 U4736 ( .A(net107134), .B(net107135), .Y(net104828) );
  OAI221X2 U4737 ( .A0(net112118), .A1(net117713), .B0(net112119), .B1(
        net117733), .C0(net112120), .Y(net105283) );
  AO21X4 U4738 ( .A0(net105288), .A1(n3953), .B0(net117625), .Y(net105269) );
  AO21X4 U4739 ( .A0(net105075), .A1(net105076), .B0(net117625), .Y(net105430)
         );
  OAI221X2 U4740 ( .A0(net111762), .A1(net117713), .B0(net111763), .B1(
        net117731), .C0(net111764), .Y(net104861) );
  NAND2X6 U4741 ( .A(n3002), .B(net105412), .Y(n4360) );
  AO21X4 U4742 ( .A0(net104866), .A1(net104867), .B0(net117625), .Y(net105412)
         );
  AO21X2 U4743 ( .A0(net105751), .A1(net105752), .B0(net117625), .Y(net105732)
         );
  OAI221X2 U4744 ( .A0(net111276), .A1(net117711), .B0(net111277), .B1(
        net117731), .C0(net111278), .Y(net106290) );
  CLKINVX3 U4745 ( .A(net111216), .Y(net105834) );
  XOR2X4 U4746 ( .A(n4356), .B(n4357), .Y(n4350) );
  CLKINVX8 U4747 ( .A(net111041), .Y(net105375) );
  AO21X2 U4748 ( .A0(net105265), .A1(net105264), .B0(net117625), .Y(net105376)
         );
  OAI221X2 U4749 ( .A0(net110953), .A1(net117711), .B0(net110954), .B1(
        net117731), .C0(net110955), .Y(net104166) );
  XOR2X4 U4750 ( .A(n4355), .B(n4354), .Y(n4351) );
  AO21X4 U4751 ( .A0(net105119), .A1(net105120), .B0(net117625), .Y(net105783)
         );
  OAI221X2 U4752 ( .A0(net110798), .A1(net117711), .B0(net110799), .B1(
        net117731), .C0(net110800), .Y(net104725) );
  XOR2X4 U4753 ( .A(n3947), .B(n10403), .Y(n4353) );
  INVX1 U4754 ( .A(net110473), .Y(net49779) );
  CLKBUFX3 U4755 ( .A(net36639), .Y(net118581) );
  NAND2X4 U4756 ( .A(net117741), .B(net105492), .Y(net105436) );
  AO21X4 U4757 ( .A0(net104698), .A1(net104699), .B0(net117625), .Y(net105195)
         );
  XOR2X4 U4758 ( .A(n4345), .B(n4344), .Y(n4338) );
  NAND2X4 U4759 ( .A(net139778), .B(net105798), .Y(n4344) );
  OAI221X2 U4760 ( .A0(net109839), .A1(net117711), .B0(net109840), .B1(
        net117731), .C0(net109841), .Y(net105003) );
  XOR2X4 U4761 ( .A(n4343), .B(n10659), .Y(n4339) );
  OAI221X2 U4762 ( .A0(net109673), .A1(net117711), .B0(net109674), .B1(
        net117731), .C0(net109675), .Y(net104934) );
  XOR2X4 U4763 ( .A(n4342), .B(n4341), .Y(n4340) );
  OAI221X2 U4764 ( .A0(net109527), .A1(net117711), .B0(net109528), .B1(
        net117731), .C0(net109529), .Y(net105227) );
  AOI22X4 U4765 ( .A0(net118215), .A1(n3616), .B0(net118227), .B1(net109447), 
        .Y(net139865) );
  XOR2X4 U4766 ( .A(n4336), .B(n3021), .Y(n4332) );
  AOI22X4 U4767 ( .A0(net118215), .A1(n3971), .B0(net118227), .B1(net109129), 
        .Y(net139777) );
  AO21X2 U4768 ( .A0(net104721), .A1(net119104), .B0(net117623), .Y(net105764)
         );
  XOR2X4 U4769 ( .A(n4334), .B(n4335), .Y(n4333) );
  AO21X2 U4770 ( .A0(net104962), .A1(n3667), .B0(net117623), .Y(net105531) );
  OAI221X2 U4771 ( .A0(net108893), .A1(net117709), .B0(net108894), .B1(
        net117731), .C0(net108895), .Y(net104957) );
  XOR2X4 U4772 ( .A(n4328), .B(n4329), .Y(n4323) );
  AOI22X4 U4773 ( .A0(net118215), .A1(net105167), .B0(net118225), .B1(
        net108579), .Y(net139866) );
  AO21X4 U4774 ( .A0(net105165), .A1(net105166), .B0(net117625), .Y(net105567)
         );
  AOI22X4 U4775 ( .A0(net118215), .A1(net104367), .B0(net118225), .B1(
        net107943), .Y(net139774) );
  OAI221X2 U4776 ( .A0(net107854), .A1(net117709), .B0(net107855), .B1(
        net117731), .C0(net107856), .Y(n4310) );
  CLKINVX3 U4777 ( .A(net104367), .Y(net107855) );
  XOR2X4 U4778 ( .A(n4322), .B(net108012), .Y(n4318) );
  INVX6 U4779 ( .A(n6488), .Y(n11026) );
  OR4X8 U4780 ( .A(n11595), .B(n11596), .C(n11597), .D(n11598), .Y(n4648) );
  AO22X4 U4781 ( .A0(n5135), .A1(n260), .B0(n5130), .B1(n429), .Y(n8352) );
  AND2X2 U4782 ( .A(n8635), .B(n126), .Y(n4726) );
  NAND2X1 U4783 ( .A(\i_MIPS/ALUin1[26] ), .B(n3973), .Y(n8635) );
  OAI221X2 U4784 ( .A0(n5324), .A1(n2024), .B0(n5353), .B1(n405), .C0(n6401), 
        .Y(n6402) );
  NAND4X4 U4785 ( .A(n8256), .B(n8255), .C(n8254), .D(n8253), .Y(n11420) );
  AOI21X4 U4786 ( .A0(n8719), .A1(n11101), .B0(n6813), .Y(n4739) );
  INVX3 U4787 ( .A(n8633), .Y(n6813) );
  NAND2X6 U4788 ( .A(\i_MIPS/ALUin1[23] ), .B(n4546), .Y(n8696) );
  OAI2BB1X4 U4789 ( .A0N(n9224), .A1N(n9223), .B0(n9222), .Y(n9227) );
  AO22X1 U4790 ( .A0(n5155), .A1(n218), .B0(n5151), .B1(n332), .Y(n6612) );
  AO22X1 U4791 ( .A0(n5154), .A1(n184), .B0(n5151), .B1(n304), .Y(n7125) );
  AO22X1 U4792 ( .A0(n5157), .A1(n185), .B0(n5151), .B1(n305), .Y(n7134) );
  AO22X1 U4793 ( .A0(n5157), .A1(n198), .B0(n5151), .B1(n306), .Y(n6894) );
  AO22X1 U4794 ( .A0(n5157), .A1(n199), .B0(n5151), .B1(n307), .Y(n7202) );
  AO22X1 U4795 ( .A0(n5157), .A1(n200), .B0(n5151), .B1(n308), .Y(n7211) );
  AO22X1 U4796 ( .A0(n5157), .A1(n216), .B0(n5151), .B1(n330), .Y(n6794) );
  AO22X1 U4797 ( .A0(n5154), .A1(n217), .B0(n5151), .B1(n331), .Y(n6803) );
  BUFX20 U4798 ( .A(n5221), .Y(n5214) );
  AO22X1 U4799 ( .A0(net118237), .A1(n771), .B0(net118255), .B1(n2363), .Y(
        n8580) );
  OA21X4 U4800 ( .A0(n3861), .A1(n5073), .B0(n7588), .Y(n6662) );
  BUFX16 U4801 ( .A(net117667), .Y(net117659) );
  CLKINVX4 U4802 ( .A(n11582), .Y(n8636) );
  AND2X4 U4803 ( .A(n6656), .B(net110423), .Y(n4700) );
  MX2XL U4804 ( .A(n3548), .B(net106031), .S0(n3595), .Y(\i_MIPS/n357 ) );
  AOI222X1 U4805 ( .A0(n5541), .A1(n11413), .B0(mem_rdata_D[37]), .B1(n129), 
        .C0(n13008), .C1(n5540), .Y(n10901) );
  OA21X4 U4806 ( .A0(\i_MIPS/ALUin1[5] ), .A1(n6712), .B0(\i_MIPS/ALUin1[4] ), 
        .Y(n4619) );
  OAI221X2 U4807 ( .A0(n5171), .A1(n2957), .B0(n5222), .B1(n1316), .C0(n6451), 
        .Y(n6452) );
  NAND4X4 U4808 ( .A(n8432), .B(n8431), .C(n8430), .D(n8429), .Y(n11396) );
  OA22X1 U4809 ( .A0(n5250), .A1(n980), .B0(n5290), .B1(n2605), .Y(n8431) );
  BUFX20 U4810 ( .A(n5186), .Y(n5174) );
  NAND2X4 U4811 ( .A(\i_MIPS/jump_addr[26] ), .B(n7739), .Y(n6769) );
  NAND2X8 U4812 ( .A(n6776), .B(n4723), .Y(net107168) );
  OA22X4 U4813 ( .A0(n5407), .A1(n2131), .B0(n5446), .B1(n506), .Y(n6441) );
  OAI221X2 U4814 ( .A0(n5326), .A1(n2025), .B0(n5354), .B1(n406), .C0(n6441), 
        .Y(n6442) );
  NAND2X4 U4815 ( .A(\i_MIPS/n202 ), .B(net144236), .Y(n4372) );
  MXI2X4 U4816 ( .A(n8293), .B(net134069), .S0(net114065), .Y(n4762) );
  CLKBUFX4 U4817 ( .A(net118243), .Y(net118237) );
  NAND2X8 U4818 ( .A(\i_MIPS/ALUin1[19] ), .B(n4578), .Y(n8683) );
  AO21X2 U4819 ( .A0(n8684), .A1(n8683), .B0(n8682), .Y(n8685) );
  OA22X4 U4820 ( .A0(n5246), .A1(n2057), .B0(n5278), .B1(n432), .Y(n9014) );
  OA22X4 U4821 ( .A0(n5246), .A1(n2134), .B0(n5296), .B1(n509), .Y(n8930) );
  OA22X4 U4822 ( .A0(n5246), .A1(n2136), .B0(n5296), .B1(n511), .Y(n9010) );
  OA22X4 U4823 ( .A0(n5256), .A1(n2137), .B0(n5298), .B1(n512), .Y(n7347) );
  BUFX20 U4824 ( .A(n5655), .Y(n5653) );
  OA22X1 U4825 ( .A0(n5653), .A1(n981), .B0(n5616), .B1(n2606), .Y(n11176) );
  OR4X8 U4826 ( .A(n11591), .B(n11592), .C(n11593), .D(n11594), .Y(n4650) );
  NAND2BX4 U4827 ( .AN(n9730), .B(net115797), .Y(n10736) );
  OAI211X2 U4828 ( .A0(n8668), .A1(n8667), .B0(n8666), .C0(n8665), .Y(n8669)
         );
  OA22X4 U4829 ( .A0(n5262), .A1(n2138), .B0(n5303), .B1(n513), .Y(n6414) );
  OAI211X2 U4830 ( .A0(n8863), .A1(n8293), .B0(n8292), .C0(n8861), .Y(n9132)
         );
  INVX4 U4831 ( .A(n8294), .Y(n8459) );
  OAI2BB2X4 U4832 ( .B0(n8462), .B1(net118601), .A0N(n8291), .A1N(net109496), 
        .Y(n8298) );
  AOI2BB1XL U4833 ( .A0N(n8639), .A1N(n8638), .B0(n4699), .Y(n8642) );
  AOI21X1 U4834 ( .A0(net108873), .A1(n3666), .B0(n8638), .Y(n4699) );
  XOR2X4 U4835 ( .A(ICACHE_addr[18]), .B(n11207), .Y(n11604) );
  INVX8 U4836 ( .A(n11360), .Y(n11207) );
  OA22X2 U4837 ( .A0(n5807), .A1(n4679), .B0(n5787), .B1(n3017), .Y(n11204) );
  OA22X4 U4838 ( .A0(n959), .A1(n5073), .B0(n3670), .B1(n5068), .Y(n7952) );
  NAND3BX4 U4839 ( .AN(n4819), .B(n7953), .C(n7952), .Y(n8037) );
  CLKBUFX2 U4840 ( .A(n4678), .Y(n5750) );
  OA22X4 U4841 ( .A0(n10307), .A1(n3766), .B0(n10310), .B1(n9536), .Y(n7920)
         );
  NAND4X2 U4842 ( .A(n7910), .B(n7909), .C(n7908), .D(n7907), .Y(n11462) );
  INVX3 U4843 ( .A(n11427), .Y(n10975) );
  CLKAND2X12 U4844 ( .A(n5043), .B(n11427), .Y(mem_wdata_D[51]) );
  AOI222X4 U4845 ( .A0(n5541), .A1(n11427), .B0(mem_rdata_D[51]), .B1(n132), 
        .C0(n12994), .C1(n5540), .Y(n10976) );
  NAND4X4 U4846 ( .A(n8346), .B(n8345), .C(n8344), .D(n8343), .Y(n11427) );
  NAND3BX4 U4847 ( .AN(n8471), .B(n7494), .C(n8044), .Y(n7765) );
  BUFX12 U4848 ( .A(n5197), .Y(n5223) );
  INVX8 U4849 ( .A(n11453), .Y(n10802) );
  NAND4X4 U4850 ( .A(n7995), .B(n7994), .C(n7993), .D(n7992), .Y(n11453) );
  AOI222X1 U4851 ( .A0(n5541), .A1(n11425), .B0(mem_rdata_D[49]), .B1(n132), 
        .C0(n12996), .C1(n5539), .Y(n10629) );
  CLKAND2X12 U4852 ( .A(n5044), .B(n11425), .Y(mem_wdata_D[49]) );
  OA22X2 U4853 ( .A0(n5831), .A1(n611), .B0(n5786), .B1(n2229), .Y(n11124) );
  NAND4X2 U4854 ( .A(n6684), .B(n6683), .C(n6682), .D(n6681), .Y(n6733) );
  CLKAND2X12 U4855 ( .A(net114065), .B(n3777), .Y(n4682) );
  NAND3BX4 U4856 ( .AN(n7239), .B(n7238), .C(n7237), .Y(net104503) );
  CLKBUFX2 U4857 ( .A(n5451), .Y(n5424) );
  CLKBUFX2 U4858 ( .A(n5451), .Y(n5425) );
  CLKBUFX2 U4859 ( .A(n5451), .Y(n5423) );
  XNOR2X4 U4860 ( .A(n6398), .B(DCACHE_addr[29]), .Y(n4366) );
  XNOR2X4 U4861 ( .A(n6413), .B(n12966), .Y(n4369) );
  BUFX20 U4862 ( .A(n5263), .Y(n5258) );
  NAND4X4 U4863 ( .A(n8428), .B(n8427), .C(n8426), .D(n8425), .Y(n11460) );
  OA22X1 U4864 ( .A0(n5174), .A1(n1241), .B0(n5213), .B1(n2860), .Y(n8428) );
  NOR2BX4 U4865 ( .AN(net105477), .B(\i_MIPS/n502 ), .Y(n4787) );
  AOI21X4 U4866 ( .A0(net108622), .A1(net108623), .B0(net108624), .Y(n4764) );
  NAND4X4 U4867 ( .A(n4656), .B(n4657), .C(n11212), .D(n11211), .Y(n11362) );
  OA22X4 U4868 ( .A0(n138), .A1(n2139), .B0(n5696), .B1(n514), .Y(n4657) );
  OA22X2 U4869 ( .A0(n5654), .A1(n612), .B0(n5608), .B1(n2230), .Y(n4656) );
  BUFX20 U4870 ( .A(n11056), .Y(n5555) );
  AOI2BB1X1 U4871 ( .A0N(\i_MIPS/PC/n19 ), .A1N(net115799), .B0(n10283), .Y(
        n10284) );
  NAND3X4 U4872 ( .A(n11603), .B(n11604), .C(n11605), .Y(n11599) );
  OA22X4 U4873 ( .A0(n5651), .A1(n2140), .B0(n5607), .B1(n515), .Y(n11117) );
  AO22X4 U4874 ( .A0(ICACHE_addr[19]), .A1(mem_read_I), .B0(mem_write_I), .B1(
        n11361), .Y(n12865) );
  NAND4X4 U4875 ( .A(n4655), .B(n11200), .C(n11199), .D(n11198), .Y(n11361) );
  OAI221X4 U4876 ( .A0(\i_MIPS/Register/register[2][25] ), .A1(net117635), 
        .B0(\i_MIPS/Register/register[10][25] ), .B1(net117653), .C0(n6876), 
        .Y(n6879) );
  BUFX20 U4877 ( .A(n4754), .Y(n5065) );
  BUFX20 U4878 ( .A(n5339), .Y(n5353) );
  AO21X4 U4879 ( .A0(n7123), .A1(n7122), .B0(n5191), .Y(net105256) );
  OA22X2 U4880 ( .A0(n10450), .A1(n3877), .B0(n10453), .B1(n4495), .Y(n7122)
         );
  NAND2X8 U4881 ( .A(n4503), .B(n1264), .Y(n8550) );
  OAI221X2 U4882 ( .A0(n5337), .A1(n2026), .B0(n5354), .B1(n407), .C0(n6493), 
        .Y(n6494) );
  AO21X4 U4883 ( .A0(net105009), .A1(net105008), .B0(net117727), .Y(net109841)
         );
  BUFX12 U4884 ( .A(n5300), .Y(n5293) );
  AOI2BB2X4 U4885 ( .B0(n3970), .B1(n9538), .A0N(n4983), .A1N(
        \i_MIPS/EX_MEM_1 ), .Y(n4982) );
  OAI221X2 U4886 ( .A0(n10699), .A1(n3767), .B0(n10702), .B1(n9536), .C0(n9535), .Y(n9538) );
  AO21X4 U4887 ( .A0(n8966), .A1(net108310), .B0(n8967), .Y(n9201) );
  AO22X4 U4888 ( .A0(n8965), .A1(n3674), .B0(n8964), .B1(n8963), .Y(n8967) );
  CLKAND2X12 U4889 ( .A(n10334), .B(net110470), .Y(n4786) );
  INVX4 U4890 ( .A(net105477), .Y(net110470) );
  OA22X1 U4891 ( .A0(n5395), .A1(n982), .B0(n5438), .B1(n2607), .Y(n7452) );
  BUFX20 U4892 ( .A(n5354), .Y(n5361) );
  BUFX20 U4893 ( .A(n3875), .Y(n5334) );
  MX2XL U4894 ( .A(n12959), .B(n4008), .S0(n3589), .Y(\i_MIPS/n373 ) );
  NOR4X4 U4895 ( .A(n8353), .B(n8352), .C(n8351), .D(n8350), .Y(n8354) );
  OA22X2 U4896 ( .A0(n8863), .A1(n8865), .B0(n6932), .B1(n8699), .Y(n6933) );
  OAI221X4 U4897 ( .A0(n300), .A1(n5072), .B0(n3744), .B1(n5067), .C0(n6840), 
        .Y(n6932) );
  INVX3 U4898 ( .A(n11444), .Y(n10750) );
  NAND4X4 U4899 ( .A(n9083), .B(n9082), .C(n9081), .D(n9080), .Y(n11476) );
  OA22X4 U4900 ( .A0(n5263), .A1(n2143), .B0(n5306), .B1(n518), .Y(n6426) );
  OA21X4 U4901 ( .A0(n2920), .A1(n5067), .B0(n8979), .Y(n7042) );
  NAND2X6 U4902 ( .A(n6708), .B(n2892), .Y(n7314) );
  OAI2BB1X2 U4903 ( .A0N(n7691), .A1N(n11097), .B0(n126), .Y(n9430) );
  INVX3 U4904 ( .A(n8635), .Y(n7691) );
  INVXL U4905 ( .A(n8211), .Y(n8212) );
  OA22X2 U4906 ( .A0(n10391), .A1(n3766), .B0(n10394), .B1(n9536), .Y(n7718)
         );
  NAND4X4 U4907 ( .A(n7708), .B(n7707), .C(n7706), .D(n7705), .Y(n11467) );
  OA22X2 U4908 ( .A0(n5180), .A1(n617), .B0(n5218), .B1(n2235), .Y(n7533) );
  OA22X2 U4909 ( .A0(n5180), .A1(n618), .B0(n5218), .B1(n2236), .Y(n7447) );
  NAND3BX2 U4910 ( .AN(n4745), .B(n8131), .C(n6657), .Y(n7583) );
  NAND3BX4 U4911 ( .AN(n7845), .B(n4718), .C(net114073), .Y(n8856) );
  INVX3 U4912 ( .A(n6471), .Y(n11042) );
  OA22X1 U4913 ( .A0(n5174), .A1(n983), .B0(n5213), .B1(n2608), .Y(n8519) );
  OA22X4 U4914 ( .A0(n5250), .A1(n2165), .B0(n5290), .B1(n546), .Y(n8427) );
  OAI221X4 U4915 ( .A0(n5169), .A1(n1304), .B0(n5209), .B1(n2990), .C0(n6392), 
        .Y(n10993) );
  AO21X4 U4916 ( .A0(n6752), .A1(n6751), .B0(n5192), .Y(net105312) );
  INVX8 U4917 ( .A(n11459), .Y(n10967) );
  NAND4X4 U4918 ( .A(n8338), .B(n8337), .C(n8336), .D(n8335), .Y(n11459) );
  OA22X2 U4919 ( .A0(n5376), .A1(n621), .B0(n5429), .B1(n2239), .Y(n8821) );
  NAND2X4 U4920 ( .A(n6712), .B(\i_MIPS/n296 ), .Y(n9298) );
  INVX2 U4921 ( .A(n8568), .Y(n8570) );
  AO21X4 U4922 ( .A0(n4710), .A1(n8566), .B0(n8565), .Y(n8568) );
  AO21X4 U4923 ( .A0(n5070), .A1(\i_MIPS/ALU/N303 ), .B0(n6842), .Y(n9314) );
  NAND2X2 U4924 ( .A(n6843), .B(n3674), .Y(n8041) );
  NAND2X4 U4925 ( .A(n3973), .B(n253), .Y(n7399) );
  AOI222X1 U4926 ( .A0(n5541), .A1(n11415), .B0(mem_rdata_D[39]), .B1(n132), 
        .C0(n13006), .C1(n5539), .Y(n10684) );
  NAND3BX4 U4927 ( .AN(n3634), .B(n11540), .C(n11343), .Y(n11346) );
  NAND2X4 U4928 ( .A(n3970), .B(n7836), .Y(n10111) );
  NAND2X2 U4929 ( .A(n5074), .B(n1264), .Y(n7104) );
  CLKMX2X4 U4930 ( .A(n6937), .B(n6936), .S0(\i_MIPS/ID_EX[81] ), .Y(n8855) );
  INVX8 U4931 ( .A(n11452), .Y(n10459) );
  NAND4X4 U4932 ( .A(n8248), .B(n8247), .C(n8246), .D(n8245), .Y(n11452) );
  BUFX3 U4933 ( .A(n5452), .Y(n5431) );
  OA22X4 U4934 ( .A0(n5394), .A1(n2167), .B0(n5431), .B1(n548), .Y(n8425) );
  NAND2X4 U4935 ( .A(n6610), .B(n4787), .Y(n4660) );
  BUFX20 U4936 ( .A(n5267), .Y(n5259) );
  OAI221X2 U4937 ( .A0(n1263), .A1(n5072), .B0(n2937), .B1(n5067), .C0(n7040), 
        .Y(n7680) );
  AOI2BB1X2 U4938 ( .A0N(n3670), .A1N(n3778), .B0(n4819), .Y(n7040) );
  NOR2BX4 U4939 ( .AN(n5066), .B(\i_MIPS/n287 ), .Y(n4819) );
  AO22X4 U4940 ( .A0(net118225), .A1(n7439), .B0(net105266), .B1(net118217), 
        .Y(net111041) );
  OAI222X2 U4941 ( .A0(n8114), .A1(n8113), .B0(n8203), .B1(n8112), .C0(n9316), 
        .C1(n8111), .Y(n8140) );
  NAND2X2 U4942 ( .A(net107652), .B(\i_MIPS/ID_EX[81] ), .Y(n8113) );
  INVX1 U4943 ( .A(n8863), .Y(n8963) );
  AO21X4 U4944 ( .A0(net105075), .A1(net105076), .B0(net117727), .Y(net111932)
         );
  OAI33X2 U4945 ( .A0(n3774), .A1(n7596), .A2(n7597), .B0(n7595), .B1(n7598), 
        .B2(n3774), .Y(n7606) );
  BUFX8 U4946 ( .A(n5197), .Y(n5224) );
  OA22X1 U4947 ( .A0(n5653), .A1(n984), .B0(n5616), .B1(n2609), .Y(n11186) );
  ACHCINX4 U4948 ( .CIN(n10567), .A(\i_MIPS/jump_addr[28] ), .B(n6016), .CO(
        n10578) );
  OAI211X2 U4949 ( .A0(\i_MIPS/IF_ID[20] ), .A1(n6016), .B0(n10332), .C0(
        n10331), .Y(n10350) );
  INVX20 U4950 ( .A(n5061), .Y(n5057) );
  BUFX20 U4951 ( .A(n4714), .Y(n5061) );
  OA22X2 U4952 ( .A0(n9316), .A1(n9201), .B0(net107988), .B1(n9205), .Y(n8972)
         );
  AOI32X2 U4953 ( .A0(n4000), .A1(n6646), .A2(n6645), .B0(n1340), .B1(n3873), 
        .Y(n6648) );
  OA22X4 U4954 ( .A0(n5652), .A1(n2146), .B0(n5585), .B1(n521), .Y(n11154) );
  NAND2X8 U4955 ( .A(n7102), .B(\i_MIPS/ID_EX[83] ), .Y(net107988) );
  AOI21X2 U4956 ( .A0(n8122), .A1(n3557), .B0(n8660), .Y(n4702) );
  OA22XL U4957 ( .A0(\i_MIPS/Register/register[6][23] ), .A1(n5081), .B0(
        \i_MIPS/Register/register[14][23] ), .B1(n5076), .Y(n7004) );
  OA22XL U4958 ( .A0(\i_MIPS/Register/register[6][6] ), .A1(n5081), .B0(
        \i_MIPS/Register/register[14][6] ), .B1(n5076), .Y(n7279) );
  BUFX20 U4959 ( .A(n5335), .Y(n5328) );
  CLKAND2X12 U4960 ( .A(n5951), .B(n11265), .Y(mem_wdata_I[47]) );
  OA22X2 U4961 ( .A0(n5334), .A1(n623), .B0(n5361), .B1(n2241), .Y(n7346) );
  BUFX20 U4962 ( .A(n5304), .Y(n5303) );
  BUFX20 U4963 ( .A(n5312), .Y(n5304) );
  AO21X4 U4964 ( .A0(n7920), .A1(n7919), .B0(n4626), .Y(net105491) );
  OA22X4 U4965 ( .A0(n10548), .A1(n3877), .B0(n10551), .B1(n4495), .Y(n7627)
         );
  INVX3 U4966 ( .A(n11436), .Y(n10551) );
  CLKAND2X12 U4967 ( .A(n5043), .B(n11436), .Y(mem_wdata_D[60]) );
  BUFX20 U4968 ( .A(n5183), .Y(n5181) );
  XNOR2X4 U4969 ( .A(ICACHE_addr[11]), .B(n11353), .Y(n11135) );
  AO22X4 U4970 ( .A0(n8463), .A1(n8462), .B0(n8461), .B1(net109196), .Y(n8474)
         );
  INVX8 U4971 ( .A(n11463), .Y(n10689) );
  AOI222X1 U4972 ( .A0(n4505), .A1(n11463), .B0(mem_rdata_D[87]), .B1(n130), 
        .C0(n12990), .C1(n5536), .Y(n10690) );
  NAND4X4 U4973 ( .A(n7068), .B(n7067), .C(n7066), .D(n7065), .Y(n11463) );
  MXI2X4 U4974 ( .A(\i_MIPS/ID_EX[113] ), .B(\i_MIPS/ID_EX[86] ), .S0(
        \i_MIPS/ID_EX_5 ), .Y(n6754) );
  INVX4 U4975 ( .A(n6754), .Y(n10849) );
  NAND4BX4 U4976 ( .AN(n4652), .B(n11158), .C(n11157), .D(n11156), .Y(n11350)
         );
  OAI22X1 U4977 ( .A0(n5653), .A1(n559), .B0(n5607), .B1(n2180), .Y(n4652) );
  NOR4X4 U4978 ( .A(n8362), .B(n8361), .C(n8360), .D(n8359), .Y(n8363) );
  BUFX20 U4979 ( .A(n5140), .Y(n5144) );
  NOR3X8 U4980 ( .A(n4648), .B(n4649), .C(n4650), .Y(n6387) );
  AOI222X4 U4981 ( .A0(n9445), .A1(n7586), .B0(net134673), .B1(n7594), .C0(
        n4715), .C1(n9442), .Y(n7610) );
  MX2X2 U4982 ( .A(n8865), .B(n8975), .S0(net114065), .Y(n8866) );
  AOI222X4 U4983 ( .A0(n3800), .A1(n11388), .B0(mem_rdata_D[12]), .B1(n129), 
        .C0(n13001), .C1(n5537), .Y(n10463) );
  AOI32X4 U4984 ( .A0(n9431), .A1(n6960), .A2(net117743), .B0(n4733), .B1(
        n11113), .Y(n6957) );
  NAND4X4 U4985 ( .A(n11196), .B(n11195), .C(n11194), .D(n11193), .Y(n11367)
         );
  NAND4X6 U4986 ( .A(n7618), .B(n7617), .C(n7616), .D(n7615), .Y(n11468) );
  OA22X4 U4987 ( .A0(n5333), .A1(n2150), .B0(n5360), .B1(n525), .Y(n7616) );
  AO21X4 U4988 ( .A0(n8348), .A1(n8347), .B0(n4626), .Y(net105663) );
  NAND2X4 U4989 ( .A(n3776), .B(n4732), .Y(n6923) );
  NAND2X4 U4990 ( .A(n9935), .B(ICACHE_addr[2]), .Y(n10051) );
  AOI222X1 U4991 ( .A0(n4534), .A1(n11494), .B0(mem_rdata_D[118]), .B1(n133), 
        .C0(n12991), .C1(n5533), .Y(n10308) );
  OR4X8 U4992 ( .A(n11599), .B(n11600), .C(n11601), .D(n11602), .Y(n4649) );
  OA22X1 U4993 ( .A0(n5653), .A1(n985), .B0(n5607), .B1(n2610), .Y(n11171) );
  OAI221X2 U4994 ( .A0(net107689), .A1(n7234), .B0(n7151), .B1(n9318), .C0(
        n7150), .Y(n7164) );
  OA21X4 U4995 ( .A0(n8574), .A1(n3967), .B0(n8572), .Y(n4633) );
  OAI211X2 U4996 ( .A0(n9438), .A1(n9437), .B0(n9436), .C0(n9435), .Y(n9439)
         );
  OA22XL U4997 ( .A0(n5333), .A1(n1278), .B0(n5358), .B1(n2910), .Y(n9178) );
  OAI211X2 U4998 ( .A0(\i_MIPS/IF_ID[23] ), .A1(n6016), .B0(n10363), .C0(
        n10362), .Y(n10373) );
  NAND3BX4 U4999 ( .AN(n4821), .B(n4804), .C(n10350), .Y(n10362) );
  INVX8 U5000 ( .A(n4546), .Y(n6686) );
  AO21X4 U5001 ( .A0(net104889), .A1(net104890), .B0(net117727), .Y(net111130)
         );
  BUFX12 U5002 ( .A(n5220), .Y(n5218) );
  AOI221X2 U5003 ( .A0(n7310), .A1(n7309), .B0(n7308), .B1(n7307), .C0(n7306), 
        .Y(n7318) );
  NAND2X4 U5004 ( .A(n4692), .B(n9301), .Y(n7488) );
  OA22X1 U5005 ( .A0(n5175), .A1(n1242), .B0(n5214), .B1(n2861), .Y(n8748) );
  OAI222X4 U5006 ( .A0(net107217), .A1(n7424), .B0(n7482), .B1(n9206), .C0(
        net117757), .C1(n7432), .Y(n7425) );
  INVX4 U5007 ( .A(n11417), .Y(n10615) );
  NAND4X2 U5008 ( .A(n8086), .B(n8085), .C(n8084), .D(n8083), .Y(n11417) );
  AO21X4 U5009 ( .A0(n8529), .A1(n8528), .B0(n4626), .Y(net119104) );
  CLKBUFX2 U5010 ( .A(n4677), .Y(n5840) );
  CLKINVX4 U5011 ( .A(n7771), .Y(n6656) );
  NAND2X4 U5012 ( .A(n8211), .B(n7956), .Y(n7771) );
  AO21X4 U5013 ( .A0(n7718), .A1(n7717), .B0(n5191), .Y(net105424) );
  OAI221X4 U5014 ( .A0(n10592), .A1(n3766), .B0(n10595), .B1(n5189), .C0(n9420), .Y(n9421) );
  OA22X4 U5015 ( .A0(n10598), .A1(n3879), .B0(n10601), .B1(n4495), .Y(n9420)
         );
  OAI221X4 U5016 ( .A0(n336), .A1(n5071), .B0(n1264), .B1(n5067), .C0(n8110), 
        .Y(n8700) );
  XOR2X4 U5017 ( .A(n11355), .B(ICACHE_addr[13]), .Y(n11598) );
  NAND4X4 U5018 ( .A(n11181), .B(n11180), .C(n11179), .D(n11178), .Y(n11355)
         );
  NAND2X4 U5019 ( .A(\i_MIPS/ALUin1[9] ), .B(n6702), .Y(n8666) );
  NAND4X4 U5020 ( .A(n8078), .B(n8077), .C(n8076), .D(n8075), .Y(n11449) );
  OA22X2 U5021 ( .A0(n5331), .A1(n712), .B0(n5359), .B1(n2334), .Y(n8076) );
  OAI2BB1X4 U5022 ( .A0N(net108847), .A1N(net108010), .B0(n9121), .Y(n8651) );
  AOI31X2 U5023 ( .A0(n8677), .A1(n8676), .A2(n8675), .B0(n8674), .Y(n8718) );
  CLKAND2X12 U5024 ( .A(n5047), .B(n11338), .Y(mem_wdata_I[123]) );
  AOI21X2 U5025 ( .A0(n6728), .A1(n8890), .B0(n6727), .Y(n6730) );
  AOI2BB2X4 U5026 ( .B0(n7500), .B1(n7499), .A0N(n7498), .A1N(n7497), .Y(n7501) );
  NAND3BX4 U5027 ( .AN(n8140), .B(n8139), .C(n8138), .Y(net104941) );
  BUFX20 U5028 ( .A(n5221), .Y(n5217) );
  BUFX20 U5029 ( .A(n5179), .Y(n5178) );
  BUFX20 U5030 ( .A(n5225), .Y(n5219) );
  OAI221X2 U5031 ( .A0(n5185), .A1(n2027), .B0(n5210), .B1(n408), .C0(n6404), 
        .Y(n6405) );
  OAI221X2 U5032 ( .A0(n3875), .A1(n412), .B0(n5354), .B1(n256), .C0(n6406), 
        .Y(n6407) );
  OAI222X4 U5033 ( .A0(n9550), .A1(n9208), .B0(n9202), .B1(n8035), .C0(n9206), 
        .C1(n8041), .Y(n6844) );
  OAI221X4 U5034 ( .A0(n343), .A1(n5064), .B0(n2920), .B1(n5056), .C0(n6833), 
        .Y(n8873) );
  OA21X2 U5035 ( .A0(n1302), .A1(n5073), .B0(n8980), .Y(n6833) );
  OA22X4 U5036 ( .A0(n10661), .A1(n3767), .B0(n10664), .B1(n9536), .Y(n9021)
         );
  MXI2X4 U5037 ( .A(n10665), .B(n10664), .S0(n5548), .Y(n10666) );
  INVX3 U5038 ( .A(n11441), .Y(n10664) );
  AOI211X4 U5039 ( .A0(n8976), .A1(n7590), .B0(net107841), .C0(n7589), .Y(
        n7609) );
  XOR2X4 U5040 ( .A(n11359), .B(ICACHE_addr[17]), .Y(n11594) );
  INVX8 U5041 ( .A(n11445), .Y(n10894) );
  NAND4X4 U5042 ( .A(n9353), .B(n9352), .C(n9351), .D(n9350), .Y(n11445) );
  AO21X4 U5043 ( .A0(net105142), .A1(net105143), .B0(net117723), .Y(n8958) );
  NAND4BX4 U5044 ( .AN(n4651), .B(n11121), .C(n11120), .D(n11119), .Y(n11353)
         );
  AOI32X2 U5045 ( .A0(net117743), .A1(n6826), .A2(n7405), .B0(n4701), .B1(
        n6825), .Y(n6852) );
  OAI211X2 U5046 ( .A0(n6964), .A1(n6963), .B0(n6962), .C0(n6961), .Y(
        net105077) );
  OR2X1 U5047 ( .A(n5557), .B(n10346), .Y(n4422) );
  OR2X1 U5048 ( .A(n5558), .B(n10382), .Y(n4418) );
  OR2XL U5049 ( .A(n5557), .B(n10369), .Y(n4416) );
  AOI211X2 U5050 ( .A0(n8215), .A1(net109168), .B0(n8214), .C0(n8213), .Y(
        n8216) );
  NAND4BX4 U5051 ( .AN(n4644), .B(n11130), .C(n11129), .D(n11128), .Y(n11357)
         );
  OAI222X1 U5052 ( .A0(net107217), .A1(net110406), .B0(n9451), .B1(net107661), 
        .C0(n351), .C1(net117757), .Y(n7792) );
  OAI221X4 U5053 ( .A0(\i_MIPS/n296 ), .A1(n5063), .B0(n1302), .B1(n5057), 
        .C0(n7232), .Y(n7788) );
  OAI31X2 U5054 ( .A0(n7), .A1(n9428), .A2(n9427), .B0(n9426), .Y(n9542) );
  OAI2BB1X2 U5055 ( .A0N(n9304), .A1N(n9303), .B0(net107680), .Y(n9305) );
  NAND4BX4 U5056 ( .AN(net109513), .B(n3857), .C(n8282), .D(net109510), .Y(
        n8779) );
  OAI221X2 U5057 ( .A0(n5186), .A1(n2028), .B0(n5210), .B1(n409), .C0(n6409), 
        .Y(n6410) );
  NAND4BX2 U5058 ( .AN(\i_MIPS/ID_EX[106] ), .B(\i_MIPS/ID_EX[105] ), .C(
        \i_MIPS/ID_EX[107] ), .D(n4672), .Y(\i_MIPS/ALU_Control/n20 ) );
  OAI21X4 U5059 ( .A0(n4834), .A1(net112555), .B0(n1340), .Y(n6644) );
  AOI222X2 U5060 ( .A0(n4688), .A1(net107992), .B0(n9546), .B1(n8976), .C0(
        n7676), .C1(n8294), .Y(n7677) );
  AOI211X4 U5061 ( .A0(net107652), .A1(n4763), .B0(n7236), .C0(n7235), .Y(
        n7237) );
  AO21X4 U5062 ( .A0(n8834), .A1(n8833), .B0(n4626), .Y(net105166) );
  NAND3BX4 U5063 ( .AN(n9325), .B(n9323), .C(n9324), .Y(net104752) );
  OAI31X2 U5064 ( .A0(n8470), .A1(n8469), .A2(n8468), .B0(n8467), .Y(n8479) );
  OAI221X4 U5065 ( .A0(n5185), .A1(n1337), .B0(n5210), .B1(n2991), .C0(n6414), 
        .Y(n6415) );
  OAI221X2 U5066 ( .A0(n3875), .A1(n413), .B0(n5354), .B1(n257), .C0(n6411), 
        .Y(n6412) );
  BUFX20 U5067 ( .A(n5183), .Y(n5182) );
  OA22X4 U5068 ( .A0(n5406), .A1(n2153), .B0(n5445), .B1(n528), .Y(n6475) );
  AO21X4 U5069 ( .A0(n6871), .A1(n6870), .B0(n5192), .Y(net105289) );
  OAI221X4 U5070 ( .A0(n10828), .A1(n5560), .B0(ICACHE_addr[0]), .B1(n5557), 
        .C0(n10827), .Y(\i_MIPS/PC/n36 ) );
  AOI211X2 U5071 ( .A0(net107652), .A1(n8710), .B0(n8709), .C0(n8708), .Y(
        n8711) );
  OAI221X2 U5072 ( .A0(n5169), .A1(n1938), .B0(n5209), .B1(n353), .C0(n6399), 
        .Y(n6400) );
  AO21X4 U5073 ( .A0(n7078), .A1(n7077), .B0(n5191), .Y(net104867) );
  OA22X2 U5074 ( .A0(n5917), .A1(n628), .B0(n5875), .B1(n2982), .Y(n11114) );
  CLKAND2X12 U5075 ( .A(n5047), .B(n11341), .Y(mem_wdata_I[126]) );
  BUFX20 U5076 ( .A(n5448), .Y(n5446) );
  OA22X4 U5077 ( .A0(n10784), .A1(n3767), .B0(n10787), .B1(n9536), .Y(n8529)
         );
  BUFX20 U5078 ( .A(n5338), .Y(n5335) );
  XOR2X4 U5079 ( .A(n6455), .B(DCACHE_addr[18]), .Y(n6456) );
  CLKINVX20 U5080 ( .A(n5044), .Y(n5040) );
  OAI211X4 U5081 ( .A0(\i_MIPS/ALUin1[15] ), .A1(n5068), .B0(n7299), .C0(n6839), .Y(n6936) );
  OAI211X2 U5082 ( .A0(n8471), .A1(n8467), .B0(n7959), .C0(n8464), .Y(n8200)
         );
  CLKAND2X12 U5083 ( .A(n5947), .B(n11376), .Y(mem_wdata_D[0]) );
  AOI2BB1X1 U5084 ( .A0N(\i_MIPS/ALUin1[14] ), .A1N(n3778), .B0(n4730), .Y(
        n7157) );
  NAND2X4 U5085 ( .A(n10138), .B(n4800), .Y(n10146) );
  CLKAND2X12 U5086 ( .A(n5043), .B(n11442), .Y(mem_wdata_D[66]) );
  NAND2X6 U5087 ( .A(n4376), .B(n4377), .Y(net144227) );
  INVXL U5088 ( .A(\i_MIPS/ID_EX[81] ), .Y(net144224) );
  OAI221X4 U5089 ( .A0(n344), .A1(n5064), .B0(n183), .B1(n5056), .C0(n7030), 
        .Y(n8462) );
  OAI221X4 U5090 ( .A0(\i_MIPS/n271 ), .A1(n5072), .B0(n2961), .B1(n5068), 
        .C0(n7031), .Y(n8293) );
  OAI2BB1X4 U5091 ( .A0N(net135772), .A1N(n3674), .B0(n7419), .Y(n7312) );
  NAND2X2 U5092 ( .A(n4505), .B(n11447), .Y(n4380) );
  NAND2XL U5093 ( .A(mem_rdata_D[71]), .B(n132), .Y(n4381) );
  NAND2XL U5094 ( .A(n13006), .B(n5536), .Y(n4382) );
  NAND4X4 U5095 ( .A(n7348), .B(n7347), .C(n7346), .D(n7345), .Y(n11447) );
  MXI2X4 U5096 ( .A(n10678), .B(n10677), .S0(n5548), .Y(n10679) );
  AND2XL U5097 ( .A(mem_rdata_D[97]), .B(n131), .Y(n4384) );
  AND2XL U5098 ( .A(n13012), .B(n5534), .Y(n4385) );
  AND2X2 U5099 ( .A(mem_rdata_D[66]), .B(n130), .Y(n4387) );
  NAND4X4 U5100 ( .A(n7192), .B(n7191), .C(n7190), .D(n7189), .Y(n11442) );
  AND2X4 U5101 ( .A(n4534), .B(n11475), .Y(n4389) );
  AND2X1 U5102 ( .A(mem_rdata_D[99]), .B(n130), .Y(n4390) );
  AND2X1 U5103 ( .A(n13010), .B(n5533), .Y(n4391) );
  NOR3X2 U5104 ( .A(n4389), .B(n4390), .C(n4391), .Y(n9800) );
  MXI2X1 U5105 ( .A(n9800), .B(n9799), .S0(n5542), .Y(n10758) );
  CLKAND2X3 U5106 ( .A(n13007), .B(n5539), .Y(n4394) );
  NOR3X4 U5107 ( .A(n4392), .B(n4393), .C(n4394), .Y(n9961) );
  MXI2X1 U5108 ( .A(n9961), .B(n9960), .S0(n5542), .Y(n9962) );
  NAND2X4 U5109 ( .A(n7222), .B(\i_MIPS/n296 ), .Y(n9308) );
  AND2XL U5110 ( .A(n5051), .B(\i_MIPS/ALU/N303 ), .Y(n4397) );
  OR2X8 U5111 ( .A(n4397), .B(n6842), .Y(n8862) );
  AO21X4 U5112 ( .A0(n5062), .A1(\i_MIPS/ALUin1[29] ), .B0(n4810), .Y(n6842)
         );
  OAI221X4 U5113 ( .A0(n5073), .A1(\i_MIPS/n301 ), .B0(\i_MIPS/n300 ), .B1(
        n5068), .C0(n7037), .Y(net107992) );
  AO22X1 U5114 ( .A0(net109168), .A1(n8482), .B0(net134673), .B1(n8481), .Y(
        n8483) );
  NAND2X4 U5115 ( .A(n7278), .B(n7277), .Y(n4406) );
  NAND2X8 U5116 ( .A(n4406), .B(n4407), .Y(net106298) );
  INVX4 U5117 ( .A(n11395), .Y(n10971) );
  OR2X1 U5118 ( .A(n10495), .B(n5560), .Y(n4413) );
  NAND3X2 U5119 ( .A(n4415), .B(n4416), .C(n10367), .Y(\i_MIPS/PC/n58 ) );
  NAND3X2 U5120 ( .A(n4417), .B(n4418), .C(n10380), .Y(\i_MIPS/PC/n60 ) );
  XOR2X2 U5121 ( .A(n10377), .B(ICACHE_addr[24]), .Y(n10382) );
  OR2X1 U5122 ( .A(n10535), .B(n5560), .Y(n4419) );
  XOR2X2 U5123 ( .A(n10532), .B(ICACHE_addr[26]), .Y(n10536) );
  AOI2BB1X1 U5124 ( .A0N(\i_MIPS/PC/n30 ), .A1N(net115789), .B0(n10533), .Y(
        n10534) );
  NAND3X2 U5125 ( .A(n4421), .B(n4422), .C(n10344), .Y(\i_MIPS/PC/n56 ) );
  OR2X1 U5126 ( .A(n9735), .B(n5560), .Y(n4423) );
  NAND3X2 U5127 ( .A(n4423), .B(n4424), .C(n9733), .Y(\i_MIPS/PC/n37 ) );
  NOR3X2 U5128 ( .A(n4461), .B(n4462), .C(n4463), .Y(n9630) );
  NOR3X2 U5129 ( .A(n4464), .B(n4466), .C(n4465), .Y(n10960) );
  NOR3X2 U5130 ( .A(n4467), .B(n4469), .C(n4468), .Y(n9682) );
  AND2X1 U5131 ( .A(net104172), .B(n11255), .Y(n4478) );
  NOR3X2 U5132 ( .A(n4490), .B(n4491), .C(n4492), .Y(n9652) );
  OR2X1 U5133 ( .A(n7420), .B(net118601), .Y(n4493) );
  NAND3X2 U5134 ( .A(n4493), .B(n4494), .C(n7419), .Y(n7481) );
  INVX3 U5135 ( .A(n7481), .Y(n7421) );
  INVX20 U5136 ( .A(n4059), .Y(n4495) );
  MXI2X4 U5137 ( .A(\i_MIPS/ID_EX[115] ), .B(\i_MIPS/ID_EX[88] ), .S0(
        \i_MIPS/ID_EX_5 ), .Y(n6633) );
  AOI2BB1X1 U5138 ( .A0N(\i_MIPS/PC/n18 ), .A1N(net115799), .B0(n10274), .Y(
        n10275) );
  AOI2BB1X1 U5139 ( .A0N(\i_MIPS/PC/n12 ), .A1N(net115789), .B0(n10169), .Y(
        n10170) );
  AOI2BB1X1 U5140 ( .A0N(\i_MIPS/PC/n31 ), .A1N(net115789), .B0(n10570), .Y(
        n10571) );
  AOI2BB1X1 U5141 ( .A0N(\i_MIPS/PC/n14 ), .A1N(net115799), .B0(n10474), .Y(
        n10475) );
  AOI2BB1X1 U5142 ( .A0N(\i_MIPS/PC/n15 ), .A1N(net115789), .B0(n10482), .Y(
        n10483) );
  OAI221X2 U5143 ( .A0(n5328), .A1(n2029), .B0(n5353), .B1(n410), .C0(n6470), 
        .Y(n6471) );
  OAI221X4 U5144 ( .A0(n5187), .A1(n1338), .B0(n5222), .B1(n2992), .C0(n6487), 
        .Y(n6488) );
  OAI221X2 U5145 ( .A0(n5170), .A1(n2354), .B0(n5212), .B1(n904), .C0(n6448), 
        .Y(n6449) );
  OAI221X2 U5146 ( .A0(n5328), .A1(n414), .B0(n5353), .B1(n258), .C0(n6475), 
        .Y(n6476) );
  CLKAND2X12 U5147 ( .A(n5947), .B(n11377), .Y(mem_wdata_D[1]) );
  AO21X4 U5148 ( .A0(n9272), .A1(n9271), .B0(n4626), .Y(net119263) );
  AO21X4 U5149 ( .A0(n9453), .A1(net108310), .B0(n3631), .Y(n8555) );
  NAND4BX4 U5150 ( .AN(n8983), .B(n8982), .C(n8981), .D(net108281), .Y(
        net104918) );
  AO21X4 U5151 ( .A0(n8005), .A1(n8004), .B0(n4626), .Y(net104699) );
  AO21X4 U5152 ( .A0(n8968), .A1(net108310), .B0(n8967), .Y(n9205) );
  OA22X2 U5153 ( .A0(n10313), .A1(n3879), .B0(n10316), .B1(n4495), .Y(n7919)
         );
  CLKINVX20 U5154 ( .A(n5027), .Y(mem_addr_D[23]) );
  INVX4 U5155 ( .A(n5011), .Y(n5027) );
  CLKINVX20 U5156 ( .A(n5031), .Y(mem_addr_D[25]) );
  INVX4 U5157 ( .A(n5013), .Y(n5031) );
  CLKINVX20 U5158 ( .A(n5033), .Y(mem_addr_D[27]) );
  INVX4 U5159 ( .A(n5015), .Y(n5033) );
  CLKINVX20 U5160 ( .A(n5035), .Y(mem_addr_D[28]) );
  INVX4 U5161 ( .A(n5016), .Y(n5035) );
  CLKINVX20 U5162 ( .A(n5038), .Y(mem_addr_D[30]) );
  INVX4 U5163 ( .A(n5018), .Y(n5038) );
  CLKINVX20 U5164 ( .A(n5039), .Y(mem_addr_D[31]) );
  INVX4 U5165 ( .A(n5019), .Y(n5039) );
  CLKINVX20 U5166 ( .A(n5028), .Y(mem_addr_D[24]) );
  INVX4 U5167 ( .A(n5012), .Y(n5028) );
  CLKINVX20 U5168 ( .A(n5032), .Y(mem_addr_D[26]) );
  INVX4 U5169 ( .A(n5014), .Y(n5032) );
  CLKINVX20 U5170 ( .A(n5037), .Y(mem_addr_D[29]) );
  INVX4 U5171 ( .A(n5017), .Y(n5037) );
  AO22X4 U5172 ( .A0(net108148), .A1(net117747), .B0(net135551), .B1(n9124), 
        .Y(n7147) );
  AOI2BB1X4 U5173 ( .A0N(n8658), .A1N(n8659), .B0(n8657), .Y(n8661) );
  OAI221X2 U5174 ( .A0(n5325), .A1(n906), .B0(n5353), .B1(n299), .C0(n6428), 
        .Y(n6429) );
  AO21X4 U5175 ( .A0(n8088), .A1(n8087), .B0(n5026), .Y(net105009) );
  AO21X4 U5176 ( .A0(n7628), .A1(n7627), .B0(n5026), .Y(net105111) );
  AO21X4 U5177 ( .A0(n7457), .A1(n7456), .B0(n4626), .Y(net105265) );
  BUFX8 U5178 ( .A(n10795), .Y(n4500) );
  BUFX8 U5179 ( .A(n10782), .Y(n4501) );
  AO22X4 U5180 ( .A0(n5062), .A1(\i_MIPS/ALUin1[1] ), .B0(\i_MIPS/ALUin1[0] ), 
        .B1(n5065), .Y(n8975) );
  BUFX8 U5181 ( .A(n10402), .Y(n4511) );
  BUFX8 U5182 ( .A(n10428), .Y(n4512) );
  BUFX8 U5183 ( .A(n10415), .Y(n4513) );
  BUFX8 U5184 ( .A(n10425), .Y(n4517) );
  BUFX8 U5185 ( .A(n10412), .Y(n4518) );
  BUFX8 U5186 ( .A(n10507), .Y(n4519) );
  BUFX8 U5187 ( .A(n10464), .Y(n4521) );
  BUFX8 U5188 ( .A(n10399), .Y(n4522) );
  BUFX8 U5189 ( .A(n10206), .Y(n4523) );
  BUFX8 U5190 ( .A(n10109), .Y(n4525) );
  BUFX8 U5191 ( .A(n9962), .Y(n4526) );
  BUFX8 U5192 ( .A(n10106), .Y(n4527) );
  BUFX8 U5193 ( .A(n9955), .Y(n4528) );
  AO21X4 U5194 ( .A0(n8258), .A1(n8257), .B0(n5026), .Y(net105233) );
  BUFX8 U5195 ( .A(n10893), .Y(n4537) );
  BUFX8 U5196 ( .A(n10786), .Y(n4542) );
  INVX3 U5197 ( .A(n8379), .Y(n6659) );
  OAI221X4 U5198 ( .A0(n2920), .A1(n5071), .B0(n300), .B1(n5068), .C0(n6658), 
        .Y(n8379) );
  BUFX8 U5199 ( .A(n10449), .Y(n4551) );
  BUFX8 U5200 ( .A(n10594), .Y(n4571) );
  BUFX8 U5201 ( .A(n10557), .Y(n4572) );
  BUFX8 U5202 ( .A(n10544), .Y(n4573) );
  BUFX8 U5203 ( .A(n10458), .Y(n4575) );
  AO21X4 U5204 ( .A0(n9363), .A1(n9362), .B0(n5191), .Y(net106038) );
  OAI31X2 U5205 ( .A0(net110424), .A1(n7777), .A2(n7776), .B0(net108873), .Y(
        n7780) );
  AOI2BB1X2 U5206 ( .A0N(n9140), .A1N(n3752), .B0(n9139), .Y(n9141) );
  OAI222X1 U5207 ( .A0(n9550), .A1(n8792), .B0(net107988), .B1(n8133), .C0(
        n8697), .C1(net107977), .Y(n8136) );
  CLKMX2X2 U5208 ( .A(n3544), .B(n3944), .S0(n3591), .Y(\i_MIPS/n327 ) );
  AO21X4 U5209 ( .A0(net105288), .A1(net105289), .B0(net117727), .Y(net112120)
         );
  OAI221X2 U5210 ( .A0(n3970), .A1(n4796), .B0(mem_ready_D), .B1(n3789), .C0(
        n9797), .Y(n9957) );
  AOI21X4 U5211 ( .A0(n8565), .A1(n8681), .B0(n8644), .Y(n4687) );
  OAI221X2 U5212 ( .A0(n5326), .A1(n2355), .B0(n5352), .B1(n905), .C0(n6437), 
        .Y(n6438) );
  AO22X1 U5213 ( .A0(n12957), .A1(mem_read_D), .B0(mem_write_D), .B1(n11530), 
        .Y(n5016) );
  CLKINVX8 U5214 ( .A(n12878), .Y(n4581) );
  INVX20 U5215 ( .A(n4581), .Y(mem_addr_I[7]) );
  CLKAND2X12 U5216 ( .A(ICACHE_addr[2]), .B(n11345), .Y(mem_addr_I[4]) );
  INVX12 U5217 ( .A(\i_MIPS/n245 ), .Y(DCACHE_wen) );
  NAND2XL U5218 ( .A(n12963), .B(\i_MIPS/n266 ), .Y(net105490) );
  AO22X2 U5219 ( .A0(n4757), .A1(n12963), .B0(n5552), .B1(n11524), .Y(n11035)
         );
  INVX12 U5220 ( .A(\i_MIPS/n181 ), .Y(DCACHE_wdata[31]) );
  INVX12 U5221 ( .A(\i_MIPS/n183 ), .Y(DCACHE_wdata[30]) );
  INVX12 U5222 ( .A(\i_MIPS/n185 ), .Y(DCACHE_wdata[29]) );
  INVX12 U5223 ( .A(\i_MIPS/n187 ), .Y(DCACHE_wdata[28]) );
  INVX12 U5224 ( .A(\i_MIPS/n195 ), .Y(DCACHE_wdata[24]) );
  INVX12 U5225 ( .A(\i_MIPS/n197 ), .Y(DCACHE_wdata[23]) );
  INVX12 U5226 ( .A(\i_MIPS/n201 ), .Y(DCACHE_wdata[21]) );
  INVX12 U5227 ( .A(\i_MIPS/n207 ), .Y(DCACHE_wdata[18]) );
  INVX12 U5228 ( .A(\i_MIPS/n209 ), .Y(DCACHE_wdata[17]) );
  INVX12 U5229 ( .A(\i_MIPS/n215 ), .Y(DCACHE_wdata[14]) );
  INVX12 U5230 ( .A(\i_MIPS/n217 ), .Y(DCACHE_wdata[13]) );
  INVX12 U5231 ( .A(\i_MIPS/n223 ), .Y(DCACHE_wdata[10]) );
  INVX12 U5232 ( .A(\i_MIPS/n225 ), .Y(DCACHE_wdata[9]) );
  INVX12 U5233 ( .A(\i_MIPS/n227 ), .Y(DCACHE_wdata[8]) );
  INVX12 U5234 ( .A(\i_MIPS/n229 ), .Y(DCACHE_wdata[7]) );
  INVX12 U5235 ( .A(\i_MIPS/n235 ), .Y(DCACHE_wdata[4]) );
  INVX12 U5236 ( .A(\i_MIPS/n241 ), .Y(DCACHE_wdata[1]) );
  INVX12 U5237 ( .A(\i_MIPS/n239 ), .Y(DCACHE_wdata[2]) );
  INVX12 U5238 ( .A(\i_MIPS/n233 ), .Y(DCACHE_wdata[5]) );
  INVX12 U5239 ( .A(\i_MIPS/n237 ), .Y(DCACHE_wdata[3]) );
  INVX12 U5240 ( .A(\i_MIPS/n213 ), .Y(DCACHE_wdata[15]) );
  INVX12 U5241 ( .A(\i_MIPS/n243 ), .Y(DCACHE_wdata[0]) );
  INVX12 U5242 ( .A(\i_MIPS/n189 ), .Y(DCACHE_wdata[27]) );
  INVX12 U5243 ( .A(\i_MIPS/n211 ), .Y(DCACHE_wdata[16]) );
  INVX12 U5244 ( .A(\i_MIPS/n193 ), .Y(DCACHE_wdata[25]) );
  INVX12 U5245 ( .A(\i_MIPS/n199 ), .Y(DCACHE_wdata[22]) );
  INVX12 U5246 ( .A(\i_MIPS/n221 ), .Y(DCACHE_wdata[11]) );
  INVX12 U5247 ( .A(\i_MIPS/n231 ), .Y(DCACHE_wdata[6]) );
  INVX12 U5248 ( .A(\i_MIPS/n219 ), .Y(DCACHE_wdata[12]) );
  INVX12 U5249 ( .A(\i_MIPS/n191 ), .Y(DCACHE_wdata[26]) );
  INVX12 U5250 ( .A(\i_MIPS/n203 ), .Y(DCACHE_wdata[20]) );
  INVX12 U5251 ( .A(\i_MIPS/n205 ), .Y(DCACHE_wdata[19]) );
  NAND2XL U5252 ( .A(n12957), .B(n5190), .Y(net105110) );
  INVX12 U5253 ( .A(n3860), .Y(DCACHE_addr[4]) );
  NAND2X1 U5254 ( .A(n9123), .B(n7145), .Y(n7146) );
  NAND2BX4 U5255 ( .AN(n3830), .B(net109519), .Y(n9218) );
  AND2XL U5256 ( .A(\i_MIPS/ALUin1[3] ), .B(n3698), .Y(n4623) );
  CLKINVX6 U5257 ( .A(n7776), .Y(n6694) );
  OAI211X2 U5258 ( .A0(net111724), .A1(net110429), .B0(n6701), .C0(n8283), .Y(
        n6820) );
  INVX2 U5259 ( .A(n8696), .Y(n8719) );
  INVXL U5260 ( .A(n9051), .Y(n8715) );
  OAI211X2 U5261 ( .A0(n8713), .A1(n8720), .B0(n8711), .C0(n8712), .Y(n8714)
         );
  BUFX8 U5262 ( .A(n5151), .Y(n5152) );
  BUFX8 U5263 ( .A(n5154), .Y(n5156) );
  BUFX4 U5264 ( .A(n5305), .Y(n5297) );
  CLKBUFX3 U5265 ( .A(n3923), .Y(n5240) );
  CLKBUFX2 U5266 ( .A(n5308), .Y(n5282) );
  BUFX8 U5267 ( .A(net117641), .Y(net117637) );
  CLKBUFX2 U5268 ( .A(n1987), .Y(n5475) );
  CLKBUFX2 U5269 ( .A(n5705), .Y(n5703) );
  CLKBUFX2 U5270 ( .A(n11210), .Y(n5928) );
  CLKBUFX2 U5271 ( .A(n4713), .Y(n5110) );
  CLKBUFX2 U5272 ( .A(n4713), .Y(n5112) );
  CLKBUFX2 U5273 ( .A(n5751), .Y(n5749) );
  CLKBUFX2 U5274 ( .A(n5841), .Y(n5839) );
  INVX3 U5275 ( .A(n144), .Y(n6824) );
  AOI21X2 U5276 ( .A0(n6914), .A1(n7399), .B0(n6913), .Y(n4736) );
  MX2X1 U5277 ( .A(n6936), .B(n8879), .S0(\i_MIPS/ID_EX[81] ), .Y(n9208) );
  OA22X1 U5278 ( .A0(n5330), .A1(n987), .B0(n5362), .B1(n2612), .Y(n7074) );
  OA22X2 U5279 ( .A0(n5807), .A1(n629), .B0(n5787), .B1(n2246), .Y(n11194) );
  OA22XL U5280 ( .A0(n5331), .A1(n1084), .B0(n5362), .B1(n2707), .Y(n7066) );
  AO22XL U5281 ( .A0(n5555), .A1(n10796), .B0(n11054), .B1(
        \i_MIPS/Sign_Extend[9] ), .Y(n10180) );
  AO22XL U5282 ( .A0(n5555), .A1(n10686), .B0(n11054), .B1(
        \i_MIPS/Sign_Extend[5] ), .Y(n10139) );
  AO22XL U5283 ( .A0(n5555), .A1(n10631), .B0(n11054), .B1(
        \i_MIPS/Sign_Extend[31] ), .Y(n10283) );
  AO22XL U5284 ( .A0(n5156), .A1(n746), .B0(n5152), .B1(n2551), .Y(n7639) );
  AO22XL U5285 ( .A0(n5156), .A1(n747), .B0(n5152), .B1(n2552), .Y(n7630) );
  AO22XL U5286 ( .A0(n5156), .A1(n748), .B0(n5152), .B1(n2553), .Y(n7729) );
  AO22XL U5287 ( .A0(n5156), .A1(n730), .B0(n5152), .B1(n2535), .Y(n7720) );
  AO22XL U5288 ( .A0(n5156), .A1(n749), .B0(n5152), .B1(n2554), .Y(n7369) );
  AO22XL U5289 ( .A0(n5156), .A1(n750), .B0(n5152), .B1(n2555), .Y(n7360) );
  AO22XL U5290 ( .A0(n5156), .A1(n751), .B0(n5152), .B1(n2556), .Y(n7289) );
  AO22XL U5291 ( .A0(n5156), .A1(n731), .B0(n5152), .B1(n2536), .Y(n7280) );
  AO22XL U5292 ( .A0(net118233), .A1(n732), .B0(net118259), .B1(n2537), .Y(
        n7384) );
  OA22XL U5293 ( .A0(\i_MIPS/Register/register[20][24] ), .A1(n5099), .B0(
        \i_MIPS/Register/register[28][24] ), .B1(n5092), .Y(n6627) );
  OA22XL U5294 ( .A0(\i_MIPS/Register/register[16][24] ), .A1(n5106), .B0(
        \i_MIPS/Register/register[24][24] ), .B1(n5105), .Y(n6626) );
  OA22XL U5295 ( .A0(\i_MIPS/Register/register[22][1] ), .A1(n5083), .B0(
        \i_MIPS/Register/register[30][1] ), .B1(n5079), .Y(n9031) );
  AND2X1 U5296 ( .A(\i_MIPS/Sign_Extend[14] ), .B(\i_MIPS/IF_ID[16] ), .Y(
        n4823) );
  AND2XL U5297 ( .A(\i_MIPS/IF_ID[15] ), .B(\i_MIPS/Sign_Extend[13] ), .Y(
        n4817) );
  NAND2XL U5298 ( .A(n3950), .B(n8567), .Y(n8574) );
  AO21X4 U5299 ( .A0(net105334), .A1(net105335), .B0(net117723), .Y(net109203)
         );
  AO22X4 U5300 ( .A0(n4711), .A1(n7602), .B0(n7601), .B1(n4682), .Y(n7603) );
  AO22X4 U5301 ( .A0(\i_MIPS/ID_EX[48] ), .A1(net143504), .B0(n5051), .B1(
        n3894), .Y(n6705) );
  CLKINVX1 U5302 ( .A(n8891), .Y(n8884) );
  OA22X2 U5303 ( .A0(n5332), .A1(n713), .B0(n5357), .B1(n2335), .Y(n9085) );
  NAND2X1 U5304 ( .A(\i_MIPS/ALUin1[4] ), .B(net111416), .Y(n9300) );
  INVX1 U5305 ( .A(n7690), .Y(n7696) );
  OA22X2 U5306 ( .A0(n5176), .A1(n714), .B0(n5215), .B1(n2336), .Y(n9087) );
  AO21X4 U5307 ( .A0(n9021), .A1(n9020), .B0(n4626), .Y(net104917) );
  BUFX8 U5308 ( .A(net117667), .Y(net117655) );
  INVX3 U5309 ( .A(n6951), .Y(n6949) );
  CLKMX2X2 U5310 ( .A(n9292), .B(n9291), .S0(net114079), .Y(n9294) );
  INVX1 U5311 ( .A(n10714), .Y(n10715) );
  INVX1 U5312 ( .A(n7867), .Y(n7865) );
  NAND2X2 U5313 ( .A(n3760), .B(n300), .Y(n7494) );
  AO21X4 U5314 ( .A0(n4762), .A1(n3673), .B0(n8298), .Y(n9133) );
  OA22X2 U5315 ( .A0(n5386), .A1(n2331), .B0(n5427), .B1(n564), .Y(n9084) );
  AO22X4 U5316 ( .A0(net118217), .A1(net104503), .B0(net118227), .B1(n7260), 
        .Y(net111364) );
  AO22X1 U5317 ( .A0(net118235), .A1(n219), .B0(net118259), .B1(n333), .Y(
        n6777) );
  AO22X1 U5318 ( .A0(net118235), .A1(n720), .B0(net118253), .B1(n2342), .Y(
        n8055) );
  OA22X1 U5319 ( .A0(\i_MIPS/Register/register[21][24] ), .A1(net118399), .B0(
        \i_MIPS/Register/register[29][24] ), .B1(net118423), .Y(n6783) );
  INVX3 U5320 ( .A(net118313), .Y(net118311) );
  INVX3 U5321 ( .A(net118337), .Y(net118335) );
  INVX1 U5322 ( .A(net110129), .Y(net110424) );
  INVX1 U5323 ( .A(n9231), .Y(n9225) );
  INVX3 U5324 ( .A(n7891), .Y(n9499) );
  INVX3 U5325 ( .A(n3977), .Y(n9443) );
  CLKMX2X2 U5326 ( .A(n8631), .B(n8630), .S0(net114079), .Y(net108893) );
  CLKMX2X2 U5327 ( .A(n8778), .B(n8777), .S0(net114079), .Y(net108640) );
  AOI211XL U5328 ( .A0(n3968), .A1(net108851), .B0(net108852), .C0(net108853), 
        .Y(n8670) );
  NAND3BX4 U5329 ( .AN(n6674), .B(n6673), .C(n6669), .Y(net112534) );
  NAND2X2 U5330 ( .A(n7423), .B(n3674), .Y(n7482) );
  OA22XL U5331 ( .A0(n5256), .A1(n1085), .B0(n5297), .B1(n2708), .Y(n7454) );
  OA22XL U5332 ( .A0(n5244), .A1(n1086), .B0(n5297), .B1(n2709), .Y(n7446) );
  INVXL U5333 ( .A(n7671), .Y(n7672) );
  INVXL U5334 ( .A(n9813), .Y(n9814) );
  AOI2BB1XL U5335 ( .A0N(n10479), .A1N(n4770), .B0(n4797), .Y(n10480) );
  NOR2BX4 U5336 ( .AN(ICACHE_addr[3]), .B(\i_MIPS/PC/n6 ), .Y(n4801) );
  OA22XL U5337 ( .A0(n5332), .A1(n2900), .B0(n5357), .B1(n1079), .Y(n9166) );
  AO22X1 U5338 ( .A0(net118271), .A1(n853), .B0(net118289), .B1(n2474), .Y(
        n7983) );
  CLKMX2X2 U5339 ( .A(\i_MIPS/ID_EX[83] ), .B(\i_MIPS/Sign_Extend[10] ), .S0(
        n3601), .Y(\i_MIPS/n438 ) );
  OA22XL U5340 ( .A0(\i_MIPS/Register/register[4][24] ), .A1(n5099), .B0(
        \i_MIPS/Register/register[12][24] ), .B1(n5092), .Y(n6618) );
  OA22XL U5341 ( .A0(\i_MIPS/Register/register[16][5] ), .A1(n5108), .B0(
        \i_MIPS/Register/register[24][5] ), .B1(n5105), .Y(n9379) );
  AO22XL U5342 ( .A0(net118239), .A1(n188), .B0(net118263), .B1(n943), .Y(
        n9331) );
  OA22XL U5343 ( .A0(\i_MIPS/Register/register[3][26] ), .A1(net118353), .B0(
        \i_MIPS/Register/register[11][26] ), .B1(net118379), .Y(n7380) );
  OA22XL U5344 ( .A0(\i_MIPS/Register/register[22][5] ), .A1(n4661), .B0(
        \i_MIPS/Register/register[30][5] ), .B1(n5079), .Y(n9373) );
  INVX3 U5345 ( .A(n8113), .Y(n8463) );
  OA22X4 U5346 ( .A0(n10620), .A1(n3767), .B0(n10622), .B1(n5189), .Y(n9272)
         );
  INVX1 U5347 ( .A(n9427), .Y(n6926) );
  INVX6 U5348 ( .A(net118365), .Y(net118355) );
  INVX6 U5349 ( .A(net118367), .Y(net118357) );
  INVX3 U5350 ( .A(net118441), .Y(net118431) );
  INVXL U5351 ( .A(n8555), .Y(n7155) );
  CLKBUFX2 U5352 ( .A(n5446), .Y(n5451) );
  NAND3BX2 U5353 ( .AN(n8884), .B(n8883), .C(n3950), .Y(n8897) );
  INVX3 U5354 ( .A(n11503), .Y(n10699) );
  INVX3 U5355 ( .A(n11470), .Y(n10595) );
  INVX3 U5356 ( .A(n11471), .Y(n10702) );
  INVX3 U5357 ( .A(n11438), .Y(n10601) );
  INVX1 U5358 ( .A(n11110), .Y(n11111) );
  INVX1 U5359 ( .A(n8855), .Y(n8858) );
  NAND2X1 U5360 ( .A(n7233), .B(n3674), .Y(n7840) );
  AND2X8 U5361 ( .A(n9544), .B(n3705), .Y(n4714) );
  INVX3 U5362 ( .A(n11502), .Y(n10592) );
  INVX1 U5363 ( .A(n7781), .Y(n7779) );
  INVX3 U5364 ( .A(n11407), .Y(n10705) );
  CLKINVX1 U5365 ( .A(n9228), .Y(n9221) );
  INVXL U5366 ( .A(n8486), .Y(n8487) );
  BUFX8 U5367 ( .A(n9499), .Y(n5116) );
  CLKBUFX3 U5368 ( .A(n10798), .Y(n5532) );
  INVX1 U5369 ( .A(n11106), .Y(n11107) );
  MX2X2 U5370 ( .A(n7584), .B(n7583), .S0(net114065), .Y(n8374) );
  INVXL U5371 ( .A(n8299), .Y(n7685) );
  CLKINVX1 U5372 ( .A(n9545), .Y(n6927) );
  AO22X1 U5373 ( .A0(net118439), .A1(n163), .B0(net118417), .B1(n178), .Y(
        n7756) );
  AO22X1 U5374 ( .A0(net118439), .A1(n242), .B0(net118409), .B1(n1994), .Y(
        n7747) );
  AO22X1 U5375 ( .A0(net118483), .A1(n363), .B0(net118457), .B1(n2001), .Y(
        n7755) );
  AO22X1 U5376 ( .A0(n4758), .A1(n362), .B0(n5112), .B1(n2000), .Y(n7897) );
  AO22X1 U5377 ( .A0(n4758), .A1(n361), .B0(n5112), .B1(n1999), .Y(n7880) );
  AO21X4 U5378 ( .A0(\i_MIPS/n520 ), .A1(\i_MIPS/n156 ), .B0(n10134), .Y(
        n10904) );
  CLKBUFX2 U5379 ( .A(n3903), .Y(net114073) );
  AND2X2 U5380 ( .A(n9730), .B(n9654), .Y(net134815) );
  AO21X1 U5381 ( .A0(\i_MIPS/n506 ), .A1(n10351), .B0(n4748), .Y(n10361) );
  AND2X1 U5382 ( .A(\i_MIPS/n506 ), .B(n10633), .Y(n4749) );
  AO22X1 U5383 ( .A0(net118439), .A1(n368), .B0(net118413), .B1(n1990), .Y(
        n9469) );
  AO22X1 U5384 ( .A0(net118439), .A1(n367), .B0(net118415), .B1(n1989), .Y(
        n9478) );
  AO22X1 U5385 ( .A0(net118441), .A1(n240), .B0(net118417), .B1(n1991), .Y(
        n9579) );
  CLKINVX1 U5386 ( .A(n9654), .Y(n9731) );
  NAND4X6 U5387 ( .A(n4663), .B(n6527), .C(n6526), .D(n6525), .Y(n11217) );
  XOR3XL U5388 ( .A(\i_MIPS/IF_ID[19] ), .B(n6016), .C(n10300), .Y(n10304) );
  INVXL U5389 ( .A(n11331), .Y(n9795) );
  INVXL U5390 ( .A(n11336), .Y(n10050) );
  NAND2XL U5391 ( .A(n4783), .B(n5559), .Y(n10587) );
  OA22X1 U5392 ( .A0(n5330), .A1(n988), .B0(n5359), .B1(n2613), .Y(n7916) );
  AO22X1 U5393 ( .A0(n5555), .A1(n10910), .B0(n11054), .B1(
        \i_MIPS/Sign_Extend[3] ), .Y(n10911) );
  OA22XL U5394 ( .A0(n5332), .A1(n1087), .B0(n5357), .B1(n2710), .Y(n9170) );
  OA22XL U5395 ( .A0(n5330), .A1(n1088), .B0(n5359), .B1(n2711), .Y(n7912) );
  OAI221XL U5396 ( .A0(\i_MIPS/Register/register[18][13] ), .A1(net117639), 
        .B0(\i_MIPS/Register/register[26][13] ), .B1(net117657), .C0(n7981), 
        .Y(n7984) );
  MXI2XL U5397 ( .A(\i_MIPS/n258 ), .B(\i_MIPS/n257 ), .S0(n3601), .Y(
        \i_MIPS/n416 ) );
  MXI2XL U5398 ( .A(\i_MIPS/n256 ), .B(\i_MIPS/n255 ), .S0(n3597), .Y(
        \i_MIPS/n415 ) );
  AO22X1 U5399 ( .A0(n5158), .A1(n772), .B0(n5153), .B1(n2364), .Y(n8531) );
  AO22X1 U5400 ( .A0(n5158), .A1(n726), .B0(n5153), .B1(n2356), .Y(n8622) );
  AO22X1 U5401 ( .A0(n5157), .A1(n773), .B0(n5153), .B1(n2365), .Y(n8613) );
  AO22X1 U5402 ( .A0(n5158), .A1(n213), .B0(n5152), .B1(n323), .Y(n6621) );
  OA22X1 U5403 ( .A0(\i_MIPS/Register/register[17][21] ), .A1(net118453), .B0(
        \i_MIPS/Register/register[25][21] ), .B1(net118477), .Y(n8911) );
  OA22X1 U5404 ( .A0(\i_MIPS/Register/register[17][9] ), .A1(net118451), .B0(
        \i_MIPS/Register/register[25][9] ), .B1(net118475), .Y(n8062) );
  OA22X1 U5405 ( .A0(\i_MIPS/Register/register[19][21] ), .A1(net118357), .B0(
        \i_MIPS/Register/register[27][21] ), .B1(net118381), .Y(n8909) );
  AO22X1 U5406 ( .A0(n5158), .A1(n378), .B0(n5153), .B1(n2366), .Y(n9374) );
  OA22X1 U5407 ( .A0(\i_MIPS/Register/register[21][9] ), .A1(net118403), .B0(
        \i_MIPS/Register/register[29][9] ), .B1(net118429), .Y(n8061) );
  OA22X1 U5408 ( .A0(\i_MIPS/Register/register[1][21] ), .A1(net118453), .B0(
        \i_MIPS/Register/register[9][21] ), .B1(net118477), .Y(n8902) );
  AO21X4 U5409 ( .A0(\i_MIPS/n513 ), .A1(\i_MIPS/n163 ), .B0(n10176), .Y(
        n10257) );
  NOR2X1 U5410 ( .A(\i_MIPS/Reg_W[4] ), .B(\i_MIPS/Reg_W[3] ), .Y(
        \i_MIPS/forward_unit/n25 ) );
  NAND2XL U5411 ( .A(\i_MIPS/IR[28] ), .B(n9600), .Y(n9813) );
  CLKINVX1 U5412 ( .A(\i_MIPS/IF_ID[18] ), .Y(n10633) );
  CLKINVX1 U5413 ( .A(\i_MIPS/IR[29] ), .Y(n9811) );
  NAND2BXL U5414 ( .AN(\i_MIPS/Sign_Extend[10] ), .B(\i_MIPS/n165 ), .Y(n10255) );
  NAND2XL U5415 ( .A(\i_MIPS/IR[26] ), .B(\i_MIPS/IR[27] ), .Y(n9823) );
  CLKINVX2 U5416 ( .A(n5177), .Y(n5165) );
  CLKINVX2 U5417 ( .A(n5375), .Y(n5373) );
  CLKINVX2 U5418 ( .A(n5355), .Y(n5348) );
  CLKINVX2 U5419 ( .A(n5333), .Y(n5322) );
  CLKINVX2 U5420 ( .A(n5210), .Y(n5206) );
  CLKINVX2 U5421 ( .A(n5179), .Y(n5166) );
  CLKINVX2 U5422 ( .A(n5378), .Y(n5370) );
  CLKINVX2 U5423 ( .A(n5360), .Y(n5346) );
  CLKINVX2 U5424 ( .A(n5325), .Y(n5319) );
  CLKINVX2 U5425 ( .A(n5381), .Y(n5367) );
  CLKINVX2 U5426 ( .A(n5352), .Y(n5343) );
  CLKINVX2 U5427 ( .A(n5327), .Y(n5316) );
  CLKINVX2 U5428 ( .A(n5284), .Y(n5271) );
  CLKINVX2 U5429 ( .A(n5215), .Y(n5201) );
  CLKINVX2 U5430 ( .A(n5384), .Y(n5364) );
  CLKINVX2 U5431 ( .A(n5353), .Y(n5340) );
  CLKINVX2 U5432 ( .A(n5328), .Y(n5313) );
  CLKINVX2 U5433 ( .A(n5216), .Y(n5198) );
  CLKINVX2 U5434 ( .A(n5172), .Y(n5159) );
  CLKINVX2 U5435 ( .A(n5383), .Y(n5365) );
  CLKINVX2 U5436 ( .A(n5353), .Y(n5341) );
  CLKINVX2 U5437 ( .A(n5328), .Y(n5314) );
  CLKINVX2 U5438 ( .A(n5216), .Y(n5199) );
  CLKINVX2 U5439 ( .A(n5172), .Y(n5160) );
  CLKINVX2 U5440 ( .A(n5377), .Y(n5371) );
  CLKINVX2 U5441 ( .A(n5355), .Y(n5347) );
  CLKINVX2 U5442 ( .A(n5325), .Y(n5320) );
  CLKINVX2 U5443 ( .A(n5171), .Y(n5161) );
  CLKINVX2 U5444 ( .A(n5333), .Y(n5321) );
  CLKINVX2 U5445 ( .A(n5382), .Y(n5366) );
  CLKINVX2 U5446 ( .A(n5352), .Y(n5342) );
  CLKINVX2 U5447 ( .A(n5327), .Y(n5315) );
  CLKINVX2 U5448 ( .A(n5215), .Y(n5200) );
  CLKINVX2 U5449 ( .A(n5380), .Y(n5368) );
  CLKINVX2 U5450 ( .A(n5358), .Y(n5344) );
  CLKINVX2 U5451 ( .A(n5326), .Y(n5317) );
  CLKINVX2 U5452 ( .A(n5212), .Y(n5202) );
  CLKINVX2 U5453 ( .A(n5170), .Y(n5162) );
  CLKINVX2 U5454 ( .A(n5379), .Y(n5369) );
  CLKINVX2 U5455 ( .A(n5326), .Y(n5318) );
  CLKINVX2 U5456 ( .A(n5212), .Y(n5203) );
  CLKINVX2 U5457 ( .A(n5170), .Y(n5163) );
  CLKINVX2 U5458 ( .A(n5351), .Y(n5350) );
  CLKINVX2 U5459 ( .A(n5324), .Y(n5323) );
  CLKINVX2 U5460 ( .A(n5209), .Y(n5208) );
  CLKINVX2 U5461 ( .A(n5169), .Y(n5168) );
  CLKINVX2 U5462 ( .A(n5420), .Y(n5414) );
  CLKINVX2 U5463 ( .A(n5420), .Y(n5412) );
  CLKINVX2 U5464 ( .A(n5425), .Y(n5409) );
  CLKINVX2 U5465 ( .A(n5424), .Y(n5410) );
  CLKINVX2 U5466 ( .A(n5423), .Y(n5411) );
  CLKINVX2 U5467 ( .A(n5421), .Y(n5413) );
  CLKINVX2 U5468 ( .A(n5422), .Y(n5415) );
  CLKINVX2 U5469 ( .A(n5896), .Y(n5892) );
  CLKINVX2 U5470 ( .A(n5673), .Y(n5670) );
  CLKINVX3 U5471 ( .A(n5896), .Y(n5891) );
  CLKINVX3 U5472 ( .A(n5673), .Y(n5669) );
  CLKINVX3 U5473 ( .A(n5896), .Y(n5885) );
  CLKINVX3 U5474 ( .A(n5905), .Y(n5893) );
  CLKINVX3 U5475 ( .A(n5690), .Y(n5671) );
  CLKINVX3 U5476 ( .A(n5896), .Y(n5886) );
  CLKINVX3 U5477 ( .A(n5896), .Y(n5887) );
  CLKINVX3 U5478 ( .A(n5897), .Y(n5889) );
  CLKINVX3 U5479 ( .A(n5687), .Y(n5666) );
  CLKINVX3 U5480 ( .A(n5894), .Y(n5890) );
  CLKINVX3 U5481 ( .A(n5681), .Y(n5668) );
  CLKINVX3 U5482 ( .A(n5673), .Y(n5665) );
  CLKINVX3 U5483 ( .A(n5689), .Y(n5667) );
  CLKINVX3 U5484 ( .A(n5895), .Y(n5888) );
  CLKINVX2 U5485 ( .A(n5432), .Y(n5419) );
  CLKINVX2 U5486 ( .A(n5421), .Y(n5416) );
  CLKINVX2 U5487 ( .A(n5420), .Y(n5417) );
  CLKINVX2 U5488 ( .A(n5242), .Y(n5229) );
  CLKBUFX2 U5489 ( .A(n5246), .Y(n5243) );
  BUFX2 U5490 ( .A(n5308), .Y(n5283) );
  CLKBUFX2 U5491 ( .A(n5308), .Y(n5284) );
  CLKBUFX2 U5492 ( .A(n3923), .Y(n5239) );
  CLKBUFX2 U5493 ( .A(n3923), .Y(n5238) );
  CLKBUFX2 U5494 ( .A(n5261), .Y(n5241) );
  CLKBUFX2 U5495 ( .A(n3984), .Y(n5242) );
  BUFX2 U5496 ( .A(n5309), .Y(n5279) );
  CLKBUFX2 U5497 ( .A(n5310), .Y(n5278) );
  CLKBUFX2 U5498 ( .A(n5309), .Y(n5280) );
  CLKBUFX2 U5499 ( .A(n5309), .Y(n5281) );
  CLKBUFX2 U5500 ( .A(n3923), .Y(n5237) );
  CLKBUFX2 U5501 ( .A(n5310), .Y(n5277) );
  CLKBUFX2 U5502 ( .A(n5129), .Y(n5130) );
  CLKBUFX2 U5503 ( .A(n10797), .Y(n5528) );
  CLKBUFX2 U5504 ( .A(n5133), .Y(n5138) );
  CLKINVX3 U5505 ( .A(n5870), .Y(n5846) );
  CLKINVX3 U5506 ( .A(n5853), .Y(n5845) );
  CLKINVX3 U5507 ( .A(n5852), .Y(n5847) );
  CLKINVX3 U5508 ( .A(n5851), .Y(n5850) );
  CLKINVX2 U5509 ( .A(n5854), .Y(n5849) );
  CLKINVX3 U5510 ( .A(n5862), .Y(n5844) );
  CLKINVX3 U5511 ( .A(n5868), .Y(n5848) );
  CLKINVX2 U5512 ( .A(n5737), .Y(n5715) );
  CLKINVX3 U5513 ( .A(n5736), .Y(n5714) );
  CLKINVX3 U5514 ( .A(n5729), .Y(n5716) );
  CLKINVX3 U5515 ( .A(n5809), .Y(n5806) );
  CLKINVX3 U5516 ( .A(n5808), .Y(n5801) );
  CLKINVX3 U5517 ( .A(n5719), .Y(n5711) );
  CLKINVX3 U5518 ( .A(n5717), .Y(n5713) );
  CLKINVX3 U5519 ( .A(n5763), .Y(n5754) );
  CLKINVX3 U5520 ( .A(n5826), .Y(n5800) );
  CLKINVX3 U5521 ( .A(n5734), .Y(n5710) );
  CLKINVX3 U5522 ( .A(n5809), .Y(n5802) );
  CLKINVX3 U5523 ( .A(n5718), .Y(n5712) );
  CLKINVX3 U5524 ( .A(n5809), .Y(n5803) );
  CLKINVX3 U5525 ( .A(n5825), .Y(n5804) );
  CLKINVX2 U5526 ( .A(n5807), .Y(n5805) );
  OA22X4 U5527 ( .A0(n10667), .A1(n3879), .B0(n10670), .B1(n4495), .Y(n9020)
         );
  OA22X4 U5528 ( .A0(n10104), .A1(n3879), .B0(n10107), .B1(n4495), .Y(n7812)
         );
  AND2X8 U5529 ( .A(n6016), .B(n3589), .Y(n4642) );
  OA22X4 U5530 ( .A0(n10790), .A1(n3878), .B0(n10793), .B1(n4495), .Y(n8528)
         );
  INVXL U5531 ( .A(n8560), .Y(n7160) );
  INVX8 U5532 ( .A(net118409), .Y(net118405) );
  INVX8 U5533 ( .A(net118413), .Y(net118403) );
  INVX8 U5534 ( .A(net118457), .Y(net118451) );
  INVX8 U5535 ( .A(net118319), .Y(net118305) );
  INVX8 U5536 ( .A(net118487), .Y(net118475) );
  CLKBUFX2 U5537 ( .A(net117665), .Y(net117663) );
  INVXL U5538 ( .A(n8133), .Y(n6666) );
  CLKINVX3 U5539 ( .A(n5462), .Y(n5460) );
  CLKBUFX2 U5540 ( .A(n5929), .Y(n5923) );
  CLKBUFX2 U5541 ( .A(n5929), .Y(n5922) );
  CLKBUFX2 U5542 ( .A(n5929), .Y(n5927) );
  CLKBUFX2 U5543 ( .A(n5707), .Y(n5697) );
  CLKBUFX2 U5544 ( .A(n5707), .Y(n5698) );
  CLKBUFX2 U5545 ( .A(n5705), .Y(n5702) );
  AOI211X1 U5546 ( .A0(net109168), .A1(n4763), .B0(n7783), .C0(n7782), .Y(
        n7794) );
  XOR2X4 U5547 ( .A(n3677), .B(n3027), .Y(net107135) );
  INVX1 U5548 ( .A(n8303), .Y(n8287) );
  MX2XL U5549 ( .A(net118597), .B(net118592), .S0(n7848), .Y(n7849) );
  INVX3 U5550 ( .A(n11476), .Y(n9804) );
  INVX3 U5551 ( .A(n11412), .Y(n10755) );
  CLKINVX3 U5552 ( .A(n7432), .Y(n7434) );
  INVXL U5553 ( .A(n8386), .Y(n8387) );
  INVX3 U5554 ( .A(n11501), .Y(n10555) );
  INVX3 U5555 ( .A(n11400), .Y(n10423) );
  INVX3 U5556 ( .A(n11482), .Y(n10771) );
  INVX3 U5557 ( .A(n11402), .Y(n10204) );
  INVX3 U5558 ( .A(n11405), .Y(n10561) );
  INVX3 U5559 ( .A(n11391), .Y(n10450) );
  INVX3 U5560 ( .A(n11499), .Y(n10391) );
  INVX3 U5561 ( .A(n11478), .Y(n9940) );
  INVX3 U5562 ( .A(n11390), .Y(n10104) );
  INVX3 U5563 ( .A(n11465), .Y(n10434) );
  INVX3 U5564 ( .A(n11462), .Y(n10310) );
  INVX3 U5565 ( .A(n11409), .Y(n10670) );
  INVX3 U5566 ( .A(n11458), .Y(n10637) );
  INVX3 U5567 ( .A(n11419), .Y(n10793) );
  INVX3 U5568 ( .A(n11455), .Y(n10447) );
  INVX3 U5569 ( .A(n11423), .Y(n10453) );
  INVX3 U5570 ( .A(n11410), .Y(n10195) );
  INVX3 U5571 ( .A(n11446), .Y(n9947) );
  INVX3 U5572 ( .A(n11442), .Y(n10189) );
  INVX3 U5573 ( .A(n11430), .Y(n10316) );
  INVX3 U5574 ( .A(n11454), .Y(n10101) );
  INVX3 U5575 ( .A(n11486), .Y(n10098) );
  INVX3 U5576 ( .A(n11498), .Y(n10198) );
  INVX3 U5577 ( .A(n11475), .Y(n9799) );
  INVX3 U5578 ( .A(n11491), .Y(n10963) );
  INVX3 U5579 ( .A(n11382), .Y(n9953) );
  INVX3 U5580 ( .A(n11404), .Y(n10548) );
  INVX3 U5581 ( .A(n11500), .Y(n10542) );
  INVX3 U5582 ( .A(n11467), .Y(n10394) );
  INVX3 U5583 ( .A(n11468), .Y(n10545) );
  INVX3 U5584 ( .A(n11464), .Y(n10420) );
  INVX3 U5585 ( .A(n11432), .Y(n10426) );
  INVXL U5586 ( .A(n8873), .Y(n8875) );
  NAND2XL U5587 ( .A(net134673), .B(n3560), .Y(n8784) );
  CLKMX2X4 U5588 ( .A(net110602), .B(n7675), .S0(net114065), .Y(n8294) );
  MX2XL U5589 ( .A(net118597), .B(net118592), .S0(n9220), .Y(n8786) );
  AOI21XL U5590 ( .A0(n8291), .A1(n7784), .B0(n4724), .Y(n4696) );
  NAND2XL U5591 ( .A(net104754), .B(net104755), .Y(n10933) );
  NAND3XL U5592 ( .A(net105449), .B(net105447), .C(net105448), .Y(n10349) );
  NAND2XL U5593 ( .A(net139778), .B(net105798), .Y(n10618) );
  NAND2XL U5594 ( .A(n2938), .B(net105396), .Y(n10429) );
  NAND2XL U5595 ( .A(net139777), .B(net105764), .Y(n10796) );
  INVX1 U5596 ( .A(net107228), .Y(net111262) );
  INVX1 U5597 ( .A(n7870), .Y(n7866) );
  INVXL U5598 ( .A(n8792), .Y(n6661) );
  INVX1 U5599 ( .A(n8893), .Y(n8888) );
  INVX1 U5600 ( .A(n7963), .Y(n7951) );
  INVX1 U5601 ( .A(net111256), .Y(net111249) );
  INVX3 U5602 ( .A(n7884), .Y(n9506) );
  INVX3 U5603 ( .A(n7888), .Y(n9502) );
  INVX3 U5604 ( .A(n7890), .Y(n9500) );
  CLKBUFX2 U5605 ( .A(n5613), .Y(n5611) );
  CLKBUFX2 U5606 ( .A(n5614), .Y(n5610) );
  CLKBUFX2 U5607 ( .A(n5751), .Y(n5744) );
  CLKBUFX2 U5608 ( .A(n5751), .Y(n5743) );
  CLKBUFX2 U5609 ( .A(n5662), .Y(n5657) );
  CLKBUFX2 U5610 ( .A(n5662), .Y(n5656) );
  CLKBUFX2 U5611 ( .A(n5884), .Y(n5880) );
  CLKBUFX2 U5612 ( .A(n5797), .Y(n5789) );
  CLKBUFX2 U5613 ( .A(n5797), .Y(n5790) );
  CLKBUFX2 U5614 ( .A(n5841), .Y(n5834) );
  CLKBUFX2 U5615 ( .A(n5750), .Y(n5748) );
  CLKBUFX2 U5616 ( .A(n5797), .Y(n5794) );
  CLKBUFX2 U5617 ( .A(n5841), .Y(n5838) );
  CLKBUFX2 U5618 ( .A(n5841), .Y(n5833) );
  CLKBUFX2 U5619 ( .A(net134682), .Y(net118395) );
  AO21X4 U5620 ( .A0(n11104), .A1(n11103), .B0(n11102), .Y(n11577) );
  NAND2X4 U5621 ( .A(n6824), .B(n2184), .Y(n7400) );
  AO21X4 U5622 ( .A0(n11113), .A1(n11112), .B0(n11111), .Y(n11573) );
  OA21XL U5623 ( .A0(n7856), .A1(n8864), .B0(n8885), .Y(n7857) );
  NAND2X4 U5624 ( .A(n6949), .B(n3861), .Y(n11097) );
  NAND2X2 U5625 ( .A(n9423), .B(n6926), .Y(n6963) );
  AO21X4 U5626 ( .A0(net104866), .A1(net104867), .B0(net117727), .Y(net111764)
         );
  AO21X4 U5627 ( .A0(net105255), .A1(net105256), .B0(net117727), .Y(net111582)
         );
  AO21X4 U5628 ( .A0(net105166), .A1(net105165), .B0(net117727), .Y(net108492)
         );
  AO21X4 U5629 ( .A0(net105119), .A1(net105120), .B0(net117723), .Y(net110800)
         );
  OAI211X2 U5630 ( .A0(n3764), .A1(net110131), .B0(net110406), .C0(net108625), 
        .Y(n8279) );
  NAND2X2 U5631 ( .A(n6693), .B(n2937), .Y(n7956) );
  NAND2XL U5632 ( .A(n8645), .B(n8666), .Y(n8033) );
  NAND2XL U5633 ( .A(n6830), .B(n4682), .Y(n6836) );
  AND2XL U5634 ( .A(n11105), .B(n9539), .Y(n9463) );
  AND2X6 U5635 ( .A(n4691), .B(n8632), .Y(net134710) );
  INVX1 U5636 ( .A(n10536), .Y(n10538) );
  NAND2XL U5637 ( .A(n9204), .B(n9222), .Y(n8640) );
  AND2XL U5638 ( .A(n8671), .B(n3857), .Y(n8641) );
  OA22XL U5639 ( .A0(n5388), .A1(n1089), .B0(n5430), .B1(n2712), .Y(n8608) );
  OA22XL U5640 ( .A0(n5248), .A1(n1090), .B0(n5288), .B1(n2713), .Y(n8610) );
  OA22XL U5641 ( .A0(n5175), .A1(n1091), .B0(n5214), .B1(n2714), .Y(n8611) );
  OA22XL U5642 ( .A0(n5176), .A1(n2862), .B0(n5215), .B1(n958), .Y(n9015) );
  OA22XL U5643 ( .A0(n5388), .A1(n1092), .B0(n5430), .B1(n2715), .Y(n8749) );
  OA22XL U5644 ( .A0(n5248), .A1(n1093), .B0(n5288), .B1(n2716), .Y(n8751) );
  OA22XL U5645 ( .A0(n5175), .A1(n1094), .B0(n5214), .B1(n2717), .Y(n8752) );
  OA22X1 U5646 ( .A0(n5174), .A1(n989), .B0(n5213), .B1(n2614), .Y(n8346) );
  OA22XL U5647 ( .A0(n5389), .A1(n1095), .B0(n5452), .B1(n2718), .Y(n8520) );
  OA22XL U5648 ( .A0(n5249), .A1(n1096), .B0(n5289), .B1(n2719), .Y(n8522) );
  OA22XL U5649 ( .A0(n5174), .A1(n1097), .B0(n5213), .B1(n2720), .Y(n8523) );
  OA22XL U5650 ( .A0(n5179), .A1(n1099), .B0(n5213), .B1(n2722), .Y(n7626) );
  NAND4X2 U5651 ( .A(n9172), .B(n9171), .C(n9170), .D(n9169), .Y(n11443) );
  OA22XL U5652 ( .A0(n5245), .A1(n1100), .B0(n5286), .B1(n2723), .Y(n9171) );
  OA22XL U5653 ( .A0(n5251), .A1(n1101), .B0(n5291), .B1(n2724), .Y(n8247) );
  OA22XL U5654 ( .A0(n5174), .A1(n1102), .B0(n5213), .B1(n2725), .Y(n8248) );
  NAND4X2 U5655 ( .A(n9011), .B(n9010), .C(n9009), .D(n9008), .Y(n11441) );
  OA22XL U5656 ( .A0(n5387), .A1(n1103), .B0(n5428), .B1(n2726), .Y(n9008) );
  OA22XL U5657 ( .A0(n5176), .A1(n1104), .B0(n5215), .B1(n2727), .Y(n9011) );
  OA22XL U5658 ( .A0(n5244), .A1(n1105), .B0(n5285), .B1(n2728), .Y(n9175) );
  OA22XL U5659 ( .A0(n5177), .A1(n1106), .B0(n5216), .B1(n2729), .Y(n9176) );
  OA22XL U5660 ( .A0(n5187), .A1(n1107), .B0(n5217), .B1(n2730), .Y(n8168) );
  OA22XL U5661 ( .A0(n3923), .A1(n1108), .B0(n5297), .B1(n2731), .Y(n7532) );
  OA22XL U5662 ( .A0(n5387), .A1(n1109), .B0(n5428), .B1(n2732), .Y(n9004) );
  OA22XL U5663 ( .A0(n5176), .A1(n1110), .B0(n5215), .B1(n2733), .Y(n9007) );
  OA22XL U5664 ( .A0(n5388), .A1(n1111), .B0(n5430), .B1(n2734), .Y(n8604) );
  OA22XL U5665 ( .A0(n5248), .A1(n1112), .B0(n5288), .B1(n2735), .Y(n8606) );
  OA22XL U5666 ( .A0(n5175), .A1(n1113), .B0(n5214), .B1(n2736), .Y(n8607) );
  OA22XL U5667 ( .A0(n5176), .A1(n1114), .B0(n5215), .B1(n2737), .Y(n8935) );
  NAND4X2 U5668 ( .A(n8744), .B(n8743), .C(n8742), .D(n8741), .Y(n11472) );
  OA22XL U5669 ( .A0(n5248), .A1(n1115), .B0(n5288), .B1(n2738), .Y(n8743) );
  OA22XL U5670 ( .A0(n5175), .A1(n1116), .B0(n5214), .B1(n2739), .Y(n8744) );
  OA22XL U5671 ( .A0(n5392), .A1(n1117), .B0(n5433), .B1(n2740), .Y(n8169) );
  OA22XL U5672 ( .A0(n5252), .A1(n1118), .B0(n5292), .B1(n2741), .Y(n8171) );
  OA22XL U5673 ( .A0(n5173), .A1(n1119), .B0(n5217), .B1(n2742), .Y(n8172) );
  OA22XL U5674 ( .A0(n5389), .A1(n1120), .B0(n5452), .B1(n2743), .Y(n8596) );
  OA22XL U5675 ( .A0(n5249), .A1(n1121), .B0(n5289), .B1(n2744), .Y(n8598) );
  OA22XL U5676 ( .A0(n5175), .A1(n1122), .B0(n5214), .B1(n2745), .Y(n8599) );
  NAND4X2 U5677 ( .A(n8252), .B(n8251), .C(n8250), .D(n8249), .Y(n11388) );
  OA22XL U5678 ( .A0(n5251), .A1(n1123), .B0(n5291), .B1(n2746), .Y(n8251) );
  OA22XL U5679 ( .A0(n5174), .A1(n1124), .B0(n5213), .B1(n2747), .Y(n8252) );
  OA22XL U5680 ( .A0(n5391), .A1(n1248), .B0(n5434), .B1(n2868), .Y(n7992) );
  OA22XL U5681 ( .A0(n5178), .A1(n1249), .B0(n5217), .B1(n2869), .Y(n7995) );
  NAND4X2 U5682 ( .A(n8828), .B(n8827), .C(n8826), .D(n8825), .Y(n11392) );
  OA22XL U5683 ( .A0(n5175), .A1(n1125), .B0(n5214), .B1(n2748), .Y(n8828) );
  OA22XL U5684 ( .A0(n5174), .A1(n1250), .B0(n5213), .B1(n2870), .Y(n8424) );
  OA22XL U5685 ( .A0(n5390), .A1(n1126), .B0(n5432), .B1(n2749), .Y(n8241) );
  OA22XL U5686 ( .A0(n5251), .A1(n1127), .B0(n5291), .B1(n2750), .Y(n8243) );
  OA22XL U5687 ( .A0(n5173), .A1(n1128), .B0(n5218), .B1(n2751), .Y(n8244) );
  OA22XL U5688 ( .A0(n5396), .A1(n1129), .B0(n5433), .B1(n2752), .Y(n8161) );
  OA22XL U5689 ( .A0(n5252), .A1(n1130), .B0(n5292), .B1(n2753), .Y(n8163) );
  OA22XL U5690 ( .A0(n5187), .A1(n1131), .B0(n5217), .B1(n2754), .Y(n8164) );
  OA22XL U5691 ( .A0(n5251), .A1(n1251), .B0(n5291), .B1(n2871), .Y(n8337) );
  OA22XL U5692 ( .A0(n5174), .A1(n1252), .B0(n5213), .B1(n2872), .Y(n8338) );
  NAND4X2 U5693 ( .A(n8820), .B(n8819), .C(n8818), .D(n8817), .Y(n11488) );
  OA22XL U5694 ( .A0(n5175), .A1(n1133), .B0(n5214), .B1(n2756), .Y(n8820) );
  OA22XL U5695 ( .A0(n5395), .A1(n1134), .B0(n5438), .B1(n2757), .Y(n7534) );
  OA22XL U5696 ( .A0(n5253), .A1(n1135), .B0(n5297), .B1(n2758), .Y(n7536) );
  OA22XL U5697 ( .A0(n5179), .A1(n1136), .B0(n5213), .B1(n2759), .Y(n7537) );
  OA22XL U5698 ( .A0(n5387), .A1(n1137), .B0(n5428), .B1(n2760), .Y(n8928) );
  OA22XL U5699 ( .A0(n5176), .A1(n1138), .B0(n5215), .B1(n2761), .Y(n8931) );
  OA22XL U5700 ( .A0(n5174), .A1(n1139), .B0(n5213), .B1(n2762), .Y(n8432) );
  OA22XL U5701 ( .A0(n5397), .A1(n1140), .B0(n5433), .B1(n2763), .Y(n8079) );
  OA22XL U5702 ( .A0(n5252), .A1(n1141), .B0(n5292), .B1(n2764), .Y(n8081) );
  OA22XL U5703 ( .A0(n5178), .A1(n1142), .B0(n5217), .B1(n2765), .Y(n8082) );
  NAND4X2 U5704 ( .A(n8923), .B(n8922), .C(n8921), .D(n8920), .Y(n11493) );
  OA22XL U5705 ( .A0(n5375), .A1(n1143), .B0(n5429), .B1(n2766), .Y(n8920) );
  OA22XL U5706 ( .A0(n5176), .A1(n1145), .B0(n5215), .B1(n2768), .Y(n8923) );
  OA22XL U5707 ( .A0(n5386), .A1(n1146), .B0(n5427), .B1(n2769), .Y(n9088) );
  OA22XL U5708 ( .A0(n5245), .A1(n2905), .B0(n5286), .B1(n1238), .Y(n9090) );
  OA22XL U5709 ( .A0(n5176), .A1(n2906), .B0(n5215), .B1(n1239), .Y(n9091) );
  OA22XL U5710 ( .A0(n3984), .A1(n1147), .B0(n5287), .B1(n2770), .Y(n6979) );
  OA22XL U5711 ( .A0(n5181), .A1(n1148), .B0(n5213), .B1(n2771), .Y(n6980) );
  OA22XL U5712 ( .A0(n5389), .A1(n1149), .B0(n5452), .B1(n2772), .Y(n8516) );
  OA22XL U5713 ( .A0(n5249), .A1(n1150), .B0(n5289), .B1(n2773), .Y(n8518) );
  OA22XL U5714 ( .A0(n5253), .A1(n1151), .B0(n5293), .B1(n2774), .Y(n7998) );
  OA22XL U5715 ( .A0(n5178), .A1(n1152), .B0(n5217), .B1(n2775), .Y(n7999) );
  OA22XL U5716 ( .A0(n5250), .A1(n954), .B0(n5290), .B1(n2578), .Y(n8341) );
  OA22XL U5717 ( .A0(n5174), .A1(n955), .B0(n5213), .B1(n2579), .Y(n8342) );
  OA22XL U5718 ( .A0(n5385), .A1(n1153), .B0(n5426), .B1(n2776), .Y(n9259) );
  OA22XL U5719 ( .A0(n5244), .A1(n1154), .B0(n5285), .B1(n2777), .Y(n9261) );
  OA22XL U5720 ( .A0(n5177), .A1(n1155), .B0(n5216), .B1(n2778), .Y(n9262) );
  OA22XL U5721 ( .A0(n5389), .A1(n1156), .B0(n5452), .B1(n2779), .Y(n8512) );
  OA22XL U5722 ( .A0(n5174), .A1(n1157), .B0(n5213), .B1(n2780), .Y(n8515) );
  OA22XL U5723 ( .A0(n5385), .A1(n1158), .B0(n5426), .B1(n2781), .Y(n9255) );
  OA22XL U5724 ( .A0(n5244), .A1(n1159), .B0(n5285), .B1(n2782), .Y(n9257) );
  OA22XL U5725 ( .A0(n5177), .A1(n1160), .B0(n5216), .B1(n2783), .Y(n9258) );
  OA22XL U5726 ( .A0(n5250), .A1(n1161), .B0(n5298), .B1(n2784), .Y(n7351) );
  OA22XL U5727 ( .A0(n5244), .A1(n1162), .B0(n5285), .B1(n2785), .Y(n9265) );
  OA22XL U5728 ( .A0(n5177), .A1(n1163), .B0(n5216), .B1(n2786), .Y(n9266) );
  NAND2X2 U5729 ( .A(n6686), .B(n183), .Y(n8692) );
  MX2XL U5730 ( .A(n9403), .B(n9402), .S0(net114079), .Y(n9466) );
  NAND2XL U5731 ( .A(net108851), .B(net109176), .Y(n8481) );
  NAND2XL U5732 ( .A(n9127), .B(n9126), .Y(n9128) );
  NAND2BX2 U5733 ( .AN(n10257), .B(n10258), .Y(n10262) );
  OA21XL U5734 ( .A0(n8690), .A1(n8688), .B0(n8859), .Y(n8689) );
  INVXL U5735 ( .A(n8029), .Y(n8034) );
  INVX3 U5736 ( .A(n6753), .Y(n10850) );
  NAND4X4 U5737 ( .A(n4654), .B(n11205), .C(n11204), .D(n11203), .Y(n11360) );
  MXI2XL U5738 ( .A(n7231), .B(n7230), .S0(net114065), .Y(n4763) );
  NAND3BXL U5739 ( .AN(n11505), .B(n11539), .C(n11504), .Y(n4996) );
  NAND2XL U5740 ( .A(n8673), .B(n8695), .Y(n7868) );
  NAND2XL U5741 ( .A(n8696), .B(n8692), .Y(n7034) );
  AO22XL U5742 ( .A0(net118395), .A1(n161), .B0(net118365), .B1(n179), .Y(
        n7757) );
  AO22XL U5743 ( .A0(net118395), .A1(n175), .B0(net118365), .B1(n247), .Y(
        n7748) );
  NAND2BX2 U5744 ( .AN(n11218), .B(n11540), .Y(n11586) );
  NAND2XL U5745 ( .A(n7669), .B(n7686), .Y(n7693) );
  NAND2XL U5746 ( .A(n9556), .B(\i_MIPS/n270 ), .Y(n9568) );
  OAI211XL U5747 ( .A0(n5051), .A1(n9446), .B0(n7588), .C0(n7587), .Y(n7590)
         );
  NAND4X8 U5748 ( .A(n4659), .B(n6361), .C(n6360), .D(n6359), .Y(n11218) );
  OA22X4 U5749 ( .A0(n5626), .A1(n2883), .B0(n5583), .B1(n1265), .Y(n4659) );
  OA22XL U5750 ( .A0(n5178), .A1(n1164), .B0(n5217), .B1(n2787), .Y(n9533) );
  INVXL U5751 ( .A(n8975), .Y(n9211) );
  INVXL U5752 ( .A(n8695), .Y(n8643) );
  INVXL U5753 ( .A(n7584), .Y(n6677) );
  INVXL U5754 ( .A(n8124), .Y(n8129) );
  OAI2BB1XL U5755 ( .A0N(n5051), .A1N(n4734), .B0(n8678), .Y(n8716) );
  OA22X4 U5756 ( .A0(n5662), .A1(n2971), .B0(n5614), .B1(n1288), .Y(n4664) );
  OA22X4 U5757 ( .A0(n5662), .A1(n534), .B0(n5613), .B1(n2931), .Y(n4665) );
  NAND4X6 U5758 ( .A(n4666), .B(n6372), .C(n6371), .D(n6370), .Y(n11371) );
  OA22X4 U5759 ( .A0(n5629), .A1(n1298), .B0(n5585), .B1(n3008), .Y(n4666) );
  AO22XL U5760 ( .A0(n5158), .A1(n239), .B0(n5153), .B1(n2007), .Y(n9394) );
  AO22XL U5761 ( .A0(n5158), .A1(n174), .B0(n5153), .B1(n375), .Y(n9385) );
  AO22XL U5762 ( .A0(net118235), .A1(n361), .B0(net118253), .B1(n1999), .Y(
        n7926) );
  AO22XL U5763 ( .A0(net118235), .A1(n362), .B0(net118253), .B1(n2000), .Y(
        n7935) );
  AO22XL U5764 ( .A0(n5157), .A1(n363), .B0(n5153), .B1(n2001), .Y(n7826) );
  AO22XL U5765 ( .A0(n5157), .A1(n360), .B0(n5153), .B1(n2006), .Y(n7817) );
  AO22XL U5766 ( .A0(net118481), .A1(n360), .B0(net118457), .B1(n2006), .Y(
        n7746) );
  CLKBUFX2 U5767 ( .A(net107195), .Y(net117727) );
  NAND4X6 U5768 ( .A(n4667), .B(n6368), .C(n6367), .D(n6366), .Y(n11369) );
  OA22X4 U5769 ( .A0(n5628), .A1(n2940), .B0(n5584), .B1(n1289), .Y(n4667) );
  NAND4X6 U5770 ( .A(n4668), .B(n6364), .C(n6363), .D(n6362), .Y(n11365) );
  OA22X4 U5771 ( .A0(n5627), .A1(n1310), .B0(n5607), .B1(n2962), .Y(n4668) );
  AND2XL U5772 ( .A(n4805), .B(n10373), .Y(n4744) );
  INVXL U5773 ( .A(n7842), .Y(n7843) );
  BUFX2 U5774 ( .A(n11214), .Y(n5938) );
  NOR3X1 U5775 ( .A(n4833), .B(n1988), .C(n223), .Y(\i_MIPS/Register/n105 ) );
  OA22XL U5776 ( .A0(n5724), .A1(n1589), .B0(n5677), .B1(n3276), .Y(n9657) );
  OA22XL U5777 ( .A0(n5900), .A1(n1590), .B0(n5858), .B1(n3277), .Y(n9655) );
  OA22XL U5778 ( .A0(n5634), .A1(n1591), .B0(n5590), .B1(n3278), .Y(n9658) );
  NAND2XL U5779 ( .A(DCACHE_addr[21]), .B(n5190), .Y(net104866) );
  NAND2XL U5780 ( .A(DCACHE_addr[0]), .B(n5190), .Y(net105751) );
  NAND2XL U5781 ( .A(n4625), .B(\i_MIPS/n266 ), .Y(net106037) );
  NAND2XL U5782 ( .A(DCACHE_addr[15]), .B(\i_MIPS/n266 ), .Y(net104985) );
  NAND2XL U5783 ( .A(DCACHE_addr[19]), .B(\i_MIPS/n266 ), .Y(net105142) );
  AO22XL U5784 ( .A0(net118395), .A1(n365), .B0(net118365), .B1(n2003), .Y(
        n9470) );
  AO22XL U5785 ( .A0(net118395), .A1(n364), .B0(net118367), .B1(n2002), .Y(
        n9479) );
  AO22XL U5786 ( .A0(net118395), .A1(n366), .B0(net118369), .B1(n2004), .Y(
        n9580) );
  NAND2XL U5787 ( .A(n11015), .B(n11014), .Y(n11513) );
  NAND2XL U5788 ( .A(n10997), .B(n10996), .Y(n11517) );
  NAND2XL U5789 ( .A(n3972), .B(n11009), .Y(n11518) );
  NAND2XL U5790 ( .A(n11029), .B(n11028), .Y(n11519) );
  NAND2XL U5791 ( .A(n11023), .B(n11024), .Y(n11515) );
  NAND2XL U5792 ( .A(n11046), .B(n11045), .Y(n11510) );
  NAND2XL U5793 ( .A(n11043), .B(n11042), .Y(n11512) );
  NAND2XL U5794 ( .A(n11040), .B(n11039), .Y(n11511) );
  NAND2XL U5795 ( .A(n3007), .B(n11007), .Y(n11516) );
  OR2XL U5796 ( .A(n10993), .B(n10994), .Y(n11509) );
  NAND2XL U5797 ( .A(n3715), .B(n11048), .Y(n11523) );
  NAND2XL U5798 ( .A(n11037), .B(n11036), .Y(n11522) );
  NAND2XL U5799 ( .A(n10988), .B(n10987), .Y(n11520) );
  NAND3BXL U5800 ( .AN(n9813), .B(n9601), .C(n9817), .Y(net110473) );
  NAND2X1 U5801 ( .A(\i_MIPS/Register/n119 ), .B(\i_MIPS/Register/n104 ), .Y(
        \i_MIPS/Register/n118 ) );
  NAND2X1 U5802 ( .A(\i_MIPS/Register/n117 ), .B(\i_MIPS/Register/n104 ), .Y(
        \i_MIPS/Register/n116 ) );
  NAND2X1 U5803 ( .A(\i_MIPS/Register/n115 ), .B(\i_MIPS/Register/n104 ), .Y(
        \i_MIPS/Register/n114 ) );
  NAND2X1 U5804 ( .A(\i_MIPS/Register/n113 ), .B(\i_MIPS/Register/n104 ), .Y(
        \i_MIPS/Register/n112 ) );
  NAND2X1 U5805 ( .A(\i_MIPS/Register/n111 ), .B(\i_MIPS/Register/n104 ), .Y(
        \i_MIPS/Register/n110 ) );
  NAND2X1 U5806 ( .A(\i_MIPS/Register/n109 ), .B(\i_MIPS/Register/n104 ), .Y(
        \i_MIPS/Register/n108 ) );
  NAND2X1 U5807 ( .A(\i_MIPS/Register/n107 ), .B(\i_MIPS/Register/n104 ), .Y(
        \i_MIPS/Register/n106 ) );
  NAND2X1 U5808 ( .A(\i_MIPS/Register/n131 ), .B(\i_MIPS/Register/n119 ), .Y(
        \i_MIPS/Register/n138 ) );
  NAND2X1 U5809 ( .A(\i_MIPS/Register/n131 ), .B(\i_MIPS/Register/n117 ), .Y(
        \i_MIPS/Register/n137 ) );
  NAND2X1 U5810 ( .A(\i_MIPS/Register/n131 ), .B(\i_MIPS/Register/n115 ), .Y(
        \i_MIPS/Register/n136 ) );
  NAND2X1 U5811 ( .A(\i_MIPS/Register/n131 ), .B(\i_MIPS/Register/n113 ), .Y(
        \i_MIPS/Register/n135 ) );
  NAND2X1 U5812 ( .A(\i_MIPS/Register/n131 ), .B(\i_MIPS/Register/n111 ), .Y(
        \i_MIPS/Register/n134 ) );
  NAND2X1 U5813 ( .A(\i_MIPS/Register/n131 ), .B(\i_MIPS/Register/n109 ), .Y(
        \i_MIPS/Register/n133 ) );
  NAND2X1 U5814 ( .A(\i_MIPS/Register/n131 ), .B(\i_MIPS/Register/n107 ), .Y(
        \i_MIPS/Register/n132 ) );
  NAND2X1 U5815 ( .A(\i_MIPS/Register/n131 ), .B(\i_MIPS/Register/n105 ), .Y(
        \i_MIPS/Register/n130 ) );
  NAND2X1 U5816 ( .A(\i_MIPS/Register/n140 ), .B(\i_MIPS/Register/n119 ), .Y(
        \i_MIPS/Register/n147 ) );
  NAND2X1 U5817 ( .A(\i_MIPS/Register/n140 ), .B(\i_MIPS/Register/n117 ), .Y(
        \i_MIPS/Register/n146 ) );
  NAND2X1 U5818 ( .A(\i_MIPS/Register/n140 ), .B(\i_MIPS/Register/n115 ), .Y(
        \i_MIPS/Register/n145 ) );
  NAND2X1 U5819 ( .A(\i_MIPS/Register/n140 ), .B(\i_MIPS/Register/n113 ), .Y(
        \i_MIPS/Register/n144 ) );
  NAND2X1 U5820 ( .A(\i_MIPS/Register/n140 ), .B(\i_MIPS/Register/n111 ), .Y(
        \i_MIPS/Register/n143 ) );
  NAND2X1 U5821 ( .A(\i_MIPS/Register/n140 ), .B(\i_MIPS/Register/n109 ), .Y(
        \i_MIPS/Register/n142 ) );
  NAND2X1 U5822 ( .A(\i_MIPS/Register/n140 ), .B(\i_MIPS/Register/n107 ), .Y(
        \i_MIPS/Register/n141 ) );
  NAND2X1 U5823 ( .A(\i_MIPS/Register/n140 ), .B(\i_MIPS/Register/n105 ), .Y(
        \i_MIPS/Register/n139 ) );
  NAND2X1 U5824 ( .A(\i_MIPS/Register/n122 ), .B(\i_MIPS/Register/n119 ), .Y(
        \i_MIPS/Register/n129 ) );
  NAND2X1 U5825 ( .A(\i_MIPS/Register/n122 ), .B(\i_MIPS/Register/n117 ), .Y(
        \i_MIPS/Register/n128 ) );
  NAND2X1 U5826 ( .A(\i_MIPS/Register/n122 ), .B(\i_MIPS/Register/n115 ), .Y(
        \i_MIPS/Register/n127 ) );
  NAND2X1 U5827 ( .A(\i_MIPS/Register/n122 ), .B(\i_MIPS/Register/n113 ), .Y(
        \i_MIPS/Register/n126 ) );
  NAND2X1 U5828 ( .A(\i_MIPS/Register/n122 ), .B(\i_MIPS/Register/n111 ), .Y(
        \i_MIPS/Register/n125 ) );
  NAND2X1 U5829 ( .A(\i_MIPS/Register/n122 ), .B(\i_MIPS/Register/n109 ), .Y(
        \i_MIPS/Register/n124 ) );
  NAND2X1 U5830 ( .A(\i_MIPS/Register/n122 ), .B(\i_MIPS/Register/n107 ), .Y(
        \i_MIPS/Register/n123 ) );
  NAND2X1 U5831 ( .A(\i_MIPS/Register/n122 ), .B(\i_MIPS/Register/n105 ), .Y(
        \i_MIPS/Register/n121 ) );
  CLKBUFX2 U5832 ( .A(net134685), .Y(net118491) );
  CLKBUFX2 U5833 ( .A(net134684), .Y(net118467) );
  AO22XL U5834 ( .A0(net118491), .A1(n176), .B0(net118457), .B1(n2005), .Y(
        n9578) );
  AO22XL U5835 ( .A0(net118487), .A1(n239), .B0(net118467), .B1(n2007), .Y(
        n9477) );
  AO22XL U5836 ( .A0(net118491), .A1(n174), .B0(net118467), .B1(n375), .Y(
        n9468) );
  AND2XL U5837 ( .A(n4804), .B(n10350), .Y(n4742) );
  AND2XL U5838 ( .A(n4809), .B(n10175), .Y(n4767) );
  AND2XL U5839 ( .A(\i_MIPS/n506 ), .B(n10513), .Y(n4748) );
  NAND2XL U5840 ( .A(\i_MIPS/n506 ), .B(n10577), .Y(n10581) );
  INVXL U5841 ( .A(n10906), .Y(n10907) );
  XNOR2XL U5842 ( .A(\i_MIPS/Sign_Extend[0] ), .B(\i_MIPS/IF_ID[2] ), .Y(
        n10828) );
  XOR3XL U5843 ( .A(\i_MIPS/IF_ID[8] ), .B(n2948), .C(n10145), .Y(n10150) );
  AOI2BB1XL U5844 ( .A0N(n10144), .A1N(n10153), .B0(n4815), .Y(n10145) );
  XOR3XL U5845 ( .A(\i_MIPS/IF_ID[10] ), .B(\i_MIPS/Sign_Extend[8] ), .C(
        n10166), .Y(n10171) );
  XOR3XL U5846 ( .A(\i_MIPS/Sign_Extend[12] ), .B(\i_MIPS/IF_ID[14] ), .C(
        n10490), .Y(n10495) );
  XOR3XL U5847 ( .A(\i_MIPS/IF_ID[13] ), .B(\i_MIPS/Sign_Extend[11] ), .C(
        n10480), .Y(n10484) );
  OA22XL U5848 ( .A0(n4694), .A1(n10736), .B0(\i_MIPS/PC/n3 ), .B1(net115799), 
        .Y(n10660) );
  XOR3XL U5849 ( .A(\i_MIPS/IF_ID[21] ), .B(n6016), .C(n4742), .Y(n10337) );
  XOR3XL U5850 ( .A(\i_MIPS/Sign_Extend[14] ), .B(\i_MIPS/IF_ID[16] ), .C(
        n10271), .Y(n10276) );
  AOI2BB1XL U5851 ( .A0N(n4816), .A1N(n4765), .B0(n4817), .Y(n10271) );
  XOR3XL U5852 ( .A(\i_MIPS/IF_ID[24] ), .B(n6016), .C(n4744), .Y(n10368) );
  INVXL U5853 ( .A(n11334), .Y(n10028) );
  INVXL U5854 ( .A(n11333), .Y(n9984) );
  INVXL U5855 ( .A(n11328), .Y(n9769) );
  INVXL U5856 ( .A(n11335), .Y(n10845) );
  INVXL U5857 ( .A(n11314), .Y(n10932) );
  INVXL U5858 ( .A(n11329), .Y(n9747) );
  INVXL U5859 ( .A(n11330), .Y(n11094) );
  INVXL U5860 ( .A(n11332), .Y(n10006) );
  XOR3XL U5861 ( .A(\i_MIPS/IF_ID[11] ), .B(\i_MIPS/Sign_Extend[9] ), .C(
        n10178), .Y(n10182) );
  AOI2BB1XL U5862 ( .A0N(n10177), .A1N(n10257), .B0(n4807), .Y(n10178) );
  XOR3XL U5863 ( .A(\i_MIPS/IF_ID[7] ), .B(\i_MIPS/Sign_Extend[5] ), .C(n10137), .Y(n10141) );
  AO22XL U5864 ( .A0(n5556), .A1(n10868), .B0(n11054), .B1(n168), .Y(n10869)
         );
  XOR3XL U5865 ( .A(\i_MIPS/IF_ID[5] ), .B(\i_MIPS/Sign_Extend[3] ), .C(n10909), .Y(n10914) );
  XOR3XL U5866 ( .A(\i_MIPS/IF_ID[17] ), .B(n6016), .C(n10281), .Y(n10285) );
  AOI2BB1XL U5867 ( .A0N(n10280), .A1N(n10289), .B0(n4823), .Y(n10281) );
  XOR3XL U5868 ( .A(\i_MIPS/IF_ID[15] ), .B(\i_MIPS/Sign_Extend[13] ), .C(
        n4765), .Y(n10268) );
  INVX3 U5869 ( .A(n6395), .Y(n10991) );
  INVX3 U5870 ( .A(n6415), .Y(n11000) );
  OAI221X2 U5871 ( .A0(n5172), .A1(n2958), .B0(n5222), .B1(n1317), .C0(n6473), 
        .Y(n6474) );
  INVX3 U5872 ( .A(n6464), .Y(n11046) );
  BUFX20 U5873 ( .A(n3859), .Y(n5055) );
  OAI221X2 U5874 ( .A0(n5186), .A1(n2959), .B0(n5211), .B1(n1318), .C0(n6426), 
        .Y(n6427) );
  OA22XL U5875 ( .A0(\i_MIPS/Register/register[6][1] ), .A1(net117685), .B0(
        \i_MIPS/Register/register[14][1] ), .B1(net117697), .Y(n8988) );
  OA22XL U5876 ( .A0(\i_MIPS/Register/register[6][19] ), .A1(net117681), .B0(
        \i_MIPS/Register/register[14][19] ), .B1(net117695), .Y(n8315) );
  OA22XL U5877 ( .A0(\i_MIPS/Register/register[6][11] ), .A1(net117685), .B0(
        \i_MIPS/Register/register[14][11] ), .B1(net117697), .Y(n8496) );
  MXI2X1 U5878 ( .A(\i_MIPS/n262 ), .B(\i_MIPS/n502 ), .S0(n3599), .Y(
        \i_MIPS/n452 ) );
  MXI2X1 U5879 ( .A(\i_MIPS/n248 ), .B(\i_MIPS/n247 ), .S0(n3590), .Y(
        \i_MIPS/n411 ) );
  OA21XL U5880 ( .A0(\i_MIPS/ALUin1[18] ), .A1(n5068), .B0(n7158), .Y(n6676)
         );
  MXI2XL U5881 ( .A(\i_MIPS/n207 ), .B(\i_MIPS/n208 ), .S0(n3593), .Y(
        \i_MIPS/n330 ) );
  MXI2XL U5882 ( .A(\i_MIPS/n181 ), .B(\i_MIPS/n182 ), .S0(n3591), .Y(
        \i_MIPS/n304 ) );
  XOR2XL U5883 ( .A(n10848), .B(n248), .Y(n6639) );
  XNOR2XL U5884 ( .A(n6753), .B(\i_MIPS/jump_addr[23] ), .Y(n4771) );
  NAND2BXL U5885 ( .AN(n11576), .B(net118581), .Y(n11588) );
  NAND2BXL U5886 ( .AN(net49779), .B(\i_MIPS/Control/n14 ), .Y(
        \i_MIPS/control_out[6] ) );
  CLKMX2X2 U5887 ( .A(\i_MIPS/ID_EX[87] ), .B(\i_MIPS/Sign_Extend[14] ), .S0(
        n3588), .Y(\i_MIPS/n434 ) );
  CLKMX2X2 U5888 ( .A(\i_MIPS/ID_EX[65] ), .B(n4987), .S0(n3593), .Y(
        \i_MIPS/n319 ) );
  CLKMX2X2 U5889 ( .A(\i_MIPS/ID_EX[63] ), .B(n10348), .S0(n3601), .Y(
        \i_MIPS/n323 ) );
  AO21X1 U5890 ( .A0(\i_MIPS/ID_EX[92] ), .A1(n3586), .B0(n4642), .Y(
        \i_MIPS/n429 ) );
  AO21X1 U5891 ( .A0(\i_MIPS/ID_EX[88] ), .A1(n3586), .B0(n4642), .Y(
        \i_MIPS/n433 ) );
  AO21X1 U5892 ( .A0(\i_MIPS/ID_EX[89] ), .A1(n3586), .B0(n4642), .Y(
        \i_MIPS/n432 ) );
  AO21X1 U5893 ( .A0(\i_MIPS/ID_EX[90] ), .A1(n3586), .B0(n4642), .Y(
        \i_MIPS/n431 ) );
  AO21X1 U5894 ( .A0(\i_MIPS/ID_EX[91] ), .A1(n3586), .B0(n4642), .Y(
        \i_MIPS/n430 ) );
  OA22XL U5895 ( .A0(n5331), .A1(n1165), .B0(n5356), .B1(n2788), .Y(n8609) );
  OA22XL U5896 ( .A0(n5332), .A1(n1166), .B0(n5357), .B1(n2789), .Y(n9009) );
  OA22XL U5897 ( .A0(n5330), .A1(n1167), .B0(n5355), .B1(n2790), .Y(n8246) );
  OA22XL U5898 ( .A0(n5330), .A1(n1168), .B0(n5355), .B1(n2791), .Y(n8517) );
  OA22XL U5899 ( .A0(n5330), .A1(n1169), .B0(n5361), .B1(n2792), .Y(n8521) );
  OA22XL U5900 ( .A0(n5333), .A1(n1170), .B0(n5360), .B1(n2793), .Y(n7624) );
  OA22XL U5901 ( .A0(n5334), .A1(n1171), .B0(n5361), .B1(n2794), .Y(n7531) );
  OA22XL U5902 ( .A0(n5333), .A1(n1172), .B0(n5362), .B1(n2795), .Y(n6978) );
  OA22XL U5903 ( .A0(n5331), .A1(n1173), .B0(n5356), .B1(n2796), .Y(n8750) );
  OA22XL U5904 ( .A0(n5330), .A1(n1174), .B0(n5361), .B1(n2797), .Y(n8250) );
  OA22XL U5905 ( .A0(n5330), .A1(n1253), .B0(n5359), .B1(n2873), .Y(n7993) );
  OA22XL U5906 ( .A0(n5333), .A1(n1175), .B0(n5360), .B1(n2798), .Y(n7535) );
  OA22XL U5907 ( .A0(n5332), .A1(n1176), .B0(n5357), .B1(n2799), .Y(n9005) );
  OA22XL U5908 ( .A0(n5334), .A1(n1177), .B0(n5361), .B1(n2800), .Y(n7441) );
  OA22XL U5909 ( .A0(n5330), .A1(n1254), .B0(n5361), .B1(n2874), .Y(n8336) );
  OA22XL U5910 ( .A0(n5330), .A1(n1178), .B0(n5355), .B1(n2801), .Y(n8430) );
  OA22XL U5911 ( .A0(n5330), .A1(n1179), .B0(n5359), .B1(n2802), .Y(n7997) );
  OA22XL U5912 ( .A0(n5332), .A1(n1180), .B0(n5357), .B1(n2803), .Y(n8929) );
  OA22XL U5913 ( .A0(n5333), .A1(n1181), .B0(n5358), .B1(n2804), .Y(n9260) );
  OA22XL U5914 ( .A0(n5330), .A1(n956), .B0(n5355), .B1(n2580), .Y(n8340) );
  OA22XL U5915 ( .A0(n5333), .A1(n1182), .B0(n5358), .B1(n2805), .Y(n9351) );
  OA22XL U5916 ( .A0(n5332), .A1(n1183), .B0(n5357), .B1(n2806), .Y(n9017) );
  OA22XL U5917 ( .A0(n5337), .A1(n1184), .B0(n5362), .B1(n2807), .Y(n7070) );
  OA22XL U5918 ( .A0(n5332), .A1(n1185), .B0(n5357), .B1(n2808), .Y(n9089) );
  OA22XL U5919 ( .A0(n5331), .A1(n1186), .B0(n5356), .B1(n2809), .Y(n8525) );
  OA22XL U5920 ( .A0(n5333), .A1(n1187), .B0(n5360), .B1(n2810), .Y(n7620) );
  OA22XL U5921 ( .A0(n5333), .A1(n1188), .B0(n5358), .B1(n2811), .Y(n9355) );
  OA22XL U5922 ( .A0(n5330), .A1(n1189), .B0(n5361), .B1(n2812), .Y(n8254) );
  OA22XL U5923 ( .A0(n5330), .A1(n1190), .B0(n5355), .B1(n2813), .Y(n8332) );
  OA22XL U5924 ( .A0(n5331), .A1(n1191), .B0(n5356), .B1(n2814), .Y(n8754) );
  OA22XL U5925 ( .A0(n5333), .A1(n1192), .B0(n5358), .B1(n2815), .Y(n9347) );
  OA22XL U5926 ( .A0(n5333), .A1(n1193), .B0(n5360), .B1(n2816), .Y(n7706) );
  OA22XL U5927 ( .A0(n5331), .A1(n1194), .B0(n5362), .B1(n2817), .Y(n7062) );
  OA22XL U5928 ( .A0(n5337), .A1(n1195), .B0(n5362), .B1(n2818), .Y(n7190) );
  OA22XL U5929 ( .A0(n5333), .A1(n1196), .B0(n5358), .B1(n2819), .Y(n9264) );
  OA22XL U5930 ( .A0(n5331), .A1(n1197), .B0(n5356), .B1(n2820), .Y(n8084) );
  OA22XL U5931 ( .A0(n5330), .A1(n1198), .B0(n5359), .B1(n2821), .Y(n8001) );
  OA22XL U5932 ( .A0(n5332), .A1(n1199), .B0(n5362), .B1(n2822), .Y(n7194) );
  OA22XL U5933 ( .A0(n5334), .A1(n1200), .B0(n5361), .B1(n2823), .Y(n7350) );
  OA22XL U5934 ( .A0(n5333), .A1(n1201), .B0(n5360), .B1(n2824), .Y(n7810) );
  OA22XL U5935 ( .A0(n5334), .A1(n1202), .B0(n5361), .B1(n2825), .Y(n7270) );
  OA22XL U5936 ( .A0(n5334), .A1(n1203), .B0(n5361), .B1(n2826), .Y(n7449) );
  OA22XL U5937 ( .A0(n5332), .A1(n1204), .B0(n5362), .B1(n2827), .Y(n7107) );
  OA22XL U5938 ( .A0(n5332), .A1(n1075), .B0(n5357), .B1(n2581), .Y(n9093) );
  OA22XL U5939 ( .A0(n5331), .A1(n1205), .B0(n5359), .B1(n2828), .Y(n8072) );
  OA22XL U5940 ( .A0(n5334), .A1(n1206), .B0(n5361), .B1(n2829), .Y(n7527) );
  OA22XL U5941 ( .A0(n5330), .A1(n1207), .B0(n5362), .B1(n2830), .Y(n7186) );
  OA22XL U5942 ( .A0(n5334), .A1(n1208), .B0(n5361), .B1(n2831), .Y(n7354) );
  OA22XL U5943 ( .A0(n5331), .A1(n1209), .B0(n5362), .B1(n2832), .Y(n7198) );
  OA22XL U5944 ( .A0(n5332), .A1(n1210), .B0(n5362), .B1(n2833), .Y(n7119) );
  OA22XL U5945 ( .A0(n5330), .A1(n1211), .B0(n5359), .B1(n2834), .Y(n7908) );
  OA22XL U5946 ( .A0(n5334), .A1(n1212), .B0(n5361), .B1(n2835), .Y(n7274) );
  OA22XL U5947 ( .A0(n5330), .A1(n1213), .B0(n5362), .B1(n2836), .Y(n7111) );
  OA22XL U5948 ( .A0(n5333), .A1(n1214), .B0(n5360), .B1(n2837), .Y(n7710) );
  OA22XL U5949 ( .A0(n5334), .A1(n1215), .B0(n5361), .B1(n2838), .Y(n7266) );
  OA22XL U5950 ( .A0(n5331), .A1(n1216), .B0(n5362), .B1(n2839), .Y(n6974) );
  OA22XL U5951 ( .A0(n5330), .A1(n1217), .B0(n5362), .B1(n2840), .Y(n7115) );
  OA22XL U5952 ( .A0(n5334), .A1(n1218), .B0(n5361), .B1(n2841), .Y(n7342) );
  OA22XL U5953 ( .A0(\i_MIPS/Register/register[22][0] ), .A1(net117681), .B0(
        \i_MIPS/Register/register[30][0] ), .B1(net117697), .Y(n8734) );
  OA22XL U5954 ( .A0(\i_MIPS/Register/register[22][1] ), .A1(net117681), .B0(
        \i_MIPS/Register/register[30][1] ), .B1(net117697), .Y(n8997) );
  OA22XL U5955 ( .A0(\i_MIPS/Register/register[22][11] ), .A1(net117685), .B0(
        \i_MIPS/Register/register[30][11] ), .B1(net117697), .Y(n8505) );
  MX2XL U5956 ( .A(\D_cache/cache[7][147] ), .B(n11004), .S0(n5416), .Y(
        \D_cache/n613 ) );
  MX2XL U5957 ( .A(\D_cache/cache[7][150] ), .B(n11022), .S0(n5417), .Y(
        \D_cache/n589 ) );
  NAND2BX1 U5958 ( .AN(n1287), .B(\i_MIPS/n162 ), .Y(n10164) );
  MX2XL U5959 ( .A(\D_cache/cache[7][46] ), .B(n4560), .S0(n5411), .Y(
        \D_cache/n1421 ) );
  MX2XL U5960 ( .A(\D_cache/cache[7][38] ), .B(n9949), .S0(n5411), .Y(
        \D_cache/n1485 ) );
  MX2XL U5961 ( .A(\D_cache/cache[7][34] ), .B(n10191), .S0(n5411), .Y(
        \D_cache/n1517 ) );
  MX2XL U5962 ( .A(\D_cache/cache[7][14] ), .B(n10100), .S0(n5411), .Y(
        \D_cache/n1677 ) );
  MX2XL U5963 ( .A(\D_cache/cache[7][6] ), .B(n9942), .S0(n5411), .Y(
        \D_cache/n1741 ) );
  MX2XL U5964 ( .A(\D_cache/cache[7][4] ), .B(n9810), .S0(n5416), .Y(
        \D_cache/n1757 ) );
  MX2XL U5965 ( .A(\D_cache/cache[7][3] ), .B(n4561), .S0(n5418), .Y(
        \D_cache/n1765 ) );
  MX2XL U5966 ( .A(\D_cache/cache[7][2] ), .B(n10188), .S0(n5411), .Y(
        \D_cache/n1773 ) );
  MX2XL U5967 ( .A(\D_cache/cache[7][110] ), .B(n4527), .S0(n5411), .Y(
        \D_cache/n909 ) );
  MX2XL U5968 ( .A(\D_cache/cache[7][102] ), .B(n4528), .S0(n5411), .Y(
        \D_cache/n973 ) );
  MX2XL U5969 ( .A(\D_cache/cache[7][78] ), .B(n4525), .S0(n5411), .Y(
        \D_cache/n1165 ) );
  MX2XL U5970 ( .A(\D_cache/cache[7][70] ), .B(n4526), .S0(n5411), .Y(
        \D_cache/n1229 ) );
  MX2XL U5971 ( .A(\D_cache/cache[7][59] ), .B(n4553), .S0(n5412), .Y(
        \D_cache/n1317 ) );
  MX2XL U5972 ( .A(\D_cache/cache[7][58] ), .B(n10203), .S0(n5412), .Y(
        \D_cache/n1325 ) );
  MX2XL U5973 ( .A(\D_cache/cache[7][57] ), .B(n4547), .S0(n5409), .Y(
        \D_cache/n1333 ) );
  MX2XL U5974 ( .A(\D_cache/cache[7][56] ), .B(n4548), .S0(n5409), .Y(
        \D_cache/n1341 ) );
  MX2XL U5975 ( .A(\D_cache/cache[7][54] ), .B(n4554), .S0(n5412), .Y(
        \D_cache/n1357 ) );
  MX2XL U5976 ( .A(\D_cache/cache[7][52] ), .B(n4549), .S0(n5409), .Y(
        \D_cache/n1373 ) );
  MX2XL U5977 ( .A(\D_cache/cache[7][48] ), .B(n4550), .S0(n5410), .Y(
        \D_cache/n1405 ) );
  MX2XL U5978 ( .A(\D_cache/cache[7][47] ), .B(n4551), .S0(n5410), .Y(
        \D_cache/n1413 ) );
  MX2XL U5979 ( .A(\D_cache/cache[7][44] ), .B(n4552), .S0(n5410), .Y(
        \D_cache/n1437 ) );
  MX2XL U5980 ( .A(\D_cache/cache[7][27] ), .B(n10393), .S0(n5412), .Y(
        \D_cache/n1573 ) );
  MX2XL U5981 ( .A(\D_cache/cache[7][26] ), .B(n10200), .S0(n5412), .Y(
        \D_cache/n1581 ) );
  MX2XL U5982 ( .A(\D_cache/cache[7][25] ), .B(n4555), .S0(n5409), .Y(
        \D_cache/n1589 ) );
  MX2XL U5983 ( .A(\D_cache/cache[7][24] ), .B(n4556), .S0(n5409), .Y(
        \D_cache/n1597 ) );
  MX2XL U5984 ( .A(\D_cache/cache[7][22] ), .B(n4559), .S0(n5412), .Y(
        \D_cache/n1613 ) );
  MX2XL U5985 ( .A(\D_cache/cache[7][20] ), .B(n4557), .S0(n5409), .Y(
        \D_cache/n1629 ) );
  MX2XL U5986 ( .A(\D_cache/cache[7][15] ), .B(n4558), .S0(n5413), .Y(
        \D_cache/n1669 ) );
  MX2XL U5987 ( .A(\D_cache/cache[7][63] ), .B(n4562), .S0(n5413), .Y(
        \D_cache/n1285 ) );
  MX2XL U5988 ( .A(\D_cache/cache[7][62] ), .B(n4563), .S0(n5414), .Y(
        \D_cache/n1293 ) );
  MX2XL U5989 ( .A(\D_cache/cache[7][61] ), .B(n4564), .S0(n5414), .Y(
        \D_cache/n1301 ) );
  MX2XL U5990 ( .A(\D_cache/cache[7][60] ), .B(n4565), .S0(n5414), .Y(
        \D_cache/n1309 ) );
  MX2XL U5991 ( .A(\D_cache/cache[7][55] ), .B(n10691), .S0(n5413), .Y(
        \D_cache/n1349 ) );
  MX2XL U5992 ( .A(\D_cache/cache[7][53] ), .B(n4566), .S0(n5410), .Y(
        \D_cache/n1365 ) );
  MX2XL U5993 ( .A(\D_cache/cache[7][50] ), .B(n4567), .S0(n5415), .Y(
        \D_cache/n1389 ) );
  MX2XL U5994 ( .A(\D_cache/cache[7][49] ), .B(n4568), .S0(n5415), .Y(
        \D_cache/n1397 ) );
  MX2XL U5995 ( .A(\D_cache/cache[7][41] ), .B(n4569), .S0(n5415), .Y(
        \D_cache/n1461 ) );
  MX2XL U5996 ( .A(\D_cache/cache[7][40] ), .B(n4570), .S0(n3561), .Y(
        \D_cache/n1469 ) );
  MX2XL U5997 ( .A(\D_cache/cache[7][39] ), .B(n10679), .S0(n5419), .Y(
        \D_cache/n1477 ) );
  MX2XL U5998 ( .A(\D_cache/cache[7][33] ), .B(n10666), .S0(n5418), .Y(
        \D_cache/n1525 ) );
  MX2XL U5999 ( .A(\D_cache/cache[7][30] ), .B(n4571), .S0(n5414), .Y(
        \D_cache/n1549 ) );
  MX2XL U6000 ( .A(\D_cache/cache[7][29] ), .B(n4572), .S0(n5414), .Y(
        \D_cache/n1557 ) );
  MX2XL U6001 ( .A(\D_cache/cache[7][28] ), .B(n4573), .S0(n5414), .Y(
        \D_cache/n1565 ) );
  MX2XL U6002 ( .A(\D_cache/cache[7][21] ), .B(n10516), .S0(n5410), .Y(
        \D_cache/n1621 ) );
  MX2XL U6003 ( .A(\D_cache/cache[7][18] ), .B(n4574), .S0(n5415), .Y(
        \D_cache/n1645 ) );
  MX2XL U6004 ( .A(\D_cache/cache[7][17] ), .B(n2995), .S0(n5415), .Y(
        \D_cache/n1653 ) );
  MX2XL U6005 ( .A(\D_cache/cache[7][16] ), .B(n146), .S0(n5410), .Y(
        \D_cache/n1661 ) );
  MX2XL U6006 ( .A(\D_cache/cache[7][12] ), .B(n4575), .S0(n5410), .Y(
        \D_cache/n1693 ) );
  MX2XL U6007 ( .A(\D_cache/cache[7][9] ), .B(n4576), .S0(n5415), .Y(
        \D_cache/n1717 ) );
  MX2XL U6008 ( .A(\D_cache/cache[7][8] ), .B(n10649), .S0(n5418), .Y(
        \D_cache/n1725 ) );
  MX2XL U6009 ( .A(\D_cache/cache[7][7] ), .B(n4577), .S0(n5418), .Y(
        \D_cache/n1733 ) );
  MX2XL U6010 ( .A(\D_cache/cache[7][1] ), .B(n10663), .S0(n3561), .Y(
        \D_cache/n1781 ) );
  MX2XL U6011 ( .A(\D_cache/cache[7][43] ), .B(n10789), .S0(n5417), .Y(
        \D_cache/n1445 ) );
  MX2XL U6012 ( .A(\D_cache/cache[7][42] ), .B(n4539), .S0(n5418), .Y(
        \D_cache/n1453 ) );
  MX2XL U6013 ( .A(\D_cache/cache[7][35] ), .B(n10761), .S0(n5418), .Y(
        \D_cache/n1509 ) );
  MX2XL U6014 ( .A(\D_cache/cache[7][32] ), .B(n4541), .S0(n5413), .Y(
        \D_cache/n1533 ) );
  MX2XL U6015 ( .A(\D_cache/cache[7][31] ), .B(n10701), .S0(n5413), .Y(
        \D_cache/n1541 ) );
  MX2XL U6016 ( .A(\D_cache/cache[7][23] ), .B(n3014), .S0(n5413), .Y(
        \D_cache/n1605 ) );
  MX2XL U6017 ( .A(\D_cache/cache[7][11] ), .B(n4542), .S0(n5418), .Y(
        \D_cache/n1701 ) );
  MX2XL U6018 ( .A(\D_cache/cache[7][10] ), .B(n4543), .S0(n5418), .Y(
        \D_cache/n1709 ) );
  MX2XL U6019 ( .A(\D_cache/cache[7][0] ), .B(n10740), .S0(n5413), .Y(
        \D_cache/n1796 ) );
  MX2XL U6020 ( .A(\D_cache/cache[7][127] ), .B(n10707), .S0(n5413), .Y(
        \D_cache/n773 ) );
  MX2XL U6021 ( .A(\D_cache/cache[7][126] ), .B(n10600), .S0(n5413), .Y(
        \D_cache/n781 ) );
  MX2XL U6022 ( .A(\D_cache/cache[7][125] ), .B(n10563), .S0(n5414), .Y(
        \D_cache/n789 ) );
  MX2XL U6023 ( .A(\D_cache/cache[7][124] ), .B(n10550), .S0(n5414), .Y(
        \D_cache/n797 ) );
  MX2XL U6024 ( .A(\D_cache/cache[7][123] ), .B(n4522), .S0(n5411), .Y(
        \D_cache/n805 ) );
  MX2XL U6025 ( .A(\D_cache/cache[7][122] ), .B(n4523), .S0(n5412), .Y(
        \D_cache/n813 ) );
  MX2XL U6026 ( .A(\D_cache/cache[7][121] ), .B(n10439), .S0(n5409), .Y(
        \D_cache/n821 ) );
  MX2XL U6027 ( .A(\D_cache/cache[7][120] ), .B(n4517), .S0(n5409), .Y(
        \D_cache/n829 ) );
  MX2XL U6028 ( .A(\D_cache/cache[7][119] ), .B(n10694), .S0(n5413), .Y(
        \D_cache/n837 ) );
  MX2XL U6029 ( .A(\D_cache/cache[7][118] ), .B(n10315), .S0(n5412), .Y(
        \D_cache/n845 ) );
  MX2XL U6030 ( .A(\D_cache/cache[7][117] ), .B(n10522), .S0(n5414), .Y(
        \D_cache/n853 ) );
  MX2XL U6031 ( .A(\D_cache/cache[7][116] ), .B(n4518), .S0(n5409), .Y(
        \D_cache/n861 ) );
  MX2XL U6032 ( .A(\D_cache/cache[7][114] ), .B(n10642), .S0(n5415), .Y(
        \D_cache/n877 ) );
  MX2XL U6033 ( .A(\D_cache/cache[7][113] ), .B(n10627), .S0(n5415), .Y(
        \D_cache/n885 ) );
  MX2XL U6034 ( .A(\D_cache/cache[7][112] ), .B(n4519), .S0(n5410), .Y(
        \D_cache/n893 ) );
  MX2XL U6035 ( .A(\D_cache/cache[7][111] ), .B(n4520), .S0(n5410), .Y(
        \D_cache/n901 ) );
  MX2XL U6036 ( .A(\D_cache/cache[7][108] ), .B(n4521), .S0(n5410), .Y(
        \D_cache/n925 ) );
  MX2XL U6037 ( .A(\D_cache/cache[7][105] ), .B(n10614), .S0(n5415), .Y(
        \D_cache/n949 ) );
  MX2XL U6038 ( .A(\D_cache/cache[7][104] ), .B(n10655), .S0(n5418), .Y(
        \D_cache/n957 ) );
  MX2XL U6039 ( .A(\D_cache/cache[7][103] ), .B(n10682), .S0(n5412), .Y(
        \D_cache/n965 ) );
  MX2XL U6040 ( .A(\D_cache/cache[7][98] ), .B(n10194), .S0(n5411), .Y(
        \D_cache/n1005 ) );
  MX2XL U6041 ( .A(\D_cache/cache[7][107] ), .B(n4497), .S0(n5409), .Y(
        \D_cache/n933 ) );
  MX2XL U6042 ( .A(\D_cache/cache[7][106] ), .B(n4498), .S0(n5418), .Y(
        \D_cache/n941 ) );
  MX2XL U6043 ( .A(\D_cache/cache[7][100] ), .B(n10754), .S0(n5418), .Y(
        \D_cache/n989 ) );
  MX2XL U6044 ( .A(\D_cache/cache[7][99] ), .B(n4499), .S0(n5418), .Y(
        \D_cache/n997 ) );
  MX2XL U6045 ( .A(\D_cache/cache[7][96] ), .B(n10746), .S0(n5413), .Y(
        \D_cache/n1021 ) );
  MX2XL U6046 ( .A(\D_cache/cache[7][95] ), .B(n10710), .S0(n5413), .Y(
        \D_cache/n1029 ) );
  MX2XL U6047 ( .A(\D_cache/cache[7][94] ), .B(n10603), .S0(n5415), .Y(
        \D_cache/n1037 ) );
  MX2XL U6048 ( .A(\D_cache/cache[7][93] ), .B(n10566), .S0(n5414), .Y(
        \D_cache/n1045 ) );
  MX2XL U6049 ( .A(\D_cache/cache[7][92] ), .B(n10553), .S0(n5414), .Y(
        \D_cache/n1053 ) );
  MX2XL U6050 ( .A(\D_cache/cache[7][91] ), .B(n4511), .S0(n5411), .Y(
        \D_cache/n1061 ) );
  MX2XL U6051 ( .A(\D_cache/cache[7][90] ), .B(n10209), .S0(n5412), .Y(
        \D_cache/n1069 ) );
  MX2XL U6052 ( .A(\D_cache/cache[7][89] ), .B(n10442), .S0(n5409), .Y(
        \D_cache/n1077 ) );
  MX2XL U6053 ( .A(\D_cache/cache[7][88] ), .B(n4512), .S0(n5409), .Y(
        \D_cache/n1085 ) );
  MX2XL U6054 ( .A(\D_cache/cache[7][87] ), .B(n10697), .S0(n5413), .Y(
        \D_cache/n1093 ) );
  MX2XL U6055 ( .A(\D_cache/cache[7][86] ), .B(n10318), .S0(n5412), .Y(
        \D_cache/n1101 ) );
  MX2XL U6056 ( .A(\D_cache/cache[7][85] ), .B(n10525), .S0(n5414), .Y(
        \D_cache/n1109 ) );
  MX2XL U6057 ( .A(\D_cache/cache[7][84] ), .B(n4513), .S0(n5409), .Y(
        \D_cache/n1117 ) );
  MX2XL U6058 ( .A(\D_cache/cache[7][82] ), .B(n10645), .S0(n5414), .Y(
        \D_cache/n1133 ) );
  MX2XL U6059 ( .A(\D_cache/cache[7][81] ), .B(n10630), .S0(n5415), .Y(
        \D_cache/n1141 ) );
  MX2XL U6060 ( .A(\D_cache/cache[7][80] ), .B(n4514), .S0(n5410), .Y(
        \D_cache/n1149 ) );
  MX2XL U6061 ( .A(\D_cache/cache[7][79] ), .B(n4515), .S0(n5410), .Y(
        \D_cache/n1157 ) );
  MX2XL U6062 ( .A(\D_cache/cache[7][76] ), .B(n4516), .S0(n5410), .Y(
        \D_cache/n1181 ) );
  MX2XL U6063 ( .A(\D_cache/cache[7][73] ), .B(n10617), .S0(n5415), .Y(
        \D_cache/n1205 ) );
  MX2XL U6064 ( .A(\D_cache/cache[7][72] ), .B(n10658), .S0(n3561), .Y(
        \D_cache/n1213 ) );
  MX2XL U6065 ( .A(\D_cache/cache[7][71] ), .B(n10685), .S0(n5412), .Y(
        \D_cache/n1221 ) );
  MX2XL U6066 ( .A(\D_cache/cache[7][66] ), .B(n10197), .S0(n5412), .Y(
        \D_cache/n1261 ) );
  MX2XL U6067 ( .A(\D_cache/cache[7][65] ), .B(n10672), .S0(n3561), .Y(
        \D_cache/n1269 ) );
  MX2XL U6068 ( .A(\D_cache/cache[7][75] ), .B(n4500), .S0(n5419), .Y(
        \D_cache/n1189 ) );
  MX2XL U6069 ( .A(\D_cache/cache[7][74] ), .B(n4501), .S0(n5418), .Y(
        \D_cache/n1197 ) );
  MX2XL U6070 ( .A(\D_cache/cache[7][68] ), .B(n10757), .S0(n5418), .Y(
        \D_cache/n1245 ) );
  MX2XL U6071 ( .A(\D_cache/cache[7][67] ), .B(n4502), .S0(n5418), .Y(
        \D_cache/n1253 ) );
  MX2XL U6072 ( .A(\D_cache/cache[7][64] ), .B(n10749), .S0(n5418), .Y(
        \D_cache/n1277 ) );
  MX2XL U6073 ( .A(\D_cache/cache[7][45] ), .B(n4538), .S0(n5419), .Y(
        \D_cache/n1429 ) );
  MX2XL U6074 ( .A(\D_cache/cache[7][37] ), .B(n10896), .S0(n5419), .Y(
        \D_cache/n1493 ) );
  MX2XL U6075 ( .A(\D_cache/cache[7][13] ), .B(n147), .S0(n5419), .Y(
        \D_cache/n1685 ) );
  MX2XL U6076 ( .A(\D_cache/cache[7][5] ), .B(n4537), .S0(n5419), .Y(
        \D_cache/n1749 ) );
  MX2XL U6077 ( .A(\D_cache/cache[7][51] ), .B(n4536), .S0(n5419), .Y(
        \D_cache/n1381 ) );
  MX2XL U6078 ( .A(\D_cache/cache[7][19] ), .B(n10965), .S0(n5419), .Y(
        \D_cache/n1637 ) );
  MX2XL U6079 ( .A(\D_cache/cache[7][109] ), .B(n10807), .S0(n5419), .Y(
        \D_cache/n917 ) );
  MX2XL U6080 ( .A(\D_cache/cache[7][101] ), .B(n10899), .S0(n5419), .Y(
        \D_cache/n981 ) );
  MX2XL U6081 ( .A(\D_cache/cache[7][83] ), .B(n10977), .S0(n5416), .Y(
        \D_cache/n1125 ) );
  MX2XL U6082 ( .A(\D_cache/cache[7][77] ), .B(n10810), .S0(n5419), .Y(
        \D_cache/n1173 ) );
  MX2XL U6083 ( .A(\D_cache/cache[7][69] ), .B(n10902), .S0(n5419), .Y(
        \D_cache/n1237 ) );
  XOR2XL U6084 ( .A(\i_MIPS/n496 ), .B(\i_MIPS/Reg_W[4] ), .Y(n6766) );
  MX2XL U6085 ( .A(\I_cache/cache[7][95] ), .B(n6577), .S0(n5848), .Y(n12078)
         );
  MX2XL U6086 ( .A(\I_cache/cache[7][81] ), .B(n6567), .S0(n5850), .Y(n12190)
         );
  MX2XL U6087 ( .A(\I_cache/cache[7][65] ), .B(n10873), .S0(n5850), .Y(n12318)
         );
  MX2XL U6088 ( .A(\I_cache/cache[7][49] ), .B(n6572), .S0(n5850), .Y(n12446)
         );
  MX2XL U6089 ( .A(\I_cache/cache[7][32] ), .B(n6557), .S0(n5844), .Y(n12582)
         );
  MX2XL U6090 ( .A(\I_cache/cache[7][94] ), .B(n9666), .S0(n5847), .Y(n12086)
         );
  MX2XL U6091 ( .A(\I_cache/cache[7][93] ), .B(n9688), .S0(n5842), .Y(n12094)
         );
  MX2XL U6092 ( .A(\I_cache/cache[7][92] ), .B(n9636), .S0(n5845), .Y(n12102)
         );
  MX2XL U6093 ( .A(\I_cache/cache[7][91] ), .B(n9614), .S0(n5847), .Y(n12110)
         );
  MX2XL U6094 ( .A(\I_cache/cache[7][90] ), .B(n6592), .S0(n5846), .Y(n12118)
         );
  MX2XL U6095 ( .A(\I_cache/cache[7][87] ), .B(n10011), .S0(n5846), .Y(n12142)
         );
  MX2XL U6096 ( .A(\I_cache/cache[7][86] ), .B(n9967), .S0(n5847), .Y(n12150)
         );
  MX2XL U6097 ( .A(\I_cache/cache[7][84] ), .B(n9778), .S0(n5843), .Y(n12166)
         );
  MX2XL U6098 ( .A(\I_cache/cache[7][74] ), .B(n9829), .S0(n5843), .Y(n12246)
         );
  MX2XL U6099 ( .A(\I_cache/cache[7][73] ), .B(n9873), .S0(n5846), .Y(n12254)
         );
  MX2XL U6100 ( .A(\I_cache/cache[7][72] ), .B(n9851), .S0(n5846), .Y(n12262)
         );
  MX2XL U6101 ( .A(\I_cache/cache[7][71] ), .B(n9895), .S0(n5846), .Y(n12270)
         );
  MX2XL U6102 ( .A(\I_cache/cache[7][70] ), .B(n9917), .S0(n5847), .Y(n12278)
         );
  MX2XL U6103 ( .A(\I_cache/cache[7][69] ), .B(n9710), .S0(n5842), .Y(n12286)
         );
  MX2XL U6104 ( .A(\I_cache/cache[7][63] ), .B(n6582), .S0(n5847), .Y(n12334)
         );
  MX2XL U6105 ( .A(\I_cache/cache[7][62] ), .B(n9671), .S0(n5848), .Y(n12342)
         );
  MX2XL U6106 ( .A(\I_cache/cache[7][61] ), .B(n3610), .S0(n5842), .Y(n12350)
         );
  MX2XL U6107 ( .A(\I_cache/cache[7][60] ), .B(n9641), .S0(n5848), .Y(n12358)
         );
  MX2XL U6108 ( .A(\I_cache/cache[7][59] ), .B(n9619), .S0(n5845), .Y(n12366)
         );
  MX2XL U6109 ( .A(\I_cache/cache[7][58] ), .B(n6597), .S0(n5845), .Y(n12374)
         );
  MX2XL U6110 ( .A(\I_cache/cache[7][54] ), .B(n9972), .S0(n5847), .Y(n12406)
         );
  MX2XL U6111 ( .A(\I_cache/cache[7][53] ), .B(n9994), .S0(n5847), .Y(n12414)
         );
  MX2XL U6112 ( .A(\I_cache/cache[7][52] ), .B(n9783), .S0(n5843), .Y(n12422)
         );
  MX2XL U6113 ( .A(\I_cache/cache[7][50] ), .B(n3615), .S0(n5843), .Y(n12438)
         );
  MX2XL U6114 ( .A(\I_cache/cache[7][48] ), .B(n3611), .S0(n5845), .Y(n12454)
         );
  MX2XL U6115 ( .A(\I_cache/cache[7][44] ), .B(n10121), .S0(n5845), .Y(n12486)
         );
  MX2XL U6116 ( .A(\I_cache/cache[7][43] ), .B(n10085), .S0(n5845), .Y(n12494)
         );
  MX2XL U6117 ( .A(\I_cache/cache[7][42] ), .B(n9834), .S0(n5843), .Y(n12502)
         );
  MX2XL U6118 ( .A(\I_cache/cache[7][41] ), .B(n9878), .S0(n5846), .Y(n12510)
         );
  MX2XL U6119 ( .A(\I_cache/cache[7][40] ), .B(n9856), .S0(n5846), .Y(n12518)
         );
  MX2XL U6120 ( .A(\I_cache/cache[7][39] ), .B(n9900), .S0(n5846), .Y(n12526)
         );
  MX2XL U6121 ( .A(\I_cache/cache[7][38] ), .B(n9922), .S0(n5847), .Y(n12534)
         );
  MX2XL U6122 ( .A(\I_cache/cache[7][37] ), .B(n3607), .S0(n5842), .Y(n12542)
         );
  MX2XL U6123 ( .A(\I_cache/cache[7][77] ), .B(n10214), .S0(n5845), .Y(n12222)
         );
  MX2XL U6124 ( .A(\I_cache/cache[7][76] ), .B(n10116), .S0(n5845), .Y(n12230)
         );
  MX2XL U6125 ( .A(\I_cache/cache[7][75] ), .B(n10080), .S0(n5844), .Y(n12238)
         );
  MX2XL U6126 ( .A(\I_cache/cache[7][56] ), .B(n10833), .S0(n5850), .Y(n12390)
         );
  MX2XL U6127 ( .A(\I_cache/cache[7][45] ), .B(n10219), .S0(n5845), .Y(n12478)
         );
  MX2XL U6128 ( .A(\I_cache/cache[7][36] ), .B(n10855), .S0(n5850), .Y(n12550)
         );
  MX2XL U6129 ( .A(\I_cache/cache[7][33] ), .B(n10878), .S0(n5850), .Y(n12574)
         );
  MX2XL U6130 ( .A(\I_cache/cache[7][68] ), .B(n6542), .S0(n5848), .Y(n12294)
         );
  MX2XL U6131 ( .A(\I_cache/cache[7][57] ), .B(n10038), .S0(n5844), .Y(n12382)
         );
  MX2XL U6132 ( .A(\I_cache/cache[7][55] ), .B(n10016), .S0(n5844), .Y(n12398)
         );
  MX2XL U6133 ( .A(\I_cache/cache[7][47] ), .B(n10062), .S0(n5844), .Y(n12462)
         );
  MX2XL U6134 ( .A(\I_cache/cache[7][89] ), .B(n10033), .S0(n5844), .Y(n12126)
         );
  MX2XL U6135 ( .A(\I_cache/cache[7][83] ), .B(n11074), .S0(n5848), .Y(n12174)
         );
  MX2XL U6136 ( .A(\I_cache/cache[7][78] ), .B(n10236), .S0(n5844), .Y(n12214)
         );
  MX2XL U6137 ( .A(\I_cache/cache[7][51] ), .B(n3614), .S0(n5848), .Y(n12430)
         );
  MX2XL U6138 ( .A(\I_cache/cache[7][46] ), .B(n10241), .S0(n5844), .Y(n12470)
         );
  MX2XL U6139 ( .A(\D_cache/cache[7][128] ), .B(n10995), .S0(n5416), .Y(
        \D_cache/n765 ) );
  MX2XL U6140 ( .A(\D_cache/cache[7][135] ), .B(n11008), .S0(n5416), .Y(
        \D_cache/n709 ) );
  MX2XL U6141 ( .A(\I_cache/cache[7][66] ), .B(n10915), .S0(n5850), .Y(n12310)
         );
  MX2XL U6142 ( .A(\I_cache/cache[7][67] ), .B(n10944), .S0(n5844), .Y(n12302)
         );
  MX2XL U6143 ( .A(\I_cache/cache[7][35] ), .B(n3618), .S0(n5847), .Y(n12558)
         );
  MX2XL U6144 ( .A(\I_cache/cache[7][34] ), .B(n3619), .S0(n5845), .Y(n12566)
         );
  NAND2XL U6145 ( .A(n12978), .B(n5190), .Y(net104889) );
  OA22XL U6146 ( .A0(\i_MIPS/Register/register[6][17] ), .A1(net117681), .B0(
        \i_MIPS/Register/register[14][17] ), .B1(net117703), .Y(n9239) );
  OA22XL U6147 ( .A0(\i_MIPS/Register/register[6][28] ), .A1(net117675), .B0(
        \i_MIPS/Register/register[14][28] ), .B1(net117697), .Y(n7567) );
  OA22XL U6148 ( .A0(\i_MIPS/Register/register[6][27] ), .A1(net117675), .B0(
        \i_MIPS/Register/register[14][27] ), .B1(net117697), .Y(n7653) );
  OA22XL U6149 ( .A0(\i_MIPS/Register/register[6][22] ), .A1(net117681), .B0(
        \i_MIPS/Register/register[14][22] ), .B1(net117695), .Y(n7925) );
  OAI221X1 U6150 ( .A0(\i_MIPS/Register/register[18][27] ), .A1(n5089), .B0(
        \i_MIPS/Register/register[26][27] ), .B1(n5085), .C0(n7728), .Y(n7736)
         );
  OAI221XL U6151 ( .A0(\i_MIPS/ALUin1[21] ), .A1(n5072), .B0(
        \i_MIPS/ALUin1[22] ), .B1(n5067), .C0(n6672), .Y(n7600) );
  XOR2XL U6152 ( .A(n10364), .B(ICACHE_addr[21]), .Y(n10359) );
  NAND2XL U6153 ( .A(n11574), .B(net118581), .Y(n11587) );
  XOR2XL U6154 ( .A(n10531), .B(ICACHE_addr[25]), .Y(n10389) );
  XOR2XL U6155 ( .A(n10376), .B(ICACHE_addr[23]), .Y(n11060) );
  OAI221XL U6156 ( .A0(\i_MIPS/ALUin1[10] ), .A1(n5071), .B0(
        \i_MIPS/ALUin1[9] ), .B1(n5068), .C0(n7311), .Y(n9137) );
  NAND2XL U6157 ( .A(n10371), .B(ICACHE_addr[21]), .Y(n10365) );
  NAND2X1 U6158 ( .A(mem_ready_I), .B(n11343), .Y(n11589) );
  NAND2XL U6159 ( .A(n10385), .B(ICACHE_addr[23]), .Y(n10377) );
  NAND2XL U6160 ( .A(\i_MIPS/ALUin1[30] ), .B(n9443), .Y(n9563) );
  MXI2XL U6161 ( .A(\i_MIPS/n209 ), .B(\i_MIPS/n210 ), .S0(n3605), .Y(
        \i_MIPS/n332 ) );
  MXI2XL U6162 ( .A(\i_MIPS/n221 ), .B(\i_MIPS/n222 ), .S0(net114325), .Y(
        \i_MIPS/n344 ) );
  MXI2XL U6163 ( .A(\i_MIPS/n217 ), .B(\i_MIPS/n218 ), .S0(n3603), .Y(
        \i_MIPS/n340 ) );
  MXI2XL U6164 ( .A(\i_MIPS/n211 ), .B(\i_MIPS/n212 ), .S0(n3601), .Y(
        \i_MIPS/n334 ) );
  MXI2XL U6165 ( .A(\i_MIPS/n201 ), .B(\i_MIPS/n202 ), .S0(n3603), .Y(
        \i_MIPS/n324 ) );
  MXI2XL U6166 ( .A(\i_MIPS/n235 ), .B(\i_MIPS/n236 ), .S0(n3593), .Y(
        \i_MIPS/n358 ) );
  MXI2XL U6167 ( .A(\i_MIPS/n233 ), .B(\i_MIPS/n234 ), .S0(n3590), .Y(
        \i_MIPS/n356 ) );
  MXI2XL U6168 ( .A(\i_MIPS/n223 ), .B(n3609), .S0(n3591), .Y(\i_MIPS/n346 )
         );
  MXI2XL U6169 ( .A(\i_MIPS/n205 ), .B(\i_MIPS/n206 ), .S0(n3595), .Y(
        \i_MIPS/n328 ) );
  MXI2XL U6170 ( .A(\i_MIPS/n213 ), .B(\i_MIPS/n214 ), .S0(n3599), .Y(
        \i_MIPS/n336 ) );
  MXI2XL U6171 ( .A(\i_MIPS/n215 ), .B(\i_MIPS/n216 ), .S0(n3595), .Y(
        \i_MIPS/n338 ) );
  XOR2XL U6172 ( .A(n7739), .B(\i_MIPS/ID_EX[113] ), .Y(n7743) );
  XOR2XL U6173 ( .A(\i_MIPS/n505 ), .B(\i_MIPS/ID_EX[111] ), .Y(n7740) );
  MXI2XL U6174 ( .A(\i_MIPS/n301 ), .B(n4695), .S0(n3599), .Y(\i_MIPS/n492 )
         );
  MXI2XL U6175 ( .A(\i_MIPS/n261 ), .B(\i_MIPS/n503 ), .S0(n3589), .Y(
        \i_MIPS/n451 ) );
  NAND2XL U6176 ( .A(\i_MIPS/IF_ID[9] ), .B(n1287), .Y(n10174) );
  OA22XL U6177 ( .A0(\i_MIPS/Register/register[4][28] ), .A1(n5099), .B0(
        \i_MIPS/Register/register[12][28] ), .B1(n5093), .Y(n7636) );
  OA22XL U6178 ( .A0(\i_MIPS/Register/register[0][28] ), .A1(n5107), .B0(
        \i_MIPS/Register/register[8][28] ), .B1(n5105), .Y(n7635) );
  OA22XL U6179 ( .A0(\i_MIPS/Register/register[4][7] ), .A1(n5099), .B0(
        \i_MIPS/Register/register[12][7] ), .B1(n5093), .Y(n7366) );
  OA22XL U6180 ( .A0(\i_MIPS/Register/register[0][7] ), .A1(n5107), .B0(
        \i_MIPS/Register/register[8][7] ), .B1(n5105), .Y(n7365) );
  OA22XL U6181 ( .A0(\i_MIPS/Register/register[4][14] ), .A1(n5099), .B0(
        \i_MIPS/Register/register[12][14] ), .B1(n5093), .Y(n7823) );
  OA22XL U6182 ( .A0(\i_MIPS/Register/register[0][14] ), .A1(n5107), .B0(
        \i_MIPS/Register/register[8][14] ), .B1(n5103), .Y(n7822) );
  OA22XL U6183 ( .A0(\i_MIPS/Register/register[5][4] ), .A1(net118405), .B0(
        \i_MIPS/Register/register[13][4] ), .B1(net118429), .Y(n9061) );
  OA22XL U6184 ( .A0(\i_MIPS/Register/register[1][4] ), .A1(net118453), .B0(
        \i_MIPS/Register/register[9][4] ), .B1(net118477), .Y(n9062) );
  OA22XL U6185 ( .A0(\i_MIPS/Register/register[7][4] ), .A1(net118303), .B0(
        \i_MIPS/Register/register[15][4] ), .B1(net118335), .Y(n9059) );
  OA22XL U6186 ( .A0(\i_MIPS/Register/register[5][17] ), .A1(net118407), .B0(
        \i_MIPS/Register/register[13][17] ), .B1(net118431), .Y(n9237) );
  OA22XL U6187 ( .A0(\i_MIPS/Register/register[1][17] ), .A1(net118455), .B0(
        \i_MIPS/Register/register[9][17] ), .B1(net118479), .Y(n9238) );
  OA22XL U6188 ( .A0(\i_MIPS/Register/register[7][17] ), .A1(net118311), .B0(
        \i_MIPS/Register/register[15][17] ), .B1(net118335), .Y(n9235) );
  OA22XL U6189 ( .A0(\i_MIPS/Register/register[5][28] ), .A1(net118401), .B0(
        \i_MIPS/Register/register[13][28] ), .B1(net118425), .Y(n7565) );
  OA22XL U6190 ( .A0(\i_MIPS/Register/register[1][28] ), .A1(net118453), .B0(
        \i_MIPS/Register/register[9][28] ), .B1(net118473), .Y(n7566) );
  OA22XL U6191 ( .A0(\i_MIPS/Register/register[5][8] ), .A1(net118403), .B0(
        \i_MIPS/Register/register[13][8] ), .B1(net118423), .Y(n8143) );
  OA22XL U6192 ( .A0(\i_MIPS/Register/register[1][8] ), .A1(net118451), .B0(
        \i_MIPS/Register/register[9][8] ), .B1(net118475), .Y(n8144) );
  OA22XL U6193 ( .A0(\i_MIPS/Register/register[5][12] ), .A1(net118403), .B0(
        \i_MIPS/Register/register[13][12] ), .B1(net118429), .Y(n8223) );
  OA22XL U6194 ( .A0(\i_MIPS/Register/register[1][12] ), .A1(net118451), .B0(
        \i_MIPS/Register/register[9][12] ), .B1(net118475), .Y(n8224) );
  OA22XL U6195 ( .A0(\i_MIPS/Register/register[5][20] ), .A1(net118403), .B0(
        \i_MIPS/Register/register[13][20] ), .B1(net118423), .Y(n8402) );
  OA22XL U6196 ( .A0(\i_MIPS/Register/register[1][20] ), .A1(net118451), .B0(
        \i_MIPS/Register/register[9][20] ), .B1(net118475), .Y(n8403) );
  OA22XL U6197 ( .A0(\i_MIPS/Register/register[7][20] ), .A1(net118307), .B0(
        \i_MIPS/Register/register[15][20] ), .B1(net118331), .Y(n8400) );
  OA22XL U6198 ( .A0(\i_MIPS/Register/register[5][21] ), .A1(net118405), .B0(
        \i_MIPS/Register/register[13][21] ), .B1(net118429), .Y(n8901) );
  OA22XL U6199 ( .A0(\i_MIPS/Register/register[7][21] ), .A1(net118305), .B0(
        \i_MIPS/Register/register[15][21] ), .B1(net118331), .Y(n8899) );
  OA22XL U6200 ( .A0(\i_MIPS/Register/register[5][26] ), .A1(net118401), .B0(
        \i_MIPS/Register/register[13][26] ), .B1(net118425), .Y(n7381) );
  OA22XL U6201 ( .A0(\i_MIPS/Register/register[1][26] ), .A1(net118453), .B0(
        \i_MIPS/Register/register[9][26] ), .B1(net118473), .Y(n7382) );
  OA22XL U6202 ( .A0(\i_MIPS/Register/register[7][26] ), .A1(net118305), .B0(
        \i_MIPS/Register/register[15][26] ), .B1(net118329), .Y(n7379) );
  OA22XL U6203 ( .A0(\i_MIPS/Register/register[1][7] ), .A1(net118453), .B0(
        \i_MIPS/Register/register[9][7] ), .B1(net118473), .Y(n7323) );
  OA22XL U6204 ( .A0(\i_MIPS/Register/register[7][7] ), .A1(net118305), .B0(
        \i_MIPS/Register/register[15][7] ), .B1(net118329), .Y(n7320) );
  OA22XL U6205 ( .A0(\i_MIPS/Register/register[21][22] ), .A1(net118401), .B0(
        \i_MIPS/Register/register[29][22] ), .B1(net118425), .Y(n7932) );
  OA22XL U6206 ( .A0(\i_MIPS/Register/register[17][22] ), .A1(net118453), .B0(
        \i_MIPS/Register/register[25][22] ), .B1(net118473), .Y(n7933) );
  OA22XL U6207 ( .A0(\i_MIPS/Register/register[23][22] ), .A1(net118305), .B0(
        \i_MIPS/Register/register[31][22] ), .B1(net118329), .Y(n7930) );
  OA22XL U6208 ( .A0(\i_MIPS/Register/register[5][22] ), .A1(net118401), .B0(
        \i_MIPS/Register/register[13][22] ), .B1(net118425), .Y(n7923) );
  OA22XL U6209 ( .A0(\i_MIPS/Register/register[1][22] ), .A1(net118453), .B0(
        \i_MIPS/Register/register[9][22] ), .B1(net118473), .Y(n7924) );
  OA22XL U6210 ( .A0(\i_MIPS/Register/register[7][22] ), .A1(net118305), .B0(
        \i_MIPS/Register/register[15][22] ), .B1(net118329), .Y(n7921) );
  OA22XL U6211 ( .A0(\i_MIPS/Register/register[20][26] ), .A1(n5101), .B0(
        \i_MIPS/Register/register[28][26] ), .B1(n5093), .Y(n7474) );
  OA22XL U6212 ( .A0(\i_MIPS/Register/register[16][26] ), .A1(n5107), .B0(
        \i_MIPS/Register/register[24][26] ), .B1(n5105), .Y(n7473) );
  OA22XL U6213 ( .A0(\i_MIPS/Register/register[20][10] ), .A1(n5099), .B0(
        \i_MIPS/Register/register[28][10] ), .B1(n5093), .Y(n7559) );
  OA22XL U6214 ( .A0(\i_MIPS/Register/register[16][10] ), .A1(n5107), .B0(
        \i_MIPS/Register/register[24][10] ), .B1(n5105), .Y(n7558) );
  OA22XL U6215 ( .A0(\i_MIPS/Register/register[20][20] ), .A1(n5100), .B0(
        \i_MIPS/Register/register[28][20] ), .B1(n5094), .Y(n8455) );
  OA22XL U6216 ( .A0(\i_MIPS/Register/register[16][17] ), .A1(n5107), .B0(
        \i_MIPS/Register/register[24][17] ), .B1(n5105), .Y(n9288) );
  OA22XL U6217 ( .A0(\i_MIPS/Register/register[20][28] ), .A1(n5100), .B0(
        \i_MIPS/Register/register[28][28] ), .B1(n5093), .Y(n7645) );
  OA22XL U6218 ( .A0(\i_MIPS/Register/register[16][28] ), .A1(n5107), .B0(
        \i_MIPS/Register/register[24][28] ), .B1(n5103), .Y(n7644) );
  OA22XL U6219 ( .A0(\i_MIPS/Register/register[20][13] ), .A1(n5100), .B0(
        \i_MIPS/Register/register[28][13] ), .B1(n5094), .Y(n8022) );
  OA22XL U6220 ( .A0(\i_MIPS/Register/register[16][13] ), .A1(n5108), .B0(
        \i_MIPS/Register/register[24][13] ), .B1(n5103), .Y(n8021) );
  OA22XL U6221 ( .A0(\i_MIPS/Register/register[20][21] ), .A1(n5101), .B0(
        \i_MIPS/Register/register[28][21] ), .B1(n5095), .Y(n8954) );
  OA22XL U6222 ( .A0(\i_MIPS/Register/register[16][21] ), .A1(n5109), .B0(
        \i_MIPS/Register/register[24][21] ), .B1(n5104), .Y(n8953) );
  OA22XL U6223 ( .A0(\i_MIPS/Register/register[20][7] ), .A1(n5099), .B0(
        \i_MIPS/Register/register[28][7] ), .B1(n5093), .Y(n7375) );
  OA22XL U6224 ( .A0(\i_MIPS/Register/register[16][7] ), .A1(n5107), .B0(
        \i_MIPS/Register/register[24][7] ), .B1(n5103), .Y(n7374) );
  OA22XL U6225 ( .A0(\i_MIPS/Register/register[20][6] ), .A1(n5099), .B0(
        \i_MIPS/Register/register[28][6] ), .B1(n5093), .Y(n7295) );
  OA22XL U6226 ( .A0(\i_MIPS/Register/register[16][6] ), .A1(n5107), .B0(
        \i_MIPS/Register/register[24][6] ), .B1(n5103), .Y(n7294) );
  OA22XL U6227 ( .A0(\i_MIPS/Register/register[20][14] ), .A1(n5101), .B0(
        \i_MIPS/Register/register[28][14] ), .B1(n5093), .Y(n7832) );
  OA22XL U6228 ( .A0(\i_MIPS/Register/register[16][14] ), .A1(n5107), .B0(
        \i_MIPS/Register/register[24][14] ), .B1(n5105), .Y(n7831) );
  OAI221X1 U6229 ( .A0(\i_MIPS/Register/register[2][27] ), .A1(n5089), .B0(
        \i_MIPS/Register/register[10][27] ), .B1(n5085), .C0(n7719), .Y(n7727)
         );
  OA22XL U6230 ( .A0(n5330), .A1(n2907), .B0(n5359), .B1(n1240), .Y(n9531) );
  AO22XL U6231 ( .A0(net118235), .A1(n733), .B0(net118253), .B1(n2538), .Y(
        n8146) );
  AO22XL U6232 ( .A0(n5158), .A1(n734), .B0(n5153), .B1(n2539), .Y(n9192) );
  AO22XL U6233 ( .A0(n5158), .A1(n735), .B0(n5153), .B1(n2540), .Y(n9183) );
  AO22XL U6234 ( .A0(net118235), .A1(n736), .B0(net118253), .B1(n2541), .Y(
        n8155) );
  AO22XL U6235 ( .A0(net118235), .A1(n737), .B0(net118253), .B1(n2542), .Y(
        n8226) );
  AO22XL U6236 ( .A0(net118235), .A1(n738), .B0(net118253), .B1(n2543), .Y(
        n8235) );
  AO22XL U6237 ( .A0(n5157), .A1(n752), .B0(n5153), .B1(n2557), .Y(n8269) );
  AO22XL U6238 ( .A0(n5157), .A1(n753), .B0(n5153), .B1(n2558), .Y(n8260) );
  AO22XL U6239 ( .A0(n5157), .A1(n754), .B0(n5153), .B1(n2559), .Y(n8189) );
  AO22XL U6240 ( .A0(n5157), .A1(n755), .B0(n5153), .B1(n2560), .Y(n8180) );
  AO22XL U6241 ( .A0(net118235), .A1(n739), .B0(net118253), .B1(n2544), .Y(
        n7973) );
  AO22XL U6242 ( .A0(net118233), .A1(n740), .B0(net118259), .B1(n2545), .Y(
        n7654) );
  AO22XL U6243 ( .A0(net118235), .A1(n756), .B0(net118253), .B1(n2561), .Y(
        n7982) );
  AO22XL U6244 ( .A0(net118233), .A1(n741), .B0(net118259), .B1(n2546), .Y(
        n7663) );
  AO22XL U6245 ( .A0(n5157), .A1(n742), .B0(n5153), .B1(n2547), .Y(n8099) );
  AO22XL U6246 ( .A0(n5157), .A1(n377), .B0(n5153), .B1(n2011), .Y(n8090) );
  AO22XL U6247 ( .A0(net118233), .A1(n757), .B0(net118259), .B1(n2562), .Y(
        n7568) );
  AO22XL U6248 ( .A0(n5158), .A1(n743), .B0(n5153), .B1(n2548), .Y(n9365) );
  AO22XL U6249 ( .A0(net118233), .A1(n758), .B0(net118259), .B1(n2563), .Y(
        n7577) );
  AO22XL U6250 ( .A0(net118233), .A1(n759), .B0(net118259), .B1(n2564), .Y(
        n7393) );
  AO22XL U6251 ( .A0(n5158), .A1(n760), .B0(n5153), .B1(n2565), .Y(n9283) );
  AO22XL U6252 ( .A0(n5158), .A1(n761), .B0(n5153), .B1(n2566), .Y(n9274) );
  AO22XL U6253 ( .A0(n5157), .A1(n744), .B0(n5153), .B1(n2549), .Y(n8007) );
  AO22XL U6254 ( .A0(n5158), .A1(n762), .B0(n5153), .B1(n2567), .Y(n9108) );
  AO22XL U6255 ( .A0(n5158), .A1(n763), .B0(n5153), .B1(n2568), .Y(n9099) );
  AO22XL U6256 ( .A0(net118233), .A1(n764), .B0(net118259), .B1(n2569), .Y(
        n7325) );
  AO22XL U6257 ( .A0(net118233), .A1(n745), .B0(net118259), .B1(n2550), .Y(
        n7245) );
  AO22XL U6258 ( .A0(net118233), .A1(n765), .B0(net118259), .B1(n2570), .Y(
        n7334) );
  AO22XL U6259 ( .A0(net118235), .A1(n189), .B0(net118259), .B1(n326), .Y(
        n6997) );
  AO22XL U6260 ( .A0(net118233), .A1(n766), .B0(net118259), .B1(n2571), .Y(
        n7254) );
  AO22XL U6261 ( .A0(net118235), .A1(n190), .B0(net118259), .B1(n327), .Y(
        n7170) );
  AO22XL U6262 ( .A0(net118235), .A1(n214), .B0(net118259), .B1(n334), .Y(
        n6877) );
  AO22XL U6263 ( .A0(net118235), .A1(n191), .B0(net118259), .B1(n328), .Y(
        n7179) );
  AO22XL U6264 ( .A0(net118235), .A1(n215), .B0(net118259), .B1(n335), .Y(
        n6786) );
  AO22XL U6265 ( .A0(net118239), .A1(n192), .B0(net118263), .B1(n944), .Y(
        n9064) );
  AO22XL U6266 ( .A0(net118239), .A1(n193), .B0(net118263), .B1(n945), .Y(
        n9150) );
  AO22XL U6267 ( .A0(net118239), .A1(n194), .B0(net118263), .B1(n946), .Y(
        n9159) );
  AO22XL U6268 ( .A0(net118239), .A1(n196), .B0(net118253), .B1(n948), .Y(
        n9340) );
  AO22XL U6269 ( .A0(net118239), .A1(n195), .B0(net118263), .B1(n947), .Y(
        n9073) );
  OA22XL U6270 ( .A0(\i_MIPS/Register/register[17][17] ), .A1(net118455), .B0(
        \i_MIPS/Register/register[25][17] ), .B1(net118479), .Y(n9247) );
  OA22XL U6271 ( .A0(n5330), .A1(n1219), .B0(n5359), .B1(n2842), .Y(n9518) );
  OA22XL U6272 ( .A0(n5332), .A1(n1256), .B0(n5359), .B1(n2876), .Y(n9522) );
  OA22XL U6273 ( .A0(n5333), .A1(n1220), .B0(n5358), .B1(n2843), .Y(n9409) );
  OA22XL U6274 ( .A0(n5333), .A1(n1221), .B0(n5358), .B1(n2844), .Y(n9405) );
  OA22XL U6275 ( .A0(n5333), .A1(n1222), .B0(n5358), .B1(n2845), .Y(n9413) );
  OA22XL U6276 ( .A0(\i_MIPS/Register/register[17][11] ), .A1(net118453), .B0(
        \i_MIPS/Register/register[25][11] ), .B1(net118477), .Y(n8504) );
  OA22XL U6277 ( .A0(\i_MIPS/Register/register[17][28] ), .A1(net118453), .B0(
        \i_MIPS/Register/register[25][28] ), .B1(net118473), .Y(n7575) );
  OA22XL U6278 ( .A0(\i_MIPS/Register/register[17][8] ), .A1(net118451), .B0(
        \i_MIPS/Register/register[25][8] ), .B1(net118475), .Y(n8153) );
  OA22XL U6279 ( .A0(\i_MIPS/Register/register[17][12] ), .A1(net118451), .B0(
        \i_MIPS/Register/register[25][12] ), .B1(net118475), .Y(n8233) );
  OA22XL U6280 ( .A0(\i_MIPS/Register/register[17][20] ), .A1(net118451), .B0(
        \i_MIPS/Register/register[25][20] ), .B1(net118475), .Y(n8412) );
  OA22XL U6281 ( .A0(\i_MIPS/Register/register[17][27] ), .A1(net118453), .B0(
        \i_MIPS/Register/register[25][27] ), .B1(net118473), .Y(n7661) );
  OA22XL U6282 ( .A0(\i_MIPS/Register/register[17][26] ), .A1(net118453), .B0(
        \i_MIPS/Register/register[25][26] ), .B1(net118473), .Y(n7391) );
  OA22XL U6283 ( .A0(\i_MIPS/Register/register[17][4] ), .A1(net118453), .B0(
        \i_MIPS/Register/register[25][4] ), .B1(net118477), .Y(n9071) );
  OA22XL U6284 ( .A0(\i_MIPS/Register/register[17][7] ), .A1(net118453), .B0(
        \i_MIPS/Register/register[25][7] ), .B1(net118473), .Y(n7332) );
  OA22XL U6285 ( .A0(\i_MIPS/Register/register[17][6] ), .A1(net118453), .B0(
        \i_MIPS/Register/register[25][6] ), .B1(net118473), .Y(n7252) );
  OA22XL U6286 ( .A0(\i_MIPS/Register/register[19][17] ), .A1(net118359), .B0(
        \i_MIPS/Register/register[27][17] ), .B1(net118379), .Y(n9245) );
  OA22XL U6287 ( .A0(\i_MIPS/Register/register[3][17] ), .A1(net118359), .B0(
        \i_MIPS/Register/register[11][17] ), .B1(net118379), .Y(n9236) );
  OA22XL U6288 ( .A0(\i_MIPS/Register/register[21][17] ), .A1(net118407), .B0(
        \i_MIPS/Register/register[29][17] ), .B1(net118431), .Y(n9246) );
  OA22XL U6289 ( .A0(\i_MIPS/Register/register[19][20] ), .A1(net118355), .B0(
        \i_MIPS/Register/register[27][20] ), .B1(net118379), .Y(n8410) );
  OA22XL U6290 ( .A0(\i_MIPS/Register/register[3][20] ), .A1(net118355), .B0(
        \i_MIPS/Register/register[11][20] ), .B1(net118379), .Y(n8401) );
  OA22XL U6291 ( .A0(\i_MIPS/Register/register[19][26] ), .A1(net118353), .B0(
        \i_MIPS/Register/register[27][26] ), .B1(net118379), .Y(n7389) );
  OA22XL U6292 ( .A0(\i_MIPS/Register/register[3][4] ), .A1(net118357), .B0(
        \i_MIPS/Register/register[11][4] ), .B1(net118381), .Y(n9060) );
  OA22XL U6293 ( .A0(\i_MIPS/Register/register[19][4] ), .A1(net118357), .B0(
        \i_MIPS/Register/register[27][4] ), .B1(net118381), .Y(n9069) );
  OA22XL U6294 ( .A0(\i_MIPS/Register/register[19][22] ), .A1(net118353), .B0(
        \i_MIPS/Register/register[27][22] ), .B1(net118375), .Y(n7931) );
  OA22XL U6295 ( .A0(\i_MIPS/Register/register[3][22] ), .A1(net118353), .B0(
        \i_MIPS/Register/register[11][22] ), .B1(net118379), .Y(n7922) );
  OA22XL U6296 ( .A0(\i_MIPS/Register/register[3][7] ), .A1(net118353), .B0(
        \i_MIPS/Register/register[11][7] ), .B1(net118381), .Y(n7321) );
  OA22XL U6297 ( .A0(\i_MIPS/Register/register[19][7] ), .A1(net118353), .B0(
        \i_MIPS/Register/register[27][7] ), .B1(net118375), .Y(n7330) );
  OA22XL U6298 ( .A0(\i_MIPS/Register/register[19][6] ), .A1(net118353), .B0(
        \i_MIPS/Register/register[27][6] ), .B1(net118379), .Y(n7250) );
  OA22XL U6299 ( .A0(\i_MIPS/Register/register[21][1] ), .A1(net118405), .B0(
        \i_MIPS/Register/register[29][1] ), .B1(net118429), .Y(n8995) );
  OA22XL U6300 ( .A0(\i_MIPS/Register/register[21][19] ), .A1(net118403), .B0(
        \i_MIPS/Register/register[29][19] ), .B1(net118429), .Y(n8322) );
  OA22XL U6301 ( .A0(\i_MIPS/Register/register[21][11] ), .A1(net118405), .B0(
        \i_MIPS/Register/register[29][11] ), .B1(net118429), .Y(n8503) );
  OA22XL U6302 ( .A0(\i_MIPS/Register/register[21][18] ), .A1(net118405), .B0(
        \i_MIPS/Register/register[29][18] ), .B1(net118429), .Y(n8586) );
  OA22XL U6303 ( .A0(\i_MIPS/Register/register[21][28] ), .A1(net118401), .B0(
        \i_MIPS/Register/register[29][28] ), .B1(net118425), .Y(n7574) );
  OA22XL U6304 ( .A0(\i_MIPS/Register/register[21][8] ), .A1(net118403), .B0(
        \i_MIPS/Register/register[29][8] ), .B1(net118429), .Y(n8152) );
  OA22XL U6305 ( .A0(\i_MIPS/Register/register[21][12] ), .A1(net118403), .B0(
        \i_MIPS/Register/register[29][12] ), .B1(net118429), .Y(n8232) );
  OA22XL U6306 ( .A0(\i_MIPS/Register/register[21][20] ), .A1(net118403), .B0(
        \i_MIPS/Register/register[29][20] ), .B1(net118429), .Y(n8411) );
  OA22XL U6307 ( .A0(\i_MIPS/Register/register[21][27] ), .A1(net118401), .B0(
        \i_MIPS/Register/register[29][27] ), .B1(net118425), .Y(n7660) );
  OA22XL U6308 ( .A0(\i_MIPS/Register/register[21][21] ), .A1(net118405), .B0(
        \i_MIPS/Register/register[29][21] ), .B1(net118429), .Y(n8910) );
  OA22XL U6309 ( .A0(\i_MIPS/Register/register[21][26] ), .A1(net118401), .B0(
        \i_MIPS/Register/register[29][26] ), .B1(net118425), .Y(n7390) );
  OA22XL U6310 ( .A0(\i_MIPS/Register/register[21][4] ), .A1(net118405), .B0(
        \i_MIPS/Register/register[29][4] ), .B1(net118429), .Y(n9070) );
  OA22XL U6311 ( .A0(\i_MIPS/Register/register[21][6] ), .A1(net118401), .B0(
        \i_MIPS/Register/register[29][6] ), .B1(net118425), .Y(n7251) );
  OA22XL U6312 ( .A0(\i_MIPS/Register/register[21][2] ), .A1(net118399), .B0(
        \i_MIPS/Register/register[29][2] ), .B1(net118423), .Y(n7176) );
  OA22XL U6313 ( .A0(\i_MIPS/Register/register[21][25] ), .A1(net118399), .B0(
        \i_MIPS/Register/register[29][25] ), .B1(net118423), .Y(n6883) );
  OA22XL U6314 ( .A0(\i_MIPS/Register/register[23][17] ), .A1(net118311), .B0(
        \i_MIPS/Register/register[31][17] ), .B1(net118335), .Y(n9244) );
  OA22XL U6315 ( .A0(\i_MIPS/Register/register[23][21] ), .A1(net118305), .B0(
        \i_MIPS/Register/register[31][21] ), .B1(net118331), .Y(n8908) );
  OA22XL U6316 ( .A0(\i_MIPS/Register/register[23][20] ), .A1(net118307), .B0(
        \i_MIPS/Register/register[31][20] ), .B1(net118331), .Y(n8409) );
  OA22XL U6317 ( .A0(\i_MIPS/Register/register[23][26] ), .A1(net118305), .B0(
        \i_MIPS/Register/register[31][26] ), .B1(net118329), .Y(n7388) );
  OA22XL U6318 ( .A0(\i_MIPS/Register/register[23][4] ), .A1(net118303), .B0(
        \i_MIPS/Register/register[31][4] ), .B1(net118329), .Y(n9068) );
  OA22XL U6319 ( .A0(\i_MIPS/Register/register[23][7] ), .A1(net118305), .B0(
        \i_MIPS/Register/register[31][7] ), .B1(net118329), .Y(n7329) );
  OA22XL U6320 ( .A0(\i_MIPS/Register/register[23][6] ), .A1(net118305), .B0(
        \i_MIPS/Register/register[31][6] ), .B1(net118329), .Y(n7249) );
  OA22XL U6321 ( .A0(\i_MIPS/Register/register[6][9] ), .A1(net117675), .B0(
        \i_MIPS/Register/register[14][9] ), .B1(net117695), .Y(n8054) );
  OA22XL U6322 ( .A0(\i_MIPS/Register/register[22][8] ), .A1(net117673), .B0(
        \i_MIPS/Register/register[30][8] ), .B1(net117695), .Y(n8154) );
  OA22XL U6323 ( .A0(\i_MIPS/Register/register[6][8] ), .A1(net117675), .B0(
        \i_MIPS/Register/register[14][8] ), .B1(net117695), .Y(n8145) );
  OA22XL U6324 ( .A0(\i_MIPS/Register/register[6][12] ), .A1(net117673), .B0(
        \i_MIPS/Register/register[14][12] ), .B1(net117695), .Y(n8225) );
  OA22XL U6325 ( .A0(\i_MIPS/Register/register[6][20] ), .A1(net117683), .B0(
        \i_MIPS/Register/register[14][20] ), .B1(net117695), .Y(n8404) );
  OA22XL U6326 ( .A0(\i_MIPS/Register/register[22][26] ), .A1(net117675), .B0(
        \i_MIPS/Register/register[30][26] ), .B1(net117697), .Y(n7392) );
  OA22XL U6327 ( .A0(\i_MIPS/Register/register[6][26] ), .A1(net117675), .B0(
        \i_MIPS/Register/register[14][26] ), .B1(net117697), .Y(n7383) );
  OA22XL U6328 ( .A0(\i_MIPS/Register/register[22][28] ), .A1(net117675), .B0(
        \i_MIPS/Register/register[30][28] ), .B1(net117697), .Y(n7576) );
  OA22XL U6329 ( .A0(\i_MIPS/Register/register[6][7] ), .A1(net117675), .B0(
        \i_MIPS/Register/register[14][7] ), .B1(net117697), .Y(n7324) );
  OA22XL U6330 ( .A0(\i_MIPS/Register/register[22][27] ), .A1(net117675), .B0(
        \i_MIPS/Register/register[30][27] ), .B1(net117697), .Y(n7662) );
  OA22XL U6331 ( .A0(\i_MIPS/Register/register[6][1] ), .A1(n5083), .B0(
        \i_MIPS/Register/register[14][1] ), .B1(n5079), .Y(n9022) );
  OA22XL U6332 ( .A0(\i_MIPS/Register/register[6][10] ), .A1(n5081), .B0(
        \i_MIPS/Register/register[14][10] ), .B1(n5077), .Y(n7543) );
  OA22XL U6333 ( .A0(\i_MIPS/Register/register[6][11] ), .A1(n5083), .B0(
        \i_MIPS/Register/register[14][11] ), .B1(n5079), .Y(n8530) );
  OA22XL U6334 ( .A0(\i_MIPS/Register/register[6][26] ), .A1(n5081), .B0(
        \i_MIPS/Register/register[14][26] ), .B1(n5077), .Y(n7458) );
  OA22XL U6335 ( .A0(\i_MIPS/Register/register[22][10] ), .A1(n5081), .B0(
        \i_MIPS/Register/register[30][10] ), .B1(n5077), .Y(n7552) );
  OA22XL U6336 ( .A0(\i_MIPS/Register/register[22][11] ), .A1(n5083), .B0(
        \i_MIPS/Register/register[30][11] ), .B1(n5079), .Y(n8539) );
  OA22XL U6337 ( .A0(\i_MIPS/Register/register[22][26] ), .A1(n5081), .B0(
        \i_MIPS/Register/register[30][26] ), .B1(n5077), .Y(n7467) );
  OA22XL U6338 ( .A0(\i_MIPS/Register/register[6][9] ), .A1(n5082), .B0(
        \i_MIPS/Register/register[14][9] ), .B1(n5078), .Y(n8089) );
  OA22XL U6339 ( .A0(\i_MIPS/Register/register[6][8] ), .A1(n5082), .B0(
        \i_MIPS/Register/register[14][8] ), .B1(n5078), .Y(n8179) );
  OA22XL U6340 ( .A0(\i_MIPS/Register/register[22][9] ), .A1(n5082), .B0(
        \i_MIPS/Register/register[30][9] ), .B1(n5078), .Y(n8098) );
  OA22XL U6341 ( .A0(\i_MIPS/Register/register[22][8] ), .A1(n5082), .B0(
        \i_MIPS/Register/register[30][8] ), .B1(n5078), .Y(n8188) );
  OA22XL U6342 ( .A0(\i_MIPS/Register/register[6][12] ), .A1(n5082), .B0(
        \i_MIPS/Register/register[14][12] ), .B1(n5078), .Y(n8259) );
  OA22XL U6343 ( .A0(\i_MIPS/Register/register[22][22] ), .A1(net117685), .B0(
        \i_MIPS/Register/register[30][22] ), .B1(net117695), .Y(n7934) );
  OA22XL U6344 ( .A0(\i_MIPS/Register/register[22][12] ), .A1(n5082), .B0(
        \i_MIPS/Register/register[30][12] ), .B1(n5078), .Y(n8268) );
  OA22XL U6345 ( .A0(\i_MIPS/Register/register[6][21] ), .A1(n5083), .B0(
        \i_MIPS/Register/register[14][21] ), .B1(n5079), .Y(n8938) );
  OA22XL U6346 ( .A0(\i_MIPS/Register/register[22][21] ), .A1(n5083), .B0(
        \i_MIPS/Register/register[30][21] ), .B1(n5079), .Y(n8947) );
  OA22XL U6347 ( .A0(\i_MIPS/Register/register[22][7] ), .A1(net117675), .B0(
        \i_MIPS/Register/register[30][7] ), .B1(net117697), .Y(n7333) );
  OA22XL U6348 ( .A0(\i_MIPS/Register/register[22][6] ), .A1(net117675), .B0(
        \i_MIPS/Register/register[30][6] ), .B1(net117697), .Y(n7253) );
  OA22XL U6349 ( .A0(\i_MIPS/Register/register[6][20] ), .A1(n5082), .B0(
        \i_MIPS/Register/register[14][20] ), .B1(n5078), .Y(n8439) );
  OA22XL U6350 ( .A0(\i_MIPS/Register/register[22][13] ), .A1(n5082), .B0(
        \i_MIPS/Register/register[30][13] ), .B1(n5078), .Y(n8015) );
  OA22XL U6351 ( .A0(\i_MIPS/Register/register[6][28] ), .A1(n5081), .B0(
        \i_MIPS/Register/register[14][28] ), .B1(n5077), .Y(n7629) );
  OA22XL U6352 ( .A0(\i_MIPS/Register/register[22][28] ), .A1(n5081), .B0(
        \i_MIPS/Register/register[30][28] ), .B1(n5077), .Y(n7638) );
  OA22XL U6353 ( .A0(\i_MIPS/Register/register[22][24] ), .A1(net117673), .B0(
        \i_MIPS/Register/register[30][24] ), .B1(net117691), .Y(n6785) );
  OA22XL U6354 ( .A0(\i_MIPS/Register/register[6][24] ), .A1(net117673), .B0(
        \i_MIPS/Register/register[14][24] ), .B1(net117691), .Y(n6775) );
  OA22XL U6355 ( .A0(\i_MIPS/Register/register[22][2] ), .A1(net117673), .B0(
        \i_MIPS/Register/register[30][2] ), .B1(net117691), .Y(n7178) );
  OA22XL U6356 ( .A0(\i_MIPS/Register/register[6][2] ), .A1(net117673), .B0(
        \i_MIPS/Register/register[14][2] ), .B1(net117691), .Y(n7169) );
  OA22XL U6357 ( .A0(\i_MIPS/Register/register[22][25] ), .A1(net117673), .B0(
        \i_MIPS/Register/register[30][25] ), .B1(net117691), .Y(n6885) );
  OA22XL U6358 ( .A0(\i_MIPS/Register/register[6][25] ), .A1(net117673), .B0(
        \i_MIPS/Register/register[14][25] ), .B1(net117691), .Y(n6876) );
  OA22XL U6359 ( .A0(\i_MIPS/Register/register[6][14] ), .A1(net117675), .B0(
        \i_MIPS/Register/register[14][14] ), .B1(net117697), .Y(n7745) );
  OA22XL U6360 ( .A0(\i_MIPS/Register/register[22][14] ), .A1(net117675), .B0(
        \i_MIPS/Register/register[30][14] ), .B1(net117697), .Y(n7754) );
  OA22XL U6361 ( .A0(\i_MIPS/Register/register[6][14] ), .A1(n5081), .B0(
        \i_MIPS/Register/register[14][14] ), .B1(n5077), .Y(n7816) );
  OA22XL U6362 ( .A0(\i_MIPS/Register/register[22][14] ), .A1(n5081), .B0(
        \i_MIPS/Register/register[30][14] ), .B1(n5077), .Y(n7825) );
  OA22XL U6363 ( .A0(\i_MIPS/Register/register[6][7] ), .A1(n5081), .B0(
        \i_MIPS/Register/register[14][7] ), .B1(n5077), .Y(n7359) );
  OA22XL U6364 ( .A0(\i_MIPS/Register/register[22][7] ), .A1(n5081), .B0(
        \i_MIPS/Register/register[30][7] ), .B1(n5077), .Y(n7368) );
  OA22XL U6365 ( .A0(\i_MIPS/Register/register[22][6] ), .A1(n5081), .B0(
        \i_MIPS/Register/register[30][6] ), .B1(n5077), .Y(n7288) );
  OA22XL U6366 ( .A0(\i_MIPS/Register/register[22][23] ), .A1(n5081), .B0(
        \i_MIPS/Register/register[30][23] ), .B1(n5076), .Y(n7013) );
  OA22XL U6367 ( .A0(\i_MIPS/Register/register[6][29] ), .A1(n5081), .B0(
        \i_MIPS/Register/register[14][29] ), .B1(n5076), .Y(n6893) );
  OA22XL U6368 ( .A0(\i_MIPS/Register/register[22][29] ), .A1(n5081), .B0(
        \i_MIPS/Register/register[30][29] ), .B1(n5076), .Y(n6902) );
  OA22XL U6369 ( .A0(\i_MIPS/Register/register[22][2] ), .A1(n5081), .B0(
        \i_MIPS/Register/register[30][2] ), .B1(n5076), .Y(n7210) );
  OA22XL U6370 ( .A0(\i_MIPS/Register/register[6][25] ), .A1(n5081), .B0(
        \i_MIPS/Register/register[14][25] ), .B1(n5076), .Y(n6793) );
  OA22XL U6371 ( .A0(\i_MIPS/Register/register[22][25] ), .A1(n5081), .B0(
        \i_MIPS/Register/register[30][25] ), .B1(n5076), .Y(n6802) );
  OA22XL U6372 ( .A0(\i_MIPS/Register/register[6][15] ), .A1(n5081), .B0(
        \i_MIPS/Register/register[14][15] ), .B1(n5076), .Y(n7124) );
  OA22XL U6373 ( .A0(\i_MIPS/Register/register[22][15] ), .A1(n5081), .B0(
        \i_MIPS/Register/register[30][15] ), .B1(n5076), .Y(n7133) );
  OA22XL U6374 ( .A0(\i_MIPS/Register/register[6][30] ), .A1(net117681), .B0(
        \i_MIPS/Register/register[14][30] ), .B1(net117703), .Y(n9467) );
  OA22XL U6375 ( .A0(\i_MIPS/Register/register[22][31] ), .A1(net117681), .B0(
        \i_MIPS/Register/register[30][31] ), .B1(net117703), .Y(n9586) );
  OA22XL U6376 ( .A0(\i_MIPS/Register/register[6][30] ), .A1(n5081), .B0(
        \i_MIPS/Register/register[14][30] ), .B1(n5079), .Y(n9384) );
  OA22XL U6377 ( .A0(\i_MIPS/Register/register[22][30] ), .A1(n5082), .B0(
        \i_MIPS/Register/register[30][30] ), .B1(n5079), .Y(n9393) );
  OA22XL U6378 ( .A0(\i_MIPS/Register/register[6][31] ), .A1(n4661), .B0(
        \i_MIPS/Register/register[14][31] ), .B1(n5079), .Y(n9489) );
  OA22XL U6379 ( .A0(\i_MIPS/Register/register[22][31] ), .A1(n4661), .B0(
        \i_MIPS/Register/register[30][31] ), .B1(n5079), .Y(n9498) );
  OA22XL U6380 ( .A0(\i_MIPS/Register/register[6][5] ), .A1(n4661), .B0(
        \i_MIPS/Register/register[14][5] ), .B1(n5079), .Y(n9364) );
  OA22XL U6381 ( .A0(\i_MIPS/Register/register[22][4] ), .A1(net117681), .B0(
        \i_MIPS/Register/register[30][4] ), .B1(net117703), .Y(n9072) );
  OA22XL U6382 ( .A0(\i_MIPS/Register/register[22][17] ), .A1(n5083), .B0(
        \i_MIPS/Register/register[30][17] ), .B1(n5079), .Y(n9282) );
  OA22XL U6383 ( .A0(\i_MIPS/Register/register[22][30] ), .A1(net117681), .B0(
        \i_MIPS/Register/register[30][30] ), .B1(net117703), .Y(n9476) );
  OA22XL U6384 ( .A0(\i_MIPS/Register/register[6][31] ), .A1(net117681), .B0(
        \i_MIPS/Register/register[14][31] ), .B1(net117703), .Y(n9577) );
  MX2XL U6385 ( .A(\I_cache/cache[7][150] ), .B(n11064), .S0(n5843), .Y(n11638) );
  MX2XL U6386 ( .A(\I_cache/cache[1][152] ), .B(n11068), .S0(n5580), .Y(n11628) );
  MX2XL U6387 ( .A(\I_cache/cache[6][152] ), .B(n11068), .S0(n5891), .Y(n11623) );
  MX2XL U6388 ( .A(\I_cache/cache[3][152] ), .B(n11068), .S0(n5669), .Y(n11626) );
  MX2XL U6389 ( .A(n5478), .B(\i_MIPS/Register/register[0][25] ), .S0(n6014), 
        .Y(\i_MIPS/Register/n1133 ) );
  MX2XL U6390 ( .A(n5479), .B(\i_MIPS/Register/register[7][25] ), .S0(n6000), 
        .Y(\i_MIPS/Register/n909 ) );
  MX2XL U6391 ( .A(n5476), .B(\i_MIPS/Register/register[0][24] ), .S0(n6014), 
        .Y(\i_MIPS/Register/n1132 ) );
  MX2XL U6392 ( .A(n5477), .B(\i_MIPS/Register/register[7][24] ), .S0(n6000), 
        .Y(\i_MIPS/Register/n908 ) );
  MX2XL U6393 ( .A(\I_cache/cache[7][144] ), .B(n11145), .S0(n5847), .Y(n11686) );
  MX2XL U6394 ( .A(\I_cache/cache[7][145] ), .B(n11065), .S0(n5850), .Y(n11678) );
  MX2XL U6395 ( .A(\D_cache/cache[7][153] ), .B(n10770), .S0(n5418), .Y(
        \D_cache/n565 ) );
  MX2XL U6396 ( .A(\I_cache/cache[7][134] ), .B(n11122), .S0(n5848), .Y(n11766) );
  MX2XL U6397 ( .A(\I_cache/cache[7][130] ), .B(n11155), .S0(n5849), .Y(n11798) );
  MX2XL U6398 ( .A(\I_cache/cache[7][140] ), .B(n11150), .S0(n5849), .Y(n11718) );
  MX2XL U6399 ( .A(\I_cache/cache[7][139] ), .B(n11140), .S0(n5848), .Y(n11726) );
  MX2XL U6400 ( .A(\I_cache/cache[7][137] ), .B(n11172), .S0(n5849), .Y(n11742) );
  MX2XL U6401 ( .A(\I_cache/cache[7][135] ), .B(n11177), .S0(n5849), .Y(n11758) );
  MX2XL U6402 ( .A(\I_cache/cache[7][131] ), .B(n11159), .S0(n5849), .Y(n11790) );
  MX2XL U6403 ( .A(\I_cache/cache[7][129] ), .B(n11164), .S0(n5849), .Y(n11806) );
  MX2XL U6404 ( .A(\I_cache/cache[7][128] ), .B(n11067), .S0(n5848), .Y(n11814) );
  MX2XL U6405 ( .A(\I_cache/cache[7][138] ), .B(n11131), .S0(n5848), .Y(n11734) );
  MX2XL U6406 ( .A(\I_cache/cache[7][152] ), .B(n11068), .S0(n5848), .Y(n11622) );
  MX2XL U6407 ( .A(\I_cache/cache[7][151] ), .B(n11066), .S0(n5848), .Y(n11630) );
  MX2XL U6408 ( .A(\I_cache/cache[7][136] ), .B(n11182), .S0(n5849), .Y(n11750) );
  MX2XL U6409 ( .A(\I_cache/cache[7][132] ), .B(n11118), .S0(n5848), .Y(n11782) );
  MX2XL U6410 ( .A(\I_cache/cache[7][149] ), .B(n11187), .S0(n5849), .Y(n11646) );
  MX2XL U6411 ( .A(\I_cache/cache[7][147] ), .B(n11192), .S0(n5849), .Y(n11662) );
  MX2XL U6412 ( .A(\I_cache/cache[7][142] ), .B(n11201), .S0(n5849), .Y(n11702) );
  MX2XL U6413 ( .A(\I_cache/cache[6][130] ), .B(n11155), .S0(n5892), .Y(n11799) );
  MX2XL U6414 ( .A(\I_cache/cache[3][130] ), .B(n11155), .S0(n5670), .Y(n11802) );
  MX2XL U6415 ( .A(\I_cache/cache[2][130] ), .B(n11155), .S0(n5715), .Y(n11803) );
  MX2XL U6416 ( .A(\I_cache/cache[1][130] ), .B(n11155), .S0(n5581), .Y(n11804) );
  MX2XL U6417 ( .A(\I_cache/cache[0][130] ), .B(n11155), .S0(n5624), .Y(n11805) );
  MX2XL U6418 ( .A(\I_cache/cache[6][140] ), .B(n11150), .S0(n5892), .Y(n11719) );
  MX2XL U6419 ( .A(\I_cache/cache[3][140] ), .B(n11150), .S0(n5670), .Y(n11722) );
  MX2XL U6420 ( .A(\I_cache/cache[2][140] ), .B(n11150), .S0(n5715), .Y(n11723) );
  MX2XL U6421 ( .A(\I_cache/cache[1][140] ), .B(n11150), .S0(n5581), .Y(n11724) );
  MX2XL U6422 ( .A(\I_cache/cache[0][140] ), .B(n11150), .S0(n5624), .Y(n11725) );
  MX2XL U6423 ( .A(\I_cache/cache[6][137] ), .B(n11172), .S0(n5892), .Y(n11743) );
  MX2XL U6424 ( .A(\I_cache/cache[3][137] ), .B(n11172), .S0(n5670), .Y(n11746) );
  MX2XL U6425 ( .A(\I_cache/cache[2][137] ), .B(n11172), .S0(n5715), .Y(n11747) );
  MX2XL U6426 ( .A(\I_cache/cache[1][137] ), .B(n11172), .S0(n5581), .Y(n11748) );
  MX2XL U6427 ( .A(\I_cache/cache[0][137] ), .B(n11172), .S0(n5624), .Y(n11749) );
  MX2XL U6428 ( .A(\I_cache/cache[6][135] ), .B(n11177), .S0(n5892), .Y(n11759) );
  MX2XL U6429 ( .A(\I_cache/cache[3][135] ), .B(n11177), .S0(n5670), .Y(n11762) );
  MX2XL U6430 ( .A(\I_cache/cache[2][135] ), .B(n11177), .S0(n5715), .Y(n11763) );
  MX2XL U6431 ( .A(\I_cache/cache[1][135] ), .B(n11177), .S0(n5581), .Y(n11764) );
  MX2XL U6432 ( .A(\I_cache/cache[0][135] ), .B(n11177), .S0(n5624), .Y(n11765) );
  MX2XL U6433 ( .A(\I_cache/cache[6][131] ), .B(n11159), .S0(n5892), .Y(n11791) );
  MX2XL U6434 ( .A(\I_cache/cache[3][131] ), .B(n11159), .S0(n5670), .Y(n11794) );
  MX2XL U6435 ( .A(\I_cache/cache[2][131] ), .B(n11159), .S0(n5715), .Y(n11795) );
  MX2XL U6436 ( .A(\I_cache/cache[1][131] ), .B(n11159), .S0(n5581), .Y(n11796) );
  MX2XL U6437 ( .A(\I_cache/cache[0][131] ), .B(n11159), .S0(n5624), .Y(n11797) );
  MX2XL U6438 ( .A(\I_cache/cache[6][129] ), .B(n11164), .S0(n5892), .Y(n11807) );
  MX2XL U6439 ( .A(\I_cache/cache[3][129] ), .B(n11164), .S0(n5670), .Y(n11810) );
  MX2XL U6440 ( .A(\I_cache/cache[2][129] ), .B(n11164), .S0(n5715), .Y(n11811) );
  MX2XL U6441 ( .A(\I_cache/cache[1][129] ), .B(n11164), .S0(n5581), .Y(n11812) );
  MX2XL U6442 ( .A(\I_cache/cache[0][129] ), .B(n11164), .S0(n5624), .Y(n11813) );
  MX2XL U6443 ( .A(\I_cache/cache[6][136] ), .B(n11182), .S0(n5892), .Y(n11751) );
  MX2XL U6444 ( .A(\I_cache/cache[3][136] ), .B(n11182), .S0(n5670), .Y(n11754) );
  MX2XL U6445 ( .A(\I_cache/cache[2][136] ), .B(n11182), .S0(n5715), .Y(n11755) );
  MX2XL U6446 ( .A(\I_cache/cache[1][136] ), .B(n11182), .S0(n5581), .Y(n11756) );
  MX2XL U6447 ( .A(\I_cache/cache[0][136] ), .B(n11182), .S0(n5624), .Y(n11757) );
  MX2XL U6448 ( .A(\I_cache/cache[6][148] ), .B(n11197), .S0(n5892), .Y(n11655) );
  MX2XL U6449 ( .A(\I_cache/cache[3][148] ), .B(n11197), .S0(n5670), .Y(n11658) );
  MX2XL U6450 ( .A(\I_cache/cache[2][148] ), .B(n11197), .S0(n5715), .Y(n11659) );
  MX2XL U6451 ( .A(\I_cache/cache[1][148] ), .B(n11197), .S0(n5581), .Y(n11660) );
  MX2XL U6452 ( .A(\I_cache/cache[0][148] ), .B(n11197), .S0(n5624), .Y(n11661) );
  MX2XL U6453 ( .A(\I_cache/cache[6][149] ), .B(n11187), .S0(n5892), .Y(n11647) );
  MX2XL U6454 ( .A(\I_cache/cache[3][149] ), .B(n11187), .S0(n5670), .Y(n11650) );
  MX2XL U6455 ( .A(\I_cache/cache[2][149] ), .B(n11187), .S0(n5715), .Y(n11651) );
  MX2XL U6456 ( .A(\I_cache/cache[1][149] ), .B(n11187), .S0(n5581), .Y(n11652) );
  MX2XL U6457 ( .A(\I_cache/cache[0][149] ), .B(n11187), .S0(n5624), .Y(n11653) );
  MX2XL U6458 ( .A(\I_cache/cache[6][147] ), .B(n11192), .S0(n5892), .Y(n11663) );
  MX2XL U6459 ( .A(\I_cache/cache[3][147] ), .B(n11192), .S0(n5670), .Y(n11666) );
  MX2XL U6460 ( .A(\I_cache/cache[2][147] ), .B(n11192), .S0(n5715), .Y(n11667) );
  MX2XL U6461 ( .A(\I_cache/cache[1][147] ), .B(n11192), .S0(n5581), .Y(n11668) );
  MX2XL U6462 ( .A(\I_cache/cache[0][147] ), .B(n11192), .S0(n5624), .Y(n11669) );
  MX2XL U6463 ( .A(\I_cache/cache[0][142] ), .B(n11201), .S0(n5624), .Y(n11709) );
  MX2XL U6464 ( .A(\I_cache/cache[2][134] ), .B(n11122), .S0(n5714), .Y(n11771) );
  MX2XL U6465 ( .A(\I_cache/cache[1][134] ), .B(n11122), .S0(n5580), .Y(n11772) );
  MX2XL U6466 ( .A(\I_cache/cache[0][134] ), .B(n11122), .S0(n5623), .Y(n11773) );
  MX2XL U6467 ( .A(\I_cache/cache[2][139] ), .B(n11140), .S0(n5714), .Y(n11731) );
  MX2XL U6468 ( .A(\I_cache/cache[1][139] ), .B(n11140), .S0(n5580), .Y(n11732) );
  MX2XL U6469 ( .A(\I_cache/cache[0][139] ), .B(n11140), .S0(n5623), .Y(n11733) );
  MX2XL U6470 ( .A(\I_cache/cache[2][133] ), .B(n11127), .S0(n5714), .Y(n11779) );
  MX2XL U6471 ( .A(\I_cache/cache[1][133] ), .B(n11127), .S0(n5580), .Y(n11780) );
  MX2XL U6472 ( .A(\I_cache/cache[0][133] ), .B(n11127), .S0(n5623), .Y(n11781) );
  MX2XL U6473 ( .A(\I_cache/cache[2][128] ), .B(n11067), .S0(n5714), .Y(n11819) );
  MX2XL U6474 ( .A(\I_cache/cache[1][128] ), .B(n11067), .S0(n5580), .Y(n11820) );
  MX2XL U6475 ( .A(\I_cache/cache[0][128] ), .B(n11067), .S0(n5623), .Y(n11821) );
  MX2XL U6476 ( .A(\I_cache/cache[2][138] ), .B(n11131), .S0(n5714), .Y(n11739) );
  MX2XL U6477 ( .A(\I_cache/cache[1][138] ), .B(n11131), .S0(n5580), .Y(n11740) );
  MX2XL U6478 ( .A(\I_cache/cache[0][138] ), .B(n11131), .S0(n5623), .Y(n11741) );
  MX2XL U6479 ( .A(\I_cache/cache[2][145] ), .B(n11065), .S0(n5716), .Y(n11683) );
  MX2XL U6480 ( .A(\I_cache/cache[0][145] ), .B(n11065), .S0(n5625), .Y(n11685) );
  MX2XL U6481 ( .A(\I_cache/cache[2][151] ), .B(n11066), .S0(n5714), .Y(n11635) );
  MX2XL U6482 ( .A(\I_cache/cache[0][151] ), .B(n11066), .S0(n5623), .Y(n11637) );
  MX2XL U6483 ( .A(\I_cache/cache[2][132] ), .B(n11118), .S0(n5714), .Y(n11787) );
  MX2XL U6484 ( .A(\I_cache/cache[1][132] ), .B(n11118), .S0(n5580), .Y(n11788) );
  MX2XL U6485 ( .A(\I_cache/cache[0][132] ), .B(n11118), .S0(n5623), .Y(n11789) );
  MX2XL U6486 ( .A(\I_cache/cache[6][134] ), .B(n11122), .S0(n5891), .Y(n11767) );
  MX2XL U6487 ( .A(\I_cache/cache[3][134] ), .B(n11122), .S0(n5669), .Y(n11770) );
  MX2XL U6488 ( .A(\I_cache/cache[6][139] ), .B(n11140), .S0(n5891), .Y(n11727) );
  MX2XL U6489 ( .A(\I_cache/cache[3][139] ), .B(n11140), .S0(n5669), .Y(n11730) );
  MX2XL U6490 ( .A(\I_cache/cache[3][133] ), .B(n11127), .S0(n5669), .Y(n11778) );
  MX2XL U6491 ( .A(\I_cache/cache[6][128] ), .B(n11067), .S0(n5891), .Y(n11815) );
  MX2XL U6492 ( .A(\I_cache/cache[3][128] ), .B(n11067), .S0(n5669), .Y(n11818) );
  MX2XL U6493 ( .A(\I_cache/cache[0][143] ), .B(n11215), .S0(n5619), .Y(n11701) );
  MX2XL U6494 ( .A(\I_cache/cache[6][138] ), .B(n11131), .S0(n5891), .Y(n11735) );
  MX2XL U6495 ( .A(\I_cache/cache[6][132] ), .B(n11118), .S0(n5891), .Y(n11783) );
  MX2XL U6496 ( .A(\I_cache/cache[3][132] ), .B(n11118), .S0(n5669), .Y(n11786) );
  MX2XL U6497 ( .A(\I_cache/cache[3][144] ), .B(n11145), .S0(n5668), .Y(n11690) );
  MX2XL U6498 ( .A(\I_cache/cache[2][144] ), .B(n11145), .S0(n5713), .Y(n11691) );
  MX2XL U6499 ( .A(\I_cache/cache[1][144] ), .B(n11145), .S0(n5579), .Y(n11692) );
  MX2XL U6500 ( .A(\I_cache/cache[0][144] ), .B(n11145), .S0(n5622), .Y(n11693) );
  MX2XL U6501 ( .A(\I_cache/cache[5][143] ), .B(n11215), .S0(n5754), .Y(n11696) );
  MX2XL U6502 ( .A(\I_cache/cache[4][143] ), .B(n11215), .S0(n5800), .Y(n11697) );
  MX2XL U6503 ( .A(\I_cache/cache[3][143] ), .B(n11215), .S0(n5665), .Y(n11698) );
  MX2XL U6504 ( .A(\I_cache/cache[2][143] ), .B(n11215), .S0(n5710), .Y(n11699) );
  MX2XL U6505 ( .A(\I_cache/cache[1][143] ), .B(n11215), .S0(n5576), .Y(n11700) );
  MX2XL U6506 ( .A(\I_cache/cache[7][146] ), .B(n11063), .S0(n5846), .Y(n11670) );
  MX2XL U6507 ( .A(\I_cache/cache[5][133] ), .B(n11127), .S0(n5758), .Y(n11776) );
  MX2XL U6508 ( .A(\I_cache/cache[4][133] ), .B(n11127), .S0(n5804), .Y(n11777) );
  MX2XL U6509 ( .A(\I_cache/cache[0][146] ), .B(n11063), .S0(n5624), .Y(n11677) );
  MX2XL U6510 ( .A(\I_cache/cache[0][150] ), .B(n11064), .S0(n5623), .Y(n11645) );
  MX2XL U6511 ( .A(\I_cache/cache[6][146] ), .B(n11063), .S0(n5888), .Y(n11671) );
  MX2XL U6512 ( .A(\I_cache/cache[5][146] ), .B(n11063), .S0(n5752), .Y(n11672) );
  MX2XL U6513 ( .A(\I_cache/cache[4][146] ), .B(n11063), .S0(n5802), .Y(n11673) );
  MX2XL U6514 ( .A(\I_cache/cache[3][146] ), .B(n11063), .S0(n5665), .Y(n11674) );
  MX2XL U6515 ( .A(\I_cache/cache[2][146] ), .B(n11063), .S0(n5708), .Y(n11675) );
  MX2XL U6516 ( .A(\I_cache/cache[1][146] ), .B(n11063), .S0(n5581), .Y(n11676) );
  MX2XL U6517 ( .A(\I_cache/cache[6][150] ), .B(n11064), .S0(n5886), .Y(n11639) );
  MX2XL U6518 ( .A(\I_cache/cache[5][150] ), .B(n11064), .S0(n5753), .Y(n11640) );
  MX2XL U6519 ( .A(\I_cache/cache[4][150] ), .B(n11064), .S0(n5800), .Y(n11641) );
  MX2XL U6520 ( .A(\I_cache/cache[3][150] ), .B(n11064), .S0(n5667), .Y(n11642) );
  MX2XL U6521 ( .A(\I_cache/cache[2][150] ), .B(n11064), .S0(n5710), .Y(n11643) );
  MX2XL U6522 ( .A(\I_cache/cache[1][150] ), .B(n11064), .S0(n5580), .Y(n11644) );
  XOR2XL U6523 ( .A(n10341), .B(ICACHE_addr[19]), .Y(n10338) );
  XOR2XL U6524 ( .A(n10481), .B(ICACHE_addr[11]), .Y(n10485) );
  XOR2XL U6525 ( .A(n10167), .B(ICACHE_addr[7]), .Y(n10162) );
  XOR2XL U6526 ( .A(n10324), .B(ICACHE_addr[18]), .Y(n10328) );
  NAND2XL U6527 ( .A(n10333), .B(ICACHE_addr[17]), .Y(n10324) );
  XOR2XL U6528 ( .A(n10472), .B(ICACHE_addr[10]), .Y(n10477) );
  XOR2XL U6529 ( .A(n10147), .B(ICACHE_addr[6]), .Y(n10151) );
  XOR2XL U6530 ( .A(n10168), .B(ICACHE_addr[8]), .Y(n10172) );
  XOR2XL U6531 ( .A(n10293), .B(ICACHE_addr[16]), .Y(n10298) );
  NAND2XL U6532 ( .A(n10301), .B(ICACHE_addr[15]), .Y(n10293) );
  XOR2XL U6533 ( .A(n10273), .B(ICACHE_addr[14]), .Y(n10277) );
  NAND2XL U6534 ( .A(n10282), .B(ICACHE_addr[13]), .Y(n10273) );
  AOI21XL U6535 ( .A0(\i_MIPS/IF_ID[23] ), .A1(\i_MIPS/Sign_Extend[31] ), .B0(
        n4811), .Y(n4805) );
  XOR2XL U6536 ( .A(n10292), .B(ICACHE_addr[15]), .Y(n10286) );
  XOR2XL U6537 ( .A(n10323), .B(ICACHE_addr[17]), .Y(n10305) );
  XOR2XL U6538 ( .A(n10272), .B(ICACHE_addr[13]), .Y(n10269) );
  XOR2XL U6539 ( .A(n10265), .B(ICACHE_addr[9]), .Y(n10183) );
  NAND2XL U6540 ( .A(n12971), .B(\i_MIPS/n266 ), .Y(n10110) );
  NAND2XL U6541 ( .A(n12961), .B(n5190), .Y(net105311) );
  NAND2XL U6542 ( .A(n12959), .B(n5190), .Y(net105264) );
  NAND2XL U6543 ( .A(n12956), .B(n5190), .Y(net105075) );
  NAND2XL U6544 ( .A(n12970), .B(n5190), .Y(net105255) );
  NAND2XL U6545 ( .A(n12969), .B(\i_MIPS/n266 ), .Y(net105165) );
  NAND2XL U6546 ( .A(n12966), .B(\i_MIPS/n266 ), .Y(net105662) );
  NAND2XL U6547 ( .A(n12973), .B(\i_MIPS/n266 ), .Y(net105232) );
  NAND2XL U6548 ( .A(n12974), .B(\i_MIPS/n266 ), .Y(net104721) );
  NAND2XL U6549 ( .A(\i_MIPS/EX_MEM[6] ), .B(\i_MIPS/n266 ), .Y(net104916) );
  OA22XL U6550 ( .A0(\i_MIPS/Register/register[4][30] ), .A1(n5099), .B0(
        \i_MIPS/Register/register[12][30] ), .B1(n5096), .Y(n9391) );
  OA22XL U6551 ( .A0(\i_MIPS/Register/register[20][30] ), .A1(n5099), .B0(
        \i_MIPS/Register/register[28][30] ), .B1(n5096), .Y(n9400) );
  OA22XL U6552 ( .A0(\i_MIPS/Register/register[4][31] ), .A1(n5101), .B0(
        \i_MIPS/Register/register[12][31] ), .B1(n5096), .Y(n9496) );
  OA22XL U6553 ( .A0(\i_MIPS/Register/register[20][31] ), .A1(n5099), .B0(
        \i_MIPS/Register/register[28][31] ), .B1(n5096), .Y(n9513) );
  OA22XL U6554 ( .A0(\i_MIPS/Register/register[0][24] ), .A1(n5106), .B0(
        \i_MIPS/Register/register[8][24] ), .B1(n5103), .Y(n6617) );
  OA22XL U6555 ( .A0(n5813), .A1(n1592), .B0(n5768), .B1(n3279), .Y(n9656) );
  OA22XL U6556 ( .A0(\i_MIPS/Register/register[0][30] ), .A1(n5107), .B0(
        \i_MIPS/Register/register[8][30] ), .B1(n5105), .Y(n9390) );
  OA22XL U6557 ( .A0(\i_MIPS/Register/register[16][30] ), .A1(n5108), .B0(
        \i_MIPS/Register/register[24][30] ), .B1(n5105), .Y(n9399) );
  OA22XL U6558 ( .A0(\i_MIPS/Register/register[0][31] ), .A1(n5107), .B0(
        \i_MIPS/Register/register[8][31] ), .B1(n5105), .Y(n9495) );
  OA22XL U6559 ( .A0(\i_MIPS/Register/register[16][31] ), .A1(n5108), .B0(
        \i_MIPS/Register/register[24][31] ), .B1(n5105), .Y(n9512) );
  AO21XL U6560 ( .A0(n5842), .A1(n11586), .B0(\I_cache/cache[7][154] ), .Y(
        n11606) );
  AO21XL U6561 ( .A0(n5624), .A1(n11586), .B0(\I_cache/cache[0][154] ), .Y(
        n11613) );
  AO21XL U6562 ( .A0(n5889), .A1(n11586), .B0(\I_cache/cache[6][154] ), .Y(
        n11607) );
  AO21XL U6563 ( .A0(n4831), .A1(n11586), .B0(\I_cache/cache[5][154] ), .Y(
        n11608) );
  AO21XL U6564 ( .A0(n5799), .A1(n11586), .B0(\I_cache/cache[4][154] ), .Y(
        n11609) );
  AO21XL U6565 ( .A0(n5663), .A1(n11586), .B0(\I_cache/cache[3][154] ), .Y(
        n11610) );
  AO21XL U6566 ( .A0(n5709), .A1(n11586), .B0(\I_cache/cache[2][154] ), .Y(
        n11611) );
  AO21XL U6567 ( .A0(n5580), .A1(n11586), .B0(\I_cache/cache[1][154] ), .Y(
        n11612) );
  AND2XL U6568 ( .A(\i_MIPS/IF_ID[19] ), .B(n6016), .Y(n4812) );
  AND2XL U6569 ( .A(\i_MIPS/IF_ID[22] ), .B(n6016), .Y(n4811) );
  AND2XL U6570 ( .A(\i_MIPS/IF_ID[24] ), .B(n6016), .Y(n4820) );
  AND2X1 U6571 ( .A(\i_MIPS/IF_ID[18] ), .B(n6016), .Y(n4822) );
  AND2XL U6572 ( .A(\i_MIPS/IF_ID[21] ), .B(n6016), .Y(n4821) );
  NAND3BXL U6573 ( .AN(n9823), .B(\i_MIPS/IR[31] ), .C(n9812), .Y(
        \i_MIPS/Control/n10 ) );
  AND3XL U6574 ( .A(n9821), .B(n9811), .C(n9820), .Y(n9812) );
  XOR2XL U6575 ( .A(n9936), .B(ICACHE_addr[4]), .Y(n10871) );
  XOR2XL U6576 ( .A(n10051), .B(ICACHE_addr[3]), .Y(n10913) );
  XOR2XL U6577 ( .A(n10146), .B(ICACHE_addr[5]), .Y(n10142) );
  XOR2XL U6578 ( .A(n9802), .B(ICACHE_addr[2]), .Y(n10936) );
  XOR2XL U6579 ( .A(\i_MIPS/n506 ), .B(\i_MIPS/jump_addr[31] ), .Y(n10724) );
  NAND4XL U6580 ( .A(n9821), .B(n9820), .C(\i_MIPS/IR[31] ), .D(
        \i_MIPS/IR[29] ), .Y(n9822) );
  NAND2XL U6581 ( .A(\i_MIPS/jump_addr[30] ), .B(n6016), .Y(n10725) );
  NAND2XL U6582 ( .A(\i_MIPS/jump_addr[29] ), .B(n6016), .Y(n10579) );
  INVXL U6583 ( .A(\i_MIPS/IR[30] ), .Y(n9821) );
  AO21XL U6584 ( .A0(n3031), .A1(n5419), .B0(\D_cache/cache[7][154] ), .Y(
        \D_cache/n557 ) );
  AO21XL U6585 ( .A0(n3031), .A1(n3574), .B0(\D_cache/cache[6][154] ), .Y(
        \D_cache/n558 ) );
  AO21XL U6586 ( .A0(n3031), .A1(n5350), .B0(\D_cache/cache[5][154] ), .Y(
        \D_cache/n559 ) );
  AO21XL U6587 ( .A0(n3031), .A1(n5323), .B0(\D_cache/cache[4][154] ), .Y(
        \D_cache/n560 ) );
  AO21XL U6588 ( .A0(n3031), .A1(n5276), .B0(\D_cache/cache[3][154] ), .Y(
        \D_cache/n561 ) );
  AO21XL U6589 ( .A0(n3031), .A1(n5236), .B0(\D_cache/cache[2][154] ), .Y(
        \D_cache/n562 ) );
  AO21XL U6590 ( .A0(n3031), .A1(n5208), .B0(\D_cache/cache[1][154] ), .Y(
        \D_cache/n563 ) );
  AO21XL U6591 ( .A0(n3031), .A1(n5168), .B0(\D_cache/cache[0][154] ), .Y(
        \D_cache/n564 ) );
  INVXL U6592 ( .A(\i_MIPS/n497 ), .Y(n10378) );
  CLKBUFX3 U6593 ( .A(net115813), .Y(net115795) );
  CLKBUFX3 U6594 ( .A(n10797), .Y(n5530) );
  CLKBUFX3 U6595 ( .A(n10797), .Y(n5529) );
  INVX3 U6596 ( .A(n5238), .Y(n5234) );
  INVX3 U6597 ( .A(n5240), .Y(n5232) );
  INVX3 U6598 ( .A(n5243), .Y(n5228) );
  INVX3 U6599 ( .A(n5242), .Y(n5233) );
  INVX3 U6600 ( .A(n5237), .Y(n5235) );
  INVX3 U6601 ( .A(n5242), .Y(n5230) );
  INVX3 U6602 ( .A(n5241), .Y(n5231) );
  INVX3 U6603 ( .A(n5673), .Y(n5664) );
  INVX3 U6604 ( .A(n5673), .Y(n5663) );
  INVX3 U6605 ( .A(n5284), .Y(n5268) );
  INVX3 U6606 ( .A(n5283), .Y(n5269) );
  INVX3 U6607 ( .A(n5279), .Y(n5274) );
  INVX3 U6608 ( .A(n5277), .Y(n5275) );
  INVX3 U6609 ( .A(n5282), .Y(n5270) );
  INVX3 U6610 ( .A(n5281), .Y(n5272) );
  INVX3 U6611 ( .A(n5280), .Y(n5273) );
  INVX3 U6612 ( .A(n5299), .Y(n5276) );
  CLKBUFX3 U6613 ( .A(n5542), .Y(n5546) );
  CLKBUFX3 U6614 ( .A(n10974), .Y(n5544) );
  CLKBUFX3 U6615 ( .A(n5542), .Y(n5547) );
  CLKBUFX3 U6616 ( .A(n10974), .Y(n5548) );
  CLKBUFX3 U6617 ( .A(n10974), .Y(n5549) );
  CLKBUFX3 U6618 ( .A(n5928), .Y(n5895) );
  CLKBUFX3 U6619 ( .A(n5928), .Y(n5894) );
  CLKBUFX3 U6620 ( .A(n5405), .Y(n5378) );
  CLKBUFX3 U6621 ( .A(n5405), .Y(n5377) );
  CLKBUFX3 U6622 ( .A(n5398), .Y(n5383) );
  CLKBUFX3 U6623 ( .A(n5394), .Y(n5382) );
  CLKBUFX3 U6624 ( .A(n5392), .Y(n5384) );
  CLKBUFX3 U6625 ( .A(n5405), .Y(n5379) );
  CLKBUFX3 U6626 ( .A(n5405), .Y(n5380) );
  CLKBUFX3 U6627 ( .A(n5406), .Y(n5375) );
  CLKBUFX3 U6628 ( .A(n5927), .Y(n5896) );
  CLKBUFX3 U6629 ( .A(n5704), .Y(n5672) );
  CLKBUFX3 U6630 ( .A(n5452), .Y(n5422) );
  CLKBUFX3 U6631 ( .A(n5702), .Y(n5673) );
  CLKBUFX3 U6632 ( .A(n5924), .Y(n5908) );
  CLKBUFX3 U6633 ( .A(n5923), .Y(n5909) );
  CLKBUFX3 U6634 ( .A(n5925), .Y(n5903) );
  CLKBUFX3 U6635 ( .A(n5923), .Y(n5910) );
  CLKBUFX3 U6636 ( .A(n5922), .Y(n5913) );
  CLKBUFX3 U6637 ( .A(n5923), .Y(n5912) );
  CLKBUFX3 U6638 ( .A(n5923), .Y(n5911) );
  CLKBUFX3 U6639 ( .A(n5925), .Y(n5904) );
  CLKBUFX3 U6640 ( .A(n5924), .Y(n5905) );
  CLKBUFX3 U6641 ( .A(n5924), .Y(n5906) );
  CLKBUFX3 U6642 ( .A(n5924), .Y(n5907) );
  CLKBUFX3 U6643 ( .A(n5925), .Y(n5902) );
  CLKBUFX3 U6644 ( .A(n5922), .Y(n5914) );
  CLKBUFX3 U6645 ( .A(n5922), .Y(n5916) );
  CLKBUFX3 U6646 ( .A(n5922), .Y(n5915) );
  CLKBUFX3 U6647 ( .A(n5926), .Y(n5897) );
  CLKBUFX3 U6648 ( .A(n5925), .Y(n5901) );
  CLKBUFX3 U6649 ( .A(n5926), .Y(n5900) );
  CLKBUFX3 U6650 ( .A(n5926), .Y(n5899) );
  CLKBUFX3 U6651 ( .A(n5926), .Y(n5898) );
  CLKBUFX3 U6652 ( .A(n5450), .Y(n5426) );
  CLKBUFX3 U6653 ( .A(n5450), .Y(n5427) );
  CLKBUFX3 U6654 ( .A(n5445), .Y(n5435) );
  CLKBUFX3 U6655 ( .A(n5448), .Y(n5434) );
  CLKBUFX3 U6656 ( .A(n5453), .Y(n5443) );
  CLKBUFX3 U6657 ( .A(n5699), .Y(n5685) );
  CLKBUFX3 U6658 ( .A(n5698), .Y(n5686) );
  CLKBUFX3 U6659 ( .A(n5700), .Y(n5680) );
  CLKBUFX3 U6660 ( .A(n5698), .Y(n5687) );
  CLKBUFX3 U6661 ( .A(n5697), .Y(n5690) );
  CLKBUFX3 U6662 ( .A(n5698), .Y(n5689) );
  CLKBUFX3 U6663 ( .A(n5698), .Y(n5688) );
  CLKBUFX3 U6664 ( .A(n5700), .Y(n5681) );
  CLKBUFX3 U6665 ( .A(n5699), .Y(n5682) );
  CLKBUFX3 U6666 ( .A(n5699), .Y(n5683) );
  CLKBUFX3 U6667 ( .A(n5699), .Y(n5684) );
  CLKBUFX3 U6668 ( .A(n5700), .Y(n5679) );
  CLKBUFX3 U6669 ( .A(n5697), .Y(n5691) );
  CLKBUFX3 U6670 ( .A(n5697), .Y(n5693) );
  CLKBUFX3 U6671 ( .A(n5697), .Y(n5692) );
  CLKBUFX3 U6672 ( .A(n5701), .Y(n5674) );
  CLKBUFX3 U6673 ( .A(n5700), .Y(n5678) );
  CLKBUFX3 U6674 ( .A(n5701), .Y(n5677) );
  CLKBUFX3 U6675 ( .A(n5701), .Y(n5676) );
  CLKBUFX3 U6676 ( .A(n5701), .Y(n5675) );
  INVX3 U6677 ( .A(n5111), .Y(n5108) );
  INVX3 U6678 ( .A(n5110), .Y(n5109) );
  INVX3 U6679 ( .A(n5111), .Y(n5107) );
  INVX3 U6680 ( .A(n5112), .Y(n5106) );
  INVX3 U6681 ( .A(n5628), .Y(n5624) );
  INVX3 U6682 ( .A(n5629), .Y(n5623) );
  INVX3 U6683 ( .A(n5809), .Y(n5799) );
  INVX3 U6684 ( .A(n5630), .Y(n5618) );
  INVX3 U6685 ( .A(n5734), .Y(n5709) );
  INVX3 U6686 ( .A(n5638), .Y(n5619) );
  INVX3 U6687 ( .A(n5630), .Y(n5620) );
  INVX3 U6688 ( .A(n5630), .Y(n5621) );
  INVX3 U6689 ( .A(n5630), .Y(n5622) );
  INVX3 U6690 ( .A(n5630), .Y(n5617) );
  INVX3 U6691 ( .A(n5823), .Y(n5798) );
  INVX3 U6692 ( .A(n5720), .Y(n5708) );
  INVX3 U6693 ( .A(n5627), .Y(n5625) );
  INVX3 U6694 ( .A(n5584), .Y(n5581) );
  INVX3 U6695 ( .A(n5760), .Y(n5758) );
  INVX3 U6696 ( .A(n5585), .Y(n5580) );
  INVX3 U6697 ( .A(n5854), .Y(n5843) );
  INVX3 U6698 ( .A(n5764), .Y(n5752) );
  INVX3 U6699 ( .A(n5764), .Y(n5753) );
  INVX3 U6700 ( .A(n5595), .Y(n5575) );
  INVX3 U6701 ( .A(n5588), .Y(n5576) );
  INVX3 U6702 ( .A(n5596), .Y(n5577) );
  INVX3 U6703 ( .A(n5762), .Y(n5756) );
  INVX3 U6704 ( .A(n5586), .Y(n5578) );
  INVX3 U6705 ( .A(n5766), .Y(n5755) );
  INVX3 U6706 ( .A(n5761), .Y(n5757) );
  INVX3 U6707 ( .A(n5587), .Y(n5579) );
  INVX3 U6708 ( .A(n5854), .Y(n5842) );
  INVX3 U6709 ( .A(n5586), .Y(n5574) );
  INVX3 U6710 ( .A(n5764), .Y(n5759) );
  INVX3 U6711 ( .A(n5594), .Y(n5582) );
  CLKBUFX3 U6712 ( .A(n6355), .Y(n6045) );
  CLKBUFX3 U6713 ( .A(n6355), .Y(n6046) );
  CLKBUFX3 U6714 ( .A(n6355), .Y(n6047) );
  CLKBUFX3 U6715 ( .A(n6355), .Y(n6048) );
  CLKBUFX3 U6716 ( .A(n6355), .Y(n6049) );
  CLKBUFX3 U6717 ( .A(n6355), .Y(n6050) );
  CLKBUFX3 U6718 ( .A(n6355), .Y(n6051) );
  CLKBUFX3 U6719 ( .A(n6355), .Y(n6052) );
  CLKBUFX3 U6720 ( .A(n6355), .Y(n6053) );
  CLKBUFX3 U6721 ( .A(n6355), .Y(n6054) );
  CLKBUFX3 U6722 ( .A(n6355), .Y(n6055) );
  CLKBUFX3 U6723 ( .A(n6355), .Y(n6056) );
  CLKBUFX3 U6724 ( .A(n6354), .Y(n6057) );
  CLKBUFX3 U6725 ( .A(n6354), .Y(n6058) );
  CLKBUFX3 U6726 ( .A(n6354), .Y(n6059) );
  CLKBUFX3 U6727 ( .A(n6354), .Y(n6060) );
  CLKBUFX3 U6728 ( .A(n6354), .Y(n6061) );
  CLKBUFX3 U6729 ( .A(n6354), .Y(n6062) );
  CLKBUFX3 U6730 ( .A(n6354), .Y(n6063) );
  CLKBUFX3 U6731 ( .A(n6354), .Y(n6064) );
  CLKBUFX3 U6732 ( .A(n6354), .Y(n6065) );
  CLKBUFX3 U6733 ( .A(n6354), .Y(n6066) );
  CLKBUFX3 U6734 ( .A(n6354), .Y(n6067) );
  CLKBUFX3 U6735 ( .A(n6354), .Y(n6068) );
  CLKBUFX3 U6736 ( .A(n6353), .Y(n6069) );
  CLKBUFX3 U6737 ( .A(n6353), .Y(n6070) );
  CLKBUFX3 U6738 ( .A(n6353), .Y(n6071) );
  CLKBUFX3 U6739 ( .A(n6353), .Y(n6072) );
  CLKBUFX3 U6740 ( .A(n6353), .Y(n6073) );
  CLKBUFX3 U6741 ( .A(n6353), .Y(n6074) );
  CLKBUFX3 U6742 ( .A(n6353), .Y(n6075) );
  CLKBUFX3 U6743 ( .A(n6353), .Y(n6076) );
  CLKBUFX3 U6744 ( .A(n6353), .Y(n6077) );
  CLKBUFX3 U6745 ( .A(n6353), .Y(n6078) );
  CLKBUFX3 U6746 ( .A(n6353), .Y(n6079) );
  CLKBUFX3 U6747 ( .A(n6353), .Y(n6080) );
  CLKBUFX3 U6748 ( .A(n6352), .Y(n6081) );
  CLKBUFX3 U6749 ( .A(n6352), .Y(n6082) );
  CLKBUFX3 U6750 ( .A(n6352), .Y(n6083) );
  CLKBUFX3 U6751 ( .A(n6352), .Y(n6084) );
  CLKBUFX3 U6752 ( .A(n6352), .Y(n6085) );
  CLKBUFX3 U6753 ( .A(n6352), .Y(n6086) );
  CLKBUFX3 U6754 ( .A(n6352), .Y(n6087) );
  CLKBUFX3 U6755 ( .A(n6352), .Y(n6088) );
  CLKBUFX3 U6756 ( .A(n6352), .Y(n6089) );
  CLKBUFX3 U6757 ( .A(n6352), .Y(n6090) );
  CLKBUFX3 U6758 ( .A(n6352), .Y(n6091) );
  CLKBUFX3 U6759 ( .A(n6352), .Y(n6092) );
  CLKBUFX3 U6760 ( .A(n6351), .Y(n6093) );
  CLKBUFX3 U6761 ( .A(n6351), .Y(n6094) );
  CLKBUFX3 U6762 ( .A(n6351), .Y(n6095) );
  CLKBUFX3 U6763 ( .A(n6351), .Y(n6096) );
  CLKBUFX3 U6764 ( .A(n6351), .Y(n6097) );
  CLKBUFX3 U6765 ( .A(n6351), .Y(n6098) );
  CLKBUFX3 U6766 ( .A(n6351), .Y(n6099) );
  CLKBUFX3 U6767 ( .A(n6351), .Y(n6100) );
  CLKBUFX3 U6768 ( .A(n6351), .Y(n6101) );
  CLKBUFX3 U6769 ( .A(n6351), .Y(n6102) );
  CLKBUFX3 U6770 ( .A(n6351), .Y(n6103) );
  CLKBUFX3 U6771 ( .A(n6351), .Y(n6104) );
  CLKBUFX3 U6772 ( .A(n6350), .Y(n6105) );
  CLKBUFX3 U6773 ( .A(n6350), .Y(n6106) );
  CLKBUFX3 U6774 ( .A(n6350), .Y(n6107) );
  CLKBUFX3 U6775 ( .A(n6350), .Y(n6108) );
  CLKBUFX3 U6776 ( .A(n6350), .Y(n6109) );
  CLKBUFX3 U6777 ( .A(n6350), .Y(n6110) );
  CLKBUFX3 U6778 ( .A(n6350), .Y(n6111) );
  CLKBUFX3 U6779 ( .A(n6350), .Y(n6112) );
  CLKBUFX3 U6780 ( .A(n6350), .Y(n6113) );
  CLKBUFX3 U6781 ( .A(n6350), .Y(n6114) );
  CLKBUFX3 U6782 ( .A(n6350), .Y(n6115) );
  CLKBUFX3 U6783 ( .A(n6350), .Y(n6116) );
  CLKBUFX3 U6784 ( .A(n6349), .Y(n6117) );
  CLKBUFX3 U6785 ( .A(n6349), .Y(n6118) );
  CLKBUFX3 U6786 ( .A(n6349), .Y(n6119) );
  CLKBUFX3 U6787 ( .A(n6341), .Y(n6224) );
  CLKBUFX3 U6788 ( .A(n6340), .Y(n6225) );
  CLKBUFX3 U6789 ( .A(n6340), .Y(n6226) );
  CLKBUFX3 U6790 ( .A(n6340), .Y(n6227) );
  CLKBUFX3 U6791 ( .A(n6340), .Y(n6228) );
  CLKBUFX3 U6792 ( .A(n6340), .Y(n6229) );
  CLKBUFX3 U6793 ( .A(n6340), .Y(n6230) );
  CLKBUFX3 U6794 ( .A(n6340), .Y(n6231) );
  CLKBUFX3 U6795 ( .A(n6340), .Y(n6232) );
  CLKBUFX3 U6796 ( .A(n6340), .Y(n6233) );
  CLKBUFX3 U6797 ( .A(n6340), .Y(n6234) );
  CLKBUFX3 U6798 ( .A(n6340), .Y(n6235) );
  CLKBUFX3 U6799 ( .A(n6340), .Y(n6236) );
  CLKBUFX3 U6800 ( .A(n6339), .Y(n6237) );
  CLKBUFX3 U6801 ( .A(n6339), .Y(n6238) );
  CLKBUFX3 U6802 ( .A(n6339), .Y(n6239) );
  CLKBUFX3 U6803 ( .A(n6339), .Y(n6240) );
  CLKBUFX3 U6804 ( .A(n6339), .Y(n6241) );
  CLKBUFX3 U6805 ( .A(n6339), .Y(n6242) );
  CLKBUFX3 U6806 ( .A(n6339), .Y(n6243) );
  CLKBUFX3 U6807 ( .A(n6339), .Y(n6244) );
  CLKBUFX3 U6808 ( .A(n6339), .Y(n6245) );
  CLKBUFX3 U6809 ( .A(n6339), .Y(n6246) );
  CLKBUFX3 U6810 ( .A(n6339), .Y(n6247) );
  CLKBUFX3 U6811 ( .A(n6339), .Y(n6248) );
  CLKBUFX3 U6812 ( .A(n6338), .Y(n6249) );
  CLKBUFX3 U6813 ( .A(n6338), .Y(n6250) );
  CLKBUFX3 U6814 ( .A(n6338), .Y(n6251) );
  CLKBUFX3 U6815 ( .A(n6338), .Y(n6252) );
  CLKBUFX3 U6816 ( .A(n6338), .Y(n6253) );
  CLKBUFX3 U6817 ( .A(n6338), .Y(n6254) );
  CLKBUFX3 U6818 ( .A(n6338), .Y(n6255) );
  CLKBUFX3 U6819 ( .A(n6338), .Y(n6256) );
  CLKBUFX3 U6820 ( .A(n6338), .Y(n6257) );
  CLKBUFX3 U6821 ( .A(n6338), .Y(n6258) );
  CLKBUFX3 U6822 ( .A(n6338), .Y(n6259) );
  CLKBUFX3 U6823 ( .A(n6338), .Y(n6260) );
  CLKBUFX3 U6824 ( .A(n6337), .Y(n6261) );
  CLKBUFX3 U6825 ( .A(n6337), .Y(n6262) );
  CLKBUFX3 U6826 ( .A(n6337), .Y(n6263) );
  CLKBUFX3 U6827 ( .A(n6337), .Y(n6264) );
  CLKBUFX3 U6828 ( .A(n6337), .Y(n6265) );
  CLKBUFX3 U6829 ( .A(n6337), .Y(n6266) );
  CLKBUFX3 U6830 ( .A(n6337), .Y(n6267) );
  CLKBUFX3 U6831 ( .A(n6337), .Y(n6268) );
  CLKBUFX3 U6832 ( .A(n6337), .Y(n6269) );
  CLKBUFX3 U6833 ( .A(n6337), .Y(n6270) );
  CLKBUFX3 U6834 ( .A(n6337), .Y(n6271) );
  CLKBUFX3 U6835 ( .A(n6337), .Y(n6272) );
  CLKBUFX3 U6836 ( .A(n6336), .Y(n6273) );
  CLKBUFX3 U6837 ( .A(n6336), .Y(n6274) );
  CLKBUFX3 U6838 ( .A(n6336), .Y(n6275) );
  CLKBUFX3 U6839 ( .A(n6336), .Y(n6276) );
  CLKBUFX3 U6840 ( .A(n6336), .Y(n6277) );
  CLKBUFX3 U6841 ( .A(n6336), .Y(n6278) );
  CLKBUFX3 U6842 ( .A(n6336), .Y(n6279) );
  CLKBUFX3 U6843 ( .A(n6336), .Y(n6280) );
  CLKBUFX3 U6844 ( .A(n6336), .Y(n6281) );
  CLKBUFX3 U6845 ( .A(n6336), .Y(n6282) );
  CLKBUFX3 U6846 ( .A(n6336), .Y(n6283) );
  CLKBUFX3 U6847 ( .A(n6336), .Y(n6284) );
  CLKBUFX3 U6848 ( .A(n6335), .Y(n6285) );
  CLKBUFX3 U6849 ( .A(n6335), .Y(n6286) );
  CLKBUFX3 U6850 ( .A(n6335), .Y(n6287) );
  CLKBUFX3 U6851 ( .A(n6335), .Y(n6288) );
  CLKBUFX3 U6852 ( .A(n6335), .Y(n6289) );
  CLKBUFX3 U6853 ( .A(n6335), .Y(n6290) );
  CLKBUFX3 U6854 ( .A(n6335), .Y(n6291) );
  CLKBUFX3 U6855 ( .A(n6335), .Y(n6292) );
  CLKBUFX3 U6856 ( .A(n6335), .Y(n6293) );
  CLKBUFX3 U6857 ( .A(n6335), .Y(n6294) );
  CLKBUFX3 U6858 ( .A(n6335), .Y(n6295) );
  CLKBUFX3 U6859 ( .A(n6335), .Y(n6296) );
  CLKBUFX3 U6860 ( .A(rst_n), .Y(n6297) );
  CLKBUFX3 U6861 ( .A(n6343), .Y(n6298) );
  CLKBUFX3 U6862 ( .A(n6336), .Y(n6299) );
  CLKBUFX3 U6863 ( .A(n6353), .Y(n6300) );
  CLKBUFX3 U6864 ( .A(n6341), .Y(n6301) );
  CLKBUFX3 U6865 ( .A(n6340), .Y(n6302) );
  CLKBUFX3 U6866 ( .A(n6337), .Y(n6303) );
  CLKBUFX3 U6867 ( .A(n6357), .Y(n6304) );
  CLKBUFX3 U6868 ( .A(n6332), .Y(n6305) );
  CLKBUFX3 U6869 ( .A(n6350), .Y(n6306) );
  CLKBUFX3 U6870 ( .A(n6343), .Y(n6307) );
  CLKBUFX3 U6871 ( .A(n6345), .Y(n6308) );
  CLKBUFX3 U6872 ( .A(n6334), .Y(n6309) );
  CLKBUFX3 U6873 ( .A(n6334), .Y(n6310) );
  CLKBUFX3 U6874 ( .A(n6349), .Y(n6120) );
  CLKBUFX3 U6875 ( .A(n6349), .Y(n6121) );
  CLKBUFX3 U6876 ( .A(n6349), .Y(n6122) );
  CLKBUFX3 U6877 ( .A(n6349), .Y(n6123) );
  CLKBUFX3 U6878 ( .A(n6349), .Y(n6124) );
  CLKBUFX3 U6879 ( .A(n6349), .Y(n6125) );
  CLKBUFX3 U6880 ( .A(n6349), .Y(n6126) );
  CLKBUFX3 U6881 ( .A(n6349), .Y(n6127) );
  CLKBUFX3 U6882 ( .A(n6349), .Y(n6128) );
  CLKBUFX3 U6883 ( .A(n6348), .Y(n6129) );
  CLKBUFX3 U6884 ( .A(n6348), .Y(n6130) );
  CLKBUFX3 U6885 ( .A(n6348), .Y(n6131) );
  CLKBUFX3 U6886 ( .A(n6348), .Y(n6132) );
  CLKBUFX3 U6887 ( .A(n6348), .Y(n6133) );
  CLKBUFX3 U6888 ( .A(n6348), .Y(n6134) );
  CLKBUFX3 U6889 ( .A(n6348), .Y(n6135) );
  CLKBUFX3 U6890 ( .A(n6348), .Y(n6136) );
  CLKBUFX3 U6891 ( .A(n6348), .Y(n6137) );
  CLKBUFX3 U6892 ( .A(n6348), .Y(n6138) );
  CLKBUFX3 U6893 ( .A(n6348), .Y(n6139) );
  CLKBUFX3 U6894 ( .A(n6348), .Y(n6140) );
  CLKBUFX3 U6895 ( .A(n6347), .Y(n6141) );
  CLKBUFX3 U6896 ( .A(n6347), .Y(n6142) );
  CLKBUFX3 U6897 ( .A(n6347), .Y(n6143) );
  CLKBUFX3 U6898 ( .A(n6347), .Y(n6144) );
  CLKBUFX3 U6899 ( .A(n6347), .Y(n6145) );
  CLKBUFX3 U6900 ( .A(n6347), .Y(n6146) );
  CLKBUFX3 U6901 ( .A(n6347), .Y(n6147) );
  CLKBUFX3 U6902 ( .A(n6347), .Y(n6148) );
  CLKBUFX3 U6903 ( .A(n6347), .Y(n6149) );
  CLKBUFX3 U6904 ( .A(n6347), .Y(n6150) );
  CLKBUFX3 U6905 ( .A(n6347), .Y(n6151) );
  CLKBUFX3 U6906 ( .A(n6347), .Y(n6152) );
  CLKBUFX3 U6907 ( .A(n6346), .Y(n6153) );
  CLKBUFX3 U6908 ( .A(n6346), .Y(n6154) );
  CLKBUFX3 U6909 ( .A(n6346), .Y(n6155) );
  CLKBUFX3 U6910 ( .A(n6346), .Y(n6156) );
  CLKBUFX3 U6911 ( .A(n6346), .Y(n6157) );
  CLKBUFX3 U6912 ( .A(n6346), .Y(n6158) );
  CLKBUFX3 U6913 ( .A(n6346), .Y(n6159) );
  CLKBUFX3 U6914 ( .A(n6346), .Y(n6160) );
  CLKBUFX3 U6915 ( .A(n6346), .Y(n6161) );
  CLKBUFX3 U6916 ( .A(n6346), .Y(n6162) );
  CLKBUFX3 U6917 ( .A(n6346), .Y(n6163) );
  CLKBUFX3 U6918 ( .A(n6346), .Y(n6164) );
  CLKBUFX3 U6919 ( .A(n6345), .Y(n6165) );
  CLKBUFX3 U6920 ( .A(n6345), .Y(n6166) );
  CLKBUFX3 U6921 ( .A(n6345), .Y(n6167) );
  CLKBUFX3 U6922 ( .A(n6345), .Y(n6168) );
  CLKBUFX3 U6923 ( .A(n6345), .Y(n6169) );
  CLKBUFX3 U6924 ( .A(n6345), .Y(n6170) );
  CLKBUFX3 U6925 ( .A(n6345), .Y(n6171) );
  CLKBUFX3 U6926 ( .A(n6345), .Y(n6172) );
  CLKBUFX3 U6927 ( .A(n6345), .Y(n6173) );
  CLKBUFX3 U6928 ( .A(n6345), .Y(n6174) );
  CLKBUFX3 U6929 ( .A(n6345), .Y(n6175) );
  CLKBUFX3 U6930 ( .A(n6345), .Y(n6176) );
  CLKBUFX3 U6931 ( .A(n6344), .Y(n6177) );
  CLKBUFX3 U6932 ( .A(n6344), .Y(n6178) );
  CLKBUFX3 U6933 ( .A(n6344), .Y(n6179) );
  CLKBUFX3 U6934 ( .A(n6344), .Y(n6180) );
  CLKBUFX3 U6935 ( .A(n6344), .Y(n6181) );
  CLKBUFX3 U6936 ( .A(n6344), .Y(n6182) );
  CLKBUFX3 U6937 ( .A(n6344), .Y(n6183) );
  CLKBUFX3 U6938 ( .A(n6344), .Y(n6184) );
  CLKBUFX3 U6939 ( .A(n6344), .Y(n6185) );
  CLKBUFX3 U6940 ( .A(n6344), .Y(n6186) );
  CLKBUFX3 U6941 ( .A(n6344), .Y(n6187) );
  CLKBUFX3 U6942 ( .A(n6344), .Y(n6188) );
  CLKBUFX3 U6943 ( .A(n6343), .Y(n6189) );
  CLKBUFX3 U6944 ( .A(n6343), .Y(n6190) );
  CLKBUFX3 U6945 ( .A(n6343), .Y(n6191) );
  CLKBUFX3 U6946 ( .A(n6343), .Y(n6192) );
  CLKBUFX3 U6947 ( .A(n6343), .Y(n6193) );
  CLKBUFX3 U6948 ( .A(n6343), .Y(n6194) );
  CLKBUFX3 U6949 ( .A(n6343), .Y(n6195) );
  CLKBUFX3 U6950 ( .A(n6343), .Y(n6196) );
  CLKBUFX3 U6951 ( .A(n6343), .Y(n6197) );
  CLKBUFX3 U6952 ( .A(n6343), .Y(n6198) );
  CLKBUFX3 U6953 ( .A(n6343), .Y(n6199) );
  CLKBUFX3 U6954 ( .A(n6343), .Y(n6200) );
  CLKBUFX3 U6955 ( .A(n6342), .Y(n6201) );
  CLKBUFX3 U6956 ( .A(n6342), .Y(n6202) );
  CLKBUFX3 U6957 ( .A(n6342), .Y(n6203) );
  CLKBUFX3 U6958 ( .A(n6342), .Y(n6204) );
  CLKBUFX3 U6959 ( .A(n6342), .Y(n6205) );
  CLKBUFX3 U6960 ( .A(n6342), .Y(n6206) );
  CLKBUFX3 U6961 ( .A(n6342), .Y(n6207) );
  CLKBUFX3 U6962 ( .A(n6342), .Y(n6208) );
  CLKBUFX3 U6963 ( .A(n6342), .Y(n6209) );
  CLKBUFX3 U6964 ( .A(n6342), .Y(n6210) );
  CLKBUFX3 U6965 ( .A(n6342), .Y(n6211) );
  CLKBUFX3 U6966 ( .A(n6342), .Y(n6212) );
  CLKBUFX3 U6967 ( .A(n6341), .Y(n6213) );
  CLKBUFX3 U6968 ( .A(n6341), .Y(n6214) );
  CLKBUFX3 U6969 ( .A(n6341), .Y(n6215) );
  CLKBUFX3 U6970 ( .A(n6341), .Y(n6216) );
  CLKBUFX3 U6971 ( .A(n6341), .Y(n6217) );
  CLKBUFX3 U6972 ( .A(n6341), .Y(n6218) );
  CLKBUFX3 U6973 ( .A(n6341), .Y(n6219) );
  CLKBUFX3 U6974 ( .A(n6341), .Y(n6220) );
  CLKBUFX3 U6975 ( .A(n6341), .Y(n6221) );
  CLKBUFX3 U6976 ( .A(n6341), .Y(n6222) );
  CLKBUFX3 U6977 ( .A(n6341), .Y(n6223) );
  CLKBUFX3 U6978 ( .A(n6334), .Y(n6311) );
  CLKBUFX3 U6979 ( .A(n6334), .Y(n6312) );
  CLKBUFX3 U6980 ( .A(n6334), .Y(n6313) );
  CLKBUFX3 U6981 ( .A(n6334), .Y(n6314) );
  CLKBUFX3 U6982 ( .A(n6334), .Y(n6315) );
  CLKBUFX3 U6983 ( .A(n6334), .Y(n6316) );
  CLKBUFX3 U6984 ( .A(n6334), .Y(n6317) );
  CLKBUFX3 U6985 ( .A(n6334), .Y(n6318) );
  CLKBUFX3 U6986 ( .A(n6334), .Y(n6319) );
  CLKBUFX3 U6987 ( .A(n6334), .Y(n6320) );
  CLKBUFX3 U6988 ( .A(n6333), .Y(n6321) );
  CLKBUFX3 U6989 ( .A(n6333), .Y(n6325) );
  CLKBUFX3 U6990 ( .A(n6333), .Y(n6326) );
  CLKBUFX3 U6991 ( .A(n6333), .Y(n6327) );
  CLKBUFX3 U6992 ( .A(n6333), .Y(n6328) );
  CLKBUFX3 U6993 ( .A(n6333), .Y(n6329) );
  CLKBUFX3 U6994 ( .A(n6333), .Y(n6330) );
  CLKBUFX3 U6995 ( .A(n6333), .Y(n6331) );
  CLKBUFX3 U6996 ( .A(n6333), .Y(n6322) );
  CLKBUFX3 U6997 ( .A(n6333), .Y(n6324) );
  CLKBUFX3 U6998 ( .A(n6333), .Y(n6323) );
  CLKBUFX3 U6999 ( .A(n6333), .Y(n6332) );
  OA22X1 U7000 ( .A0(n10423), .A1(n3877), .B0(n10426), .B1(n4495), .Y(n6751)
         );
  INVX12 U7001 ( .A(n4935), .Y(mem_wdata_D[14]) );
  OR2XL U7002 ( .A(n5040), .B(n10104), .Y(n4935) );
  INVX12 U7003 ( .A(n4943), .Y(mem_wdata_D[15]) );
  OR2XL U7004 ( .A(n5040), .B(n10450), .Y(n4943) );
  INVX12 U7005 ( .A(n4974), .Y(mem_wdata_D[24]) );
  OR2XL U7006 ( .A(n5040), .B(n10423), .Y(n4974) );
  INVX12 U7007 ( .A(n4976), .Y(mem_wdata_D[25]) );
  OR2XL U7008 ( .A(n5040), .B(n10437), .Y(n4976) );
  INVX12 U7009 ( .A(n4978), .Y(mem_wdata_D[26]) );
  OR2XL U7010 ( .A(n5040), .B(n10204), .Y(n4978) );
  INVX12 U7011 ( .A(n4979), .Y(mem_wdata_D[27]) );
  OR2XL U7012 ( .A(n5040), .B(n10397), .Y(n4979) );
  INVX12 U7013 ( .A(n4984), .Y(mem_wdata_D[29]) );
  OR2XL U7014 ( .A(n5040), .B(n10561), .Y(n4984) );
  INVX12 U7015 ( .A(n4985), .Y(mem_wdata_D[30]) );
  OR2XL U7016 ( .A(n5040), .B(n10598), .Y(n4985) );
  INVX12 U7017 ( .A(n4986), .Y(mem_wdata_D[31]) );
  OR2XL U7018 ( .A(n5040), .B(n10705), .Y(n4986) );
  INVX12 U7019 ( .A(n4988), .Y(mem_wdata_D[32]) );
  OR2XL U7020 ( .A(n5040), .B(n10747), .Y(n4988) );
  INVX12 U7021 ( .A(n4989), .Y(mem_wdata_D[33]) );
  OR2XL U7022 ( .A(n5040), .B(n10670), .Y(n4989) );
  INVX12 U7023 ( .A(n4990), .Y(mem_wdata_D[34]) );
  OR2XL U7024 ( .A(n5040), .B(n10195), .Y(n4990) );
  INVX12 U7025 ( .A(n4991), .Y(mem_wdata_D[35]) );
  OR2XL U7026 ( .A(n5040), .B(n10765), .Y(n4991) );
  INVX12 U7027 ( .A(n4992), .Y(mem_wdata_D[36]) );
  OR2XL U7028 ( .A(n5040), .B(n10755), .Y(n4992) );
  INVX12 U7029 ( .A(n4993), .Y(mem_wdata_D[37]) );
  OR2XL U7030 ( .A(n5040), .B(n10900), .Y(n4993) );
  INVX12 U7031 ( .A(n4994), .Y(mem_wdata_D[38]) );
  INVX12 U7032 ( .A(n4995), .Y(mem_wdata_D[39]) );
  OR2XL U7033 ( .A(n5040), .B(n10683), .Y(n4995) );
  INVX12 U7034 ( .A(n4997), .Y(mem_wdata_D[40]) );
  OR2XL U7035 ( .A(n5040), .B(n10656), .Y(n4997) );
  INVX12 U7036 ( .A(n4998), .Y(mem_wdata_D[41]) );
  OR2XL U7037 ( .A(n5040), .B(n10615), .Y(n4998) );
  INVX12 U7038 ( .A(n4999), .Y(mem_wdata_D[42]) );
  OR2XL U7039 ( .A(n5040), .B(n10780), .Y(n4999) );
  INVX12 U7040 ( .A(n5000), .Y(mem_wdata_D[43]) );
  OR2XL U7041 ( .A(n5040), .B(n10793), .Y(n5000) );
  INVX12 U7042 ( .A(n5001), .Y(mem_wdata_D[44]) );
  OR2XL U7043 ( .A(n5040), .B(n10465), .Y(n5001) );
  INVX12 U7044 ( .A(n5002), .Y(mem_wdata_D[45]) );
  OR2XL U7045 ( .A(n5040), .B(n10808), .Y(n5002) );
  INVX12 U7046 ( .A(n5003), .Y(mem_wdata_D[46]) );
  OR2XL U7047 ( .A(n5040), .B(n10107), .Y(n5003) );
  INVX12 U7048 ( .A(n5004), .Y(mem_wdata_D[47]) );
  OR2XL U7049 ( .A(n5040), .B(n10453), .Y(n5004) );
  INVX12 U7050 ( .A(n4922), .Y(mem_wdata_D[70]) );
  OR2XL U7051 ( .A(n5040), .B(n9947), .Y(n4922) );
  INVX12 U7052 ( .A(n4936), .Y(mem_wdata_D[79]) );
  OR2XL U7053 ( .A(n5040), .B(n10447), .Y(n4936) );
  INVX12 U7054 ( .A(n4944), .Y(mem_wdata_D[82]) );
  OR2XL U7055 ( .A(n5040), .B(n10637), .Y(n4944) );
  INVX12 U7056 ( .A(n4933), .Y(mem_wdata_D[86]) );
  OR2XL U7057 ( .A(n5040), .B(n10310), .Y(n4933) );
  INVX12 U7058 ( .A(n4939), .Y(mem_wdata_D[89]) );
  OR2XL U7059 ( .A(n5040), .B(n10434), .Y(n4939) );
  INVX12 U7060 ( .A(n4973), .Y(mem_wdata_D[100]) );
  OR2XL U7061 ( .A(n5040), .B(n9804), .Y(n4973) );
  INVX12 U7062 ( .A(n4975), .Y(mem_wdata_D[103]) );
  OR2XL U7063 ( .A(n5040), .B(n10674), .Y(n4975) );
  INVX12 U7064 ( .A(n4938), .Y(mem_wdata_D[105]) );
  OR2XL U7065 ( .A(n5040), .B(n10606), .Y(n4938) );
  INVX12 U7066 ( .A(n4981), .Y(mem_wdata_D[106]) );
  OR2XL U7067 ( .A(n5040), .B(n10771), .Y(n4981) );
  INVX12 U7068 ( .A(n4971), .Y(mem_wdata_D[120]) );
  OR2XL U7069 ( .A(n5040), .B(n10417), .Y(n4971) );
  INVX12 U7070 ( .A(n4980), .Y(mem_wdata_D[125]) );
  OR2XL U7071 ( .A(n5040), .B(n10555), .Y(n4980) );
  CLKINVX1 U7072 ( .A(n8856), .Y(n8857) );
  CLKBUFX3 U7073 ( .A(n10974), .Y(n5543) );
  CLKINVX1 U7074 ( .A(n9433), .Y(n9436) );
  CLKBUFX3 U7075 ( .A(n5660), .Y(n5626) );
  CLKBUFX3 U7076 ( .A(n5749), .Y(n5719) );
  CLKBUFX3 U7077 ( .A(n5749), .Y(n5718) );
  CLKBUFX3 U7078 ( .A(n5749), .Y(n5717) );
  CLKBUFX3 U7079 ( .A(n5660), .Y(n5629) );
  CLKBUFX3 U7080 ( .A(n5660), .Y(n5628) );
  CLKBUFX3 U7081 ( .A(n5660), .Y(n5627) );
  CLKBUFX3 U7082 ( .A(n5839), .Y(n5808) );
  CLKBUFX3 U7083 ( .A(n5841), .Y(n5807) );
  CLKBUFX3 U7084 ( .A(n5748), .Y(n5720) );
  CLKBUFX3 U7085 ( .A(n5838), .Y(n5809) );
  CLKBUFX3 U7086 ( .A(n5658), .Y(n5630) );
  CLKBUFX3 U7087 ( .A(n5795), .Y(n5763) );
  CLKBUFX3 U7088 ( .A(n5878), .Y(n5853) );
  CLKBUFX3 U7089 ( .A(n5876), .Y(n5852) );
  CLKBUFX3 U7090 ( .A(n5615), .Y(n5585) );
  CLKBUFX3 U7091 ( .A(n5615), .Y(n5584) );
  CLKBUFX3 U7092 ( .A(n5795), .Y(n5762) );
  CLKBUFX3 U7093 ( .A(n5795), .Y(n5761) );
  CLKBUFX3 U7094 ( .A(n5796), .Y(n5760) );
  CLKBUFX3 U7095 ( .A(n5612), .Y(n5586) );
  CLKBUFX3 U7096 ( .A(n5867), .Y(n5854) );
  CLKBUFX3 U7097 ( .A(n5794), .Y(n5764) );
  CLKBUFX3 U7098 ( .A(n5745), .Y(n5732) );
  CLKBUFX3 U7099 ( .A(n5835), .Y(n5821) );
  CLKBUFX3 U7100 ( .A(n5658), .Y(n5642) );
  CLKBUFX3 U7101 ( .A(n5744), .Y(n5733) );
  CLKBUFX3 U7102 ( .A(n5834), .Y(n5822) );
  CLKBUFX3 U7103 ( .A(n5657), .Y(n5643) );
  CLKBUFX3 U7104 ( .A(n5746), .Y(n5727) );
  CLKBUFX3 U7105 ( .A(n5836), .Y(n5816) );
  CLKBUFX3 U7106 ( .A(n5659), .Y(n5637) );
  CLKBUFX3 U7107 ( .A(n5744), .Y(n5734) );
  CLKBUFX3 U7108 ( .A(n5834), .Y(n5823) );
  CLKBUFX3 U7109 ( .A(n5657), .Y(n5644) );
  CLKBUFX3 U7110 ( .A(n5743), .Y(n5737) );
  CLKBUFX3 U7111 ( .A(n5833), .Y(n5826) );
  CLKBUFX3 U7112 ( .A(n5656), .Y(n5647) );
  CLKBUFX3 U7113 ( .A(n5744), .Y(n5736) );
  CLKBUFX3 U7114 ( .A(n5834), .Y(n5825) );
  CLKBUFX3 U7115 ( .A(n5657), .Y(n5646) );
  CLKBUFX3 U7116 ( .A(n5744), .Y(n5735) );
  CLKBUFX3 U7117 ( .A(n5834), .Y(n5824) );
  CLKBUFX3 U7118 ( .A(n5657), .Y(n5645) );
  CLKBUFX3 U7119 ( .A(n5746), .Y(n5728) );
  CLKBUFX3 U7120 ( .A(n5836), .Y(n5817) );
  CLKBUFX3 U7121 ( .A(n5659), .Y(n5638) );
  CLKBUFX3 U7122 ( .A(n5745), .Y(n5729) );
  CLKBUFX3 U7123 ( .A(n5835), .Y(n5818) );
  CLKBUFX3 U7124 ( .A(n5658), .Y(n5639) );
  CLKBUFX3 U7125 ( .A(n5745), .Y(n5730) );
  CLKBUFX3 U7126 ( .A(n5835), .Y(n5819) );
  CLKBUFX3 U7127 ( .A(n5658), .Y(n5640) );
  CLKBUFX3 U7128 ( .A(n5745), .Y(n5731) );
  CLKBUFX3 U7129 ( .A(n5835), .Y(n5820) );
  CLKBUFX3 U7130 ( .A(n5658), .Y(n5641) );
  CLKBUFX3 U7131 ( .A(n5746), .Y(n5726) );
  CLKBUFX3 U7132 ( .A(n5836), .Y(n5815) );
  CLKBUFX3 U7133 ( .A(n5659), .Y(n5636) );
  CLKBUFX3 U7134 ( .A(n5743), .Y(n5738) );
  CLKBUFX3 U7135 ( .A(n5833), .Y(n5827) );
  CLKBUFX3 U7136 ( .A(n5656), .Y(n5648) );
  CLKBUFX3 U7137 ( .A(n5743), .Y(n5740) );
  CLKBUFX3 U7138 ( .A(n5833), .Y(n5829) );
  CLKBUFX3 U7139 ( .A(n5656), .Y(n5650) );
  CLKBUFX3 U7140 ( .A(n5743), .Y(n5739) );
  CLKBUFX3 U7141 ( .A(n5833), .Y(n5828) );
  CLKBUFX3 U7142 ( .A(n5656), .Y(n5649) );
  CLKBUFX3 U7143 ( .A(n5747), .Y(n5721) );
  CLKBUFX3 U7144 ( .A(n5837), .Y(n5810) );
  CLKBUFX3 U7145 ( .A(n5659), .Y(n5631) );
  CLKBUFX3 U7146 ( .A(n5746), .Y(n5725) );
  CLKBUFX3 U7147 ( .A(n5836), .Y(n5814) );
  CLKBUFX3 U7148 ( .A(n5659), .Y(n5635) );
  CLKBUFX3 U7149 ( .A(n5747), .Y(n5724) );
  CLKBUFX3 U7150 ( .A(n5837), .Y(n5813) );
  CLKBUFX3 U7151 ( .A(n5658), .Y(n5634) );
  CLKBUFX3 U7152 ( .A(n5747), .Y(n5723) );
  CLKBUFX3 U7153 ( .A(n5837), .Y(n5812) );
  CLKBUFX3 U7154 ( .A(n5659), .Y(n5633) );
  CLKBUFX3 U7155 ( .A(n5747), .Y(n5722) );
  CLKBUFX3 U7156 ( .A(n5837), .Y(n5811) );
  CLKBUFX3 U7157 ( .A(n5658), .Y(n5632) );
  CLKBUFX3 U7158 ( .A(n5881), .Y(n5866) );
  CLKBUFX3 U7159 ( .A(n5791), .Y(n5776) );
  CLKBUFX3 U7160 ( .A(n5612), .Y(n5598) );
  CLKBUFX3 U7161 ( .A(n5880), .Y(n5867) );
  CLKBUFX3 U7162 ( .A(n5790), .Y(n5777) );
  CLKBUFX3 U7163 ( .A(n5611), .Y(n5599) );
  CLKBUFX3 U7164 ( .A(n5882), .Y(n5861) );
  CLKBUFX3 U7165 ( .A(n5792), .Y(n5771) );
  CLKBUFX3 U7166 ( .A(n5613), .Y(n5593) );
  CLKBUFX3 U7167 ( .A(n5880), .Y(n5868) );
  CLKBUFX3 U7168 ( .A(n5790), .Y(n5778) );
  CLKBUFX3 U7169 ( .A(n5611), .Y(n5600) );
  CLKBUFX3 U7170 ( .A(n5879), .Y(n5871) );
  CLKBUFX3 U7171 ( .A(n5789), .Y(n5781) );
  CLKBUFX3 U7172 ( .A(n5610), .Y(n5603) );
  CLKBUFX3 U7173 ( .A(n5880), .Y(n5870) );
  CLKBUFX3 U7174 ( .A(n5790), .Y(n5780) );
  CLKBUFX3 U7175 ( .A(n5611), .Y(n5602) );
  CLKBUFX3 U7176 ( .A(n5880), .Y(n5869) );
  CLKBUFX3 U7177 ( .A(n5790), .Y(n5779) );
  CLKBUFX3 U7178 ( .A(n5611), .Y(n5601) );
  CLKBUFX3 U7179 ( .A(n5882), .Y(n5862) );
  CLKBUFX3 U7180 ( .A(n5792), .Y(n5772) );
  CLKBUFX3 U7181 ( .A(n5613), .Y(n5594) );
  CLKBUFX3 U7182 ( .A(n5881), .Y(n5863) );
  CLKBUFX3 U7183 ( .A(n5791), .Y(n5773) );
  CLKBUFX3 U7184 ( .A(n5612), .Y(n5595) );
  CLKBUFX3 U7185 ( .A(n5881), .Y(n5864) );
  CLKBUFX3 U7186 ( .A(n5791), .Y(n5774) );
  CLKBUFX3 U7187 ( .A(n5612), .Y(n5596) );
  CLKBUFX3 U7188 ( .A(n5881), .Y(n5865) );
  CLKBUFX3 U7189 ( .A(n5791), .Y(n5775) );
  CLKBUFX3 U7190 ( .A(n5612), .Y(n5597) );
  CLKBUFX3 U7191 ( .A(n5882), .Y(n5860) );
  CLKBUFX3 U7192 ( .A(n5792), .Y(n5770) );
  CLKBUFX3 U7193 ( .A(n5613), .Y(n5592) );
  CLKBUFX3 U7194 ( .A(n5879), .Y(n5872) );
  CLKBUFX3 U7195 ( .A(n5789), .Y(n5782) );
  CLKBUFX3 U7196 ( .A(n5610), .Y(n5604) );
  CLKBUFX3 U7197 ( .A(n5879), .Y(n5874) );
  CLKBUFX3 U7198 ( .A(n5789), .Y(n5784) );
  CLKBUFX3 U7199 ( .A(n5610), .Y(n5606) );
  CLKBUFX3 U7200 ( .A(n5879), .Y(n5873) );
  CLKBUFX3 U7201 ( .A(n5789), .Y(n5783) );
  CLKBUFX3 U7202 ( .A(n5610), .Y(n5605) );
  CLKBUFX3 U7203 ( .A(n5883), .Y(n5855) );
  CLKBUFX3 U7204 ( .A(n5793), .Y(n5765) );
  CLKBUFX3 U7205 ( .A(n5614), .Y(n5587) );
  CLKBUFX3 U7206 ( .A(n5882), .Y(n5859) );
  CLKBUFX3 U7207 ( .A(n5792), .Y(n5769) );
  CLKBUFX3 U7208 ( .A(n5613), .Y(n5591) );
  CLKBUFX3 U7209 ( .A(n5883), .Y(n5858) );
  CLKBUFX3 U7210 ( .A(n5793), .Y(n5768) );
  CLKBUFX3 U7211 ( .A(n5614), .Y(n5590) );
  CLKBUFX3 U7212 ( .A(n5883), .Y(n5857) );
  CLKBUFX3 U7213 ( .A(n5793), .Y(n5767) );
  CLKBUFX3 U7214 ( .A(n5614), .Y(n5589) );
  CLKBUFX3 U7215 ( .A(n5883), .Y(n5856) );
  CLKBUFX3 U7216 ( .A(n5793), .Y(n5766) );
  CLKBUFX3 U7217 ( .A(n5614), .Y(n5588) );
  CLKMX2X2 U7218 ( .A(net107656), .B(net107657), .S0(n149), .Y(n7235) );
  CLKMX2X2 U7219 ( .A(net107656), .B(net107657), .S0(n3764), .Y(n7782) );
  CLKMX2X2 U7220 ( .A(net107656), .B(net107657), .S0(n8119), .Y(n7315) );
  CLKMX2X2 U7221 ( .A(net107656), .B(net107657), .S0(n9138), .Y(n9139) );
  CLKINVX1 U7222 ( .A(n8887), .Y(n8883) );
  INVX3 U7223 ( .A(n5462), .Y(n5461) );
  INVX3 U7224 ( .A(n1937), .Y(n5471) );
  INVX3 U7225 ( .A(n1937), .Y(n5472) );
  INVX3 U7226 ( .A(n1986), .Y(n5195) );
  INVX3 U7227 ( .A(n1986), .Y(n5196) );
  INVX3 U7228 ( .A(n2896), .Y(n5478) );
  INVX3 U7229 ( .A(n2896), .Y(n5479) );
  INVX3 U7230 ( .A(n1933), .Y(n5518) );
  INVX3 U7231 ( .A(n338), .Y(n5492) );
  INVX3 U7232 ( .A(n5475), .Y(n5473) );
  INVX3 U7233 ( .A(n5510), .Y(n5508) );
  INVX3 U7234 ( .A(n5507), .Y(n5505) );
  CLKBUFX3 U7235 ( .A(n339), .Y(n5507) );
  INVX3 U7236 ( .A(n152), .Y(n5526) );
  INVX3 U7237 ( .A(n5496), .Y(n5494) );
  INVX3 U7238 ( .A(n5504), .Y(n5502) );
  CLKBUFX3 U7239 ( .A(n1936), .Y(n5504) );
  INVX3 U7240 ( .A(n154), .Y(n5511) );
  INVX3 U7241 ( .A(n5457), .Y(n5455) );
  INVX3 U7242 ( .A(n157), .Y(n5226) );
  INVX3 U7243 ( .A(n5465), .Y(n5463) );
  CLKBUFX3 U7244 ( .A(n1934), .Y(n5465) );
  INVX3 U7245 ( .A(n1933), .Y(n5519) );
  INVX3 U7246 ( .A(n338), .Y(n5493) );
  INVX3 U7247 ( .A(n5475), .Y(n5474) );
  INVX3 U7248 ( .A(n5510), .Y(n5509) );
  INVX3 U7249 ( .A(n5507), .Y(n5506) );
  INVX3 U7250 ( .A(n152), .Y(n5527) );
  INVX3 U7251 ( .A(n5496), .Y(n5495) );
  INVX3 U7252 ( .A(n5504), .Y(n5503) );
  INVX3 U7253 ( .A(n154), .Y(n5512) );
  INVX3 U7254 ( .A(n5457), .Y(n5456) );
  INVX3 U7255 ( .A(n157), .Y(n5227) );
  INVX3 U7256 ( .A(n5465), .Y(n5464) );
  INVX3 U7257 ( .A(n341), .Y(n5458) );
  INVX3 U7258 ( .A(n341), .Y(n5459) );
  INVX3 U7259 ( .A(net134682), .Y(net118381) );
  CLKBUFX3 U7260 ( .A(net107619), .Y(net118281) );
  CLKBUFX2 U7261 ( .A(n3633), .Y(net115813) );
  CLKBUFX3 U7262 ( .A(n5929), .Y(n5924) );
  CLKBUFX3 U7263 ( .A(n5706), .Y(n5699) );
  CLKBUFX3 U7264 ( .A(n5929), .Y(n5925) );
  CLKBUFX3 U7265 ( .A(n5706), .Y(n5700) );
  CLKBUFX3 U7266 ( .A(n5929), .Y(n5926) );
  CLKBUFX3 U7267 ( .A(n5706), .Y(n5701) );
  CLKBUFX3 U7268 ( .A(n5116), .Y(n5113) );
  CLKBUFX3 U7269 ( .A(n5142), .Y(n5141) );
  CLKBUFX3 U7270 ( .A(n9502), .Y(n5133) );
  CLKBUFX3 U7271 ( .A(n5116), .Y(n5115) );
  CLKBUFX3 U7272 ( .A(n5142), .Y(n5139) );
  NAND2X1 U7273 ( .A(n5532), .B(n5953), .Y(n10797) );
  CLKINVX1 U7274 ( .A(n10469), .Y(n10177) );
  CLKBUFX3 U7275 ( .A(n6345), .Y(n6017) );
  CLKBUFX3 U7276 ( .A(n6358), .Y(n6018) );
  CLKBUFX3 U7277 ( .A(n6358), .Y(n6019) );
  CLKBUFX3 U7278 ( .A(n6333), .Y(n6020) );
  CLKBUFX3 U7279 ( .A(n6357), .Y(n6021) );
  CLKBUFX3 U7280 ( .A(n6357), .Y(n6022) );
  CLKBUFX3 U7281 ( .A(n6357), .Y(n6023) );
  CLKBUFX3 U7282 ( .A(n6357), .Y(n6024) );
  CLKBUFX3 U7283 ( .A(n6357), .Y(n6025) );
  CLKBUFX3 U7284 ( .A(n6357), .Y(n6026) );
  CLKBUFX3 U7285 ( .A(n6357), .Y(n6027) );
  CLKBUFX3 U7286 ( .A(n6357), .Y(n6028) );
  CLKBUFX3 U7287 ( .A(n6357), .Y(n6029) );
  CLKBUFX3 U7288 ( .A(n6357), .Y(n6030) );
  CLKBUFX3 U7289 ( .A(n6357), .Y(n6031) );
  CLKBUFX3 U7290 ( .A(n6357), .Y(n6032) );
  CLKBUFX3 U7291 ( .A(n6356), .Y(n6033) );
  CLKBUFX3 U7292 ( .A(n6356), .Y(n6034) );
  CLKBUFX3 U7293 ( .A(n6356), .Y(n6035) );
  CLKBUFX3 U7294 ( .A(n6356), .Y(n6036) );
  CLKBUFX3 U7295 ( .A(n6356), .Y(n6037) );
  CLKBUFX3 U7296 ( .A(n6356), .Y(n6038) );
  CLKBUFX3 U7297 ( .A(n6356), .Y(n6039) );
  CLKBUFX3 U7298 ( .A(n6356), .Y(n6040) );
  CLKBUFX3 U7299 ( .A(n6356), .Y(n6041) );
  CLKBUFX3 U7300 ( .A(n6356), .Y(n6042) );
  CLKBUFX3 U7301 ( .A(n6356), .Y(n6043) );
  CLKBUFX3 U7302 ( .A(n6356), .Y(n6044) );
  CLKBUFX3 U7303 ( .A(n6358), .Y(n6355) );
  CLKBUFX3 U7304 ( .A(n6358), .Y(n6354) );
  CLKBUFX3 U7305 ( .A(n6358), .Y(n6353) );
  CLKBUFX3 U7306 ( .A(rst_n), .Y(n6352) );
  CLKBUFX3 U7307 ( .A(n6346), .Y(n6351) );
  CLKBUFX3 U7308 ( .A(rst_n), .Y(n6350) );
  CLKBUFX3 U7309 ( .A(n6338), .Y(n6340) );
  CLKBUFX3 U7310 ( .A(n6358), .Y(n6339) );
  CLKBUFX3 U7311 ( .A(n6358), .Y(n6338) );
  CLKBUFX3 U7312 ( .A(n6342), .Y(n6337) );
  CLKBUFX3 U7313 ( .A(n6332), .Y(n6336) );
  CLKBUFX3 U7314 ( .A(n6358), .Y(n6335) );
  CLKBUFX3 U7315 ( .A(n6358), .Y(n6349) );
  CLKBUFX3 U7316 ( .A(n6358), .Y(n6348) );
  CLKBUFX3 U7317 ( .A(n6358), .Y(n6347) );
  CLKBUFX3 U7318 ( .A(rst_n), .Y(n6346) );
  CLKBUFX3 U7319 ( .A(rst_n), .Y(n6345) );
  CLKBUFX3 U7320 ( .A(n6358), .Y(n6344) );
  CLKBUFX3 U7321 ( .A(n6350), .Y(n6343) );
  CLKBUFX3 U7322 ( .A(n6358), .Y(n6342) );
  CLKBUFX3 U7323 ( .A(n6335), .Y(n6341) );
  CLKBUFX3 U7324 ( .A(rst_n), .Y(n6334) );
  CLKBUFX3 U7325 ( .A(n6352), .Y(n6333) );
  INVX12 U7326 ( .A(n1861), .Y(mem_wdata_D[6]) );
  INVX12 U7327 ( .A(n1862), .Y(mem_wdata_D[7]) );
  INVX12 U7328 ( .A(n1863), .Y(mem_wdata_D[8]) );
  INVX12 U7329 ( .A(n1864), .Y(mem_wdata_D[9]) );
  INVX12 U7330 ( .A(n1865), .Y(mem_wdata_D[10]) );
  INVX12 U7331 ( .A(n1866), .Y(mem_wdata_D[12]) );
  INVX12 U7332 ( .A(n1867), .Y(mem_wdata_D[13]) );
  INVX12 U7333 ( .A(n1868), .Y(mem_wdata_D[16]) );
  INVX12 U7334 ( .A(n1869), .Y(mem_wdata_D[17]) );
  INVX12 U7335 ( .A(n1870), .Y(mem_wdata_D[18]) );
  INVX12 U7336 ( .A(n1871), .Y(mem_wdata_D[19]) );
  INVX12 U7337 ( .A(n1872), .Y(mem_wdata_D[20]) );
  INVX12 U7338 ( .A(n1873), .Y(mem_wdata_D[21]) );
  INVX12 U7339 ( .A(n1874), .Y(mem_wdata_D[22]) );
  INVX12 U7340 ( .A(n1875), .Y(mem_wdata_D[23]) );
  INVX12 U7341 ( .A(n1876), .Y(mem_wdata_D[28]) );
  CLKINVX1 U7342 ( .A(n8673), .Y(n8674) );
  AO21X1 U7343 ( .A0(n8673), .A1(n7025), .B0(n8643), .Y(n7058) );
  NAND2XL U7344 ( .A(net117747), .B(n7047), .Y(n7060) );
  CLKINVX1 U7345 ( .A(n7593), .Y(n7596) );
  INVX12 U7346 ( .A(n1857), .Y(mem_wdata_D[2]) );
  INVX12 U7347 ( .A(n1858), .Y(mem_wdata_D[3]) );
  INVX12 U7348 ( .A(n1859), .Y(mem_wdata_D[4]) );
  INVX12 U7349 ( .A(n1860), .Y(mem_wdata_D[5]) );
  INVX12 U7350 ( .A(n1877), .Y(mem_wdata_D[53]) );
  INVX12 U7351 ( .A(n1878), .Y(mem_wdata_D[56]) );
  INVX12 U7352 ( .A(n1879), .Y(mem_wdata_D[58]) );
  INVX12 U7353 ( .A(n1880), .Y(mem_wdata_D[59]) );
  INVX12 U7354 ( .A(n1881), .Y(mem_wdata_D[61]) );
  INVX12 U7355 ( .A(n1883), .Y(mem_wdata_D[64]) );
  INVX12 U7356 ( .A(n1885), .Y(mem_wdata_D[69]) );
  INVX12 U7357 ( .A(n1887), .Y(mem_wdata_D[72]) );
  INVX12 U7358 ( .A(n1890), .Y(mem_wdata_D[75]) );
  INVX12 U7359 ( .A(n1893), .Y(mem_wdata_D[78]) );
  CLKINVX1 U7360 ( .A(n7847), .Y(n7851) );
  CLKINVX1 U7361 ( .A(n7861), .Y(n7848) );
  NOR4X1 U7362 ( .A(n8889), .B(n8644), .C(n8680), .D(n8643), .Y(n8676) );
  CLKINVX1 U7363 ( .A(n9050), .Y(n8215) );
  CLKINVX1 U7364 ( .A(n9604), .Y(n9605) );
  INVXL U7365 ( .A(n8381), .Y(n8377) );
  INVX12 U7366 ( .A(n1882), .Y(mem_wdata_D[62]) );
  INVX12 U7367 ( .A(n1884), .Y(mem_wdata_D[65]) );
  INVX12 U7368 ( .A(n4893), .Y(mem_wdata_D[67]) );
  INVX1 U7369 ( .A(n12853), .Y(n4893) );
  INVX12 U7370 ( .A(n4902), .Y(mem_wdata_D[68]) );
  INVX1 U7371 ( .A(n12852), .Y(n4902) );
  INVX12 U7372 ( .A(n1886), .Y(mem_wdata_D[71]) );
  INVX12 U7373 ( .A(n1888), .Y(mem_wdata_D[73]) );
  INVX12 U7374 ( .A(n1889), .Y(mem_wdata_D[74]) );
  INVX12 U7375 ( .A(n1891), .Y(mem_wdata_D[76]) );
  INVX12 U7376 ( .A(n1892), .Y(mem_wdata_D[77]) );
  INVX12 U7377 ( .A(n1894), .Y(mem_wdata_D[80]) );
  INVX12 U7378 ( .A(n1895), .Y(mem_wdata_D[81]) );
  INVX12 U7379 ( .A(n1896), .Y(mem_wdata_D[83]) );
  INVX12 U7380 ( .A(n1897), .Y(mem_wdata_D[84]) );
  INVX12 U7381 ( .A(n1898), .Y(mem_wdata_D[85]) );
  INVX12 U7382 ( .A(n1899), .Y(mem_wdata_D[87]) );
  INVX12 U7383 ( .A(n1900), .Y(mem_wdata_D[88]) );
  INVX12 U7384 ( .A(n4907), .Y(mem_wdata_D[90]) );
  INVX1 U7385 ( .A(n12851), .Y(n4907) );
  INVX12 U7386 ( .A(n1901), .Y(mem_wdata_D[91]) );
  INVX12 U7387 ( .A(n1902), .Y(mem_wdata_D[92]) );
  INVX12 U7388 ( .A(n1903), .Y(mem_wdata_D[93]) );
  INVX12 U7389 ( .A(n1904), .Y(mem_wdata_D[94]) );
  INVX12 U7390 ( .A(n1905), .Y(mem_wdata_D[95]) );
  INVX12 U7391 ( .A(n1906), .Y(mem_wdata_D[96]) );
  INVX12 U7392 ( .A(n1907), .Y(mem_wdata_D[97]) );
  INVX12 U7393 ( .A(n1908), .Y(mem_wdata_D[98]) );
  INVX12 U7394 ( .A(n1909), .Y(mem_wdata_D[99]) );
  INVX12 U7395 ( .A(n1910), .Y(mem_wdata_D[101]) );
  INVX12 U7396 ( .A(n1911), .Y(mem_wdata_D[104]) );
  INVX12 U7397 ( .A(n1912), .Y(mem_wdata_D[107]) );
  INVX12 U7398 ( .A(n1913), .Y(mem_wdata_D[108]) );
  INVX12 U7399 ( .A(n1914), .Y(mem_wdata_D[109]) );
  INVX12 U7400 ( .A(n1915), .Y(mem_wdata_D[110]) );
  INVX12 U7401 ( .A(n1916), .Y(mem_wdata_D[111]) );
  INVX12 U7402 ( .A(n1917), .Y(mem_wdata_D[112]) );
  INVX12 U7403 ( .A(n1918), .Y(mem_wdata_D[113]) );
  INVX12 U7404 ( .A(n1919), .Y(mem_wdata_D[114]) );
  INVX12 U7405 ( .A(n1920), .Y(mem_wdata_D[115]) );
  INVX12 U7406 ( .A(n1921), .Y(mem_wdata_D[116]) );
  INVX12 U7407 ( .A(n4954), .Y(mem_wdata_D[117]) );
  INVX1 U7408 ( .A(n12850), .Y(n4954) );
  INVX12 U7409 ( .A(n1922), .Y(mem_wdata_D[119]) );
  INVX12 U7410 ( .A(n1923), .Y(mem_wdata_D[121]) );
  INVX12 U7411 ( .A(n1924), .Y(mem_wdata_D[122]) );
  INVX12 U7412 ( .A(n1925), .Y(mem_wdata_D[124]) );
  INVX12 U7413 ( .A(n1926), .Y(mem_wdata_D[126]) );
  NAND2X1 U7414 ( .A(n11217), .B(n11218), .Y(n11343) );
  CLKINVX1 U7415 ( .A(n8886), .Y(n8864) );
  NAND3BX1 U7416 ( .AN(n4753), .B(n8481), .C(net117745), .Y(n8490) );
  INVXL U7417 ( .A(net107992), .Y(net107991) );
  NAND2XL U7418 ( .A(n3733), .B(net105549), .Y(n10631) );
  NAND2XL U7419 ( .A(net105834), .B(net105835), .Y(n10686) );
  NAND2XL U7420 ( .A(net106040), .B(net106041), .Y(n10868) );
  NAND2XL U7421 ( .A(net105731), .B(net105732), .Y(n10825) );
  NAND2XL U7422 ( .A(n3023), .B(net105430), .Y(n10569) );
  NAND2XL U7423 ( .A(n3015), .B(net105269), .Y(n11055) );
  NAND2X1 U7424 ( .A(n7669), .B(n7591), .Y(n9427) );
  CLKINVX1 U7425 ( .A(n11394), .Y(n10640) );
  CLKINVX1 U7426 ( .A(n11473), .Y(n10661) );
  CLKINVX1 U7427 ( .A(n11493), .Y(n10514) );
  CLKINVX1 U7428 ( .A(n11492), .Y(n10404) );
  CLKINVX1 U7429 ( .A(n11488), .Y(n10499) );
  CLKINVX1 U7430 ( .A(n11385), .Y(n10612) );
  CLKINVX1 U7431 ( .A(n11440), .Y(n10741) );
  CLKINVX1 U7432 ( .A(n11460), .Y(n10407) );
  CLKINVX1 U7433 ( .A(n11456), .Y(n10502) );
  CLKINVX1 U7434 ( .A(n11466), .Y(n10201) );
  CLKINVX1 U7435 ( .A(n11449), .Y(n10609) );
  CLKINVX1 U7436 ( .A(n11447), .Y(n10677) );
  CLKINVX1 U7437 ( .A(n8122), .Y(n7304) );
  CLKINVX1 U7438 ( .A(net109176), .Y(net108852) );
  CLKINVX1 U7439 ( .A(n9308), .Y(n9319) );
  CLKINVX1 U7440 ( .A(n7494), .Y(n8469) );
  CLKINVX1 U7441 ( .A(n7399), .Y(n7407) );
  CLKINVX1 U7442 ( .A(n7400), .Y(n11102) );
  NAND3BXL U7443 ( .AN(n6825), .B(n6838), .C(net135551), .Y(n6821) );
  INVXL U7444 ( .A(n9206), .Y(n6665) );
  OA22X1 U7445 ( .A0(n10687), .A1(n3767), .B0(n10689), .B1(n9536), .Y(n7078)
         );
  OA22X1 U7446 ( .A0(n10561), .A1(n3877), .B0(n10564), .B1(n4495), .Y(n6981)
         );
  AND3XL U7447 ( .A(n6730), .B(n6729), .C(net117747), .Y(n6732) );
  AND2XL U7448 ( .A(net135551), .B(n6826), .Y(n4701) );
  CLKINVX1 U7449 ( .A(n7669), .Y(n7670) );
  AND2X2 U7450 ( .A(n8886), .B(n7861), .Y(n4709) );
  CLKINVX1 U7451 ( .A(n9541), .Y(n9449) );
  CLKINVX1 U7452 ( .A(n11369), .Y(n6369) );
  CLKINVX1 U7453 ( .A(n11365), .Y(n6365) );
  CLKINVX1 U7454 ( .A(n11097), .Y(n11098) );
  NAND2BXL U7455 ( .AN(n9444), .B(n9445), .Y(n9459) );
  NAND2XL U7456 ( .A(n4733), .B(n7595), .Y(n6958) );
  INVXL U7457 ( .A(n8288), .Y(n8289) );
  CLKINVX1 U7458 ( .A(n6919), .Y(n6828) );
  CLKINVX1 U7459 ( .A(n7961), .Y(n7942) );
  CLKINVX1 U7460 ( .A(n8692), .Y(n8693) );
  CLKINVX1 U7461 ( .A(n7034), .Y(n7035) );
  CLKINVX1 U7462 ( .A(n11105), .Y(n11109) );
  CLKBUFX3 U7463 ( .A(net134685), .Y(net118483) );
  CLKBUFX3 U7464 ( .A(net134685), .Y(net118487) );
  CLKBUFX3 U7465 ( .A(net134679), .Y(net118339) );
  CLKBUFX3 U7466 ( .A(net134683), .Y(net118441) );
  CLKBUFX3 U7467 ( .A(net134679), .Y(net118345) );
  CLKBUFX3 U7468 ( .A(net134683), .Y(net118439) );
  CLKBUFX3 U7469 ( .A(net134679), .Y(net118343) );
  CLKBUFX3 U7470 ( .A(net134679), .Y(net118341) );
  CLKBUFX3 U7471 ( .A(net134679), .Y(net118337) );
  CLKBUFX3 U7472 ( .A(net134681), .Y(net118365) );
  AND2X2 U7473 ( .A(n4722), .B(n4721), .Y(n4713) );
  CLKINVX1 U7474 ( .A(n10362), .Y(n10352) );
  CLKINVX1 U7475 ( .A(n10331), .Y(n10321) );
  CLKINVX1 U7476 ( .A(n10632), .Y(n5510) );
  NAND2XL U7477 ( .A(net104962), .B(n3667), .Y(n10632) );
  INVX1 U7478 ( .A(n10527), .Y(n5496) );
  NAND2XL U7479 ( .A(net105119), .B(net105120), .Y(n10527) );
  INVX1 U7480 ( .A(n9938), .Y(n5457) );
  CLKINVX1 U7481 ( .A(n11096), .Y(n11100) );
  CLKINVX1 U7482 ( .A(n8374), .Y(n7586) );
  MX2XL U7483 ( .A(net118592), .B(net118597), .S0(n7041), .Y(n7044) );
  MX2XL U7484 ( .A(net118597), .B(net118592), .S0(n9209), .Y(n9213) );
  MX2XL U7485 ( .A(net118597), .B(net118592), .S0(n7407), .Y(n7415) );
  CLKINVX1 U7486 ( .A(n8697), .Y(n8710) );
  CLKINVX1 U7487 ( .A(n9317), .Y(n8868) );
  CLKINVX1 U7488 ( .A(n6960), .Y(n6940) );
  CLKINVX1 U7489 ( .A(n7482), .Y(n7483) );
  CLKBUFX3 U7490 ( .A(n4759), .Y(n5098) );
  CLKBUFX3 U7491 ( .A(n4760), .Y(n5102) );
  INVX3 U7492 ( .A(n5499), .Y(n5497) );
  INVX3 U7493 ( .A(n5499), .Y(n5498) );
  INVX3 U7494 ( .A(n153), .Y(n5500) );
  INVX3 U7495 ( .A(n156), .Y(n5480) );
  INVX3 U7496 ( .A(n5468), .Y(n5466) );
  CLKBUFX3 U7497 ( .A(n337), .Y(n5468) );
  INVX3 U7498 ( .A(n5491), .Y(n5489) );
  INVX3 U7499 ( .A(n151), .Y(n5482) );
  INVX3 U7500 ( .A(n354), .Y(n5487) );
  INVX3 U7501 ( .A(n5486), .Y(n5484) );
  CLKBUFX3 U7502 ( .A(n340), .Y(n5486) );
  INVX3 U7503 ( .A(n4716), .Y(n5524) );
  INVX3 U7504 ( .A(n153), .Y(n5501) );
  INVX3 U7505 ( .A(n156), .Y(n5481) );
  INVX3 U7506 ( .A(n5468), .Y(n5467) );
  INVX3 U7507 ( .A(n5491), .Y(n5490) );
  INVX3 U7508 ( .A(n151), .Y(n5483) );
  INVX3 U7509 ( .A(n354), .Y(n5488) );
  INVX3 U7510 ( .A(n5486), .Y(n5485) );
  INVX3 U7511 ( .A(n4716), .Y(n5525) );
  INVX3 U7512 ( .A(n166), .Y(n5476) );
  INVX3 U7513 ( .A(n166), .Y(n5477) );
  INVX3 U7514 ( .A(n1935), .Y(n5469) );
  INVX3 U7515 ( .A(n155), .Y(n5516) );
  INVX3 U7516 ( .A(n5515), .Y(n5513) );
  CLKBUFX3 U7517 ( .A(n357), .Y(n5515) );
  INVX3 U7518 ( .A(n342), .Y(n5522) );
  INVX3 U7519 ( .A(n1935), .Y(n5470) );
  INVX3 U7520 ( .A(n155), .Y(n5517) );
  INVX3 U7521 ( .A(n5515), .Y(n5514) );
  INVX3 U7522 ( .A(n342), .Y(n5523) );
  CLKINVX1 U7523 ( .A(n9134), .Y(n8482) );
  CLKBUFX3 U7524 ( .A(n5851), .Y(n5881) );
  CLKBUFX3 U7525 ( .A(n5750), .Y(n5745) );
  CLKBUFX3 U7526 ( .A(n5797), .Y(n5791) );
  CLKBUFX3 U7527 ( .A(n5840), .Y(n5835) );
  CLKBUFX3 U7528 ( .A(n5616), .Y(n5612) );
  CLKBUFX3 U7529 ( .A(n5662), .Y(n5658) );
  CLKBUFX3 U7530 ( .A(n5879), .Y(n5882) );
  CLKBUFX3 U7531 ( .A(n5750), .Y(n5746) );
  CLKBUFX3 U7532 ( .A(n5797), .Y(n5792) );
  CLKBUFX3 U7533 ( .A(n5840), .Y(n5836) );
  CLKBUFX3 U7534 ( .A(n5616), .Y(n5613) );
  CLKBUFX3 U7535 ( .A(n5662), .Y(n5659) );
  CLKBUFX3 U7536 ( .A(n5874), .Y(n5883) );
  CLKBUFX3 U7537 ( .A(n5750), .Y(n5747) );
  CLKBUFX3 U7538 ( .A(n5797), .Y(n5793) );
  CLKBUFX3 U7539 ( .A(n5840), .Y(n5837) );
  CLKBUFX3 U7540 ( .A(n5616), .Y(n5614) );
  CLKBUFX3 U7541 ( .A(n11210), .Y(n5929) );
  CLKBUFX3 U7542 ( .A(net139718), .Y(net117665) );
  CLKBUFX3 U7543 ( .A(net139718), .Y(net117667) );
  CLKBUFX3 U7544 ( .A(n5937), .Y(n5932) );
  CLKBUFX3 U7545 ( .A(net107606), .Y(net118223) );
  CLKBUFX3 U7546 ( .A(net134679), .Y(net118347) );
  NAND2BX1 U7547 ( .AN(n10259), .B(n10175), .Y(n10469) );
  CLKINVX1 U7548 ( .A(n10290), .Y(n10280) );
  CLKBUFX3 U7549 ( .A(\i_MIPS/Register/n147 ), .Y(n6014) );
  CLKBUFX3 U7550 ( .A(\i_MIPS/Register/n147 ), .Y(n6015) );
  CLKBUFX3 U7551 ( .A(\i_MIPS/Register/n146 ), .Y(n6012) );
  CLKBUFX3 U7552 ( .A(\i_MIPS/Register/n146 ), .Y(n6013) );
  CLKBUFX3 U7553 ( .A(\i_MIPS/Register/n145 ), .Y(n6010) );
  CLKBUFX3 U7554 ( .A(\i_MIPS/Register/n145 ), .Y(n6011) );
  CLKBUFX3 U7555 ( .A(\i_MIPS/Register/n144 ), .Y(n6008) );
  CLKBUFX3 U7556 ( .A(\i_MIPS/Register/n144 ), .Y(n6009) );
  CLKBUFX3 U7557 ( .A(\i_MIPS/Register/n143 ), .Y(n6006) );
  CLKBUFX3 U7558 ( .A(\i_MIPS/Register/n143 ), .Y(n6007) );
  CLKBUFX3 U7559 ( .A(\i_MIPS/Register/n142 ), .Y(n6004) );
  CLKBUFX3 U7560 ( .A(\i_MIPS/Register/n142 ), .Y(n6005) );
  CLKBUFX3 U7561 ( .A(\i_MIPS/Register/n141 ), .Y(n6002) );
  CLKBUFX3 U7562 ( .A(\i_MIPS/Register/n141 ), .Y(n6003) );
  CLKBUFX3 U7563 ( .A(\i_MIPS/Register/n139 ), .Y(n6000) );
  CLKBUFX3 U7564 ( .A(\i_MIPS/Register/n139 ), .Y(n6001) );
  CLKBUFX3 U7565 ( .A(\i_MIPS/Register/n138 ), .Y(n5998) );
  CLKBUFX3 U7566 ( .A(\i_MIPS/Register/n138 ), .Y(n5999) );
  CLKBUFX3 U7567 ( .A(\i_MIPS/Register/n137 ), .Y(n5996) );
  CLKBUFX3 U7568 ( .A(\i_MIPS/Register/n137 ), .Y(n5997) );
  CLKBUFX3 U7569 ( .A(\i_MIPS/Register/n136 ), .Y(n5994) );
  CLKBUFX3 U7570 ( .A(\i_MIPS/Register/n136 ), .Y(n5995) );
  CLKBUFX3 U7571 ( .A(\i_MIPS/Register/n135 ), .Y(n5992) );
  CLKBUFX3 U7572 ( .A(\i_MIPS/Register/n135 ), .Y(n5993) );
  CLKBUFX3 U7573 ( .A(\i_MIPS/Register/n134 ), .Y(n5990) );
  CLKBUFX3 U7574 ( .A(\i_MIPS/Register/n134 ), .Y(n5991) );
  CLKBUFX3 U7575 ( .A(\i_MIPS/Register/n133 ), .Y(n5988) );
  CLKBUFX3 U7576 ( .A(\i_MIPS/Register/n133 ), .Y(n5989) );
  CLKBUFX3 U7577 ( .A(\i_MIPS/Register/n132 ), .Y(n5986) );
  CLKBUFX3 U7578 ( .A(\i_MIPS/Register/n132 ), .Y(n5987) );
  CLKBUFX3 U7579 ( .A(\i_MIPS/Register/n130 ), .Y(n5984) );
  CLKBUFX3 U7580 ( .A(\i_MIPS/Register/n130 ), .Y(n5985) );
  CLKBUFX3 U7581 ( .A(\i_MIPS/Register/n129 ), .Y(n5982) );
  CLKBUFX3 U7582 ( .A(\i_MIPS/Register/n129 ), .Y(n5983) );
  CLKBUFX3 U7583 ( .A(\i_MIPS/Register/n128 ), .Y(n5980) );
  CLKBUFX3 U7584 ( .A(\i_MIPS/Register/n128 ), .Y(n5981) );
  CLKBUFX3 U7585 ( .A(\i_MIPS/Register/n127 ), .Y(n5978) );
  CLKBUFX3 U7586 ( .A(\i_MIPS/Register/n127 ), .Y(n5979) );
  CLKBUFX3 U7587 ( .A(\i_MIPS/Register/n126 ), .Y(n5976) );
  CLKBUFX3 U7588 ( .A(\i_MIPS/Register/n126 ), .Y(n5977) );
  CLKBUFX3 U7589 ( .A(\i_MIPS/Register/n125 ), .Y(n5974) );
  CLKBUFX3 U7590 ( .A(\i_MIPS/Register/n125 ), .Y(n5975) );
  CLKBUFX3 U7591 ( .A(\i_MIPS/Register/n124 ), .Y(n5972) );
  CLKBUFX3 U7592 ( .A(\i_MIPS/Register/n124 ), .Y(n5973) );
  CLKBUFX3 U7593 ( .A(\i_MIPS/Register/n123 ), .Y(n5970) );
  CLKBUFX3 U7594 ( .A(\i_MIPS/Register/n123 ), .Y(n5971) );
  CLKBUFX3 U7595 ( .A(\i_MIPS/Register/n121 ), .Y(n5968) );
  CLKBUFX3 U7596 ( .A(\i_MIPS/Register/n121 ), .Y(n5969) );
  CLKBUFX3 U7597 ( .A(\i_MIPS/Register/n112 ), .Y(n5960) );
  CLKBUFX3 U7598 ( .A(\i_MIPS/Register/n112 ), .Y(n5961) );
  CLKBUFX3 U7599 ( .A(\i_MIPS/Register/n108 ), .Y(n5956) );
  CLKBUFX3 U7600 ( .A(\i_MIPS/Register/n108 ), .Y(n5957) );
  CLKBUFX3 U7601 ( .A(\i_MIPS/Register/n106 ), .Y(n5954) );
  CLKBUFX3 U7602 ( .A(\i_MIPS/Register/n106 ), .Y(n5955) );
  CLKBUFX3 U7603 ( .A(\i_MIPS/Register/n116 ), .Y(n5964) );
  CLKBUFX3 U7604 ( .A(\i_MIPS/Register/n116 ), .Y(n5965) );
  CLKBUFX3 U7605 ( .A(\i_MIPS/Register/n114 ), .Y(n5962) );
  CLKBUFX3 U7606 ( .A(\i_MIPS/Register/n114 ), .Y(n5963) );
  CLKBUFX3 U7607 ( .A(\i_MIPS/Register/n110 ), .Y(n5958) );
  CLKBUFX3 U7608 ( .A(\i_MIPS/Register/n110 ), .Y(n5959) );
  CLKBUFX3 U7609 ( .A(\i_MIPS/Register/n118 ), .Y(n5966) );
  CLKBUFX3 U7610 ( .A(\i_MIPS/Register/n118 ), .Y(n5967) );
  CLKBUFX3 U7611 ( .A(n10798), .Y(n5531) );
  CLKINVX1 U7612 ( .A(n10903), .Y(n10908) );
  CLKBUFX3 U7613 ( .A(n6354), .Y(n6357) );
  CLKBUFX3 U7614 ( .A(n6339), .Y(n6356) );
  CLKBUFX3 U7615 ( .A(n6334), .Y(n6358) );
  CLKINVX1 U7616 ( .A(n11589), .Y(n11062) );
  OA22XL U7617 ( .A0(n5258), .A1(n1279), .B0(n5291), .B1(n2911), .Y(n6560) );
  AO22X1 U7618 ( .A0(DCACHE_addr[19]), .A1(n11534), .B0(n5947), .B1(n11523), 
        .Y(n12846) );
  INVX12 U7619 ( .A(n350), .Y(mem_addr_D[4]) );
  NAND4BX1 U7620 ( .AN(n9392), .B(n9391), .C(n9390), .D(n9389), .Y(n9403) );
  NAND4BX1 U7621 ( .AN(n9401), .B(n9400), .C(n9399), .D(n9398), .Y(n9402) );
  CLKMX2X2 U7622 ( .A(n9516), .B(n9515), .S0(net114079), .Y(n9576) );
  NAND4BX1 U7623 ( .AN(n9497), .B(n9496), .C(n9495), .D(n9494), .Y(n9516) );
  NAND4BX1 U7624 ( .AN(n9514), .B(n9513), .C(n9512), .D(n9511), .Y(n9515) );
  CLKMX2X2 U7625 ( .A(n8108), .B(n8107), .S0(net114081), .Y(net109839) );
  CLKMX2X2 U7626 ( .A(n8854), .B(n8853), .S0(net114079), .Y(net108490) );
  CLKMX2X2 U7627 ( .A(n8025), .B(n8024), .S0(net114081), .Y(net109989) );
  CLKMX2X2 U7628 ( .A(n7764), .B(n7763), .S0(net114087), .Y(n7815) );
  NAND4BX1 U7629 ( .AN(n7753), .B(n7752), .C(n7751), .D(n7750), .Y(n7764) );
  CLKMX2X2 U7630 ( .A(n6912), .B(n6911), .S0(\i_MIPS/jump_addr[22] ), .Y(
        net111930) );
  NOR2BX1 U7631 ( .AN(net104721), .B(n4717), .Y(n4716) );
  AOI21XL U7632 ( .A0(n8529), .A1(n8528), .B0(n3969), .Y(n4717) );
  CLKMX2X2 U7633 ( .A(n8458), .B(n8457), .S0(net114079), .Y(net109201) );
  CLKMX2X2 U7634 ( .A(n8198), .B(n8197), .S0(net114081), .Y(net109673) );
  CLKMX2X2 U7635 ( .A(n7378), .B(n7377), .S0(net114081), .Y(net111128) );
  CLKMX2X2 U7636 ( .A(n8278), .B(n8277), .S0(net114081), .Y(net109527) );
  CLKMX2X2 U7637 ( .A(n7562), .B(n7561), .S0(net114081), .Y(net110798) );
  OA22X2 U7638 ( .A0(n5239), .A1(n634), .B0(n5278), .B1(n2251), .Y(n9519) );
  OA22X1 U7639 ( .A0(n5254), .A1(n990), .B0(n5294), .B1(n2615), .Y(n7905) );
  NAND4X1 U7640 ( .A(n9601), .B(n9820), .C(n9600), .D(n9817), .Y(n11576) );
  OAI222XL U7641 ( .A0(net107217), .A1(n9569), .B0(n9568), .B1(net118592), 
        .C0(n9557), .C1(net117757), .Y(n9558) );
  CLKINVX1 U7642 ( .A(n8567), .Y(n8554) );
  OA22X2 U7643 ( .A0(n5250), .A1(n644), .B0(n5290), .B1(n2261), .Y(n8345) );
  OA22X2 U7644 ( .A0(n5392), .A1(n645), .B0(n5435), .B1(n2262), .Y(n7915) );
  OA22X2 U7645 ( .A0(n5178), .A1(n646), .B0(n5217), .B1(n2263), .Y(n7918) );
  OA22X1 U7646 ( .A0(n5257), .A1(n991), .B0(n5301), .B1(n2616), .Y(n6868) );
  OA22XL U7647 ( .A0(n5182), .A1(n1223), .B0(n5219), .B1(n2846), .Y(n6869) );
  OAI222XL U7648 ( .A0(n5531), .A1(n352), .B0(n5462), .B1(n5530), .C0(n5952), 
        .C1(n10723), .Y(n11542) );
  OAI222XL U7649 ( .A0(n5531), .A1(n233), .B0(n153), .B1(n5530), .C0(n5952), 
        .C1(n10577), .Y(n11543) );
  OAI222XL U7650 ( .A0(n5531), .A1(n230), .B0(n338), .B1(n5530), .C0(n5953), 
        .C1(n10513), .Y(n11551) );
  OAI222XL U7651 ( .A0(n5532), .A1(n158), .B0(n5468), .B1(n5529), .C0(n5953), 
        .C1(n10320), .Y(n11553) );
  OAI222XL U7652 ( .A0(n5531), .A1(n225), .B0(n5510), .B1(n5530), .C0(n5952), 
        .C1(n10633), .Y(n11554) );
  OAI222XL U7653 ( .A0(n5531), .A1(n169), .B0(n5507), .B1(n5530), .C0(n5952), 
        .C1(\i_MIPS/n170 ), .Y(n11555) );
  OAI222XL U7654 ( .A0(n5531), .A1(n229), .B0(n5491), .B1(n5530), .C0(n5953), 
        .C1(\i_MIPS/n169 ), .Y(n11556) );
  OAI222XL U7655 ( .A0(n5531), .A1(n160), .B0(n151), .B1(n5530), .C0(n5953), 
        .C1(\i_MIPS/n168 ), .Y(n11557) );
  OAI222XL U7656 ( .A0(n5531), .A1(n159), .B0(n152), .B1(n5528), .C0(n5952), 
        .C1(\i_MIPS/n166 ), .Y(n11559) );
  OAI222XL U7657 ( .A0(n5531), .A1(n171), .B0(n5486), .B1(n5530), .C0(n5953), 
        .C1(\i_MIPS/n165 ), .Y(n11560) );
  OAI222XL U7658 ( .A0(n5531), .A1(n172), .B0(n4716), .B1(n5528), .C0(n5952), 
        .C1(\i_MIPS/n164 ), .Y(n11561) );
  OAI222XL U7659 ( .A0(n5531), .A1(n164), .B0(n5496), .B1(n5530), .C0(n5952), 
        .C1(\i_MIPS/n163 ), .Y(n11562) );
  OAI222XL U7660 ( .A0(n5531), .A1(n165), .B0(n5504), .B1(n5530), .C0(n5952), 
        .C1(\i_MIPS/n162 ), .Y(n11563) );
  OAI222XL U7661 ( .A0(n5531), .A1(n173), .B0(n154), .B1(n5528), .C0(n5952), 
        .C1(\i_MIPS/n161 ), .Y(n11564) );
  OAI222XL U7662 ( .A0(n5531), .A1(n231), .B0(n155), .B1(n5528), .C0(n5952), 
        .C1(\i_MIPS/n160 ), .Y(n11565) );
  OAI222XL U7663 ( .A0(n5532), .A1(n232), .B0(n5457), .B1(n5529), .C0(n5953), 
        .C1(\i_MIPS/n159 ), .Y(n11566) );
  OAI222XL U7664 ( .A0(n5532), .A1(n226), .B0(n341), .B1(n5529), .C0(n5953), 
        .C1(\i_MIPS/n158 ), .Y(n11567) );
  OAI222XL U7665 ( .A0(n5532), .A1(n359), .B0(n157), .B1(n5529), .C0(n5952), 
        .C1(\i_MIPS/n157 ), .Y(n11568) );
  OAI222XL U7666 ( .A0(n5532), .A1(n228), .B0(n1986), .B1(n5529), .C0(n5952), 
        .C1(\i_MIPS/n156 ), .Y(n11569) );
  OAI222XL U7667 ( .A0(n5531), .A1(n170), .B0(n357), .B1(n5528), .C0(n5953), 
        .C1(\i_MIPS/n154 ), .Y(n11571) );
  OAI222XL U7668 ( .A0(n5531), .A1(n227), .B0(n342), .B1(n5528), .C0(n5952), 
        .C1(\i_MIPS/n153 ), .Y(n11572) );
  OAI222XL U7669 ( .A0(n5531), .A1(n224), .B0(n166), .B1(n5529), .C0(n5953), 
        .C1(\i_MIPS/n177 ), .Y(n11548) );
  OAI222XL U7670 ( .A0(n5531), .A1(n167), .B0(n354), .B1(n5530), .C0(n5953), 
        .C1(\i_MIPS/n167 ), .Y(n11558) );
  OA22X1 U7671 ( .A0(n5648), .A1(n1347), .B0(n5604), .B1(n3034), .Y(n10816) );
  OA22X1 U7672 ( .A0(n5827), .A1(n1348), .B0(n5782), .B1(n3035), .Y(n10814) );
  OA22X1 U7673 ( .A0(n5738), .A1(n1349), .B0(n5691), .B1(n3036), .Y(n10815) );
  OA22X1 U7674 ( .A0(n5644), .A1(n1350), .B0(n5600), .B1(n3037), .Y(n10042) );
  OA22X1 U7675 ( .A0(n5823), .A1(n1351), .B0(n5778), .B1(n3038), .Y(n10040) );
  OA22X1 U7676 ( .A0(n5734), .A1(n1352), .B0(n5687), .B1(n3039), .Y(n10041) );
  NAND4X1 U7677 ( .A(n10837), .B(n10836), .C(n10835), .D(n10834), .Y(n11242)
         );
  OA22X1 U7678 ( .A0(n5648), .A1(n1353), .B0(n5604), .B1(n3040), .Y(n10837) );
  OA22X1 U7679 ( .A0(n5827), .A1(n1354), .B0(n5782), .B1(n3041), .Y(n10835) );
  OA22X1 U7680 ( .A0(n5738), .A1(n1355), .B0(n5691), .B1(n3042), .Y(n10836) );
  NAND4X1 U7681 ( .A(n10020), .B(n10019), .C(n10018), .D(n10017), .Y(n11241)
         );
  OA22X1 U7682 ( .A0(n5643), .A1(n1356), .B0(n5599), .B1(n3043), .Y(n10020) );
  OA22X1 U7683 ( .A0(n5822), .A1(n1357), .B0(n5777), .B1(n3044), .Y(n10018) );
  OA22X1 U7684 ( .A0(n5733), .A1(n1358), .B0(n5686), .B1(n3045), .Y(n10019) );
  NAND4X1 U7685 ( .A(n9976), .B(n9975), .C(n9974), .D(n9973), .Y(n11240) );
  OA22X1 U7686 ( .A0(n5642), .A1(n1359), .B0(n5598), .B1(n3046), .Y(n9976) );
  OA22X1 U7687 ( .A0(n5821), .A1(n1360), .B0(n5776), .B1(n3047), .Y(n9974) );
  OA22X1 U7688 ( .A0(n5732), .A1(n1361), .B0(n5685), .B1(n3048), .Y(n9975) );
  NAND4X1 U7689 ( .A(n9998), .B(n9997), .C(n9996), .D(n9995), .Y(n11239) );
  OA22X1 U7690 ( .A0(n5643), .A1(n1362), .B0(n5599), .B1(n3049), .Y(n9998) );
  OA22X1 U7691 ( .A0(n5822), .A1(n1363), .B0(n5777), .B1(n3050), .Y(n9996) );
  OA22X1 U7692 ( .A0(n5733), .A1(n1364), .B0(n5686), .B1(n3051), .Y(n9997) );
  OA22X1 U7693 ( .A0(n5638), .A1(n1365), .B0(n5594), .B1(n3052), .Y(n9787) );
  OA22X1 U7694 ( .A0(n5817), .A1(n1366), .B0(n5772), .B1(n3053), .Y(n9785) );
  OA22X1 U7695 ( .A0(n5728), .A1(n1367), .B0(n5681), .B1(n3054), .Y(n9786) );
  NAND4X1 U7696 ( .A(n11084), .B(n11083), .C(n11082), .D(n11081), .Y(n11237)
         );
  OA22XL U7697 ( .A0(n5651), .A1(n1593), .B0(n5607), .B1(n3280), .Y(n11084) );
  OA22XL U7698 ( .A0(n5830), .A1(n1594), .B0(n5785), .B1(n3281), .Y(n11082) );
  OA22XL U7699 ( .A0(n5741), .A1(n1595), .B0(n5702), .B1(n3282), .Y(n11083) );
  OA22X1 U7700 ( .A0(n5637), .A1(n1368), .B0(n5593), .B1(n3055), .Y(net106692)
         );
  OA22X1 U7701 ( .A0(n5816), .A1(n1369), .B0(n5771), .B1(n3056), .Y(net106694)
         );
  OA22X1 U7702 ( .A0(n5727), .A1(n1370), .B0(n5680), .B1(n3057), .Y(net106693)
         );
  OA22X1 U7703 ( .A0(n5636), .A1(n3033), .B0(n5592), .B1(n1345), .Y(n9739) );
  OA22X1 U7704 ( .A0(n5815), .A1(n1371), .B0(n5770), .B1(n3058), .Y(n9737) );
  OA22X1 U7705 ( .A0(n5726), .A1(n1372), .B0(n5679), .B1(n3059), .Y(n9738) );
  NAND4X1 U7706 ( .A(n9761), .B(n9760), .C(n9759), .D(n9758), .Y(n11235) );
  OA22X1 U7707 ( .A0(n5637), .A1(n1373), .B0(n5593), .B1(n3060), .Y(n9761) );
  OA22X1 U7708 ( .A0(n5816), .A1(n1374), .B0(n5771), .B1(n3061), .Y(n9759) );
  OA22X1 U7709 ( .A0(n5727), .A1(n1375), .B0(n5680), .B1(n3062), .Y(n9760) );
  OA22X1 U7710 ( .A0(n5645), .A1(n1376), .B0(n5601), .B1(n3063), .Y(n10066) );
  OA22X1 U7711 ( .A0(n5824), .A1(n1377), .B0(n5779), .B1(n3064), .Y(n10064) );
  OA22X1 U7712 ( .A0(n5735), .A1(n1378), .B0(n5688), .B1(n3065), .Y(n10065) );
  OA22X1 U7713 ( .A0(n5647), .A1(n1379), .B0(n5603), .B1(n3066), .Y(n10245) );
  OA22X1 U7714 ( .A0(n5826), .A1(n1380), .B0(n5781), .B1(n3067), .Y(n10243) );
  OA22X1 U7715 ( .A0(n5737), .A1(n1381), .B0(n5690), .B1(n3068), .Y(n10244) );
  OA22X1 U7716 ( .A0(n5647), .A1(n1382), .B0(n5603), .B1(n3069), .Y(n10223) );
  OA22X1 U7717 ( .A0(n5826), .A1(n1383), .B0(n5781), .B1(n3070), .Y(n10221) );
  OA22X1 U7718 ( .A0(n5737), .A1(n1384), .B0(n5690), .B1(n3071), .Y(n10222) );
  OA22X1 U7719 ( .A0(n5646), .A1(n1385), .B0(n5602), .B1(n3072), .Y(n10125) );
  OA22X1 U7720 ( .A0(n5825), .A1(n1386), .B0(n5780), .B1(n3073), .Y(n10123) );
  OA22X1 U7721 ( .A0(n5736), .A1(n1387), .B0(n5689), .B1(n3074), .Y(n10124) );
  OA22X1 U7722 ( .A0(n5645), .A1(n1388), .B0(n5601), .B1(n3075), .Y(n10089) );
  OA22X1 U7723 ( .A0(n5824), .A1(n1389), .B0(n5779), .B1(n3076), .Y(n10087) );
  OA22X1 U7724 ( .A0(n5735), .A1(n1390), .B0(n5688), .B1(n3077), .Y(n10088) );
  OA22X1 U7725 ( .A0(n5639), .A1(n1391), .B0(n5595), .B1(n3078), .Y(n9838) );
  OA22X1 U7726 ( .A0(n5818), .A1(n1392), .B0(n5773), .B1(n3079), .Y(n9836) );
  OA22X1 U7727 ( .A0(n5729), .A1(n1393), .B0(n5682), .B1(n3080), .Y(n9837) );
  OA22X1 U7728 ( .A0(n5640), .A1(n1394), .B0(n5596), .B1(n3081), .Y(n9882) );
  OA22X1 U7729 ( .A0(n5819), .A1(n1395), .B0(n5774), .B1(n3082), .Y(n9880) );
  OA22X1 U7730 ( .A0(n5730), .A1(n1396), .B0(n5683), .B1(n3083), .Y(n9881) );
  OA22X1 U7731 ( .A0(n5639), .A1(n1397), .B0(n5595), .B1(n3084), .Y(n9860) );
  OA22X1 U7732 ( .A0(n5818), .A1(n1398), .B0(n5773), .B1(n3085), .Y(n9858) );
  OA22X1 U7733 ( .A0(n5729), .A1(n1399), .B0(n5682), .B1(n3086), .Y(n9859) );
  OA22X1 U7734 ( .A0(n5641), .A1(n1400), .B0(n5597), .B1(n3087), .Y(n9904) );
  OA22X1 U7735 ( .A0(n5820), .A1(n1401), .B0(n5775), .B1(n3088), .Y(n9902) );
  OA22X1 U7736 ( .A0(n5731), .A1(n1402), .B0(n5684), .B1(n3089), .Y(n9903) );
  OA22X1 U7737 ( .A0(n5641), .A1(n1403), .B0(n5597), .B1(n3090), .Y(n9926) );
  OA22X1 U7738 ( .A0(n5820), .A1(n1404), .B0(n5775), .B1(n3091), .Y(n9924) );
  OA22X1 U7739 ( .A0(n5731), .A1(n1405), .B0(n5684), .B1(n3092), .Y(n9925) );
  OA22X1 U7740 ( .A0(n5636), .A1(n1406), .B0(n5592), .B1(n3093), .Y(n9719) );
  OA22X1 U7741 ( .A0(n5815), .A1(n1407), .B0(n5770), .B1(n3094), .Y(n9717) );
  OA22X1 U7742 ( .A0(n5726), .A1(n1408), .B0(n5679), .B1(n3095), .Y(n9718) );
  OA22X1 U7743 ( .A0(n5649), .A1(n1409), .B0(n5605), .B1(n3096), .Y(n10859) );
  OA22X1 U7744 ( .A0(n5828), .A1(n1410), .B0(n5783), .B1(n3097), .Y(n10857) );
  OA22X1 U7745 ( .A0(n5739), .A1(n1411), .B0(n5692), .B1(n3098), .Y(n10858) );
  OA22X1 U7746 ( .A0(n5650), .A1(n1412), .B0(n5606), .B1(n3099), .Y(n10953) );
  OA22X1 U7747 ( .A0(n5829), .A1(n1413), .B0(n5784), .B1(n3100), .Y(n10951) );
  OA22X1 U7748 ( .A0(n5740), .A1(n1414), .B0(n5693), .B1(n3101), .Y(n10952) );
  NAND4X1 U7749 ( .A(n10924), .B(n10923), .C(n10922), .D(n10921), .Y(n11221)
         );
  OA22X1 U7750 ( .A0(n5650), .A1(n1415), .B0(n5606), .B1(n3102), .Y(n10924) );
  OA22X1 U7751 ( .A0(n5829), .A1(n1416), .B0(n5784), .B1(n3103), .Y(n10922) );
  OA22X1 U7752 ( .A0(n5740), .A1(n1417), .B0(n5693), .B1(n3104), .Y(n10923) );
  OA22X1 U7753 ( .A0(n5649), .A1(n1418), .B0(n5605), .B1(n3105), .Y(n10882) );
  OA22X1 U7754 ( .A0(n5828), .A1(n1419), .B0(n5783), .B1(n3106), .Y(n10880) );
  OA22X1 U7755 ( .A0(n5739), .A1(n1420), .B0(n5692), .B1(n3107), .Y(n10881) );
  OA22X1 U7756 ( .A0(n5632), .A1(n1421), .B0(n5588), .B1(n3108), .Y(n6586) );
  OA22X1 U7757 ( .A0(n5811), .A1(n1422), .B0(n5766), .B1(n3109), .Y(n6584) );
  OA22X1 U7758 ( .A0(n5722), .A1(n1423), .B0(n5675), .B1(n3110), .Y(n6585) );
  OA22X1 U7759 ( .A0(n5634), .A1(n1424), .B0(n5590), .B1(n3111), .Y(n9675) );
  OA22X1 U7760 ( .A0(n5813), .A1(n1425), .B0(n5768), .B1(n3112), .Y(n9673) );
  OA22X1 U7761 ( .A0(n5724), .A1(n1426), .B0(n5677), .B1(n3113), .Y(n9674) );
  OA22X1 U7762 ( .A0(n5635), .A1(n1427), .B0(n5591), .B1(n3114), .Y(n9697) );
  OA22X1 U7763 ( .A0(n5814), .A1(n1428), .B0(n5769), .B1(n3115), .Y(n9695) );
  OA22X1 U7764 ( .A0(n5725), .A1(n1429), .B0(n5678), .B1(n3116), .Y(n9696) );
  OA22X1 U7765 ( .A0(n5633), .A1(n1430), .B0(n5589), .B1(n3117), .Y(n9645) );
  OA22X1 U7766 ( .A0(n5812), .A1(n1431), .B0(n5767), .B1(n3118), .Y(n9643) );
  OA22X1 U7767 ( .A0(n5723), .A1(n1432), .B0(n5676), .B1(n3119), .Y(n9644) );
  OA22X1 U7768 ( .A0(n5633), .A1(n1433), .B0(n5589), .B1(n3120), .Y(n9623) );
  OA22X1 U7769 ( .A0(n5812), .A1(n1434), .B0(n5767), .B1(n3121), .Y(n9621) );
  OA22X1 U7770 ( .A0(n5723), .A1(n1435), .B0(n5676), .B1(n3122), .Y(n9622) );
  OA22X1 U7771 ( .A0(n5632), .A1(n1436), .B0(n5588), .B1(n3123), .Y(n6601) );
  OA22X1 U7772 ( .A0(n5811), .A1(n1437), .B0(n5766), .B1(n3124), .Y(n6599) );
  OA22X1 U7773 ( .A0(n5722), .A1(n1438), .B0(n5675), .B1(n3125), .Y(n6600) );
  OA22X1 U7774 ( .A0(n5631), .A1(n1601), .B0(n5587), .B1(n3289), .Y(n6551) );
  OA22X1 U7775 ( .A0(n5810), .A1(n1602), .B0(n5765), .B1(n3290), .Y(n6549) );
  OA22X1 U7776 ( .A0(n5721), .A1(n1603), .B0(n5674), .B1(n3291), .Y(n6550) );
  OA22X1 U7777 ( .A0(n5644), .A1(n1604), .B0(n5600), .B1(n3292), .Y(n10032) );
  OA22X1 U7778 ( .A0(n5823), .A1(n1605), .B0(n5778), .B1(n3293), .Y(n10030) );
  OA22X1 U7779 ( .A0(n5734), .A1(n1606), .B0(n5687), .B1(n3294), .Y(n10031) );
  OA22X1 U7780 ( .A0(n5631), .A1(n1607), .B0(n5586), .B1(n3295), .Y(n6546) );
  OA22X1 U7781 ( .A0(n5809), .A1(n1608), .B0(n5764), .B1(n3296), .Y(n6544) );
  OA22X1 U7782 ( .A0(n5720), .A1(n1609), .B0(n5702), .B1(n3297), .Y(n6545) );
  NAND4X1 U7783 ( .A(n10010), .B(n10009), .C(n10008), .D(n10007), .Y(n11272)
         );
  OA22X1 U7784 ( .A0(n5643), .A1(n1610), .B0(n5599), .B1(n3298), .Y(n10010) );
  OA22X1 U7785 ( .A0(n5822), .A1(n1611), .B0(n5777), .B1(n3299), .Y(n10008) );
  OA22X1 U7786 ( .A0(n5733), .A1(n1612), .B0(n5686), .B1(n3300), .Y(n10009) );
  NAND4X1 U7787 ( .A(n9966), .B(n9965), .C(n9964), .D(n9963), .Y(n11271) );
  OA22X1 U7788 ( .A0(n5642), .A1(n1613), .B0(n5598), .B1(n3301), .Y(n9966) );
  OA22X1 U7789 ( .A0(n5821), .A1(n1614), .B0(n5776), .B1(n3302), .Y(n9964) );
  OA22X1 U7790 ( .A0(n5732), .A1(n1615), .B0(n5685), .B1(n3303), .Y(n9965) );
  NAND4X1 U7791 ( .A(n9988), .B(n9987), .C(n9986), .D(n9985), .Y(n11270) );
  OA22X1 U7792 ( .A0(n5642), .A1(n1616), .B0(n5598), .B1(n3304), .Y(n9988) );
  OA22X1 U7793 ( .A0(n5821), .A1(n1617), .B0(n5776), .B1(n3305), .Y(n9986) );
  OA22X1 U7794 ( .A0(n5732), .A1(n1618), .B0(n5685), .B1(n3306), .Y(n9987) );
  OA22X1 U7795 ( .A0(n5638), .A1(n1619), .B0(n5594), .B1(n3307), .Y(n9777) );
  OA22X1 U7796 ( .A0(n5817), .A1(n1620), .B0(n5772), .B1(n3308), .Y(n9775) );
  OA22X1 U7797 ( .A0(n5728), .A1(n1621), .B0(n5681), .B1(n3309), .Y(n9776) );
  NAND4X1 U7798 ( .A(n11072), .B(n11071), .C(n11070), .D(n11069), .Y(n11268)
         );
  OA22XL U7799 ( .A0(n5651), .A1(n1847), .B0(n5607), .B1(n3535), .Y(n11072) );
  OA22XL U7800 ( .A0(n5830), .A1(n1848), .B0(n5785), .B1(n3536), .Y(n11070) );
  OA22XL U7801 ( .A0(n5741), .A1(n1849), .B0(n5702), .B1(n3537), .Y(n11071) );
  OA22X1 U7802 ( .A0(n5637), .A1(n1622), .B0(n5593), .B1(n3310), .Y(net106718)
         );
  OA22X1 U7803 ( .A0(n5816), .A1(n1623), .B0(n5771), .B1(n3311), .Y(net106720)
         );
  OA22X1 U7804 ( .A0(n5727), .A1(n1624), .B0(n5680), .B1(n3312), .Y(net106719)
         );
  NAND4X1 U7805 ( .A(n6566), .B(n6565), .C(n6564), .D(n6563), .Y(n11267) );
  OA22X1 U7806 ( .A0(n5631), .A1(n1625), .B0(n5587), .B1(n3313), .Y(n6566) );
  OA22X1 U7807 ( .A0(n5810), .A1(n1626), .B0(n5765), .B1(n3314), .Y(n6564) );
  OA22X1 U7808 ( .A0(n5721), .A1(n1627), .B0(n5674), .B1(n3315), .Y(n6565) );
  OA22X1 U7809 ( .A0(n5636), .A1(n1346), .B0(n5592), .B1(n3316), .Y(n9751) );
  OA22X1 U7810 ( .A0(n5815), .A1(n1628), .B0(n5770), .B1(n3317), .Y(n9749) );
  OA22X1 U7811 ( .A0(n5726), .A1(n1629), .B0(n5679), .B1(n3318), .Y(n9750) );
  OA22X1 U7812 ( .A0(n5644), .A1(n1630), .B0(n5600), .B1(n3319), .Y(n10056) );
  OA22X1 U7813 ( .A0(n5823), .A1(n1631), .B0(n5778), .B1(n3320), .Y(n10054) );
  OA22X1 U7814 ( .A0(n5734), .A1(n1632), .B0(n5687), .B1(n3321), .Y(n10055) );
  OA22X1 U7815 ( .A0(n5647), .A1(n1633), .B0(n5603), .B1(n3322), .Y(n10235) );
  OA22X1 U7816 ( .A0(n5826), .A1(n1634), .B0(n5781), .B1(n3323), .Y(n10233) );
  OA22X1 U7817 ( .A0(n5737), .A1(n1635), .B0(n5690), .B1(n3324), .Y(n10234) );
  OA22X1 U7818 ( .A0(n5646), .A1(n1636), .B0(n5602), .B1(n3325), .Y(n10213) );
  OA22X1 U7819 ( .A0(n5825), .A1(n1637), .B0(n5780), .B1(n3326), .Y(n10211) );
  OA22X1 U7820 ( .A0(n5736), .A1(n1638), .B0(n5689), .B1(n3327), .Y(n10212) );
  OA22X1 U7821 ( .A0(n5646), .A1(n1639), .B0(n5602), .B1(n3328), .Y(n10115) );
  OA22X1 U7822 ( .A0(n5825), .A1(n1640), .B0(n5780), .B1(n3329), .Y(n10113) );
  OA22X1 U7823 ( .A0(n5736), .A1(n1641), .B0(n5689), .B1(n3330), .Y(n10114) );
  OA22X1 U7824 ( .A0(n5645), .A1(n1642), .B0(n5601), .B1(n3331), .Y(n10079) );
  OA22X1 U7825 ( .A0(n5824), .A1(n1643), .B0(n5779), .B1(n3332), .Y(n10077) );
  OA22X1 U7826 ( .A0(n5735), .A1(n1644), .B0(n5688), .B1(n3333), .Y(n10078) );
  OA22X1 U7827 ( .A0(n5638), .A1(n1645), .B0(n5594), .B1(n3334), .Y(n9828) );
  OA22X1 U7828 ( .A0(n5817), .A1(n1646), .B0(n5772), .B1(n3335), .Y(n9826) );
  OA22X1 U7829 ( .A0(n5728), .A1(n1647), .B0(n5681), .B1(n3336), .Y(n9827) );
  OA22X1 U7830 ( .A0(n5640), .A1(n1648), .B0(n5596), .B1(n3337), .Y(n9872) );
  OA22X1 U7831 ( .A0(n5819), .A1(n1649), .B0(n5774), .B1(n3338), .Y(n9870) );
  OA22X1 U7832 ( .A0(n5730), .A1(n1650), .B0(n5683), .B1(n3339), .Y(n9871) );
  OA22X1 U7833 ( .A0(n5639), .A1(n1651), .B0(n5595), .B1(n3340), .Y(n9850) );
  OA22X1 U7834 ( .A0(n5818), .A1(n1652), .B0(n5773), .B1(n3341), .Y(n9848) );
  OA22X1 U7835 ( .A0(n5729), .A1(n1653), .B0(n5682), .B1(n3342), .Y(n9849) );
  OA22X1 U7836 ( .A0(n5640), .A1(n1654), .B0(n5596), .B1(n3343), .Y(n9894) );
  OA22X1 U7837 ( .A0(n5819), .A1(n1655), .B0(n5774), .B1(n3344), .Y(n9892) );
  OA22X1 U7838 ( .A0(n5730), .A1(n1656), .B0(n5683), .B1(n3345), .Y(n9893) );
  OA22X1 U7839 ( .A0(n5641), .A1(n1657), .B0(n5597), .B1(n3346), .Y(n9916) );
  OA22X1 U7840 ( .A0(n5820), .A1(n1658), .B0(n5775), .B1(n3347), .Y(n9914) );
  OA22X1 U7841 ( .A0(n5731), .A1(n1659), .B0(n5684), .B1(n3348), .Y(n9915) );
  OA22X1 U7842 ( .A0(n5635), .A1(n1660), .B0(n5591), .B1(n3349), .Y(n9709) );
  OA22X1 U7843 ( .A0(n5814), .A1(n1661), .B0(n5769), .B1(n3350), .Y(n9707) );
  OA22X1 U7844 ( .A0(n5725), .A1(n1662), .B0(n5678), .B1(n3351), .Y(n9708) );
  OA22X1 U7845 ( .A0(n5630), .A1(n1663), .B0(n5586), .B1(n3352), .Y(n6541) );
  OA22X1 U7846 ( .A0(n5809), .A1(n1664), .B0(n5764), .B1(n3353), .Y(n6539) );
  OA22X1 U7847 ( .A0(n5720), .A1(n1665), .B0(n5673), .B1(n3354), .Y(n6540) );
  OA22X1 U7848 ( .A0(n5650), .A1(n1666), .B0(n5606), .B1(n3355), .Y(n10943) );
  OA22X1 U7849 ( .A0(n5829), .A1(n1667), .B0(n5784), .B1(n3356), .Y(n10941) );
  OA22X1 U7850 ( .A0(n5740), .A1(n1668), .B0(n5693), .B1(n3357), .Y(n10942) );
  OA22X1 U7851 ( .A0(n5636), .A1(n1669), .B0(n5612), .B1(n3358), .Y(n6533) );
  OA22X1 U7852 ( .A0(n5838), .A1(n1670), .B0(n5794), .B1(n3359), .Y(n6531) );
  OA22X1 U7853 ( .A0(n5720), .A1(n1671), .B0(n5702), .B1(n3360), .Y(n6532) );
  OA22X1 U7854 ( .A0(n5630), .A1(n221), .B0(n5586), .B1(n1850), .Y(n6537) );
  OA22X1 U7855 ( .A0(n5809), .A1(n1672), .B0(n5764), .B1(n3361), .Y(n6535) );
  OA22X1 U7856 ( .A0(n5720), .A1(n1673), .B0(n5673), .B1(n349), .Y(n6536) );
  OA22X1 U7857 ( .A0(n5631), .A1(n1674), .B0(n5587), .B1(n3362), .Y(n6576) );
  OA22X1 U7858 ( .A0(n5810), .A1(n1675), .B0(n5765), .B1(n3363), .Y(n6574) );
  OA22X1 U7859 ( .A0(n5721), .A1(n1676), .B0(n5674), .B1(n3364), .Y(n6575) );
  OA22X1 U7860 ( .A0(n5634), .A1(n1677), .B0(n5590), .B1(n3365), .Y(n9665) );
  OA22X1 U7861 ( .A0(n5813), .A1(n1678), .B0(n5768), .B1(n3366), .Y(n9663) );
  OA22X1 U7862 ( .A0(n5724), .A1(n1679), .B0(n5677), .B1(n3367), .Y(n9664) );
  OA22X1 U7863 ( .A0(n5635), .A1(n1680), .B0(n5591), .B1(n3368), .Y(n9687) );
  OA22X1 U7864 ( .A0(n5814), .A1(n1681), .B0(n5769), .B1(n3369), .Y(n9685) );
  OA22X1 U7865 ( .A0(n5725), .A1(n1682), .B0(n5678), .B1(n3370), .Y(n9686) );
  OA22X1 U7866 ( .A0(n5633), .A1(n1683), .B0(n5589), .B1(n3371), .Y(n9635) );
  OA22X1 U7867 ( .A0(n5812), .A1(n1684), .B0(n5767), .B1(n3372), .Y(n9633) );
  OA22X1 U7868 ( .A0(n5723), .A1(n1685), .B0(n5676), .B1(n3373), .Y(n9634) );
  OA22X1 U7869 ( .A0(n5632), .A1(n1686), .B0(n5588), .B1(n3374), .Y(n9613) );
  OA22X1 U7870 ( .A0(n5811), .A1(n1687), .B0(n5766), .B1(n3375), .Y(n9611) );
  OA22X1 U7871 ( .A0(n5722), .A1(n1688), .B0(n5675), .B1(n3376), .Y(n9612) );
  OA22X1 U7872 ( .A0(n5632), .A1(n1689), .B0(n5588), .B1(n3377), .Y(n6591) );
  OA22X1 U7873 ( .A0(n5811), .A1(n1690), .B0(n5766), .B1(n3378), .Y(n6589) );
  OA22X1 U7874 ( .A0(n5722), .A1(n1691), .B0(n5675), .B1(n3379), .Y(n6590) );
  OA22X1 U7875 ( .A0(n5631), .A1(n1692), .B0(n5587), .B1(n3380), .Y(n6556) );
  OA22X1 U7876 ( .A0(n5810), .A1(n1693), .B0(n5765), .B1(n3381), .Y(n6554) );
  OA22X1 U7877 ( .A0(n5721), .A1(n1694), .B0(n5674), .B1(n3382), .Y(n6555) );
  OA22X1 U7878 ( .A0(n5644), .A1(n1695), .B0(n5600), .B1(n3383), .Y(n10037) );
  OA22X1 U7879 ( .A0(n5823), .A1(n1696), .B0(n5778), .B1(n3384), .Y(n10035) );
  OA22X1 U7880 ( .A0(n5734), .A1(n1697), .B0(n5687), .B1(n3385), .Y(n10036) );
  NAND4X1 U7881 ( .A(n10832), .B(n10831), .C(n10830), .D(n10829), .Y(n11304)
         );
  OA22X1 U7882 ( .A0(n5648), .A1(n1698), .B0(n5604), .B1(n3386), .Y(n10832) );
  OA22X1 U7883 ( .A0(n5827), .A1(n1699), .B0(n5782), .B1(n3387), .Y(n10830) );
  OA22X1 U7884 ( .A0(n5738), .A1(n1700), .B0(n5691), .B1(n3388), .Y(n10831) );
  NAND4X1 U7885 ( .A(n10015), .B(n10014), .C(n10013), .D(n10012), .Y(n11303)
         );
  OA22X1 U7886 ( .A0(n5643), .A1(n1701), .B0(n5599), .B1(n3389), .Y(n10015) );
  OA22X1 U7887 ( .A0(n5822), .A1(n1702), .B0(n5777), .B1(n3390), .Y(n10013) );
  OA22X1 U7888 ( .A0(n5733), .A1(n1703), .B0(n5686), .B1(n3391), .Y(n10014) );
  NAND4X1 U7889 ( .A(n9971), .B(n9970), .C(n9969), .D(n9968), .Y(n11302) );
  OA22X1 U7890 ( .A0(n5642), .A1(n1704), .B0(n5598), .B1(n3392), .Y(n9971) );
  OA22X1 U7891 ( .A0(n5821), .A1(n1705), .B0(n5776), .B1(n3393), .Y(n9969) );
  OA22X1 U7892 ( .A0(n5732), .A1(n1706), .B0(n5685), .B1(n3394), .Y(n9970) );
  NAND4X1 U7893 ( .A(n9993), .B(n9992), .C(n9991), .D(n9990), .Y(n11301) );
  OA22X1 U7894 ( .A0(n5642), .A1(n1707), .B0(n5598), .B1(n3395), .Y(n9993) );
  OA22X1 U7895 ( .A0(n5821), .A1(n1708), .B0(n5776), .B1(n3396), .Y(n9991) );
  OA22X1 U7896 ( .A0(n5732), .A1(n1709), .B0(n5685), .B1(n3397), .Y(n9992) );
  OA22X1 U7897 ( .A0(n5638), .A1(n1710), .B0(n5594), .B1(n3398), .Y(n9782) );
  OA22X1 U7898 ( .A0(n5817), .A1(n1711), .B0(n5772), .B1(n3399), .Y(n9780) );
  OA22X1 U7899 ( .A0(n5728), .A1(n1712), .B0(n5681), .B1(n3400), .Y(n9781) );
  NAND4X1 U7900 ( .A(n11078), .B(n11077), .C(n11076), .D(n11075), .Y(n11299)
         );
  OA22XL U7901 ( .A0(n5651), .A1(n1851), .B0(n5607), .B1(n3538), .Y(n11078) );
  OA22XL U7902 ( .A0(n5830), .A1(n1852), .B0(n5785), .B1(n3539), .Y(n11076) );
  OA22XL U7903 ( .A0(n5741), .A1(n1853), .B0(n5702), .B1(n3540), .Y(n11077) );
  OA22X1 U7904 ( .A0(n5637), .A1(n1713), .B0(n5593), .B1(n3401), .Y(net106705)
         );
  OA22X1 U7905 ( .A0(n5816), .A1(n1714), .B0(n5771), .B1(n3402), .Y(net106707)
         );
  OA22X1 U7906 ( .A0(n5727), .A1(n1715), .B0(n5680), .B1(n3403), .Y(net106706)
         );
  NAND4X1 U7907 ( .A(n6571), .B(n6570), .C(n6569), .D(n6568), .Y(n11298) );
  OA22X1 U7908 ( .A0(n5631), .A1(n1716), .B0(n5587), .B1(n3404), .Y(n6571) );
  OA22X1 U7909 ( .A0(n5810), .A1(n1717), .B0(n5765), .B1(n3405), .Y(n6569) );
  OA22X1 U7910 ( .A0(n5721), .A1(n1718), .B0(n5674), .B1(n3406), .Y(n6570) );
  NAND4X1 U7911 ( .A(n9756), .B(n9755), .C(n9754), .D(n9753), .Y(n11297) );
  OA22X1 U7912 ( .A0(n5636), .A1(n1719), .B0(n5592), .B1(n3407), .Y(n9756) );
  OA22X1 U7913 ( .A0(n5815), .A1(n1720), .B0(n5770), .B1(n3408), .Y(n9754) );
  OA22X1 U7914 ( .A0(n5726), .A1(n1721), .B0(n5679), .B1(n3409), .Y(n9755) );
  OA22X1 U7915 ( .A0(n5644), .A1(n1722), .B0(n5600), .B1(n3410), .Y(n10061) );
  OA22X1 U7916 ( .A0(n5823), .A1(n1723), .B0(n5778), .B1(n3411), .Y(n10059) );
  OA22X1 U7917 ( .A0(n5734), .A1(n1724), .B0(n5687), .B1(n3412), .Y(n10060) );
  OA22X1 U7918 ( .A0(n5647), .A1(n1725), .B0(n5603), .B1(n3413), .Y(n10240) );
  OA22X1 U7919 ( .A0(n5826), .A1(n1726), .B0(n5781), .B1(n3414), .Y(n10238) );
  OA22X1 U7920 ( .A0(n5737), .A1(n1727), .B0(n5690), .B1(n3415), .Y(n10239) );
  OA22X1 U7921 ( .A0(n5646), .A1(n1728), .B0(n5602), .B1(n3416), .Y(n10218) );
  OA22X1 U7922 ( .A0(n5825), .A1(n1729), .B0(n5780), .B1(n3417), .Y(n10216) );
  OA22X1 U7923 ( .A0(n5736), .A1(n1730), .B0(n5689), .B1(n3418), .Y(n10217) );
  OA22X1 U7924 ( .A0(n5646), .A1(n1731), .B0(n5602), .B1(n3419), .Y(n10120) );
  OA22X1 U7925 ( .A0(n5825), .A1(n1732), .B0(n5780), .B1(n3420), .Y(n10118) );
  OA22X1 U7926 ( .A0(n5736), .A1(n1733), .B0(n5689), .B1(n3421), .Y(n10119) );
  OA22X1 U7927 ( .A0(n5645), .A1(n1734), .B0(n5601), .B1(n3422), .Y(n10084) );
  OA22X1 U7928 ( .A0(n5824), .A1(n1735), .B0(n5779), .B1(n3423), .Y(n10082) );
  OA22X1 U7929 ( .A0(n5735), .A1(n1736), .B0(n5688), .B1(n3424), .Y(n10083) );
  OA22X1 U7930 ( .A0(n5638), .A1(n1737), .B0(n5594), .B1(n3425), .Y(n9833) );
  OA22X1 U7931 ( .A0(n5817), .A1(n1738), .B0(n5772), .B1(n3426), .Y(n9831) );
  OA22X1 U7932 ( .A0(n5728), .A1(n1739), .B0(n5681), .B1(n3427), .Y(n9832) );
  OA22X1 U7933 ( .A0(n5640), .A1(n1740), .B0(n5596), .B1(n3428), .Y(n9877) );
  OA22X1 U7934 ( .A0(n5819), .A1(n1741), .B0(n5774), .B1(n3429), .Y(n9875) );
  OA22X1 U7935 ( .A0(n5730), .A1(n1742), .B0(n5683), .B1(n3430), .Y(n9876) );
  OA22X1 U7936 ( .A0(n5639), .A1(n1743), .B0(n5595), .B1(n3431), .Y(n9855) );
  OA22X1 U7937 ( .A0(n5818), .A1(n1744), .B0(n5773), .B1(n3432), .Y(n9853) );
  OA22X1 U7938 ( .A0(n5729), .A1(n1745), .B0(n5682), .B1(n3433), .Y(n9854) );
  OA22X1 U7939 ( .A0(n5640), .A1(n1746), .B0(n5596), .B1(n3434), .Y(n9899) );
  OA22X1 U7940 ( .A0(n5819), .A1(n1747), .B0(n5774), .B1(n3435), .Y(n9897) );
  OA22X1 U7941 ( .A0(n5730), .A1(n1748), .B0(n5683), .B1(n3436), .Y(n9898) );
  OA22X1 U7942 ( .A0(n5641), .A1(n1749), .B0(n5597), .B1(n3437), .Y(n9921) );
  OA22X1 U7943 ( .A0(n5820), .A1(n1750), .B0(n5775), .B1(n3438), .Y(n9919) );
  OA22X1 U7944 ( .A0(n5731), .A1(n1751), .B0(n5684), .B1(n3439), .Y(n9920) );
  OA22X1 U7945 ( .A0(n5635), .A1(n1752), .B0(n5591), .B1(n3440), .Y(n9714) );
  OA22X1 U7946 ( .A0(n5814), .A1(n1753), .B0(n5769), .B1(n3441), .Y(n9712) );
  OA22X1 U7947 ( .A0(n5725), .A1(n1754), .B0(n5678), .B1(n3442), .Y(n9713) );
  OA22X1 U7948 ( .A0(n5648), .A1(n1755), .B0(n5604), .B1(n3443), .Y(n10854) );
  OA22X1 U7949 ( .A0(n5827), .A1(n1756), .B0(n5782), .B1(n3444), .Y(n10852) );
  OA22X1 U7950 ( .A0(n5738), .A1(n1757), .B0(n5691), .B1(n3445), .Y(n10853) );
  OA22X1 U7951 ( .A0(n5650), .A1(n1758), .B0(n5606), .B1(n3446), .Y(n10948) );
  OA22X1 U7952 ( .A0(n5829), .A1(n1759), .B0(n5784), .B1(n3447), .Y(n10946) );
  OA22X1 U7953 ( .A0(n5740), .A1(n1760), .B0(n5693), .B1(n3448), .Y(n10947) );
  NAND4X1 U7954 ( .A(n10919), .B(n10918), .C(n10917), .D(n10916), .Y(n11283)
         );
  OA22X1 U7955 ( .A0(n5649), .A1(n1761), .B0(n5605), .B1(n3449), .Y(n10919) );
  OA22X1 U7956 ( .A0(n5828), .A1(n1762), .B0(n5783), .B1(n3450), .Y(n10917) );
  OA22X1 U7957 ( .A0(n5739), .A1(n1763), .B0(n5692), .B1(n3451), .Y(n10918) );
  OA22X1 U7958 ( .A0(n5649), .A1(n1764), .B0(n5605), .B1(n3452), .Y(n10877) );
  OA22X1 U7959 ( .A0(n5828), .A1(n1765), .B0(n5783), .B1(n3453), .Y(n10875) );
  OA22X1 U7960 ( .A0(n5739), .A1(n1766), .B0(n5692), .B1(n3454), .Y(n10876) );
  OA22X1 U7961 ( .A0(n5631), .A1(n1767), .B0(n5587), .B1(n3455), .Y(n6581) );
  OA22X1 U7962 ( .A0(n5810), .A1(n1768), .B0(n5765), .B1(n3456), .Y(n6579) );
  OA22X1 U7963 ( .A0(n5721), .A1(n1769), .B0(n5674), .B1(n3457), .Y(n6580) );
  OA22X1 U7964 ( .A0(n5634), .A1(n1770), .B0(n5590), .B1(n3458), .Y(n9670) );
  OA22X1 U7965 ( .A0(n5813), .A1(n1771), .B0(n5768), .B1(n3459), .Y(n9668) );
  OA22X1 U7966 ( .A0(n5724), .A1(n1772), .B0(n5677), .B1(n3460), .Y(n9669) );
  OA22X1 U7967 ( .A0(n5635), .A1(n1773), .B0(n5591), .B1(n3461), .Y(n9692) );
  OA22X1 U7968 ( .A0(n5814), .A1(n1774), .B0(n5769), .B1(n3462), .Y(n9690) );
  OA22X1 U7969 ( .A0(n5725), .A1(n1775), .B0(n5678), .B1(n3463), .Y(n9691) );
  OA22X1 U7970 ( .A0(n5633), .A1(n1776), .B0(n5589), .B1(n3464), .Y(n9640) );
  OA22X1 U7971 ( .A0(n5812), .A1(n1777), .B0(n5767), .B1(n3465), .Y(n9638) );
  OA22X1 U7972 ( .A0(n5723), .A1(n1778), .B0(n5676), .B1(n3466), .Y(n9639) );
  OA22X1 U7973 ( .A0(n5633), .A1(n1779), .B0(n5589), .B1(n3467), .Y(n9618) );
  OA22X1 U7974 ( .A0(n5812), .A1(n1780), .B0(n5767), .B1(n3468), .Y(n9616) );
  OA22X1 U7975 ( .A0(n5723), .A1(n1781), .B0(n5676), .B1(n3469), .Y(n9617) );
  OA22X1 U7976 ( .A0(n5632), .A1(n1782), .B0(n5588), .B1(n3470), .Y(n6596) );
  OA22X1 U7977 ( .A0(n5811), .A1(n1783), .B0(n5766), .B1(n3471), .Y(n6594) );
  OA22X1 U7978 ( .A0(n5722), .A1(n1784), .B0(n5675), .B1(n3472), .Y(n6595) );
  OA22X2 U7979 ( .A0(n5241), .A1(n650), .B0(n5279), .B1(n2267), .Y(n9418) );
  OA22X2 U7980 ( .A0(n5386), .A1(n652), .B0(n5427), .B1(n2269), .Y(n9169) );
  OA22X2 U7981 ( .A0(n5176), .A1(n653), .B0(n5215), .B1(n2270), .Y(n9172) );
  OA22X2 U7982 ( .A0(n5375), .A1(n715), .B0(n5421), .B1(n2337), .Y(n9521) );
  OA22X2 U7983 ( .A0(n5238), .A1(n716), .B0(n5289), .B1(n2338), .Y(n9523) );
  OA22X2 U7984 ( .A0(n5241), .A1(n655), .B0(n5280), .B1(n2272), .Y(n9410) );
  OA22X2 U7985 ( .A0(n5380), .A1(n659), .B0(n5439), .B1(n2276), .Y(n9404) );
  OA22X2 U7986 ( .A0(n5242), .A1(n660), .B0(n5281), .B1(n2277), .Y(n9406) );
  OA22X2 U7987 ( .A0(n5177), .A1(n661), .B0(n5216), .B1(n2278), .Y(n9407) );
  OA22X2 U7988 ( .A0(n5386), .A1(n565), .B0(n5427), .B1(n2280), .Y(n9165) );
  OA22X1 U7989 ( .A0(n5245), .A1(n992), .B0(n5286), .B1(n2617), .Y(n9167) );
  OA22X2 U7990 ( .A0(n5390), .A1(n664), .B0(n5432), .B1(n2282), .Y(n8331) );
  OA22X1 U7991 ( .A0(n5257), .A1(n993), .B0(n5287), .B1(n2618), .Y(n7067) );
  OA22X1 U7992 ( .A0(n5253), .A1(n994), .B0(n5293), .B1(n2619), .Y(n7990) );
  OA22X2 U7993 ( .A0(n5394), .A1(n670), .B0(n5437), .B1(n2288), .Y(n7615) );
  OA22X1 U7994 ( .A0(n5256), .A1(n995), .B0(n5296), .B1(n2620), .Y(n7617) );
  OA22X2 U7995 ( .A0(n5179), .A1(n671), .B0(n5213), .B1(n2289), .Y(n7618) );
  OA22X1 U7996 ( .A0(n5254), .A1(n996), .B0(n5287), .B1(n2621), .Y(n6971) );
  OA22XL U7997 ( .A0(n5182), .A1(n1224), .B0(n5219), .B1(n2847), .Y(n6972) );
  OA22X1 U7998 ( .A0(n5254), .A1(n997), .B0(n5287), .B1(n2622), .Y(n7071) );
  OA22X2 U7999 ( .A0(n5383), .A1(n675), .B0(n5424), .B1(n2293), .Y(n9350) );
  OA22X1 U8000 ( .A0(n5266), .A1(n998), .B0(n5283), .B1(n2623), .Y(n9352) );
  OA22X2 U8001 ( .A0(n5394), .A1(n677), .B0(n5437), .B1(n2295), .Y(n7619) );
  OA22X1 U8002 ( .A0(n5255), .A1(n999), .B0(n5296), .B1(n2624), .Y(n7621) );
  OA22X2 U8003 ( .A0(n5179), .A1(n678), .B0(n5213), .B1(n2296), .Y(n7622) );
  OA22X2 U8004 ( .A0(n5382), .A1(n679), .B0(n5423), .B1(n2297), .Y(n9354) );
  OA22X2 U8005 ( .A0(n5177), .A1(n680), .B0(n5216), .B1(n2298), .Y(n9357) );
  OA22X2 U8006 ( .A0(n5393), .A1(n681), .B0(n5436), .B1(n2299), .Y(n7705) );
  OA22X1 U8007 ( .A0(n5255), .A1(n1000), .B0(n5295), .B1(n2625), .Y(n7707) );
  OA22X1 U8008 ( .A0(n5254), .A1(n1001), .B0(n5309), .B1(n2626), .Y(n7063) );
  OA22X2 U8009 ( .A0(n5384), .A1(n687), .B0(n5425), .B1(n2305), .Y(n9346) );
  OA22X2 U8010 ( .A0(n5177), .A1(n688), .B0(n5216), .B1(n2306), .Y(n9349) );
  OA22X2 U8011 ( .A0(n5394), .A1(n691), .B0(n5437), .B1(n2309), .Y(n7611) );
  OA22X1 U8012 ( .A0(n5266), .A1(n1002), .B0(n5296), .B1(n2627), .Y(n7613) );
  OA22X1 U8013 ( .A0(n5392), .A1(n1003), .B0(n5435), .B1(n2628), .Y(n7911) );
  OA22X1 U8014 ( .A0(n5254), .A1(n1004), .B0(n5294), .B1(n2629), .Y(n7913) );
  OA22X1 U8015 ( .A0(n5178), .A1(n1005), .B0(n5217), .B1(n2630), .Y(n7914) );
  OA22X1 U8016 ( .A0(n5397), .A1(n1006), .B0(n5441), .B1(n2631), .Y(n7106) );
  OA22X1 U8017 ( .A0(n3984), .A1(n1007), .B0(n5300), .B1(n2632), .Y(n7108) );
  OA22X1 U8018 ( .A0(n5181), .A1(n1008), .B0(n5218), .B1(n2633), .Y(n7109) );
  OA22X1 U8019 ( .A0(n5397), .A1(n1009), .B0(n5441), .B1(n2634), .Y(n7185) );
  OA22X1 U8020 ( .A0(n5250), .A1(n1010), .B0(n5300), .B1(n2635), .Y(n7187) );
  OA22X1 U8021 ( .A0(n5181), .A1(n949), .B0(n5218), .B1(n2636), .Y(n7188) );
  OA22X1 U8022 ( .A0(n5393), .A1(n1011), .B0(n5436), .B1(n2637), .Y(n7801) );
  OA22X1 U8023 ( .A0(n5179), .A1(n1012), .B0(n5218), .B1(n2638), .Y(n7804) );
  OA22X1 U8024 ( .A0(n5399), .A1(n1013), .B0(n5443), .B1(n2639), .Y(n6747) );
  OA22X1 U8025 ( .A0(n5257), .A1(n1014), .B0(n5301), .B1(n2640), .Y(n6749) );
  OA22XL U8026 ( .A0(n5182), .A1(n1225), .B0(n5219), .B1(n2848), .Y(n6750) );
  NAND4X1 U8027 ( .A(n6857), .B(n6856), .C(n6855), .D(n6854), .Y(n11497) );
  OA22X1 U8028 ( .A0(n5399), .A1(n1243), .B0(n5443), .B1(n2863), .Y(n6854) );
  OA22X1 U8029 ( .A0(n5257), .A1(n1244), .B0(n5301), .B1(n2864), .Y(n6856) );
  OA22XL U8030 ( .A0(n5182), .A1(n1257), .B0(n5219), .B1(n2877), .Y(n6857) );
  OA22X1 U8031 ( .A0(n5393), .A1(n1015), .B0(n5436), .B1(n2641), .Y(n7797) );
  OA22X1 U8032 ( .A0(n5179), .A1(n1016), .B0(n5213), .B1(n2642), .Y(n7800) );
  OA22XL U8033 ( .A0(n5258), .A1(n1258), .B0(n5291), .B1(n2878), .Y(n6741) );
  OA22XL U8034 ( .A0(n5182), .A1(n1259), .B0(n5219), .B1(n2879), .Y(n6742) );
  OA22XL U8035 ( .A0(n5751), .A1(n1226), .B0(n5695), .B1(n2849), .Y(n11170) );
  NAND4X1 U8036 ( .A(n10821), .B(n10820), .C(n10819), .D(n10818), .Y(n11312)
         );
  OA22X1 U8037 ( .A0(n5648), .A1(n1439), .B0(n5604), .B1(n3126), .Y(n10821) );
  OA22X1 U8038 ( .A0(n5827), .A1(n1440), .B0(n5782), .B1(n3127), .Y(n10819) );
  OA22X1 U8039 ( .A0(n5738), .A1(n1441), .B0(n5691), .B1(n3128), .Y(n10820) );
  NAND4X1 U8040 ( .A(n10047), .B(n10046), .C(n10045), .D(n10044), .Y(n11336)
         );
  OA22X1 U8041 ( .A0(n5644), .A1(n1442), .B0(n5600), .B1(n3129), .Y(n10047) );
  OA22X1 U8042 ( .A0(n5823), .A1(n1443), .B0(n5778), .B1(n3130), .Y(n10045) );
  OA22X1 U8043 ( .A0(n5734), .A1(n1444), .B0(n5687), .B1(n3131), .Y(n10046) );
  NAND4X1 U8044 ( .A(n10842), .B(n10841), .C(n10840), .D(n10839), .Y(n11335)
         );
  OA22X1 U8045 ( .A0(n5648), .A1(n1445), .B0(n5604), .B1(n3132), .Y(n10842) );
  OA22X1 U8046 ( .A0(n5827), .A1(n1446), .B0(n5782), .B1(n3133), .Y(n10840) );
  OA22X1 U8047 ( .A0(n5738), .A1(n1447), .B0(n5691), .B1(n3134), .Y(n10841) );
  NAND4X1 U8048 ( .A(n10025), .B(n10024), .C(n10023), .D(n10022), .Y(n11334)
         );
  OA22X1 U8049 ( .A0(n5643), .A1(n1448), .B0(n5599), .B1(n3135), .Y(n10025) );
  OA22X1 U8050 ( .A0(n5822), .A1(n1449), .B0(n5777), .B1(n3136), .Y(n10023) );
  OA22X1 U8051 ( .A0(n5733), .A1(n1450), .B0(n5686), .B1(n3137), .Y(n10024) );
  NAND4X1 U8052 ( .A(n9981), .B(n9980), .C(n9979), .D(n9978), .Y(n11333) );
  OA22X1 U8053 ( .A0(n5642), .A1(n1451), .B0(n5598), .B1(n3138), .Y(n9981) );
  OA22X1 U8054 ( .A0(n5821), .A1(n1452), .B0(n5776), .B1(n3139), .Y(n9979) );
  OA22X1 U8055 ( .A0(n5732), .A1(n1453), .B0(n5685), .B1(n3140), .Y(n9980) );
  NAND4X1 U8056 ( .A(n10003), .B(n10002), .C(n10001), .D(n10000), .Y(n11332)
         );
  OA22X1 U8057 ( .A0(n5643), .A1(n1454), .B0(n5599), .B1(n3141), .Y(n10003) );
  OA22X1 U8058 ( .A0(n5822), .A1(n1455), .B0(n5777), .B1(n3142), .Y(n10001) );
  OA22X1 U8059 ( .A0(n5733), .A1(n1456), .B0(n5686), .B1(n3143), .Y(n10002) );
  NAND4X1 U8060 ( .A(n9792), .B(n9791), .C(n9790), .D(n9789), .Y(n11331) );
  OA22X1 U8061 ( .A0(n5638), .A1(n1457), .B0(n5594), .B1(n3144), .Y(n9792) );
  OA22X1 U8062 ( .A0(n5817), .A1(n1458), .B0(n5772), .B1(n3145), .Y(n9790) );
  OA22X1 U8063 ( .A0(n5728), .A1(n1459), .B0(n5681), .B1(n3146), .Y(n9791) );
  NAND4X1 U8064 ( .A(n11090), .B(n11089), .C(n11088), .D(n11087), .Y(n11330)
         );
  OA22XL U8065 ( .A0(n5651), .A1(n1596), .B0(n5607), .B1(n3283), .Y(n11090) );
  OA22XL U8066 ( .A0(n5830), .A1(n1597), .B0(n5785), .B1(n3284), .Y(n11088) );
  OA22XL U8067 ( .A0(n5741), .A1(n1598), .B0(n5702), .B1(n3285), .Y(n11089) );
  OA22X1 U8068 ( .A0(n5637), .A1(n1460), .B0(n5593), .B1(n3147), .Y(net106679)
         );
  OA22X1 U8069 ( .A0(n5816), .A1(n1461), .B0(n5771), .B1(n3148), .Y(net106681)
         );
  OA22X1 U8070 ( .A0(n5727), .A1(n1462), .B0(n5680), .B1(n3149), .Y(net106680)
         );
  NAND4X1 U8071 ( .A(n9744), .B(n9743), .C(n9742), .D(n9741), .Y(n11329) );
  OA22X1 U8072 ( .A0(n5636), .A1(n1463), .B0(n5592), .B1(n3150), .Y(n9744) );
  OA22X1 U8073 ( .A0(n5815), .A1(n1464), .B0(n5770), .B1(n3151), .Y(n9742) );
  OA22X1 U8074 ( .A0(n5726), .A1(n1465), .B0(n5679), .B1(n3152), .Y(n9743) );
  NAND4X1 U8075 ( .A(n9766), .B(n9765), .C(n9764), .D(n9763), .Y(n11328) );
  OA22X1 U8076 ( .A0(n5637), .A1(n1466), .B0(n5593), .B1(n3153), .Y(n9766) );
  OA22X1 U8077 ( .A0(n5816), .A1(n1467), .B0(n5771), .B1(n3154), .Y(n9764) );
  OA22X1 U8078 ( .A0(n5727), .A1(n1468), .B0(n5680), .B1(n3155), .Y(n9765) );
  NAND4X1 U8079 ( .A(n10071), .B(n10070), .C(n10069), .D(n10068), .Y(n11327)
         );
  OA22X1 U8080 ( .A0(n5645), .A1(n1469), .B0(n5601), .B1(n3156), .Y(n10071) );
  OA22X1 U8081 ( .A0(n5824), .A1(n1470), .B0(n5779), .B1(n3157), .Y(n10069) );
  OA22X1 U8082 ( .A0(n5735), .A1(n1471), .B0(n5688), .B1(n3158), .Y(n10070) );
  NAND4X1 U8083 ( .A(n10250), .B(n10249), .C(n10248), .D(n10247), .Y(n11326)
         );
  OA22X1 U8084 ( .A0(n5647), .A1(n1472), .B0(n5603), .B1(n3159), .Y(n10250) );
  OA22X1 U8085 ( .A0(n5826), .A1(n1473), .B0(n5781), .B1(n3160), .Y(n10248) );
  OA22X1 U8086 ( .A0(n5737), .A1(n1474), .B0(n5690), .B1(n3161), .Y(n10249) );
  NAND4X1 U8087 ( .A(n10228), .B(n10227), .C(n10226), .D(n10225), .Y(n11325)
         );
  OA22X1 U8088 ( .A0(n5647), .A1(n1475), .B0(n5603), .B1(n3162), .Y(n10228) );
  OA22X1 U8089 ( .A0(n5826), .A1(n1476), .B0(n5781), .B1(n3163), .Y(n10226) );
  OA22X1 U8090 ( .A0(n5737), .A1(n1477), .B0(n5690), .B1(n3164), .Y(n10227) );
  NAND4X1 U8091 ( .A(n10130), .B(n10129), .C(n10128), .D(n10127), .Y(n11324)
         );
  OA22X1 U8092 ( .A0(n5646), .A1(n1478), .B0(n5602), .B1(n3165), .Y(n10130) );
  OA22X1 U8093 ( .A0(n5825), .A1(n1479), .B0(n5780), .B1(n3166), .Y(n10128) );
  OA22X1 U8094 ( .A0(n5736), .A1(n1480), .B0(n5689), .B1(n3167), .Y(n10129) );
  NAND4X1 U8095 ( .A(n10094), .B(n10093), .C(n10092), .D(n10091), .Y(n11323)
         );
  OA22X1 U8096 ( .A0(n5645), .A1(n1481), .B0(n5601), .B1(n3168), .Y(n10094) );
  OA22X1 U8097 ( .A0(n5824), .A1(n1482), .B0(n5779), .B1(n3169), .Y(n10092) );
  OA22X1 U8098 ( .A0(n5735), .A1(n1483), .B0(n5688), .B1(n3170), .Y(n10093) );
  NAND4X1 U8099 ( .A(n9843), .B(n9842), .C(n9841), .D(n9840), .Y(n11322) );
  OA22X1 U8100 ( .A0(n5639), .A1(n1484), .B0(n5595), .B1(n3171), .Y(n9843) );
  OA22X1 U8101 ( .A0(n5818), .A1(n1485), .B0(n5773), .B1(n3172), .Y(n9841) );
  OA22X1 U8102 ( .A0(n5729), .A1(n1486), .B0(n5682), .B1(n3173), .Y(n9842) );
  NAND4X1 U8103 ( .A(n9887), .B(n9886), .C(n9885), .D(n9884), .Y(n11321) );
  OA22X1 U8104 ( .A0(n5640), .A1(n1487), .B0(n5596), .B1(n3174), .Y(n9887) );
  OA22X1 U8105 ( .A0(n5819), .A1(n1488), .B0(n5774), .B1(n3175), .Y(n9885) );
  OA22X1 U8106 ( .A0(n5730), .A1(n1489), .B0(n5683), .B1(n3176), .Y(n9886) );
  NAND4X1 U8107 ( .A(n9865), .B(n9864), .C(n9863), .D(n9862), .Y(n11320) );
  OA22X1 U8108 ( .A0(n5639), .A1(n1490), .B0(n5595), .B1(n3177), .Y(n9865) );
  OA22X1 U8109 ( .A0(n5818), .A1(n1491), .B0(n5773), .B1(n3178), .Y(n9863) );
  OA22X1 U8110 ( .A0(n5729), .A1(n1492), .B0(n5682), .B1(n3179), .Y(n9864) );
  NAND4X1 U8111 ( .A(n9909), .B(n9908), .C(n9907), .D(n9906), .Y(n11319) );
  OA22X1 U8112 ( .A0(n5641), .A1(n1493), .B0(n5597), .B1(n3180), .Y(n9909) );
  OA22X1 U8113 ( .A0(n5820), .A1(n1494), .B0(n5775), .B1(n3181), .Y(n9907) );
  OA22X1 U8114 ( .A0(n5731), .A1(n1495), .B0(n5684), .B1(n3182), .Y(n9908) );
  NAND4X1 U8115 ( .A(n9931), .B(n9930), .C(n9929), .D(n9928), .Y(n11318) );
  OA22X1 U8116 ( .A0(n5641), .A1(n1496), .B0(n5597), .B1(n3183), .Y(n9931) );
  OA22X1 U8117 ( .A0(n5820), .A1(n1497), .B0(n5775), .B1(n3184), .Y(n9929) );
  OA22X1 U8118 ( .A0(n5731), .A1(n1498), .B0(n5684), .B1(n3185), .Y(n9930) );
  NAND4X1 U8119 ( .A(n9724), .B(n9723), .C(n9722), .D(n9721), .Y(n11317) );
  OA22X1 U8120 ( .A0(n5636), .A1(n1499), .B0(n5592), .B1(n3186), .Y(n9724) );
  OA22X1 U8121 ( .A0(n5815), .A1(n1500), .B0(n5770), .B1(n3187), .Y(n9722) );
  OA22X1 U8122 ( .A0(n5726), .A1(n1501), .B0(n5679), .B1(n3188), .Y(n9723) );
  NAND4X1 U8123 ( .A(n10864), .B(n10863), .C(n10862), .D(n10861), .Y(n11316)
         );
  OA22X1 U8124 ( .A0(n5649), .A1(n1502), .B0(n5605), .B1(n3189), .Y(n10864) );
  OA22X1 U8125 ( .A0(n5828), .A1(n1503), .B0(n5783), .B1(n3190), .Y(n10862) );
  OA22X1 U8126 ( .A0(n5739), .A1(n1504), .B0(n5692), .B1(n3191), .Y(n10863) );
  NAND4X1 U8127 ( .A(n10958), .B(n10957), .C(n10956), .D(n10955), .Y(n11315)
         );
  OA22X1 U8128 ( .A0(n5650), .A1(n1505), .B0(n5606), .B1(n3192), .Y(n10958) );
  OA22X1 U8129 ( .A0(n5829), .A1(n1506), .B0(n5784), .B1(n3193), .Y(n10956) );
  OA22X1 U8130 ( .A0(n5740), .A1(n1507), .B0(n5693), .B1(n3194), .Y(n10957) );
  NAND4X1 U8131 ( .A(n10929), .B(n10928), .C(n10927), .D(n10926), .Y(n11314)
         );
  OA22X1 U8132 ( .A0(n5650), .A1(n1508), .B0(n5606), .B1(n3195), .Y(n10929) );
  OA22X1 U8133 ( .A0(n5829), .A1(n1509), .B0(n5784), .B1(n3196), .Y(n10927) );
  OA22X1 U8134 ( .A0(n5740), .A1(n1510), .B0(n5693), .B1(n3197), .Y(n10928) );
  NAND4X1 U8135 ( .A(n10887), .B(n10886), .C(n10885), .D(n10884), .Y(n11313)
         );
  OA22X1 U8136 ( .A0(n5649), .A1(n1511), .B0(n5605), .B1(n3198), .Y(n10887) );
  OA22X1 U8137 ( .A0(n5828), .A1(n1512), .B0(n5783), .B1(n3199), .Y(n10885) );
  OA22X1 U8138 ( .A0(n5739), .A1(n1513), .B0(n5692), .B1(n3200), .Y(n10886) );
  NAND4X1 U8139 ( .A(n9680), .B(n9679), .C(n9678), .D(n9677), .Y(n11341) );
  OA22X1 U8140 ( .A0(n5634), .A1(n1514), .B0(n5590), .B1(n3201), .Y(n9680) );
  OA22X1 U8141 ( .A0(n5813), .A1(n1515), .B0(n5768), .B1(n3202), .Y(n9678) );
  OA22X1 U8142 ( .A0(n5724), .A1(n1516), .B0(n5677), .B1(n3203), .Y(n9679) );
  NAND4X1 U8143 ( .A(n9702), .B(n9701), .C(n9700), .D(n9699), .Y(n11340) );
  OA22X1 U8144 ( .A0(n5635), .A1(n1517), .B0(n5591), .B1(n3204), .Y(n9702) );
  OA22X1 U8145 ( .A0(n5814), .A1(n1518), .B0(n5769), .B1(n3205), .Y(n9700) );
  OA22X1 U8146 ( .A0(n5725), .A1(n1519), .B0(n5678), .B1(n3206), .Y(n9701) );
  NAND4X1 U8147 ( .A(n9650), .B(n9649), .C(n9648), .D(n9647), .Y(n11339) );
  OA22X1 U8148 ( .A0(n5634), .A1(n1520), .B0(n5590), .B1(n3207), .Y(n9650) );
  OA22X1 U8149 ( .A0(n5813), .A1(n1521), .B0(n5768), .B1(n3208), .Y(n9648) );
  OA22X1 U8150 ( .A0(n5724), .A1(n1522), .B0(n5677), .B1(n3209), .Y(n9649) );
  NAND4X1 U8151 ( .A(n9628), .B(n9627), .C(n9626), .D(n9625), .Y(n11338) );
  OA22X1 U8152 ( .A0(n5633), .A1(n1523), .B0(n5589), .B1(n3210), .Y(n9628) );
  OA22X1 U8153 ( .A0(n5812), .A1(n1524), .B0(n5767), .B1(n3211), .Y(n9626) );
  OA22X1 U8154 ( .A0(n5723), .A1(n1525), .B0(n5676), .B1(n3212), .Y(n9627) );
  NAND4X1 U8155 ( .A(n6606), .B(n6605), .C(n6604), .D(n6603), .Y(n11337) );
  OA22X1 U8156 ( .A0(n5632), .A1(n1526), .B0(n5588), .B1(n3213), .Y(n6606) );
  OA22X1 U8157 ( .A0(n5811), .A1(n1527), .B0(n5766), .B1(n3214), .Y(n6604) );
  OA22X1 U8158 ( .A0(n5722), .A1(n1528), .B0(n5675), .B1(n3215), .Y(n6605) );
  AO22X2 U8159 ( .A0(n5554), .A1(DCACHE_addr[29]), .B0(n5551), .B1(n11533), 
        .Y(n10992) );
  AO22X2 U8160 ( .A0(n5554), .A1(DCACHE_addr[21]), .B0(n5551), .B1(n11525), 
        .Y(n10986) );
  AO22X2 U8161 ( .A0(n5554), .A1(DCACHE_addr[16]), .B0(n5551), .B1(n11520), 
        .Y(n10989) );
  AO22X2 U8162 ( .A0(n5553), .A1(DCACHE_addr[7]), .B0(n5552), .B1(n11511), .Y(
        n11041) );
  AO22X2 U8163 ( .A0(n5554), .A1(DCACHE_addr[8]), .B0(n5552), .B1(n11512), .Y(
        n11044) );
  AO22X2 U8164 ( .A0(n5554), .A1(DCACHE_addr[6]), .B0(n5552), .B1(n11510), .Y(
        n11047) );
  AO22X2 U8165 ( .A0(n5553), .A1(DCACHE_addr[19]), .B0(n5552), .B1(n11523), 
        .Y(n11051) );
  AOI211XL U8166 ( .A0(n4734), .A1(n9544), .B0(n4795), .C0(n4792), .Y(n7151)
         );
  NAND2XL U8167 ( .A(n3637), .B(n3867), .Y(n7149) );
  NOR4X1 U8168 ( .A(n9397), .B(n9396), .C(n9395), .D(n9394), .Y(n9398) );
  AO22X1 U8169 ( .A0(n5124), .A1(n352), .B0(n5120), .B1(n1992), .Y(n9397) );
  AO22X1 U8170 ( .A0(n5137), .A1(n364), .B0(n5128), .B1(n2002), .Y(n9396) );
  AO22X1 U8171 ( .A0(n5150), .A1(n367), .B0(n5145), .B1(n1989), .Y(n9395) );
  NOR4X1 U8172 ( .A(n9388), .B(n9387), .C(n9386), .D(n9385), .Y(n9389) );
  AO22X1 U8173 ( .A0(n5124), .A1(n243), .B0(n5120), .B1(n1995), .Y(n9388) );
  AO22X1 U8174 ( .A0(n5137), .A1(n365), .B0(n5125), .B1(n2003), .Y(n9387) );
  AO22X1 U8175 ( .A0(n5150), .A1(n368), .B0(n5145), .B1(n1990), .Y(n9386) );
  NOR4X1 U8176 ( .A(n9510), .B(n9509), .C(n9508), .D(n9507), .Y(n9511) );
  AO22X1 U8177 ( .A0(n5124), .A1(n222), .B0(n5120), .B1(n373), .Y(n9510) );
  AO22X1 U8178 ( .A0(n5138), .A1(n241), .B0(n5130), .B1(n374), .Y(n9509) );
  AO22X1 U8179 ( .A0(n5148), .A1(n162), .B0(n5145), .B1(n244), .Y(n9508) );
  NOR4X1 U8180 ( .A(n9493), .B(n9492), .C(n9491), .D(n9490), .Y(n9494) );
  AO22X1 U8181 ( .A0(n5122), .A1(n369), .B0(n5120), .B1(n1993), .Y(n9493) );
  AO22X1 U8182 ( .A0(n5138), .A1(n366), .B0(n5130), .B1(n2004), .Y(n9492) );
  AO22X1 U8183 ( .A0(n5148), .A1(n240), .B0(n5145), .B1(n1991), .Y(n9491) );
  NOR4X1 U8184 ( .A(n9590), .B(n9589), .C(n9588), .D(n9587), .Y(n9591) );
  AO22X1 U8185 ( .A0(net118347), .A1(n222), .B0(net118319), .B1(n373), .Y(
        n9590) );
  AO22X1 U8186 ( .A0(net118395), .A1(n241), .B0(net118369), .B1(n374), .Y(
        n9589) );
  AO22X1 U8187 ( .A0(net118441), .A1(n162), .B0(net118417), .B1(n244), .Y(
        n9588) );
  NOR4X1 U8188 ( .A(n6624), .B(n6623), .C(n6622), .D(n6621), .Y(n6625) );
  AO22X1 U8189 ( .A0(n9500), .A1(n224), .B0(n5117), .B1(n2367), .Y(n6624) );
  AO22X1 U8190 ( .A0(n5134), .A1(n774), .B0(n5127), .B1(n2368), .Y(n6623) );
  AO22X1 U8191 ( .A0(n5147), .A1(n775), .B0(n5143), .B1(n2369), .Y(n6622) );
  NOR4X1 U8192 ( .A(n6615), .B(n6614), .C(n6613), .D(n6612), .Y(n6616) );
  AO22X1 U8193 ( .A0(n9500), .A1(n391), .B0(n5117), .B1(n2572), .Y(n6615) );
  AO22X1 U8194 ( .A0(n5134), .A1(n907), .B0(n5127), .B1(n2573), .Y(n6614) );
  AO22X1 U8195 ( .A0(n5147), .A1(n908), .B0(n5143), .B1(n2574), .Y(n6613) );
  NOR4X1 U8196 ( .A(n9480), .B(n9479), .C(n9478), .D(n9477), .Y(n9481) );
  AO22X1 U8197 ( .A0(net118343), .A1(n352), .B0(net118319), .B1(n1992), .Y(
        n9480) );
  NOR4X1 U8198 ( .A(n9581), .B(n9580), .C(n9579), .D(n9578), .Y(n9582) );
  AO22X1 U8199 ( .A0(net118345), .A1(n369), .B0(net118321), .B1(n1993), .Y(
        n9581) );
  NOR4X1 U8200 ( .A(n7758), .B(n7757), .C(n7756), .D(n7755), .Y(n7759) );
  AO22X1 U8201 ( .A0(net118339), .A1(n167), .B0(net118315), .B1(n245), .Y(
        n7758) );
  NOR4X1 U8202 ( .A(n7749), .B(n7748), .C(n7747), .D(n7746), .Y(n7750) );
  AO22X1 U8203 ( .A0(net118337), .A1(n177), .B0(net118313), .B1(n246), .Y(
        n7749) );
  NOR4X1 U8204 ( .A(n9286), .B(n9285), .C(n9284), .D(n9283), .Y(n9287) );
  AO22X1 U8205 ( .A0(n5124), .A1(n169), .B0(n5120), .B1(n2475), .Y(n9286) );
  AO22X1 U8206 ( .A0(n5137), .A1(n854), .B0(n5127), .B1(n2476), .Y(n9285) );
  AO22X1 U8207 ( .A0(n5150), .A1(n855), .B0(n5145), .B1(n2477), .Y(n9284) );
  AO22X1 U8208 ( .A0(n5124), .A1(n856), .B0(n5120), .B1(n2478), .Y(n9277) );
  AO22X1 U8209 ( .A0(n5137), .A1(n857), .B0(n5125), .B1(n2479), .Y(n9276) );
  AO22X1 U8210 ( .A0(n5150), .A1(n858), .B0(n5145), .B1(n2480), .Y(n9275) );
  NOR4X1 U8211 ( .A(n9035), .B(n9034), .C(n9033), .D(n9032), .Y(n9036) );
  AO22X1 U8212 ( .A0(n5124), .A1(n170), .B0(n5120), .B1(n2370), .Y(n9035) );
  AO22X1 U8213 ( .A0(n5137), .A1(n776), .B0(n5127), .B1(n2371), .Y(n9034) );
  AO22X1 U8214 ( .A0(n5150), .A1(n859), .B0(n5145), .B1(n2481), .Y(n9033) );
  NOR4X1 U8215 ( .A(n8272), .B(n8271), .C(n8270), .D(n8269), .Y(n8273) );
  AO22X1 U8216 ( .A0(n5121), .A1(n171), .B0(n5119), .B1(n309), .Y(n8272) );
  AO22X1 U8217 ( .A0(n5135), .A1(n270), .B0(n5127), .B1(n915), .Y(n8271) );
  AO22X1 U8218 ( .A0(n5148), .A1(n860), .B0(n5144), .B1(n2482), .Y(n8270) );
  NOR4X1 U8219 ( .A(n9026), .B(n9025), .C(n9024), .D(n9023), .Y(n9027) );
  AO22X1 U8220 ( .A0(n5124), .A1(n777), .B0(n5120), .B1(n2372), .Y(n9026) );
  AO22X1 U8221 ( .A0(n5137), .A1(n778), .B0(n5128), .B1(n2373), .Y(n9025) );
  AO22X1 U8222 ( .A0(n5150), .A1(n779), .B0(n5145), .B1(n2374), .Y(n9024) );
  NOR4X1 U8223 ( .A(n8263), .B(n8262), .C(n8261), .D(n8260), .Y(n8264) );
  AO22X1 U8224 ( .A0(n5121), .A1(n201), .B0(n5119), .B1(n310), .Y(n8263) );
  AO22X1 U8225 ( .A0(n5135), .A1(n271), .B0(n5127), .B1(n916), .Y(n8262) );
  AO22X1 U8226 ( .A0(n5148), .A1(n861), .B0(n5144), .B1(n2483), .Y(n8261) );
  NOR4X1 U8227 ( .A(n8625), .B(n8624), .C(n8623), .D(n8622), .Y(n8626) );
  AO22X1 U8228 ( .A0(n5123), .A1(n225), .B0(n5119), .B1(n2375), .Y(n8625) );
  AO22X1 U8229 ( .A0(n5136), .A1(n780), .B0(n5129), .B1(n2376), .Y(n8624) );
  AO22X1 U8230 ( .A0(n5149), .A1(n293), .B0(n5140), .B1(n937), .Y(n8623) );
  NOR4X1 U8231 ( .A(n9377), .B(n9376), .C(n9375), .D(n9374), .Y(n9378) );
  AO22X1 U8232 ( .A0(n5124), .A1(n226), .B0(n5120), .B1(n2377), .Y(n9377) );
  AO22X1 U8233 ( .A0(n5137), .A1(n781), .B0(n5128), .B1(n2378), .Y(n9376) );
  AO22X1 U8234 ( .A0(n5150), .A1(n782), .B0(n5145), .B1(n2379), .Y(n9375) );
  AO22X1 U8235 ( .A0(n5123), .A1(n227), .B0(n5119), .B1(n2380), .Y(n8772) );
  AO22X1 U8236 ( .A0(n5136), .A1(n783), .B0(n5129), .B1(n2381), .Y(n8771) );
  AO22X1 U8237 ( .A0(n5149), .A1(n272), .B0(n5140), .B1(n917), .Y(n8770) );
  NOR4X1 U8238 ( .A(n8616), .B(n8615), .C(n8614), .D(n8613), .Y(n8617) );
  AO22X1 U8239 ( .A0(n5123), .A1(n784), .B0(n5119), .B1(n2382), .Y(n8616) );
  AO22X1 U8240 ( .A0(n5136), .A1(n785), .B0(n5129), .B1(n2383), .Y(n8615) );
  AO22X1 U8241 ( .A0(n5149), .A1(n273), .B0(n5140), .B1(n918), .Y(n8614) );
  NOR4X1 U8242 ( .A(n9368), .B(n9367), .C(n9366), .D(n9365), .Y(n9369) );
  AO22X1 U8243 ( .A0(n5124), .A1(n786), .B0(n5120), .B1(n2384), .Y(n9368) );
  AO22X1 U8244 ( .A0(n5137), .A1(n787), .B0(n5128), .B1(n2385), .Y(n9367) );
  AO22X1 U8245 ( .A0(n5150), .A1(n788), .B0(n5145), .B1(n2386), .Y(n9366) );
  AO22X1 U8246 ( .A0(n5123), .A1(n789), .B0(n5119), .B1(n2387), .Y(n8763) );
  AO22X1 U8247 ( .A0(n5136), .A1(n790), .B0(n5129), .B1(n2388), .Y(n8762) );
  AO22X1 U8248 ( .A0(n5149), .A1(n274), .B0(n5140), .B1(n919), .Y(n8761) );
  AO22X1 U8249 ( .A0(n5124), .A1(n228), .B0(n5120), .B1(n2389), .Y(n9195) );
  AO22X1 U8250 ( .A0(n5137), .A1(n791), .B0(n5128), .B1(n2390), .Y(n9194) );
  AO22X1 U8251 ( .A0(n5150), .A1(n792), .B0(n5145), .B1(n2391), .Y(n9193) );
  AO22X1 U8252 ( .A0(n5124), .A1(n793), .B0(n5120), .B1(n2392), .Y(n9186) );
  AO22X1 U8253 ( .A0(n5137), .A1(n794), .B0(n5128), .B1(n2393), .Y(n9185) );
  AO22X1 U8254 ( .A0(n5150), .A1(n795), .B0(n5145), .B1(n2394), .Y(n9184) );
  NOR4X1 U8255 ( .A(n8543), .B(n8542), .C(n8541), .D(n8540), .Y(n8544) );
  AO22X1 U8256 ( .A0(n5123), .A1(n172), .B0(n5119), .B1(n2395), .Y(n8543) );
  AO22X1 U8257 ( .A0(n5136), .A1(n796), .B0(n5129), .B1(n2396), .Y(n8542) );
  AO22X1 U8258 ( .A0(n5149), .A1(n294), .B0(n5140), .B1(n938), .Y(n8541) );
  NOR4X1 U8259 ( .A(n8848), .B(n8847), .C(n8846), .D(n8845), .Y(n8849) );
  AO22X1 U8260 ( .A0(n5123), .A1(n229), .B0(n5119), .B1(n2397), .Y(n8848) );
  AO22X1 U8261 ( .A0(n5136), .A1(n797), .B0(n5129), .B1(n2398), .Y(n8847) );
  AO22X1 U8262 ( .A0(n5149), .A1(n275), .B0(n5140), .B1(n920), .Y(n8846) );
  NOR4X1 U8263 ( .A(n8534), .B(n8533), .C(n8532), .D(n8531), .Y(n8535) );
  AO22X1 U8264 ( .A0(n5123), .A1(n798), .B0(n5119), .B1(n2399), .Y(n8534) );
  AO22X1 U8265 ( .A0(n5136), .A1(n799), .B0(n5129), .B1(n2400), .Y(n8533) );
  AO22X1 U8266 ( .A0(n5149), .A1(n276), .B0(n5140), .B1(n921), .Y(n8532) );
  AO22X1 U8267 ( .A0(n5136), .A1(n862), .B0(n5129), .B1(n2484), .Y(n8451) );
  AO22X1 U8268 ( .A0(n5149), .A1(n295), .B0(n5140), .B1(n939), .Y(n8450) );
  NOR4X1 U8269 ( .A(n8839), .B(n8838), .C(n8837), .D(n8836), .Y(n8840) );
  AO22X1 U8270 ( .A0(n5123), .A1(n800), .B0(n5119), .B1(n2401), .Y(n8839) );
  AO22X1 U8271 ( .A0(n5136), .A1(n801), .B0(n5129), .B1(n2402), .Y(n8838) );
  AO22X1 U8272 ( .A0(n5149), .A1(n277), .B0(n5140), .B1(n922), .Y(n8837) );
  AO22X1 U8273 ( .A0(n5121), .A1(n158), .B0(n5120), .B1(n311), .Y(n8362) );
  AO22X1 U8274 ( .A0(n5135), .A1(n278), .B0(n5125), .B1(n923), .Y(n8361) );
  AO22X1 U8275 ( .A0(n5148), .A1(n863), .B0(n5144), .B1(n2485), .Y(n8360) );
  AO22X1 U8276 ( .A0(n5123), .A1(n864), .B0(n5119), .B1(n2486), .Y(n8443) );
  AO22X1 U8277 ( .A0(n5136), .A1(n865), .B0(n5129), .B1(n2487), .Y(n8442) );
  AO22X1 U8278 ( .A0(n5149), .A1(n296), .B0(n5140), .B1(n940), .Y(n8441) );
  AO22X1 U8279 ( .A0(n5123), .A1(n230), .B0(n5119), .B1(n2488), .Y(n8951) );
  AO22X1 U8280 ( .A0(n5136), .A1(n802), .B0(n5129), .B1(n2403), .Y(n8950) );
  AO22X1 U8281 ( .A0(n5149), .A1(n297), .B0(n5140), .B1(n941), .Y(n8949) );
  AO22X1 U8282 ( .A0(n5121), .A1(n202), .B0(n5114), .B1(n312), .Y(n8353) );
  NOR4X1 U8283 ( .A(n8942), .B(n8941), .C(n8940), .D(n8939), .Y(n8943) );
  AO22X1 U8284 ( .A0(n5123), .A1(n866), .B0(n5119), .B1(n2489), .Y(n8942) );
  AO22X1 U8285 ( .A0(n5136), .A1(n803), .B0(n5129), .B1(n2404), .Y(n8941) );
  AO22X1 U8286 ( .A0(n5149), .A1(n298), .B0(n5140), .B1(n942), .Y(n8940) );
  NOR4X1 U8287 ( .A(n8192), .B(n8191), .C(n8190), .D(n8189), .Y(n8193) );
  AO22X1 U8288 ( .A0(n5123), .A1(n173), .B0(n5119), .B1(n313), .Y(n8192) );
  AO22X1 U8289 ( .A0(n5135), .A1(n279), .B0(n5127), .B1(n924), .Y(n8191) );
  AO22X1 U8290 ( .A0(n5148), .A1(n867), .B0(n5144), .B1(n2490), .Y(n8190) );
  NOR4X1 U8291 ( .A(n8183), .B(n8182), .C(n8181), .D(n8180), .Y(n8184) );
  AO22X1 U8292 ( .A0(n5121), .A1(n203), .B0(n5119), .B1(n314), .Y(n8183) );
  AO22X1 U8293 ( .A0(n5135), .A1(n280), .B0(n5127), .B1(n925), .Y(n8182) );
  AO22X1 U8294 ( .A0(n5148), .A1(n868), .B0(n5144), .B1(n2491), .Y(n8181) );
  NOR4X1 U8295 ( .A(n7471), .B(n7470), .C(n7469), .D(n7468), .Y(n7472) );
  AO22X1 U8296 ( .A0(n5122), .A1(n235), .B0(n5118), .B1(n2492), .Y(n7471) );
  AO22X1 U8297 ( .A0(n5131), .A1(n869), .B0(n5128), .B1(n2493), .Y(n7470) );
  AO22X1 U8298 ( .A0(n5149), .A1(n870), .B0(n5143), .B1(n2494), .Y(n7469) );
  NOR4X1 U8299 ( .A(n7462), .B(n7461), .C(n7460), .D(n7459), .Y(n7463) );
  AO22X1 U8300 ( .A0(n5122), .A1(n871), .B0(n5118), .B1(n2495), .Y(n7462) );
  AO22X1 U8301 ( .A0(n5131), .A1(n872), .B0(n5128), .B1(n2496), .Y(n7461) );
  AO22X1 U8302 ( .A0(n5150), .A1(n873), .B0(n5143), .B1(n2497), .Y(n7460) );
  NOR4X1 U8303 ( .A(n7556), .B(n7555), .C(n7554), .D(n7553), .Y(n7557) );
  AO22X1 U8304 ( .A0(n5122), .A1(n164), .B0(n5118), .B1(n2405), .Y(n7556) );
  AO22X1 U8305 ( .A0(n5131), .A1(n379), .B0(n5128), .B1(n2406), .Y(n7555) );
  AO22X1 U8306 ( .A0(n5150), .A1(n380), .B0(n5143), .B1(n2407), .Y(n7554) );
  NOR4X1 U8307 ( .A(n7547), .B(n7546), .C(n7545), .D(n7544), .Y(n7548) );
  AO22X1 U8308 ( .A0(n5122), .A1(n381), .B0(n5118), .B1(n2408), .Y(n7547) );
  AO22X1 U8309 ( .A0(n5131), .A1(n382), .B0(n5128), .B1(n2409), .Y(n7546) );
  AO22X1 U8310 ( .A0(n5149), .A1(n383), .B0(n5139), .B1(n2410), .Y(n7545) );
  AO22X1 U8311 ( .A0(n5124), .A1(n359), .B0(n5120), .B1(n2498), .Y(n9111) );
  AO22X1 U8312 ( .A0(n5137), .A1(n874), .B0(n5125), .B1(n2499), .Y(n9110) );
  AO22X1 U8313 ( .A0(n5150), .A1(n875), .B0(n5145), .B1(n2500), .Y(n9109) );
  AO22X1 U8314 ( .A0(n5124), .A1(n876), .B0(n5120), .B1(n2501), .Y(n9102) );
  AO22X1 U8315 ( .A0(n5137), .A1(n877), .B0(n5127), .B1(n2502), .Y(n9101) );
  AO22X1 U8316 ( .A0(n5150), .A1(n878), .B0(n5145), .B1(n2503), .Y(n9100) );
  NOR4X1 U8317 ( .A(n8102), .B(n8101), .C(n8100), .D(n8099), .Y(n8103) );
  AO22X1 U8318 ( .A0(n5121), .A1(n165), .B0(n5119), .B1(n251), .Y(n8102) );
  AO22X1 U8319 ( .A0(n5135), .A1(n249), .B0(n5127), .B1(n392), .Y(n8101) );
  AO22X1 U8320 ( .A0(n5148), .A1(n384), .B0(n5144), .B1(n2009), .Y(n8100) );
  NOR4X1 U8321 ( .A(n7372), .B(n7371), .C(n7370), .D(n7369), .Y(n7373) );
  AO22X1 U8322 ( .A0(n5122), .A1(n231), .B0(n5118), .B1(n2504), .Y(n7372) );
  AO22X1 U8323 ( .A0(n5131), .A1(n879), .B0(n5128), .B1(n2505), .Y(n7371) );
  AO22X1 U8324 ( .A0(n5149), .A1(n880), .B0(n5143), .B1(n2506), .Y(n7370) );
  NOR4X1 U8325 ( .A(n8093), .B(n8092), .C(n8091), .D(n8090), .Y(n8094) );
  AO22X1 U8326 ( .A0(n5121), .A1(n180), .B0(n5114), .B1(n252), .Y(n8093) );
  AO22X1 U8327 ( .A0(n5135), .A1(n250), .B0(n5127), .B1(n393), .Y(n8092) );
  AO22X1 U8328 ( .A0(n5148), .A1(n385), .B0(n5144), .B1(n2010), .Y(n8091) );
  AO22X1 U8329 ( .A0(n5135), .A1(n281), .B0(n5125), .B1(n926), .Y(n8018) );
  AO22X1 U8330 ( .A0(n5148), .A1(n804), .B0(n5144), .B1(n2411), .Y(n8017) );
  NOR4X1 U8331 ( .A(n7363), .B(n7362), .C(n7361), .D(n7360), .Y(n7364) );
  AO22X1 U8332 ( .A0(n5122), .A1(n390), .B0(n5118), .B1(n2507), .Y(n7363) );
  AO22X1 U8333 ( .A0(n5131), .A1(n881), .B0(n5128), .B1(n2508), .Y(n7362) );
  AO22X1 U8334 ( .A0(n5150), .A1(n882), .B0(n5143), .B1(n2509), .Y(n7361) );
  AO22X1 U8335 ( .A0(n5121), .A1(n181), .B0(n5114), .B1(n316), .Y(n8010) );
  AO22X1 U8336 ( .A0(n5135), .A1(n282), .B0(n5125), .B1(n927), .Y(n8009) );
  AO22X1 U8337 ( .A0(n5148), .A1(n805), .B0(n5144), .B1(n2412), .Y(n8008) );
  NOR4X1 U8338 ( .A(n7292), .B(n7291), .C(n7290), .D(n7289), .Y(n7293) );
  AO22X1 U8339 ( .A0(n5122), .A1(n232), .B0(n5118), .B1(n2510), .Y(n7292) );
  AO22X1 U8340 ( .A0(n5134), .A1(n883), .B0(n5128), .B1(n2511), .Y(n7291) );
  AO22X1 U8341 ( .A0(n5150), .A1(n884), .B0(n5143), .B1(n2512), .Y(n7290) );
  NOR4X1 U8342 ( .A(n7283), .B(n7282), .C(n7281), .D(n7280), .Y(n7284) );
  AO22X1 U8343 ( .A0(n5122), .A1(n806), .B0(n5118), .B1(n2413), .Y(n7283) );
  AO22X1 U8344 ( .A0(n5131), .A1(n807), .B0(n5128), .B1(n2414), .Y(n7282) );
  AO22X1 U8345 ( .A0(n5150), .A1(n808), .B0(n5143), .B1(n2415), .Y(n7281) );
  NOR4X1 U8346 ( .A(n7642), .B(n7641), .C(n7640), .D(n7639), .Y(n7643) );
  AO22X1 U8347 ( .A0(n5122), .A1(n234), .B0(n5118), .B1(n2416), .Y(n7642) );
  AO22X1 U8348 ( .A0(n5131), .A1(n809), .B0(n5128), .B1(n2417), .Y(n7641) );
  AO22X1 U8349 ( .A0(n5149), .A1(n885), .B0(n5143), .B1(n2513), .Y(n7640) );
  NOR4X1 U8350 ( .A(n7633), .B(n7632), .C(n7631), .D(n7630), .Y(n7634) );
  AO22X1 U8351 ( .A0(n5122), .A1(n386), .B0(n5118), .B1(n2418), .Y(n7633) );
  AO22X1 U8352 ( .A0(n5131), .A1(n810), .B0(n5128), .B1(n2419), .Y(n7632) );
  AO22X1 U8353 ( .A0(n5150), .A1(n886), .B0(n5143), .B1(n2514), .Y(n7631) );
  NOR4X1 U8354 ( .A(n7017), .B(n7016), .C(n7015), .D(n7014), .Y(n7018) );
  AO22X1 U8355 ( .A0(n5124), .A1(n236), .B0(n5117), .B1(n2420), .Y(n7017) );
  AO22X1 U8356 ( .A0(n5134), .A1(n811), .B0(n5127), .B1(n2421), .Y(n7016) );
  AO22X1 U8357 ( .A0(n5147), .A1(n812), .B0(n5143), .B1(n2422), .Y(n7015) );
  NOR4X1 U8358 ( .A(n7008), .B(n7007), .C(n7006), .D(n7005), .Y(n7009) );
  AO22X1 U8359 ( .A0(n5122), .A1(n813), .B0(n5117), .B1(n2423), .Y(n7008) );
  AO22X1 U8360 ( .A0(n5134), .A1(n814), .B0(n5127), .B1(n2424), .Y(n7007) );
  AO22X1 U8361 ( .A0(n5147), .A1(n815), .B0(n5143), .B1(n2425), .Y(n7006) );
  NOR4X1 U8362 ( .A(n7214), .B(n7213), .C(n7212), .D(n7211), .Y(n7215) );
  AO22X1 U8363 ( .A0(n5122), .A1(n237), .B0(n5117), .B1(n2426), .Y(n7214) );
  AO22X1 U8364 ( .A0(n5134), .A1(n816), .B0(n5127), .B1(n2427), .Y(n7213) );
  AO22X1 U8365 ( .A0(n5147), .A1(n887), .B0(n5143), .B1(n2515), .Y(n7212) );
  NOR4X1 U8366 ( .A(n7205), .B(n7204), .C(n7203), .D(n7202), .Y(n7206) );
  AO22X1 U8367 ( .A0(n5124), .A1(n817), .B0(n5117), .B1(n2428), .Y(n7205) );
  AO22X1 U8368 ( .A0(n5134), .A1(n818), .B0(n5127), .B1(n2429), .Y(n7204) );
  AO22X1 U8369 ( .A0(n5147), .A1(n819), .B0(n5143), .B1(n2430), .Y(n7203) );
  NOR4X1 U8370 ( .A(n6906), .B(n6905), .C(n6904), .D(n6903), .Y(n6907) );
  AO22X1 U8371 ( .A0(n5122), .A1(n233), .B0(n5117), .B1(n2431), .Y(n6906) );
  AO22X1 U8372 ( .A0(n5134), .A1(n387), .B0(n5127), .B1(n2432), .Y(n6905) );
  AO22X1 U8373 ( .A0(n5147), .A1(n820), .B0(n5143), .B1(n2433), .Y(n6904) );
  NOR4X1 U8374 ( .A(n6897), .B(n6896), .C(n6895), .D(n6894), .Y(n6898) );
  AO22X1 U8375 ( .A0(n5124), .A1(n388), .B0(n5117), .B1(n2434), .Y(n6897) );
  AO22X1 U8376 ( .A0(n5134), .A1(n389), .B0(n5127), .B1(n2435), .Y(n6896) );
  AO22X1 U8377 ( .A0(n5147), .A1(n821), .B0(n5143), .B1(n2436), .Y(n6895) );
  NOR4X1 U8378 ( .A(n7137), .B(n7136), .C(n7135), .D(n7134), .Y(n7138) );
  AO22X1 U8379 ( .A0(n5124), .A1(n160), .B0(n5117), .B1(n2516), .Y(n7137) );
  AO22X1 U8380 ( .A0(n5134), .A1(n888), .B0(n5127), .B1(n2517), .Y(n7136) );
  AO22X1 U8381 ( .A0(n5147), .A1(n889), .B0(n5143), .B1(n2518), .Y(n7135) );
  NOR4X1 U8382 ( .A(n7128), .B(n7127), .C(n7126), .D(n7125), .Y(n7129) );
  AO22X1 U8383 ( .A0(n5122), .A1(n890), .B0(n5117), .B1(n2519), .Y(n7128) );
  AO22X1 U8384 ( .A0(n5134), .A1(n891), .B0(n5127), .B1(n2520), .Y(n7127) );
  AO22X1 U8385 ( .A0(n5147), .A1(n892), .B0(n5143), .B1(n2521), .Y(n7126) );
  NOR4X1 U8386 ( .A(n6806), .B(n6805), .C(n6804), .D(n6803), .Y(n6807) );
  AO22X1 U8387 ( .A0(n5122), .A1(n238), .B0(n5117), .B1(n2437), .Y(n6806) );
  AO22X1 U8388 ( .A0(n5134), .A1(n822), .B0(n5127), .B1(n2438), .Y(n6805) );
  AO22X1 U8389 ( .A0(n5147), .A1(n893), .B0(n5143), .B1(n2522), .Y(n6804) );
  NOR4X1 U8390 ( .A(n6797), .B(n6796), .C(n6795), .D(n6794), .Y(n6798) );
  AO22X1 U8391 ( .A0(n5122), .A1(n909), .B0(n5117), .B1(n2575), .Y(n6797) );
  AO22X1 U8392 ( .A0(n5134), .A1(n910), .B0(n5127), .B1(n2576), .Y(n6796) );
  AO22X1 U8393 ( .A0(n5147), .A1(n911), .B0(n5143), .B1(n2577), .Y(n6795) );
  NOR4X1 U8394 ( .A(n7829), .B(n7828), .C(n7827), .D(n7826), .Y(n7830) );
  AO22X1 U8395 ( .A0(n5124), .A1(n167), .B0(n5114), .B1(n245), .Y(n7829) );
  AO22X1 U8396 ( .A0(n5135), .A1(n161), .B0(n5125), .B1(n179), .Y(n7828) );
  AO22X1 U8397 ( .A0(n5148), .A1(n163), .B0(n5144), .B1(n178), .Y(n7827) );
  NOR4X1 U8398 ( .A(n7820), .B(n7819), .C(n7818), .D(n7817), .Y(n7821) );
  AO22X1 U8399 ( .A0(n5121), .A1(n177), .B0(n5114), .B1(n246), .Y(n7820) );
  AO22X1 U8400 ( .A0(n5135), .A1(n175), .B0(n5125), .B1(n247), .Y(n7819) );
  AO22X1 U8401 ( .A0(n5148), .A1(n242), .B0(n5144), .B1(n1994), .Y(n7818) );
  NOR4X1 U8402 ( .A(n7732), .B(n7731), .C(n7730), .D(n7729), .Y(n7733) );
  AO22X1 U8403 ( .A0(n5122), .A1(n259), .B0(n5118), .B1(n2439), .Y(n7732) );
  AO22X1 U8404 ( .A0(n5131), .A1(n823), .B0(n5128), .B1(n2440), .Y(n7731) );
  AO22X1 U8405 ( .A0(n5149), .A1(n894), .B0(n5139), .B1(n2523), .Y(n7730) );
  NOR4X1 U8406 ( .A(n7723), .B(n7722), .C(n7721), .D(n7720), .Y(n7724) );
  AO22X1 U8407 ( .A0(n5122), .A1(n824), .B0(n5118), .B1(n2441), .Y(n7723) );
  AO22X1 U8408 ( .A0(n5131), .A1(n825), .B0(n5128), .B1(n2442), .Y(n7722) );
  AO22X1 U8409 ( .A0(n5150), .A1(n826), .B0(n5139), .B1(n2443), .Y(n7721) );
  NOR4X1 U8410 ( .A(n9471), .B(n9470), .C(n9469), .D(n9468), .Y(n9472) );
  AO22X1 U8411 ( .A0(net118341), .A1(n243), .B0(net118321), .B1(n1995), .Y(
        n9471) );
  CLKINVX1 U8412 ( .A(n8385), .Y(n8371) );
  INVX12 U8413 ( .A(n4877), .Y(mem_addr_D[5]) );
  INVX1 U8414 ( .A(n12849), .Y(n4877) );
  NAND2X1 U8415 ( .A(n10712), .B(n10724), .Y(n10720) );
  NAND2X1 U8416 ( .A(n7424), .B(n7399), .Y(n7432) );
  NAND2X1 U8417 ( .A(DCACHE_addr[7]), .B(n5190), .Y(net105008) );
  AOI32XL U8418 ( .A0(n3024), .A1(net108631), .A2(net108632), .B0(n8783), .B1(
        net107404), .Y(n8785) );
  NAND2X1 U8419 ( .A(DCACHE_addr[6]), .B(n5190), .Y(net104939) );
  AOI211XL U8420 ( .A0(n6927), .A1(n9544), .B0(n4794), .C0(n4793), .Y(n6930)
         );
  INVXL U8421 ( .A(n8550), .Y(n8551) );
  INVXL U8422 ( .A(n9303), .Y(n7223) );
  OA22XL U8423 ( .A0(n3670), .A1(n5073), .B0(n959), .B1(n5067), .Y(n7416) );
  MX2XL U8424 ( .A(net118597), .B(net118592), .S0(net108299), .Y(n8982) );
  OAI2BB2XL U8425 ( .B0(n9548), .B1(n9547), .A0N(n9546), .A1N(n4682), .Y(n9561) );
  AOI2BB1XL U8426 ( .A0N(n9545), .A1N(n9544), .B0(n4810), .Y(n9548) );
  NAND2X1 U8427 ( .A(n6666), .B(n6665), .Y(n6683) );
  INVXL U8428 ( .A(n11101), .Y(n11104) );
  AND2XL U8429 ( .A(n7494), .B(n8467), .Y(n7498) );
  NAND2XL U8430 ( .A(net109179), .B(n8648), .Y(n7500) );
  NAND2XL U8431 ( .A(n8382), .B(n8381), .Y(n8393) );
  NAND2XL U8432 ( .A(n8886), .B(n8885), .Y(n8893) );
  NAND2XL U8433 ( .A(n8860), .B(n8859), .Y(n8891) );
  NAND2XL U8434 ( .A(n8550), .B(n8556), .Y(n8569) );
  CLKINVX1 U8435 ( .A(n7686), .Y(n7602) );
  NAND2XL U8436 ( .A(n5075), .B(\i_MIPS/n287 ), .Y(n7299) );
  NAND2X1 U8437 ( .A(n7591), .B(n9425), .Y(n7593) );
  NAND2XL U8438 ( .A(net110131), .B(n7956), .Y(n7963) );
  NAND2XL U8439 ( .A(n9217), .B(n9216), .Y(n9228) );
  NAND2XL U8440 ( .A(n11097), .B(n126), .Y(n7690) );
  NAND2BXL U8441 ( .AN(net108851), .B(net108874), .Y(n7949) );
  NAND2XL U8442 ( .A(n7862), .B(n7861), .Y(n7870) );
  NAND2XL U8443 ( .A(n7024), .B(n7041), .Y(n7047) );
  NAND2XL U8444 ( .A(n3697), .B(n8464), .Y(n8486) );
  NAND2X1 U8445 ( .A(\i_MIPS/n519 ), .B(\i_MIPS/n157 ), .Y(n10903) );
  NAND2X1 U8446 ( .A(\i_MIPS/n506 ), .B(\i_MIPS/n170 ), .Y(n10288) );
  NAND2BXL U8447 ( .AN(net108869), .B(n124), .Y(n8671) );
  CLKMX2X2 U8448 ( .A(n7902), .B(n7901), .S0(net114081), .Y(net110227) );
  NOR4X1 U8449 ( .A(n7883), .B(n7882), .C(n7881), .D(n7880), .Y(n7902) );
  NOR4X1 U8450 ( .A(n7900), .B(n7899), .C(n7898), .D(n7897), .Y(n7901) );
  NAND2XL U8451 ( .A(net110406), .B(net110423), .Y(n7781) );
  NOR4X1 U8452 ( .A(n7929), .B(n7928), .C(n7927), .D(n7926), .Y(n7940) );
  NOR4X1 U8453 ( .A(n7938), .B(n7937), .C(n7936), .D(n7935), .Y(n7939) );
  MX2XL U8454 ( .A(net118597), .B(net118592), .S0(n7670), .Y(n7679) );
  NAND2X1 U8455 ( .A(n7672), .B(n4682), .Y(n7678) );
  NAND2X1 U8456 ( .A(n11026), .B(n3005), .Y(n11514) );
  MX2XL U8457 ( .A(net118597), .B(net118592), .S0(n6828), .Y(n6837) );
  AOI2BB1XL U8458 ( .A0N(n8649), .A1N(n8662), .B0(n4699), .Y(n8672) );
  NAND2XL U8459 ( .A(n3868), .B(n7486), .Y(n7226) );
  CLKINVX1 U8460 ( .A(n7844), .Y(n7409) );
  NAND4X1 U8461 ( .A(n9019), .B(n9018), .C(n9017), .D(n9016), .Y(n11409) );
  OA22X2 U8462 ( .A0(n5390), .A1(n695), .B0(n5432), .B1(n2313), .Y(n8253) );
  OA22X1 U8463 ( .A0(n5251), .A1(n1017), .B0(n5291), .B1(n2643), .Y(n8255) );
  OA22X1 U8464 ( .A0(n5244), .A1(n1018), .B0(n5285), .B1(n2644), .Y(n9179) );
  OA22X1 U8465 ( .A0(n5248), .A1(n1019), .B0(n5288), .B1(n2645), .Y(n8755) );
  OA22X2 U8466 ( .A0(n5386), .A1(n566), .B0(n5427), .B1(n2318), .Y(n9092) );
  OA22X1 U8467 ( .A0(n5249), .A1(n1020), .B0(n5289), .B1(n2646), .Y(n8526) );
  OA22X2 U8468 ( .A0(n5378), .A1(n702), .B0(n5420), .B1(n2322), .Y(n9412) );
  OA22X1 U8469 ( .A0(n5240), .A1(n1021), .B0(n5290), .B1(n2647), .Y(n9414) );
  OA22X1 U8470 ( .A0(n5177), .A1(n1022), .B0(n5216), .B1(n2648), .Y(n9415) );
  OA22X2 U8471 ( .A0(n5389), .A1(n718), .B0(n5436), .B1(n2340), .Y(n8600) );
  OA22X1 U8472 ( .A0(n5237), .A1(n1023), .B0(n5277), .B1(n2649), .Y(n9527) );
  OA22X1 U8473 ( .A0(n5252), .A1(n1024), .B0(n5292), .B1(n2650), .Y(n8175) );
  OA22X1 U8474 ( .A0(n5405), .A1(n1025), .B0(n5433), .B1(n2651), .Y(n8083) );
  OA22X1 U8475 ( .A0(n5252), .A1(n1026), .B0(n5292), .B1(n2652), .Y(n8085) );
  OA22X1 U8476 ( .A0(n5175), .A1(n1027), .B0(n5214), .B1(n2653), .Y(n8086) );
  OA22X1 U8477 ( .A0(n5391), .A1(n1028), .B0(n5434), .B1(n2654), .Y(n8000) );
  OA22X1 U8478 ( .A0(n5253), .A1(n1029), .B0(n5293), .B1(n2655), .Y(n8002) );
  OA22X1 U8479 ( .A0(n5178), .A1(n1030), .B0(n5217), .B1(n2656), .Y(n8003) );
  OA22X1 U8480 ( .A0(n5395), .A1(n1031), .B0(n5439), .B1(n2657), .Y(n7353) );
  OA22X1 U8481 ( .A0(n5266), .A1(n1032), .B0(n5298), .B1(n2658), .Y(n7355) );
  OA22X1 U8482 ( .A0(n5180), .A1(n1033), .B0(n5218), .B1(n2659), .Y(n7356) );
  OA22X1 U8483 ( .A0(n5256), .A1(n1034), .B0(n5285), .B1(n2660), .Y(n9360) );
  OA22X1 U8484 ( .A0(n5177), .A1(n1035), .B0(n5216), .B1(n2661), .Y(n9361) );
  OA22X1 U8485 ( .A0(n5395), .A1(n1036), .B0(n5438), .B1(n2662), .Y(n7448) );
  OA22X1 U8486 ( .A0(n5250), .A1(n1037), .B0(n5297), .B1(n2663), .Y(n7450) );
  OA22X1 U8487 ( .A0(n5395), .A1(n1038), .B0(n5438), .B1(n2664), .Y(n7526) );
  OA22X1 U8488 ( .A0(n5255), .A1(n1039), .B0(n5297), .B1(n2665), .Y(n7528) );
  OA22X1 U8489 ( .A0(n5180), .A1(n1040), .B0(n5218), .B1(n2666), .Y(n7529) );
  OA22X1 U8490 ( .A0(n5245), .A1(n1041), .B0(n5286), .B1(n2667), .Y(n9082) );
  OA22X1 U8491 ( .A0(n5176), .A1(n950), .B0(n5215), .B1(n2668), .Y(n9083) );
  OA22X1 U8492 ( .A0(n5181), .A1(n1042), .B0(n5218), .B1(n2669), .Y(n7200) );
  OA22X1 U8493 ( .A0(n5178), .A1(n1045), .B0(n5217), .B1(n2672), .Y(n8074) );
  OA22X1 U8494 ( .A0(n5253), .A1(n1046), .B0(n5298), .B1(n2673), .Y(n7275) );
  OA22X1 U8495 ( .A0(n5180), .A1(n1047), .B0(n5218), .B1(n2674), .Y(n7276) );
  OA22X1 U8496 ( .A0(n5395), .A1(n1048), .B0(n5439), .B1(n2675), .Y(n7341) );
  OA22X1 U8497 ( .A0(n5253), .A1(n1050), .B0(n5300), .B1(n2677), .Y(n7120) );
  OA22X1 U8498 ( .A0(n5181), .A1(n1051), .B0(n5218), .B1(n2678), .Y(n7121) );
  OA22X1 U8499 ( .A0(n5396), .A1(n1052), .B0(n5440), .B1(n2679), .Y(n7265) );
  OA22X1 U8500 ( .A0(n5392), .A1(n1053), .B0(n5435), .B1(n2680), .Y(n7809) );
  OA22X1 U8501 ( .A0(n5254), .A1(n1054), .B0(n5294), .B1(n2681), .Y(n7811) );
  OA22X1 U8502 ( .A0(n5397), .A1(n1055), .B0(n5441), .B1(n2682), .Y(n7110) );
  OA22X1 U8503 ( .A0(n5250), .A1(n1056), .B0(n5300), .B1(n2683), .Y(n7112) );
  OA22X1 U8504 ( .A0(n5181), .A1(n1057), .B0(n5218), .B1(n2684), .Y(n7113) );
  OA22X1 U8505 ( .A0(n5179), .A1(n1059), .B0(n5213), .B1(n2686), .Y(n7712) );
  OA22XL U8506 ( .A0(n5392), .A1(n1228), .B0(n5435), .B1(n2851), .Y(n7907) );
  OA22XL U8507 ( .A0(n5178), .A1(n1229), .B0(n5217), .B1(n2852), .Y(n7910) );
  OA22X1 U8508 ( .A0(n5396), .A1(n1061), .B0(n5440), .B1(n2688), .Y(n7261) );
  OA22X1 U8509 ( .A0(n5180), .A1(n957), .B0(n5218), .B1(n2689), .Y(n7264) );
  OA22X1 U8510 ( .A0(n5398), .A1(n1062), .B0(n5442), .B1(n2690), .Y(n6973) );
  OA22X1 U8511 ( .A0(n5257), .A1(n1063), .B0(n5309), .B1(n2691), .Y(n6975) );
  OA22X1 U8512 ( .A0(n5181), .A1(n1064), .B0(n5218), .B1(n2692), .Y(n6976) );
  OA22X1 U8513 ( .A0(n5179), .A1(n1066), .B0(n5218), .B1(n2694), .Y(n7808) );
  OA22X1 U8514 ( .A0(n5394), .A1(n1067), .B0(n5437), .B1(n2695), .Y(n7701) );
  OA22X1 U8515 ( .A0(n5179), .A1(n2893), .B0(n5213), .B1(n1230), .Y(n7704) );
  OA22X1 U8516 ( .A0(n5266), .A1(n1068), .B0(n5296), .B1(n2696), .Y(n7703) );
  OA22X1 U8517 ( .A0(n5397), .A1(n1069), .B0(n5441), .B1(n2697), .Y(n7114) );
  OA22X1 U8518 ( .A0(n5251), .A1(n1070), .B0(n5300), .B1(n2698), .Y(n7116) );
  OA22X1 U8519 ( .A0(n5181), .A1(n1071), .B0(n5218), .B1(n2699), .Y(n7117) );
  OA22X1 U8520 ( .A0(n5257), .A1(n1072), .B0(n5301), .B1(n2700), .Y(n6967) );
  OA22XL U8521 ( .A0(n5182), .A1(n1231), .B0(n5219), .B1(n2853), .Y(n6968) );
  OA22X1 U8522 ( .A0(n5257), .A1(n1245), .B0(n5301), .B1(n2865), .Y(n6860) );
  OA22XL U8523 ( .A0(n5182), .A1(n1260), .B0(n5219), .B1(n2880), .Y(n6861) );
  OA22X1 U8524 ( .A0(n5399), .A1(n1073), .B0(n5443), .B1(n2701), .Y(n6862) );
  OA22X1 U8525 ( .A0(n5257), .A1(n1074), .B0(n5301), .B1(n2702), .Y(n6864) );
  OA22XL U8526 ( .A0(n5182), .A1(n1232), .B0(n5219), .B1(n2854), .Y(n6865) );
  NAND4X1 U8527 ( .A(n6746), .B(n6745), .C(n6744), .D(n6743), .Y(n11400) );
  OA22XL U8528 ( .A0(n5258), .A1(n1233), .B0(n5291), .B1(n2855), .Y(n6745) );
  OA22XL U8529 ( .A0(n5182), .A1(n1234), .B0(n5219), .B1(n2856), .Y(n6746) );
  NAND4X1 U8530 ( .A(n6738), .B(n6737), .C(n6736), .D(n6735), .Y(n11496) );
  OA22XL U8531 ( .A0(n5258), .A1(n1261), .B0(n5289), .B1(n2881), .Y(n6737) );
  OA22XL U8532 ( .A0(n5177), .A1(n1262), .B0(n5219), .B1(n2882), .Y(n6738) );
  NAND3BX1 U8533 ( .AN(n10583), .B(n10582), .C(n10581), .Y(n10584) );
  NAND2XL U8534 ( .A(n8124), .B(n8134), .Y(n8125) );
  CLKINVX1 U8535 ( .A(n7431), .Y(n6914) );
  INVXL U8536 ( .A(n3789), .Y(n9796) );
  CLKINVX1 U8537 ( .A(n7680), .Y(n7681) );
  CLKINVX1 U8538 ( .A(n7145), .Y(n9122) );
  NAND2XL U8539 ( .A(n8117), .B(n7314), .Y(n7309) );
  CLKMX2X2 U8540 ( .A(n7002), .B(n7001), .S0(net114085), .Y(n7003) );
  NOR4X1 U8541 ( .A(n6991), .B(n6990), .C(n6989), .D(n6988), .Y(n7002) );
  NAND2X1 U8542 ( .A(DCACHE_addr[16]), .B(\i_MIPS/n266 ), .Y(net104962) );
  NAND2X1 U8543 ( .A(DCACHE_addr[11]), .B(n5190), .Y(net104698) );
  NAND2X1 U8544 ( .A(DCACHE_addr[18]), .B(n5190), .Y(net105334) );
  OA21XL U8545 ( .A0(n8647), .A1(n8646), .B0(n8645), .Y(n8649) );
  NAND2XL U8546 ( .A(n9299), .B(n9298), .Y(n9313) );
  AOI2BB1XL U8547 ( .A0N(n9135), .A1N(n9544), .B0(n4799), .Y(n8973) );
  NAND2XL U8548 ( .A(n9303), .B(net107680), .Y(n9048) );
  CLKINVX1 U8549 ( .A(n9603), .Y(n9601) );
  NAND2XL U8550 ( .A(n8646), .B(n8663), .Y(n8128) );
  INVX1 U8551 ( .A(n9606), .Y(n9607) );
  NAND2XL U8552 ( .A(n9309), .B(n9308), .Y(n9310) );
  CLKINVX1 U8553 ( .A(n7600), .Y(n7601) );
  NAND2XL U8554 ( .A(n3557), .B(n8120), .Y(n7308) );
  NAND2X1 U8555 ( .A(DCACHE_addr[8]), .B(n5190), .Y(net105119) );
  MXI2XL U8556 ( .A(\i_MIPS/n299 ), .B(n2928), .S0(n5050), .Y(n4734) );
  NAND2XL U8557 ( .A(n7301), .B(n3727), .Y(n7229) );
  MX2XL U8558 ( .A(\i_MIPS/n296 ), .B(n1302), .S0(n5050), .Y(n9136) );
  CLKMX2X2 U8559 ( .A(n7098), .B(n7097), .S0(net114087), .Y(n7099) );
  NOR4X1 U8560 ( .A(n7087), .B(n7086), .C(n7085), .D(n7084), .Y(n7098) );
  NOR4X1 U8561 ( .A(n7173), .B(n7172), .C(n7171), .D(n7170), .Y(n7184) );
  CLKMX2X2 U8562 ( .A(n7259), .B(n7258), .S0(net114087), .Y(n7260) );
  NOR4X1 U8563 ( .A(n7248), .B(n7247), .C(n7246), .D(n7245), .Y(n7259) );
  CLKMX2X2 U8564 ( .A(n6791), .B(n6790), .S0(net114087), .Y(n6792) );
  NOR4X1 U8565 ( .A(n7513), .B(n7512), .C(n7511), .D(n7510), .Y(n7524) );
  NOR4X1 U8566 ( .A(n8408), .B(n8407), .C(n8406), .D(n8405), .Y(n8419) );
  NOR4X1 U8567 ( .A(n8907), .B(n8906), .C(n8905), .D(n8904), .Y(n8918) );
  CLKMX2X2 U8568 ( .A(n8740), .B(n8739), .S0(net114085), .Y(net108729) );
  NOR4X1 U8569 ( .A(n8729), .B(n8728), .C(n8727), .D(n8726), .Y(n8740) );
  CLKMX2X2 U8570 ( .A(n7398), .B(n7397), .S0(net114087), .Y(n7439) );
  NOR4X1 U8571 ( .A(n7387), .B(n7386), .C(n7385), .D(n7384), .Y(n7398) );
  CLKMX2X2 U8572 ( .A(n8511), .B(n8510), .S0(net114085), .Y(net109129) );
  NOR4X1 U8573 ( .A(n8500), .B(n8499), .C(n8498), .D(n8497), .Y(n8511) );
  CLKMX2X2 U8574 ( .A(n8330), .B(n8329), .S0(net114085), .Y(net109447) );
  NOR4X1 U8575 ( .A(n8319), .B(n8318), .C(n8317), .D(n8316), .Y(n8330) );
  CLKMX2X2 U8576 ( .A(n7582), .B(n7581), .S0(net114087), .Y(net110729) );
  NOR4X1 U8577 ( .A(n7571), .B(n7570), .C(n7569), .D(n7568), .Y(n7582) );
  CLKMX2X2 U8578 ( .A(n8240), .B(n8239), .S0(net114087), .Y(net109616) );
  NOR4X1 U8579 ( .A(n8229), .B(n8228), .C(n8227), .D(n8226), .Y(n8240) );
  CLKMX2X2 U8580 ( .A(n9003), .B(n9002), .S0(net114085), .Y(net108249) );
  NOR4X1 U8581 ( .A(n8992), .B(n8991), .C(n8990), .D(n8989), .Y(n9003) );
  CLKMX2X2 U8582 ( .A(n8816), .B(n8815), .S0(net114085), .Y(net108579) );
  NOR4X1 U8583 ( .A(n8805), .B(n8804), .C(n8803), .D(n8802), .Y(n8816) );
  CLKMX2X2 U8584 ( .A(n7668), .B(n7667), .S0(net114087), .Y(net110569) );
  NOR4X1 U8585 ( .A(n7657), .B(n7656), .C(n7655), .D(n7654), .Y(n7668) );
  AND2XL U8586 ( .A(n4803), .B(n10319), .Y(n4743) );
  MX2XL U8587 ( .A(n347), .B(n3861), .S0(n5050), .Y(n9446) );
  MX2XL U8588 ( .A(n2961), .B(n347), .S0(n5050), .Y(n9545) );
  AND2X2 U8589 ( .A(\i_MIPS/n517 ), .B(\i_MIPS/n159 ), .Y(n4747) );
  MX2XL U8590 ( .A(n2928), .B(\i_MIPS/n297 ), .S0(n5050), .Y(n9135) );
  AND4XL U8591 ( .A(n8634), .B(n11103), .C(n8633), .D(n8632), .Y(n4751) );
  CLKINVX1 U8592 ( .A(n10110), .Y(n7813) );
  CLKMX2X2 U8593 ( .A(n6812), .B(n6811), .S0(\i_MIPS/jump_addr[22] ), .Y(
        net112118) );
  CLKMX2X2 U8594 ( .A(n8957), .B(n8956), .S0(net114081), .Y(n8960) );
  AO21X1 U8595 ( .A0(\i_MIPS/n506 ), .A1(n10320), .B0(n4749), .Y(n10330) );
  CLKMX2X2 U8596 ( .A(n7835), .B(n7834), .S0(net114081), .Y(n7839) );
  CLKINVX1 U8597 ( .A(n9563), .Y(n9564) );
  AND2XL U8598 ( .A(n8211), .B(n8199), .Y(n8220) );
  AND2XL U8599 ( .A(n8202), .B(n3666), .Y(n8217) );
  INVX1 U8600 ( .A(n10539), .Y(n5499) );
  NAND2XL U8601 ( .A(net105165), .B(net105166), .Y(n10498) );
  MX3XL U8602 ( .A(n9135), .B(n9136), .C(n9137), .S0(n5051), .S1(net114065), 
        .Y(n9140) );
  CLKBUFX3 U8603 ( .A(\i_MIPS/n266 ), .Y(n5190) );
  CLKMX2X2 U8604 ( .A(net107657), .B(net107656), .S0(n4761), .Y(n8708) );
  NAND2XL U8605 ( .A(n3852), .B(\i_MIPS/n301 ), .Y(n4761) );
  MX2XL U8606 ( .A(DCACHE_addr[1]), .B(n3759), .S0(n3599), .Y(\i_MIPS/n396 )
         );
  MX2XL U8607 ( .A(DCACHE_addr[23]), .B(net105290), .S0(n3588), .Y(
        \i_MIPS/n374 ) );
  MX2XL U8608 ( .A(DCACHE_addr[25]), .B(net105425), .S0(n3597), .Y(
        \i_MIPS/n372 ) );
  AND4X2 U8609 ( .A(n9456), .B(net107389), .C(n9455), .D(n9454), .Y(n9457) );
  MX2XL U8610 ( .A(net118597), .B(net118592), .S0(n9449), .Y(n9456) );
  NAND2XL U8611 ( .A(n9450), .B(n4682), .Y(n9455) );
  AO22X1 U8612 ( .A0(n5158), .A1(n372), .B0(n5151), .B1(n1998), .Y(n9507) );
  AO22X1 U8613 ( .A0(n5158), .A1(n176), .B0(n5153), .B1(n2005), .Y(n9490) );
  AO22X1 U8614 ( .A0(net118271), .A1(n370), .B0(net118289), .B1(n1996), .Y(
        n7936) );
  AO22X1 U8615 ( .A0(net118271), .A1(n371), .B0(net118289), .B1(n1997), .Y(
        n7927) );
  AO22X1 U8616 ( .A0(n5098), .A1(n370), .B0(n5102), .B1(n1996), .Y(n7898) );
  AO22X1 U8617 ( .A0(n5098), .A1(n371), .B0(n5102), .B1(n1997), .Y(n7881) );
  MX2XL U8618 ( .A(DCACHE_addr[0]), .B(net104765), .S0(n3605), .Y(
        \i_MIPS/n397 ) );
  OA22XL U8619 ( .A0(n9448), .A1(n3617), .B0(n3617), .B1(n9447), .Y(n9458) );
  AOI2BB1XL U8620 ( .A0N(n9446), .A1N(n9544), .B0(n4798), .Y(n9448) );
  INVXL U8621 ( .A(n7941), .Y(n7948) );
  AO22X1 U8622 ( .A0(n7945), .A1(n7790), .B0(net107652), .B1(n7789), .Y(n7791)
         );
  MX2XL U8623 ( .A(n5055), .B(n3886), .S0(n3590), .Y(\i_MIPS/n393 ) );
  MX2XL U8624 ( .A(DCACHE_addr[2]), .B(n3734), .S0(n3603), .Y(\i_MIPS/n395 )
         );
  CLKINVX1 U8625 ( .A(n10582), .Y(n10580) );
  CLKINVX1 U8626 ( .A(n8662), .Y(n8664) );
  MX2XL U8627 ( .A(DCACHE_addr[28]), .B(n4020), .S0(n3589), .Y(\i_MIPS/n369 )
         );
  AO22XL U8628 ( .A0(n8976), .A1(n8975), .B0(n4735), .B1(net107652), .Y(n8977)
         );
  NOR4X1 U8629 ( .A(n7328), .B(n7327), .C(n7326), .D(n7325), .Y(n7339) );
  AND3XL U8630 ( .A(net111262), .B(n3673), .C(net109965), .Y(n7306) );
  MX2XL U8631 ( .A(DCACHE_addr[19]), .B(n3836), .S0(n3597), .Y(\i_MIPS/n378 )
         );
  MX2XL U8632 ( .A(DCACHE_addr[6]), .B(n3639), .S0(n3595), .Y(\i_MIPS/n391 )
         );
  INVXL U8633 ( .A(n8681), .Y(n8684) );
  OAI221XL U8634 ( .A0(\i_MIPS/n270 ), .A1(net118597), .B0(n9556), .B1(
        net118597), .C0(n9554), .Y(n9559) );
  AO22X1 U8635 ( .A0(DCACHE_addr[28]), .A1(mem_read_D), .B0(mem_write_D), .B1(
        n11532), .Y(n5018) );
  AO22X1 U8636 ( .A0(DCACHE_addr[29]), .A1(mem_read_D), .B0(mem_write_D), .B1(
        n11533), .Y(n5019) );
  INVX1 U8637 ( .A(n7959), .Y(n7773) );
  NAND3BX1 U8638 ( .AN(n11574), .B(\i_MIPS/Control/n10 ), .C(
        \i_MIPS/Control/n14 ), .Y(n9824) );
  CLKBUFX3 U8639 ( .A(n11208), .Y(n5616) );
  CLKBUFX3 U8640 ( .A(n135), .Y(n5662) );
  AO22X1 U8641 ( .A0(net118491), .A1(n372), .B0(net118467), .B1(n1998), .Y(
        n9587) );
  NAND4X1 U8642 ( .A(n9658), .B(n9657), .C(n9656), .D(n9655), .Y(n11342) );
  AO21X2 U8643 ( .A0(\i_MIPS/Register/n104 ), .A1(\i_MIPS/Register/n105 ), 
        .B0(n4837), .Y(n10798) );
  NAND2X1 U8644 ( .A(\i_MIPS/PC/n4 ), .B(\i_MIPS/PC/n5 ), .Y(n9604) );
  NAND2X1 U8645 ( .A(\i_MIPS/Control/n14 ), .B(n11576), .Y(
        \i_MIPS/control_out[7] ) );
  AND2XL U8646 ( .A(n4802), .B(n10279), .Y(n4765) );
  AND2XL U8647 ( .A(n10155), .B(n10156), .Y(n4766) );
  AND2XL U8648 ( .A(n10905), .B(n10904), .Y(n4768) );
  AND2X2 U8649 ( .A(\i_MIPS/n506 ), .B(\i_MIPS/n177 ), .Y(n4769) );
  AOI21XL U8650 ( .A0(n10470), .A1(n10469), .B0(n10468), .Y(n4770) );
  INVX3 U8651 ( .A(n4837), .Y(n5953) );
  INVX3 U8652 ( .A(\i_MIPS/n496 ), .Y(net114085) );
  INVX3 U8653 ( .A(\i_MIPS/n496 ), .Y(net114087) );
  INVX3 U8654 ( .A(n4837), .Y(n5952) );
  AND3XL U8655 ( .A(n10157), .B(n10156), .C(n10155), .Y(n10144) );
  CLKINVX1 U8656 ( .A(\i_MIPS/Control/n10 ), .Y(n11538) );
  CLKINVX1 U8657 ( .A(n10724), .Y(n10728) );
  CLKINVX1 U8658 ( .A(n10157), .Y(n10136) );
  CLKINVX1 U8659 ( .A(n10174), .Y(n10165) );
  CLKINVX1 U8660 ( .A(n10725), .Y(n10712) );
  NAND4BX4 U8661 ( .AN(n4771), .B(n6760), .C(\i_MIPS/ID_EX_0 ), .D(n6759), .Y(
        net107141) );
  MXI2X2 U8662 ( .A(n10706), .B(n10705), .S0(n5549), .Y(n10707) );
  MXI2X2 U8663 ( .A(n10599), .B(n10598), .S0(n5547), .Y(n10600) );
  MXI2X2 U8664 ( .A(n10398), .B(n10397), .S0(n5543), .Y(n10399) );
  MXI2X2 U8665 ( .A(n10205), .B(n10204), .S0(n5543), .Y(n10206) );
  MXI2X2 U8666 ( .A(n10438), .B(n10437), .S0(n5544), .Y(n10439) );
  MXI2X2 U8667 ( .A(n10424), .B(n10423), .S0(n5544), .Y(n10425) );
  AOI222XL U8668 ( .A0(n3800), .A1(n11400), .B0(mem_rdata_D[24]), .B1(n133), 
        .C0(n12989), .C1(n5537), .Y(n10424) );
  MXI2X2 U8669 ( .A(n10693), .B(n10692), .S0(n5549), .Y(n10694) );
  MXI2X2 U8670 ( .A(n10314), .B(n10313), .S0(n5543), .Y(n10315) );
  MXI2X2 U8671 ( .A(n10411), .B(n10410), .S0(n5544), .Y(n10412) );
  AOI222XL U8672 ( .A0(n3800), .A1(n11396), .B0(mem_rdata_D[20]), .B1(n129), 
        .C0(n12993), .C1(n5537), .Y(n10411) );
  MXI2X2 U8673 ( .A(n10641), .B(n10640), .S0(n5547), .Y(n10642) );
  MXI2X2 U8674 ( .A(n10105), .B(n10104), .S0(n5542), .Y(n10106) );
  AOI222XL U8675 ( .A0(n3800), .A1(n11390), .B0(mem_rdata_D[14]), .B1(n130), 
        .C0(n12999), .C1(n5537), .Y(n10105) );
  MXI2X2 U8676 ( .A(n10613), .B(n10612), .S0(n5547), .Y(n10614) );
  MXI2X2 U8677 ( .A(n10654), .B(n10653), .S0(n5548), .Y(n10655) );
  MXI2X2 U8678 ( .A(n10681), .B(n10680), .S0(n5548), .Y(n10682) );
  MXI2X2 U8679 ( .A(n9954), .B(n9953), .S0(n5542), .Y(n9955) );
  AOI222XL U8680 ( .A0(n3800), .A1(n11382), .B0(mem_rdata_D[6]), .B1(n131), 
        .C0(n13007), .C1(n5537), .Y(n9954) );
  MXI2X2 U8681 ( .A(n10193), .B(n10192), .S0(n5543), .Y(n10194) );
  MXI2X2 U8682 ( .A(n10668), .B(n10667), .S0(n5548), .Y(n10669) );
  MXI2X2 U8683 ( .A(n10703), .B(n10702), .S0(n5549), .Y(n10704) );
  MXI2X2 U8684 ( .A(n10596), .B(n10595), .S0(n5546), .Y(n10597) );
  MXI2X2 U8685 ( .A(n10559), .B(n10558), .S0(n5546), .Y(n10560) );
  MXI2X2 U8686 ( .A(n10546), .B(n10545), .S0(n5546), .Y(n10547) );
  MXI2X2 U8687 ( .A(n10395), .B(n10394), .S0(n5543), .Y(n10396) );
  MXI2X2 U8688 ( .A(n10421), .B(n10420), .S0(n5544), .Y(n10422) );
  MXI2X2 U8689 ( .A(n10311), .B(n10310), .S0(n5543), .Y(n10312) );
  MXI2X2 U8690 ( .A(n10638), .B(n10637), .S0(n5547), .Y(n10639) );
  MXI2X2 U8691 ( .A(n10623), .B(n10622), .S0(n5547), .Y(n10624) );
  MXI2X2 U8692 ( .A(n10102), .B(n10101), .S0(n5542), .Y(n10103) );
  MXI2X2 U8693 ( .A(n10460), .B(n10459), .S0(n5545), .Y(n10461) );
  MXI2X2 U8694 ( .A(n10610), .B(n10609), .S0(n5547), .Y(n10611) );
  AOI222XL U8695 ( .A0(n4505), .A1(n11449), .B0(mem_rdata_D[73]), .B1(n131), 
        .C0(n13004), .C1(n5536), .Y(n10610) );
  MXI2X2 U8696 ( .A(n10651), .B(n10650), .S0(n5548), .Y(n10652) );
  MXI2X2 U8697 ( .A(n10593), .B(n10592), .S0(n5546), .Y(n10594) );
  MXI2X2 U8698 ( .A(n10556), .B(n10555), .S0(n5546), .Y(n10557) );
  MXI2X2 U8699 ( .A(n10543), .B(n10542), .S0(n5546), .Y(n10544) );
  AOI222XL U8700 ( .A0(n4535), .A1(n11497), .B0(mem_rdata_D[121]), .B1(n133), 
        .C0(n12988), .C1(n5533), .Y(n10432) );
  AOI222XL U8701 ( .A0(n4535), .A1(n11496), .B0(mem_rdata_D[120]), .B1(n133), 
        .C0(n12989), .C1(n5533), .Y(n10418) );
  MXI2X2 U8702 ( .A(n10308), .B(n10307), .S0(n5543), .Y(n10309) );
  MXI2X2 U8703 ( .A(n10635), .B(n10634), .S0(n5547), .Y(n10636) );
  MXI2X2 U8704 ( .A(n10445), .B(n10444), .S0(n5545), .Y(n10446) );
  MXI2X2 U8705 ( .A(n10457), .B(n10456), .S0(n5545), .Y(n10458) );
  MXI2X2 U8706 ( .A(n10607), .B(n10606), .S0(n5547), .Y(n10608) );
  MXI2X2 U8707 ( .A(n10675), .B(n10674), .S0(n5548), .Y(n10676) );
  AOI222XL U8708 ( .A0(n4535), .A1(n11478), .B0(mem_rdata_D[102]), .B1(n132), 
        .C0(n13007), .C1(n5533), .Y(n9941) );
  AOI222XL U8709 ( .A0(n4535), .A1(n11474), .B0(mem_rdata_D[98]), .B1(n131), 
        .C0(n13011), .C1(n5533), .Y(n10187) );
  MXI2X2 U8710 ( .A(n10401), .B(n10400), .S0(n5544), .Y(n10402) );
  AOI222XL U8711 ( .A0(n5541), .A1(n11435), .B0(mem_rdata_D[59]), .B1(n130), 
        .C0(n12986), .C1(n5539), .Y(n10401) );
  MXI2X2 U8712 ( .A(n10441), .B(n10440), .S0(n5544), .Y(n10442) );
  MXI2X2 U8713 ( .A(n10427), .B(n10426), .S0(n5544), .Y(n10428) );
  AOI222XL U8714 ( .A0(n5541), .A1(n11432), .B0(mem_rdata_D[56]), .B1(n132), 
        .C0(n12989), .C1(n5539), .Y(n10427) );
  MXI2X2 U8715 ( .A(n10317), .B(n10316), .S0(n5543), .Y(n10318) );
  AOI222XL U8716 ( .A0(n5541), .A1(n11428), .B0(mem_rdata_D[52]), .B1(n131), 
        .C0(n12993), .C1(n5539), .Y(n10414) );
  MXI2X2 U8717 ( .A(n10629), .B(n10628), .S0(n5547), .Y(n10630) );
  MXI2X2 U8718 ( .A(n10108), .B(n10107), .S0(n5542), .Y(n10109) );
  AOI222XL U8719 ( .A0(n5541), .A1(n11422), .B0(mem_rdata_D[46]), .B1(n132), 
        .C0(n12999), .C1(n5539), .Y(n10108) );
  MXI2X2 U8720 ( .A(n10616), .B(n10615), .S0(n5547), .Y(n10617) );
  MXI2X2 U8721 ( .A(n10684), .B(n10683), .S0(n5548), .Y(n10685) );
  AOI222XL U8722 ( .A0(n5541), .A1(n11410), .B0(mem_rdata_D[34]), .B1(n133), 
        .C0(n13011), .C1(n5539), .Y(n10196) );
  MXI2X2 U8723 ( .A(n10809), .B(n10808), .S0(n5544), .Y(n10810) );
  MXI2X2 U8724 ( .A(n10794), .B(n10793), .S0(n5550), .Y(n10795) );
  MXI2X2 U8725 ( .A(n10781), .B(n10780), .S0(n5550), .Y(n10782) );
  AOI222XL U8726 ( .A0(n5541), .A1(n11418), .B0(mem_rdata_D[42]), .B1(n132), 
        .C0(n13003), .C1(n5540), .Y(n10781) );
  MXI2X2 U8727 ( .A(n10901), .B(n10900), .S0(n5550), .Y(n10902) );
  AOI222XL U8728 ( .A0(n5541), .A1(n11412), .B0(mem_rdata_D[36]), .B1(n129), 
        .C0(n13009), .C1(n5540), .Y(n10756) );
  MXI2X2 U8729 ( .A(n10748), .B(n10747), .S0(n5549), .Y(n10749) );
  MXI2X2 U8730 ( .A(n10806), .B(n10805), .S0(n5543), .Y(n10807) );
  MXI2X2 U8731 ( .A(n10791), .B(n10790), .S0(n5550), .Y(n10792) );
  MXI2X2 U8732 ( .A(n10898), .B(n10897), .S0(n5548), .Y(n10899) );
  MXI2X2 U8733 ( .A(n10745), .B(n10744), .S0(n5549), .Y(n10746) );
  MXI2X2 U8734 ( .A(n10803), .B(n10802), .S0(n5547), .Y(n10804) );
  AOI222XL U8735 ( .A0(n4506), .A1(n11453), .B0(mem_rdata_D[77]), .B1(n132), 
        .C0(n13000), .C1(n5536), .Y(n10803) );
  MXI2X2 U8736 ( .A(n10775), .B(n10774), .S0(n5550), .Y(n10776) );
  MXI2X2 U8737 ( .A(n10751), .B(n10750), .S0(n5549), .Y(n10752) );
  MXI2X2 U8738 ( .A(n10742), .B(n10741), .S0(n5549), .Y(n10743) );
  MXI2X2 U8739 ( .A(n10785), .B(n10784), .S0(n5550), .Y(n10786) );
  MXI2X2 U8740 ( .A(n10892), .B(n10891), .S0(n5547), .Y(n10893) );
  MXI2X2 U8741 ( .A(n10968), .B(n10967), .S0(n5547), .Y(n10969) );
  MXI2X2 U8742 ( .A(n10964), .B(n10963), .S0(n5548), .Y(n10965) );
  OA22XL U8743 ( .A0(\i_MIPS/ALUin1[5] ), .A1(n5063), .B0(\i_MIPS/ALUin1[4] ), 
        .B1(n5059), .Y(n8679) );
  AOI2BB1XL U8744 ( .A0N(\i_MIPS/ALUin1[12] ), .A1N(n5068), .B0(n4745), .Y(
        n7156) );
  OAI2BB1XL U8745 ( .A0N(mem_ready_I), .A1N(net36572), .B0(n11217), .Y(n10938)
         );
  OA22XL U8746 ( .A0(\i_MIPS/ALUin1[22] ), .A1(n5064), .B0(\i_MIPS/ALUin1[23] ), .B1(n3778), .Y(n7032) );
  NAND2X1 U8747 ( .A(n10568), .B(ICACHE_addr[25]), .Y(n10532) );
  CLKINVX1 U8748 ( .A(n10330), .Y(n10332) );
  CLKINVX1 U8749 ( .A(n10361), .Y(n10363) );
  OAI222XL U8750 ( .A0(n5532), .A1(n234), .B0(n5499), .B1(n5530), .C0(n5952), 
        .C1(n10540), .Y(n11544) );
  CLKINVX1 U8751 ( .A(\i_MIPS/jump_addr[28] ), .Y(n10540) );
  OAI222XL U8752 ( .A0(n5532), .A1(n259), .B0(n1937), .B1(n5529), .C0(n5953), 
        .C1(\i_MIPS/n180 ), .Y(n11545) );
  OAI222XL U8753 ( .A0(n10798), .A1(n235), .B0(n156), .B1(n5529), .C0(n5953), 
        .C1(\i_MIPS/n179 ), .Y(n11546) );
  OAI222XL U8754 ( .A0(n5531), .A1(n236), .B0(n1933), .B1(n5528), .C0(n5952), 
        .C1(\i_MIPS/n176 ), .Y(n11549) );
  OAI222XL U8755 ( .A0(n5532), .A1(n3546), .B0(n1935), .B1(n5529), .C0(n5953), 
        .C1(n10351), .Y(n11550) );
  OAI222XL U8756 ( .A0(n10798), .A1(n356), .B0(n5475), .B1(n5529), .C0(n5953), 
        .C1(\i_MIPS/n173 ), .Y(n11552) );
  OAI222XL U8757 ( .A0(n5532), .A1(n237), .B0(n1934), .B1(n5529), .C0(n5953), 
        .C1(\i_MIPS/n155 ), .Y(n11570) );
  OAI222XL U8758 ( .A0(n10798), .A1(n238), .B0(n2896), .B1(n5529), .C0(n5953), 
        .C1(\i_MIPS/n178 ), .Y(n11547) );
  OAI222XL U8759 ( .A0(n5531), .A1(n222), .B0(n4982), .B1(n5528), .C0(n5952), 
        .C1(n10734), .Y(n11541) );
  CLKINVX1 U8760 ( .A(\i_MIPS/jump_addr[31] ), .Y(n10734) );
  AO22X2 U8761 ( .A0(n5554), .A1(DCACHE_addr[5]), .B0(n5551), .B1(n11509), .Y(
        n10995) );
  AO22X2 U8762 ( .A0(n5937), .A1(ICACHE_addr[9]), .B0(n5931), .B1(n11351), .Y(
        n11118) );
  AO22X2 U8763 ( .A0(mem_rdata_I[127]), .A1(n5943), .B0(n5573), .B1(n11342), 
        .Y(n9659) );
  AO22X2 U8764 ( .A0(n6562), .A1(n11373), .B0(n4719), .B1(n10979), .Y(n10770)
         );
  NAND2XL U8765 ( .A(mem_ready_D), .B(n10980), .Y(n6562) );
  AO22X2 U8766 ( .A0(mem_rdata_I[31]), .A1(n5944), .B0(n5570), .B1(n11249), 
        .Y(n6587) );
  AO22X2 U8767 ( .A0(mem_rdata_I[30]), .A1(n5943), .B0(n5570), .B1(n11248), 
        .Y(n9676) );
  AO22X2 U8768 ( .A0(mem_rdata_I[29]), .A1(n5943), .B0(n5570), .B1(n11247), 
        .Y(n9698) );
  AO22X2 U8769 ( .A0(mem_rdata_I[28]), .A1(n5943), .B0(n5570), .B1(n11246), 
        .Y(n9646) );
  AO22X2 U8770 ( .A0(mem_rdata_I[27]), .A1(n5944), .B0(n5570), .B1(n11245), 
        .Y(n9624) );
  AO22X2 U8771 ( .A0(mem_rdata_I[26]), .A1(n5944), .B0(n5570), .B1(n11244), 
        .Y(n6602) );
  AO22X2 U8772 ( .A0(mem_rdata_I[25]), .A1(n5940), .B0(n5571), .B1(n11243), 
        .Y(n10043) );
  AO22X2 U8773 ( .A0(mem_rdata_I[24]), .A1(n5939), .B0(n11085), .B1(n11242), 
        .Y(n10838) );
  AO22X2 U8774 ( .A0(mem_rdata_I[23]), .A1(n5940), .B0(n5571), .B1(n11241), 
        .Y(n10021) );
  AO22X2 U8775 ( .A0(mem_rdata_I[22]), .A1(n5944), .B0(n5571), .B1(n11240), 
        .Y(n9977) );
  AO22X2 U8776 ( .A0(mem_rdata_I[20]), .A1(n5941), .B0(n5570), .B1(n11238), 
        .Y(n9788) );
  AO22X2 U8777 ( .A0(mem_rdata_I[19]), .A1(n5944), .B0(n11085), .B1(n11237), 
        .Y(n11086) );
  AO22X2 U8778 ( .A0(mem_rdata_I[18]), .A1(n5942), .B0(n5570), .B1(net103849), 
        .Y(n9772) );
  AO22X2 U8779 ( .A0(mem_rdata_I[16]), .A1(n5942), .B0(n5570), .B1(n11235), 
        .Y(n9762) );
  AO22X2 U8780 ( .A0(mem_rdata_I[14]), .A1(n5939), .B0(n11085), .B1(n11233), 
        .Y(n10246) );
  AO22X2 U8781 ( .A0(mem_rdata_I[13]), .A1(n5940), .B0(n5571), .B1(n11232), 
        .Y(n10224) );
  AO22X2 U8782 ( .A0(mem_rdata_I[12]), .A1(n5940), .B0(n5571), .B1(n11231), 
        .Y(n10126) );
  AO22X2 U8783 ( .A0(mem_rdata_I[11]), .A1(n5940), .B0(n5571), .B1(n11230), 
        .Y(n10090) );
  AO22X2 U8784 ( .A0(mem_rdata_I[10]), .A1(n5941), .B0(n5570), .B1(n11229), 
        .Y(n9839) );
  AO22X2 U8785 ( .A0(mem_rdata_I[9]), .A1(n5933), .B0(n5571), .B1(n11228), .Y(
        n9883) );
  AO22X2 U8786 ( .A0(mem_rdata_I[8]), .A1(n5941), .B0(n5571), .B1(n11227), .Y(
        n9861) );
  AO22X2 U8787 ( .A0(mem_rdata_I[7]), .A1(n5933), .B0(n5571), .B1(n11226), .Y(
        n9905) );
  AO22X2 U8788 ( .A0(mem_rdata_I[6]), .A1(n5941), .B0(n5571), .B1(n11225), .Y(
        n9927) );
  AO22X2 U8789 ( .A0(mem_rdata_I[4]), .A1(n5939), .B0(n11085), .B1(n11223), 
        .Y(n10860) );
  AO22X2 U8790 ( .A0(mem_rdata_I[3]), .A1(n5941), .B0(n11085), .B1(n11222), 
        .Y(n10954) );
  AO22X2 U8791 ( .A0(mem_rdata_I[2]), .A1(n5941), .B0(n11085), .B1(n11221), 
        .Y(n10925) );
  AO22X2 U8792 ( .A0(mem_rdata_I[1]), .A1(n5939), .B0(n11085), .B1(n11220), 
        .Y(n10883) );
  AO22X2 U8793 ( .A0(mem_rdata_I[0]), .A1(n5939), .B0(n11085), .B1(n11219), 
        .Y(n10817) );
  AO22X2 U8794 ( .A0(n4757), .A1(n12956), .B0(n5552), .B1(n11531), .Y(n11022)
         );
  AO22X2 U8795 ( .A0(n4757), .A1(n12961), .B0(n5552), .B1(n11526), .Y(n11019)
         );
  AO22X2 U8796 ( .A0(n5939), .A1(ICACHE_addr[18]), .B0(n5930), .B1(n11360), 
        .Y(n11206) );
  AO22X2 U8797 ( .A0(n5937), .A1(ICACHE_addr[13]), .B0(n5930), .B1(n11355), 
        .Y(n11182) );
  AO22X2 U8798 ( .A0(n5939), .A1(ICACHE_addr[5]), .B0(n5931), .B1(n11347), .Y(
        n11067) );
  AO22X2 U8799 ( .A0(mem_rdata_I[126]), .A1(n5943), .B0(n5573), .B1(n11341), 
        .Y(n9681) );
  AO22X2 U8800 ( .A0(mem_rdata_I[125]), .A1(n5943), .B0(n5573), .B1(n11340), 
        .Y(n9703) );
  AO22X2 U8801 ( .A0(mem_rdata_I[124]), .A1(n5943), .B0(n5573), .B1(n11339), 
        .Y(n9651) );
  AO22X2 U8802 ( .A0(mem_rdata_I[122]), .A1(n5944), .B0(n5573), .B1(n11337), 
        .Y(n6607) );
  AO22X2 U8803 ( .A0(mem_rdata_I[121]), .A1(n5940), .B0(n5572), .B1(n11336), 
        .Y(n10048) );
  AO22X2 U8804 ( .A0(mem_rdata_I[120]), .A1(n5939), .B0(n5573), .B1(n11335), 
        .Y(n10843) );
  AO22X2 U8805 ( .A0(mem_rdata_I[119]), .A1(n5940), .B0(n5572), .B1(n11334), 
        .Y(n10026) );
  AO22X2 U8806 ( .A0(mem_rdata_I[118]), .A1(n5944), .B0(n5572), .B1(n11333), 
        .Y(n9982) );
  AO22X2 U8807 ( .A0(mem_rdata_I[117]), .A1(n5944), .B0(n5572), .B1(n11332), 
        .Y(n10004) );
  AO22X2 U8808 ( .A0(mem_rdata_I[116]), .A1(n5941), .B0(n5573), .B1(n11331), 
        .Y(n9793) );
  AO22X2 U8809 ( .A0(mem_rdata_I[115]), .A1(n5944), .B0(n5573), .B1(n11330), 
        .Y(n11092) );
  AO22X2 U8810 ( .A0(mem_rdata_I[114]), .A1(n5941), .B0(n5573), .B1(net103753), 
        .Y(n9773) );
  AO22X2 U8811 ( .A0(mem_rdata_I[113]), .A1(n5942), .B0(n5573), .B1(n11329), 
        .Y(n9745) );
  AO22X2 U8812 ( .A0(mem_rdata_I[112]), .A1(n5942), .B0(n5573), .B1(n11328), 
        .Y(n9767) );
  AO22X2 U8813 ( .A0(mem_rdata_I[111]), .A1(n5940), .B0(n5572), .B1(n11327), 
        .Y(n10072) );
  AO22X2 U8814 ( .A0(mem_rdata_I[110]), .A1(n5939), .B0(n5573), .B1(n11326), 
        .Y(n10251) );
  AO22X2 U8815 ( .A0(mem_rdata_I[109]), .A1(n5940), .B0(n5572), .B1(n11325), 
        .Y(n10229) );
  AO22X2 U8816 ( .A0(mem_rdata_I[108]), .A1(n5940), .B0(n5572), .B1(n11324), 
        .Y(n10131) );
  AO22X2 U8817 ( .A0(mem_rdata_I[107]), .A1(n5940), .B0(n5572), .B1(n11323), 
        .Y(n10095) );
  AO22X2 U8818 ( .A0(mem_rdata_I[106]), .A1(n5941), .B0(n5573), .B1(n11322), 
        .Y(n9844) );
  AO22X2 U8819 ( .A0(mem_rdata_I[105]), .A1(n5933), .B0(n5572), .B1(n11321), 
        .Y(n9888) );
  AO22X2 U8820 ( .A0(mem_rdata_I[104]), .A1(n5933), .B0(n5572), .B1(n11320), 
        .Y(n9866) );
  AO22X2 U8821 ( .A0(mem_rdata_I[102]), .A1(n5944), .B0(n5572), .B1(n11318), 
        .Y(n9932) );
  AO22X2 U8822 ( .A0(mem_rdata_I[101]), .A1(n5942), .B0(n5573), .B1(n11317), 
        .Y(n9725) );
  AO22X2 U8823 ( .A0(mem_rdata_I[100]), .A1(n5939), .B0(n5573), .B1(n11316), 
        .Y(n10865) );
  AO22X2 U8824 ( .A0(mem_rdata_I[98]), .A1(n5941), .B0(n5573), .B1(n11314), 
        .Y(n10930) );
  AO22X2 U8825 ( .A0(mem_rdata_I[97]), .A1(n5939), .B0(n5573), .B1(n11313), 
        .Y(n10888) );
  AO22X2 U8826 ( .A0(mem_rdata_I[96]), .A1(n5939), .B0(n5573), .B1(n11312), 
        .Y(n10822) );
  AO22X2 U8827 ( .A0(n5936), .A1(ICACHE_addr[25]), .B0(n5930), .B1(n11367), 
        .Y(n11197) );
  AO22X2 U8828 ( .A0(n5554), .A1(n12969), .B0(n5551), .B1(n11518), .Y(n11010)
         );
  AO22X2 U8829 ( .A0(n4757), .A1(n12973), .B0(n5552), .B1(n11514), .Y(n11027)
         );
  AO22X2 U8830 ( .A0(n4757), .A1(n12974), .B0(n5552), .B1(n11513), .Y(n11016)
         );
  AO22X2 U8831 ( .A0(n5554), .A1(n12970), .B0(n5551), .B1(n11517), .Y(n10998)
         );
  AO22X2 U8832 ( .A0(n5554), .A1(n12971), .B0(n5551), .B1(n11516), .Y(n11008)
         );
  AO22X2 U8833 ( .A0(n5554), .A1(n12966), .B0(n5551), .B1(n11521), .Y(n10983)
         );
  OAI221XL U8834 ( .A0(\i_MIPS/Register/register[2][6] ), .A1(net117635), .B0(
        \i_MIPS/Register/register[10][6] ), .B1(net117655), .C0(n7244), .Y(
        n7247) );
  OA22X1 U8835 ( .A0(\i_MIPS/Register/register[6][6] ), .A1(net117673), .B0(
        \i_MIPS/Register/register[14][6] ), .B1(net117691), .Y(n7244) );
  OAI221XL U8836 ( .A0(\i_MIPS/Register/register[2][7] ), .A1(net117637), .B0(
        \i_MIPS/Register/register[10][7] ), .B1(net117655), .C0(n7324), .Y(
        n7327) );
  OAI221XL U8837 ( .A0(\i_MIPS/Register/register[2][23] ), .A1(net117635), 
        .B0(\i_MIPS/Register/register[10][23] ), .B1(net117653), .C0(n7083), 
        .Y(n7086) );
  OA22X1 U8838 ( .A0(\i_MIPS/Register/register[6][23] ), .A1(net117673), .B0(
        \i_MIPS/Register/register[14][23] ), .B1(net117691), .Y(n7083) );
  OAI221XL U8839 ( .A0(\i_MIPS/Register/register[2][10] ), .A1(net117637), 
        .B0(\i_MIPS/Register/register[10][10] ), .B1(net117655), .C0(n7509), 
        .Y(n7512) );
  OA22X1 U8840 ( .A0(\i_MIPS/Register/register[6][10] ), .A1(net117675), .B0(
        \i_MIPS/Register/register[14][10] ), .B1(net117697), .Y(n7509) );
  OAI221XL U8841 ( .A0(\i_MIPS/Register/register[2][26] ), .A1(net117637), 
        .B0(\i_MIPS/Register/register[10][26] ), .B1(net117655), .C0(n7383), 
        .Y(n7386) );
  OAI221XL U8842 ( .A0(\i_MIPS/Register/register[2][11] ), .A1(net117641), 
        .B0(\i_MIPS/Register/register[10][11] ), .B1(net117659), .C0(n8496), 
        .Y(n8499) );
  OAI221XL U8843 ( .A0(\i_MIPS/Register/register[2][19] ), .A1(net117639), 
        .B0(\i_MIPS/Register/register[10][19] ), .B1(net117659), .C0(n8315), 
        .Y(n8318) );
  OAI221XL U8844 ( .A0(\i_MIPS/Register/register[2][13] ), .A1(net117639), 
        .B0(\i_MIPS/Register/register[10][13] ), .B1(net117657), .C0(n7972), 
        .Y(n7975) );
  OA22X1 U8845 ( .A0(\i_MIPS/Register/register[6][13] ), .A1(net117675), .B0(
        \i_MIPS/Register/register[14][13] ), .B1(net117695), .Y(n7972) );
  OAI221XL U8846 ( .A0(\i_MIPS/Register/register[2][12] ), .A1(net117639), 
        .B0(\i_MIPS/Register/register[10][12] ), .B1(net117657), .C0(n8225), 
        .Y(n8228) );
  OAI221XL U8847 ( .A0(\i_MIPS/Register/register[2][17] ), .A1(net117643), 
        .B0(\i_MIPS/Register/register[10][17] ), .B1(net117661), .C0(n9239), 
        .Y(n9242) );
  OAI221XL U8848 ( .A0(\i_MIPS/Register/register[2][5] ), .A1(net117643), .B0(
        \i_MIPS/Register/register[10][5] ), .B1(net117661), .C0(n9330), .Y(
        n9333) );
  OA22X1 U8849 ( .A0(\i_MIPS/Register/register[6][5] ), .A1(net117681), .B0(
        \i_MIPS/Register/register[14][5] ), .B1(net117703), .Y(n9330) );
  OAI221XL U8850 ( .A0(\i_MIPS/Register/register[2][21] ), .A1(net117641), 
        .B0(\i_MIPS/Register/register[10][21] ), .B1(net117661), .C0(n8903), 
        .Y(n8906) );
  OA22X1 U8851 ( .A0(\i_MIPS/Register/register[6][0] ), .A1(net117681), .B0(
        \i_MIPS/Register/register[14][0] ), .B1(net117697), .Y(n8725) );
  OAI221XL U8852 ( .A0(\i_MIPS/Register/register[2][1] ), .A1(net117641), .B0(
        \i_MIPS/Register/register[10][1] ), .B1(net117661), .C0(n8988), .Y(
        n8991) );
  OAI221XL U8853 ( .A0(\i_MIPS/Register/register[2][16] ), .A1(net117641), 
        .B0(\i_MIPS/Register/register[10][16] ), .B1(net117659), .C0(n8801), 
        .Y(n8804) );
  OA22X1 U8854 ( .A0(\i_MIPS/Register/register[6][16] ), .A1(net117685), .B0(
        \i_MIPS/Register/register[14][16] ), .B1(net117697), .Y(n8801) );
  OAI221XL U8855 ( .A0(\i_MIPS/Register/register[2][28] ), .A1(net117637), 
        .B0(\i_MIPS/Register/register[10][28] ), .B1(net117655), .C0(n7567), 
        .Y(n7570) );
  OAI221XL U8856 ( .A0(\i_MIPS/Register/register[2][27] ), .A1(net117637), 
        .B0(\i_MIPS/Register/register[10][27] ), .B1(net117655), .C0(n7653), 
        .Y(n7656) );
  OAI221XL U8857 ( .A0(\i_MIPS/Register/register[2][29] ), .A1(net117635), 
        .B0(\i_MIPS/Register/register[10][29] ), .B1(net117653), .C0(n6987), 
        .Y(n6990) );
  OA22X1 U8858 ( .A0(\i_MIPS/Register/register[6][29] ), .A1(net117673), .B0(
        \i_MIPS/Register/register[14][29] ), .B1(net117691), .Y(n6987) );
  OAI221XL U8859 ( .A0(\i_MIPS/Register/register[2][24] ), .A1(net117635), 
        .B0(\i_MIPS/Register/register[10][24] ), .B1(net117653), .C0(n6775), 
        .Y(n6779) );
  OAI221XL U8860 ( .A0(\i_MIPS/Register/register[2][2] ), .A1(net117635), .B0(
        \i_MIPS/Register/register[10][2] ), .B1(net117653), .C0(n7169), .Y(
        n7172) );
  OAI221XL U8861 ( .A0(\i_MIPS/Register/register[2][22] ), .A1(net117639), 
        .B0(\i_MIPS/Register/register[10][22] ), .B1(net117657), .C0(n7925), 
        .Y(n7928) );
  XOR2XL U8862 ( .A(\i_MIPS/Reg_W[0] ), .B(\i_MIPS/jump_addr[23] ), .Y(n6763)
         );
  XOR2XL U8863 ( .A(\i_MIPS/Reg_W[1] ), .B(n254), .Y(n6762) );
  XOR2XL U8864 ( .A(\i_MIPS/Reg_W[2] ), .B(n11053), .Y(n6761) );
  XOR2X1 U8865 ( .A(\i_MIPS/jump_addr[22] ), .B(n10846), .Y(n6637) );
  XOR2X1 U8866 ( .A(n11053), .B(n10849), .Y(n6758) );
  CLKINVX1 U8867 ( .A(\i_MIPS/n188 ), .Y(n10541) );
  OAI221XL U8868 ( .A0(\i_MIPS/Register/register[18][4] ), .A1(net117643), 
        .B0(\i_MIPS/Register/register[26][4] ), .B1(net117661), .C0(n9072), 
        .Y(n9075) );
  NAND4X1 U8869 ( .A(n9071), .B(n9070), .C(n9069), .D(n9068), .Y(n9076) );
  AO22X1 U8870 ( .A0(net118275), .A1(n283), .B0(net118291), .B1(n2444), .Y(
        n9074) );
  NOR4X1 U8871 ( .A(n8916), .B(n8915), .C(n8914), .D(n8913), .Y(n8917) );
  OAI221XL U8872 ( .A0(\i_MIPS/Register/register[18][21] ), .A1(net117641), 
        .B0(\i_MIPS/Register/register[26][21] ), .B1(net117661), .C0(n8912), 
        .Y(n8915) );
  NAND4X1 U8873 ( .A(n8911), .B(n8910), .C(n8909), .D(n8908), .Y(n8916) );
  AO22X1 U8874 ( .A0(net118275), .A1(n262), .B0(net118291), .B1(n2348), .Y(
        n9250) );
  AO22X1 U8875 ( .A0(net118275), .A1(n266), .B0(net118291), .B1(n2357), .Y(
        n9160) );
  NOR4X1 U8876 ( .A(n8509), .B(n8508), .C(n8507), .D(n8506), .Y(n8510) );
  OAI221XL U8877 ( .A0(\i_MIPS/Register/register[18][11] ), .A1(net117641), 
        .B0(\i_MIPS/Register/register[26][11] ), .B1(net117659), .C0(n8505), 
        .Y(n8508) );
  NAND4X1 U8878 ( .A(n8504), .B(n8503), .C(n8502), .D(n8501), .Y(n8509) );
  AO22X1 U8879 ( .A0(net118273), .A1(n827), .B0(net118291), .B1(n2445), .Y(
        n8507) );
  NOR4X1 U8880 ( .A(n8417), .B(n8416), .C(n8415), .D(n8414), .Y(n8418) );
  NAND4X1 U8881 ( .A(n8412), .B(n8411), .C(n8410), .D(n8409), .Y(n8417) );
  AO22X1 U8882 ( .A0(net118273), .A1(n895), .B0(net118291), .B1(n2524), .Y(
        n8415) );
  NOR4X1 U8883 ( .A(n8328), .B(n8327), .C(n8326), .D(n8325), .Y(n8329) );
  NAND4X1 U8884 ( .A(n8323), .B(n8322), .C(n8321), .D(n8320), .Y(n8328) );
  AO22X1 U8885 ( .A0(net118271), .A1(n828), .B0(net118289), .B1(n2446), .Y(
        n8326) );
  OAI221XL U8886 ( .A0(\i_MIPS/Register/register[18][5] ), .A1(net117643), 
        .B0(\i_MIPS/Register/register[26][5] ), .B1(net117661), .C0(n9339), 
        .Y(n9342) );
  NAND4X1 U8887 ( .A(n9338), .B(n9337), .C(n9336), .D(n9335), .Y(n9343) );
  AO22X1 U8888 ( .A0(net118275), .A1(n263), .B0(net118291), .B1(n2349), .Y(
        n9341) );
  NOR4X1 U8889 ( .A(n8814), .B(n8813), .C(n8812), .D(n8811), .Y(n8815) );
  NAND4X1 U8890 ( .A(n8809), .B(n8808), .C(n8807), .D(n8806), .Y(n8814) );
  AO22X1 U8891 ( .A0(net118273), .A1(n829), .B0(net118291), .B1(n2447), .Y(
        n8812) );
  NOR4X1 U8892 ( .A(n8738), .B(n8737), .C(n8736), .D(n8735), .Y(n8739) );
  NAND4X1 U8893 ( .A(n8733), .B(n8732), .C(n8731), .D(n8730), .Y(n8738) );
  AO22X1 U8894 ( .A0(net118273), .A1(n830), .B0(net118291), .B1(n2448), .Y(
        n8736) );
  NOR4X1 U8895 ( .A(n7096), .B(n7095), .C(n7094), .D(n7093), .Y(n7097) );
  NAND4X1 U8896 ( .A(n7091), .B(n7090), .C(n7089), .D(n7088), .Y(n7096) );
  AO22X1 U8897 ( .A0(net118267), .A1(n284), .B0(net118295), .B1(n928), .Y(
        n7094) );
  NOR4X1 U8898 ( .A(n8238), .B(n8237), .C(n8236), .D(n8235), .Y(n8239) );
  NAND4X1 U8899 ( .A(n8233), .B(n8232), .C(n8231), .D(n8230), .Y(n8238) );
  AO22X1 U8900 ( .A0(net118271), .A1(n831), .B0(net118289), .B1(n2449), .Y(
        n8236) );
  NAND4X1 U8901 ( .A(n8996), .B(n8995), .C(n8994), .D(n8993), .Y(n9001) );
  AO22X1 U8902 ( .A0(net118275), .A1(n285), .B0(net118291), .B1(n2450), .Y(
        n8999) );
  NOR4X1 U8903 ( .A(n8158), .B(n8157), .C(n8156), .D(n8155), .Y(n8159) );
  OAI221XL U8904 ( .A0(\i_MIPS/Register/register[18][8] ), .A1(net117639), 
        .B0(\i_MIPS/Register/register[26][8] ), .B1(net117657), .C0(n8154), 
        .Y(n8157) );
  NAND4X1 U8905 ( .A(n8153), .B(n8152), .C(n8151), .D(n8150), .Y(n8158) );
  AO22X1 U8906 ( .A0(net118271), .A1(n832), .B0(net118289), .B1(n2451), .Y(
        n8156) );
  NOR4X1 U8907 ( .A(n7337), .B(n7336), .C(n7335), .D(n7334), .Y(n7338) );
  OAI221XL U8908 ( .A0(\i_MIPS/Register/register[18][7] ), .A1(net117637), 
        .B0(\i_MIPS/Register/register[26][7] ), .B1(net117655), .C0(n7333), 
        .Y(n7336) );
  NAND4X1 U8909 ( .A(n7332), .B(n7331), .C(n7330), .D(n7329), .Y(n7337) );
  AO22X1 U8910 ( .A0(net118269), .A1(n896), .B0(net118295), .B1(n2525), .Y(
        n7335) );
  NOR4X1 U8911 ( .A(n7522), .B(n7521), .C(n7520), .D(n7519), .Y(n7523) );
  NAND4X1 U8912 ( .A(n7517), .B(n7516), .C(n7515), .D(n7514), .Y(n7522) );
  AO22X1 U8913 ( .A0(net118269), .A1(n723), .B0(net118295), .B1(n2345), .Y(
        n7520) );
  NOR4X1 U8914 ( .A(n7257), .B(n7256), .C(n7255), .D(n7254), .Y(n7258) );
  OAI221XL U8915 ( .A0(\i_MIPS/Register/register[18][6] ), .A1(net117637), 
        .B0(\i_MIPS/Register/register[26][6] ), .B1(net117655), .C0(n7253), 
        .Y(n7256) );
  NAND4X1 U8916 ( .A(n7252), .B(n7251), .C(n7250), .D(n7249), .Y(n7257) );
  AO22X1 U8917 ( .A0(net118269), .A1(n897), .B0(net118295), .B1(n2526), .Y(
        n7255) );
  NOR4X1 U8918 ( .A(n7396), .B(n7395), .C(n7394), .D(n7393), .Y(n7397) );
  OAI221XL U8919 ( .A0(\i_MIPS/Register/register[18][26] ), .A1(net117637), 
        .B0(\i_MIPS/Register/register[26][26] ), .B1(net117655), .C0(n7392), 
        .Y(n7395) );
  NAND4X1 U8920 ( .A(n7391), .B(n7390), .C(n7389), .D(n7388), .Y(n7396) );
  AO22X1 U8921 ( .A0(net118269), .A1(n898), .B0(net118295), .B1(n2527), .Y(
        n7394) );
  NOR4X1 U8922 ( .A(n7000), .B(n6999), .C(n6998), .D(n6997), .Y(n7001) );
  NAND4X1 U8923 ( .A(n6995), .B(n6994), .C(n6993), .D(n6992), .Y(n7000) );
  AO22X1 U8924 ( .A0(net118267), .A1(n286), .B0(net118295), .B1(n929), .Y(
        n6998) );
  NAND4X1 U8925 ( .A(n8062), .B(n8061), .C(n8060), .D(n8059), .Y(n8067) );
  NAND4X1 U8926 ( .A(n7980), .B(n7979), .C(n7978), .D(n7977), .Y(n7985) );
  NOR4X1 U8927 ( .A(n7182), .B(n7181), .C(n7180), .D(n7179), .Y(n7183) );
  OAI221XL U8928 ( .A0(\i_MIPS/Register/register[18][2] ), .A1(net117635), 
        .B0(\i_MIPS/Register/register[26][2] ), .B1(net117653), .C0(n7178), 
        .Y(n7181) );
  NAND4X1 U8929 ( .A(n7177), .B(n7176), .C(n7175), .D(n7174), .Y(n7182) );
  AO22X1 U8930 ( .A0(net118267), .A1(n287), .B0(net118295), .B1(n930), .Y(
        n7180) );
  NOR4X1 U8931 ( .A(n7666), .B(n7665), .C(n7664), .D(n7663), .Y(n7667) );
  OAI221XL U8932 ( .A0(\i_MIPS/Register/register[18][27] ), .A1(net117637), 
        .B0(\i_MIPS/Register/register[26][27] ), .B1(net117655), .C0(n7662), 
        .Y(n7665) );
  NAND4X1 U8933 ( .A(n7661), .B(n7660), .C(n7659), .D(n7658), .Y(n7666) );
  AO22X1 U8934 ( .A0(net118269), .A1(n833), .B0(net118295), .B1(n2452), .Y(
        n7664) );
  NOR4X1 U8935 ( .A(n7580), .B(n7579), .C(n7578), .D(n7577), .Y(n7581) );
  OAI221XL U8936 ( .A0(\i_MIPS/Register/register[18][28] ), .A1(net117637), 
        .B0(\i_MIPS/Register/register[26][28] ), .B1(net117655), .C0(n7576), 
        .Y(n7579) );
  NAND4X1 U8937 ( .A(n7575), .B(n7574), .C(n7573), .D(n7572), .Y(n7580) );
  AO22X1 U8938 ( .A0(net118269), .A1(n899), .B0(net118295), .B1(n2528), .Y(
        n7578) );
  NAND4X1 U8939 ( .A(n6884), .B(n6883), .C(n6882), .D(n6881), .Y(n6889) );
  AO22X1 U8940 ( .A0(net118267), .A1(n301), .B0(net118295), .B1(n951), .Y(
        n6887) );
  NOR4X1 U8941 ( .A(n6789), .B(n6788), .C(n6787), .D(n6786), .Y(n6790) );
  OAI221XL U8942 ( .A0(\i_MIPS/Register/register[18][24] ), .A1(net117635), 
        .B0(\i_MIPS/Register/register[26][24] ), .B1(net117653), .C0(n6785), 
        .Y(n6788) );
  NAND4X1 U8943 ( .A(n6784), .B(n6783), .C(n6782), .D(n6781), .Y(n6789) );
  AO22X1 U8944 ( .A0(net118267), .A1(n303), .B0(net118295), .B1(n953), .Y(
        n6787) );
  AOI2BB1X1 U8945 ( .A0N(n10908), .A1N(n4768), .B0(n10907), .Y(n10909) );
  XOR3X1 U8946 ( .A(\i_MIPS/IF_ID[23] ), .B(n6016), .C(n10353), .Y(n10358) );
  AOI2BB1X1 U8947 ( .A0N(n10352), .A1N(n10361), .B0(n4811), .Y(n10353) );
  AOI2BB1X1 U8948 ( .A0N(n4749), .A1N(n4743), .B0(n4822), .Y(n10300) );
  AOI2BB1X1 U8949 ( .A0N(n4747), .A1N(n4766), .B0(n10136), .Y(n10137) );
  XOR3X1 U8950 ( .A(\i_MIPS/IF_ID[25] ), .B(n6016), .C(n11052), .Y(n11061) );
  AOI2BB1X1 U8951 ( .A0N(n4744), .A1N(n4769), .B0(n4820), .Y(n11052) );
  CLKINVX1 U8952 ( .A(n11327), .Y(n10074) );
  CLKINVX1 U8953 ( .A(n11325), .Y(n10231) );
  CLKINVX1 U8954 ( .A(n11324), .Y(n10133) );
  CLKINVX1 U8955 ( .A(n11323), .Y(n10097) );
  CLKINVX1 U8956 ( .A(n11322), .Y(n9846) );
  CLKINVX1 U8957 ( .A(n11321), .Y(n9890) );
  CLKINVX1 U8958 ( .A(n11320), .Y(n9868) );
  CLKINVX1 U8959 ( .A(n11318), .Y(n9934) );
  CLKINVX1 U8960 ( .A(n11342), .Y(n9661) );
  CLKINVX1 U8961 ( .A(n11341), .Y(n9683) );
  CLKINVX1 U8962 ( .A(n11339), .Y(n9653) );
  CLKINVX1 U8963 ( .A(n11338), .Y(n9631) );
  CLKINVX1 U8964 ( .A(n11337), .Y(n9609) );
  CLKINVX1 U8965 ( .A(n11312), .Y(n10824) );
  CLKINVX1 U8966 ( .A(n11316), .Y(n10867) );
  CLKINVX1 U8967 ( .A(n11315), .Y(n10961) );
  CLKINVX1 U8968 ( .A(n11313), .Y(n10890) );
  AOI2BB1X1 U8969 ( .A0N(n10489), .A1N(n10488), .B0(n4806), .Y(n10490) );
  XOR3X1 U8970 ( .A(\i_MIPS/IF_ID[22] ), .B(\i_MIPS/Sign_Extend[31] ), .C(
        n10340), .Y(n10345) );
  AOI2BB1XL U8971 ( .A0N(\i_MIPS/PC/n24 ), .A1N(net115799), .B0(n10343), .Y(
        n10344) );
  AOI2BB1X1 U8972 ( .A0N(n4748), .A1N(n4742), .B0(n4821), .Y(n10340) );
  AOI2BB1X1 U8973 ( .A0N(n10176), .A1N(n4767), .B0(n10165), .Y(n10166) );
  XOR3X1 U8974 ( .A(\i_MIPS/jump_addr[28] ), .B(n6016), .C(n10567), .Y(n10535)
         );
  AO22X1 U8975 ( .A0(n5556), .A1(n10554), .B0(n11054), .B1(n10537), .Y(n10533)
         );
  XOR3X1 U8976 ( .A(\i_MIPS/IF_ID[20] ), .B(n6016), .C(n10322), .Y(n10327) );
  AOI2BB1X1 U8977 ( .A0N(n10321), .A1N(n10330), .B0(n4812), .Y(n10322) );
  XOR3X1 U8978 ( .A(\i_MIPS/IF_ID[18] ), .B(n6016), .C(n4743), .Y(n10297) );
  AO22X1 U8979 ( .A0(n5555), .A1(n10646), .B0(n11054), .B1(n10294), .Y(n10295)
         );
  OAI221XL U8980 ( .A0(\i_MIPS/Register/register[18][3] ), .A1(n5088), .B0(
        \i_MIPS/Register/register[26][3] ), .B1(n5086), .C0(n9191), .Y(n9199)
         );
  OA22X1 U8981 ( .A0(\i_MIPS/Register/register[22][3] ), .A1(n5083), .B0(
        \i_MIPS/Register/register[30][3] ), .B1(n5079), .Y(n9191) );
  OAI221XL U8982 ( .A0(\i_MIPS/Register/register[2][3] ), .A1(n5088), .B0(
        \i_MIPS/Register/register[10][3] ), .B1(n5086), .C0(n9182), .Y(n9190)
         );
  OA22X1 U8983 ( .A0(\i_MIPS/Register/register[6][3] ), .A1(n5083), .B0(
        \i_MIPS/Register/register[14][3] ), .B1(n5079), .Y(n9182) );
  OAI221XL U8984 ( .A0(\i_MIPS/Register/register[2][14] ), .A1(net117637), 
        .B0(\i_MIPS/Register/register[10][14] ), .B1(net117657), .C0(n7745), 
        .Y(n7753) );
  OAI221XL U8985 ( .A0(\i_MIPS/Register/register[18][24] ), .A1(n5089), .B0(
        \i_MIPS/Register/register[26][24] ), .B1(n5084), .C0(n6620), .Y(n6628)
         );
  OAI221XL U8986 ( .A0(\i_MIPS/Register/register[2][24] ), .A1(n5091), .B0(
        \i_MIPS/Register/register[10][24] ), .B1(n5084), .C0(n6611), .Y(n6619)
         );
  OAI221XL U8987 ( .A0(\i_MIPS/Register/register[18][31] ), .A1(n5090), .B0(
        \i_MIPS/Register/register[26][31] ), .B1(n5086), .C0(n9498), .Y(n9514)
         );
  OAI221XL U8988 ( .A0(\i_MIPS/Register/register[2][31] ), .A1(n5090), .B0(
        \i_MIPS/Register/register[10][31] ), .B1(n5086), .C0(n9489), .Y(n9497)
         );
  OAI221XL U8989 ( .A0(\i_MIPS/Register/register[18][30] ), .A1(n5091), .B0(
        \i_MIPS/Register/register[26][30] ), .B1(n5084), .C0(n9393), .Y(n9401)
         );
  OAI221XL U8990 ( .A0(\i_MIPS/Register/register[2][30] ), .A1(n5091), .B0(
        \i_MIPS/Register/register[10][30] ), .B1(n5084), .C0(n9384), .Y(n9392)
         );
  OAI221XL U8991 ( .A0(\i_MIPS/Register/register[18][31] ), .A1(net117643), 
        .B0(\i_MIPS/Register/register[26][31] ), .B1(net117663), .C0(n9586), 
        .Y(n9594) );
  OAI221XL U8992 ( .A0(\i_MIPS/Register/register[2][30] ), .A1(net117643), 
        .B0(\i_MIPS/Register/register[10][30] ), .B1(net117663), .C0(n9467), 
        .Y(n9475) );
  XOR2XL U8993 ( .A(net110470), .B(\i_MIPS/ID_EX[113] ), .Y(n7741) );
  NAND2X1 U8994 ( .A(\i_MIPS/EX_MEM[5] ), .B(n5190), .Y(net104792) );
  AOI32XL U8995 ( .A0(net107404), .A1(\i_MIPS/ALUin1[30] ), .A2(n9443), .B0(
        n4696), .B1(n9442), .Y(n9460) );
  XNOR2X1 U8996 ( .A(net114079), .B(\i_MIPS/Reg_W[4] ), .Y(n6642) );
  XNOR2XL U8997 ( .A(\i_MIPS/Reg_W[3] ), .B(n10334), .Y(n6631) );
  AOI2BB1XL U8998 ( .A0N(\i_MIPS/ALUin1[15] ), .A1N(n5059), .B0(n4731), .Y(
        n7103) );
  XNOR2XL U8999 ( .A(\i_MIPS/Reg_W[1] ), .B(n248), .Y(n6632) );
  XNOR2XL U9000 ( .A(\i_MIPS/Reg_W[2] ), .B(net105477), .Y(n6629) );
  XNOR2XL U9001 ( .A(\i_MIPS/Reg_W[0] ), .B(\i_MIPS/jump_addr[18] ), .Y(n6630)
         );
  NAND2X1 U9002 ( .A(\i_MIPS/IF_ID[4] ), .B(\i_MIPS/Sign_Extend[2] ), .Y(
        n10906) );
  NAND2XL U9003 ( .A(n4755), .B(\i_MIPS/ALUin1[7] ), .Y(n8980) );
  NAND2XL U9004 ( .A(\i_MIPS/ALU/N303 ), .B(n9555), .Y(n9569) );
  NAND4BX1 U9005 ( .AN(n7727), .B(n7726), .C(n7725), .D(n7724), .Y(n7738) );
  OA22X1 U9006 ( .A0(\i_MIPS/Register/register[4][27] ), .A1(n5101), .B0(
        \i_MIPS/Register/register[12][27] ), .B1(n5093), .Y(n7726) );
  OA22X1 U9007 ( .A0(\i_MIPS/Register/register[0][27] ), .A1(n5107), .B0(
        \i_MIPS/Register/register[8][27] ), .B1(n5105), .Y(n7725) );
  NAND4BX1 U9008 ( .AN(n7736), .B(n7735), .C(n7734), .D(n7733), .Y(n7737) );
  OA22X1 U9009 ( .A0(\i_MIPS/Register/register[20][27] ), .A1(n5099), .B0(
        \i_MIPS/Register/register[28][27] ), .B1(n5093), .Y(n7735) );
  OA22X1 U9010 ( .A0(\i_MIPS/Register/register[16][27] ), .A1(n5107), .B0(
        \i_MIPS/Register/register[24][27] ), .B1(n5105), .Y(n7734) );
  OAI2BB2XL U9011 ( .B0(\i_MIPS/n154 ), .B1(net115795), .A0N(\i_MIPS/PC_o[1] ), 
        .A1N(n4544), .Y(\i_MIPS/N18 ) );
  OAI2BB2XL U9012 ( .B0(\i_MIPS/n165 ), .B1(net115795), .A0N(n10478), .A1N(
        n4545), .Y(\i_MIPS/N29 ) );
  CLKINVX1 U9013 ( .A(n10477), .Y(n10478) );
  OAI2BB2XL U9014 ( .B0(\i_MIPS/n166 ), .B1(net115795), .A0N(n10486), .A1N(
        n4544), .Y(\i_MIPS/N30 ) );
  CLKINVX1 U9015 ( .A(n10485), .Y(n10486) );
  OAI2BB2XL U9016 ( .B0(\i_MIPS/n167 ), .B1(net115795), .A0N(n10497), .A1N(
        n4545), .Y(\i_MIPS/N31 ) );
  CLKINVX1 U9017 ( .A(n10496), .Y(n10497) );
  OAI2BB2XL U9018 ( .B0(\i_MIPS/n174 ), .B1(net115797), .A0N(n10339), .A1N(
        n4544), .Y(\i_MIPS/N38 ) );
  CLKINVX1 U9019 ( .A(n10338), .Y(n10339) );
  OAI2BB2XL U9020 ( .B0(\i_MIPS/n175 ), .B1(net115797), .A0N(n10347), .A1N(
        n4545), .Y(\i_MIPS/N39 ) );
  CLKINVX1 U9021 ( .A(n10346), .Y(n10347) );
  OAI2BB2XL U9022 ( .B0(\i_MIPS/n176 ), .B1(net115797), .A0N(n10360), .A1N(
        n4544), .Y(\i_MIPS/N40 ) );
  CLKINVX1 U9023 ( .A(n10359), .Y(n10360) );
  OAI2BB2XL U9024 ( .B0(\i_MIPS/n177 ), .B1(net115797), .A0N(n10370), .A1N(
        n4545), .Y(\i_MIPS/N41 ) );
  CLKINVX1 U9025 ( .A(n10369), .Y(n10370) );
  OAI2BB2XL U9026 ( .B0(\i_MIPS/n179 ), .B1(net115797), .A0N(n10383), .A1N(
        n4544), .Y(\i_MIPS/N43 ) );
  CLKINVX1 U9027 ( .A(n10382), .Y(n10383) );
  OAI2BB2XL U9028 ( .B0(\i_MIPS/n180 ), .B1(net115795), .A0N(n10390), .A1N(
        n4544), .Y(\i_MIPS/N44 ) );
  CLKINVX1 U9029 ( .A(n10389), .Y(n10390) );
  OAI2BB2XL U9030 ( .B0(\i_MIPS/n178 ), .B1(net115797), .A0N(n4544), .A1N(
        n10372), .Y(\i_MIPS/N42 ) );
  INVXL U9031 ( .A(n11060), .Y(n10372) );
  OAI2BB2XL U9032 ( .B0(\i_MIPS/n158 ), .B1(net115795), .A0N(n4545), .A1N(
        n10052), .Y(\i_MIPS/N22 ) );
  CLKINVX1 U9033 ( .A(n10913), .Y(n10052) );
  OAI2BB2XL U9034 ( .B0(\i_MIPS/n153 ), .B1(net115793), .A0N(
        \i_MIPS/PC_add4[0] ), .A1N(n4545), .Y(\i_MIPS/N17 ) );
  OAI2BB2XL U9035 ( .B0(\i_MIPS/n160 ), .B1(net115795), .A0N(n10143), .A1N(
        n4545), .Y(\i_MIPS/N24 ) );
  CLKINVX1 U9036 ( .A(n10142), .Y(n10143) );
  CLKINVX1 U9037 ( .A(n10151), .Y(n10152) );
  OAI2BB2XL U9038 ( .B0(\i_MIPS/n162 ), .B1(net115795), .A0N(n10163), .A1N(
        n4544), .Y(\i_MIPS/N26 ) );
  CLKINVX1 U9039 ( .A(n10162), .Y(n10163) );
  OAI2BB2XL U9040 ( .B0(\i_MIPS/n163 ), .B1(net115795), .A0N(n10173), .A1N(
        n4545), .Y(\i_MIPS/N27 ) );
  CLKINVX1 U9041 ( .A(n10172), .Y(n10173) );
  OAI2BB2XL U9042 ( .B0(\i_MIPS/n164 ), .B1(net115795), .A0N(n10184), .A1N(
        n4544), .Y(\i_MIPS/N28 ) );
  CLKINVX1 U9043 ( .A(n10183), .Y(n10184) );
  OAI2BB2XL U9044 ( .B0(\i_MIPS/n168 ), .B1(net115795), .A0N(n10270), .A1N(
        n4545), .Y(\i_MIPS/N32 ) );
  CLKINVX1 U9045 ( .A(n10269), .Y(n10270) );
  OAI2BB2XL U9046 ( .B0(\i_MIPS/n169 ), .B1(net115795), .A0N(n10278), .A1N(
        n4544), .Y(\i_MIPS/N33 ) );
  CLKINVX1 U9047 ( .A(n10277), .Y(n10278) );
  OAI2BB2XL U9048 ( .B0(\i_MIPS/n170 ), .B1(net115795), .A0N(n10287), .A1N(
        n4545), .Y(\i_MIPS/N34 ) );
  CLKINVX1 U9049 ( .A(n10286), .Y(n10287) );
  OAI2BB2XL U9050 ( .B0(\i_MIPS/n171 ), .B1(net115797), .A0N(n10299), .A1N(
        n4545), .Y(\i_MIPS/N35 ) );
  CLKINVX1 U9051 ( .A(n10298), .Y(n10299) );
  OAI2BB2XL U9052 ( .B0(\i_MIPS/n172 ), .B1(net115797), .A0N(n10306), .A1N(
        n4544), .Y(\i_MIPS/N36 ) );
  CLKINVX1 U9053 ( .A(n10305), .Y(n10306) );
  OAI2BB2XL U9054 ( .B0(\i_MIPS/n173 ), .B1(net115797), .A0N(n10329), .A1N(
        n4545), .Y(\i_MIPS/N37 ) );
  CLKINVX1 U9055 ( .A(n10328), .Y(n10329) );
  OAI2BB2XL U9056 ( .B0(\i_MIPS/n155 ), .B1(net115793), .A0N(n4544), .A1N(
        \i_MIPS/PC/n4 ), .Y(\i_MIPS/N19 ) );
  OAI2BB2XL U9057 ( .B0(\i_MIPS/n156 ), .B1(net115793), .A0N(n4545), .A1N(
        n9728), .Y(\i_MIPS/N20 ) );
  CLKINVX1 U9058 ( .A(n9734), .Y(n9728) );
  OAI2BB2XL U9059 ( .B0(\i_MIPS/n157 ), .B1(net115793), .A0N(n4544), .A1N(
        n9803), .Y(\i_MIPS/N21 ) );
  CLKINVX1 U9060 ( .A(n10936), .Y(n9803) );
  OAI2BB2XL U9061 ( .B0(\i_MIPS/n159 ), .B1(net115793), .A0N(n4545), .A1N(
        n9937), .Y(\i_MIPS/N23 ) );
  CLKINVX1 U9062 ( .A(n10871), .Y(n9937) );
  NAND2BX1 U9063 ( .AN(\i_MIPS/Sign_Extend[9] ), .B(\i_MIPS/n164 ), .Y(n10258)
         );
  NAND2X1 U9064 ( .A(\i_MIPS/n167 ), .B(\i_MIPS/n509 ), .Y(n10254) );
  AND2X2 U9065 ( .A(n6529), .B(mem_ready_I), .Y(n11214) );
  NAND4X1 U9066 ( .A(n9062), .B(n9061), .C(n9060), .D(n9059), .Y(n9067) );
  NAND4X1 U9067 ( .A(n6986), .B(n6985), .C(n6984), .D(n6983), .Y(n6991) );
  OA22X1 U9068 ( .A0(\i_MIPS/Register/register[5][29] ), .A1(net118399), .B0(
        \i_MIPS/Register/register[13][29] ), .B1(net118423), .Y(n6985) );
  OA22X1 U9069 ( .A0(\i_MIPS/Register/register[1][29] ), .A1(net118453), .B0(
        \i_MIPS/Register/register[9][29] ), .B1(net118479), .Y(n6986) );
  OA22X1 U9070 ( .A0(\i_MIPS/Register/register[7][29] ), .A1(net118303), .B0(
        \i_MIPS/Register/register[15][29] ), .B1(net118327), .Y(n6983) );
  NAND4X1 U9071 ( .A(n7243), .B(n7242), .C(n7241), .D(n7240), .Y(n7248) );
  OA22X1 U9072 ( .A0(\i_MIPS/Register/register[5][6] ), .A1(net118399), .B0(
        \i_MIPS/Register/register[13][6] ), .B1(net118423), .Y(n7242) );
  OA22X1 U9073 ( .A0(\i_MIPS/Register/register[1][6] ), .A1(net118453), .B0(
        \i_MIPS/Register/register[9][6] ), .B1(net118479), .Y(n7243) );
  OA22X1 U9074 ( .A0(\i_MIPS/Register/register[7][6] ), .A1(net118303), .B0(
        \i_MIPS/Register/register[15][6] ), .B1(net118327), .Y(n7240) );
  NAND4X1 U9075 ( .A(n7082), .B(n7081), .C(n7080), .D(n7079), .Y(n7087) );
  OA22X1 U9076 ( .A0(\i_MIPS/Register/register[5][23] ), .A1(net118399), .B0(
        \i_MIPS/Register/register[13][23] ), .B1(net118423), .Y(n7081) );
  OA22X1 U9077 ( .A0(\i_MIPS/Register/register[1][23] ), .A1(net118453), .B0(
        \i_MIPS/Register/register[9][23] ), .B1(net118479), .Y(n7082) );
  OA22X1 U9078 ( .A0(\i_MIPS/Register/register[7][23] ), .A1(net118303), .B0(
        \i_MIPS/Register/register[15][23] ), .B1(net118327), .Y(n7079) );
  NAND4X1 U9079 ( .A(n7168), .B(n7167), .C(n7166), .D(n7165), .Y(n7173) );
  OA22X1 U9080 ( .A0(\i_MIPS/Register/register[5][2] ), .A1(net118399), .B0(
        \i_MIPS/Register/register[13][2] ), .B1(net118423), .Y(n7167) );
  OA22X1 U9081 ( .A0(\i_MIPS/Register/register[1][2] ), .A1(net118453), .B0(
        \i_MIPS/Register/register[9][2] ), .B1(net118479), .Y(n7168) );
  OA22X1 U9082 ( .A0(\i_MIPS/Register/register[7][2] ), .A1(net118303), .B0(
        \i_MIPS/Register/register[15][2] ), .B1(net118327), .Y(n7165) );
  NAND4X1 U9083 ( .A(n6875), .B(n6874), .C(n6873), .D(n6872), .Y(n6880) );
  OA22X1 U9084 ( .A0(\i_MIPS/Register/register[5][25] ), .A1(net118399), .B0(
        \i_MIPS/Register/register[13][25] ), .B1(net118423), .Y(n6874) );
  OA22X1 U9085 ( .A0(\i_MIPS/Register/register[1][25] ), .A1(net118453), .B0(
        \i_MIPS/Register/register[9][25] ), .B1(net118479), .Y(n6875) );
  OA22X1 U9086 ( .A0(\i_MIPS/Register/register[7][25] ), .A1(net118303), .B0(
        \i_MIPS/Register/register[15][25] ), .B1(net118327), .Y(n6872) );
  NAND4X1 U9087 ( .A(n7566), .B(n7565), .C(n7564), .D(n7563), .Y(n7571) );
  OA22X1 U9088 ( .A0(\i_MIPS/Register/register[7][28] ), .A1(net118305), .B0(
        \i_MIPS/Register/register[15][28] ), .B1(net118329), .Y(n7563) );
  NAND4X1 U9089 ( .A(n7508), .B(n7507), .C(n7506), .D(n7505), .Y(n7513) );
  OA22X1 U9090 ( .A0(\i_MIPS/Register/register[5][10] ), .A1(net118401), .B0(
        \i_MIPS/Register/register[13][10] ), .B1(net118425), .Y(n7507) );
  OA22X1 U9091 ( .A0(\i_MIPS/Register/register[1][10] ), .A1(net118453), .B0(
        \i_MIPS/Register/register[9][10] ), .B1(net118473), .Y(n7508) );
  OA22X1 U9092 ( .A0(\i_MIPS/Register/register[7][10] ), .A1(net118305), .B0(
        \i_MIPS/Register/register[15][10] ), .B1(net118329), .Y(n7505) );
  NAND4X1 U9093 ( .A(n7382), .B(n7381), .C(n7380), .D(n7379), .Y(n7387) );
  NAND4X1 U9094 ( .A(n7652), .B(n7651), .C(n7650), .D(n7649), .Y(n7657) );
  OA22X1 U9095 ( .A0(\i_MIPS/Register/register[5][27] ), .A1(net118401), .B0(
        \i_MIPS/Register/register[13][27] ), .B1(net118425), .Y(n7651) );
  OA22X1 U9096 ( .A0(\i_MIPS/Register/register[1][27] ), .A1(net118453), .B0(
        \i_MIPS/Register/register[9][27] ), .B1(net118473), .Y(n7652) );
  OA22X1 U9097 ( .A0(\i_MIPS/Register/register[7][27] ), .A1(net118305), .B0(
        \i_MIPS/Register/register[15][27] ), .B1(net118329), .Y(n7649) );
  NAND4X1 U9098 ( .A(n8495), .B(n8494), .C(n8493), .D(n8492), .Y(n8500) );
  OA22X1 U9099 ( .A0(\i_MIPS/Register/register[5][11] ), .A1(net118403), .B0(
        \i_MIPS/Register/register[13][11] ), .B1(net118423), .Y(n8494) );
  OA22X1 U9100 ( .A0(\i_MIPS/Register/register[1][11] ), .A1(net118451), .B0(
        \i_MIPS/Register/register[9][11] ), .B1(net118475), .Y(n8495) );
  OA22X1 U9101 ( .A0(\i_MIPS/Register/register[7][11] ), .A1(net118307), .B0(
        \i_MIPS/Register/register[15][11] ), .B1(net118331), .Y(n8492) );
  NAND4X1 U9102 ( .A(n8314), .B(n8313), .C(n8312), .D(n8311), .Y(n8319) );
  OA22X1 U9103 ( .A0(\i_MIPS/Register/register[5][19] ), .A1(net118403), .B0(
        \i_MIPS/Register/register[13][19] ), .B1(net118429), .Y(n8313) );
  OA22X1 U9104 ( .A0(\i_MIPS/Register/register[1][19] ), .A1(net118451), .B0(
        \i_MIPS/Register/register[9][19] ), .B1(net118475), .Y(n8314) );
  OA22X1 U9105 ( .A0(\i_MIPS/Register/register[7][19] ), .A1(net118307), .B0(
        \i_MIPS/Register/register[15][19] ), .B1(net118331), .Y(n8311) );
  NAND4X1 U9106 ( .A(n8578), .B(n8577), .C(n8576), .D(n8575), .Y(n8583) );
  OA22X1 U9107 ( .A0(\i_MIPS/Register/register[5][18] ), .A1(net118405), .B0(
        \i_MIPS/Register/register[13][18] ), .B1(net118429), .Y(n8577) );
  OA22X1 U9108 ( .A0(\i_MIPS/Register/register[1][18] ), .A1(net118453), .B0(
        \i_MIPS/Register/register[9][18] ), .B1(net118477), .Y(n8578) );
  OA22X1 U9109 ( .A0(\i_MIPS/Register/register[7][18] ), .A1(net118303), .B0(
        \i_MIPS/Register/register[15][18] ), .B1(net118329), .Y(n8575) );
  NAND4X1 U9110 ( .A(n7971), .B(n7970), .C(n7969), .D(n7968), .Y(n7976) );
  OA22X1 U9111 ( .A0(\i_MIPS/Register/register[5][13] ), .A1(net118403), .B0(
        \i_MIPS/Register/register[13][13] ), .B1(net118429), .Y(n7970) );
  OA22X1 U9112 ( .A0(\i_MIPS/Register/register[1][13] ), .A1(net118451), .B0(
        \i_MIPS/Register/register[9][13] ), .B1(net118475), .Y(n7971) );
  OA22X1 U9113 ( .A0(\i_MIPS/Register/register[7][13] ), .A1(net118307), .B0(
        \i_MIPS/Register/register[15][13] ), .B1(net118331), .Y(n7968) );
  NAND4X1 U9114 ( .A(n8224), .B(n8223), .C(n8222), .D(n8221), .Y(n8229) );
  OA22X1 U9115 ( .A0(\i_MIPS/Register/register[7][12] ), .A1(net118307), .B0(
        \i_MIPS/Register/register[15][12] ), .B1(net118331), .Y(n8221) );
  OA22X1 U9116 ( .A0(\i_MIPS/Register/register[7][8] ), .A1(net118307), .B0(
        \i_MIPS/Register/register[15][8] ), .B1(net118331), .Y(n8141) );
  NAND4X1 U9117 ( .A(n8053), .B(n8052), .C(n8051), .D(n8050), .Y(n8058) );
  OA22X1 U9118 ( .A0(\i_MIPS/Register/register[5][9] ), .A1(net118403), .B0(
        \i_MIPS/Register/register[13][9] ), .B1(net118429), .Y(n8052) );
  OA22X1 U9119 ( .A0(\i_MIPS/Register/register[1][9] ), .A1(net118451), .B0(
        \i_MIPS/Register/register[9][9] ), .B1(net118475), .Y(n8053) );
  OA22X1 U9120 ( .A0(\i_MIPS/Register/register[7][9] ), .A1(net118307), .B0(
        \i_MIPS/Register/register[15][9] ), .B1(net118331), .Y(n8050) );
  OA22X1 U9121 ( .A0(\i_MIPS/Register/register[5][5] ), .A1(net118407), .B0(
        \i_MIPS/Register/register[13][5] ), .B1(net118431), .Y(n9328) );
  OA22X1 U9122 ( .A0(\i_MIPS/Register/register[1][5] ), .A1(net118455), .B0(
        \i_MIPS/Register/register[9][5] ), .B1(net118479), .Y(n9329) );
  OA22X1 U9123 ( .A0(\i_MIPS/Register/register[7][5] ), .A1(net118311), .B0(
        \i_MIPS/Register/register[15][5] ), .B1(net118335), .Y(n9326) );
  OA22X1 U9124 ( .A0(\i_MIPS/Register/register[5][3] ), .A1(net118407), .B0(
        \i_MIPS/Register/register[13][3] ), .B1(net118431), .Y(n9147) );
  OA22X1 U9125 ( .A0(\i_MIPS/Register/register[1][3] ), .A1(net118455), .B0(
        \i_MIPS/Register/register[9][3] ), .B1(net118479), .Y(n9148) );
  OA22X1 U9126 ( .A0(\i_MIPS/Register/register[7][3] ), .A1(net118311), .B0(
        \i_MIPS/Register/register[15][3] ), .B1(net118335), .Y(n9145) );
  NAND4X1 U9127 ( .A(n8902), .B(n8901), .C(n8900), .D(n8899), .Y(n8907) );
  NAND4X1 U9128 ( .A(n8724), .B(n8723), .C(n8722), .D(n8721), .Y(n8729) );
  OA22X1 U9129 ( .A0(\i_MIPS/Register/register[5][0] ), .A1(net118405), .B0(
        \i_MIPS/Register/register[13][0] ), .B1(net118429), .Y(n8723) );
  OA22X1 U9130 ( .A0(\i_MIPS/Register/register[1][0] ), .A1(net118453), .B0(
        \i_MIPS/Register/register[9][0] ), .B1(net118477), .Y(n8724) );
  OA22X1 U9131 ( .A0(\i_MIPS/Register/register[7][0] ), .A1(net118311), .B0(
        \i_MIPS/Register/register[15][0] ), .B1(net118329), .Y(n8721) );
  NAND4X1 U9132 ( .A(n8987), .B(n8986), .C(n8985), .D(n8984), .Y(n8992) );
  OA22X1 U9133 ( .A0(\i_MIPS/Register/register[5][1] ), .A1(net118405), .B0(
        \i_MIPS/Register/register[13][1] ), .B1(net118429), .Y(n8986) );
  OA22X1 U9134 ( .A0(\i_MIPS/Register/register[1][1] ), .A1(net118453), .B0(
        \i_MIPS/Register/register[9][1] ), .B1(net118477), .Y(n8987) );
  OA22X1 U9135 ( .A0(\i_MIPS/Register/register[7][1] ), .A1(net118307), .B0(
        \i_MIPS/Register/register[15][1] ), .B1(net118327), .Y(n8984) );
  NAND4X1 U9136 ( .A(n8800), .B(n8799), .C(n8798), .D(n8797), .Y(n8805) );
  OA22X1 U9137 ( .A0(\i_MIPS/Register/register[5][16] ), .A1(net118405), .B0(
        \i_MIPS/Register/register[13][16] ), .B1(net118429), .Y(n8799) );
  OA22X1 U9138 ( .A0(\i_MIPS/Register/register[1][16] ), .A1(net118453), .B0(
        \i_MIPS/Register/register[9][16] ), .B1(net118477), .Y(n8800) );
  OA22X1 U9139 ( .A0(\i_MIPS/Register/register[7][16] ), .A1(net118307), .B0(
        \i_MIPS/Register/register[15][16] ), .B1(net118331), .Y(n8797) );
  OA22X1 U9140 ( .A0(\i_MIPS/Register/register[5][24] ), .A1(net118399), .B0(
        \i_MIPS/Register/register[13][24] ), .B1(net118423), .Y(n6773) );
  OA22X1 U9141 ( .A0(\i_MIPS/Register/register[7][24] ), .A1(net118303), .B0(
        \i_MIPS/Register/register[15][24] ), .B1(net118327), .Y(n6771) );
  NAND4X1 U9142 ( .A(n7933), .B(n7932), .C(n7931), .D(n7930), .Y(n7938) );
  NAND4X1 U9143 ( .A(n7924), .B(n7923), .C(n7922), .D(n7921), .Y(n7929) );
  NAND4X1 U9144 ( .A(n7895), .B(n7894), .C(n7893), .D(n7892), .Y(n7900) );
  OA22XL U9145 ( .A0(\i_MIPS/Register/register[21][22] ), .A1(n7887), .B0(
        \i_MIPS/Register/register[29][22] ), .B1(n7886), .Y(n7894) );
  OA22XL U9146 ( .A0(\i_MIPS/Register/register[17][22] ), .A1(n7885), .B0(
        \i_MIPS/Register/register[25][22] ), .B1(n7884), .Y(n7895) );
  OA22XL U9147 ( .A0(\i_MIPS/Register/register[23][22] ), .A1(n7891), .B0(
        \i_MIPS/Register/register[31][22] ), .B1(n7890), .Y(n7892) );
  NAND4X1 U9148 ( .A(n7878), .B(n7877), .C(n7876), .D(n7875), .Y(n7883) );
  OA22XL U9149 ( .A0(\i_MIPS/Register/register[5][22] ), .A1(n7887), .B0(
        \i_MIPS/Register/register[13][22] ), .B1(n7886), .Y(n7877) );
  OA22XL U9150 ( .A0(\i_MIPS/Register/register[1][22] ), .A1(n7885), .B0(
        \i_MIPS/Register/register[9][22] ), .B1(n7884), .Y(n7878) );
  OA22XL U9151 ( .A0(\i_MIPS/Register/register[7][22] ), .A1(n7891), .B0(
        \i_MIPS/Register/register[15][22] ), .B1(n7890), .Y(n7875) );
  OAI22XL U9152 ( .A0(n3586), .A1(n5952), .B0(\i_MIPS/n269 ), .B1(n3597), .Y(
        \i_MIPS/n460 ) );
  OAI22XL U9153 ( .A0(\i_MIPS/n302 ), .A1(n3586), .B0(\i_MIPS/n303 ), .B1(
        n3601), .Y(\i_MIPS/n493 ) );
  OAI22XL U9154 ( .A0(\i_MIPS/n269 ), .A1(n3586), .B0(\i_MIPS/n268 ), .B1(
        n3590), .Y(\i_MIPS/n459 ) );
  OAI22XL U9155 ( .A0(\i_MIPS/n246 ), .A1(n3586), .B0(\i_MIPS/n245 ), .B1(
        n3589), .Y(\i_MIPS/n409 ) );
  NAND4BX1 U9156 ( .AN(n9585), .B(n9584), .C(n9583), .D(n9582), .Y(n9596) );
  OA22XL U9157 ( .A0(\i_MIPS/Register/register[4][31] ), .A1(net107169), .B0(
        \i_MIPS/Register/register[12][31] ), .B1(net107170), .Y(n9584) );
  OA22XL U9158 ( .A0(\i_MIPS/Register/register[0][31] ), .A1(net107167), .B0(
        \i_MIPS/Register/register[8][31] ), .B1(net107168), .Y(n9583) );
  OAI221XL U9159 ( .A0(\i_MIPS/Register/register[2][31] ), .A1(net117643), 
        .B0(\i_MIPS/Register/register[10][31] ), .B1(net117663), .C0(n9577), 
        .Y(n9585) );
  OA22X1 U9160 ( .A0(\i_MIPS/Register/register[0][17] ), .A1(n5107), .B0(
        \i_MIPS/Register/register[8][17] ), .B1(n5105), .Y(n9279) );
  NAND4BX1 U9161 ( .AN(n9030), .B(n9029), .C(n9028), .D(n9027), .Y(n9041) );
  OA22X1 U9162 ( .A0(\i_MIPS/Register/register[4][1] ), .A1(n5101), .B0(
        \i_MIPS/Register/register[12][1] ), .B1(n5095), .Y(n9029) );
  OA22X1 U9163 ( .A0(\i_MIPS/Register/register[0][1] ), .A1(n5109), .B0(
        \i_MIPS/Register/register[8][1] ), .B1(n5104), .Y(n9028) );
  OAI221XL U9164 ( .A0(\i_MIPS/Register/register[2][1] ), .A1(n5091), .B0(
        \i_MIPS/Register/register[10][1] ), .B1(n5086), .C0(n9022), .Y(n9030)
         );
  NAND4BX1 U9165 ( .AN(n8267), .B(n8266), .C(n8265), .D(n8264), .Y(n8278) );
  OA22X1 U9166 ( .A0(\i_MIPS/Register/register[4][12] ), .A1(n5100), .B0(
        \i_MIPS/Register/register[12][12] ), .B1(n5094), .Y(n8266) );
  OA22X1 U9167 ( .A0(\i_MIPS/Register/register[0][12] ), .A1(n5108), .B0(
        \i_MIPS/Register/register[8][12] ), .B1(n5103), .Y(n8265) );
  OAI221XL U9168 ( .A0(\i_MIPS/Register/register[2][12] ), .A1(n5090), .B0(
        \i_MIPS/Register/register[10][12] ), .B1(n5085), .C0(n8259), .Y(n8267)
         );
  NAND4BX1 U9169 ( .AN(n8620), .B(n8619), .C(n8618), .D(n8617), .Y(n8631) );
  OA22X1 U9170 ( .A0(\i_MIPS/Register/register[4][18] ), .A1(n5101), .B0(
        \i_MIPS/Register/register[12][18] ), .B1(n5095), .Y(n8619) );
  OA22X1 U9171 ( .A0(\i_MIPS/Register/register[0][18] ), .A1(n5109), .B0(
        \i_MIPS/Register/register[8][18] ), .B1(n5104), .Y(n8618) );
  OAI221XL U9172 ( .A0(\i_MIPS/Register/register[2][18] ), .A1(n5091), .B0(
        \i_MIPS/Register/register[10][18] ), .B1(n4669), .C0(n8612), .Y(n8620)
         );
  OA22X1 U9173 ( .A0(\i_MIPS/Register/register[0][5] ), .A1(n5109), .B0(
        \i_MIPS/Register/register[8][5] ), .B1(n5105), .Y(n9370) );
  OAI221XL U9174 ( .A0(\i_MIPS/Register/register[2][5] ), .A1(n5091), .B0(
        \i_MIPS/Register/register[10][5] ), .B1(n5086), .C0(n9364), .Y(n9372)
         );
  OA22X1 U9175 ( .A0(\i_MIPS/Register/register[4][0] ), .A1(n5101), .B0(
        \i_MIPS/Register/register[12][0] ), .B1(n5095), .Y(n8766) );
  OA22X1 U9176 ( .A0(\i_MIPS/Register/register[0][0] ), .A1(n5109), .B0(
        \i_MIPS/Register/register[8][0] ), .B1(n5104), .Y(n8765) );
  NAND4BX1 U9177 ( .AN(n8538), .B(n8537), .C(n8536), .D(n8535), .Y(n8549) );
  OA22X1 U9178 ( .A0(\i_MIPS/Register/register[4][11] ), .A1(n5100), .B0(
        \i_MIPS/Register/register[12][11] ), .B1(n5094), .Y(n8537) );
  OA22X1 U9179 ( .A0(\i_MIPS/Register/register[0][11] ), .A1(n5108), .B0(
        \i_MIPS/Register/register[8][11] ), .B1(n5103), .Y(n8536) );
  OAI221XL U9180 ( .A0(\i_MIPS/Register/register[2][11] ), .A1(n5091), .B0(
        \i_MIPS/Register/register[10][11] ), .B1(n4669), .C0(n8530), .Y(n8538)
         );
  NAND4BX1 U9181 ( .AN(n8843), .B(n8842), .C(n8841), .D(n8840), .Y(n8854) );
  OA22X1 U9182 ( .A0(\i_MIPS/Register/register[4][16] ), .A1(n5101), .B0(
        \i_MIPS/Register/register[12][16] ), .B1(n5095), .Y(n8842) );
  OA22X1 U9183 ( .A0(\i_MIPS/Register/register[0][16] ), .A1(n5109), .B0(
        \i_MIPS/Register/register[8][16] ), .B1(n5104), .Y(n8841) );
  OAI221XL U9184 ( .A0(\i_MIPS/Register/register[2][16] ), .A1(n5091), .B0(
        \i_MIPS/Register/register[10][16] ), .B1(n5087), .C0(n8835), .Y(n8843)
         );
  NAND4BX1 U9185 ( .AN(n8447), .B(n8446), .C(n8445), .D(n8444), .Y(n8458) );
  OA22X1 U9186 ( .A0(\i_MIPS/Register/register[4][20] ), .A1(n5100), .B0(
        \i_MIPS/Register/register[12][20] ), .B1(n5094), .Y(n8446) );
  OA22X1 U9187 ( .A0(\i_MIPS/Register/register[0][20] ), .A1(n5108), .B0(
        \i_MIPS/Register/register[8][20] ), .B1(n5103), .Y(n8445) );
  OAI221XL U9188 ( .A0(\i_MIPS/Register/register[2][20] ), .A1(n5090), .B0(
        \i_MIPS/Register/register[10][20] ), .B1(n4669), .C0(n8439), .Y(n8447)
         );
  NAND4BX1 U9189 ( .AN(n8357), .B(n8356), .C(n8355), .D(n8354), .Y(n8368) );
  OA22X1 U9190 ( .A0(\i_MIPS/Register/register[4][19] ), .A1(n5100), .B0(
        \i_MIPS/Register/register[12][19] ), .B1(n5094), .Y(n8356) );
  OA22X1 U9191 ( .A0(\i_MIPS/Register/register[0][19] ), .A1(n5108), .B0(
        \i_MIPS/Register/register[8][19] ), .B1(n5103), .Y(n8355) );
  NAND4BX1 U9192 ( .AN(n8946), .B(n8945), .C(n8944), .D(n8943), .Y(n8957) );
  OA22X1 U9193 ( .A0(\i_MIPS/Register/register[4][21] ), .A1(n5101), .B0(
        \i_MIPS/Register/register[12][21] ), .B1(n5095), .Y(n8945) );
  OA22X1 U9194 ( .A0(\i_MIPS/Register/register[0][21] ), .A1(n5109), .B0(
        \i_MIPS/Register/register[8][21] ), .B1(n5104), .Y(n8944) );
  OAI221XL U9195 ( .A0(\i_MIPS/Register/register[2][21] ), .A1(n5091), .B0(
        \i_MIPS/Register/register[10][21] ), .B1(n5086), .C0(n8938), .Y(n8946)
         );
  NAND4BX1 U9196 ( .AN(n8187), .B(n8186), .C(n8185), .D(n8184), .Y(n8198) );
  OA22X1 U9197 ( .A0(\i_MIPS/Register/register[4][8] ), .A1(n5100), .B0(
        \i_MIPS/Register/register[12][8] ), .B1(n5094), .Y(n8186) );
  OA22X1 U9198 ( .A0(\i_MIPS/Register/register[0][8] ), .A1(n5108), .B0(
        \i_MIPS/Register/register[8][8] ), .B1(n5103), .Y(n8185) );
  OAI221XL U9199 ( .A0(\i_MIPS/Register/register[2][8] ), .A1(n5090), .B0(
        \i_MIPS/Register/register[10][8] ), .B1(n5085), .C0(n8179), .Y(n8187)
         );
  NAND4BX1 U9200 ( .AN(n7466), .B(n7465), .C(n7464), .D(n7463), .Y(n7477) );
  OA22X1 U9201 ( .A0(\i_MIPS/Register/register[4][26] ), .A1(n5099), .B0(
        \i_MIPS/Register/register[12][26] ), .B1(n5093), .Y(n7465) );
  OA22X1 U9202 ( .A0(\i_MIPS/Register/register[0][26] ), .A1(n5107), .B0(
        \i_MIPS/Register/register[8][26] ), .B1(n5105), .Y(n7464) );
  OAI221XL U9203 ( .A0(\i_MIPS/Register/register[2][26] ), .A1(n5089), .B0(
        \i_MIPS/Register/register[10][26] ), .B1(n5085), .C0(n7458), .Y(n7466)
         );
  NAND4BX1 U9204 ( .AN(n7551), .B(n7550), .C(n7549), .D(n7548), .Y(n7562) );
  OA22X1 U9205 ( .A0(\i_MIPS/Register/register[4][10] ), .A1(n5101), .B0(
        \i_MIPS/Register/register[12][10] ), .B1(n5093), .Y(n7550) );
  OA22X1 U9206 ( .A0(\i_MIPS/Register/register[0][10] ), .A1(n5107), .B0(
        \i_MIPS/Register/register[8][10] ), .B1(n5105), .Y(n7549) );
  OAI221XL U9207 ( .A0(\i_MIPS/Register/register[2][10] ), .A1(n5089), .B0(
        \i_MIPS/Register/register[10][10] ), .B1(n5085), .C0(n7543), .Y(n7551)
         );
  OA22X1 U9208 ( .A0(\i_MIPS/Register/register[4][4] ), .A1(n5101), .B0(
        \i_MIPS/Register/register[12][4] ), .B1(n5095), .Y(n9105) );
  OA22X1 U9209 ( .A0(\i_MIPS/Register/register[0][4] ), .A1(n5109), .B0(
        \i_MIPS/Register/register[8][4] ), .B1(n5104), .Y(n9104) );
  OAI221XL U9210 ( .A0(\i_MIPS/Register/register[2][4] ), .A1(n5088), .B0(
        \i_MIPS/Register/register[10][4] ), .B1(n5086), .C0(n9098), .Y(n9106)
         );
  NAND4BX1 U9211 ( .AN(n8097), .B(n8096), .C(n8095), .D(n8094), .Y(n8108) );
  OA22X1 U9212 ( .A0(\i_MIPS/Register/register[4][9] ), .A1(n5100), .B0(
        \i_MIPS/Register/register[12][9] ), .B1(n5094), .Y(n8096) );
  OA22X1 U9213 ( .A0(\i_MIPS/Register/register[0][9] ), .A1(n5108), .B0(
        \i_MIPS/Register/register[8][9] ), .B1(n5103), .Y(n8095) );
  OAI221XL U9214 ( .A0(\i_MIPS/Register/register[2][9] ), .A1(n5090), .B0(
        \i_MIPS/Register/register[10][9] ), .B1(n5085), .C0(n8089), .Y(n8097)
         );
  NAND4BX1 U9215 ( .AN(n7367), .B(n7366), .C(n7365), .D(n7364), .Y(n7378) );
  OAI221XL U9216 ( .A0(\i_MIPS/Register/register[2][7] ), .A1(n5089), .B0(
        \i_MIPS/Register/register[10][7] ), .B1(n5085), .C0(n7359), .Y(n7367)
         );
  NAND4BX1 U9217 ( .AN(n8014), .B(n8013), .C(n8012), .D(n8011), .Y(n8025) );
  OA22X1 U9218 ( .A0(\i_MIPS/Register/register[4][13] ), .A1(n5100), .B0(
        \i_MIPS/Register/register[12][13] ), .B1(n5094), .Y(n8013) );
  OA22X1 U9219 ( .A0(\i_MIPS/Register/register[0][13] ), .A1(n5108), .B0(
        \i_MIPS/Register/register[8][13] ), .B1(n5103), .Y(n8012) );
  OAI221XL U9220 ( .A0(\i_MIPS/Register/register[2][13] ), .A1(n5090), .B0(
        \i_MIPS/Register/register[10][13] ), .B1(n5085), .C0(n8006), .Y(n8014)
         );
  NAND4BX1 U9221 ( .AN(n7287), .B(n7286), .C(n7285), .D(n7284), .Y(n7298) );
  OA22X1 U9222 ( .A0(\i_MIPS/Register/register[4][6] ), .A1(n5099), .B0(
        \i_MIPS/Register/register[12][6] ), .B1(n5092), .Y(n7286) );
  OA22X1 U9223 ( .A0(\i_MIPS/Register/register[0][6] ), .A1(n5106), .B0(
        \i_MIPS/Register/register[8][6] ), .B1(n5103), .Y(n7285) );
  OAI221XL U9224 ( .A0(\i_MIPS/Register/register[2][6] ), .A1(n5089), .B0(
        \i_MIPS/Register/register[10][6] ), .B1(n5085), .C0(n7279), .Y(n7287)
         );
  NAND4BX1 U9225 ( .AN(n7637), .B(n7636), .C(n7635), .D(n7634), .Y(n7648) );
  OAI221XL U9226 ( .A0(\i_MIPS/Register/register[2][28] ), .A1(n5089), .B0(
        \i_MIPS/Register/register[10][28] ), .B1(n5085), .C0(n7629), .Y(n7637)
         );
  NAND4BX1 U9227 ( .AN(n7012), .B(n7011), .C(n7010), .D(n7009), .Y(n7023) );
  OA22X1 U9228 ( .A0(\i_MIPS/Register/register[4][23] ), .A1(n5099), .B0(
        \i_MIPS/Register/register[12][23] ), .B1(n5092), .Y(n7011) );
  OA22X1 U9229 ( .A0(\i_MIPS/Register/register[0][23] ), .A1(n5106), .B0(
        \i_MIPS/Register/register[8][23] ), .B1(n5103), .Y(n7010) );
  OAI221XL U9230 ( .A0(\i_MIPS/Register/register[2][23] ), .A1(n5089), .B0(
        \i_MIPS/Register/register[10][23] ), .B1(n5084), .C0(n7004), .Y(n7012)
         );
  NAND4BX1 U9231 ( .AN(n7209), .B(n7208), .C(n7207), .D(n7206), .Y(n7220) );
  OA22X1 U9232 ( .A0(\i_MIPS/Register/register[4][2] ), .A1(n5099), .B0(
        \i_MIPS/Register/register[12][2] ), .B1(n5092), .Y(n7208) );
  OA22X1 U9233 ( .A0(\i_MIPS/Register/register[0][2] ), .A1(n5106), .B0(
        \i_MIPS/Register/register[8][2] ), .B1(n5103), .Y(n7207) );
  NAND4BX1 U9234 ( .AN(n6901), .B(n6900), .C(n6899), .D(n6898), .Y(n6912) );
  OA22X1 U9235 ( .A0(\i_MIPS/Register/register[4][29] ), .A1(n5099), .B0(
        \i_MIPS/Register/register[12][29] ), .B1(n5092), .Y(n6900) );
  OA22X1 U9236 ( .A0(\i_MIPS/Register/register[0][29] ), .A1(n5106), .B0(
        \i_MIPS/Register/register[8][29] ), .B1(n5105), .Y(n6899) );
  OAI221XL U9237 ( .A0(\i_MIPS/Register/register[2][29] ), .A1(n5091), .B0(
        \i_MIPS/Register/register[10][29] ), .B1(n5084), .C0(n6893), .Y(n6901)
         );
  NAND4BX1 U9238 ( .AN(n7132), .B(n7131), .C(n7130), .D(n7129), .Y(n7143) );
  OA22X1 U9239 ( .A0(\i_MIPS/Register/register[4][15] ), .A1(n5099), .B0(
        \i_MIPS/Register/register[12][15] ), .B1(n5092), .Y(n7131) );
  OA22X1 U9240 ( .A0(\i_MIPS/Register/register[0][15] ), .A1(n5106), .B0(
        \i_MIPS/Register/register[8][15] ), .B1(n5103), .Y(n7130) );
  OAI221XL U9241 ( .A0(\i_MIPS/Register/register[2][15] ), .A1(n5091), .B0(
        \i_MIPS/Register/register[10][15] ), .B1(n5084), .C0(n7124), .Y(n7132)
         );
  NAND4BX1 U9242 ( .AN(n6801), .B(n6800), .C(n6799), .D(n6798), .Y(n6812) );
  OA22X1 U9243 ( .A0(\i_MIPS/Register/register[4][25] ), .A1(n5099), .B0(
        \i_MIPS/Register/register[12][25] ), .B1(n5092), .Y(n6800) );
  OA22X1 U9244 ( .A0(\i_MIPS/Register/register[0][25] ), .A1(n5106), .B0(
        \i_MIPS/Register/register[8][25] ), .B1(n5105), .Y(n6799) );
  OAI221XL U9245 ( .A0(\i_MIPS/Register/register[2][25] ), .A1(n5089), .B0(
        \i_MIPS/Register/register[10][25] ), .B1(n5084), .C0(n6793), .Y(n6801)
         );
  NAND4BX1 U9246 ( .AN(n7824), .B(n7823), .C(n7822), .D(n7821), .Y(n7835) );
  OAI221XL U9247 ( .A0(\i_MIPS/Register/register[2][14] ), .A1(n5089), .B0(
        \i_MIPS/Register/register[10][14] ), .B1(n5085), .C0(n7816), .Y(n7824)
         );
  NAND4BX1 U9248 ( .AN(n9484), .B(n9483), .C(n9482), .D(n9481), .Y(n9485) );
  OA22XL U9249 ( .A0(\i_MIPS/Register/register[20][30] ), .A1(net107169), .B0(
        \i_MIPS/Register/register[28][30] ), .B1(net107170), .Y(n9483) );
  OA22XL U9250 ( .A0(\i_MIPS/Register/register[16][30] ), .A1(net107167), .B0(
        \i_MIPS/Register/register[24][30] ), .B1(net107168), .Y(n9482) );
  OAI221XL U9251 ( .A0(\i_MIPS/Register/register[18][30] ), .A1(net117643), 
        .B0(\i_MIPS/Register/register[26][30] ), .B1(net117663), .C0(n9476), 
        .Y(n9484) );
  NAND4BX1 U9252 ( .AN(n7762), .B(n7761), .C(n7760), .D(n7759), .Y(n7763) );
  OA22XL U9253 ( .A0(\i_MIPS/Register/register[20][14] ), .A1(net107169), .B0(
        \i_MIPS/Register/register[28][14] ), .B1(net107170), .Y(n7761) );
  OA22XL U9254 ( .A0(\i_MIPS/Register/register[16][14] ), .A1(net107167), .B0(
        \i_MIPS/Register/register[24][14] ), .B1(net107168), .Y(n7760) );
  OAI221XL U9255 ( .A0(\i_MIPS/Register/register[18][14] ), .A1(net117637), 
        .B0(\i_MIPS/Register/register[26][14] ), .B1(net117657), .C0(n7754), 
        .Y(n7762) );
  OAI221XL U9256 ( .A0(\i_MIPS/Register/register[18][17] ), .A1(n5088), .B0(
        \i_MIPS/Register/register[26][17] ), .B1(n5086), .C0(n9282), .Y(n9290)
         );
  OA22X1 U9257 ( .A0(\i_MIPS/Register/register[20][1] ), .A1(n5101), .B0(
        \i_MIPS/Register/register[28][1] ), .B1(n5095), .Y(n9038) );
  OA22X1 U9258 ( .A0(\i_MIPS/Register/register[16][1] ), .A1(n5109), .B0(
        \i_MIPS/Register/register[24][1] ), .B1(n5104), .Y(n9037) );
  OAI221XL U9259 ( .A0(\i_MIPS/Register/register[18][1] ), .A1(n5091), .B0(
        \i_MIPS/Register/register[26][1] ), .B1(n5086), .C0(n9031), .Y(n9039)
         );
  NAND4BX1 U9260 ( .AN(n8276), .B(n8275), .C(n8274), .D(n8273), .Y(n8277) );
  OA22X1 U9261 ( .A0(\i_MIPS/Register/register[20][12] ), .A1(n5100), .B0(
        \i_MIPS/Register/register[28][12] ), .B1(n5094), .Y(n8275) );
  OA22X1 U9262 ( .A0(\i_MIPS/Register/register[16][12] ), .A1(n5108), .B0(
        \i_MIPS/Register/register[24][12] ), .B1(n5103), .Y(n8274) );
  OAI221XL U9263 ( .A0(\i_MIPS/Register/register[18][12] ), .A1(n5090), .B0(
        \i_MIPS/Register/register[26][12] ), .B1(n5085), .C0(n8268), .Y(n8276)
         );
  NAND4BX1 U9264 ( .AN(n8629), .B(n8628), .C(n8627), .D(n8626), .Y(n8630) );
  OA22X1 U9265 ( .A0(\i_MIPS/Register/register[20][18] ), .A1(n5101), .B0(
        \i_MIPS/Register/register[28][18] ), .B1(n5095), .Y(n8628) );
  OA22X1 U9266 ( .A0(\i_MIPS/Register/register[16][18] ), .A1(n5109), .B0(
        \i_MIPS/Register/register[24][18] ), .B1(n5104), .Y(n8627) );
  OAI221XL U9267 ( .A0(\i_MIPS/Register/register[18][18] ), .A1(n5091), .B0(
        \i_MIPS/Register/register[26][18] ), .B1(n4669), .C0(n8621), .Y(n8629)
         );
  OAI221XL U9268 ( .A0(\i_MIPS/Register/register[18][5] ), .A1(n5088), .B0(
        \i_MIPS/Register/register[26][5] ), .B1(n5086), .C0(n9373), .Y(n9381)
         );
  OA22X1 U9269 ( .A0(\i_MIPS/Register/register[20][0] ), .A1(n5101), .B0(
        \i_MIPS/Register/register[28][0] ), .B1(n5095), .Y(n8775) );
  OA22X1 U9270 ( .A0(\i_MIPS/Register/register[16][0] ), .A1(n5109), .B0(
        \i_MIPS/Register/register[24][0] ), .B1(n5104), .Y(n8774) );
  NAND4BX1 U9271 ( .AN(n8547), .B(n8546), .C(n8545), .D(n8544), .Y(n8548) );
  OA22X1 U9272 ( .A0(\i_MIPS/Register/register[20][11] ), .A1(n5101), .B0(
        \i_MIPS/Register/register[28][11] ), .B1(n5095), .Y(n8546) );
  OA22X1 U9273 ( .A0(\i_MIPS/Register/register[16][11] ), .A1(n5109), .B0(
        \i_MIPS/Register/register[24][11] ), .B1(n5104), .Y(n8545) );
  OAI221XL U9274 ( .A0(\i_MIPS/Register/register[18][11] ), .A1(n5091), .B0(
        \i_MIPS/Register/register[26][11] ), .B1(n4669), .C0(n8539), .Y(n8547)
         );
  NAND4BX1 U9275 ( .AN(n8852), .B(n8851), .C(n8850), .D(n8849), .Y(n8853) );
  OA22X1 U9276 ( .A0(\i_MIPS/Register/register[20][16] ), .A1(n5101), .B0(
        \i_MIPS/Register/register[28][16] ), .B1(n5095), .Y(n8851) );
  OA22X1 U9277 ( .A0(\i_MIPS/Register/register[16][16] ), .A1(n5109), .B0(
        \i_MIPS/Register/register[24][16] ), .B1(n5104), .Y(n8850) );
  OAI221XL U9278 ( .A0(\i_MIPS/Register/register[18][16] ), .A1(n5091), .B0(
        \i_MIPS/Register/register[26][16] ), .B1(n5087), .C0(n8844), .Y(n8852)
         );
  NAND4BX1 U9279 ( .AN(n8456), .B(n8455), .C(n8454), .D(n8453), .Y(n8457) );
  OA22X1 U9280 ( .A0(\i_MIPS/Register/register[16][20] ), .A1(n5108), .B0(
        \i_MIPS/Register/register[24][20] ), .B1(n5103), .Y(n8454) );
  OAI221XL U9281 ( .A0(\i_MIPS/Register/register[18][20] ), .A1(n5091), .B0(
        \i_MIPS/Register/register[26][20] ), .B1(n4669), .C0(n8448), .Y(n8456)
         );
  OA22X1 U9282 ( .A0(\i_MIPS/Register/register[20][19] ), .A1(n5100), .B0(
        \i_MIPS/Register/register[28][19] ), .B1(n5094), .Y(n8365) );
  OA22X1 U9283 ( .A0(\i_MIPS/Register/register[16][19] ), .A1(n5108), .B0(
        \i_MIPS/Register/register[24][19] ), .B1(n5103), .Y(n8364) );
  NAND4BX1 U9284 ( .AN(n8955), .B(n8954), .C(n8953), .D(n8952), .Y(n8956) );
  OAI221XL U9285 ( .A0(\i_MIPS/Register/register[18][21] ), .A1(n5091), .B0(
        \i_MIPS/Register/register[26][21] ), .B1(n5086), .C0(n8947), .Y(n8955)
         );
  NAND4BX1 U9286 ( .AN(n8196), .B(n8195), .C(n8194), .D(n8193), .Y(n8197) );
  OA22X1 U9287 ( .A0(\i_MIPS/Register/register[20][8] ), .A1(n5100), .B0(
        \i_MIPS/Register/register[28][8] ), .B1(n5094), .Y(n8195) );
  OA22X1 U9288 ( .A0(\i_MIPS/Register/register[16][8] ), .A1(n5108), .B0(
        \i_MIPS/Register/register[24][8] ), .B1(n5103), .Y(n8194) );
  OAI221XL U9289 ( .A0(\i_MIPS/Register/register[18][8] ), .A1(n5090), .B0(
        \i_MIPS/Register/register[26][8] ), .B1(n5085), .C0(n8188), .Y(n8196)
         );
  OAI221XL U9290 ( .A0(\i_MIPS/Register/register[18][26] ), .A1(n5089), .B0(
        \i_MIPS/Register/register[26][26] ), .B1(n5085), .C0(n7467), .Y(n7475)
         );
  NAND4BX1 U9291 ( .AN(n7560), .B(n7559), .C(n7558), .D(n7557), .Y(n7561) );
  OAI221XL U9292 ( .A0(\i_MIPS/Register/register[18][10] ), .A1(n5089), .B0(
        \i_MIPS/Register/register[26][10] ), .B1(n5085), .C0(n7552), .Y(n7560)
         );
  OA22X1 U9293 ( .A0(\i_MIPS/Register/register[20][4] ), .A1(n5101), .B0(
        \i_MIPS/Register/register[28][4] ), .B1(n5095), .Y(n9114) );
  OA22X1 U9294 ( .A0(\i_MIPS/Register/register[16][4] ), .A1(n5109), .B0(
        \i_MIPS/Register/register[24][4] ), .B1(n5104), .Y(n9113) );
  NAND4BX1 U9295 ( .AN(n8106), .B(n8105), .C(n8104), .D(n8103), .Y(n8107) );
  OA22X1 U9296 ( .A0(\i_MIPS/Register/register[20][9] ), .A1(n5100), .B0(
        \i_MIPS/Register/register[28][9] ), .B1(n5094), .Y(n8105) );
  OA22X1 U9297 ( .A0(\i_MIPS/Register/register[16][9] ), .A1(n5108), .B0(
        \i_MIPS/Register/register[24][9] ), .B1(n5103), .Y(n8104) );
  OAI221XL U9298 ( .A0(\i_MIPS/Register/register[18][9] ), .A1(n5090), .B0(
        \i_MIPS/Register/register[26][9] ), .B1(n5085), .C0(n8098), .Y(n8106)
         );
  NAND4BX1 U9299 ( .AN(n7376), .B(n7375), .C(n7374), .D(n7373), .Y(n7377) );
  OAI221XL U9300 ( .A0(\i_MIPS/Register/register[18][7] ), .A1(n5089), .B0(
        \i_MIPS/Register/register[26][7] ), .B1(n5085), .C0(n7368), .Y(n7376)
         );
  NAND4BX1 U9301 ( .AN(n8023), .B(n8022), .C(n8021), .D(n8020), .Y(n8024) );
  OAI221XL U9302 ( .A0(\i_MIPS/Register/register[18][13] ), .A1(n5090), .B0(
        \i_MIPS/Register/register[26][13] ), .B1(n5085), .C0(n8015), .Y(n8023)
         );
  NAND4BX1 U9303 ( .AN(n7296), .B(n7295), .C(n7294), .D(n7293), .Y(n7297) );
  OAI221XL U9304 ( .A0(\i_MIPS/Register/register[18][6] ), .A1(n5089), .B0(
        \i_MIPS/Register/register[26][6] ), .B1(n5085), .C0(n7288), .Y(n7296)
         );
  OAI221XL U9305 ( .A0(\i_MIPS/Register/register[18][28] ), .A1(n5089), .B0(
        \i_MIPS/Register/register[26][28] ), .B1(n5085), .C0(n7638), .Y(n7646)
         );
  NAND4BX1 U9306 ( .AN(n7021), .B(n7020), .C(n7019), .D(n7018), .Y(n7022) );
  OA22X1 U9307 ( .A0(\i_MIPS/Register/register[20][23] ), .A1(n5099), .B0(
        \i_MIPS/Register/register[28][23] ), .B1(n5092), .Y(n7020) );
  OA22X1 U9308 ( .A0(\i_MIPS/Register/register[16][23] ), .A1(n5106), .B0(
        \i_MIPS/Register/register[24][23] ), .B1(n5105), .Y(n7019) );
  OAI221XL U9309 ( .A0(\i_MIPS/Register/register[18][23] ), .A1(n5089), .B0(
        \i_MIPS/Register/register[26][23] ), .B1(n5084), .C0(n7013), .Y(n7021)
         );
  NAND4BX1 U9310 ( .AN(n7218), .B(n7217), .C(n7216), .D(n7215), .Y(n7219) );
  OA22X1 U9311 ( .A0(\i_MIPS/Register/register[20][2] ), .A1(n5099), .B0(
        \i_MIPS/Register/register[28][2] ), .B1(n5092), .Y(n7217) );
  OA22X1 U9312 ( .A0(\i_MIPS/Register/register[16][2] ), .A1(n5106), .B0(
        \i_MIPS/Register/register[24][2] ), .B1(n5105), .Y(n7216) );
  NAND4BX1 U9313 ( .AN(n6910), .B(n6909), .C(n6908), .D(n6907), .Y(n6911) );
  OA22X1 U9314 ( .A0(\i_MIPS/Register/register[20][29] ), .A1(n5099), .B0(
        \i_MIPS/Register/register[28][29] ), .B1(n5092), .Y(n6909) );
  OA22X1 U9315 ( .A0(\i_MIPS/Register/register[16][29] ), .A1(n5106), .B0(
        \i_MIPS/Register/register[24][29] ), .B1(n5103), .Y(n6908) );
  OAI221XL U9316 ( .A0(\i_MIPS/Register/register[18][29] ), .A1(n5089), .B0(
        \i_MIPS/Register/register[26][29] ), .B1(n5084), .C0(n6902), .Y(n6910)
         );
  NAND4BX1 U9317 ( .AN(n7141), .B(n7140), .C(n7139), .D(n7138), .Y(n7142) );
  OA22X1 U9318 ( .A0(\i_MIPS/Register/register[20][15] ), .A1(n5099), .B0(
        \i_MIPS/Register/register[28][15] ), .B1(n5092), .Y(n7140) );
  OA22X1 U9319 ( .A0(\i_MIPS/Register/register[16][15] ), .A1(n5106), .B0(
        \i_MIPS/Register/register[24][15] ), .B1(n5105), .Y(n7139) );
  OAI221XL U9320 ( .A0(\i_MIPS/Register/register[18][15] ), .A1(n5091), .B0(
        \i_MIPS/Register/register[26][15] ), .B1(n5084), .C0(n7133), .Y(n7141)
         );
  NAND4BX1 U9321 ( .AN(n6810), .B(n6809), .C(n6808), .D(n6807), .Y(n6811) );
  OA22X1 U9322 ( .A0(\i_MIPS/Register/register[20][25] ), .A1(n5099), .B0(
        \i_MIPS/Register/register[28][25] ), .B1(n5092), .Y(n6809) );
  OA22X1 U9323 ( .A0(\i_MIPS/Register/register[16][25] ), .A1(n5106), .B0(
        \i_MIPS/Register/register[24][25] ), .B1(n5103), .Y(n6808) );
  OAI221XL U9324 ( .A0(\i_MIPS/Register/register[18][25] ), .A1(n5089), .B0(
        \i_MIPS/Register/register[26][25] ), .B1(n5084), .C0(n6802), .Y(n6810)
         );
  NAND4BX1 U9325 ( .AN(n7833), .B(n7832), .C(n7831), .D(n7830), .Y(n7834) );
  OAI221XL U9326 ( .A0(\i_MIPS/Register/register[18][14] ), .A1(n5089), .B0(
        \i_MIPS/Register/register[26][14] ), .B1(n5085), .C0(n7825), .Y(n7833)
         );
  NAND3X2 U9327 ( .A(ICACHE_addr[24]), .B(ICACHE_addr[23]), .C(n10385), .Y(
        n10531) );
  INVX1 U9328 ( .A(n7411), .Y(n9450) );
  OAI221XL U9329 ( .A0(\i_MIPS/ALUin1[22] ), .A1(n5072), .B0(
        \i_MIPS/ALUin1[23] ), .B1(n5068), .C0(n6831), .Y(n6832) );
  INVX1 U9330 ( .A(n7674), .Y(n9546) );
  OAI221XL U9331 ( .A0(\i_MIPS/ALUin1[24] ), .A1(n5071), .B0(
        \i_MIPS/ALUin1[25] ), .B1(n5068), .C0(n7673), .Y(n7674) );
  MXI2XL U9332 ( .A(\i_MIPS/n270 ), .B(n3027), .S0(n3601), .Y(\i_MIPS/n461 )
         );
  MXI2XL U9333 ( .A(\i_MIPS/n287 ), .B(n3690), .S0(n3593), .Y(\i_MIPS/n478 )
         );
  MXI2X1 U9334 ( .A(\i_MIPS/n300 ), .B(n4694), .S0(n3597), .Y(\i_MIPS/n491 )
         );
  MXI2XL U9335 ( .A(\i_MIPS/n271 ), .B(n3675), .S0(n3590), .Y(\i_MIPS/n462 )
         );
  MXI2X1 U9336 ( .A(\i_MIPS/n263 ), .B(\i_MIPS/n501 ), .S0(n3597), .Y(
        \i_MIPS/n453 ) );
  MXI2XL U9337 ( .A(\i_MIPS/n260 ), .B(\i_MIPS/n504 ), .S0(n3605), .Y(
        \i_MIPS/n450 ) );
  MXI2XL U9338 ( .A(\i_MIPS/n259 ), .B(\i_MIPS/n505 ), .S0(n3605), .Y(
        \i_MIPS/n449 ) );
  MX2XL U9339 ( .A(\i_MIPS/ALUin1[22] ), .B(n10349), .S0(n3589), .Y(
        \i_MIPS/n470 ) );
  MXI2XL U9340 ( .A(\i_MIPS/n264 ), .B(\i_MIPS/n265 ), .S0(n3590), .Y(
        \i_MIPS/n454 ) );
  MXI2XL U9341 ( .A(\i_MIPS/n266 ), .B(\i_MIPS/n267 ), .S0(n3599), .Y(
        \i_MIPS/n456 ) );
  MX2XL U9342 ( .A(\i_MIPS/ALUin1[2] ), .B(n10825), .S0(n3595), .Y(
        \i_MIPS/n490 ) );
  MX2XL U9343 ( .A(\i_MIPS/ALUin1[3] ), .B(n10768), .S0(n3588), .Y(
        \i_MIPS/n489 ) );
  MX2XL U9344 ( .A(\i_MIPS/ALUin1[4] ), .B(n10933), .S0(n3595), .Y(
        \i_MIPS/n488 ) );
  MX2XL U9345 ( .A(\i_MIPS/ALUin1[5] ), .B(n10910), .S0(n3599), .Y(
        \i_MIPS/n487 ) );
  MX2XL U9346 ( .A(\i_MIPS/ALUin1[6] ), .B(n10868), .S0(n3591), .Y(
        \i_MIPS/n486 ) );
  MX2XL U9347 ( .A(\i_MIPS/ALUin1[7] ), .B(n10686), .S0(n3593), .Y(
        \i_MIPS/n485 ) );
  MX2XL U9348 ( .A(\i_MIPS/ALUin1[9] ), .B(n10618), .S0(n3601), .Y(
        \i_MIPS/n483 ) );
  MX2XL U9349 ( .A(\i_MIPS/ALUin1[10] ), .B(n10528), .S0(n3595), .Y(
        \i_MIPS/n482 ) );
  MX2XL U9350 ( .A(\i_MIPS/ALUin1[11] ), .B(n10796), .S0(n3593), .Y(
        \i_MIPS/n481 ) );
  MX2XL U9351 ( .A(\i_MIPS/ALUin1[12] ), .B(n10473), .S0(n3599), .Y(
        \i_MIPS/n480 ) );
  MX2XL U9352 ( .A(\i_MIPS/ALUin1[13] ), .B(n10811), .S0(n3605), .Y(
        \i_MIPS/n479 ) );
  MX2XL U9353 ( .A(\i_MIPS/ALUin1[15] ), .B(net105236), .S0(n3588), .Y(
        \i_MIPS/n477 ) );
  MX2XL U9354 ( .A(\i_MIPS/ALUin1[16] ), .B(n10511), .S0(n3601), .Y(
        \i_MIPS/n476 ) );
  MX2XL U9355 ( .A(\i_MIPS/ALUin1[19] ), .B(n10978), .S0(n3588), .Y(
        \i_MIPS/n473 ) );
  MX2XL U9356 ( .A(\i_MIPS/ALUin1[20] ), .B(n10416), .S0(n3601), .Y(
        \i_MIPS/n472 ) );
  MX2XL U9357 ( .A(\i_MIPS/ALUin1[21] ), .B(n10526), .S0(n3590), .Y(
        \i_MIPS/n471 ) );
  MX2XL U9358 ( .A(\i_MIPS/ALUin1[24] ), .B(n10429), .S0(n3591), .Y(
        \i_MIPS/n468 ) );
  MX2XL U9359 ( .A(\i_MIPS/ALUin1[25] ), .B(n11055), .S0(n3591), .Y(
        \i_MIPS/n467 ) );
  MX2XL U9360 ( .A(\i_MIPS/ALUin1[26] ), .B(n10443), .S0(n3603), .Y(
        \i_MIPS/n466 ) );
  MX2XL U9361 ( .A(\i_MIPS/ALUin1[27] ), .B(n3888), .S0(n3601), .Y(
        \i_MIPS/n465 ) );
  MX2XL U9362 ( .A(\i_MIPS/ALUin1[28] ), .B(n10554), .S0(n3603), .Y(
        \i_MIPS/n464 ) );
  MX2XL U9363 ( .A(\i_MIPS/ALUin1[29] ), .B(n10569), .S0(n3588), .Y(
        \i_MIPS/n463 ) );
  MX2XL U9364 ( .A(\i_MIPS/ALUin1[8] ), .B(n10659), .S0(n3595), .Y(
        \i_MIPS/n484 ) );
  MX2XL U9365 ( .A(\i_MIPS/ALUin1[17] ), .B(n10631), .S0(n3599), .Y(
        \i_MIPS/n475 ) );
  MX2XL U9366 ( .A(\i_MIPS/ALUin1[18] ), .B(n10646), .S0(n3597), .Y(
        \i_MIPS/n474 ) );
  MX2XL U9367 ( .A(\i_MIPS/ALUin1[23] ), .B(n10698), .S0(n3601), .Y(
        \i_MIPS/n469 ) );
  MXI2XL U9368 ( .A(\i_MIPS/n254 ), .B(\i_MIPS/n253 ), .S0(n3603), .Y(
        \i_MIPS/n414 ) );
  MXI2XL U9369 ( .A(\i_MIPS/n250 ), .B(\i_MIPS/n249 ), .S0(n3588), .Y(
        \i_MIPS/n412 ) );
  MXI2XL U9370 ( .A(\i_MIPS/n252 ), .B(\i_MIPS/n251 ), .S0(n3599), .Y(
        \i_MIPS/n413 ) );
  MXI2X1 U9371 ( .A(\i_MIPS/n237 ), .B(n3559), .S0(n3605), .Y(\i_MIPS/n360 )
         );
  MXI2X1 U9372 ( .A(\i_MIPS/n231 ), .B(\i_MIPS/n232 ), .S0(n3599), .Y(
        \i_MIPS/n354 ) );
  MXI2X1 U9373 ( .A(\i_MIPS/n243 ), .B(n6713), .S0(n3597), .Y(\i_MIPS/n366 )
         );
  MXI2X1 U9374 ( .A(\i_MIPS/n239 ), .B(\i_MIPS/n240 ), .S0(n3588), .Y(
        \i_MIPS/n362 ) );
  MXI2X1 U9375 ( .A(\i_MIPS/n225 ), .B(\i_MIPS/n226 ), .S0(n3591), .Y(
        \i_MIPS/n348 ) );
  MXI2X1 U9376 ( .A(\i_MIPS/n199 ), .B(\i_MIPS/n200 ), .S0(n3599), .Y(
        \i_MIPS/n322 ) );
  MXI2X1 U9377 ( .A(\i_MIPS/n195 ), .B(\i_MIPS/n196 ), .S0(n3603), .Y(
        \i_MIPS/n318 ) );
  MXI2X1 U9378 ( .A(\i_MIPS/n193 ), .B(\i_MIPS/n194 ), .S0(n3597), .Y(
        \i_MIPS/n316 ) );
  MXI2X1 U9379 ( .A(\i_MIPS/n191 ), .B(\i_MIPS/n192 ), .S0(n3601), .Y(
        \i_MIPS/n314 ) );
  MXI2X1 U9380 ( .A(\i_MIPS/n189 ), .B(\i_MIPS/n190 ), .S0(n3591), .Y(
        \i_MIPS/n312 ) );
  MXI2X1 U9381 ( .A(\i_MIPS/n187 ), .B(\i_MIPS/n188 ), .S0(n3593), .Y(
        \i_MIPS/n310 ) );
  MXI2X1 U9382 ( .A(\i_MIPS/n185 ), .B(\i_MIPS/n186 ), .S0(n3599), .Y(
        \i_MIPS/n308 ) );
  MXI2X1 U9383 ( .A(\i_MIPS/n183 ), .B(\i_MIPS/n184 ), .S0(n3590), .Y(
        \i_MIPS/n306 ) );
  MXI2X1 U9384 ( .A(\i_MIPS/n241 ), .B(\i_MIPS/n242 ), .S0(n3589), .Y(
        \i_MIPS/n364 ) );
  MXI2X1 U9385 ( .A(\i_MIPS/n229 ), .B(\i_MIPS/n230 ), .S0(n3605), .Y(
        \i_MIPS/n352 ) );
  MXI2X1 U9386 ( .A(\i_MIPS/n227 ), .B(\i_MIPS/n228 ), .S0(n3590), .Y(
        \i_MIPS/n350 ) );
  MXI2X1 U9387 ( .A(\i_MIPS/n197 ), .B(\i_MIPS/n198 ), .S0(n3599), .Y(
        \i_MIPS/n320 ) );
  NOR3X1 U9388 ( .A(\i_MIPS/Hazard_detection/n8 ), .B(
        \i_MIPS/Hazard_detection/n9 ), .C(\i_MIPS/Hazard_detection/n10 ), .Y(
        \i_MIPS/Hazard_detection/n7 ) );
  XOR2XL U9389 ( .A(\i_MIPS/ID_EX[114] ), .B(\i_MIPS/jump_addr[26] ), .Y(
        \i_MIPS/Hazard_detection/n8 ) );
  XOR2XL U9390 ( .A(\i_MIPS/ID_EX[115] ), .B(n3001), .Y(
        \i_MIPS/Hazard_detection/n10 ) );
  NOR3X1 U9391 ( .A(\i_MIPS/Hazard_detection/n11 ), .B(
        \i_MIPS/Hazard_detection/n12 ), .C(\i_MIPS/Hazard_detection/n13 ), .Y(
        \i_MIPS/Hazard_detection/n4 ) );
  XOR2XL U9392 ( .A(\i_MIPS/ID_EX[115] ), .B(\i_MIPS/jump_addr[22] ), .Y(
        \i_MIPS/Hazard_detection/n13 ) );
  CLKINVX1 U9393 ( .A(\i_MIPS/IF_ID[21] ), .Y(n10513) );
  CLKINVX1 U9394 ( .A(\i_MIPS/IF_ID[22] ), .Y(n10351) );
  CLKINVX1 U9395 ( .A(\i_MIPS/IF_ID[19] ), .Y(n10320) );
  AOI22X1 U9396 ( .A0(n4806), .A1(n10254), .B0(\i_MIPS/Sign_Extend[12] ), .B1(
        \i_MIPS/IF_ID[14] ), .Y(n4802) );
  AOI22X1 U9397 ( .A0(n4823), .A1(n10288), .B0(\i_MIPS/IF_ID[17] ), .B1(n6016), 
        .Y(n4803) );
  AOI21X1 U9398 ( .A0(\i_MIPS/IF_ID[20] ), .A1(\i_MIPS/Sign_Extend[31] ), .B0(
        n4812), .Y(n4804) );
  OA22XL U9399 ( .A0(\i_MIPS/n522 ), .A1(n10721), .B0(\i_MIPS/PC/n33 ), .B1(
        net115799), .Y(n10731) );
  OAI2BB2XL U9400 ( .B0(n3605), .B1(\i_MIPS/n302 ), .A0N(n2899), .A1N(n3588), 
        .Y(\i_MIPS/n458 ) );
  NAND3BX1 U9401 ( .AN(\i_MIPS/control_out[7] ), .B(n5952), .C(
        \i_MIPS/Control/n10 ), .Y(\i_MIPS/control_out[0] ) );
  OAI22XL U9402 ( .A0(n3593), .A1(\i_MIPS/n246 ), .B0(n11587), .B1(n3586), .Y(
        \i_MIPS/n410 ) );
  OAI2BB2XL U9403 ( .B0(n3589), .B1(\i_MIPS/n267 ), .A0N(n428), .A1N(n3593), 
        .Y(\i_MIPS/n457 ) );
  OAI2BB2XL U9404 ( .B0(n3595), .B1(\i_MIPS/n265 ), .A0N(n428), .A1N(n3589), 
        .Y(\i_MIPS/n455 ) );
  NOR2BX1 U9405 ( .AN(\i_MIPS/IF_ID[7] ), .B(\i_MIPS/n516 ), .Y(n4815) );
  AND2X2 U9406 ( .A(\i_MIPS/n508 ), .B(\i_MIPS/n168 ), .Y(n4816) );
  NAND2XL U9407 ( .A(n10354), .B(ICACHE_addr[19]), .Y(n10342) );
  NAND4BX1 U9408 ( .AN(n9190), .B(n9189), .C(n9188), .D(n9187), .Y(net107857)
         );
  AO22X1 U9409 ( .A0(n4807), .A1(n10258), .B0(\i_MIPS/IF_ID[11] ), .B1(
        \i_MIPS/Sign_Extend[9] ), .Y(n10468) );
  OA22X1 U9410 ( .A0(n5333), .A1(n1276), .B0(n5360), .B1(n2908), .Y(n7539) );
  OA22XL U9411 ( .A0(n5329), .A1(n1280), .B0(n5362), .B1(n2912), .Y(n9526) );
  OA22XL U9412 ( .A0(n5335), .A1(n1306), .B0(n5359), .B1(n2944), .Y(n6859) );
  OA22XL U9413 ( .A0(n5335), .A1(n1281), .B0(n5359), .B1(n2913), .Y(n6966) );
  OA22XL U9414 ( .A0(n5335), .A1(n1282), .B0(n5355), .B1(n2914), .Y(n6863) );
  OA22XL U9415 ( .A0(n5335), .A1(n1283), .B0(n5358), .B1(n2915), .Y(n6744) );
  OA22XL U9416 ( .A0(n5335), .A1(n1307), .B0(n5358), .B1(n2945), .Y(n6736) );
  MX2XL U9417 ( .A(\D_cache/cache[7][149] ), .B(n11006), .S0(n5416), .Y(
        \D_cache/n597 ) );
  MX2XL U9418 ( .A(\D_cache/cache[5][149] ), .B(n11006), .S0(n5349), .Y(
        \D_cache/n599 ) );
  MX2XL U9419 ( .A(\D_cache/cache[4][149] ), .B(n11006), .S0(n5321), .Y(
        \D_cache/n600 ) );
  MX2XL U9420 ( .A(\D_cache/cache[3][149] ), .B(n11006), .S0(n5276), .Y(
        \D_cache/n601 ) );
  MX2XL U9421 ( .A(\D_cache/cache[2][149] ), .B(n11006), .S0(n5233), .Y(
        \D_cache/n602 ) );
  MX2XL U9422 ( .A(\D_cache/cache[1][149] ), .B(n11006), .S0(n5207), .Y(
        \D_cache/n603 ) );
  MX2XL U9423 ( .A(\D_cache/cache[0][149] ), .B(n11006), .S0(n5165), .Y(
        \D_cache/n604 ) );
  MX2XL U9424 ( .A(\D_cache/cache[7][143] ), .B(n11035), .S0(n5417), .Y(
        \D_cache/n645 ) );
  MX2XL U9425 ( .A(\D_cache/cache[6][143] ), .B(n11035), .S0(n5373), .Y(
        \D_cache/n646 ) );
  MX2XL U9426 ( .A(\D_cache/cache[5][143] ), .B(n11035), .S0(n5348), .Y(
        \D_cache/n647 ) );
  MX2XL U9427 ( .A(\D_cache/cache[4][143] ), .B(n11035), .S0(n5322), .Y(
        \D_cache/n648 ) );
  MX2XL U9428 ( .A(\D_cache/cache[3][143] ), .B(n11035), .S0(n5270), .Y(
        \D_cache/n649 ) );
  MX2XL U9429 ( .A(\D_cache/cache[2][143] ), .B(n11035), .S0(n5234), .Y(
        \D_cache/n650 ) );
  MX2XL U9430 ( .A(\D_cache/cache[1][143] ), .B(n11035), .S0(n5206), .Y(
        \D_cache/n651 ) );
  MX2XL U9431 ( .A(\D_cache/cache[0][143] ), .B(n11035), .S0(n5166), .Y(
        \D_cache/n652 ) );
  MX2XL U9432 ( .A(\D_cache/cache[7][148] ), .B(n11013), .S0(n5415), .Y(
        \D_cache/n605 ) );
  MX2XL U9433 ( .A(\D_cache/cache[6][148] ), .B(n11013), .S0(n5371), .Y(
        \D_cache/n606 ) );
  MX2XL U9434 ( .A(\D_cache/cache[5][148] ), .B(n11013), .S0(n5347), .Y(
        \D_cache/n607 ) );
  MX2XL U9435 ( .A(\D_cache/cache[4][148] ), .B(n11013), .S0(n5320), .Y(
        \D_cache/n608 ) );
  MX2XL U9436 ( .A(\D_cache/cache[3][148] ), .B(n11013), .S0(n5274), .Y(
        \D_cache/n609 ) );
  MX2XL U9437 ( .A(\D_cache/cache[2][148] ), .B(n11013), .S0(n5233), .Y(
        \D_cache/n610 ) );
  MX2XL U9438 ( .A(\D_cache/cache[1][148] ), .B(n11013), .S0(n5205), .Y(
        \D_cache/n611 ) );
  MX2XL U9439 ( .A(\D_cache/cache[0][148] ), .B(n11013), .S0(n5164), .Y(
        \D_cache/n612 ) );
  MX2XL U9440 ( .A(\D_cache/cache[7][146] ), .B(n11033), .S0(n5417), .Y(
        \D_cache/n621 ) );
  MX2XL U9441 ( .A(\D_cache/cache[6][146] ), .B(n11033), .S0(n5373), .Y(
        \D_cache/n622 ) );
  MX2XL U9442 ( .A(\D_cache/cache[5][146] ), .B(n11033), .S0(n5348), .Y(
        \D_cache/n623 ) );
  MX2XL U9443 ( .A(\D_cache/cache[4][146] ), .B(n11033), .S0(n5322), .Y(
        \D_cache/n624 ) );
  MX2XL U9444 ( .A(\D_cache/cache[3][146] ), .B(n11033), .S0(n5274), .Y(
        \D_cache/n625 ) );
  MX2XL U9445 ( .A(\D_cache/cache[2][146] ), .B(n11033), .S0(n5234), .Y(
        \D_cache/n626 ) );
  MX2XL U9446 ( .A(\D_cache/cache[1][146] ), .B(n11033), .S0(n5206), .Y(
        \D_cache/n627 ) );
  MX2XL U9447 ( .A(\D_cache/cache[0][146] ), .B(n11033), .S0(n5166), .Y(
        \D_cache/n628 ) );
  AND4X1 U9448 ( .A(n6632), .B(n6631), .C(n6630), .D(n6629), .Y(n4826) );
  AO22X1 U9449 ( .A0(n4783), .A1(n4544), .B0(net104801), .B1(n10589), .Y(
        \i_MIPS/N47 ) );
  CLKINVX1 U9450 ( .A(\i_MIPS/n523 ), .Y(n10589) );
  AO22X1 U9451 ( .A0(n4676), .A1(n4545), .B0(net104801), .B1(n10733), .Y(
        \i_MIPS/N48 ) );
  CLKINVX1 U9452 ( .A(\i_MIPS/n522 ), .Y(n10733) );
  OAI222XL U9453 ( .A0(\i_MIPS/n523 ), .A1(n10721), .B0(n3675), .B1(n10736), 
        .C0(\i_MIPS/PC/n32 ), .C1(net115789), .Y(n10588) );
  CLKINVX1 U9454 ( .A(\i_MIPS/n192 ), .Y(n11095) );
  MXI2XL U9455 ( .A(\i_MIPS/n216 ), .B(n3025), .S0(n3601), .Y(\i_MIPS/n339 )
         );
  MX2XL U9456 ( .A(\i_MIPS/ID_EX[76] ), .B(\i_MIPS/Sign_Extend[3] ), .S0(n3601), .Y(\i_MIPS/n445 ) );
  OA22XL U9457 ( .A0(\i_MIPS/Register/register[0][14] ), .A1(net107167), .B0(
        \i_MIPS/Register/register[8][14] ), .B1(net107168), .Y(n7751) );
  OA22XL U9458 ( .A0(\i_MIPS/Register/register[16][31] ), .A1(net107167), .B0(
        \i_MIPS/Register/register[24][31] ), .B1(net107168), .Y(n9592) );
  OA22XL U9459 ( .A0(\i_MIPS/Register/register[0][30] ), .A1(net107167), .B0(
        \i_MIPS/Register/register[8][30] ), .B1(net107168), .Y(n9473) );
  CLKMX2X2 U9460 ( .A(\I_cache/cache[7][153] ), .B(n10939), .S0(n5842), .Y(
        n11614) );
  CLKMX2X2 U9461 ( .A(\I_cache/cache[6][153] ), .B(n10939), .S0(n5885), .Y(
        n11615) );
  CLKMX2X2 U9462 ( .A(\I_cache/cache[5][153] ), .B(n10939), .S0(n4831), .Y(
        n11616) );
  CLKMX2X2 U9463 ( .A(\I_cache/cache[4][153] ), .B(n10939), .S0(n5798), .Y(
        n11617) );
  CLKMX2X2 U9464 ( .A(\I_cache/cache[3][153] ), .B(n10939), .S0(n5667), .Y(
        n11618) );
  CLKMX2X2 U9465 ( .A(\I_cache/cache[2][153] ), .B(n10939), .S0(n5710), .Y(
        n11619) );
  CLKMX2X2 U9466 ( .A(\I_cache/cache[1][153] ), .B(n10939), .S0(n5578), .Y(
        n11620) );
  CLKMX2X2 U9467 ( .A(\I_cache/cache[0][153] ), .B(n10939), .S0(n5623), .Y(
        n11621) );
  OA22X1 U9468 ( .A0(\i_MIPS/Register/register[23][5] ), .A1(net118311), .B0(
        \i_MIPS/Register/register[31][5] ), .B1(net118335), .Y(n9335) );
  OA22X1 U9469 ( .A0(\i_MIPS/Register/register[23][3] ), .A1(net118311), .B0(
        \i_MIPS/Register/register[31][3] ), .B1(net118335), .Y(n9154) );
  OA22X1 U9470 ( .A0(\i_MIPS/Register/register[23][28] ), .A1(net118305), .B0(
        \i_MIPS/Register/register[31][28] ), .B1(net118329), .Y(n7572) );
  OA22X1 U9471 ( .A0(\i_MIPS/Register/register[23][10] ), .A1(net118305), .B0(
        \i_MIPS/Register/register[31][10] ), .B1(net118329), .Y(n7514) );
  OA22X1 U9472 ( .A0(\i_MIPS/Register/register[23][27] ), .A1(net118305), .B0(
        \i_MIPS/Register/register[31][27] ), .B1(net118329), .Y(n7658) );
  OA22X1 U9473 ( .A0(\i_MIPS/Register/register[23][11] ), .A1(net118307), .B0(
        \i_MIPS/Register/register[31][11] ), .B1(net118331), .Y(n8501) );
  OA22X1 U9474 ( .A0(\i_MIPS/Register/register[23][19] ), .A1(net118307), .B0(
        \i_MIPS/Register/register[31][19] ), .B1(net118331), .Y(n8320) );
  OA22X1 U9475 ( .A0(\i_MIPS/Register/register[23][18] ), .A1(net118307), .B0(
        \i_MIPS/Register/register[31][18] ), .B1(net118327), .Y(n8584) );
  OA22X1 U9476 ( .A0(\i_MIPS/Register/register[23][13] ), .A1(net118307), .B0(
        \i_MIPS/Register/register[31][13] ), .B1(net118331), .Y(n7977) );
  OA22X1 U9477 ( .A0(\i_MIPS/Register/register[23][12] ), .A1(net118307), .B0(
        \i_MIPS/Register/register[31][12] ), .B1(net118331), .Y(n8230) );
  OA22X1 U9478 ( .A0(\i_MIPS/Register/register[23][8] ), .A1(net118307), .B0(
        \i_MIPS/Register/register[31][8] ), .B1(net118331), .Y(n8150) );
  OA22X1 U9479 ( .A0(\i_MIPS/Register/register[23][9] ), .A1(net118307), .B0(
        \i_MIPS/Register/register[31][9] ), .B1(net118331), .Y(n8059) );
  OA22X1 U9480 ( .A0(\i_MIPS/Register/register[23][0] ), .A1(net118307), .B0(
        \i_MIPS/Register/register[31][0] ), .B1(net118327), .Y(n8730) );
  OA22X1 U9481 ( .A0(\i_MIPS/Register/register[23][1] ), .A1(net118303), .B0(
        \i_MIPS/Register/register[31][1] ), .B1(net118327), .Y(n8993) );
  OA22X1 U9482 ( .A0(\i_MIPS/Register/register[23][16] ), .A1(net118311), .B0(
        \i_MIPS/Register/register[31][16] ), .B1(net118327), .Y(n8806) );
  OA22X1 U9483 ( .A0(\i_MIPS/Register/register[23][23] ), .A1(net118303), .B0(
        \i_MIPS/Register/register[31][23] ), .B1(net118327), .Y(n7088) );
  OA22X1 U9484 ( .A0(\i_MIPS/Register/register[23][25] ), .A1(net118303), .B0(
        \i_MIPS/Register/register[31][25] ), .B1(net118327), .Y(n6881) );
  OA22X1 U9485 ( .A0(\i_MIPS/Register/register[23][29] ), .A1(net118303), .B0(
        \i_MIPS/Register/register[31][29] ), .B1(net118327), .Y(n6992) );
  OA22X1 U9486 ( .A0(\i_MIPS/Register/register[23][24] ), .A1(net118303), .B0(
        \i_MIPS/Register/register[31][24] ), .B1(net118327), .Y(n6781) );
  OA22X1 U9487 ( .A0(\i_MIPS/Register/register[23][2] ), .A1(net118303), .B0(
        \i_MIPS/Register/register[31][2] ), .B1(net118327), .Y(n7174) );
  OA22X1 U9488 ( .A0(n5927), .A1(n1785), .B0(n5871), .B1(n3473), .Y(n6543) );
  OA22X1 U9489 ( .A0(n5896), .A1(n1786), .B0(n5854), .B1(n3474), .Y(n6538) );
  OA22X1 U9490 ( .A0(n5927), .A1(n1787), .B0(n5873), .B1(n3475), .Y(n6530) );
  OA22X1 U9491 ( .A0(n5896), .A1(n1788), .B0(n5871), .B1(n3476), .Y(n6534) );
  OA22X1 U9492 ( .A0(n5914), .A1(n1529), .B0(n5872), .B1(n3216), .Y(n10813) );
  OA22X1 U9493 ( .A0(n5897), .A1(n1789), .B0(n5855), .B1(n3477), .Y(n6548) );
  OA22X1 U9494 ( .A0(n5897), .A1(n1790), .B0(n5855), .B1(n3478), .Y(n6553) );
  OA22X1 U9495 ( .A0(n5914), .A1(n1530), .B0(n5872), .B1(n3217), .Y(n10818) );
  OA22X1 U9496 ( .A0(n5910), .A1(n1531), .B0(n5868), .B1(n3218), .Y(n10039) );
  OA22X1 U9497 ( .A0(n5910), .A1(n1791), .B0(n5868), .B1(n3479), .Y(n10029) );
  OA22X1 U9498 ( .A0(n5910), .A1(n1792), .B0(n5868), .B1(n3480), .Y(n10034) );
  OA22X1 U9499 ( .A0(n5910), .A1(n1532), .B0(n5868), .B1(n3219), .Y(n10044) );
  OA22X1 U9500 ( .A0(n5914), .A1(n1533), .B0(n5872), .B1(n3220), .Y(n10834) );
  OA22X1 U9501 ( .A0(n5914), .A1(n1793), .B0(n5872), .B1(n3481), .Y(n10829) );
  OA22X1 U9502 ( .A0(n5914), .A1(n1534), .B0(n5872), .B1(n3221), .Y(n10839) );
  OA22X1 U9503 ( .A0(n5909), .A1(n1535), .B0(n5867), .B1(n3222), .Y(n10017) );
  OA22X1 U9504 ( .A0(n5909), .A1(n1794), .B0(n5867), .B1(n3482), .Y(n10007) );
  OA22X1 U9505 ( .A0(n5909), .A1(n1795), .B0(n5867), .B1(n3483), .Y(n10012) );
  OA22X1 U9506 ( .A0(n5909), .A1(n1536), .B0(n5867), .B1(n3223), .Y(n10022) );
  OA22X1 U9507 ( .A0(n5908), .A1(n1537), .B0(n5866), .B1(n3224), .Y(n9973) );
  OA22X1 U9508 ( .A0(n5908), .A1(n1796), .B0(n5866), .B1(n3484), .Y(n9963) );
  OA22X1 U9509 ( .A0(n5908), .A1(n1797), .B0(n5866), .B1(n3485), .Y(n9968) );
  OA22X1 U9510 ( .A0(n5908), .A1(n1538), .B0(n5866), .B1(n3225), .Y(n9978) );
  OA22X1 U9511 ( .A0(n5909), .A1(n1539), .B0(n5867), .B1(n3226), .Y(n9995) );
  OA22X1 U9512 ( .A0(n5908), .A1(n1798), .B0(n5866), .B1(n3486), .Y(n9985) );
  OA22X1 U9513 ( .A0(n5908), .A1(n1799), .B0(n5866), .B1(n3487), .Y(n9990) );
  OA22X1 U9514 ( .A0(n5909), .A1(n1540), .B0(n5867), .B1(n3227), .Y(n10000) );
  OA22X1 U9515 ( .A0(n5904), .A1(n1541), .B0(n5862), .B1(n3228), .Y(n9784) );
  OA22X1 U9516 ( .A0(n5904), .A1(n1800), .B0(n5862), .B1(n3488), .Y(n9774) );
  OA22X1 U9517 ( .A0(n5904), .A1(n1801), .B0(n5862), .B1(n3489), .Y(n9779) );
  OA22X1 U9518 ( .A0(n5904), .A1(n1542), .B0(n5862), .B1(n3229), .Y(n9789) );
  OA22XL U9519 ( .A0(n5917), .A1(n1599), .B0(n5875), .B1(n3286), .Y(n11081) );
  OA22XL U9520 ( .A0(n5917), .A1(n1854), .B0(n5875), .B1(n3541), .Y(n11069) );
  OA22XL U9521 ( .A0(n5917), .A1(n1855), .B0(n5875), .B1(n3542), .Y(n11075) );
  OA22XL U9522 ( .A0(n5917), .A1(n1600), .B0(n5875), .B1(n3287), .Y(n11087) );
  OA22X1 U9523 ( .A0(n5903), .A1(n1543), .B0(n5861), .B1(n3230), .Y(net106695)
         );
  OA22X1 U9524 ( .A0(n5903), .A1(n1802), .B0(n5861), .B1(n3490), .Y(net106721)
         );
  OA22X1 U9525 ( .A0(n5903), .A1(n1803), .B0(n5861), .B1(n3491), .Y(net106708)
         );
  OA22X1 U9526 ( .A0(n5903), .A1(n1544), .B0(n5861), .B1(n3231), .Y(net106682)
         );
  OA22X1 U9527 ( .A0(n5902), .A1(n1344), .B0(n5860), .B1(n3232), .Y(n9736) );
  OA22X1 U9528 ( .A0(n5897), .A1(n1804), .B0(n5855), .B1(n3492), .Y(n6563) );
  OA22X1 U9529 ( .A0(n5897), .A1(n1805), .B0(n5855), .B1(n3493), .Y(n6568) );
  OA22X1 U9530 ( .A0(n5902), .A1(n1545), .B0(n5860), .B1(n3233), .Y(n9741) );
  OA22X1 U9531 ( .A0(n5903), .A1(n1546), .B0(n5861), .B1(n3234), .Y(n9758) );
  OA22X1 U9532 ( .A0(n5902), .A1(n1806), .B0(n5860), .B1(n3494), .Y(n9748) );
  OA22X1 U9533 ( .A0(n5902), .A1(n1807), .B0(n5860), .B1(n3495), .Y(n9753) );
  OA22X1 U9534 ( .A0(n5903), .A1(n1547), .B0(n5861), .B1(n3235), .Y(n9763) );
  OA22X1 U9535 ( .A0(n5911), .A1(n1548), .B0(n5869), .B1(n3236), .Y(n10063) );
  OA22X1 U9536 ( .A0(n5910), .A1(n1808), .B0(n5868), .B1(n3496), .Y(n10053) );
  OA22X1 U9537 ( .A0(n5910), .A1(n1809), .B0(n5868), .B1(n3497), .Y(n10058) );
  OA22X1 U9538 ( .A0(n5911), .A1(n1549), .B0(n5869), .B1(n3237), .Y(n10068) );
  OA22X1 U9539 ( .A0(n5913), .A1(n1550), .B0(n5871), .B1(n3238), .Y(n10242) );
  OA22X1 U9540 ( .A0(n5913), .A1(n1810), .B0(n5871), .B1(n3498), .Y(n10232) );
  OA22X1 U9541 ( .A0(n5913), .A1(n1811), .B0(n5871), .B1(n3499), .Y(n10237) );
  OA22X1 U9542 ( .A0(n5913), .A1(n1551), .B0(n5871), .B1(n3239), .Y(n10247) );
  OA22X1 U9543 ( .A0(n5913), .A1(n1552), .B0(n5871), .B1(n3240), .Y(n10220) );
  OA22X1 U9544 ( .A0(n5912), .A1(n1812), .B0(n5870), .B1(n3500), .Y(n10210) );
  OA22X1 U9545 ( .A0(n5912), .A1(n1813), .B0(n5870), .B1(n3501), .Y(n10215) );
  OA22X1 U9546 ( .A0(n5913), .A1(n1553), .B0(n5871), .B1(n3241), .Y(n10225) );
  OA22X1 U9547 ( .A0(n5912), .A1(n1554), .B0(n5870), .B1(n3242), .Y(n10122) );
  OA22X1 U9548 ( .A0(n5912), .A1(n1814), .B0(n5870), .B1(n3502), .Y(n10112) );
  OA22X1 U9549 ( .A0(n5912), .A1(n1815), .B0(n5870), .B1(n3503), .Y(n10117) );
  OA22X1 U9550 ( .A0(n5912), .A1(n1555), .B0(n5870), .B1(n3243), .Y(n10127) );
  OA22X1 U9551 ( .A0(n5911), .A1(n1556), .B0(n5869), .B1(n3244), .Y(n10086) );
  OA22X1 U9552 ( .A0(n5911), .A1(n1816), .B0(n5869), .B1(n3504), .Y(n10076) );
  OA22X1 U9553 ( .A0(n5911), .A1(n1817), .B0(n5869), .B1(n3505), .Y(n10081) );
  OA22X1 U9554 ( .A0(n5911), .A1(n1557), .B0(n5869), .B1(n3245), .Y(n10091) );
  OA22X1 U9555 ( .A0(n5905), .A1(n1558), .B0(n5863), .B1(n3246), .Y(n9835) );
  OA22X1 U9556 ( .A0(n5904), .A1(n1818), .B0(n5862), .B1(n3506), .Y(n9825) );
  OA22X1 U9557 ( .A0(n5904), .A1(n1819), .B0(n5862), .B1(n3507), .Y(n9830) );
  OA22X1 U9558 ( .A0(n5905), .A1(n1559), .B0(n5863), .B1(n3247), .Y(n9840) );
  OA22X1 U9559 ( .A0(n5906), .A1(n1560), .B0(n5864), .B1(n3248), .Y(n9879) );
  OA22X1 U9560 ( .A0(n5906), .A1(n1820), .B0(n5864), .B1(n3508), .Y(n9869) );
  OA22X1 U9561 ( .A0(n5906), .A1(n1821), .B0(n5864), .B1(n3509), .Y(n9874) );
  OA22X1 U9562 ( .A0(n5906), .A1(n1561), .B0(n5864), .B1(n3249), .Y(n9884) );
  OA22X1 U9563 ( .A0(n5905), .A1(n1562), .B0(n5863), .B1(n3250), .Y(n9857) );
  OA22X1 U9564 ( .A0(n5905), .A1(n1822), .B0(n5863), .B1(n3510), .Y(n9847) );
  OA22X1 U9565 ( .A0(n5905), .A1(n1823), .B0(n5863), .B1(n3511), .Y(n9852) );
  OA22X1 U9566 ( .A0(n5905), .A1(n1563), .B0(n5863), .B1(n3251), .Y(n9862) );
  OA22X1 U9567 ( .A0(n5907), .A1(n1564), .B0(n5865), .B1(n3252), .Y(n9901) );
  OA22X1 U9568 ( .A0(n5906), .A1(n1824), .B0(n5864), .B1(n3512), .Y(n9891) );
  OA22X1 U9569 ( .A0(n5906), .A1(n1825), .B0(n5864), .B1(n3513), .Y(n9896) );
  OA22X1 U9570 ( .A0(n5907), .A1(n1565), .B0(n5865), .B1(n3253), .Y(n9906) );
  OA22X1 U9571 ( .A0(n5907), .A1(n1566), .B0(n5865), .B1(n3254), .Y(n9923) );
  OA22X1 U9572 ( .A0(n5907), .A1(n1826), .B0(n5865), .B1(n3514), .Y(n9913) );
  OA22X1 U9573 ( .A0(n5907), .A1(n1827), .B0(n5865), .B1(n3515), .Y(n9918) );
  OA22X1 U9574 ( .A0(n5907), .A1(n1567), .B0(n5865), .B1(n3255), .Y(n9928) );
  OA22X1 U9575 ( .A0(n5902), .A1(n1568), .B0(n5860), .B1(n3256), .Y(n9716) );
  OA22X1 U9576 ( .A0(n5901), .A1(n1828), .B0(n5859), .B1(n3516), .Y(n9706) );
  OA22X1 U9577 ( .A0(n5901), .A1(n1829), .B0(n5859), .B1(n3517), .Y(n9711) );
  OA22X1 U9578 ( .A0(n5902), .A1(n1569), .B0(n5860), .B1(n3257), .Y(n9721) );
  OA22X1 U9579 ( .A0(n5915), .A1(n1570), .B0(n5873), .B1(n3258), .Y(n10856) );
  OA22X1 U9580 ( .A0(n5914), .A1(n1830), .B0(n5872), .B1(n3518), .Y(n10851) );
  OA22X1 U9581 ( .A0(n5915), .A1(n1571), .B0(n5873), .B1(n3259), .Y(n10861) );
  OA22X1 U9582 ( .A0(n5916), .A1(n1572), .B0(n5874), .B1(n3260), .Y(n10950) );
  OA22X1 U9583 ( .A0(n5916), .A1(n1831), .B0(n5874), .B1(n3519), .Y(n10940) );
  OA22X1 U9584 ( .A0(n5916), .A1(n1832), .B0(n5874), .B1(n3520), .Y(n10945) );
  OA22X1 U9585 ( .A0(n5916), .A1(n1573), .B0(n5874), .B1(n3261), .Y(n10955) );
  OA22X1 U9586 ( .A0(n5916), .A1(n1574), .B0(n5874), .B1(n3262), .Y(n10921) );
  OA22X1 U9587 ( .A0(n5915), .A1(n1833), .B0(n5873), .B1(n3521), .Y(n10916) );
  OA22X1 U9588 ( .A0(n5916), .A1(n1575), .B0(n5874), .B1(n3263), .Y(n10926) );
  OA22X1 U9589 ( .A0(n5915), .A1(n1576), .B0(n5873), .B1(n3288), .Y(n10879) );
  OA22X1 U9590 ( .A0(n5915), .A1(n1834), .B0(n5873), .B1(n3522), .Y(n10874) );
  OA22X1 U9591 ( .A0(n5915), .A1(n1577), .B0(n5873), .B1(n3264), .Y(n10884) );
  OA22X1 U9592 ( .A0(n5898), .A1(n1578), .B0(n5856), .B1(n3265), .Y(n6583) );
  OA22X1 U9593 ( .A0(n5897), .A1(n1835), .B0(n5855), .B1(n3523), .Y(n6573) );
  OA22X1 U9594 ( .A0(n5897), .A1(n1836), .B0(n5855), .B1(n3524), .Y(n6578) );
  OA22X1 U9595 ( .A0(n5900), .A1(n1579), .B0(n5858), .B1(n3266), .Y(n9672) );
  OA22X1 U9596 ( .A0(n5900), .A1(n1837), .B0(n5858), .B1(n3525), .Y(n9662) );
  OA22X1 U9597 ( .A0(n5900), .A1(n1838), .B0(n5858), .B1(n3526), .Y(n9667) );
  OA22X1 U9598 ( .A0(n5900), .A1(n1580), .B0(n5858), .B1(n3267), .Y(n9677) );
  OA22X1 U9599 ( .A0(n5901), .A1(n1581), .B0(n5859), .B1(n3268), .Y(n9694) );
  OA22X1 U9600 ( .A0(n5901), .A1(n1839), .B0(n5859), .B1(n3527), .Y(n9684) );
  OA22X1 U9601 ( .A0(n5901), .A1(n1840), .B0(n5859), .B1(n3528), .Y(n9689) );
  OA22X1 U9602 ( .A0(n5901), .A1(n1582), .B0(n5859), .B1(n3269), .Y(n9699) );
  OA22X1 U9603 ( .A0(n5899), .A1(n1583), .B0(n5857), .B1(n3270), .Y(n9642) );
  OA22X1 U9604 ( .A0(n5899), .A1(n1841), .B0(n5857), .B1(n3529), .Y(n9632) );
  OA22X1 U9605 ( .A0(n5899), .A1(n1842), .B0(n5857), .B1(n3530), .Y(n9637) );
  OA22X1 U9606 ( .A0(n5900), .A1(n1584), .B0(n5858), .B1(n3271), .Y(n9647) );
  OA22X1 U9607 ( .A0(n5899), .A1(n1585), .B0(n5857), .B1(n3272), .Y(n9620) );
  OA22X1 U9608 ( .A0(n5898), .A1(n1843), .B0(n5856), .B1(n3531), .Y(n9610) );
  OA22X1 U9609 ( .A0(n5899), .A1(n1844), .B0(n5857), .B1(n3532), .Y(n9615) );
  OA22X1 U9610 ( .A0(n5899), .A1(n1586), .B0(n5857), .B1(n3273), .Y(n9625) );
  OA22X1 U9611 ( .A0(n5898), .A1(n1587), .B0(n5856), .B1(n3274), .Y(n6598) );
  OA22X1 U9612 ( .A0(n5898), .A1(n1845), .B0(n5856), .B1(n3533), .Y(n6588) );
  OA22X1 U9613 ( .A0(n5898), .A1(n1846), .B0(n5856), .B1(n3534), .Y(n6593) );
  OA22X1 U9614 ( .A0(n5898), .A1(n1588), .B0(n5856), .B1(n3275), .Y(n6603) );
  OA22XL U9615 ( .A0(\i_MIPS/Register/register[4][14] ), .A1(net107169), .B0(
        \i_MIPS/Register/register[12][14] ), .B1(net107170), .Y(n7752) );
  OA22XL U9616 ( .A0(\i_MIPS/Register/register[20][31] ), .A1(net107169), .B0(
        \i_MIPS/Register/register[28][31] ), .B1(net107170), .Y(n9593) );
  OA22XL U9617 ( .A0(\i_MIPS/Register/register[4][30] ), .A1(net107169), .B0(
        \i_MIPS/Register/register[12][30] ), .B1(net107170), .Y(n9474) );
  AO22X1 U9618 ( .A0(n5556), .A1(n4071), .B0(n11054), .B1(
        \i_MIPS/Sign_Extend[12] ), .Y(n10493) );
  OA22X1 U9619 ( .A0(\i_MIPS/Register/register[16][3] ), .A1(n5108), .B0(
        \i_MIPS/Register/register[24][3] ), .B1(n5105), .Y(n9197) );
  OA22X1 U9620 ( .A0(\i_MIPS/Register/register[0][3] ), .A1(n5107), .B0(
        \i_MIPS/Register/register[8][3] ), .B1(n5105), .Y(n9188) );
  OA22XL U9621 ( .A0(\i_MIPS/Register/register[19][22] ), .A1(n7889), .B0(
        \i_MIPS/Register/register[27][22] ), .B1(n7888), .Y(n7893) );
  OA22XL U9622 ( .A0(\i_MIPS/Register/register[3][22] ), .A1(n7889), .B0(
        \i_MIPS/Register/register[11][22] ), .B1(n7888), .Y(n7876) );
  OA22X1 U9623 ( .A0(\i_MIPS/Register/register[19][28] ), .A1(net118353), .B0(
        \i_MIPS/Register/register[27][28] ), .B1(net118381), .Y(n7573) );
  OA22X1 U9624 ( .A0(\i_MIPS/Register/register[3][28] ), .A1(net118353), .B0(
        \i_MIPS/Register/register[11][28] ), .B1(net118379), .Y(n7564) );
  OA22X1 U9625 ( .A0(\i_MIPS/Register/register[19][10] ), .A1(net118353), .B0(
        \i_MIPS/Register/register[27][10] ), .B1(net118379), .Y(n7515) );
  OA22X1 U9626 ( .A0(\i_MIPS/Register/register[3][10] ), .A1(net118353), .B0(
        \i_MIPS/Register/register[11][10] ), .B1(net118379), .Y(n7506) );
  OA22X1 U9627 ( .A0(\i_MIPS/Register/register[19][27] ), .A1(net118353), .B0(
        \i_MIPS/Register/register[27][27] ), .B1(net118379), .Y(n7659) );
  OA22X1 U9628 ( .A0(\i_MIPS/Register/register[3][27] ), .A1(net118353), .B0(
        \i_MIPS/Register/register[11][27] ), .B1(net118375), .Y(n7650) );
  OA22X1 U9629 ( .A0(\i_MIPS/Register/register[19][11] ), .A1(net118357), .B0(
        \i_MIPS/Register/register[27][11] ), .B1(net118381), .Y(n8502) );
  OA22X1 U9630 ( .A0(\i_MIPS/Register/register[3][11] ), .A1(net118355), .B0(
        \i_MIPS/Register/register[11][11] ), .B1(net118379), .Y(n8493) );
  OA22X1 U9631 ( .A0(\i_MIPS/Register/register[19][19] ), .A1(net118355), .B0(
        \i_MIPS/Register/register[27][19] ), .B1(net118379), .Y(n8321) );
  OA22X1 U9632 ( .A0(\i_MIPS/Register/register[3][19] ), .A1(net118355), .B0(
        \i_MIPS/Register/register[11][19] ), .B1(net118379), .Y(n8312) );
  OA22X1 U9633 ( .A0(\i_MIPS/Register/register[19][18] ), .A1(net118357), .B0(
        \i_MIPS/Register/register[27][18] ), .B1(net118381), .Y(n8585) );
  OA22X1 U9634 ( .A0(\i_MIPS/Register/register[3][18] ), .A1(net118357), .B0(
        \i_MIPS/Register/register[11][18] ), .B1(net118381), .Y(n8576) );
  OA22X1 U9635 ( .A0(\i_MIPS/Register/register[19][13] ), .A1(net118355), .B0(
        \i_MIPS/Register/register[27][13] ), .B1(net118379), .Y(n7978) );
  OA22X1 U9636 ( .A0(\i_MIPS/Register/register[3][13] ), .A1(net118355), .B0(
        \i_MIPS/Register/register[11][13] ), .B1(net118379), .Y(n7969) );
  OA22X1 U9637 ( .A0(\i_MIPS/Register/register[19][12] ), .A1(net118355), .B0(
        \i_MIPS/Register/register[27][12] ), .B1(net118379), .Y(n8231) );
  OA22X1 U9638 ( .A0(\i_MIPS/Register/register[3][12] ), .A1(net118355), .B0(
        \i_MIPS/Register/register[11][12] ), .B1(net118379), .Y(n8222) );
  OA22X1 U9639 ( .A0(\i_MIPS/Register/register[19][8] ), .A1(net118355), .B0(
        \i_MIPS/Register/register[27][8] ), .B1(net118379), .Y(n8151) );
  OA22X1 U9640 ( .A0(\i_MIPS/Register/register[3][8] ), .A1(net118355), .B0(
        \i_MIPS/Register/register[11][8] ), .B1(net118379), .Y(n8142) );
  OA22X1 U9641 ( .A0(\i_MIPS/Register/register[19][9] ), .A1(net118355), .B0(
        \i_MIPS/Register/register[27][9] ), .B1(net118379), .Y(n8060) );
  OA22X1 U9642 ( .A0(\i_MIPS/Register/register[3][9] ), .A1(net118355), .B0(
        \i_MIPS/Register/register[11][9] ), .B1(net118379), .Y(n8051) );
  OA22X1 U9643 ( .A0(\i_MIPS/Register/register[19][5] ), .A1(net118359), .B0(
        \i_MIPS/Register/register[27][5] ), .B1(net118379), .Y(n9336) );
  OA22X1 U9644 ( .A0(\i_MIPS/Register/register[3][5] ), .A1(net118359), .B0(
        \i_MIPS/Register/register[11][5] ), .B1(net118379), .Y(n9327) );
  OA22X1 U9645 ( .A0(\i_MIPS/Register/register[19][3] ), .A1(net118359), .B0(
        \i_MIPS/Register/register[27][3] ), .B1(net118379), .Y(n9155) );
  OA22X1 U9646 ( .A0(\i_MIPS/Register/register[3][3] ), .A1(net118359), .B0(
        \i_MIPS/Register/register[11][3] ), .B1(net118379), .Y(n9146) );
  OA22X1 U9647 ( .A0(\i_MIPS/Register/register[3][21] ), .A1(net118357), .B0(
        \i_MIPS/Register/register[11][21] ), .B1(net118381), .Y(n8900) );
  OA22X1 U9648 ( .A0(\i_MIPS/Register/register[19][0] ), .A1(net118357), .B0(
        \i_MIPS/Register/register[27][0] ), .B1(net118381), .Y(n8731) );
  OA22X1 U9649 ( .A0(\i_MIPS/Register/register[3][0] ), .A1(net118357), .B0(
        \i_MIPS/Register/register[11][0] ), .B1(net118381), .Y(n8722) );
  OA22X1 U9650 ( .A0(\i_MIPS/Register/register[19][1] ), .A1(net118357), .B0(
        \i_MIPS/Register/register[27][1] ), .B1(net118381), .Y(n8994) );
  OA22X1 U9651 ( .A0(\i_MIPS/Register/register[3][1] ), .A1(net118357), .B0(
        \i_MIPS/Register/register[11][1] ), .B1(net118381), .Y(n8985) );
  OA22X1 U9652 ( .A0(\i_MIPS/Register/register[19][16] ), .A1(net118357), .B0(
        \i_MIPS/Register/register[27][16] ), .B1(net118381), .Y(n8807) );
  OA22X1 U9653 ( .A0(\i_MIPS/Register/register[3][16] ), .A1(net118357), .B0(
        \i_MIPS/Register/register[11][16] ), .B1(net118381), .Y(n8798) );
  OA22X1 U9654 ( .A0(\i_MIPS/Register/register[19][23] ), .A1(net118351), .B0(
        \i_MIPS/Register/register[27][23] ), .B1(net118375), .Y(n7089) );
  OA22X1 U9655 ( .A0(\i_MIPS/Register/register[3][23] ), .A1(net118351), .B0(
        \i_MIPS/Register/register[11][23] ), .B1(net118375), .Y(n7080) );
  OA22X1 U9656 ( .A0(\i_MIPS/Register/register[19][25] ), .A1(net118351), .B0(
        \i_MIPS/Register/register[27][25] ), .B1(net118375), .Y(n6882) );
  OA22X1 U9657 ( .A0(\i_MIPS/Register/register[3][25] ), .A1(net118351), .B0(
        \i_MIPS/Register/register[11][25] ), .B1(net118375), .Y(n6873) );
  OA22X1 U9658 ( .A0(\i_MIPS/Register/register[19][29] ), .A1(net118351), .B0(
        \i_MIPS/Register/register[27][29] ), .B1(net118375), .Y(n6993) );
  OA22X1 U9659 ( .A0(\i_MIPS/Register/register[3][29] ), .A1(net118351), .B0(
        \i_MIPS/Register/register[11][29] ), .B1(net118375), .Y(n6984) );
  OA22X1 U9660 ( .A0(\i_MIPS/Register/register[19][24] ), .A1(net118351), .B0(
        \i_MIPS/Register/register[27][24] ), .B1(net118375), .Y(n6782) );
  OA22X1 U9661 ( .A0(\i_MIPS/Register/register[3][24] ), .A1(net118351), .B0(
        \i_MIPS/Register/register[11][24] ), .B1(net118375), .Y(n6772) );
  OA22X1 U9662 ( .A0(\i_MIPS/Register/register[3][6] ), .A1(net118351), .B0(
        \i_MIPS/Register/register[11][6] ), .B1(net118375), .Y(n7241) );
  OA22X1 U9663 ( .A0(\i_MIPS/Register/register[19][2] ), .A1(net118351), .B0(
        \i_MIPS/Register/register[27][2] ), .B1(net118375), .Y(n7175) );
  OA22X1 U9664 ( .A0(\i_MIPS/Register/register[3][2] ), .A1(net118351), .B0(
        \i_MIPS/Register/register[11][2] ), .B1(net118375), .Y(n7166) );
  OA22X1 U9665 ( .A0(n5330), .A1(n1277), .B0(n5355), .B1(n2909), .Y(n8344) );
  OA22XL U9666 ( .A0(n5329), .A1(n1235), .B0(n5354), .B1(n2857), .Y(n8242) );
  OA22XL U9667 ( .A0(n5329), .A1(n1236), .B0(n5354), .B1(n2858), .Y(n8170) );
  OA22XL U9668 ( .A0(n5329), .A1(n1237), .B0(n5354), .B1(n2859), .Y(n8162) );
  OA22XL U9669 ( .A0(n5335), .A1(n1284), .B0(n5359), .B1(n2916), .Y(n6970) );
  OA22XL U9670 ( .A0(n5335), .A1(n1285), .B0(n5359), .B1(n2917), .Y(n6748) );
  OA22XL U9671 ( .A0(n5335), .A1(n1308), .B0(n5359), .B1(n2946), .Y(n6855) );
  OA22XL U9672 ( .A0(n5335), .A1(n1309), .B0(n5359), .B1(n2947), .Y(n6740) );
  AO22X1 U9673 ( .A0(net118235), .A1(n834), .B0(net118253), .B1(n2453), .Y(
        n8325) );
  AO22X1 U9674 ( .A0(net118235), .A1(n835), .B0(net118253), .B1(n2454), .Y(
        n8316) );
  AO22X1 U9675 ( .A0(n5158), .A1(n836), .B0(n5153), .B1(n2455), .Y(n9032) );
  AO22X1 U9676 ( .A0(n5158), .A1(n837), .B0(n5153), .B1(n2456), .Y(n9023) );
  AO22X1 U9677 ( .A0(net118237), .A1(n838), .B0(net118255), .B1(n2457), .Y(
        n8735) );
  AO22X1 U9678 ( .A0(net118237), .A1(n839), .B0(net118255), .B1(n2458), .Y(
        n8726) );
  AO22X1 U9679 ( .A0(net118239), .A1(n204), .B0(net118261), .B1(n931), .Y(
        n8998) );
  AO22X1 U9680 ( .A0(net118235), .A1(n205), .B0(net118259), .B1(n317), .Y(
        n7084) );
  AO22X1 U9681 ( .A0(net118239), .A1(n206), .B0(net118261), .B1(n932), .Y(
        n8989) );
  AO22X1 U9682 ( .A0(net118233), .A1(n724), .B0(net118259), .B1(n2346), .Y(
        n7519) );
  AO22X1 U9683 ( .A0(net118233), .A1(n721), .B0(net118259), .B1(n2343), .Y(
        n7510) );
  AO22X1 U9684 ( .A0(n5157), .A1(n840), .B0(n5153), .B1(n2459), .Y(n8359) );
  AO22X1 U9685 ( .A0(net118235), .A1(n207), .B0(net118259), .B1(n318), .Y(
        n7093) );
  AO22X1 U9686 ( .A0(net118235), .A1(n208), .B0(net118259), .B1(n319), .Y(
        n6988) );
  AO22X1 U9687 ( .A0(n5156), .A1(n725), .B0(n5152), .B1(n2347), .Y(n7468) );
  AO22X1 U9688 ( .A0(n5156), .A1(n900), .B0(n5152), .B1(n2529), .Y(n7459) );
  AO22X1 U9689 ( .A0(n5156), .A1(n841), .B0(n5152), .B1(n2460), .Y(n7553) );
  AO22X1 U9690 ( .A0(n5156), .A1(n842), .B0(n5152), .B1(n2461), .Y(n7544) );
  AO22X1 U9691 ( .A0(n5154), .A1(n209), .B0(n5151), .B1(n320), .Y(n7014) );
  AO22X1 U9692 ( .A0(n5157), .A1(n210), .B0(n5151), .B1(n321), .Y(n7005) );
  AO22X1 U9693 ( .A0(n5154), .A1(n211), .B0(n5151), .B1(n322), .Y(n6903) );
  AOI2BB2X4 U9694 ( .B0(n4828), .B1(\I_cache/cache[5][145] ), .A0N(n5808), 
        .A1N(n2922), .Y(n6380) );
  OA22X2 U9695 ( .A0(n5831), .A1(n708), .B0(n5786), .B1(n2328), .Y(n11147) );
  OA22X2 U9696 ( .A0(n5831), .A1(n709), .B0(n5786), .B1(n2329), .Y(n11137) );
  OA22X1 U9697 ( .A0(\i_MIPS/Register/register[22][10] ), .A1(net117675), .B0(
        \i_MIPS/Register/register[30][10] ), .B1(net117697), .Y(n7518) );
  OA22X1 U9698 ( .A0(\i_MIPS/Register/register[22][13] ), .A1(net117675), .B0(
        \i_MIPS/Register/register[30][13] ), .B1(net117695), .Y(n7981) );
  OA22X1 U9699 ( .A0(\i_MIPS/Register/register[22][5] ), .A1(net117681), .B0(
        \i_MIPS/Register/register[30][5] ), .B1(net117703), .Y(n9339) );
  OA22X1 U9700 ( .A0(\i_MIPS/Register/register[22][16] ), .A1(net117685), .B0(
        \i_MIPS/Register/register[30][16] ), .B1(net117697), .Y(n8810) );
  OA22X1 U9701 ( .A0(\i_MIPS/Register/register[22][19] ), .A1(n5082), .B0(
        \i_MIPS/Register/register[30][19] ), .B1(n5078), .Y(n8358) );
  OA22X1 U9702 ( .A0(\i_MIPS/Register/register[6][19] ), .A1(n5082), .B0(
        \i_MIPS/Register/register[14][19] ), .B1(n5078), .Y(n8349) );
  OA22X1 U9703 ( .A0(\i_MIPS/Register/register[22][16] ), .A1(n5083), .B0(
        \i_MIPS/Register/register[30][16] ), .B1(n5079), .Y(n8844) );
  OA22X1 U9704 ( .A0(\i_MIPS/Register/register[6][16] ), .A1(n5083), .B0(
        \i_MIPS/Register/register[14][16] ), .B1(n5079), .Y(n8835) );
  OA22X1 U9705 ( .A0(\i_MIPS/Register/register[22][23] ), .A1(net117673), .B0(
        \i_MIPS/Register/register[30][23] ), .B1(net117691), .Y(n7092) );
  OA22X1 U9706 ( .A0(\i_MIPS/Register/register[22][27] ), .A1(n5081), .B0(
        \i_MIPS/Register/register[30][27] ), .B1(n5077), .Y(n7728) );
  OA22X1 U9707 ( .A0(\i_MIPS/Register/register[6][27] ), .A1(n5081), .B0(
        \i_MIPS/Register/register[14][27] ), .B1(n5077), .Y(n7719) );
  OA22X1 U9708 ( .A0(\i_MIPS/Register/register[22][29] ), .A1(net117673), .B0(
        \i_MIPS/Register/register[30][29] ), .B1(net117691), .Y(n6996) );
  OA22X1 U9709 ( .A0(\i_MIPS/Register/register[21][10] ), .A1(net118401), .B0(
        \i_MIPS/Register/register[29][10] ), .B1(net118425), .Y(n7516) );
  OA22X1 U9710 ( .A0(\i_MIPS/Register/register[21][13] ), .A1(net118403), .B0(
        \i_MIPS/Register/register[29][13] ), .B1(net118429), .Y(n7979) );
  OA22X1 U9711 ( .A0(\i_MIPS/Register/register[21][5] ), .A1(net118407), .B0(
        \i_MIPS/Register/register[29][5] ), .B1(net118431), .Y(n9337) );
  OA22X1 U9712 ( .A0(\i_MIPS/Register/register[21][3] ), .A1(net118407), .B0(
        \i_MIPS/Register/register[29][3] ), .B1(net118431), .Y(n9156) );
  OA22X1 U9713 ( .A0(\i_MIPS/Register/register[21][0] ), .A1(net118405), .B0(
        \i_MIPS/Register/register[29][0] ), .B1(net118429), .Y(n8732) );
  OA22X1 U9714 ( .A0(\i_MIPS/Register/register[21][16] ), .A1(net118405), .B0(
        \i_MIPS/Register/register[29][16] ), .B1(net118429), .Y(n8808) );
  OA22X1 U9715 ( .A0(\i_MIPS/Register/register[21][23] ), .A1(net118399), .B0(
        \i_MIPS/Register/register[29][23] ), .B1(net118423), .Y(n7090) );
  OA22X1 U9716 ( .A0(\i_MIPS/Register/register[21][29] ), .A1(net118399), .B0(
        \i_MIPS/Register/register[29][29] ), .B1(net118423), .Y(n6994) );
  AO22X1 U9717 ( .A0(net118275), .A1(n288), .B0(net118291), .B1(n2462), .Y(
        n9065) );
  AO22X1 U9718 ( .A0(net118275), .A1(n264), .B0(net118291), .B1(n2350), .Y(
        n9241) );
  AO22X1 U9719 ( .A0(net118275), .A1(n267), .B0(net118291), .B1(n2358), .Y(
        n9151) );
  AO22X1 U9720 ( .A0(net118273), .A1(n843), .B0(net118291), .B1(n2463), .Y(
        n8498) );
  AO22X1 U9721 ( .A0(net118271), .A1(n844), .B0(net118289), .B1(n2464), .Y(
        n8317) );
  AO22X1 U9722 ( .A0(net118275), .A1(n265), .B0(net118291), .B1(n2351), .Y(
        n9332) );
  AO22X1 U9723 ( .A0(net118273), .A1(n845), .B0(net118291), .B1(n2465), .Y(
        n8803) );
  AO22X1 U9724 ( .A0(net118273), .A1(n846), .B0(net118291), .B1(n2466), .Y(
        n8727) );
  AO22X1 U9725 ( .A0(net118271), .A1(n847), .B0(net118289), .B1(n2467), .Y(
        n8227) );
  AO22X1 U9726 ( .A0(net118275), .A1(n289), .B0(net118291), .B1(n2468), .Y(
        n8990) );
  AO22X1 U9727 ( .A0(net118271), .A1(n848), .B0(net118289), .B1(n2469), .Y(
        n8147) );
  AO22X1 U9728 ( .A0(net118267), .A1(n290), .B0(net118295), .B1(n933), .Y(
        n7085) );
  AO22X1 U9729 ( .A0(net118269), .A1(n722), .B0(net118295), .B1(n2344), .Y(
        n7511) );
  AO22X1 U9730 ( .A0(net118269), .A1(n901), .B0(net118295), .B1(n2530), .Y(
        n7326) );
  AO22X1 U9731 ( .A0(net118269), .A1(n849), .B0(net118295), .B1(n2470), .Y(
        n7246) );
  AO22X1 U9732 ( .A0(net118269), .A1(n850), .B0(net118295), .B1(n2471), .Y(
        n7385) );
  AO22X1 U9733 ( .A0(net118267), .A1(n291), .B0(net118295), .B1(n934), .Y(
        n6989) );
  AO22X1 U9734 ( .A0(net118271), .A1(n851), .B0(net118289), .B1(n2472), .Y(
        n7974) );
  AO22X1 U9735 ( .A0(net118267), .A1(n292), .B0(net118295), .B1(n935), .Y(
        n7171) );
  AO22X1 U9736 ( .A0(net118269), .A1(n852), .B0(net118295), .B1(n2473), .Y(
        n7655) );
  AO22X1 U9737 ( .A0(net118269), .A1(n902), .B0(net118295), .B1(n2531), .Y(
        n7569) );
  AO22X1 U9738 ( .A0(net118267), .A1(n302), .B0(net118295), .B1(n952), .Y(
        n6878) );
  AO22X1 U9739 ( .A0(net118267), .A1(n220), .B0(net118291), .B1(n329), .Y(
        n6778) );
  MX2XL U9740 ( .A(\D_cache/cache[6][51] ), .B(n4536), .S0(n3574), .Y(
        \D_cache/n1382 ) );
  MX2XL U9741 ( .A(\D_cache/cache[5][51] ), .B(n4536), .S0(n5350), .Y(
        \D_cache/n1383 ) );
  MX2XL U9742 ( .A(\D_cache/cache[4][51] ), .B(n4536), .S0(n5323), .Y(
        \D_cache/n1384 ) );
  MX2XL U9743 ( .A(\D_cache/cache[3][51] ), .B(n4536), .S0(n5276), .Y(
        \D_cache/n1385 ) );
  MX2XL U9744 ( .A(\D_cache/cache[2][51] ), .B(n4536), .S0(n5236), .Y(
        \D_cache/n1386 ) );
  MX2XL U9745 ( .A(\D_cache/cache[1][51] ), .B(n4536), .S0(n5208), .Y(
        \D_cache/n1387 ) );
  MX2XL U9746 ( .A(\D_cache/cache[0][51] ), .B(n4536), .S0(n5168), .Y(
        \D_cache/n1388 ) );
  MX2XL U9747 ( .A(\D_cache/cache[6][19] ), .B(n10965), .S0(n3574), .Y(
        \D_cache/n1638 ) );
  MX2XL U9748 ( .A(\D_cache/cache[5][19] ), .B(n10965), .S0(n5350), .Y(
        \D_cache/n1639 ) );
  MX2XL U9749 ( .A(\D_cache/cache[4][19] ), .B(n10965), .S0(n5323), .Y(
        \D_cache/n1640 ) );
  MX2XL U9750 ( .A(\D_cache/cache[3][19] ), .B(n10965), .S0(n5276), .Y(
        \D_cache/n1641 ) );
  MX2XL U9751 ( .A(\D_cache/cache[2][19] ), .B(n10965), .S0(n5236), .Y(
        \D_cache/n1642 ) );
  MX2XL U9752 ( .A(\D_cache/cache[1][19] ), .B(n10965), .S0(n5208), .Y(
        \D_cache/n1643 ) );
  MX2XL U9753 ( .A(\D_cache/cache[0][19] ), .B(n10965), .S0(n5168), .Y(
        \D_cache/n1644 ) );
  MX2XL U9754 ( .A(\D_cache/cache[6][127] ), .B(n10707), .S0(n5369), .Y(
        \D_cache/n774 ) );
  MX2XL U9755 ( .A(\D_cache/cache[5][127] ), .B(n10707), .S0(n3575), .Y(
        \D_cache/n775 ) );
  MX2XL U9756 ( .A(\D_cache/cache[4][127] ), .B(n10707), .S0(n5318), .Y(
        \D_cache/n776 ) );
  MX2XL U9757 ( .A(\D_cache/cache[3][127] ), .B(n10707), .S0(n5273), .Y(
        \D_cache/n777 ) );
  MX2XL U9758 ( .A(\D_cache/cache[2][127] ), .B(n10707), .S0(n5231), .Y(
        \D_cache/n778 ) );
  MX2XL U9759 ( .A(\D_cache/cache[1][127] ), .B(n10707), .S0(n5203), .Y(
        \D_cache/n779 ) );
  MX2XL U9760 ( .A(\D_cache/cache[0][127] ), .B(n10707), .S0(n5163), .Y(
        \D_cache/n780 ) );
  MX2XL U9761 ( .A(\D_cache/cache[6][126] ), .B(n10600), .S0(n5369), .Y(
        \D_cache/n782 ) );
  MX2XL U9762 ( .A(\D_cache/cache[5][126] ), .B(n10600), .S0(n3575), .Y(
        \D_cache/n783 ) );
  MX2XL U9763 ( .A(\D_cache/cache[4][126] ), .B(n10600), .S0(n5318), .Y(
        \D_cache/n784 ) );
  MX2XL U9764 ( .A(\D_cache/cache[3][126] ), .B(n10600), .S0(n5273), .Y(
        \D_cache/n785 ) );
  MX2XL U9765 ( .A(\D_cache/cache[2][126] ), .B(n10600), .S0(n5231), .Y(
        \D_cache/n786 ) );
  MX2XL U9766 ( .A(\D_cache/cache[1][126] ), .B(n10600), .S0(n5205), .Y(
        \D_cache/n787 ) );
  MX2XL U9767 ( .A(\D_cache/cache[0][126] ), .B(n10600), .S0(n5164), .Y(
        \D_cache/n788 ) );
  MX2XL U9768 ( .A(\D_cache/cache[6][125] ), .B(n10563), .S0(n5370), .Y(
        \D_cache/n790 ) );
  MX2XL U9769 ( .A(\D_cache/cache[5][125] ), .B(n10563), .S0(n5346), .Y(
        \D_cache/n791 ) );
  MX2XL U9770 ( .A(\D_cache/cache[4][125] ), .B(n10563), .S0(n5319), .Y(
        \D_cache/n792 ) );
  MX2XL U9771 ( .A(\D_cache/cache[3][125] ), .B(n10563), .S0(n5274), .Y(
        \D_cache/n793 ) );
  MX2XL U9772 ( .A(\D_cache/cache[2][125] ), .B(n10563), .S0(n5232), .Y(
        \D_cache/n794 ) );
  MX2XL U9773 ( .A(\D_cache/cache[1][125] ), .B(n10563), .S0(n5204), .Y(
        \D_cache/n795 ) );
  MX2XL U9774 ( .A(\D_cache/cache[0][125] ), .B(n10563), .S0(n5164), .Y(
        \D_cache/n796 ) );
  MX2XL U9775 ( .A(\D_cache/cache[6][124] ), .B(n10550), .S0(n5370), .Y(
        \D_cache/n798 ) );
  MX2XL U9776 ( .A(\D_cache/cache[5][124] ), .B(n10550), .S0(n5346), .Y(
        \D_cache/n799 ) );
  MX2XL U9777 ( .A(\D_cache/cache[4][124] ), .B(n10550), .S0(n5319), .Y(
        \D_cache/n800 ) );
  MX2XL U9778 ( .A(\D_cache/cache[3][124] ), .B(n10550), .S0(n5269), .Y(
        \D_cache/n801 ) );
  MX2XL U9779 ( .A(\D_cache/cache[2][124] ), .B(n10550), .S0(n5232), .Y(
        \D_cache/n802 ) );
  MX2XL U9780 ( .A(\D_cache/cache[1][124] ), .B(n10550), .S0(n5204), .Y(
        \D_cache/n803 ) );
  MX2XL U9781 ( .A(\D_cache/cache[0][124] ), .B(n10550), .S0(n5164), .Y(
        \D_cache/n804 ) );
  MX2XL U9782 ( .A(\D_cache/cache[6][123] ), .B(n4522), .S0(n5366), .Y(
        \D_cache/n806 ) );
  MX2XL U9783 ( .A(\D_cache/cache[5][123] ), .B(n4522), .S0(n5342), .Y(
        \D_cache/n807 ) );
  MX2XL U9784 ( .A(\D_cache/cache[4][123] ), .B(n4522), .S0(n5315), .Y(
        \D_cache/n808 ) );
  MX2XL U9785 ( .A(\D_cache/cache[3][123] ), .B(n4522), .S0(n5270), .Y(
        \D_cache/n809 ) );
  MX2XL U9786 ( .A(\D_cache/cache[2][123] ), .B(n4522), .S0(n5230), .Y(
        \D_cache/n810 ) );
  MX2XL U9787 ( .A(\D_cache/cache[1][123] ), .B(n4522), .S0(n5200), .Y(
        \D_cache/n811 ) );
  MX2XL U9788 ( .A(\D_cache/cache[0][123] ), .B(n4522), .S0(n5159), .Y(
        \D_cache/n812 ) );
  MX2XL U9789 ( .A(\D_cache/cache[6][122] ), .B(n4523), .S0(n5367), .Y(
        \D_cache/n814 ) );
  MX2XL U9790 ( .A(\D_cache/cache[5][122] ), .B(n4523), .S0(n5343), .Y(
        \D_cache/n815 ) );
  MX2XL U9791 ( .A(\D_cache/cache[4][122] ), .B(n4523), .S0(n5316), .Y(
        \D_cache/n816 ) );
  MX2XL U9792 ( .A(\D_cache/cache[3][122] ), .B(n4523), .S0(n5271), .Y(
        \D_cache/n817 ) );
  MX2XL U9793 ( .A(\D_cache/cache[2][122] ), .B(n4523), .S0(n5229), .Y(
        \D_cache/n818 ) );
  MX2XL U9794 ( .A(\D_cache/cache[1][122] ), .B(n4523), .S0(n5201), .Y(
        \D_cache/n819 ) );
  MX2XL U9795 ( .A(\D_cache/cache[0][122] ), .B(n4523), .S0(n5161), .Y(
        \D_cache/n820 ) );
  MX2XL U9796 ( .A(\D_cache/cache[6][121] ), .B(n10439), .S0(n5364), .Y(
        \D_cache/n822 ) );
  MX2XL U9797 ( .A(\D_cache/cache[5][121] ), .B(n10439), .S0(n5340), .Y(
        \D_cache/n823 ) );
  MX2XL U9798 ( .A(\D_cache/cache[4][121] ), .B(n10439), .S0(n5313), .Y(
        \D_cache/n824 ) );
  MX2XL U9799 ( .A(\D_cache/cache[3][121] ), .B(n10439), .S0(n5268), .Y(
        \D_cache/n825 ) );
  MX2XL U9800 ( .A(\D_cache/cache[2][121] ), .B(n10439), .S0(n5228), .Y(
        \D_cache/n826 ) );
  MX2XL U9801 ( .A(\D_cache/cache[1][121] ), .B(n10439), .S0(n5198), .Y(
        \D_cache/n827 ) );
  MX2XL U9802 ( .A(\D_cache/cache[0][121] ), .B(n10439), .S0(n5163), .Y(
        \D_cache/n828 ) );
  MX2XL U9803 ( .A(\D_cache/cache[6][120] ), .B(n4517), .S0(n5364), .Y(
        \D_cache/n830 ) );
  MX2XL U9804 ( .A(\D_cache/cache[5][120] ), .B(n4517), .S0(n5340), .Y(
        \D_cache/n831 ) );
  MX2XL U9805 ( .A(\D_cache/cache[4][120] ), .B(n4517), .S0(n5313), .Y(
        \D_cache/n832 ) );
  MX2XL U9806 ( .A(\D_cache/cache[3][120] ), .B(n4517), .S0(n5268), .Y(
        \D_cache/n833 ) );
  MX2XL U9807 ( .A(\D_cache/cache[2][120] ), .B(n4517), .S0(n5228), .Y(
        \D_cache/n834 ) );
  MX2XL U9808 ( .A(\D_cache/cache[1][120] ), .B(n4517), .S0(n5198), .Y(
        \D_cache/n835 ) );
  MX2XL U9809 ( .A(\D_cache/cache[0][120] ), .B(n4517), .S0(n5159), .Y(
        \D_cache/n836 ) );
  MX2XL U9810 ( .A(\D_cache/cache[6][119] ), .B(n10694), .S0(n5369), .Y(
        \D_cache/n838 ) );
  MX2XL U9811 ( .A(\D_cache/cache[5][119] ), .B(n10694), .S0(n3575), .Y(
        \D_cache/n839 ) );
  MX2XL U9812 ( .A(\D_cache/cache[4][119] ), .B(n10694), .S0(n5318), .Y(
        \D_cache/n840 ) );
  MX2XL U9813 ( .A(\D_cache/cache[3][119] ), .B(n10694), .S0(n5273), .Y(
        \D_cache/n841 ) );
  MX2XL U9814 ( .A(\D_cache/cache[2][119] ), .B(n10694), .S0(n5231), .Y(
        \D_cache/n842 ) );
  MX2XL U9815 ( .A(\D_cache/cache[1][119] ), .B(n10694), .S0(n5203), .Y(
        \D_cache/n843 ) );
  MX2XL U9816 ( .A(\D_cache/cache[0][119] ), .B(n10694), .S0(n5163), .Y(
        \D_cache/n844 ) );
  MX2XL U9817 ( .A(\D_cache/cache[6][118] ), .B(n10315), .S0(n5367), .Y(
        \D_cache/n846 ) );
  MX2XL U9818 ( .A(\D_cache/cache[5][118] ), .B(n10315), .S0(n5343), .Y(
        \D_cache/n847 ) );
  MX2XL U9819 ( .A(\D_cache/cache[4][118] ), .B(n10315), .S0(n5316), .Y(
        \D_cache/n848 ) );
  MX2XL U9820 ( .A(\D_cache/cache[3][118] ), .B(n10315), .S0(n5271), .Y(
        \D_cache/n849 ) );
  MX2XL U9821 ( .A(\D_cache/cache[2][118] ), .B(n10315), .S0(n5229), .Y(
        \D_cache/n850 ) );
  MX2XL U9822 ( .A(\D_cache/cache[1][118] ), .B(n10315), .S0(n5201), .Y(
        \D_cache/n851 ) );
  MX2XL U9823 ( .A(\D_cache/cache[0][118] ), .B(n10315), .S0(n5161), .Y(
        \D_cache/n852 ) );
  MX2XL U9824 ( .A(\D_cache/cache[6][117] ), .B(n10522), .S0(n5370), .Y(
        \D_cache/n854 ) );
  MX2XL U9825 ( .A(\D_cache/cache[5][117] ), .B(n10522), .S0(n5346), .Y(
        \D_cache/n855 ) );
  MX2XL U9826 ( .A(\D_cache/cache[4][117] ), .B(n10522), .S0(n5319), .Y(
        \D_cache/n856 ) );
  MX2XL U9827 ( .A(\D_cache/cache[3][117] ), .B(n10522), .S0(n5275), .Y(
        \D_cache/n857 ) );
  MX2XL U9828 ( .A(\D_cache/cache[2][117] ), .B(n10522), .S0(n5232), .Y(
        \D_cache/n858 ) );
  MX2XL U9829 ( .A(\D_cache/cache[1][117] ), .B(n10522), .S0(n5204), .Y(
        \D_cache/n859 ) );
  MX2XL U9830 ( .A(\D_cache/cache[0][117] ), .B(n10522), .S0(n3564), .Y(
        \D_cache/n860 ) );
  MX2XL U9831 ( .A(\D_cache/cache[6][116] ), .B(n4518), .S0(n5364), .Y(
        \D_cache/n862 ) );
  MX2XL U9832 ( .A(\D_cache/cache[5][116] ), .B(n4518), .S0(n5340), .Y(
        \D_cache/n863 ) );
  MX2XL U9833 ( .A(\D_cache/cache[4][116] ), .B(n4518), .S0(n5313), .Y(
        \D_cache/n864 ) );
  MX2XL U9834 ( .A(\D_cache/cache[3][116] ), .B(n4518), .S0(n5268), .Y(
        \D_cache/n865 ) );
  MX2XL U9835 ( .A(\D_cache/cache[2][116] ), .B(n4518), .S0(n5228), .Y(
        \D_cache/n866 ) );
  MX2XL U9836 ( .A(\D_cache/cache[1][116] ), .B(n4518), .S0(n5198), .Y(
        \D_cache/n867 ) );
  MX2XL U9837 ( .A(\D_cache/cache[0][116] ), .B(n4518), .S0(n5159), .Y(
        \D_cache/n868 ) );
  MX2XL U9838 ( .A(\D_cache/cache[6][114] ), .B(n10642), .S0(n5371), .Y(
        \D_cache/n878 ) );
  MX2XL U9839 ( .A(\D_cache/cache[5][114] ), .B(n10642), .S0(n5347), .Y(
        \D_cache/n879 ) );
  MX2XL U9840 ( .A(\D_cache/cache[4][114] ), .B(n10642), .S0(n5320), .Y(
        \D_cache/n880 ) );
  MX2XL U9841 ( .A(\D_cache/cache[3][114] ), .B(n10642), .S0(n5274), .Y(
        \D_cache/n881 ) );
  MX2XL U9842 ( .A(\D_cache/cache[2][114] ), .B(n10642), .S0(n5233), .Y(
        \D_cache/n882 ) );
  MX2XL U9843 ( .A(\D_cache/cache[1][114] ), .B(n10642), .S0(n5204), .Y(
        \D_cache/n883 ) );
  MX2XL U9844 ( .A(\D_cache/cache[0][114] ), .B(n10642), .S0(n5162), .Y(
        \D_cache/n884 ) );
  MX2XL U9845 ( .A(\D_cache/cache[6][113] ), .B(n10627), .S0(n5371), .Y(
        \D_cache/n886 ) );
  MX2XL U9846 ( .A(\D_cache/cache[5][113] ), .B(n10627), .S0(n5347), .Y(
        \D_cache/n887 ) );
  MX2XL U9847 ( .A(\D_cache/cache[4][113] ), .B(n10627), .S0(n5320), .Y(
        \D_cache/n888 ) );
  MX2XL U9848 ( .A(\D_cache/cache[3][113] ), .B(n10627), .S0(n5274), .Y(
        \D_cache/n889 ) );
  MX2XL U9849 ( .A(\D_cache/cache[2][113] ), .B(n10627), .S0(n5233), .Y(
        \D_cache/n890 ) );
  MX2XL U9850 ( .A(\D_cache/cache[1][113] ), .B(n10627), .S0(n5205), .Y(
        \D_cache/n891 ) );
  MX2XL U9851 ( .A(\D_cache/cache[0][113] ), .B(n10627), .S0(n5164), .Y(
        \D_cache/n892 ) );
  MX2XL U9852 ( .A(\D_cache/cache[6][112] ), .B(n4519), .S0(n5365), .Y(
        \D_cache/n894 ) );
  MX2XL U9853 ( .A(\D_cache/cache[5][112] ), .B(n4519), .S0(n5341), .Y(
        \D_cache/n895 ) );
  MX2XL U9854 ( .A(\D_cache/cache[4][112] ), .B(n4519), .S0(n5314), .Y(
        \D_cache/n896 ) );
  MX2XL U9855 ( .A(\D_cache/cache[3][112] ), .B(n4519), .S0(n5269), .Y(
        \D_cache/n897 ) );
  MX2XL U9856 ( .A(\D_cache/cache[2][112] ), .B(n4519), .S0(n5231), .Y(
        \D_cache/n898 ) );
  MX2XL U9857 ( .A(\D_cache/cache[1][112] ), .B(n4519), .S0(n5199), .Y(
        \D_cache/n899 ) );
  MX2XL U9858 ( .A(\D_cache/cache[0][112] ), .B(n4519), .S0(n5160), .Y(
        \D_cache/n900 ) );
  MX2XL U9859 ( .A(\D_cache/cache[6][111] ), .B(n4520), .S0(n5365), .Y(
        \D_cache/n902 ) );
  MX2XL U9860 ( .A(\D_cache/cache[5][111] ), .B(n4520), .S0(n5341), .Y(
        \D_cache/n903 ) );
  MX2XL U9861 ( .A(\D_cache/cache[4][111] ), .B(n4520), .S0(n5314), .Y(
        \D_cache/n904 ) );
  MX2XL U9862 ( .A(\D_cache/cache[3][111] ), .B(n4520), .S0(n5269), .Y(
        \D_cache/n905 ) );
  MX2XL U9863 ( .A(\D_cache/cache[2][111] ), .B(n4520), .S0(n5235), .Y(
        \D_cache/n906 ) );
  MX2XL U9864 ( .A(\D_cache/cache[1][111] ), .B(n4520), .S0(n5199), .Y(
        \D_cache/n907 ) );
  MX2XL U9865 ( .A(\D_cache/cache[0][111] ), .B(n4520), .S0(n5160), .Y(
        \D_cache/n908 ) );
  MX2XL U9866 ( .A(\D_cache/cache[6][110] ), .B(n4527), .S0(n5366), .Y(
        \D_cache/n910 ) );
  MX2XL U9867 ( .A(\D_cache/cache[5][110] ), .B(n4527), .S0(n5342), .Y(
        \D_cache/n911 ) );
  MX2XL U9868 ( .A(\D_cache/cache[4][110] ), .B(n4527), .S0(n5315), .Y(
        \D_cache/n912 ) );
  MX2XL U9869 ( .A(\D_cache/cache[3][110] ), .B(n4527), .S0(n5270), .Y(
        \D_cache/n913 ) );
  MX2XL U9870 ( .A(\D_cache/cache[2][110] ), .B(n4527), .S0(n5228), .Y(
        \D_cache/n914 ) );
  MX2XL U9871 ( .A(\D_cache/cache[1][110] ), .B(n4527), .S0(n5200), .Y(
        \D_cache/n915 ) );
  MX2XL U9872 ( .A(\D_cache/cache[0][110] ), .B(n4527), .S0(n5167), .Y(
        \D_cache/n916 ) );
  MX2XL U9873 ( .A(\D_cache/cache[6][108] ), .B(n4521), .S0(n5365), .Y(
        \D_cache/n926 ) );
  MX2XL U9874 ( .A(\D_cache/cache[5][108] ), .B(n4521), .S0(n5341), .Y(
        \D_cache/n927 ) );
  MX2XL U9875 ( .A(\D_cache/cache[4][108] ), .B(n4521), .S0(n5314), .Y(
        \D_cache/n928 ) );
  MX2XL U9876 ( .A(\D_cache/cache[3][108] ), .B(n4521), .S0(n5269), .Y(
        \D_cache/n929 ) );
  MX2XL U9877 ( .A(\D_cache/cache[2][108] ), .B(n4521), .S0(n5232), .Y(
        \D_cache/n930 ) );
  MX2XL U9878 ( .A(\D_cache/cache[1][108] ), .B(n4521), .S0(n5199), .Y(
        \D_cache/n931 ) );
  MX2XL U9879 ( .A(\D_cache/cache[0][108] ), .B(n4521), .S0(n5160), .Y(
        \D_cache/n932 ) );
  MX2XL U9880 ( .A(\D_cache/cache[6][105] ), .B(n10614), .S0(n5371), .Y(
        \D_cache/n950 ) );
  MX2XL U9881 ( .A(\D_cache/cache[5][105] ), .B(n10614), .S0(n5347), .Y(
        \D_cache/n951 ) );
  MX2XL U9882 ( .A(\D_cache/cache[4][105] ), .B(n10614), .S0(n5320), .Y(
        \D_cache/n952 ) );
  MX2XL U9883 ( .A(\D_cache/cache[3][105] ), .B(n10614), .S0(n5274), .Y(
        \D_cache/n953 ) );
  MX2XL U9884 ( .A(\D_cache/cache[2][105] ), .B(n10614), .S0(n5233), .Y(
        \D_cache/n954 ) );
  MX2XL U9885 ( .A(\D_cache/cache[1][105] ), .B(n10614), .S0(n5205), .Y(
        \D_cache/n955 ) );
  MX2XL U9886 ( .A(\D_cache/cache[0][105] ), .B(n10614), .S0(n5164), .Y(
        \D_cache/n956 ) );
  MX2XL U9887 ( .A(\D_cache/cache[6][104] ), .B(n10655), .S0(n5368), .Y(
        \D_cache/n958 ) );
  MX2XL U9888 ( .A(\D_cache/cache[5][104] ), .B(n10655), .S0(n5344), .Y(
        \D_cache/n959 ) );
  MX2XL U9889 ( .A(\D_cache/cache[4][104] ), .B(n10655), .S0(n5317), .Y(
        \D_cache/n960 ) );
  MX2XL U9890 ( .A(\D_cache/cache[3][104] ), .B(n10655), .S0(n5272), .Y(
        \D_cache/n961 ) );
  MX2XL U9891 ( .A(\D_cache/cache[2][104] ), .B(n10655), .S0(n5230), .Y(
        \D_cache/n962 ) );
  MX2XL U9892 ( .A(\D_cache/cache[1][104] ), .B(n10655), .S0(n5202), .Y(
        \D_cache/n963 ) );
  MX2XL U9893 ( .A(\D_cache/cache[0][104] ), .B(n10655), .S0(n5162), .Y(
        \D_cache/n964 ) );
  MX2XL U9894 ( .A(\D_cache/cache[6][103] ), .B(n10682), .S0(n5367), .Y(
        \D_cache/n966 ) );
  MX2XL U9895 ( .A(\D_cache/cache[5][103] ), .B(n10682), .S0(n5343), .Y(
        \D_cache/n967 ) );
  MX2XL U9896 ( .A(\D_cache/cache[4][103] ), .B(n10682), .S0(n5316), .Y(
        \D_cache/n968 ) );
  MX2XL U9897 ( .A(\D_cache/cache[3][103] ), .B(n10682), .S0(n5271), .Y(
        \D_cache/n969 ) );
  MX2XL U9898 ( .A(\D_cache/cache[2][103] ), .B(n10682), .S0(n5229), .Y(
        \D_cache/n970 ) );
  MX2XL U9899 ( .A(\D_cache/cache[1][103] ), .B(n10682), .S0(n5201), .Y(
        \D_cache/n971 ) );
  MX2XL U9900 ( .A(\D_cache/cache[0][103] ), .B(n10682), .S0(n5163), .Y(
        \D_cache/n972 ) );
  MX2XL U9901 ( .A(\D_cache/cache[6][102] ), .B(n4528), .S0(n5366), .Y(
        \D_cache/n974 ) );
  MX2XL U9902 ( .A(\D_cache/cache[5][102] ), .B(n4528), .S0(n5342), .Y(
        \D_cache/n975 ) );
  MX2XL U9903 ( .A(\D_cache/cache[4][102] ), .B(n4528), .S0(n5315), .Y(
        \D_cache/n976 ) );
  MX2XL U9904 ( .A(\D_cache/cache[3][102] ), .B(n4528), .S0(n5270), .Y(
        \D_cache/n977 ) );
  MX2XL U9905 ( .A(\D_cache/cache[2][102] ), .B(n4528), .S0(n5231), .Y(
        \D_cache/n978 ) );
  MX2XL U9906 ( .A(\D_cache/cache[1][102] ), .B(n4528), .S0(n5200), .Y(
        \D_cache/n979 ) );
  MX2XL U9907 ( .A(\D_cache/cache[0][102] ), .B(n4528), .S0(n5167), .Y(
        \D_cache/n980 ) );
  MX2XL U9908 ( .A(\D_cache/cache[6][98] ), .B(n10194), .S0(n5366), .Y(
        \D_cache/n1006 ) );
  MX2XL U9909 ( .A(\D_cache/cache[5][98] ), .B(n10194), .S0(n5342), .Y(
        \D_cache/n1007 ) );
  MX2XL U9910 ( .A(\D_cache/cache[4][98] ), .B(n10194), .S0(n5315), .Y(
        \D_cache/n1008 ) );
  MX2XL U9911 ( .A(\D_cache/cache[3][98] ), .B(n10194), .S0(n5270), .Y(
        \D_cache/n1009 ) );
  MX2XL U9912 ( .A(\D_cache/cache[2][98] ), .B(n10194), .S0(n5233), .Y(
        \D_cache/n1010 ) );
  MX2XL U9913 ( .A(\D_cache/cache[1][98] ), .B(n10194), .S0(n5201), .Y(
        \D_cache/n1011 ) );
  MX2XL U9914 ( .A(\D_cache/cache[0][98] ), .B(n10194), .S0(n5161), .Y(
        \D_cache/n1012 ) );
  MX2XL U9915 ( .A(\D_cache/cache[6][63] ), .B(n4562), .S0(n5369), .Y(
        \D_cache/n1286 ) );
  MX2XL U9916 ( .A(\D_cache/cache[5][63] ), .B(n4562), .S0(n3575), .Y(
        \D_cache/n1287 ) );
  MX2XL U9917 ( .A(\D_cache/cache[4][63] ), .B(n4562), .S0(n5318), .Y(
        \D_cache/n1288 ) );
  MX2XL U9918 ( .A(\D_cache/cache[3][63] ), .B(n4562), .S0(n5273), .Y(
        \D_cache/n1289 ) );
  MX2XL U9919 ( .A(\D_cache/cache[2][63] ), .B(n4562), .S0(n5231), .Y(
        \D_cache/n1290 ) );
  MX2XL U9920 ( .A(\D_cache/cache[1][63] ), .B(n4562), .S0(n5203), .Y(
        \D_cache/n1291 ) );
  MX2XL U9921 ( .A(\D_cache/cache[0][63] ), .B(n4562), .S0(n5163), .Y(
        \D_cache/n1292 ) );
  MX2XL U9922 ( .A(\D_cache/cache[6][62] ), .B(n4563), .S0(n5370), .Y(
        \D_cache/n1294 ) );
  MX2XL U9923 ( .A(\D_cache/cache[5][62] ), .B(n4563), .S0(n5346), .Y(
        \D_cache/n1295 ) );
  MX2XL U9924 ( .A(\D_cache/cache[4][62] ), .B(n4563), .S0(n5319), .Y(
        \D_cache/n1296 ) );
  MX2XL U9925 ( .A(\D_cache/cache[3][62] ), .B(n4563), .S0(n5274), .Y(
        \D_cache/n1297 ) );
  MX2XL U9926 ( .A(\D_cache/cache[2][62] ), .B(n4563), .S0(n5232), .Y(
        \D_cache/n1298 ) );
  MX2XL U9927 ( .A(\D_cache/cache[1][62] ), .B(n4563), .S0(n5203), .Y(
        \D_cache/n1299 ) );
  MX2XL U9928 ( .A(\D_cache/cache[0][62] ), .B(n4563), .S0(n5164), .Y(
        \D_cache/n1300 ) );
  MX2XL U9929 ( .A(\D_cache/cache[6][61] ), .B(n4564), .S0(n5370), .Y(
        \D_cache/n1302 ) );
  MX2XL U9930 ( .A(\D_cache/cache[5][61] ), .B(n4564), .S0(n5346), .Y(
        \D_cache/n1303 ) );
  MX2XL U9931 ( .A(\D_cache/cache[4][61] ), .B(n4564), .S0(n5319), .Y(
        \D_cache/n1304 ) );
  MX2XL U9932 ( .A(\D_cache/cache[3][61] ), .B(n4564), .S0(n5276), .Y(
        \D_cache/n1305 ) );
  MX2XL U9933 ( .A(\D_cache/cache[2][61] ), .B(n4564), .S0(n5232), .Y(
        \D_cache/n1306 ) );
  MX2XL U9934 ( .A(\D_cache/cache[1][61] ), .B(n4564), .S0(n5204), .Y(
        \D_cache/n1307 ) );
  MX2XL U9935 ( .A(\D_cache/cache[0][61] ), .B(n4564), .S0(n3565), .Y(
        \D_cache/n1308 ) );
  MX2XL U9936 ( .A(\D_cache/cache[6][60] ), .B(n4565), .S0(n5370), .Y(
        \D_cache/n1310 ) );
  MX2XL U9937 ( .A(\D_cache/cache[5][60] ), .B(n4565), .S0(n5346), .Y(
        \D_cache/n1311 ) );
  MX2XL U9938 ( .A(\D_cache/cache[4][60] ), .B(n4565), .S0(n5319), .Y(
        \D_cache/n1312 ) );
  MX2XL U9939 ( .A(\D_cache/cache[3][60] ), .B(n4565), .S0(n5273), .Y(
        \D_cache/n1313 ) );
  MX2XL U9940 ( .A(\D_cache/cache[2][60] ), .B(n4565), .S0(n5232), .Y(
        \D_cache/n1314 ) );
  MX2XL U9941 ( .A(\D_cache/cache[1][60] ), .B(n4565), .S0(n5204), .Y(
        \D_cache/n1315 ) );
  MX2XL U9942 ( .A(\D_cache/cache[0][60] ), .B(n4565), .S0(n3565), .Y(
        \D_cache/n1316 ) );
  MX2XL U9943 ( .A(\D_cache/cache[6][59] ), .B(n4553), .S0(n5367), .Y(
        \D_cache/n1318 ) );
  MX2XL U9944 ( .A(\D_cache/cache[5][59] ), .B(n4553), .S0(n5343), .Y(
        \D_cache/n1319 ) );
  MX2XL U9945 ( .A(\D_cache/cache[4][59] ), .B(n4553), .S0(n5316), .Y(
        \D_cache/n1320 ) );
  MX2XL U9946 ( .A(\D_cache/cache[3][59] ), .B(n4553), .S0(n5271), .Y(
        \D_cache/n1321 ) );
  MX2XL U9947 ( .A(\D_cache/cache[2][59] ), .B(n4553), .S0(n5229), .Y(
        \D_cache/n1322 ) );
  MX2XL U9948 ( .A(\D_cache/cache[1][59] ), .B(n4553), .S0(n5200), .Y(
        \D_cache/n1323 ) );
  MX2XL U9949 ( .A(\D_cache/cache[0][59] ), .B(n4553), .S0(n5167), .Y(
        \D_cache/n1324 ) );
  MX2XL U9950 ( .A(\D_cache/cache[6][58] ), .B(n10203), .S0(n5367), .Y(
        \D_cache/n1326 ) );
  MX2XL U9951 ( .A(\D_cache/cache[5][58] ), .B(n10203), .S0(n5343), .Y(
        \D_cache/n1327 ) );
  MX2XL U9952 ( .A(\D_cache/cache[4][58] ), .B(n10203), .S0(n5316), .Y(
        \D_cache/n1328 ) );
  MX2XL U9953 ( .A(\D_cache/cache[3][58] ), .B(n10203), .S0(n5271), .Y(
        \D_cache/n1329 ) );
  MX2XL U9954 ( .A(\D_cache/cache[2][58] ), .B(n10203), .S0(n5229), .Y(
        \D_cache/n1330 ) );
  MX2XL U9955 ( .A(\D_cache/cache[1][58] ), .B(n10203), .S0(n5201), .Y(
        \D_cache/n1331 ) );
  MX2XL U9956 ( .A(\D_cache/cache[0][58] ), .B(n10203), .S0(n5161), .Y(
        \D_cache/n1332 ) );
  MX2XL U9957 ( .A(\D_cache/cache[6][57] ), .B(n4547), .S0(n5364), .Y(
        \D_cache/n1334 ) );
  MX2XL U9958 ( .A(\D_cache/cache[5][57] ), .B(n4547), .S0(n5340), .Y(
        \D_cache/n1335 ) );
  MX2XL U9959 ( .A(\D_cache/cache[4][57] ), .B(n4547), .S0(n5313), .Y(
        \D_cache/n1336 ) );
  MX2XL U9960 ( .A(\D_cache/cache[3][57] ), .B(n4547), .S0(n5268), .Y(
        \D_cache/n1337 ) );
  MX2XL U9961 ( .A(\D_cache/cache[2][57] ), .B(n4547), .S0(n5228), .Y(
        \D_cache/n1338 ) );
  MX2XL U9962 ( .A(\D_cache/cache[1][57] ), .B(n4547), .S0(n5198), .Y(
        \D_cache/n1339 ) );
  MX2XL U9963 ( .A(\D_cache/cache[0][57] ), .B(n4547), .S0(n5159), .Y(
        \D_cache/n1340 ) );
  MX2XL U9964 ( .A(\D_cache/cache[6][56] ), .B(n4548), .S0(n5364), .Y(
        \D_cache/n1342 ) );
  MX2XL U9965 ( .A(\D_cache/cache[5][56] ), .B(n4548), .S0(n5340), .Y(
        \D_cache/n1343 ) );
  MX2XL U9966 ( .A(\D_cache/cache[4][56] ), .B(n4548), .S0(n5313), .Y(
        \D_cache/n1344 ) );
  MX2XL U9967 ( .A(\D_cache/cache[3][56] ), .B(n4548), .S0(n5268), .Y(
        \D_cache/n1345 ) );
  MX2XL U9968 ( .A(\D_cache/cache[2][56] ), .B(n4548), .S0(n5228), .Y(
        \D_cache/n1346 ) );
  MX2XL U9969 ( .A(\D_cache/cache[1][56] ), .B(n4548), .S0(n5198), .Y(
        \D_cache/n1347 ) );
  MX2XL U9970 ( .A(\D_cache/cache[0][56] ), .B(n4548), .S0(n5159), .Y(
        \D_cache/n1348 ) );
  MX2XL U9971 ( .A(\D_cache/cache[6][55] ), .B(n10691), .S0(n5369), .Y(
        \D_cache/n1350 ) );
  MX2XL U9972 ( .A(\D_cache/cache[5][55] ), .B(n10691), .S0(n3575), .Y(
        \D_cache/n1351 ) );
  MX2XL U9973 ( .A(\D_cache/cache[4][55] ), .B(n10691), .S0(n5318), .Y(
        \D_cache/n1352 ) );
  MX2XL U9974 ( .A(\D_cache/cache[3][55] ), .B(n10691), .S0(n5273), .Y(
        \D_cache/n1353 ) );
  MX2XL U9975 ( .A(\D_cache/cache[2][55] ), .B(n10691), .S0(n5231), .Y(
        \D_cache/n1354 ) );
  MX2XL U9976 ( .A(\D_cache/cache[1][55] ), .B(n10691), .S0(n5203), .Y(
        \D_cache/n1355 ) );
  MX2XL U9977 ( .A(\D_cache/cache[0][55] ), .B(n10691), .S0(n5163), .Y(
        \D_cache/n1356 ) );
  MX2XL U9978 ( .A(\D_cache/cache[6][54] ), .B(n4554), .S0(n5367), .Y(
        \D_cache/n1358 ) );
  MX2XL U9979 ( .A(\D_cache/cache[5][54] ), .B(n4554), .S0(n5343), .Y(
        \D_cache/n1359 ) );
  MX2XL U9980 ( .A(\D_cache/cache[4][54] ), .B(n4554), .S0(n5316), .Y(
        \D_cache/n1360 ) );
  MX2XL U9981 ( .A(\D_cache/cache[3][54] ), .B(n4554), .S0(n5271), .Y(
        \D_cache/n1361 ) );
  MX2XL U9982 ( .A(\D_cache/cache[2][54] ), .B(n4554), .S0(n5229), .Y(
        \D_cache/n1362 ) );
  MX2XL U9983 ( .A(\D_cache/cache[1][54] ), .B(n4554), .S0(n5201), .Y(
        \D_cache/n1363 ) );
  MX2XL U9984 ( .A(\D_cache/cache[0][54] ), .B(n4554), .S0(n5161), .Y(
        \D_cache/n1364 ) );
  MX2XL U9985 ( .A(\D_cache/cache[6][53] ), .B(n4566), .S0(n5365), .Y(
        \D_cache/n1366 ) );
  MX2XL U9986 ( .A(\D_cache/cache[5][53] ), .B(n4566), .S0(n5341), .Y(
        \D_cache/n1367 ) );
  MX2XL U9987 ( .A(\D_cache/cache[4][53] ), .B(n4566), .S0(n5314), .Y(
        \D_cache/n1368 ) );
  MX2XL U9988 ( .A(\D_cache/cache[3][53] ), .B(n4566), .S0(n5269), .Y(
        \D_cache/n1369 ) );
  MX2XL U9989 ( .A(\D_cache/cache[2][53] ), .B(n4566), .S0(n5230), .Y(
        \D_cache/n1370 ) );
  MX2XL U9990 ( .A(\D_cache/cache[1][53] ), .B(n4566), .S0(n5204), .Y(
        \D_cache/n1371 ) );
  MX2XL U9991 ( .A(\D_cache/cache[0][53] ), .B(n4566), .S0(n3564), .Y(
        \D_cache/n1372 ) );
  MX2XL U9992 ( .A(\D_cache/cache[6][52] ), .B(n4549), .S0(n5364), .Y(
        \D_cache/n1374 ) );
  MX2XL U9993 ( .A(\D_cache/cache[5][52] ), .B(n4549), .S0(n5340), .Y(
        \D_cache/n1375 ) );
  MX2XL U9994 ( .A(\D_cache/cache[4][52] ), .B(n4549), .S0(n5313), .Y(
        \D_cache/n1376 ) );
  MX2XL U9995 ( .A(\D_cache/cache[3][52] ), .B(n4549), .S0(n5268), .Y(
        \D_cache/n1377 ) );
  MX2XL U9996 ( .A(\D_cache/cache[2][52] ), .B(n4549), .S0(n5228), .Y(
        \D_cache/n1378 ) );
  MX2XL U9997 ( .A(\D_cache/cache[1][52] ), .B(n4549), .S0(n5198), .Y(
        \D_cache/n1379 ) );
  MX2XL U9998 ( .A(\D_cache/cache[0][52] ), .B(n4549), .S0(n5159), .Y(
        \D_cache/n1380 ) );
  MX2XL U9999 ( .A(\D_cache/cache[6][50] ), .B(n4567), .S0(n5371), .Y(
        \D_cache/n1390 ) );
  MX2XL U10000 ( .A(\D_cache/cache[5][50] ), .B(n4567), .S0(n5347), .Y(
        \D_cache/n1391 ) );
  MX2XL U10001 ( .A(\D_cache/cache[4][50] ), .B(n4567), .S0(n5320), .Y(
        \D_cache/n1392 ) );
  MX2XL U10002 ( .A(\D_cache/cache[3][50] ), .B(n4567), .S0(n5274), .Y(
        \D_cache/n1393 ) );
  MX2XL U10003 ( .A(\D_cache/cache[2][50] ), .B(n4567), .S0(n5233), .Y(
        \D_cache/n1394 ) );
  MX2XL U10004 ( .A(\D_cache/cache[1][50] ), .B(n4567), .S0(n5205), .Y(
        \D_cache/n1395 ) );
  MX2XL U10005 ( .A(\D_cache/cache[0][50] ), .B(n4567), .S0(n3995), .Y(
        \D_cache/n1396 ) );
  MX2XL U10006 ( .A(\D_cache/cache[6][49] ), .B(n4568), .S0(n5371), .Y(
        \D_cache/n1398 ) );
  MX2XL U10007 ( .A(\D_cache/cache[5][49] ), .B(n4568), .S0(n5347), .Y(
        \D_cache/n1399 ) );
  MX2XL U10008 ( .A(\D_cache/cache[4][49] ), .B(n4568), .S0(n5320), .Y(
        \D_cache/n1400 ) );
  MX2XL U10009 ( .A(\D_cache/cache[3][49] ), .B(n4568), .S0(n5274), .Y(
        \D_cache/n1401 ) );
  MX2XL U10010 ( .A(\D_cache/cache[2][49] ), .B(n4568), .S0(n5233), .Y(
        \D_cache/n1402 ) );
  MX2XL U10011 ( .A(\D_cache/cache[1][49] ), .B(n4568), .S0(n5205), .Y(
        \D_cache/n1403 ) );
  MX2XL U10012 ( .A(\D_cache/cache[0][49] ), .B(n4568), .S0(n5164), .Y(
        \D_cache/n1404 ) );
  MX2XL U10013 ( .A(\D_cache/cache[6][48] ), .B(n4550), .S0(n5365), .Y(
        \D_cache/n1406 ) );
  MX2XL U10014 ( .A(\D_cache/cache[5][48] ), .B(n4550), .S0(n5341), .Y(
        \D_cache/n1407 ) );
  MX2XL U10015 ( .A(\D_cache/cache[4][48] ), .B(n4550), .S0(n5314), .Y(
        \D_cache/n1408 ) );
  MX2XL U10016 ( .A(\D_cache/cache[3][48] ), .B(n4550), .S0(n5269), .Y(
        \D_cache/n1409 ) );
  MX2XL U10017 ( .A(\D_cache/cache[2][48] ), .B(n4550), .S0(n5234), .Y(
        \D_cache/n1410 ) );
  MX2XL U10018 ( .A(\D_cache/cache[1][48] ), .B(n4550), .S0(n5199), .Y(
        \D_cache/n1411 ) );
  MX2XL U10019 ( .A(\D_cache/cache[0][48] ), .B(n4550), .S0(n5160), .Y(
        \D_cache/n1412 ) );
  MX2XL U10020 ( .A(\D_cache/cache[6][47] ), .B(n4551), .S0(n5365), .Y(
        \D_cache/n1414 ) );
  MX2XL U10021 ( .A(\D_cache/cache[5][47] ), .B(n4551), .S0(n5341), .Y(
        \D_cache/n1415 ) );
  MX2XL U10022 ( .A(\D_cache/cache[4][47] ), .B(n4551), .S0(n5314), .Y(
        \D_cache/n1416 ) );
  MX2XL U10023 ( .A(\D_cache/cache[3][47] ), .B(n4551), .S0(n5269), .Y(
        \D_cache/n1417 ) );
  MX2XL U10024 ( .A(\D_cache/cache[2][47] ), .B(n4551), .S0(n5231), .Y(
        \D_cache/n1418 ) );
  MX2XL U10025 ( .A(\D_cache/cache[1][47] ), .B(n4551), .S0(n5199), .Y(
        \D_cache/n1419 ) );
  MX2XL U10026 ( .A(\D_cache/cache[0][47] ), .B(n4551), .S0(n5160), .Y(
        \D_cache/n1420 ) );
  MX2XL U10027 ( .A(\D_cache/cache[6][46] ), .B(n4560), .S0(n5366), .Y(
        \D_cache/n1422 ) );
  MX2XL U10028 ( .A(\D_cache/cache[5][46] ), .B(n4560), .S0(n5342), .Y(
        \D_cache/n1423 ) );
  MX2XL U10029 ( .A(\D_cache/cache[4][46] ), .B(n4560), .S0(n5315), .Y(
        \D_cache/n1424 ) );
  MX2XL U10030 ( .A(\D_cache/cache[3][46] ), .B(n4560), .S0(n5270), .Y(
        \D_cache/n1425 ) );
  MX2XL U10031 ( .A(\D_cache/cache[2][46] ), .B(n4560), .S0(n5234), .Y(
        \D_cache/n1426 ) );
  MX2XL U10032 ( .A(\D_cache/cache[1][46] ), .B(n4560), .S0(n5200), .Y(
        \D_cache/n1427 ) );
  MX2XL U10033 ( .A(\D_cache/cache[0][46] ), .B(n4560), .S0(n5164), .Y(
        \D_cache/n1428 ) );
  MX2XL U10034 ( .A(\D_cache/cache[6][44] ), .B(n4552), .S0(n5365), .Y(
        \D_cache/n1438 ) );
  MX2XL U10035 ( .A(\D_cache/cache[5][44] ), .B(n4552), .S0(n5341), .Y(
        \D_cache/n1439 ) );
  MX2XL U10036 ( .A(\D_cache/cache[4][44] ), .B(n4552), .S0(n5314), .Y(
        \D_cache/n1440 ) );
  MX2XL U10037 ( .A(\D_cache/cache[3][44] ), .B(n4552), .S0(n5269), .Y(
        \D_cache/n1441 ) );
  MX2XL U10038 ( .A(\D_cache/cache[2][44] ), .B(n4552), .S0(n5235), .Y(
        \D_cache/n1442 ) );
  MX2XL U10039 ( .A(\D_cache/cache[1][44] ), .B(n4552), .S0(n5199), .Y(
        \D_cache/n1443 ) );
  MX2XL U10040 ( .A(\D_cache/cache[0][44] ), .B(n4552), .S0(n5160), .Y(
        \D_cache/n1444 ) );
  MX2XL U10041 ( .A(\D_cache/cache[6][41] ), .B(n4569), .S0(n5371), .Y(
        \D_cache/n1462 ) );
  MX2XL U10042 ( .A(\D_cache/cache[5][41] ), .B(n4569), .S0(n5347), .Y(
        \D_cache/n1463 ) );
  MX2XL U10043 ( .A(\D_cache/cache[4][41] ), .B(n4569), .S0(n5320), .Y(
        \D_cache/n1464 ) );
  MX2XL U10044 ( .A(\D_cache/cache[3][41] ), .B(n4569), .S0(n5274), .Y(
        \D_cache/n1465 ) );
  MX2XL U10045 ( .A(\D_cache/cache[2][41] ), .B(n4569), .S0(n5233), .Y(
        \D_cache/n1466 ) );
  MX2XL U10046 ( .A(\D_cache/cache[1][41] ), .B(n4569), .S0(n5205), .Y(
        \D_cache/n1467 ) );
  MX2XL U10047 ( .A(\D_cache/cache[6][40] ), .B(n4570), .S0(n5368), .Y(
        \D_cache/n1470 ) );
  MX2XL U10048 ( .A(\D_cache/cache[5][40] ), .B(n4570), .S0(n5344), .Y(
        \D_cache/n1471 ) );
  MX2XL U10049 ( .A(\D_cache/cache[4][40] ), .B(n4570), .S0(n5317), .Y(
        \D_cache/n1472 ) );
  MX2XL U10050 ( .A(\D_cache/cache[3][40] ), .B(n4570), .S0(n5272), .Y(
        \D_cache/n1473 ) );
  MX2XL U10051 ( .A(\D_cache/cache[2][40] ), .B(n4570), .S0(n5230), .Y(
        \D_cache/n1474 ) );
  MX2XL U10052 ( .A(\D_cache/cache[1][40] ), .B(n4570), .S0(n5202), .Y(
        \D_cache/n1475 ) );
  MX2XL U10053 ( .A(\D_cache/cache[0][40] ), .B(n4570), .S0(n5162), .Y(
        \D_cache/n1476 ) );
  MX2XL U10054 ( .A(\D_cache/cache[6][39] ), .B(n10679), .S0(n5368), .Y(
        \D_cache/n1478 ) );
  MX2XL U10055 ( .A(\D_cache/cache[5][39] ), .B(n10679), .S0(n5344), .Y(
        \D_cache/n1479 ) );
  MX2XL U10056 ( .A(\D_cache/cache[4][39] ), .B(n10679), .S0(n5317), .Y(
        \D_cache/n1480 ) );
  MX2XL U10057 ( .A(\D_cache/cache[3][39] ), .B(n10679), .S0(n5272), .Y(
        \D_cache/n1481 ) );
  MX2XL U10058 ( .A(\D_cache/cache[2][39] ), .B(n10679), .S0(n5230), .Y(
        \D_cache/n1482 ) );
  MX2XL U10059 ( .A(\D_cache/cache[1][39] ), .B(n10679), .S0(n5201), .Y(
        \D_cache/n1483 ) );
  MX2XL U10060 ( .A(\D_cache/cache[0][39] ), .B(n10679), .S0(n5161), .Y(
        \D_cache/n1484 ) );
  MX2XL U10061 ( .A(\D_cache/cache[6][38] ), .B(n9949), .S0(n5366), .Y(
        \D_cache/n1486 ) );
  MX2XL U10062 ( .A(\D_cache/cache[5][38] ), .B(n9949), .S0(n5342), .Y(
        \D_cache/n1487 ) );
  MX2XL U10063 ( .A(\D_cache/cache[4][38] ), .B(n9949), .S0(n5315), .Y(
        \D_cache/n1488 ) );
  MX2XL U10064 ( .A(\D_cache/cache[3][38] ), .B(n9949), .S0(n5270), .Y(
        \D_cache/n1489 ) );
  MX2XL U10065 ( .A(\D_cache/cache[2][38] ), .B(n9949), .S0(n5235), .Y(
        \D_cache/n1490 ) );
  MX2XL U10066 ( .A(\D_cache/cache[1][38] ), .B(n9949), .S0(n5200), .Y(
        \D_cache/n1491 ) );
  MX2XL U10067 ( .A(\D_cache/cache[0][38] ), .B(n9949), .S0(n3564), .Y(
        \D_cache/n1492 ) );
  MX2XL U10068 ( .A(\D_cache/cache[6][34] ), .B(n10191), .S0(n5366), .Y(
        \D_cache/n1518 ) );
  MX2XL U10069 ( .A(\D_cache/cache[5][34] ), .B(n10191), .S0(n5342), .Y(
        \D_cache/n1519 ) );
  MX2XL U10070 ( .A(\D_cache/cache[4][34] ), .B(n10191), .S0(n5315), .Y(
        \D_cache/n1520 ) );
  MX2XL U10071 ( .A(\D_cache/cache[3][34] ), .B(n10191), .S0(n5270), .Y(
        \D_cache/n1521 ) );
  MX2XL U10072 ( .A(\D_cache/cache[2][34] ), .B(n10191), .S0(n5230), .Y(
        \D_cache/n1522 ) );
  MX2XL U10073 ( .A(\D_cache/cache[1][34] ), .B(n10191), .S0(n5200), .Y(
        \D_cache/n1523 ) );
  MX2XL U10074 ( .A(\D_cache/cache[0][34] ), .B(n10191), .S0(n5161), .Y(
        \D_cache/n1524 ) );
  MX2XL U10075 ( .A(\D_cache/cache[6][33] ), .B(n10666), .S0(n5368), .Y(
        \D_cache/n1526 ) );
  MX2XL U10076 ( .A(\D_cache/cache[5][33] ), .B(n10666), .S0(n5344), .Y(
        \D_cache/n1527 ) );
  MX2XL U10077 ( .A(\D_cache/cache[4][33] ), .B(n10666), .S0(n5317), .Y(
        \D_cache/n1528 ) );
  MX2XL U10078 ( .A(\D_cache/cache[3][33] ), .B(n10666), .S0(n5272), .Y(
        \D_cache/n1529 ) );
  MX2XL U10079 ( .A(\D_cache/cache[2][33] ), .B(n10666), .S0(n5230), .Y(
        \D_cache/n1530 ) );
  MX2XL U10080 ( .A(\D_cache/cache[1][33] ), .B(n10666), .S0(n5202), .Y(
        \D_cache/n1531 ) );
  MX2XL U10081 ( .A(\D_cache/cache[0][33] ), .B(n10666), .S0(n5162), .Y(
        \D_cache/n1532 ) );
  MX2XL U10082 ( .A(\D_cache/cache[6][30] ), .B(n4571), .S0(n5370), .Y(
        \D_cache/n1550 ) );
  MX2XL U10083 ( .A(\D_cache/cache[5][30] ), .B(n4571), .S0(n5346), .Y(
        \D_cache/n1551 ) );
  MX2XL U10084 ( .A(\D_cache/cache[4][30] ), .B(n4571), .S0(n5319), .Y(
        \D_cache/n1552 ) );
  MX2XL U10085 ( .A(\D_cache/cache[3][30] ), .B(n4571), .S0(n5272), .Y(
        \D_cache/n1553 ) );
  MX2XL U10086 ( .A(\D_cache/cache[2][30] ), .B(n4571), .S0(n5232), .Y(
        \D_cache/n1554 ) );
  MX2XL U10087 ( .A(\D_cache/cache[1][30] ), .B(n4571), .S0(n5204), .Y(
        \D_cache/n1555 ) );
  MX2XL U10088 ( .A(\D_cache/cache[0][30] ), .B(n4571), .S0(n5163), .Y(
        \D_cache/n1556 ) );
  MX2XL U10089 ( .A(\D_cache/cache[6][29] ), .B(n4572), .S0(n5370), .Y(
        \D_cache/n1558 ) );
  MX2XL U10090 ( .A(\D_cache/cache[5][29] ), .B(n4572), .S0(n5346), .Y(
        \D_cache/n1559 ) );
  MX2XL U10091 ( .A(\D_cache/cache[4][29] ), .B(n4572), .S0(n5319), .Y(
        \D_cache/n1560 ) );
  MX2XL U10092 ( .A(\D_cache/cache[3][29] ), .B(n4572), .S0(n5273), .Y(
        \D_cache/n1561 ) );
  MX2XL U10093 ( .A(\D_cache/cache[2][29] ), .B(n4572), .S0(n5232), .Y(
        \D_cache/n1562 ) );
  MX2XL U10094 ( .A(\D_cache/cache[1][29] ), .B(n4572), .S0(n5204), .Y(
        \D_cache/n1563 ) );
  MX2XL U10095 ( .A(\D_cache/cache[0][29] ), .B(n4572), .S0(n3565), .Y(
        \D_cache/n1564 ) );
  MX2XL U10096 ( .A(\D_cache/cache[6][28] ), .B(n4573), .S0(n5370), .Y(
        \D_cache/n1566 ) );
  MX2XL U10097 ( .A(\D_cache/cache[5][28] ), .B(n4573), .S0(n5346), .Y(
        \D_cache/n1567 ) );
  MX2XL U10098 ( .A(\D_cache/cache[4][28] ), .B(n4573), .S0(n5319), .Y(
        \D_cache/n1568 ) );
  MX2XL U10099 ( .A(\D_cache/cache[3][28] ), .B(n4573), .S0(n5270), .Y(
        \D_cache/n1569 ) );
  MX2XL U10100 ( .A(\D_cache/cache[2][28] ), .B(n4573), .S0(n5232), .Y(
        \D_cache/n1570 ) );
  MX2XL U10101 ( .A(\D_cache/cache[1][28] ), .B(n4573), .S0(n5204), .Y(
        \D_cache/n1571 ) );
  MX2XL U10102 ( .A(\D_cache/cache[0][28] ), .B(n4573), .S0(n3995), .Y(
        \D_cache/n1572 ) );
  MX2XL U10103 ( .A(\D_cache/cache[6][27] ), .B(n10393), .S0(n5367), .Y(
        \D_cache/n1574 ) );
  MX2XL U10104 ( .A(\D_cache/cache[5][27] ), .B(n10393), .S0(n5343), .Y(
        \D_cache/n1575 ) );
  MX2XL U10105 ( .A(\D_cache/cache[4][27] ), .B(n10393), .S0(n5316), .Y(
        \D_cache/n1576 ) );
  MX2XL U10106 ( .A(\D_cache/cache[3][27] ), .B(n10393), .S0(n5271), .Y(
        \D_cache/n1577 ) );
  MX2XL U10107 ( .A(\D_cache/cache[2][27] ), .B(n10393), .S0(n5229), .Y(
        \D_cache/n1578 ) );
  MX2XL U10108 ( .A(\D_cache/cache[1][27] ), .B(n10393), .S0(n5201), .Y(
        \D_cache/n1579 ) );
  MX2XL U10109 ( .A(\D_cache/cache[6][26] ), .B(n10200), .S0(n5367), .Y(
        \D_cache/n1582 ) );
  MX2XL U10110 ( .A(\D_cache/cache[5][26] ), .B(n10200), .S0(n5343), .Y(
        \D_cache/n1583 ) );
  MX2XL U10111 ( .A(\D_cache/cache[4][26] ), .B(n10200), .S0(n5316), .Y(
        \D_cache/n1584 ) );
  MX2XL U10112 ( .A(\D_cache/cache[3][26] ), .B(n10200), .S0(n5271), .Y(
        \D_cache/n1585 ) );
  MX2XL U10113 ( .A(\D_cache/cache[2][26] ), .B(n10200), .S0(n5229), .Y(
        \D_cache/n1586 ) );
  MX2XL U10114 ( .A(\D_cache/cache[1][26] ), .B(n10200), .S0(n5201), .Y(
        \D_cache/n1587 ) );
  MX2XL U10115 ( .A(\D_cache/cache[0][26] ), .B(n10200), .S0(n5161), .Y(
        \D_cache/n1588 ) );
  MX2XL U10116 ( .A(\D_cache/cache[6][25] ), .B(n4555), .S0(n5364), .Y(
        \D_cache/n1590 ) );
  MX2XL U10117 ( .A(\D_cache/cache[5][25] ), .B(n4555), .S0(n5340), .Y(
        \D_cache/n1591 ) );
  MX2XL U10118 ( .A(\D_cache/cache[4][25] ), .B(n4555), .S0(n5313), .Y(
        \D_cache/n1592 ) );
  MX2XL U10119 ( .A(\D_cache/cache[3][25] ), .B(n4555), .S0(n5268), .Y(
        \D_cache/n1593 ) );
  MX2XL U10120 ( .A(\D_cache/cache[2][25] ), .B(n4555), .S0(n5228), .Y(
        \D_cache/n1594 ) );
  MX2XL U10121 ( .A(\D_cache/cache[1][25] ), .B(n4555), .S0(n5198), .Y(
        \D_cache/n1595 ) );
  MX2XL U10122 ( .A(\D_cache/cache[0][25] ), .B(n4555), .S0(n5159), .Y(
        \D_cache/n1596 ) );
  MX2XL U10123 ( .A(\D_cache/cache[6][24] ), .B(n4556), .S0(n5364), .Y(
        \D_cache/n1598 ) );
  MX2XL U10124 ( .A(\D_cache/cache[5][24] ), .B(n4556), .S0(n5340), .Y(
        \D_cache/n1599 ) );
  MX2XL U10125 ( .A(\D_cache/cache[4][24] ), .B(n4556), .S0(n5313), .Y(
        \D_cache/n1600 ) );
  MX2XL U10126 ( .A(\D_cache/cache[3][24] ), .B(n4556), .S0(n5268), .Y(
        \D_cache/n1601 ) );
  MX2XL U10127 ( .A(\D_cache/cache[2][24] ), .B(n4556), .S0(n5228), .Y(
        \D_cache/n1602 ) );
  MX2XL U10128 ( .A(\D_cache/cache[1][24] ), .B(n4556), .S0(n5198), .Y(
        \D_cache/n1603 ) );
  MX2XL U10129 ( .A(\D_cache/cache[0][24] ), .B(n4556), .S0(n5159), .Y(
        \D_cache/n1604 ) );
  MX2XL U10130 ( .A(\D_cache/cache[6][22] ), .B(n4559), .S0(n5367), .Y(
        \D_cache/n1614 ) );
  MX2XL U10131 ( .A(\D_cache/cache[5][22] ), .B(n4559), .S0(n5343), .Y(
        \D_cache/n1615 ) );
  MX2XL U10132 ( .A(\D_cache/cache[4][22] ), .B(n4559), .S0(n5316), .Y(
        \D_cache/n1616 ) );
  MX2XL U10133 ( .A(\D_cache/cache[3][22] ), .B(n4559), .S0(n5271), .Y(
        \D_cache/n1617 ) );
  MX2XL U10134 ( .A(\D_cache/cache[2][22] ), .B(n4559), .S0(n5229), .Y(
        \D_cache/n1618 ) );
  MX2XL U10135 ( .A(\D_cache/cache[1][22] ), .B(n4559), .S0(n5201), .Y(
        \D_cache/n1619 ) );
  MX2XL U10136 ( .A(\D_cache/cache[0][22] ), .B(n4559), .S0(n5161), .Y(
        \D_cache/n1620 ) );
  MX2XL U10137 ( .A(\D_cache/cache[6][21] ), .B(n10516), .S0(n5365), .Y(
        \D_cache/n1622 ) );
  MX2XL U10138 ( .A(\D_cache/cache[5][21] ), .B(n10516), .S0(n5341), .Y(
        \D_cache/n1623 ) );
  MX2XL U10139 ( .A(\D_cache/cache[4][21] ), .B(n10516), .S0(n5314), .Y(
        \D_cache/n1624 ) );
  MX2XL U10140 ( .A(\D_cache/cache[3][21] ), .B(n10516), .S0(n5269), .Y(
        \D_cache/n1625 ) );
  MX2XL U10141 ( .A(\D_cache/cache[2][21] ), .B(n10516), .S0(n5230), .Y(
        \D_cache/n1626 ) );
  MX2XL U10142 ( .A(\D_cache/cache[1][21] ), .B(n10516), .S0(n5199), .Y(
        \D_cache/n1627 ) );
  MX2XL U10143 ( .A(\D_cache/cache[0][21] ), .B(n10516), .S0(n5164), .Y(
        \D_cache/n1628 ) );
  MX2XL U10144 ( .A(\D_cache/cache[6][20] ), .B(n4557), .S0(n5364), .Y(
        \D_cache/n1630 ) );
  MX2XL U10145 ( .A(\D_cache/cache[5][20] ), .B(n4557), .S0(n5340), .Y(
        \D_cache/n1631 ) );
  MX2XL U10146 ( .A(\D_cache/cache[4][20] ), .B(n4557), .S0(n5313), .Y(
        \D_cache/n1632 ) );
  MX2XL U10147 ( .A(\D_cache/cache[3][20] ), .B(n4557), .S0(n5268), .Y(
        \D_cache/n1633 ) );
  MX2XL U10148 ( .A(\D_cache/cache[2][20] ), .B(n4557), .S0(n5228), .Y(
        \D_cache/n1634 ) );
  MX2XL U10149 ( .A(\D_cache/cache[1][20] ), .B(n4557), .S0(n5198), .Y(
        \D_cache/n1635 ) );
  MX2XL U10150 ( .A(\D_cache/cache[0][20] ), .B(n4557), .S0(n5159), .Y(
        \D_cache/n1636 ) );
  MX2XL U10151 ( .A(\D_cache/cache[6][18] ), .B(n4574), .S0(n5371), .Y(
        \D_cache/n1646 ) );
  MX2XL U10152 ( .A(\D_cache/cache[5][18] ), .B(n4574), .S0(n5347), .Y(
        \D_cache/n1647 ) );
  MX2XL U10153 ( .A(\D_cache/cache[4][18] ), .B(n4574), .S0(n5320), .Y(
        \D_cache/n1648 ) );
  MX2XL U10154 ( .A(\D_cache/cache[3][18] ), .B(n4574), .S0(n5274), .Y(
        \D_cache/n1649 ) );
  MX2XL U10155 ( .A(\D_cache/cache[2][18] ), .B(n4574), .S0(n5233), .Y(
        \D_cache/n1650 ) );
  MX2XL U10156 ( .A(\D_cache/cache[1][18] ), .B(n4574), .S0(n5205), .Y(
        \D_cache/n1651 ) );
  MX2XL U10157 ( .A(\D_cache/cache[0][18] ), .B(n4574), .S0(n5164), .Y(
        \D_cache/n1652 ) );
  MX2XL U10158 ( .A(\D_cache/cache[6][17] ), .B(n2995), .S0(n5371), .Y(
        \D_cache/n1654 ) );
  MX2XL U10159 ( .A(\D_cache/cache[5][17] ), .B(n2995), .S0(n5347), .Y(
        \D_cache/n1655 ) );
  MX2XL U10160 ( .A(\D_cache/cache[4][17] ), .B(n2995), .S0(n5320), .Y(
        \D_cache/n1656 ) );
  MX2XL U10161 ( .A(\D_cache/cache[3][17] ), .B(n2995), .S0(n5274), .Y(
        \D_cache/n1657 ) );
  MX2XL U10162 ( .A(\D_cache/cache[2][17] ), .B(n2995), .S0(n5233), .Y(
        \D_cache/n1658 ) );
  MX2XL U10163 ( .A(\D_cache/cache[1][17] ), .B(n2995), .S0(n5205), .Y(
        \D_cache/n1659 ) );
  MX2XL U10164 ( .A(\D_cache/cache[0][17] ), .B(n2995), .S0(n5164), .Y(
        \D_cache/n1660 ) );
  MX2XL U10165 ( .A(\D_cache/cache[6][16] ), .B(n146), .S0(n5365), .Y(
        \D_cache/n1662 ) );
  MX2XL U10166 ( .A(\D_cache/cache[5][16] ), .B(n146), .S0(n5341), .Y(
        \D_cache/n1663 ) );
  MX2XL U10167 ( .A(\D_cache/cache[4][16] ), .B(n146), .S0(n5314), .Y(
        \D_cache/n1664 ) );
  MX2XL U10168 ( .A(\D_cache/cache[3][16] ), .B(n146), .S0(n5269), .Y(
        \D_cache/n1665 ) );
  MX2XL U10169 ( .A(\D_cache/cache[2][16] ), .B(n146), .S0(n5234), .Y(
        \D_cache/n1666 ) );
  MX2XL U10170 ( .A(\D_cache/cache[1][16] ), .B(n146), .S0(n5199), .Y(
        \D_cache/n1667 ) );
  MX2XL U10171 ( .A(\D_cache/cache[0][16] ), .B(n146), .S0(n5160), .Y(
        \D_cache/n1668 ) );
  MX2XL U10172 ( .A(\D_cache/cache[6][15] ), .B(n4558), .S0(n5369), .Y(
        \D_cache/n1670 ) );
  MX2XL U10173 ( .A(\D_cache/cache[5][15] ), .B(n4558), .S0(n3575), .Y(
        \D_cache/n1671 ) );
  MX2XL U10174 ( .A(\D_cache/cache[4][15] ), .B(n4558), .S0(n5318), .Y(
        \D_cache/n1672 ) );
  MX2XL U10175 ( .A(\D_cache/cache[3][15] ), .B(n4558), .S0(n5273), .Y(
        \D_cache/n1673 ) );
  MX2XL U10176 ( .A(\D_cache/cache[2][15] ), .B(n4558), .S0(n5231), .Y(
        \D_cache/n1674 ) );
  MX2XL U10177 ( .A(\D_cache/cache[1][15] ), .B(n4558), .S0(n5199), .Y(
        \D_cache/n1675 ) );
  MX2XL U10178 ( .A(\D_cache/cache[0][15] ), .B(n4558), .S0(n5160), .Y(
        \D_cache/n1676 ) );
  MX2XL U10179 ( .A(\D_cache/cache[6][14] ), .B(n10100), .S0(n5366), .Y(
        \D_cache/n1678 ) );
  MX2XL U10180 ( .A(\D_cache/cache[5][14] ), .B(n10100), .S0(n5342), .Y(
        \D_cache/n1679 ) );
  MX2XL U10181 ( .A(\D_cache/cache[4][14] ), .B(n10100), .S0(n5315), .Y(
        \D_cache/n1680 ) );
  MX2XL U10182 ( .A(\D_cache/cache[3][14] ), .B(n10100), .S0(n5270), .Y(
        \D_cache/n1681 ) );
  MX2XL U10183 ( .A(\D_cache/cache[2][14] ), .B(n10100), .S0(n5228), .Y(
        \D_cache/n1682 ) );
  MX2XL U10184 ( .A(\D_cache/cache[1][14] ), .B(n10100), .S0(n5200), .Y(
        \D_cache/n1683 ) );
  MX2XL U10185 ( .A(\D_cache/cache[0][14] ), .B(n10100), .S0(n5164), .Y(
        \D_cache/n1684 ) );
  MX2XL U10186 ( .A(\D_cache/cache[6][12] ), .B(n4575), .S0(n5365), .Y(
        \D_cache/n1694 ) );
  MX2XL U10187 ( .A(\D_cache/cache[5][12] ), .B(n4575), .S0(n5341), .Y(
        \D_cache/n1695 ) );
  MX2XL U10188 ( .A(\D_cache/cache[4][12] ), .B(n4575), .S0(n5314), .Y(
        \D_cache/n1696 ) );
  MX2XL U10189 ( .A(\D_cache/cache[3][12] ), .B(n4575), .S0(n5269), .Y(
        \D_cache/n1697 ) );
  MX2XL U10190 ( .A(\D_cache/cache[2][12] ), .B(n4575), .S0(n5233), .Y(
        \D_cache/n1698 ) );
  MX2XL U10191 ( .A(\D_cache/cache[1][12] ), .B(n4575), .S0(n5199), .Y(
        \D_cache/n1699 ) );
  MX2XL U10192 ( .A(\D_cache/cache[0][12] ), .B(n4575), .S0(n5160), .Y(
        \D_cache/n1700 ) );
  MX2XL U10193 ( .A(\D_cache/cache[6][9] ), .B(n4576), .S0(n5371), .Y(
        \D_cache/n1718 ) );
  MX2XL U10194 ( .A(\D_cache/cache[5][9] ), .B(n4576), .S0(n5347), .Y(
        \D_cache/n1719 ) );
  MX2XL U10195 ( .A(\D_cache/cache[4][9] ), .B(n4576), .S0(n5320), .Y(
        \D_cache/n1720 ) );
  MX2XL U10196 ( .A(\D_cache/cache[3][9] ), .B(n4576), .S0(n5274), .Y(
        \D_cache/n1721 ) );
  MX2XL U10197 ( .A(\D_cache/cache[2][9] ), .B(n4576), .S0(n5233), .Y(
        \D_cache/n1722 ) );
  MX2XL U10198 ( .A(\D_cache/cache[1][9] ), .B(n4576), .S0(n5205), .Y(
        \D_cache/n1723 ) );
  MX2XL U10199 ( .A(\D_cache/cache[0][9] ), .B(n4576), .S0(n5164), .Y(
        \D_cache/n1724 ) );
  MX2XL U10200 ( .A(\D_cache/cache[6][8] ), .B(n10649), .S0(n5368), .Y(
        \D_cache/n1726 ) );
  MX2XL U10201 ( .A(\D_cache/cache[5][8] ), .B(n10649), .S0(n5344), .Y(
        \D_cache/n1727 ) );
  MX2XL U10202 ( .A(\D_cache/cache[4][8] ), .B(n10649), .S0(n5317), .Y(
        \D_cache/n1728 ) );
  MX2XL U10203 ( .A(\D_cache/cache[3][8] ), .B(n10649), .S0(n5272), .Y(
        \D_cache/n1729 ) );
  MX2XL U10204 ( .A(\D_cache/cache[2][8] ), .B(n10649), .S0(n5230), .Y(
        \D_cache/n1730 ) );
  MX2XL U10205 ( .A(\D_cache/cache[1][8] ), .B(n10649), .S0(n5202), .Y(
        \D_cache/n1731 ) );
  MX2XL U10206 ( .A(\D_cache/cache[0][8] ), .B(n10649), .S0(n5162), .Y(
        \D_cache/n1732 ) );
  MX2XL U10207 ( .A(\D_cache/cache[6][7] ), .B(n4577), .S0(n5368), .Y(
        \D_cache/n1734 ) );
  MX2XL U10208 ( .A(\D_cache/cache[5][7] ), .B(n4577), .S0(n5344), .Y(
        \D_cache/n1735 ) );
  MX2XL U10209 ( .A(\D_cache/cache[4][7] ), .B(n4577), .S0(n5317), .Y(
        \D_cache/n1736 ) );
  MX2XL U10210 ( .A(\D_cache/cache[3][7] ), .B(n4577), .S0(n5272), .Y(
        \D_cache/n1737 ) );
  MX2XL U10211 ( .A(\D_cache/cache[2][7] ), .B(n4577), .S0(n5230), .Y(
        \D_cache/n1738 ) );
  MX2XL U10212 ( .A(\D_cache/cache[1][7] ), .B(n4577), .S0(n5202), .Y(
        \D_cache/n1739 ) );
  MX2XL U10213 ( .A(\D_cache/cache[0][7] ), .B(n4577), .S0(n5161), .Y(
        \D_cache/n1740 ) );
  MX2XL U10214 ( .A(\D_cache/cache[6][6] ), .B(n9942), .S0(n5366), .Y(
        \D_cache/n1742 ) );
  MX2XL U10215 ( .A(\D_cache/cache[5][6] ), .B(n9942), .S0(n5342), .Y(
        \D_cache/n1743 ) );
  MX2XL U10216 ( .A(\D_cache/cache[4][6] ), .B(n9942), .S0(n5315), .Y(
        \D_cache/n1744 ) );
  MX2XL U10217 ( .A(\D_cache/cache[3][6] ), .B(n9942), .S0(n5270), .Y(
        \D_cache/n1745 ) );
  MX2XL U10218 ( .A(\D_cache/cache[2][6] ), .B(n9942), .S0(n5231), .Y(
        \D_cache/n1746 ) );
  MX2XL U10219 ( .A(\D_cache/cache[1][6] ), .B(n9942), .S0(n5200), .Y(
        \D_cache/n1747 ) );
  MX2XL U10220 ( .A(\D_cache/cache[6][4] ), .B(n9810), .S0(n5372), .Y(
        \D_cache/n1758 ) );
  MX2XL U10221 ( .A(\D_cache/cache[5][4] ), .B(n9810), .S0(n5349), .Y(
        \D_cache/n1759 ) );
  MX2XL U10222 ( .A(\D_cache/cache[4][4] ), .B(n9810), .S0(n5321), .Y(
        \D_cache/n1760 ) );
  MX2XL U10223 ( .A(\D_cache/cache[3][4] ), .B(n9810), .S0(n5276), .Y(
        \D_cache/n1761 ) );
  MX2XL U10224 ( .A(\D_cache/cache[2][4] ), .B(n9810), .S0(n5232), .Y(
        \D_cache/n1762 ) );
  MX2XL U10225 ( .A(\D_cache/cache[1][4] ), .B(n9810), .S0(n5200), .Y(
        \D_cache/n1763 ) );
  MX2XL U10226 ( .A(\D_cache/cache[3][3] ), .B(n4561), .S0(n5275), .Y(
        \D_cache/n1769 ) );
  MX2XL U10227 ( .A(\D_cache/cache[2][3] ), .B(n4561), .S0(n5235), .Y(
        \D_cache/n1770 ) );
  MX2XL U10228 ( .A(\D_cache/cache[1][3] ), .B(n4561), .S0(n5204), .Y(
        \D_cache/n1771 ) );
  MX2XL U10229 ( .A(\D_cache/cache[0][3] ), .B(n4561), .S0(n3565), .Y(
        \D_cache/n1772 ) );
  MX2XL U10230 ( .A(\D_cache/cache[6][2] ), .B(n10188), .S0(n5366), .Y(
        \D_cache/n1774 ) );
  MX2XL U10231 ( .A(\D_cache/cache[5][2] ), .B(n10188), .S0(n5342), .Y(
        \D_cache/n1775 ) );
  MX2XL U10232 ( .A(\D_cache/cache[4][2] ), .B(n10188), .S0(n5315), .Y(
        \D_cache/n1776 ) );
  MX2XL U10233 ( .A(\D_cache/cache[3][2] ), .B(n10188), .S0(n5270), .Y(
        \D_cache/n1777 ) );
  MX2XL U10234 ( .A(\D_cache/cache[2][2] ), .B(n10188), .S0(n5234), .Y(
        \D_cache/n1778 ) );
  MX2XL U10235 ( .A(\D_cache/cache[1][2] ), .B(n10188), .S0(n5200), .Y(
        \D_cache/n1779 ) );
  MX2XL U10236 ( .A(\D_cache/cache[6][1] ), .B(n10663), .S0(n5368), .Y(
        \D_cache/n1782 ) );
  MX2XL U10237 ( .A(\D_cache/cache[5][1] ), .B(n10663), .S0(n5344), .Y(
        \D_cache/n1783 ) );
  MX2XL U10238 ( .A(\D_cache/cache[4][1] ), .B(n10663), .S0(n5317), .Y(
        \D_cache/n1784 ) );
  MX2XL U10239 ( .A(\D_cache/cache[3][1] ), .B(n10663), .S0(n5272), .Y(
        \D_cache/n1785 ) );
  MX2XL U10240 ( .A(\D_cache/cache[2][1] ), .B(n10663), .S0(n5230), .Y(
        \D_cache/n1786 ) );
  MX2XL U10241 ( .A(\D_cache/cache[1][1] ), .B(n10663), .S0(n5202), .Y(
        \D_cache/n1787 ) );
  MX2XL U10242 ( .A(\D_cache/cache[0][1] ), .B(n10663), .S0(n5162), .Y(
        \D_cache/n1788 ) );
  MX2XL U10243 ( .A(\D_cache/cache[6][95] ), .B(n10710), .S0(n5369), .Y(
        \D_cache/n1030 ) );
  MX2XL U10244 ( .A(\D_cache/cache[5][95] ), .B(n10710), .S0(n3575), .Y(
        \D_cache/n1031 ) );
  MX2XL U10245 ( .A(\D_cache/cache[4][95] ), .B(n10710), .S0(n5318), .Y(
        \D_cache/n1032 ) );
  MX2XL U10246 ( .A(\D_cache/cache[3][95] ), .B(n10710), .S0(n5273), .Y(
        \D_cache/n1033 ) );
  MX2XL U10247 ( .A(\D_cache/cache[2][95] ), .B(n10710), .S0(n5231), .Y(
        \D_cache/n1034 ) );
  MX2XL U10248 ( .A(\D_cache/cache[1][95] ), .B(n10710), .S0(n5203), .Y(
        \D_cache/n1035 ) );
  MX2XL U10249 ( .A(\D_cache/cache[0][95] ), .B(n10710), .S0(n5163), .Y(
        \D_cache/n1036 ) );
  MX2XL U10250 ( .A(\D_cache/cache[6][94] ), .B(n10603), .S0(n5371), .Y(
        \D_cache/n1038 ) );
  MX2XL U10251 ( .A(\D_cache/cache[5][94] ), .B(n10603), .S0(n5347), .Y(
        \D_cache/n1039 ) );
  MX2XL U10252 ( .A(\D_cache/cache[4][94] ), .B(n10603), .S0(n5320), .Y(
        \D_cache/n1040 ) );
  MX2XL U10253 ( .A(\D_cache/cache[3][94] ), .B(n10603), .S0(n5274), .Y(
        \D_cache/n1041 ) );
  MX2XL U10254 ( .A(\D_cache/cache[2][94] ), .B(n10603), .S0(n5233), .Y(
        \D_cache/n1042 ) );
  MX2XL U10255 ( .A(\D_cache/cache[1][94] ), .B(n10603), .S0(n5205), .Y(
        \D_cache/n1043 ) );
  MX2XL U10256 ( .A(\D_cache/cache[0][94] ), .B(n10603), .S0(n5164), .Y(
        \D_cache/n1044 ) );
  MX2XL U10257 ( .A(\D_cache/cache[6][93] ), .B(n10566), .S0(n5370), .Y(
        \D_cache/n1046 ) );
  MX2XL U10258 ( .A(\D_cache/cache[5][93] ), .B(n10566), .S0(n5346), .Y(
        \D_cache/n1047 ) );
  MX2XL U10259 ( .A(\D_cache/cache[4][93] ), .B(n10566), .S0(n5319), .Y(
        \D_cache/n1048 ) );
  MX2XL U10260 ( .A(\D_cache/cache[3][93] ), .B(n10566), .S0(n5268), .Y(
        \D_cache/n1049 ) );
  MX2XL U10261 ( .A(\D_cache/cache[2][93] ), .B(n10566), .S0(n5232), .Y(
        \D_cache/n1050 ) );
  MX2XL U10262 ( .A(\D_cache/cache[1][93] ), .B(n10566), .S0(n5204), .Y(
        \D_cache/n1051 ) );
  MX2XL U10263 ( .A(\D_cache/cache[0][93] ), .B(n10566), .S0(n3995), .Y(
        \D_cache/n1052 ) );
  MX2XL U10264 ( .A(\D_cache/cache[6][92] ), .B(n10553), .S0(n5370), .Y(
        \D_cache/n1054 ) );
  MX2XL U10265 ( .A(\D_cache/cache[5][92] ), .B(n10553), .S0(n5346), .Y(
        \D_cache/n1055 ) );
  MX2XL U10266 ( .A(\D_cache/cache[4][92] ), .B(n10553), .S0(n5319), .Y(
        \D_cache/n1056 ) );
  MX2XL U10267 ( .A(\D_cache/cache[3][92] ), .B(n10553), .S0(n5269), .Y(
        \D_cache/n1057 ) );
  MX2XL U10268 ( .A(\D_cache/cache[2][92] ), .B(n10553), .S0(n5232), .Y(
        \D_cache/n1058 ) );
  MX2XL U10269 ( .A(\D_cache/cache[1][92] ), .B(n10553), .S0(n5204), .Y(
        \D_cache/n1059 ) );
  MX2XL U10270 ( .A(\D_cache/cache[0][92] ), .B(n10553), .S0(n5168), .Y(
        \D_cache/n1060 ) );
  MX2XL U10271 ( .A(\D_cache/cache[6][91] ), .B(n4511), .S0(n5366), .Y(
        \D_cache/n1062 ) );
  MX2XL U10272 ( .A(\D_cache/cache[5][91] ), .B(n4511), .S0(n5342), .Y(
        \D_cache/n1063 ) );
  MX2XL U10273 ( .A(\D_cache/cache[4][91] ), .B(n4511), .S0(n5315), .Y(
        \D_cache/n1064 ) );
  MX2XL U10274 ( .A(\D_cache/cache[3][91] ), .B(n4511), .S0(n5270), .Y(
        \D_cache/n1065 ) );
  MX2XL U10275 ( .A(\D_cache/cache[2][91] ), .B(n4511), .S0(n5235), .Y(
        \D_cache/n1066 ) );
  MX2XL U10276 ( .A(\D_cache/cache[1][91] ), .B(n4511), .S0(n5198), .Y(
        \D_cache/n1067 ) );
  MX2XL U10277 ( .A(\D_cache/cache[0][91] ), .B(n4511), .S0(n5159), .Y(
        \D_cache/n1068 ) );
  MX2XL U10278 ( .A(\D_cache/cache[6][90] ), .B(n10209), .S0(n5367), .Y(
        \D_cache/n1070 ) );
  MX2XL U10279 ( .A(\D_cache/cache[5][90] ), .B(n10209), .S0(n5343), .Y(
        \D_cache/n1071 ) );
  MX2XL U10280 ( .A(\D_cache/cache[4][90] ), .B(n10209), .S0(n5316), .Y(
        \D_cache/n1072 ) );
  MX2XL U10281 ( .A(\D_cache/cache[3][90] ), .B(n10209), .S0(n5271), .Y(
        \D_cache/n1073 ) );
  MX2XL U10282 ( .A(\D_cache/cache[2][90] ), .B(n10209), .S0(n5229), .Y(
        \D_cache/n1074 ) );
  MX2XL U10283 ( .A(\D_cache/cache[1][90] ), .B(n10209), .S0(n5201), .Y(
        \D_cache/n1075 ) );
  MX2XL U10284 ( .A(\D_cache/cache[0][90] ), .B(n10209), .S0(n5161), .Y(
        \D_cache/n1076 ) );
  MX2XL U10285 ( .A(\D_cache/cache[6][89] ), .B(n10442), .S0(n5364), .Y(
        \D_cache/n1078 ) );
  MX2XL U10286 ( .A(\D_cache/cache[5][89] ), .B(n10442), .S0(n5340), .Y(
        \D_cache/n1079 ) );
  MX2XL U10287 ( .A(\D_cache/cache[4][89] ), .B(n10442), .S0(n5313), .Y(
        \D_cache/n1080 ) );
  MX2XL U10288 ( .A(\D_cache/cache[3][89] ), .B(n10442), .S0(n5268), .Y(
        \D_cache/n1081 ) );
  MX2XL U10289 ( .A(\D_cache/cache[2][89] ), .B(n10442), .S0(n5228), .Y(
        \D_cache/n1082 ) );
  MX2XL U10290 ( .A(\D_cache/cache[1][89] ), .B(n10442), .S0(n5203), .Y(
        \D_cache/n1083 ) );
  MX2XL U10291 ( .A(\D_cache/cache[0][89] ), .B(n10442), .S0(n5160), .Y(
        \D_cache/n1084 ) );
  MX2XL U10292 ( .A(\D_cache/cache[6][88] ), .B(n4512), .S0(n5364), .Y(
        \D_cache/n1086 ) );
  MX2XL U10293 ( .A(\D_cache/cache[5][88] ), .B(n4512), .S0(n5340), .Y(
        \D_cache/n1087 ) );
  MX2XL U10294 ( .A(\D_cache/cache[4][88] ), .B(n4512), .S0(n5313), .Y(
        \D_cache/n1088 ) );
  MX2XL U10295 ( .A(\D_cache/cache[3][88] ), .B(n4512), .S0(n5268), .Y(
        \D_cache/n1089 ) );
  MX2XL U10296 ( .A(\D_cache/cache[2][88] ), .B(n4512), .S0(n5228), .Y(
        \D_cache/n1090 ) );
  MX2XL U10297 ( .A(\D_cache/cache[1][88] ), .B(n4512), .S0(n5198), .Y(
        \D_cache/n1091 ) );
  MX2XL U10298 ( .A(\D_cache/cache[0][88] ), .B(n4512), .S0(n5159), .Y(
        \D_cache/n1092 ) );
  MX2XL U10299 ( .A(\D_cache/cache[6][87] ), .B(n10697), .S0(n5369), .Y(
        \D_cache/n1094 ) );
  MX2XL U10300 ( .A(\D_cache/cache[5][87] ), .B(n10697), .S0(n3575), .Y(
        \D_cache/n1095 ) );
  MX2XL U10301 ( .A(\D_cache/cache[4][87] ), .B(n10697), .S0(n5318), .Y(
        \D_cache/n1096 ) );
  MX2XL U10302 ( .A(\D_cache/cache[3][87] ), .B(n10697), .S0(n5273), .Y(
        \D_cache/n1097 ) );
  MX2XL U10303 ( .A(\D_cache/cache[2][87] ), .B(n10697), .S0(n5231), .Y(
        \D_cache/n1098 ) );
  MX2XL U10304 ( .A(\D_cache/cache[1][87] ), .B(n10697), .S0(n5203), .Y(
        \D_cache/n1099 ) );
  MX2XL U10305 ( .A(\D_cache/cache[0][87] ), .B(n10697), .S0(n5163), .Y(
        \D_cache/n1100 ) );
  MX2XL U10306 ( .A(\D_cache/cache[6][86] ), .B(n10318), .S0(n5367), .Y(
        \D_cache/n1102 ) );
  MX2XL U10307 ( .A(\D_cache/cache[5][86] ), .B(n10318), .S0(n5343), .Y(
        \D_cache/n1103 ) );
  MX2XL U10308 ( .A(\D_cache/cache[4][86] ), .B(n10318), .S0(n5316), .Y(
        \D_cache/n1104 ) );
  MX2XL U10309 ( .A(\D_cache/cache[3][86] ), .B(n10318), .S0(n5271), .Y(
        \D_cache/n1105 ) );
  MX2XL U10310 ( .A(\D_cache/cache[2][86] ), .B(n10318), .S0(n5229), .Y(
        \D_cache/n1106 ) );
  MX2XL U10311 ( .A(\D_cache/cache[1][86] ), .B(n10318), .S0(n5201), .Y(
        \D_cache/n1107 ) );
  MX2XL U10312 ( .A(\D_cache/cache[0][86] ), .B(n10318), .S0(n5161), .Y(
        \D_cache/n1108 ) );
  MX2XL U10313 ( .A(\D_cache/cache[6][85] ), .B(n10525), .S0(n5370), .Y(
        \D_cache/n1110 ) );
  MX2XL U10314 ( .A(\D_cache/cache[5][85] ), .B(n10525), .S0(n5346), .Y(
        \D_cache/n1111 ) );
  MX2XL U10315 ( .A(\D_cache/cache[4][85] ), .B(n10525), .S0(n5319), .Y(
        \D_cache/n1112 ) );
  MX2XL U10316 ( .A(\D_cache/cache[3][85] ), .B(n10525), .S0(n5274), .Y(
        \D_cache/n1113 ) );
  MX2XL U10317 ( .A(\D_cache/cache[2][85] ), .B(n10525), .S0(n5232), .Y(
        \D_cache/n1114 ) );
  MX2XL U10318 ( .A(\D_cache/cache[1][85] ), .B(n10525), .S0(n5204), .Y(
        \D_cache/n1115 ) );
  MX2XL U10319 ( .A(\D_cache/cache[0][85] ), .B(n10525), .S0(n5167), .Y(
        \D_cache/n1116 ) );
  MX2XL U10320 ( .A(\D_cache/cache[6][84] ), .B(n4513), .S0(n5364), .Y(
        \D_cache/n1118 ) );
  MX2XL U10321 ( .A(\D_cache/cache[5][84] ), .B(n4513), .S0(n5340), .Y(
        \D_cache/n1119 ) );
  MX2XL U10322 ( .A(\D_cache/cache[4][84] ), .B(n4513), .S0(n5313), .Y(
        \D_cache/n1120 ) );
  MX2XL U10323 ( .A(\D_cache/cache[3][84] ), .B(n4513), .S0(n5268), .Y(
        \D_cache/n1121 ) );
  MX2XL U10324 ( .A(\D_cache/cache[2][84] ), .B(n4513), .S0(n5228), .Y(
        \D_cache/n1122 ) );
  MX2XL U10325 ( .A(\D_cache/cache[1][84] ), .B(n4513), .S0(n5198), .Y(
        \D_cache/n1123 ) );
  MX2XL U10326 ( .A(\D_cache/cache[0][84] ), .B(n4513), .S0(n5159), .Y(
        \D_cache/n1124 ) );
  MX2XL U10327 ( .A(\D_cache/cache[6][82] ), .B(n10645), .S0(n5370), .Y(
        \D_cache/n1134 ) );
  MX2XL U10328 ( .A(\D_cache/cache[5][82] ), .B(n10645), .S0(n5346), .Y(
        \D_cache/n1135 ) );
  MX2XL U10329 ( .A(\D_cache/cache[4][82] ), .B(n10645), .S0(n5319), .Y(
        \D_cache/n1136 ) );
  MX2XL U10330 ( .A(\D_cache/cache[3][82] ), .B(n10645), .S0(n5269), .Y(
        \D_cache/n1137 ) );
  MX2XL U10331 ( .A(\D_cache/cache[2][82] ), .B(n10645), .S0(n5232), .Y(
        \D_cache/n1138 ) );
  MX2XL U10332 ( .A(\D_cache/cache[1][82] ), .B(n10645), .S0(n5202), .Y(
        \D_cache/n1139 ) );
  MX2XL U10333 ( .A(\D_cache/cache[0][82] ), .B(n10645), .S0(n5162), .Y(
        \D_cache/n1140 ) );
  MX2XL U10334 ( .A(\D_cache/cache[6][81] ), .B(n10630), .S0(n5371), .Y(
        \D_cache/n1142 ) );
  MX2XL U10335 ( .A(\D_cache/cache[5][81] ), .B(n10630), .S0(n5347), .Y(
        \D_cache/n1143 ) );
  MX2XL U10336 ( .A(\D_cache/cache[4][81] ), .B(n10630), .S0(n5320), .Y(
        \D_cache/n1144 ) );
  MX2XL U10337 ( .A(\D_cache/cache[3][81] ), .B(n10630), .S0(n5274), .Y(
        \D_cache/n1145 ) );
  MX2XL U10338 ( .A(\D_cache/cache[2][81] ), .B(n10630), .S0(n5233), .Y(
        \D_cache/n1146 ) );
  MX2XL U10339 ( .A(\D_cache/cache[1][81] ), .B(n10630), .S0(n5205), .Y(
        \D_cache/n1147 ) );
  MX2XL U10340 ( .A(\D_cache/cache[0][81] ), .B(n10630), .S0(n5164), .Y(
        \D_cache/n1148 ) );
  MX2XL U10341 ( .A(\D_cache/cache[6][80] ), .B(n4514), .S0(n5365), .Y(
        \D_cache/n1150 ) );
  MX2XL U10342 ( .A(\D_cache/cache[5][80] ), .B(n4514), .S0(n5341), .Y(
        \D_cache/n1151 ) );
  MX2XL U10343 ( .A(\D_cache/cache[4][80] ), .B(n4514), .S0(n5314), .Y(
        \D_cache/n1152 ) );
  MX2XL U10344 ( .A(\D_cache/cache[3][80] ), .B(n4514), .S0(n5269), .Y(
        \D_cache/n1153 ) );
  MX2XL U10345 ( .A(\D_cache/cache[2][80] ), .B(n4514), .S0(n5231), .Y(
        \D_cache/n1154 ) );
  MX2XL U10346 ( .A(\D_cache/cache[1][80] ), .B(n4514), .S0(n5199), .Y(
        \D_cache/n1155 ) );
  MX2XL U10347 ( .A(\D_cache/cache[0][80] ), .B(n4514), .S0(n5160), .Y(
        \D_cache/n1156 ) );
  MX2XL U10348 ( .A(\D_cache/cache[6][79] ), .B(n4515), .S0(n5365), .Y(
        \D_cache/n1158 ) );
  MX2XL U10349 ( .A(\D_cache/cache[5][79] ), .B(n4515), .S0(n5341), .Y(
        \D_cache/n1159 ) );
  MX2XL U10350 ( .A(\D_cache/cache[4][79] ), .B(n4515), .S0(n5314), .Y(
        \D_cache/n1160 ) );
  MX2XL U10351 ( .A(\D_cache/cache[3][79] ), .B(n4515), .S0(n5269), .Y(
        \D_cache/n1161 ) );
  MX2XL U10352 ( .A(\D_cache/cache[2][79] ), .B(n4515), .S0(n5232), .Y(
        \D_cache/n1162 ) );
  MX2XL U10353 ( .A(\D_cache/cache[1][79] ), .B(n4515), .S0(n5199), .Y(
        \D_cache/n1163 ) );
  MX2XL U10354 ( .A(\D_cache/cache[0][79] ), .B(n4515), .S0(n5160), .Y(
        \D_cache/n1164 ) );
  MX2XL U10355 ( .A(\D_cache/cache[6][78] ), .B(n4525), .S0(n5366), .Y(
        \D_cache/n1166 ) );
  MX2XL U10356 ( .A(\D_cache/cache[5][78] ), .B(n4525), .S0(n5342), .Y(
        \D_cache/n1167 ) );
  MX2XL U10357 ( .A(\D_cache/cache[4][78] ), .B(n4525), .S0(n5315), .Y(
        \D_cache/n1168 ) );
  MX2XL U10358 ( .A(\D_cache/cache[3][78] ), .B(n4525), .S0(n5270), .Y(
        \D_cache/n1169 ) );
  MX2XL U10359 ( .A(\D_cache/cache[2][78] ), .B(n4525), .S0(n5228), .Y(
        \D_cache/n1170 ) );
  MX2XL U10360 ( .A(\D_cache/cache[1][78] ), .B(n4525), .S0(n5200), .Y(
        \D_cache/n1171 ) );
  MX2XL U10361 ( .A(\D_cache/cache[0][78] ), .B(n4525), .S0(n3564), .Y(
        \D_cache/n1172 ) );
  MX2XL U10362 ( .A(\D_cache/cache[6][76] ), .B(n4516), .S0(n5365), .Y(
        \D_cache/n1182 ) );
  MX2XL U10363 ( .A(\D_cache/cache[5][76] ), .B(n4516), .S0(n5341), .Y(
        \D_cache/n1183 ) );
  MX2XL U10364 ( .A(\D_cache/cache[4][76] ), .B(n4516), .S0(n5314), .Y(
        \D_cache/n1184 ) );
  MX2XL U10365 ( .A(\D_cache/cache[3][76] ), .B(n4516), .S0(n5269), .Y(
        \D_cache/n1185 ) );
  MX2XL U10366 ( .A(\D_cache/cache[2][76] ), .B(n4516), .S0(n5230), .Y(
        \D_cache/n1186 ) );
  MX2XL U10367 ( .A(\D_cache/cache[1][76] ), .B(n4516), .S0(n5199), .Y(
        \D_cache/n1187 ) );
  MX2XL U10368 ( .A(\D_cache/cache[0][76] ), .B(n4516), .S0(n5160), .Y(
        \D_cache/n1188 ) );
  MX2XL U10369 ( .A(\D_cache/cache[6][73] ), .B(n10617), .S0(n5371), .Y(
        \D_cache/n1206 ) );
  MX2XL U10370 ( .A(\D_cache/cache[5][73] ), .B(n10617), .S0(n5347), .Y(
        \D_cache/n1207 ) );
  MX2XL U10371 ( .A(\D_cache/cache[4][73] ), .B(n10617), .S0(n5320), .Y(
        \D_cache/n1208 ) );
  MX2XL U10372 ( .A(\D_cache/cache[3][73] ), .B(n10617), .S0(n5274), .Y(
        \D_cache/n1209 ) );
  MX2XL U10373 ( .A(\D_cache/cache[2][73] ), .B(n10617), .S0(n5233), .Y(
        \D_cache/n1210 ) );
  MX2XL U10374 ( .A(\D_cache/cache[1][73] ), .B(n10617), .S0(n5205), .Y(
        \D_cache/n1211 ) );
  MX2XL U10375 ( .A(\D_cache/cache[0][73] ), .B(n10617), .S0(n5164), .Y(
        \D_cache/n1212 ) );
  MX2XL U10376 ( .A(\D_cache/cache[6][72] ), .B(n10658), .S0(n5368), .Y(
        \D_cache/n1214 ) );
  MX2XL U10377 ( .A(\D_cache/cache[5][72] ), .B(n10658), .S0(n5344), .Y(
        \D_cache/n1215 ) );
  MX2XL U10378 ( .A(\D_cache/cache[4][72] ), .B(n10658), .S0(n5317), .Y(
        \D_cache/n1216 ) );
  MX2XL U10379 ( .A(\D_cache/cache[3][72] ), .B(n10658), .S0(n5272), .Y(
        \D_cache/n1217 ) );
  MX2XL U10380 ( .A(\D_cache/cache[2][72] ), .B(n10658), .S0(n5230), .Y(
        \D_cache/n1218 ) );
  MX2XL U10381 ( .A(\D_cache/cache[1][72] ), .B(n10658), .S0(n5202), .Y(
        \D_cache/n1219 ) );
  MX2XL U10382 ( .A(\D_cache/cache[0][72] ), .B(n10658), .S0(n5162), .Y(
        \D_cache/n1220 ) );
  MX2XL U10383 ( .A(\D_cache/cache[6][71] ), .B(n10685), .S0(n5367), .Y(
        \D_cache/n1222 ) );
  MX2XL U10384 ( .A(\D_cache/cache[5][71] ), .B(n10685), .S0(n5343), .Y(
        \D_cache/n1223 ) );
  MX2XL U10385 ( .A(\D_cache/cache[4][71] ), .B(n10685), .S0(n5316), .Y(
        \D_cache/n1224 ) );
  MX2XL U10386 ( .A(\D_cache/cache[3][71] ), .B(n10685), .S0(n5271), .Y(
        \D_cache/n1225 ) );
  MX2XL U10387 ( .A(\D_cache/cache[2][71] ), .B(n10685), .S0(n5229), .Y(
        \D_cache/n1226 ) );
  MX2XL U10388 ( .A(\D_cache/cache[1][71] ), .B(n10685), .S0(n5203), .Y(
        \D_cache/n1227 ) );
  MX2XL U10389 ( .A(\D_cache/cache[0][71] ), .B(n10685), .S0(n5163), .Y(
        \D_cache/n1228 ) );
  MX2XL U10390 ( .A(\D_cache/cache[6][70] ), .B(n4526), .S0(n5366), .Y(
        \D_cache/n1230 ) );
  MX2XL U10391 ( .A(\D_cache/cache[5][70] ), .B(n4526), .S0(n5342), .Y(
        \D_cache/n1231 ) );
  MX2XL U10392 ( .A(\D_cache/cache[4][70] ), .B(n4526), .S0(n5315), .Y(
        \D_cache/n1232 ) );
  MX2XL U10393 ( .A(\D_cache/cache[3][70] ), .B(n4526), .S0(n5270), .Y(
        \D_cache/n1233 ) );
  MX2XL U10394 ( .A(\D_cache/cache[2][70] ), .B(n4526), .S0(n5234), .Y(
        \D_cache/n1234 ) );
  MX2XL U10395 ( .A(\D_cache/cache[1][70] ), .B(n4526), .S0(n5200), .Y(
        \D_cache/n1235 ) );
  MX2XL U10396 ( .A(\D_cache/cache[0][70] ), .B(n4526), .S0(n5164), .Y(
        \D_cache/n1236 ) );
  MX2XL U10397 ( .A(\D_cache/cache[6][66] ), .B(n10197), .S0(n5367), .Y(
        \D_cache/n1262 ) );
  MX2XL U10398 ( .A(\D_cache/cache[5][66] ), .B(n10197), .S0(n5343), .Y(
        \D_cache/n1263 ) );
  MX2XL U10399 ( .A(\D_cache/cache[4][66] ), .B(n10197), .S0(n5316), .Y(
        \D_cache/n1264 ) );
  MX2XL U10400 ( .A(\D_cache/cache[3][66] ), .B(n10197), .S0(n5271), .Y(
        \D_cache/n1265 ) );
  MX2XL U10401 ( .A(\D_cache/cache[2][66] ), .B(n10197), .S0(n5229), .Y(
        \D_cache/n1266 ) );
  MX2XL U10402 ( .A(\D_cache/cache[1][66] ), .B(n10197), .S0(n5201), .Y(
        \D_cache/n1267 ) );
  MX2XL U10403 ( .A(\D_cache/cache[0][66] ), .B(n10197), .S0(n5161), .Y(
        \D_cache/n1268 ) );
  MX2XL U10404 ( .A(\D_cache/cache[6][65] ), .B(n10672), .S0(n5368), .Y(
        \D_cache/n1270 ) );
  MX2XL U10405 ( .A(\D_cache/cache[5][65] ), .B(n10672), .S0(n5344), .Y(
        \D_cache/n1271 ) );
  MX2XL U10406 ( .A(\D_cache/cache[4][65] ), .B(n10672), .S0(n5317), .Y(
        \D_cache/n1272 ) );
  MX2XL U10407 ( .A(\D_cache/cache[3][65] ), .B(n10672), .S0(n5272), .Y(
        \D_cache/n1273 ) );
  MX2XL U10408 ( .A(\D_cache/cache[2][65] ), .B(n10672), .S0(n5230), .Y(
        \D_cache/n1274 ) );
  MX2XL U10409 ( .A(\D_cache/cache[1][65] ), .B(n10672), .S0(n5202), .Y(
        \D_cache/n1275 ) );
  MX2XL U10410 ( .A(\D_cache/cache[0][65] ), .B(n10672), .S0(n5162), .Y(
        \D_cache/n1276 ) );
  MX2XL U10411 ( .A(\D_cache/cache[6][83] ), .B(n10977), .S0(n5372), .Y(
        \D_cache/n1126 ) );
  MX2XL U10412 ( .A(\D_cache/cache[5][83] ), .B(n10977), .S0(n5349), .Y(
        \D_cache/n1127 ) );
  MX2XL U10413 ( .A(\D_cache/cache[4][83] ), .B(n10977), .S0(n5321), .Y(
        \D_cache/n1128 ) );
  MX2XL U10414 ( .A(\D_cache/cache[3][83] ), .B(n10977), .S0(n5276), .Y(
        \D_cache/n1129 ) );
  MX2XL U10415 ( .A(\D_cache/cache[2][83] ), .B(n10977), .S0(n5232), .Y(
        \D_cache/n1130 ) );
  MX2XL U10416 ( .A(\D_cache/cache[1][83] ), .B(n10977), .S0(n5207), .Y(
        \D_cache/n1131 ) );
  MX2XL U10417 ( .A(\D_cache/cache[0][83] ), .B(n10977), .S0(n5165), .Y(
        \D_cache/n1132 ) );
  MX2XL U10418 ( .A(\D_cache/cache[6][77] ), .B(n10810), .S0(n3574), .Y(
        \D_cache/n1174 ) );
  MX2XL U10419 ( .A(\D_cache/cache[5][77] ), .B(n10810), .S0(n5350), .Y(
        \D_cache/n1175 ) );
  MX2XL U10420 ( .A(\D_cache/cache[4][77] ), .B(n10810), .S0(n5323), .Y(
        \D_cache/n1176 ) );
  MX2XL U10421 ( .A(\D_cache/cache[3][77] ), .B(n10810), .S0(n5276), .Y(
        \D_cache/n1177 ) );
  MX2XL U10422 ( .A(\D_cache/cache[2][77] ), .B(n10810), .S0(n5236), .Y(
        \D_cache/n1178 ) );
  MX2XL U10423 ( .A(\D_cache/cache[1][77] ), .B(n10810), .S0(n5208), .Y(
        \D_cache/n1179 ) );
  MX2XL U10424 ( .A(\D_cache/cache[0][77] ), .B(n10810), .S0(n5168), .Y(
        \D_cache/n1180 ) );
  MX2XL U10425 ( .A(\D_cache/cache[6][75] ), .B(n4500), .S0(n3574), .Y(
        \D_cache/n1190 ) );
  MX2XL U10426 ( .A(\D_cache/cache[5][75] ), .B(n4500), .S0(n5350), .Y(
        \D_cache/n1191 ) );
  MX2XL U10427 ( .A(\D_cache/cache[4][75] ), .B(n4500), .S0(n5323), .Y(
        \D_cache/n1192 ) );
  MX2XL U10428 ( .A(\D_cache/cache[3][75] ), .B(n4500), .S0(n5276), .Y(
        \D_cache/n1193 ) );
  MX2XL U10429 ( .A(\D_cache/cache[2][75] ), .B(n4500), .S0(n5236), .Y(
        \D_cache/n1194 ) );
  MX2XL U10430 ( .A(\D_cache/cache[1][75] ), .B(n4500), .S0(n5208), .Y(
        \D_cache/n1195 ) );
  MX2XL U10431 ( .A(\D_cache/cache[0][75] ), .B(n4500), .S0(n5168), .Y(
        \D_cache/n1196 ) );
  MX2XL U10432 ( .A(\D_cache/cache[6][74] ), .B(n4501), .S0(n5372), .Y(
        \D_cache/n1198 ) );
  MX2XL U10433 ( .A(\D_cache/cache[5][74] ), .B(n4501), .S0(n5349), .Y(
        \D_cache/n1199 ) );
  MX2XL U10434 ( .A(\D_cache/cache[4][74] ), .B(n4501), .S0(n3763), .Y(
        \D_cache/n1200 ) );
  MX2XL U10435 ( .A(\D_cache/cache[3][74] ), .B(n4501), .S0(n5275), .Y(
        \D_cache/n1201 ) );
  MX2XL U10436 ( .A(\D_cache/cache[2][74] ), .B(n4501), .S0(n5235), .Y(
        \D_cache/n1202 ) );
  MX2XL U10437 ( .A(\D_cache/cache[1][74] ), .B(n4501), .S0(n5207), .Y(
        \D_cache/n1203 ) );
  MX2XL U10438 ( .A(\D_cache/cache[0][74] ), .B(n4501), .S0(n5167), .Y(
        \D_cache/n1204 ) );
  MX2XL U10439 ( .A(\D_cache/cache[6][69] ), .B(n10902), .S0(n3574), .Y(
        \D_cache/n1238 ) );
  MX2XL U10440 ( .A(\D_cache/cache[5][69] ), .B(n10902), .S0(n5350), .Y(
        \D_cache/n1239 ) );
  MX2XL U10441 ( .A(\D_cache/cache[4][69] ), .B(n10902), .S0(n5323), .Y(
        \D_cache/n1240 ) );
  MX2XL U10442 ( .A(\D_cache/cache[3][69] ), .B(n10902), .S0(n5276), .Y(
        \D_cache/n1241 ) );
  MX2XL U10443 ( .A(\D_cache/cache[2][69] ), .B(n10902), .S0(n5236), .Y(
        \D_cache/n1242 ) );
  MX2XL U10444 ( .A(\D_cache/cache[1][69] ), .B(n10902), .S0(n5208), .Y(
        \D_cache/n1243 ) );
  MX2XL U10445 ( .A(\D_cache/cache[0][69] ), .B(n10902), .S0(n5168), .Y(
        \D_cache/n1244 ) );
  MX2XL U10446 ( .A(\D_cache/cache[3][68] ), .B(n10757), .S0(n5275), .Y(
        \D_cache/n1249 ) );
  MX2XL U10447 ( .A(\D_cache/cache[2][68] ), .B(n10757), .S0(n5235), .Y(
        \D_cache/n1250 ) );
  MX2XL U10448 ( .A(\D_cache/cache[1][68] ), .B(n10757), .S0(n5207), .Y(
        \D_cache/n1251 ) );
  MX2XL U10449 ( .A(\D_cache/cache[6][67] ), .B(n4502), .S0(n5372), .Y(
        \D_cache/n1254 ) );
  MX2XL U10450 ( .A(\D_cache/cache[5][67] ), .B(n4502), .S0(n5349), .Y(
        \D_cache/n1255 ) );
  MX2XL U10451 ( .A(\D_cache/cache[4][67] ), .B(n4502), .S0(n3763), .Y(
        \D_cache/n1256 ) );
  MX2XL U10452 ( .A(\D_cache/cache[3][67] ), .B(n4502), .S0(n5275), .Y(
        \D_cache/n1257 ) );
  MX2XL U10453 ( .A(\D_cache/cache[2][67] ), .B(n4502), .S0(n5235), .Y(
        \D_cache/n1258 ) );
  MX2XL U10454 ( .A(\D_cache/cache[1][67] ), .B(n4502), .S0(n5207), .Y(
        \D_cache/n1259 ) );
  MX2XL U10455 ( .A(\D_cache/cache[0][67] ), .B(n4502), .S0(n5167), .Y(
        \D_cache/n1260 ) );
  MX2XL U10456 ( .A(\D_cache/cache[6][64] ), .B(n10749), .S0(n5368), .Y(
        \D_cache/n1278 ) );
  MX2XL U10457 ( .A(\D_cache/cache[5][64] ), .B(n10749), .S0(n5344), .Y(
        \D_cache/n1279 ) );
  MX2XL U10458 ( .A(\D_cache/cache[4][64] ), .B(n10749), .S0(n5317), .Y(
        \D_cache/n1280 ) );
  MX2XL U10459 ( .A(\D_cache/cache[3][64] ), .B(n10749), .S0(n5272), .Y(
        \D_cache/n1281 ) );
  MX2XL U10460 ( .A(\D_cache/cache[2][64] ), .B(n10749), .S0(n5230), .Y(
        \D_cache/n1282 ) );
  MX2XL U10461 ( .A(\D_cache/cache[1][64] ), .B(n10749), .S0(n5202), .Y(
        \D_cache/n1283 ) );
  MX2XL U10462 ( .A(\D_cache/cache[0][64] ), .B(n10749), .S0(n5167), .Y(
        \D_cache/n1284 ) );
  MX2XL U10463 ( .A(\D_cache/cache[6][109] ), .B(n10807), .S0(n3574), .Y(
        \D_cache/n918 ) );
  MX2XL U10464 ( .A(\D_cache/cache[5][109] ), .B(n10807), .S0(n5350), .Y(
        \D_cache/n919 ) );
  MX2XL U10465 ( .A(\D_cache/cache[4][109] ), .B(n10807), .S0(n5323), .Y(
        \D_cache/n920 ) );
  MX2XL U10466 ( .A(\D_cache/cache[3][109] ), .B(n10807), .S0(n5276), .Y(
        \D_cache/n921 ) );
  MX2XL U10467 ( .A(\D_cache/cache[2][109] ), .B(n10807), .S0(n5236), .Y(
        \D_cache/n922 ) );
  MX2XL U10468 ( .A(\D_cache/cache[1][109] ), .B(n10807), .S0(n5208), .Y(
        \D_cache/n923 ) );
  MX2XL U10469 ( .A(\D_cache/cache[0][109] ), .B(n10807), .S0(n5168), .Y(
        \D_cache/n924 ) );
  MX2XL U10470 ( .A(\D_cache/cache[6][107] ), .B(n4497), .S0(n5364), .Y(
        \D_cache/n934 ) );
  MX2XL U10471 ( .A(\D_cache/cache[5][107] ), .B(n4497), .S0(n5340), .Y(
        \D_cache/n935 ) );
  MX2XL U10472 ( .A(\D_cache/cache[4][107] ), .B(n4497), .S0(n5313), .Y(
        \D_cache/n936 ) );
  MX2XL U10473 ( .A(\D_cache/cache[3][107] ), .B(n4497), .S0(n5268), .Y(
        \D_cache/n937 ) );
  MX2XL U10474 ( .A(\D_cache/cache[2][107] ), .B(n4497), .S0(n5228), .Y(
        \D_cache/n938 ) );
  MX2XL U10475 ( .A(\D_cache/cache[1][107] ), .B(n4497), .S0(n5198), .Y(
        \D_cache/n939 ) );
  MX2XL U10476 ( .A(\D_cache/cache[0][107] ), .B(n4497), .S0(n5159), .Y(
        \D_cache/n940 ) );
  MX2XL U10477 ( .A(\D_cache/cache[6][106] ), .B(n4498), .S0(n5372), .Y(
        \D_cache/n942 ) );
  MX2XL U10478 ( .A(\D_cache/cache[5][106] ), .B(n4498), .S0(n5349), .Y(
        \D_cache/n943 ) );
  MX2XL U10479 ( .A(\D_cache/cache[4][106] ), .B(n4498), .S0(n3763), .Y(
        \D_cache/n944 ) );
  MX2XL U10480 ( .A(\D_cache/cache[3][106] ), .B(n4498), .S0(n5275), .Y(
        \D_cache/n945 ) );
  MX2XL U10481 ( .A(\D_cache/cache[2][106] ), .B(n4498), .S0(n5235), .Y(
        \D_cache/n946 ) );
  MX2XL U10482 ( .A(\D_cache/cache[1][106] ), .B(n4498), .S0(n5207), .Y(
        \D_cache/n947 ) );
  MX2XL U10483 ( .A(\D_cache/cache[0][106] ), .B(n4498), .S0(n5167), .Y(
        \D_cache/n948 ) );
  MX2XL U10484 ( .A(\D_cache/cache[6][101] ), .B(n10899), .S0(n3574), .Y(
        \D_cache/n982 ) );
  MX2XL U10485 ( .A(\D_cache/cache[5][101] ), .B(n10899), .S0(n5350), .Y(
        \D_cache/n983 ) );
  MX2XL U10486 ( .A(\D_cache/cache[4][101] ), .B(n10899), .S0(n5323), .Y(
        \D_cache/n984 ) );
  MX2XL U10487 ( .A(\D_cache/cache[3][101] ), .B(n10899), .S0(n5276), .Y(
        \D_cache/n985 ) );
  MX2XL U10488 ( .A(\D_cache/cache[2][101] ), .B(n10899), .S0(n5236), .Y(
        \D_cache/n986 ) );
  MX2XL U10489 ( .A(\D_cache/cache[1][101] ), .B(n10899), .S0(n5208), .Y(
        \D_cache/n987 ) );
  MX2XL U10490 ( .A(\D_cache/cache[0][101] ), .B(n10899), .S0(n5168), .Y(
        \D_cache/n988 ) );
  MX2XL U10491 ( .A(\D_cache/cache[6][100] ), .B(n10754), .S0(n5372), .Y(
        \D_cache/n990 ) );
  MX2XL U10492 ( .A(\D_cache/cache[5][100] ), .B(n10754), .S0(n5349), .Y(
        \D_cache/n991 ) );
  MX2XL U10493 ( .A(\D_cache/cache[4][100] ), .B(n10754), .S0(n3763), .Y(
        \D_cache/n992 ) );
  MX2XL U10494 ( .A(\D_cache/cache[3][100] ), .B(n10754), .S0(n5275), .Y(
        \D_cache/n993 ) );
  MX2XL U10495 ( .A(\D_cache/cache[2][100] ), .B(n10754), .S0(n5235), .Y(
        \D_cache/n994 ) );
  MX2XL U10496 ( .A(\D_cache/cache[1][100] ), .B(n10754), .S0(n5207), .Y(
        \D_cache/n995 ) );
  MX2XL U10497 ( .A(\D_cache/cache[0][100] ), .B(n10754), .S0(n5167), .Y(
        \D_cache/n996 ) );
  MX2XL U10498 ( .A(\D_cache/cache[6][99] ), .B(n4499), .S0(n5372), .Y(
        \D_cache/n998 ) );
  MX2XL U10499 ( .A(\D_cache/cache[5][99] ), .B(n4499), .S0(n5349), .Y(
        \D_cache/n999 ) );
  MX2XL U10500 ( .A(\D_cache/cache[4][99] ), .B(n4499), .S0(n3763), .Y(
        \D_cache/n1000 ) );
  MX2XL U10501 ( .A(\D_cache/cache[3][99] ), .B(n4499), .S0(n5275), .Y(
        \D_cache/n1001 ) );
  MX2XL U10502 ( .A(\D_cache/cache[2][99] ), .B(n4499), .S0(n5235), .Y(
        \D_cache/n1002 ) );
  MX2XL U10503 ( .A(\D_cache/cache[1][99] ), .B(n4499), .S0(n5207), .Y(
        \D_cache/n1003 ) );
  MX2XL U10504 ( .A(\D_cache/cache[0][99] ), .B(n4499), .S0(n5167), .Y(
        \D_cache/n1004 ) );
  MX2XL U10505 ( .A(\D_cache/cache[6][96] ), .B(n10746), .S0(n5369), .Y(
        \D_cache/n1022 ) );
  MX2XL U10506 ( .A(\D_cache/cache[5][96] ), .B(n10746), .S0(n3575), .Y(
        \D_cache/n1023 ) );
  MX2XL U10507 ( .A(\D_cache/cache[4][96] ), .B(n10746), .S0(n5318), .Y(
        \D_cache/n1024 ) );
  MX2XL U10508 ( .A(\D_cache/cache[3][96] ), .B(n10746), .S0(n5273), .Y(
        \D_cache/n1025 ) );
  MX2XL U10509 ( .A(\D_cache/cache[2][96] ), .B(n10746), .S0(n5231), .Y(
        \D_cache/n1026 ) );
  MX2XL U10510 ( .A(\D_cache/cache[1][96] ), .B(n10746), .S0(n5202), .Y(
        \D_cache/n1027 ) );
  MX2XL U10511 ( .A(\D_cache/cache[0][96] ), .B(n10746), .S0(n5162), .Y(
        \D_cache/n1028 ) );
  MX2XL U10512 ( .A(\D_cache/cache[5][45] ), .B(n4538), .S0(n5350), .Y(
        \D_cache/n1431 ) );
  MX2XL U10513 ( .A(\D_cache/cache[4][45] ), .B(n4538), .S0(n5323), .Y(
        \D_cache/n1432 ) );
  MX2XL U10514 ( .A(\D_cache/cache[3][45] ), .B(n4538), .S0(n5276), .Y(
        \D_cache/n1433 ) );
  MX2XL U10515 ( .A(\D_cache/cache[2][45] ), .B(n4538), .S0(n5236), .Y(
        \D_cache/n1434 ) );
  MX2XL U10516 ( .A(\D_cache/cache[1][45] ), .B(n4538), .S0(n5208), .Y(
        \D_cache/n1435 ) );
  MX2XL U10517 ( .A(\D_cache/cache[0][45] ), .B(n4538), .S0(n5168), .Y(
        \D_cache/n1436 ) );
  MX2XL U10518 ( .A(\D_cache/cache[6][43] ), .B(n10789), .S0(n5373), .Y(
        \D_cache/n1446 ) );
  MX2XL U10519 ( .A(\D_cache/cache[5][43] ), .B(n10789), .S0(n5348), .Y(
        \D_cache/n1447 ) );
  MX2XL U10520 ( .A(\D_cache/cache[4][43] ), .B(n10789), .S0(n5322), .Y(
        \D_cache/n1448 ) );
  MX2XL U10521 ( .A(\D_cache/cache[3][43] ), .B(n10789), .S0(n5268), .Y(
        \D_cache/n1449 ) );
  MX2XL U10522 ( .A(\D_cache/cache[2][43] ), .B(n10789), .S0(n5234), .Y(
        \D_cache/n1450 ) );
  MX2XL U10523 ( .A(\D_cache/cache[1][43] ), .B(n10789), .S0(n5206), .Y(
        \D_cache/n1451 ) );
  MX2XL U10524 ( .A(\D_cache/cache[0][43] ), .B(n10789), .S0(n5166), .Y(
        \D_cache/n1452 ) );
  MX2XL U10525 ( .A(\D_cache/cache[6][42] ), .B(n4539), .S0(n3574), .Y(
        \D_cache/n1454 ) );
  MX2XL U10526 ( .A(\D_cache/cache[5][42] ), .B(n4539), .S0(n5349), .Y(
        \D_cache/n1455 ) );
  MX2XL U10527 ( .A(\D_cache/cache[4][42] ), .B(n4539), .S0(n3763), .Y(
        \D_cache/n1456 ) );
  MX2XL U10528 ( .A(\D_cache/cache[3][42] ), .B(n4539), .S0(n5275), .Y(
        \D_cache/n1457 ) );
  MX2XL U10529 ( .A(\D_cache/cache[2][42] ), .B(n4539), .S0(n5235), .Y(
        \D_cache/n1458 ) );
  MX2XL U10530 ( .A(\D_cache/cache[1][42] ), .B(n4539), .S0(n5207), .Y(
        \D_cache/n1459 ) );
  MX2XL U10531 ( .A(\D_cache/cache[0][42] ), .B(n4539), .S0(n5167), .Y(
        \D_cache/n1460 ) );
  MX2XL U10532 ( .A(\D_cache/cache[6][37] ), .B(n10896), .S0(n3574), .Y(
        \D_cache/n1494 ) );
  MX2XL U10533 ( .A(\D_cache/cache[5][37] ), .B(n10896), .S0(n5350), .Y(
        \D_cache/n1495 ) );
  MX2XL U10534 ( .A(\D_cache/cache[4][37] ), .B(n10896), .S0(n5323), .Y(
        \D_cache/n1496 ) );
  MX2XL U10535 ( .A(\D_cache/cache[3][37] ), .B(n10896), .S0(n5276), .Y(
        \D_cache/n1497 ) );
  MX2XL U10536 ( .A(\D_cache/cache[2][37] ), .B(n10896), .S0(n5236), .Y(
        \D_cache/n1498 ) );
  MX2XL U10537 ( .A(\D_cache/cache[1][37] ), .B(n10896), .S0(n5208), .Y(
        \D_cache/n1499 ) );
  MX2XL U10538 ( .A(\D_cache/cache[0][37] ), .B(n10896), .S0(n5168), .Y(
        \D_cache/n1500 ) );
  MX2XL U10539 ( .A(\D_cache/cache[6][36] ), .B(n4540), .S0(n5368), .Y(
        \D_cache/n1502 ) );
  MX2XL U10540 ( .A(\D_cache/cache[5][36] ), .B(n4540), .S0(n5344), .Y(
        \D_cache/n1503 ) );
  MX2XL U10541 ( .A(\D_cache/cache[4][36] ), .B(n4540), .S0(n5317), .Y(
        \D_cache/n1504 ) );
  MX2XL U10542 ( .A(\D_cache/cache[3][36] ), .B(n4540), .S0(n5272), .Y(
        \D_cache/n1505 ) );
  MX2XL U10543 ( .A(\D_cache/cache[2][36] ), .B(n4540), .S0(n5230), .Y(
        \D_cache/n1506 ) );
  MX2XL U10544 ( .A(\D_cache/cache[1][36] ), .B(n4540), .S0(n5207), .Y(
        \D_cache/n1507 ) );
  MX2XL U10545 ( .A(\D_cache/cache[0][36] ), .B(n4540), .S0(n5167), .Y(
        \D_cache/n1508 ) );
  MX2XL U10546 ( .A(\D_cache/cache[6][35] ), .B(n10761), .S0(n3574), .Y(
        \D_cache/n1510 ) );
  MX2XL U10547 ( .A(\D_cache/cache[5][35] ), .B(n10761), .S0(n5349), .Y(
        \D_cache/n1511 ) );
  MX2XL U10548 ( .A(\D_cache/cache[4][35] ), .B(n10761), .S0(n3763), .Y(
        \D_cache/n1512 ) );
  MX2XL U10549 ( .A(\D_cache/cache[3][35] ), .B(n10761), .S0(n5275), .Y(
        \D_cache/n1513 ) );
  MX2XL U10550 ( .A(\D_cache/cache[2][35] ), .B(n10761), .S0(n5235), .Y(
        \D_cache/n1514 ) );
  MX2XL U10551 ( .A(\D_cache/cache[1][35] ), .B(n10761), .S0(n5207), .Y(
        \D_cache/n1515 ) );
  MX2XL U10552 ( .A(\D_cache/cache[0][35] ), .B(n10761), .S0(n5167), .Y(
        \D_cache/n1516 ) );
  MX2XL U10553 ( .A(\D_cache/cache[6][32] ), .B(n4541), .S0(n5369), .Y(
        \D_cache/n1534 ) );
  MX2XL U10554 ( .A(\D_cache/cache[5][32] ), .B(n4541), .S0(n3575), .Y(
        \D_cache/n1535 ) );
  MX2XL U10555 ( .A(\D_cache/cache[4][32] ), .B(n4541), .S0(n5318), .Y(
        \D_cache/n1536 ) );
  MX2XL U10556 ( .A(\D_cache/cache[3][32] ), .B(n4541), .S0(n5273), .Y(
        \D_cache/n1537 ) );
  MX2XL U10557 ( .A(\D_cache/cache[2][32] ), .B(n4541), .S0(n5231), .Y(
        \D_cache/n1538 ) );
  MX2XL U10558 ( .A(\D_cache/cache[1][32] ), .B(n4541), .S0(n5203), .Y(
        \D_cache/n1539 ) );
  MX2XL U10559 ( .A(\D_cache/cache[0][32] ), .B(n4541), .S0(n5162), .Y(
        \D_cache/n1540 ) );
  MX2XL U10560 ( .A(\D_cache/cache[6][31] ), .B(n10701), .S0(n5369), .Y(
        \D_cache/n1542 ) );
  MX2XL U10561 ( .A(\D_cache/cache[5][31] ), .B(n10701), .S0(n3575), .Y(
        \D_cache/n1543 ) );
  MX2XL U10562 ( .A(\D_cache/cache[4][31] ), .B(n10701), .S0(n5318), .Y(
        \D_cache/n1544 ) );
  MX2XL U10563 ( .A(\D_cache/cache[3][31] ), .B(n10701), .S0(n5273), .Y(
        \D_cache/n1545 ) );
  MX2XL U10564 ( .A(\D_cache/cache[2][31] ), .B(n10701), .S0(n5231), .Y(
        \D_cache/n1546 ) );
  MX2XL U10565 ( .A(\D_cache/cache[1][31] ), .B(n10701), .S0(n5203), .Y(
        \D_cache/n1547 ) );
  MX2XL U10566 ( .A(\D_cache/cache[0][31] ), .B(n10701), .S0(n5163), .Y(
        \D_cache/n1548 ) );
  MX2XL U10567 ( .A(\D_cache/cache[6][23] ), .B(n3014), .S0(n5369), .Y(
        \D_cache/n1606 ) );
  MX2XL U10568 ( .A(\D_cache/cache[5][23] ), .B(n3014), .S0(n3575), .Y(
        \D_cache/n1607 ) );
  MX2XL U10569 ( .A(\D_cache/cache[4][23] ), .B(n3014), .S0(n5318), .Y(
        \D_cache/n1608 ) );
  MX2XL U10570 ( .A(\D_cache/cache[3][23] ), .B(n3014), .S0(n5273), .Y(
        \D_cache/n1609 ) );
  MX2XL U10571 ( .A(\D_cache/cache[2][23] ), .B(n3014), .S0(n5231), .Y(
        \D_cache/n1610 ) );
  MX2XL U10572 ( .A(\D_cache/cache[1][23] ), .B(n3014), .S0(n5203), .Y(
        \D_cache/n1611 ) );
  MX2XL U10573 ( .A(\D_cache/cache[0][23] ), .B(n3014), .S0(n5163), .Y(
        \D_cache/n1612 ) );
  MX2XL U10574 ( .A(\D_cache/cache[6][13] ), .B(n147), .S0(n3574), .Y(
        \D_cache/n1686 ) );
  MX2XL U10575 ( .A(\D_cache/cache[5][13] ), .B(n147), .S0(n5350), .Y(
        \D_cache/n1687 ) );
  MX2XL U10576 ( .A(\D_cache/cache[4][13] ), .B(n147), .S0(n5323), .Y(
        \D_cache/n1688 ) );
  MX2XL U10577 ( .A(\D_cache/cache[3][13] ), .B(n147), .S0(n5276), .Y(
        \D_cache/n1689 ) );
  MX2XL U10578 ( .A(\D_cache/cache[2][13] ), .B(n147), .S0(n5236), .Y(
        \D_cache/n1690 ) );
  MX2XL U10579 ( .A(\D_cache/cache[1][13] ), .B(n147), .S0(n5208), .Y(
        \D_cache/n1691 ) );
  MX2XL U10580 ( .A(\D_cache/cache[0][13] ), .B(n147), .S0(n5168), .Y(
        \D_cache/n1692 ) );
  MX2XL U10581 ( .A(\D_cache/cache[6][11] ), .B(n4542), .S0(n3574), .Y(
        \D_cache/n1702 ) );
  MX2XL U10582 ( .A(\D_cache/cache[5][11] ), .B(n4542), .S0(n5349), .Y(
        \D_cache/n1703 ) );
  MX2XL U10583 ( .A(\D_cache/cache[4][11] ), .B(n4542), .S0(n3763), .Y(
        \D_cache/n1704 ) );
  MX2XL U10584 ( .A(\D_cache/cache[3][11] ), .B(n4542), .S0(n5275), .Y(
        \D_cache/n1705 ) );
  MX2XL U10585 ( .A(\D_cache/cache[2][11] ), .B(n4542), .S0(n5235), .Y(
        \D_cache/n1706 ) );
  MX2XL U10586 ( .A(\D_cache/cache[1][11] ), .B(n4542), .S0(n5207), .Y(
        \D_cache/n1707 ) );
  MX2XL U10587 ( .A(\D_cache/cache[0][11] ), .B(n4542), .S0(n5167), .Y(
        \D_cache/n1708 ) );
  MX2XL U10588 ( .A(\D_cache/cache[6][10] ), .B(n4543), .S0(n3574), .Y(
        \D_cache/n1710 ) );
  MX2XL U10589 ( .A(\D_cache/cache[5][10] ), .B(n4543), .S0(n5349), .Y(
        \D_cache/n1711 ) );
  MX2XL U10590 ( .A(\D_cache/cache[4][10] ), .B(n4543), .S0(n3763), .Y(
        \D_cache/n1712 ) );
  MX2XL U10591 ( .A(\D_cache/cache[3][10] ), .B(n4543), .S0(n5275), .Y(
        \D_cache/n1713 ) );
  MX2XL U10592 ( .A(\D_cache/cache[2][10] ), .B(n4543), .S0(n5235), .Y(
        \D_cache/n1714 ) );
  MX2XL U10593 ( .A(\D_cache/cache[1][10] ), .B(n4543), .S0(n5207), .Y(
        \D_cache/n1715 ) );
  MX2XL U10594 ( .A(\D_cache/cache[0][10] ), .B(n4543), .S0(n5167), .Y(
        \D_cache/n1716 ) );
  MX2XL U10595 ( .A(\D_cache/cache[6][5] ), .B(n4537), .S0(n3574), .Y(
        \D_cache/n1750 ) );
  MX2XL U10596 ( .A(\D_cache/cache[5][5] ), .B(n4537), .S0(n5350), .Y(
        \D_cache/n1751 ) );
  MX2XL U10597 ( .A(\D_cache/cache[4][5] ), .B(n4537), .S0(n5323), .Y(
        \D_cache/n1752 ) );
  MX2XL U10598 ( .A(\D_cache/cache[3][5] ), .B(n4537), .S0(n5276), .Y(
        \D_cache/n1753 ) );
  MX2XL U10599 ( .A(\D_cache/cache[2][5] ), .B(n4537), .S0(n5236), .Y(
        \D_cache/n1754 ) );
  MX2XL U10600 ( .A(\D_cache/cache[1][5] ), .B(n4537), .S0(n5208), .Y(
        \D_cache/n1755 ) );
  MX2XL U10601 ( .A(\D_cache/cache[0][5] ), .B(n4537), .S0(n5168), .Y(
        \D_cache/n1756 ) );
  MX2XL U10602 ( .A(\D_cache/cache[6][0] ), .B(n10740), .S0(n5369), .Y(
        \D_cache/n1789 ) );
  MX2XL U10603 ( .A(\D_cache/cache[5][0] ), .B(n10740), .S0(n3575), .Y(
        \D_cache/n1790 ) );
  MX2XL U10604 ( .A(\D_cache/cache[4][0] ), .B(n10740), .S0(n5318), .Y(
        \D_cache/n1791 ) );
  MX2XL U10605 ( .A(\D_cache/cache[3][0] ), .B(n10740), .S0(n5273), .Y(
        \D_cache/n1792 ) );
  MX2XL U10606 ( .A(\D_cache/cache[2][0] ), .B(n10740), .S0(n5231), .Y(
        \D_cache/n1793 ) );
  MX2XL U10607 ( .A(\D_cache/cache[1][0] ), .B(n10740), .S0(n5203), .Y(
        \D_cache/n1794 ) );
  MX2XL U10608 ( .A(\D_cache/cache[0][0] ), .B(n10740), .S0(n5163), .Y(
        \D_cache/n1795 ) );
  OA22X1 U10609 ( .A0(\i_MIPS/Register/register[17][10] ), .A1(net118453), 
        .B0(\i_MIPS/Register/register[25][10] ), .B1(net118473), .Y(n7517) );
  OA22X1 U10610 ( .A0(\i_MIPS/Register/register[17][19] ), .A1(net118451), 
        .B0(\i_MIPS/Register/register[25][19] ), .B1(net118475), .Y(n8323) );
  OA22X1 U10611 ( .A0(\i_MIPS/Register/register[17][13] ), .A1(net118451), 
        .B0(\i_MIPS/Register/register[25][13] ), .B1(net118475), .Y(n7980) );
  OA22X1 U10612 ( .A0(\i_MIPS/Register/register[17][5] ), .A1(net118455), .B0(
        \i_MIPS/Register/register[25][5] ), .B1(net118479), .Y(n9338) );
  OA22X1 U10613 ( .A0(\i_MIPS/Register/register[17][3] ), .A1(net118455), .B0(
        \i_MIPS/Register/register[25][3] ), .B1(net118479), .Y(n9157) );
  OA22X1 U10614 ( .A0(\i_MIPS/Register/register[17][0] ), .A1(net118453), .B0(
        \i_MIPS/Register/register[25][0] ), .B1(net118477), .Y(n8733) );
  OA22X1 U10615 ( .A0(\i_MIPS/Register/register[17][1] ), .A1(net118453), .B0(
        \i_MIPS/Register/register[25][1] ), .B1(net118477), .Y(n8996) );
  OA22X1 U10616 ( .A0(\i_MIPS/Register/register[17][16] ), .A1(net118453), 
        .B0(\i_MIPS/Register/register[25][16] ), .B1(net118477), .Y(n8809) );
  OA22X1 U10617 ( .A0(\i_MIPS/Register/register[17][23] ), .A1(net118453), 
        .B0(\i_MIPS/Register/register[25][23] ), .B1(net118479), .Y(n7091) );
  OA22X1 U10618 ( .A0(\i_MIPS/Register/register[17][29] ), .A1(net118453), 
        .B0(\i_MIPS/Register/register[25][29] ), .B1(net118479), .Y(n6995) );
  MX2XL U10619 ( .A(n3558), .B(n4937), .S0(n3601), .Y(\i_MIPS/n361 ) );
  MX2XL U10620 ( .A(n10605), .B(n4091), .S0(n3605), .Y(\i_MIPS/n349 ) );
  CLKINVX1 U10621 ( .A(\i_MIPS/n226 ), .Y(n10605) );
  MX2XL U10622 ( .A(n3549), .B(n4093), .S0(n3589), .Y(\i_MIPS/n335 ) );
  MX2XL U10623 ( .A(n10591), .B(n140), .S0(n3590), .Y(\i_MIPS/n307 ) );
  CLKINVX1 U10624 ( .A(\i_MIPS/n184 ), .Y(n10591) );
  MX2XL U10625 ( .A(\D_cache/cache[6][128] ), .B(n10995), .S0(n5372), .Y(
        \D_cache/n766 ) );
  MX2XL U10626 ( .A(\D_cache/cache[5][128] ), .B(n10995), .S0(n5349), .Y(
        \D_cache/n767 ) );
  MX2XL U10627 ( .A(\D_cache/cache[4][128] ), .B(n10995), .S0(n5321), .Y(
        \D_cache/n768 ) );
  MX2XL U10628 ( .A(\D_cache/cache[3][128] ), .B(n10995), .S0(n5276), .Y(
        \D_cache/n769 ) );
  MX2XL U10629 ( .A(\D_cache/cache[2][128] ), .B(n10995), .S0(n5233), .Y(
        \D_cache/n770 ) );
  MX2XL U10630 ( .A(\D_cache/cache[1][128] ), .B(n10995), .S0(n5204), .Y(
        \D_cache/n771 ) );
  MX2XL U10631 ( .A(\D_cache/cache[0][128] ), .B(n10995), .S0(n5165), .Y(
        \D_cache/n772 ) );
  MX2XL U10632 ( .A(n3883), .B(n4081), .S0(n3588), .Y(\i_MIPS/n367 ) );
  MX2XL U10633 ( .A(net104905), .B(net104906), .S0(n3593), .Y(\i_MIPS/n365 )
         );
  CLKINVX1 U10634 ( .A(\i_MIPS/n242 ), .Y(net104905) );
  MX2XL U10635 ( .A(\i_MIPS/Reg_W[4] ), .B(n10846), .S0(n3593), .Y(
        \i_MIPS/n403 ) );
  MX2XL U10636 ( .A(\i_MIPS/Reg_W[3] ), .B(n10847), .S0(n3603), .Y(
        \i_MIPS/n404 ) );
  MX2XL U10637 ( .A(\i_MIPS/Reg_W[2] ), .B(n10849), .S0(n3590), .Y(
        \i_MIPS/n405 ) );
  MXI2XL U10638 ( .A(n4833), .B(n10848), .S0(n3601), .Y(\i_MIPS/n406 ) );
  MX2XL U10639 ( .A(\i_MIPS/Reg_W[0] ), .B(n10850), .S0(n3605), .Y(
        \i_MIPS/n407 ) );
  MX2XL U10640 ( .A(\D_cache/cache[6][153] ), .B(n10770), .S0(n5372), .Y(
        \D_cache/n566 ) );
  MX2XL U10641 ( .A(\D_cache/cache[5][153] ), .B(n10770), .S0(n5349), .Y(
        \D_cache/n567 ) );
  MX2XL U10642 ( .A(\D_cache/cache[4][153] ), .B(n10770), .S0(n5323), .Y(
        \D_cache/n568 ) );
  MX2XL U10643 ( .A(\D_cache/cache[3][153] ), .B(n10770), .S0(n5275), .Y(
        \D_cache/n569 ) );
  MX2XL U10644 ( .A(\D_cache/cache[2][153] ), .B(n10770), .S0(n5235), .Y(
        \D_cache/n570 ) );
  MX2XL U10645 ( .A(\D_cache/cache[1][153] ), .B(n10770), .S0(n5207), .Y(
        \D_cache/n571 ) );
  MX2XL U10646 ( .A(\D_cache/cache[0][153] ), .B(n10770), .S0(n5165), .Y(
        \D_cache/n572 ) );
  MX2XL U10647 ( .A(\D_cache/cache[7][139] ), .B(n10989), .S0(n5416), .Y(
        \D_cache/n677 ) );
  MX2XL U10648 ( .A(\D_cache/cache[6][139] ), .B(n10989), .S0(n5372), .Y(
        \D_cache/n678 ) );
  MX2XL U10649 ( .A(\D_cache/cache[5][139] ), .B(n10989), .S0(n5349), .Y(
        \D_cache/n679 ) );
  MX2XL U10650 ( .A(\D_cache/cache[4][139] ), .B(n10989), .S0(n5321), .Y(
        \D_cache/n680 ) );
  MX2XL U10651 ( .A(\D_cache/cache[3][139] ), .B(n10989), .S0(n5276), .Y(
        \D_cache/n681 ) );
  MX2XL U10652 ( .A(\D_cache/cache[2][139] ), .B(n10989), .S0(n5232), .Y(
        \D_cache/n682 ) );
  MX2XL U10653 ( .A(\D_cache/cache[1][139] ), .B(n10989), .S0(n5207), .Y(
        \D_cache/n683 ) );
  MX2XL U10654 ( .A(\D_cache/cache[0][139] ), .B(n10989), .S0(n5165), .Y(
        \D_cache/n684 ) );
  MX2XL U10655 ( .A(\D_cache/cache[7][151] ), .B(n3794), .S0(n5416), .Y(
        \D_cache/n581 ) );
  MX2XL U10656 ( .A(\D_cache/cache[6][151] ), .B(n11001), .S0(n5372), .Y(
        \D_cache/n582 ) );
  MX2XL U10657 ( .A(\D_cache/cache[5][151] ), .B(n11001), .S0(n5349), .Y(
        \D_cache/n583 ) );
  MX2XL U10658 ( .A(\D_cache/cache[4][151] ), .B(n11001), .S0(n5321), .Y(
        \D_cache/n584 ) );
  MX2XL U10659 ( .A(\D_cache/cache[3][151] ), .B(n3794), .S0(n5275), .Y(
        \D_cache/n585 ) );
  MX2XL U10660 ( .A(\D_cache/cache[2][151] ), .B(n3794), .S0(n5234), .Y(
        \D_cache/n586 ) );
  MX2XL U10661 ( .A(\D_cache/cache[1][151] ), .B(n3794), .S0(n5204), .Y(
        \D_cache/n587 ) );
  MX2XL U10662 ( .A(\D_cache/cache[0][151] ), .B(n11001), .S0(n5165), .Y(
        \D_cache/n588 ) );
  MX2XL U10663 ( .A(\D_cache/cache[7][144] ), .B(n10986), .S0(n5416), .Y(
        \D_cache/n637 ) );
  MX2XL U10664 ( .A(\D_cache/cache[6][144] ), .B(n10986), .S0(n5372), .Y(
        \D_cache/n638 ) );
  MX2XL U10665 ( .A(\D_cache/cache[5][144] ), .B(n10986), .S0(n5350), .Y(
        \D_cache/n639 ) );
  MX2XL U10666 ( .A(\D_cache/cache[4][144] ), .B(n10986), .S0(n5321), .Y(
        \D_cache/n640 ) );
  MX2XL U10667 ( .A(\D_cache/cache[3][144] ), .B(n10986), .S0(n5275), .Y(
        \D_cache/n641 ) );
  MX2XL U10668 ( .A(\D_cache/cache[2][144] ), .B(n10986), .S0(n5233), .Y(
        \D_cache/n642 ) );
  MX2XL U10669 ( .A(\D_cache/cache[1][144] ), .B(n10986), .S0(n5207), .Y(
        \D_cache/n643 ) );
  MX2XL U10670 ( .A(\D_cache/cache[0][144] ), .B(n10986), .S0(n5165), .Y(
        \D_cache/n644 ) );
  MX2XL U10671 ( .A(\D_cache/cache[7][130] ), .B(n11041), .S0(n5417), .Y(
        \D_cache/n749 ) );
  MX2XL U10672 ( .A(\D_cache/cache[6][130] ), .B(n11041), .S0(n5373), .Y(
        \D_cache/n750 ) );
  MX2XL U10673 ( .A(\D_cache/cache[5][130] ), .B(n11041), .S0(n5348), .Y(
        \D_cache/n751 ) );
  MX2XL U10674 ( .A(\D_cache/cache[4][130] ), .B(n11041), .S0(n5322), .Y(
        \D_cache/n752 ) );
  MX2XL U10675 ( .A(\D_cache/cache[3][130] ), .B(n11041), .S0(n5269), .Y(
        \D_cache/n753 ) );
  MX2XL U10676 ( .A(\D_cache/cache[2][130] ), .B(n11041), .S0(n5234), .Y(
        \D_cache/n754 ) );
  MX2XL U10677 ( .A(\D_cache/cache[1][130] ), .B(n11041), .S0(n5206), .Y(
        \D_cache/n755 ) );
  MX2XL U10678 ( .A(\D_cache/cache[0][130] ), .B(n11041), .S0(n5166), .Y(
        \D_cache/n756 ) );
  MX2XL U10679 ( .A(\D_cache/cache[7][152] ), .B(n10992), .S0(n5416), .Y(
        \D_cache/n573 ) );
  MX2XL U10680 ( .A(\D_cache/cache[6][152] ), .B(n10992), .S0(n5372), .Y(
        \D_cache/n574 ) );
  MX2XL U10681 ( .A(\D_cache/cache[5][152] ), .B(n10992), .S0(n3575), .Y(
        \D_cache/n575 ) );
  MX2XL U10682 ( .A(\D_cache/cache[4][152] ), .B(n10992), .S0(n5321), .Y(
        \D_cache/n576 ) );
  MX2XL U10683 ( .A(\D_cache/cache[3][152] ), .B(n10992), .S0(n5275), .Y(
        \D_cache/n577 ) );
  MX2XL U10684 ( .A(\D_cache/cache[2][152] ), .B(n10992), .S0(n5232), .Y(
        \D_cache/n578 ) );
  MX2XL U10685 ( .A(\D_cache/cache[1][152] ), .B(n10992), .S0(n5204), .Y(
        \D_cache/n579 ) );
  MX2XL U10686 ( .A(\D_cache/cache[0][152] ), .B(n10992), .S0(n5165), .Y(
        \D_cache/n580 ) );
  MX2XL U10687 ( .A(\D_cache/cache[7][138] ), .B(n11030), .S0(n5417), .Y(
        \D_cache/n685 ) );
  MX2XL U10688 ( .A(\D_cache/cache[6][138] ), .B(n11030), .S0(n5373), .Y(
        \D_cache/n686 ) );
  MX2XL U10689 ( .A(\D_cache/cache[5][138] ), .B(n11030), .S0(n5348), .Y(
        \D_cache/n687 ) );
  MX2XL U10690 ( .A(\D_cache/cache[4][138] ), .B(n11030), .S0(n5322), .Y(
        \D_cache/n688 ) );
  MX2XL U10691 ( .A(\D_cache/cache[3][138] ), .B(n11030), .S0(n5274), .Y(
        \D_cache/n689 ) );
  MX2XL U10692 ( .A(\D_cache/cache[2][138] ), .B(n11030), .S0(n5234), .Y(
        \D_cache/n690 ) );
  MX2XL U10693 ( .A(\D_cache/cache[1][138] ), .B(n11030), .S0(n5206), .Y(
        \D_cache/n691 ) );
  MX2XL U10694 ( .A(\D_cache/cache[0][138] ), .B(n11030), .S0(n5166), .Y(
        \D_cache/n692 ) );
  MX2XL U10695 ( .A(\D_cache/cache[7][134] ), .B(n11025), .S0(n5417), .Y(
        \D_cache/n717 ) );
  MX2XL U10696 ( .A(\D_cache/cache[6][134] ), .B(n11025), .S0(n5373), .Y(
        \D_cache/n718 ) );
  MX2XL U10697 ( .A(\D_cache/cache[5][134] ), .B(n11025), .S0(n5348), .Y(
        \D_cache/n719 ) );
  MX2XL U10698 ( .A(\D_cache/cache[4][134] ), .B(n11025), .S0(n5322), .Y(
        \D_cache/n720 ) );
  MX2XL U10699 ( .A(\D_cache/cache[3][134] ), .B(n11025), .S0(n5273), .Y(
        \D_cache/n721 ) );
  MX2XL U10700 ( .A(\D_cache/cache[2][134] ), .B(n11025), .S0(n5234), .Y(
        \D_cache/n722 ) );
  MX2XL U10701 ( .A(\D_cache/cache[1][134] ), .B(n11025), .S0(n5206), .Y(
        \D_cache/n723 ) );
  MX2XL U10702 ( .A(\D_cache/cache[0][134] ), .B(n11025), .S0(n5166), .Y(
        \D_cache/n724 ) );
  MX2XL U10703 ( .A(\D_cache/cache[7][131] ), .B(n11044), .S0(n5417), .Y(
        \D_cache/n741 ) );
  MX2XL U10704 ( .A(\D_cache/cache[6][131] ), .B(n11044), .S0(n5373), .Y(
        \D_cache/n742 ) );
  MX2XL U10705 ( .A(\D_cache/cache[5][131] ), .B(n11044), .S0(n5348), .Y(
        \D_cache/n743 ) );
  MX2XL U10706 ( .A(\D_cache/cache[4][131] ), .B(n11044), .S0(n5322), .Y(
        \D_cache/n744 ) );
  MX2XL U10707 ( .A(\D_cache/cache[3][131] ), .B(n11044), .S0(n5272), .Y(
        \D_cache/n745 ) );
  MX2XL U10708 ( .A(\D_cache/cache[2][131] ), .B(n11044), .S0(n5234), .Y(
        \D_cache/n746 ) );
  MX2XL U10709 ( .A(\D_cache/cache[1][131] ), .B(n11044), .S0(n5206), .Y(
        \D_cache/n747 ) );
  MX2XL U10710 ( .A(\D_cache/cache[0][131] ), .B(n11044), .S0(n5166), .Y(
        \D_cache/n748 ) );
  MX2XL U10711 ( .A(\i_MIPS/ID_EX[64] ), .B(n3904), .S0(n3601), .Y(
        \i_MIPS/n321 ) );
  MX2XL U10712 ( .A(\D_cache/cache[7][141] ), .B(n11038), .S0(n5417), .Y(
        \D_cache/n661 ) );
  MX2XL U10713 ( .A(\D_cache/cache[6][141] ), .B(n11038), .S0(n5373), .Y(
        \D_cache/n662 ) );
  MX2XL U10714 ( .A(\D_cache/cache[5][141] ), .B(n11038), .S0(n5348), .Y(
        \D_cache/n663 ) );
  MX2XL U10715 ( .A(\D_cache/cache[4][141] ), .B(n11038), .S0(n5322), .Y(
        \D_cache/n664 ) );
  MX2XL U10716 ( .A(\D_cache/cache[3][141] ), .B(n11038), .S0(n5275), .Y(
        \D_cache/n665 ) );
  MX2XL U10717 ( .A(\D_cache/cache[2][141] ), .B(n11038), .S0(n5234), .Y(
        \D_cache/n666 ) );
  MX2XL U10718 ( .A(\D_cache/cache[1][141] ), .B(n11038), .S0(n5206), .Y(
        \D_cache/n667 ) );
  MX2XL U10719 ( .A(\D_cache/cache[0][141] ), .B(n11038), .S0(n5166), .Y(
        \D_cache/n668 ) );
  MX2XL U10720 ( .A(\D_cache/cache[7][129] ), .B(n11047), .S0(n5417), .Y(
        \D_cache/n757 ) );
  MX2XL U10721 ( .A(\D_cache/cache[6][129] ), .B(n11047), .S0(n5373), .Y(
        \D_cache/n758 ) );
  MX2XL U10722 ( .A(\D_cache/cache[5][129] ), .B(n11047), .S0(n5348), .Y(
        \D_cache/n759 ) );
  MX2XL U10723 ( .A(\D_cache/cache[4][129] ), .B(n11047), .S0(n5322), .Y(
        \D_cache/n760 ) );
  MX2XL U10724 ( .A(\D_cache/cache[3][129] ), .B(n11047), .S0(n5272), .Y(
        \D_cache/n761 ) );
  MX2XL U10725 ( .A(\D_cache/cache[2][129] ), .B(n11047), .S0(n5234), .Y(
        \D_cache/n762 ) );
  MX2XL U10726 ( .A(\D_cache/cache[1][129] ), .B(n11047), .S0(n5206), .Y(
        \D_cache/n763 ) );
  MX2XL U10727 ( .A(\D_cache/cache[0][129] ), .B(n11047), .S0(n5166), .Y(
        \D_cache/n764 ) );
  MX2XL U10728 ( .A(\D_cache/cache[7][137] ), .B(n11010), .S0(n5416), .Y(
        \D_cache/n693 ) );
  MX2XL U10729 ( .A(\D_cache/cache[6][137] ), .B(n11010), .S0(n5372), .Y(
        \D_cache/n694 ) );
  MX2XL U10730 ( .A(\D_cache/cache[5][137] ), .B(n11010), .S0(n3575), .Y(
        \D_cache/n695 ) );
  MX2XL U10731 ( .A(\D_cache/cache[4][137] ), .B(n11010), .S0(n5321), .Y(
        \D_cache/n696 ) );
  MX2XL U10732 ( .A(\D_cache/cache[3][137] ), .B(n11010), .S0(n5269), .Y(
        \D_cache/n697 ) );
  MX2XL U10733 ( .A(\D_cache/cache[2][137] ), .B(n11010), .S0(n5233), .Y(
        \D_cache/n698 ) );
  MX2XL U10734 ( .A(\D_cache/cache[1][137] ), .B(n11010), .S0(n5208), .Y(
        \D_cache/n699 ) );
  MX2XL U10735 ( .A(\D_cache/cache[0][137] ), .B(n11010), .S0(n5165), .Y(
        \D_cache/n700 ) );
  MX2XL U10736 ( .A(\D_cache/cache[7][133] ), .B(n11027), .S0(n5417), .Y(
        \D_cache/n725 ) );
  MX2XL U10737 ( .A(\D_cache/cache[6][133] ), .B(n11027), .S0(n5373), .Y(
        \D_cache/n726 ) );
  MX2XL U10738 ( .A(\D_cache/cache[5][133] ), .B(n11027), .S0(n5348), .Y(
        \D_cache/n727 ) );
  MX2XL U10739 ( .A(\D_cache/cache[4][133] ), .B(n11027), .S0(n5322), .Y(
        \D_cache/n728 ) );
  MX2XL U10740 ( .A(\D_cache/cache[3][133] ), .B(n11027), .S0(n5270), .Y(
        \D_cache/n729 ) );
  MX2XL U10741 ( .A(\D_cache/cache[2][133] ), .B(n11027), .S0(n5234), .Y(
        \D_cache/n730 ) );
  MX2XL U10742 ( .A(\D_cache/cache[1][133] ), .B(n11027), .S0(n5206), .Y(
        \D_cache/n731 ) );
  MX2XL U10743 ( .A(\D_cache/cache[0][133] ), .B(n11027), .S0(n5166), .Y(
        \D_cache/n732 ) );
  MX2XL U10744 ( .A(\D_cache/cache[7][132] ), .B(n11016), .S0(n5417), .Y(
        \D_cache/n733 ) );
  MX2XL U10745 ( .A(\D_cache/cache[6][132] ), .B(n11016), .S0(n5373), .Y(
        \D_cache/n734 ) );
  MX2XL U10746 ( .A(\D_cache/cache[5][132] ), .B(n11016), .S0(n5348), .Y(
        \D_cache/n735 ) );
  MX2XL U10747 ( .A(\D_cache/cache[4][132] ), .B(n11016), .S0(n5322), .Y(
        \D_cache/n736 ) );
  MX2XL U10748 ( .A(\D_cache/cache[3][132] ), .B(n11016), .S0(n5268), .Y(
        \D_cache/n737 ) );
  MX2XL U10749 ( .A(\D_cache/cache[2][132] ), .B(n11016), .S0(n5234), .Y(
        \D_cache/n738 ) );
  MX2XL U10750 ( .A(\D_cache/cache[1][132] ), .B(n11016), .S0(n5206), .Y(
        \D_cache/n739 ) );
  MX2XL U10751 ( .A(\D_cache/cache[0][132] ), .B(n11016), .S0(n5166), .Y(
        \D_cache/n740 ) );
  MX2XL U10752 ( .A(\D_cache/cache[7][136] ), .B(n10998), .S0(n5416), .Y(
        \D_cache/n701 ) );
  MX2XL U10753 ( .A(\D_cache/cache[6][136] ), .B(n10998), .S0(n5372), .Y(
        \D_cache/n702 ) );
  MX2XL U10754 ( .A(\D_cache/cache[5][136] ), .B(n10998), .S0(n3575), .Y(
        \D_cache/n703 ) );
  MX2XL U10755 ( .A(\D_cache/cache[4][136] ), .B(n10998), .S0(n5321), .Y(
        \D_cache/n704 ) );
  MX2XL U10756 ( .A(\D_cache/cache[3][136] ), .B(n10998), .S0(n5276), .Y(
        \D_cache/n705 ) );
  MX2XL U10757 ( .A(\D_cache/cache[2][136] ), .B(n10998), .S0(n5235), .Y(
        \D_cache/n706 ) );
  MX2XL U10758 ( .A(\D_cache/cache[1][136] ), .B(n10998), .S0(n5207), .Y(
        \D_cache/n707 ) );
  MX2XL U10759 ( .A(\D_cache/cache[0][136] ), .B(n10998), .S0(n5165), .Y(
        \D_cache/n708 ) );
  MX2XL U10760 ( .A(\D_cache/cache[7][140] ), .B(n10983), .S0(n5416), .Y(
        \D_cache/n669 ) );
  MX2XL U10761 ( .A(\D_cache/cache[6][140] ), .B(n10983), .S0(n5372), .Y(
        \D_cache/n670 ) );
  MX2XL U10762 ( .A(\D_cache/cache[5][140] ), .B(n10983), .S0(n3575), .Y(
        \D_cache/n671 ) );
  MX2XL U10763 ( .A(\D_cache/cache[4][140] ), .B(n10983), .S0(n5321), .Y(
        \D_cache/n672 ) );
  MX2XL U10764 ( .A(\D_cache/cache[3][140] ), .B(n10983), .S0(n5274), .Y(
        \D_cache/n673 ) );
  MX2XL U10765 ( .A(\D_cache/cache[2][140] ), .B(n10983), .S0(n5230), .Y(
        \D_cache/n674 ) );
  MX2XL U10766 ( .A(\D_cache/cache[1][140] ), .B(n10983), .S0(n5204), .Y(
        \D_cache/n675 ) );
  MX2XL U10767 ( .A(\D_cache/cache[0][140] ), .B(n10983), .S0(n5165), .Y(
        \D_cache/n676 ) );
  MX2XL U10768 ( .A(\D_cache/cache[6][150] ), .B(n11022), .S0(n5373), .Y(
        \D_cache/n590 ) );
  MX2XL U10769 ( .A(\D_cache/cache[5][150] ), .B(n11022), .S0(n5348), .Y(
        \D_cache/n591 ) );
  MX2XL U10770 ( .A(\D_cache/cache[4][150] ), .B(n11022), .S0(n5322), .Y(
        \D_cache/n592 ) );
  MX2XL U10771 ( .A(\D_cache/cache[3][150] ), .B(n11022), .S0(n5269), .Y(
        \D_cache/n593 ) );
  MX2XL U10772 ( .A(\D_cache/cache[2][150] ), .B(n11022), .S0(n5234), .Y(
        \D_cache/n594 ) );
  MX2XL U10773 ( .A(\D_cache/cache[1][150] ), .B(n11022), .S0(n5206), .Y(
        \D_cache/n595 ) );
  MX2XL U10774 ( .A(\D_cache/cache[0][150] ), .B(n11022), .S0(n5166), .Y(
        \D_cache/n596 ) );
  MX2XL U10775 ( .A(\D_cache/cache[6][147] ), .B(n11004), .S0(n5372), .Y(
        \D_cache/n614 ) );
  MX2XL U10776 ( .A(\D_cache/cache[5][147] ), .B(n11004), .S0(n5345), .Y(
        \D_cache/n615 ) );
  MX2XL U10777 ( .A(\D_cache/cache[4][147] ), .B(n11004), .S0(n5321), .Y(
        \D_cache/n616 ) );
  MX2XL U10778 ( .A(\D_cache/cache[3][147] ), .B(n11004), .S0(n5272), .Y(
        \D_cache/n617 ) );
  MX2XL U10779 ( .A(\D_cache/cache[2][147] ), .B(n11004), .S0(n5231), .Y(
        \D_cache/n618 ) );
  MX2XL U10780 ( .A(\D_cache/cache[1][147] ), .B(n11004), .S0(n5207), .Y(
        \D_cache/n619 ) );
  MX2XL U10781 ( .A(\D_cache/cache[0][147] ), .B(n11004), .S0(n5165), .Y(
        \D_cache/n620 ) );
  MX2XL U10782 ( .A(\D_cache/cache[7][145] ), .B(n11019), .S0(n5417), .Y(
        \D_cache/n629 ) );
  MX2XL U10783 ( .A(\D_cache/cache[6][145] ), .B(n11019), .S0(n5373), .Y(
        \D_cache/n630 ) );
  MX2XL U10784 ( .A(\D_cache/cache[5][145] ), .B(n11019), .S0(n5348), .Y(
        \D_cache/n631 ) );
  MX2XL U10785 ( .A(\D_cache/cache[4][145] ), .B(n11019), .S0(n5322), .Y(
        \D_cache/n632 ) );
  MX2XL U10786 ( .A(\D_cache/cache[3][145] ), .B(n11019), .S0(n5273), .Y(
        \D_cache/n633 ) );
  MX2XL U10787 ( .A(\D_cache/cache[2][145] ), .B(n11019), .S0(n5234), .Y(
        \D_cache/n634 ) );
  MX2XL U10788 ( .A(\D_cache/cache[1][145] ), .B(n11019), .S0(n5206), .Y(
        \D_cache/n635 ) );
  MX2XL U10789 ( .A(\D_cache/cache[0][145] ), .B(n11019), .S0(n5166), .Y(
        \D_cache/n636 ) );
  MX2XL U10790 ( .A(\D_cache/cache[6][135] ), .B(n11008), .S0(n5372), .Y(
        \D_cache/n710 ) );
  MX2XL U10791 ( .A(\D_cache/cache[5][135] ), .B(n11008), .S0(n5345), .Y(
        \D_cache/n711 ) );
  MX2XL U10792 ( .A(\D_cache/cache[4][135] ), .B(n11008), .S0(n5321), .Y(
        \D_cache/n712 ) );
  MX2XL U10793 ( .A(\D_cache/cache[3][135] ), .B(n11008), .S0(n5275), .Y(
        \D_cache/n713 ) );
  MX2XL U10794 ( .A(\D_cache/cache[2][135] ), .B(n11008), .S0(n5235), .Y(
        \D_cache/n714 ) );
  MX2XL U10795 ( .A(\D_cache/cache[1][135] ), .B(n11008), .S0(n5204), .Y(
        \D_cache/n715 ) );
  MX2XL U10796 ( .A(\D_cache/cache[0][135] ), .B(n11008), .S0(n5165), .Y(
        \D_cache/n716 ) );
  MX2XL U10797 ( .A(\I_cache/cache[5][152] ), .B(n11068), .S0(n5758), .Y(
        n11624) );
  MX2XL U10798 ( .A(\I_cache/cache[4][152] ), .B(n11068), .S0(n5804), .Y(
        n11625) );
  MX2XL U10799 ( .A(\I_cache/cache[2][152] ), .B(n11068), .S0(n5714), .Y(
        n11627) );
  MX2XL U10800 ( .A(\I_cache/cache[0][152] ), .B(n11068), .S0(n5623), .Y(
        n11629) );
  MX2XL U10801 ( .A(\I_cache/cache[6][151] ), .B(n11066), .S0(n5891), .Y(
        n11631) );
  MX2XL U10802 ( .A(\I_cache/cache[5][151] ), .B(n11066), .S0(n5758), .Y(
        n11632) );
  MX2XL U10803 ( .A(\I_cache/cache[4][151] ), .B(n11066), .S0(n5804), .Y(
        n11633) );
  MX2XL U10804 ( .A(\I_cache/cache[3][151] ), .B(n11066), .S0(n5669), .Y(
        n11634) );
  MX2XL U10805 ( .A(\I_cache/cache[1][151] ), .B(n11066), .S0(n5580), .Y(
        n11636) );
  MX2XL U10806 ( .A(\I_cache/cache[5][149] ), .B(n11187), .S0(n5758), .Y(
        n11648) );
  MX2XL U10807 ( .A(\I_cache/cache[4][149] ), .B(n11187), .S0(n5805), .Y(
        n11649) );
  MX2XL U10808 ( .A(\I_cache/cache[5][148] ), .B(n11197), .S0(n5758), .Y(
        n11656) );
  MX2XL U10809 ( .A(\I_cache/cache[4][148] ), .B(n11197), .S0(n5805), .Y(
        n11657) );
  MX2XL U10810 ( .A(\I_cache/cache[5][147] ), .B(n11192), .S0(n5759), .Y(
        n11664) );
  MX2XL U10811 ( .A(\I_cache/cache[4][147] ), .B(n11192), .S0(n5805), .Y(
        n11665) );
  MX2XL U10812 ( .A(\I_cache/cache[6][145] ), .B(n11065), .S0(n5893), .Y(
        n11679) );
  MX2XL U10813 ( .A(\I_cache/cache[5][145] ), .B(n11065), .S0(n5759), .Y(
        n11680) );
  MX2XL U10814 ( .A(\I_cache/cache[4][145] ), .B(n11065), .S0(n5806), .Y(
        n11681) );
  MX2XL U10815 ( .A(\I_cache/cache[3][145] ), .B(n11065), .S0(n5671), .Y(
        n11682) );
  MX2XL U10816 ( .A(\I_cache/cache[1][145] ), .B(n11065), .S0(n5582), .Y(
        n11684) );
  MX2XL U10817 ( .A(\I_cache/cache[5][144] ), .B(n11145), .S0(n5757), .Y(
        n11688) );
  MX2XL U10818 ( .A(\I_cache/cache[4][144] ), .B(n11145), .S0(n5803), .Y(
        n11689) );
  MX2XL U10819 ( .A(\I_cache/cache[7][143] ), .B(n11215), .S0(n5844), .Y(
        n11694) );
  MX2XL U10820 ( .A(\I_cache/cache[6][143] ), .B(n11215), .S0(n5888), .Y(
        n11695) );
  MX2XL U10821 ( .A(\I_cache/cache[6][142] ), .B(n11201), .S0(n5892), .Y(
        n11703) );
  MX2XL U10822 ( .A(\I_cache/cache[5][142] ), .B(n11201), .S0(n5758), .Y(
        n11704) );
  MX2XL U10823 ( .A(\I_cache/cache[4][142] ), .B(n11201), .S0(n5805), .Y(
        n11705) );
  MX2XL U10824 ( .A(\I_cache/cache[3][142] ), .B(n11201), .S0(n5670), .Y(
        n11706) );
  MX2XL U10825 ( .A(\I_cache/cache[2][142] ), .B(n11201), .S0(n5715), .Y(
        n11707) );
  MX2XL U10826 ( .A(\I_cache/cache[1][142] ), .B(n11201), .S0(n5581), .Y(
        n11708) );
  MX2XL U10827 ( .A(\I_cache/cache[7][141] ), .B(n11206), .S0(n5849), .Y(
        n11710) );
  MX2XL U10828 ( .A(\I_cache/cache[6][141] ), .B(n11206), .S0(n5892), .Y(
        n11711) );
  MX2XL U10829 ( .A(\I_cache/cache[5][141] ), .B(n11206), .S0(n5756), .Y(
        n11712) );
  MX2XL U10830 ( .A(\I_cache/cache[4][141] ), .B(n11206), .S0(n5805), .Y(
        n11713) );
  MX2XL U10831 ( .A(\I_cache/cache[3][141] ), .B(n11206), .S0(n5670), .Y(
        n11714) );
  MX2XL U10832 ( .A(\I_cache/cache[2][141] ), .B(n11206), .S0(n5715), .Y(
        n11715) );
  MX2XL U10833 ( .A(\I_cache/cache[1][141] ), .B(n11206), .S0(n5581), .Y(
        n11716) );
  MX2XL U10834 ( .A(\I_cache/cache[0][141] ), .B(n11206), .S0(n5624), .Y(
        n11717) );
  MX2XL U10835 ( .A(\I_cache/cache[5][140] ), .B(n11150), .S0(n5759), .Y(
        n11720) );
  MX2XL U10836 ( .A(\I_cache/cache[4][140] ), .B(n11150), .S0(n5805), .Y(
        n11721) );
  MX2XL U10837 ( .A(\I_cache/cache[5][139] ), .B(n11140), .S0(n5758), .Y(
        n11728) );
  MX2XL U10838 ( .A(\I_cache/cache[4][139] ), .B(n11140), .S0(n5804), .Y(
        n11729) );
  MX2XL U10839 ( .A(\I_cache/cache[5][138] ), .B(n11131), .S0(n5758), .Y(
        n11736) );
  MX2XL U10840 ( .A(\I_cache/cache[4][138] ), .B(n11131), .S0(n5804), .Y(
        n11737) );
  MX2XL U10841 ( .A(\I_cache/cache[3][138] ), .B(n11131), .S0(n5669), .Y(
        n11738) );
  MX2XL U10842 ( .A(\I_cache/cache[5][137] ), .B(n11172), .S0(n5758), .Y(
        n11744) );
  MX2XL U10843 ( .A(\I_cache/cache[4][137] ), .B(n11172), .S0(n5805), .Y(
        n11745) );
  MX2XL U10844 ( .A(\I_cache/cache[5][136] ), .B(n11182), .S0(n5759), .Y(
        n11752) );
  MX2XL U10845 ( .A(\I_cache/cache[4][136] ), .B(n11182), .S0(n5805), .Y(
        n11753) );
  MX2XL U10846 ( .A(\I_cache/cache[5][135] ), .B(n11177), .S0(n5758), .Y(
        n11760) );
  MX2XL U10847 ( .A(\I_cache/cache[4][135] ), .B(n11177), .S0(n5805), .Y(
        n11761) );
  MX2XL U10848 ( .A(\I_cache/cache[5][134] ), .B(n11122), .S0(n5758), .Y(
        n11768) );
  MX2XL U10849 ( .A(\I_cache/cache[4][134] ), .B(n11122), .S0(n5804), .Y(
        n11769) );
  MX2XL U10850 ( .A(\I_cache/cache[5][132] ), .B(n11118), .S0(n5758), .Y(
        n11784) );
  MX2XL U10851 ( .A(\I_cache/cache[4][132] ), .B(n11118), .S0(n5804), .Y(
        n11785) );
  MX2XL U10852 ( .A(\I_cache/cache[5][129] ), .B(n11164), .S0(n5759), .Y(
        n11808) );
  MX2XL U10853 ( .A(\I_cache/cache[4][129] ), .B(n11164), .S0(n5805), .Y(
        n11809) );
  MX2XL U10854 ( .A(\I_cache/cache[7][133] ), .B(n11127), .S0(n5848), .Y(
        n11774) );
  MX2XL U10855 ( .A(\I_cache/cache[6][133] ), .B(n11127), .S0(n5891), .Y(
        n11775) );
  MX2XL U10856 ( .A(\I_cache/cache[5][131] ), .B(n11159), .S0(n5758), .Y(
        n11792) );
  MX2XL U10857 ( .A(\I_cache/cache[4][131] ), .B(n11159), .S0(n5805), .Y(
        n11793) );
  MX2XL U10858 ( .A(\I_cache/cache[5][130] ), .B(n11155), .S0(n5759), .Y(
        n11800) );
  MX2XL U10859 ( .A(\I_cache/cache[4][130] ), .B(n11155), .S0(n5805), .Y(
        n11801) );
  MX2XL U10860 ( .A(\I_cache/cache[5][128] ), .B(n11067), .S0(n5758), .Y(
        n11816) );
  MX2XL U10861 ( .A(\I_cache/cache[4][128] ), .B(n11067), .S0(n5804), .Y(
        n11817) );
  CLKMX2X2 U10862 ( .A(\I_cache/cache[7][127] ), .B(n6587), .S0(n5850), .Y(
        n11822) );
  CLKMX2X2 U10863 ( .A(\I_cache/cache[6][127] ), .B(n6587), .S0(n5893), .Y(
        n11823) );
  CLKMX2X2 U10864 ( .A(\I_cache/cache[5][127] ), .B(n6587), .S0(n5752), .Y(
        n11824) );
  CLKMX2X2 U10865 ( .A(\I_cache/cache[4][127] ), .B(n6587), .S0(n5806), .Y(
        n11825) );
  CLKMX2X2 U10866 ( .A(\I_cache/cache[3][127] ), .B(n6587), .S0(n5665), .Y(
        n11826) );
  CLKMX2X2 U10867 ( .A(\I_cache/cache[2][127] ), .B(n6587), .S0(n5716), .Y(
        n11827) );
  CLKMX2X2 U10868 ( .A(\I_cache/cache[1][127] ), .B(n6587), .S0(n5577), .Y(
        n11828) );
  CLKMX2X2 U10869 ( .A(\I_cache/cache[0][127] ), .B(n6587), .S0(n5623), .Y(
        n11829) );
  CLKMX2X2 U10870 ( .A(\I_cache/cache[7][126] ), .B(n9676), .S0(n5844), .Y(
        n11830) );
  CLKMX2X2 U10871 ( .A(\I_cache/cache[6][126] ), .B(n9676), .S0(n5888), .Y(
        n11831) );
  CLKMX2X2 U10872 ( .A(\I_cache/cache[5][126] ), .B(n9676), .S0(n5753), .Y(
        n11832) );
  CLKMX2X2 U10873 ( .A(\I_cache/cache[4][126] ), .B(n9676), .S0(n5802), .Y(
        n11833) );
  CLKMX2X2 U10874 ( .A(\I_cache/cache[3][126] ), .B(n9676), .S0(n5667), .Y(
        n11834) );
  CLKMX2X2 U10875 ( .A(\I_cache/cache[2][126] ), .B(n9676), .S0(n5709), .Y(
        n11835) );
  CLKMX2X2 U10876 ( .A(\I_cache/cache[1][126] ), .B(n9676), .S0(n5574), .Y(
        n11836) );
  CLKMX2X2 U10877 ( .A(\I_cache/cache[0][126] ), .B(n9676), .S0(n5617), .Y(
        n11837) );
  CLKMX2X2 U10878 ( .A(\I_cache/cache[7][125] ), .B(n9698), .S0(n5842), .Y(
        n11838) );
  CLKMX2X2 U10879 ( .A(\I_cache/cache[6][125] ), .B(n9698), .S0(n5885), .Y(
        n11839) );
  CLKMX2X2 U10880 ( .A(\I_cache/cache[5][125] ), .B(n9698), .S0(n5754), .Y(
        n11840) );
  CLKMX2X2 U10881 ( .A(\I_cache/cache[4][125] ), .B(n9698), .S0(n5798), .Y(
        n11841) );
  CLKMX2X2 U10882 ( .A(\I_cache/cache[3][125] ), .B(n9698), .S0(n5663), .Y(
        n11842) );
  CLKMX2X2 U10883 ( .A(\I_cache/cache[2][125] ), .B(n9698), .S0(n5708), .Y(
        n11843) );
  CLKMX2X2 U10884 ( .A(\I_cache/cache[1][125] ), .B(n9698), .S0(n5574), .Y(
        n11844) );
  CLKMX2X2 U10885 ( .A(\I_cache/cache[0][125] ), .B(n9698), .S0(n5617), .Y(
        n11845) );
  CLKMX2X2 U10886 ( .A(\I_cache/cache[7][124] ), .B(n9646), .S0(n5850), .Y(
        n11846) );
  CLKMX2X2 U10887 ( .A(\I_cache/cache[6][124] ), .B(n9646), .S0(n5887), .Y(
        n11847) );
  CLKMX2X2 U10888 ( .A(\I_cache/cache[5][124] ), .B(n9646), .S0(n5753), .Y(
        n11848) );
  CLKMX2X2 U10889 ( .A(\I_cache/cache[4][124] ), .B(n9646), .S0(n5799), .Y(
        n11849) );
  CLKMX2X2 U10890 ( .A(\I_cache/cache[3][124] ), .B(n9646), .S0(n5663), .Y(
        n11850) );
  CLKMX2X2 U10891 ( .A(\I_cache/cache[2][124] ), .B(n9646), .S0(n5709), .Y(
        n11851) );
  CLKMX2X2 U10892 ( .A(\I_cache/cache[1][124] ), .B(n9646), .S0(n5575), .Y(
        n11852) );
  CLKMX2X2 U10893 ( .A(\I_cache/cache[0][124] ), .B(n9646), .S0(n5619), .Y(
        n11853) );
  CLKMX2X2 U10894 ( .A(\I_cache/cache[7][123] ), .B(n9624), .S0(n5846), .Y(
        n11854) );
  CLKMX2X2 U10895 ( .A(\I_cache/cache[6][123] ), .B(n9624), .S0(n5887), .Y(
        n11855) );
  CLKMX2X2 U10896 ( .A(\I_cache/cache[5][123] ), .B(n9624), .S0(n5753), .Y(
        n11856) );
  CLKMX2X2 U10897 ( .A(\I_cache/cache[4][123] ), .B(n9624), .S0(n5802), .Y(
        n11857) );
  CLKMX2X2 U10898 ( .A(\I_cache/cache[3][123] ), .B(n9624), .S0(n5665), .Y(
        n11858) );
  CLKMX2X2 U10899 ( .A(\I_cache/cache[2][123] ), .B(n9624), .S0(n5709), .Y(
        n11859) );
  CLKMX2X2 U10900 ( .A(\I_cache/cache[1][123] ), .B(n9624), .S0(n5575), .Y(
        n11860) );
  CLKMX2X2 U10901 ( .A(\I_cache/cache[0][123] ), .B(n9624), .S0(n5617), .Y(
        n11861) );
  CLKMX2X2 U10902 ( .A(\I_cache/cache[7][122] ), .B(n6602), .S0(n5847), .Y(
        n11862) );
  CLKMX2X2 U10903 ( .A(\I_cache/cache[6][122] ), .B(n6602), .S0(n5887), .Y(
        n11863) );
  CLKMX2X2 U10904 ( .A(\I_cache/cache[5][122] ), .B(n6602), .S0(n5753), .Y(
        n11864) );
  CLKMX2X2 U10905 ( .A(\I_cache/cache[4][122] ), .B(n6602), .S0(n5800), .Y(
        n11865) );
  CLKMX2X2 U10906 ( .A(\I_cache/cache[3][122] ), .B(n6602), .S0(n5667), .Y(
        n11866) );
  CLKMX2X2 U10907 ( .A(\I_cache/cache[2][122] ), .B(n6602), .S0(n5709), .Y(
        n11867) );
  CLKMX2X2 U10908 ( .A(\I_cache/cache[1][122] ), .B(n6602), .S0(n5579), .Y(
        n11868) );
  CLKMX2X2 U10909 ( .A(\I_cache/cache[0][122] ), .B(n6602), .S0(n5620), .Y(
        n11869) );
  CLKMX2X2 U10910 ( .A(\I_cache/cache[7][121] ), .B(n10043), .S0(n5844), .Y(
        n11870) );
  CLKMX2X2 U10911 ( .A(\I_cache/cache[6][121] ), .B(n10043), .S0(n5888), .Y(
        n11871) );
  CLKMX2X2 U10912 ( .A(\I_cache/cache[5][121] ), .B(n10043), .S0(n5754), .Y(
        n11872) );
  CLKMX2X2 U10913 ( .A(\I_cache/cache[4][121] ), .B(n10043), .S0(n5800), .Y(
        n11873) );
  CLKMX2X2 U10914 ( .A(\I_cache/cache[3][121] ), .B(n10043), .S0(n5665), .Y(
        n11874) );
  CLKMX2X2 U10915 ( .A(\I_cache/cache[2][121] ), .B(n10043), .S0(n5710), .Y(
        n11875) );
  CLKMX2X2 U10916 ( .A(\I_cache/cache[1][121] ), .B(n10043), .S0(n5576), .Y(
        n11876) );
  CLKMX2X2 U10917 ( .A(\I_cache/cache[0][121] ), .B(n10043), .S0(n5619), .Y(
        n11877) );
  CLKMX2X2 U10918 ( .A(\I_cache/cache[7][120] ), .B(n10838), .S0(n5850), .Y(
        n11878) );
  CLKMX2X2 U10919 ( .A(\I_cache/cache[6][120] ), .B(n10838), .S0(n5893), .Y(
        n11879) );
  CLKMX2X2 U10920 ( .A(\I_cache/cache[5][120] ), .B(n10838), .S0(n5759), .Y(
        n11880) );
  CLKMX2X2 U10921 ( .A(\I_cache/cache[4][120] ), .B(n10838), .S0(n5806), .Y(
        n11881) );
  CLKMX2X2 U10922 ( .A(\I_cache/cache[3][120] ), .B(n10838), .S0(n5671), .Y(
        n11882) );
  CLKMX2X2 U10923 ( .A(\I_cache/cache[2][120] ), .B(n10838), .S0(n5716), .Y(
        n11883) );
  CLKMX2X2 U10924 ( .A(\I_cache/cache[1][120] ), .B(n10838), .S0(n5582), .Y(
        n11884) );
  CLKMX2X2 U10925 ( .A(\I_cache/cache[0][120] ), .B(n10838), .S0(n5625), .Y(
        n11885) );
  CLKMX2X2 U10926 ( .A(\I_cache/cache[7][119] ), .B(n10021), .S0(n5844), .Y(
        n11886) );
  CLKMX2X2 U10927 ( .A(\I_cache/cache[6][119] ), .B(n10021), .S0(n5888), .Y(
        n11887) );
  CLKMX2X2 U10928 ( .A(\I_cache/cache[5][119] ), .B(n10021), .S0(n5754), .Y(
        n11888) );
  CLKMX2X2 U10929 ( .A(\I_cache/cache[4][119] ), .B(n10021), .S0(n5800), .Y(
        n11889) );
  CLKMX2X2 U10930 ( .A(\I_cache/cache[3][119] ), .B(n10021), .S0(n5665), .Y(
        n11890) );
  CLKMX2X2 U10931 ( .A(\I_cache/cache[2][119] ), .B(n10021), .S0(n5710), .Y(
        n11891) );
  CLKMX2X2 U10932 ( .A(\I_cache/cache[1][119] ), .B(n10021), .S0(n5576), .Y(
        n11892) );
  CLKMX2X2 U10933 ( .A(\I_cache/cache[0][119] ), .B(n10021), .S0(n5619), .Y(
        n11893) );
  CLKMX2X2 U10934 ( .A(\I_cache/cache[7][118] ), .B(n9977), .S0(n5847), .Y(
        n11894) );
  CLKMX2X2 U10935 ( .A(\I_cache/cache[6][118] ), .B(n9977), .S0(n5890), .Y(
        n11895) );
  CLKMX2X2 U10936 ( .A(\I_cache/cache[5][118] ), .B(n9977), .S0(n5757), .Y(
        n11896) );
  CLKMX2X2 U10937 ( .A(\I_cache/cache[4][118] ), .B(n9977), .S0(n5803), .Y(
        n11897) );
  CLKMX2X2 U10938 ( .A(\I_cache/cache[3][118] ), .B(n9977), .S0(n5668), .Y(
        n11898) );
  CLKMX2X2 U10939 ( .A(\I_cache/cache[2][118] ), .B(n9977), .S0(n5713), .Y(
        n11899) );
  CLKMX2X2 U10940 ( .A(\I_cache/cache[1][118] ), .B(n9977), .S0(n5579), .Y(
        n11900) );
  CLKMX2X2 U10941 ( .A(\I_cache/cache[0][118] ), .B(n9977), .S0(n5622), .Y(
        n11901) );
  CLKMX2X2 U10942 ( .A(\I_cache/cache[7][117] ), .B(n9999), .S0(n5847), .Y(
        n11902) );
  CLKMX2X2 U10943 ( .A(\I_cache/cache[6][117] ), .B(n9999), .S0(n5890), .Y(
        n11903) );
  CLKMX2X2 U10944 ( .A(\I_cache/cache[5][117] ), .B(n9999), .S0(n5757), .Y(
        n11904) );
  CLKMX2X2 U10945 ( .A(\I_cache/cache[4][117] ), .B(n9999), .S0(n5803), .Y(
        n11905) );
  CLKMX2X2 U10946 ( .A(\I_cache/cache[3][117] ), .B(n9999), .S0(n5668), .Y(
        n11906) );
  CLKMX2X2 U10947 ( .A(\I_cache/cache[2][117] ), .B(n9999), .S0(n5713), .Y(
        n11907) );
  CLKMX2X2 U10948 ( .A(\I_cache/cache[1][117] ), .B(n9999), .S0(n5579), .Y(
        n11908) );
  CLKMX2X2 U10949 ( .A(\I_cache/cache[0][117] ), .B(n9999), .S0(n5621), .Y(
        n11909) );
  CLKMX2X2 U10950 ( .A(\I_cache/cache[7][116] ), .B(n9788), .S0(n5843), .Y(
        n11910) );
  CLKMX2X2 U10951 ( .A(\I_cache/cache[6][116] ), .B(n9788), .S0(n5886), .Y(
        n11911) );
  CLKMX2X2 U10952 ( .A(\I_cache/cache[5][116] ), .B(n9788), .S0(n5752), .Y(
        n11912) );
  CLKMX2X2 U10953 ( .A(\I_cache/cache[4][116] ), .B(n9788), .S0(n5799), .Y(
        n11913) );
  CLKMX2X2 U10954 ( .A(\I_cache/cache[3][116] ), .B(n9788), .S0(n5664), .Y(
        n11914) );
  CLKMX2X2 U10955 ( .A(\I_cache/cache[2][116] ), .B(n9788), .S0(n5709), .Y(
        n11915) );
  CLKMX2X2 U10956 ( .A(\I_cache/cache[1][116] ), .B(n9788), .S0(n5578), .Y(
        n11916) );
  CLKMX2X2 U10957 ( .A(\I_cache/cache[0][116] ), .B(n9788), .S0(n5618), .Y(
        n11917) );
  CLKMX2X2 U10958 ( .A(\I_cache/cache[7][115] ), .B(n11086), .S0(n5848), .Y(
        n11918) );
  CLKMX2X2 U10959 ( .A(\I_cache/cache[6][115] ), .B(n11086), .S0(n5891), .Y(
        n11919) );
  CLKMX2X2 U10960 ( .A(\I_cache/cache[5][115] ), .B(n11086), .S0(n5758), .Y(
        n11920) );
  CLKMX2X2 U10961 ( .A(\I_cache/cache[4][115] ), .B(n11086), .S0(n5804), .Y(
        n11921) );
  CLKMX2X2 U10962 ( .A(\I_cache/cache[3][115] ), .B(n11086), .S0(n5669), .Y(
        n11922) );
  CLKMX2X2 U10963 ( .A(\I_cache/cache[2][115] ), .B(n11086), .S0(n5714), .Y(
        n11923) );
  CLKMX2X2 U10964 ( .A(\I_cache/cache[1][115] ), .B(n11086), .S0(n5580), .Y(
        n11924) );
  CLKMX2X2 U10965 ( .A(\I_cache/cache[0][115] ), .B(n11086), .S0(n5623), .Y(
        n11925) );
  CLKMX2X2 U10966 ( .A(\I_cache/cache[7][114] ), .B(n9772), .S0(n5843), .Y(
        n11926) );
  CLKMX2X2 U10967 ( .A(\I_cache/cache[6][114] ), .B(n9772), .S0(n5886), .Y(
        n11927) );
  CLKMX2X2 U10968 ( .A(\I_cache/cache[5][114] ), .B(n9772), .S0(n5752), .Y(
        n11928) );
  CLKMX2X2 U10969 ( .A(\I_cache/cache[4][114] ), .B(n9772), .S0(n5799), .Y(
        n11929) );
  CLKMX2X2 U10970 ( .A(\I_cache/cache[3][114] ), .B(n9772), .S0(n5664), .Y(
        n11930) );
  CLKMX2X2 U10971 ( .A(\I_cache/cache[2][114] ), .B(n9772), .S0(n5708), .Y(
        n11931) );
  CLKMX2X2 U10972 ( .A(\I_cache/cache[1][114] ), .B(n9772), .S0(n5580), .Y(
        n11932) );
  CLKMX2X2 U10973 ( .A(\I_cache/cache[0][114] ), .B(n9772), .S0(n5618), .Y(
        n11933) );
  CLKMX2X2 U10974 ( .A(\I_cache/cache[7][113] ), .B(n9740), .S0(n5842), .Y(
        n11934) );
  CLKMX2X2 U10975 ( .A(\I_cache/cache[5][113] ), .B(n9740), .S0(n5755), .Y(
        n11936) );
  CLKMX2X2 U10976 ( .A(\I_cache/cache[4][113] ), .B(n9740), .S0(n5798), .Y(
        n11937) );
  CLKMX2X2 U10977 ( .A(\I_cache/cache[3][113] ), .B(n9740), .S0(n5663), .Y(
        n11938) );
  CLKMX2X2 U10978 ( .A(\I_cache/cache[2][113] ), .B(n9740), .S0(n5708), .Y(
        n11939) );
  CLKMX2X2 U10979 ( .A(\I_cache/cache[0][113] ), .B(n9740), .S0(n5617), .Y(
        n11941) );
  CLKMX2X2 U10980 ( .A(\I_cache/cache[7][112] ), .B(n9762), .S0(n5843), .Y(
        n11942) );
  CLKMX2X2 U10981 ( .A(\I_cache/cache[6][112] ), .B(n9762), .S0(n5886), .Y(
        n11943) );
  CLKMX2X2 U10982 ( .A(\I_cache/cache[5][112] ), .B(n9762), .S0(n5752), .Y(
        n11944) );
  CLKMX2X2 U10983 ( .A(\I_cache/cache[4][112] ), .B(n9762), .S0(n5799), .Y(
        n11945) );
  CLKMX2X2 U10984 ( .A(\I_cache/cache[3][112] ), .B(n9762), .S0(n5664), .Y(
        n11946) );
  CLKMX2X2 U10985 ( .A(\I_cache/cache[2][112] ), .B(n9762), .S0(n5710), .Y(
        n11947) );
  CLKMX2X2 U10986 ( .A(\I_cache/cache[1][112] ), .B(n9762), .S0(n5577), .Y(
        n11948) );
  CLKMX2X2 U10987 ( .A(\I_cache/cache[0][112] ), .B(n9762), .S0(n5618), .Y(
        n11949) );
  CLKMX2X2 U10988 ( .A(\I_cache/cache[7][111] ), .B(n10067), .S0(n5844), .Y(
        n11950) );
  CLKMX2X2 U10989 ( .A(\I_cache/cache[6][111] ), .B(n10067), .S0(n5888), .Y(
        n11951) );
  CLKMX2X2 U10990 ( .A(\I_cache/cache[5][111] ), .B(n10067), .S0(n5754), .Y(
        n11952) );
  CLKMX2X2 U10991 ( .A(\I_cache/cache[4][111] ), .B(n10067), .S0(n5800), .Y(
        n11953) );
  CLKMX2X2 U10992 ( .A(\I_cache/cache[3][111] ), .B(n10067), .S0(n5665), .Y(
        n11954) );
  CLKMX2X2 U10993 ( .A(\I_cache/cache[2][111] ), .B(n10067), .S0(n5710), .Y(
        n11955) );
  CLKMX2X2 U10994 ( .A(\I_cache/cache[1][111] ), .B(n10067), .S0(n5575), .Y(
        n11956) );
  CLKMX2X2 U10995 ( .A(\I_cache/cache[0][111] ), .B(n10067), .S0(n5621), .Y(
        n11957) );
  CLKMX2X2 U10996 ( .A(\I_cache/cache[7][110] ), .B(n10246), .S0(n5850), .Y(
        n11958) );
  CLKMX2X2 U10997 ( .A(\I_cache/cache[6][110] ), .B(n10246), .S0(n5893), .Y(
        n11959) );
  CLKMX2X2 U10998 ( .A(\I_cache/cache[5][110] ), .B(n10246), .S0(n5759), .Y(
        n11960) );
  CLKMX2X2 U10999 ( .A(\I_cache/cache[4][110] ), .B(n10246), .S0(n5806), .Y(
        n11961) );
  CLKMX2X2 U11000 ( .A(\I_cache/cache[3][110] ), .B(n10246), .S0(n5671), .Y(
        n11962) );
  CLKMX2X2 U11001 ( .A(\I_cache/cache[2][110] ), .B(n10246), .S0(n5716), .Y(
        n11963) );
  CLKMX2X2 U11002 ( .A(\I_cache/cache[1][110] ), .B(n10246), .S0(n5582), .Y(
        n11964) );
  CLKMX2X2 U11003 ( .A(\I_cache/cache[0][110] ), .B(n10246), .S0(n5625), .Y(
        n11965) );
  CLKMX2X2 U11004 ( .A(\I_cache/cache[7][109] ), .B(n10224), .S0(n5845), .Y(
        n11966) );
  CLKMX2X2 U11005 ( .A(\I_cache/cache[6][109] ), .B(n10224), .S0(n5889), .Y(
        n11967) );
  CLKMX2X2 U11006 ( .A(\I_cache/cache[5][109] ), .B(n10224), .S0(n5755), .Y(
        n11968) );
  CLKMX2X2 U11007 ( .A(\I_cache/cache[4][109] ), .B(n10224), .S0(n5801), .Y(
        n11969) );
  CLKMX2X2 U11008 ( .A(\I_cache/cache[3][109] ), .B(n10224), .S0(n5666), .Y(
        n11970) );
  CLKMX2X2 U11009 ( .A(\I_cache/cache[2][109] ), .B(n10224), .S0(n5711), .Y(
        n11971) );
  CLKMX2X2 U11010 ( .A(\I_cache/cache[1][109] ), .B(n10224), .S0(n5577), .Y(
        n11972) );
  CLKMX2X2 U11011 ( .A(\I_cache/cache[0][109] ), .B(n10224), .S0(n5619), .Y(
        n11973) );
  CLKMX2X2 U11012 ( .A(\I_cache/cache[7][108] ), .B(n10126), .S0(n5845), .Y(
        n11974) );
  CLKMX2X2 U11013 ( .A(\I_cache/cache[6][108] ), .B(n10126), .S0(n5889), .Y(
        n11975) );
  CLKMX2X2 U11014 ( .A(\I_cache/cache[5][108] ), .B(n10126), .S0(n5755), .Y(
        n11976) );
  CLKMX2X2 U11015 ( .A(\I_cache/cache[4][108] ), .B(n10126), .S0(n5801), .Y(
        n11977) );
  CLKMX2X2 U11016 ( .A(\I_cache/cache[3][108] ), .B(n10126), .S0(n5666), .Y(
        n11978) );
  CLKMX2X2 U11017 ( .A(\I_cache/cache[2][108] ), .B(n10126), .S0(n5711), .Y(
        n11979) );
  CLKMX2X2 U11018 ( .A(\I_cache/cache[1][108] ), .B(n10126), .S0(n5577), .Y(
        n11980) );
  CLKMX2X2 U11019 ( .A(\I_cache/cache[0][108] ), .B(n10126), .S0(n5620), .Y(
        n11981) );
  CLKMX2X2 U11020 ( .A(\I_cache/cache[7][107] ), .B(n10090), .S0(n5845), .Y(
        n11982) );
  CLKMX2X2 U11021 ( .A(\I_cache/cache[6][107] ), .B(n10090), .S0(n5889), .Y(
        n11983) );
  CLKMX2X2 U11022 ( .A(\I_cache/cache[5][107] ), .B(n10090), .S0(n5755), .Y(
        n11984) );
  CLKMX2X2 U11023 ( .A(\I_cache/cache[4][107] ), .B(n10090), .S0(n5801), .Y(
        n11985) );
  CLKMX2X2 U11024 ( .A(\I_cache/cache[3][107] ), .B(n10090), .S0(n5666), .Y(
        n11986) );
  CLKMX2X2 U11025 ( .A(\I_cache/cache[2][107] ), .B(n10090), .S0(n5711), .Y(
        n11987) );
  CLKMX2X2 U11026 ( .A(\I_cache/cache[1][107] ), .B(n10090), .S0(n5577), .Y(
        n11988) );
  CLKMX2X2 U11027 ( .A(\I_cache/cache[0][107] ), .B(n10090), .S0(n5620), .Y(
        n11989) );
  CLKMX2X2 U11028 ( .A(\I_cache/cache[7][106] ), .B(n9839), .S0(n5843), .Y(
        n11990) );
  CLKMX2X2 U11029 ( .A(\I_cache/cache[6][106] ), .B(n9839), .S0(n5886), .Y(
        n11991) );
  CLKMX2X2 U11030 ( .A(\I_cache/cache[5][106] ), .B(n9839), .S0(n5752), .Y(
        n11992) );
  CLKMX2X2 U11031 ( .A(\I_cache/cache[4][106] ), .B(n9839), .S0(n5799), .Y(
        n11993) );
  CLKMX2X2 U11032 ( .A(\I_cache/cache[3][106] ), .B(n9839), .S0(n5664), .Y(
        n11994) );
  CLKMX2X2 U11033 ( .A(\I_cache/cache[2][106] ), .B(n9839), .S0(n5712), .Y(
        n11995) );
  CLKMX2X2 U11034 ( .A(\I_cache/cache[1][106] ), .B(n9839), .S0(n5578), .Y(
        n11996) );
  CLKMX2X2 U11035 ( .A(\I_cache/cache[0][106] ), .B(n9839), .S0(n5621), .Y(
        n11997) );
  CLKMX2X2 U11036 ( .A(\I_cache/cache[7][105] ), .B(n9883), .S0(n5846), .Y(
        n11998) );
  CLKMX2X2 U11037 ( .A(\I_cache/cache[6][105] ), .B(n9883), .S0(n5890), .Y(
        n11999) );
  CLKMX2X2 U11038 ( .A(\I_cache/cache[5][105] ), .B(n9883), .S0(n5756), .Y(
        n12000) );
  CLKMX2X2 U11039 ( .A(\I_cache/cache[4][105] ), .B(n9883), .S0(n5802), .Y(
        n12001) );
  CLKMX2X2 U11040 ( .A(\I_cache/cache[3][105] ), .B(n9883), .S0(n5667), .Y(
        n12002) );
  CLKMX2X2 U11041 ( .A(\I_cache/cache[2][105] ), .B(n9883), .S0(n5712), .Y(
        n12003) );
  CLKMX2X2 U11042 ( .A(\I_cache/cache[1][105] ), .B(n9883), .S0(n5578), .Y(
        n12004) );
  CLKMX2X2 U11043 ( .A(\I_cache/cache[0][105] ), .B(n9883), .S0(n5621), .Y(
        n12005) );
  CLKMX2X2 U11044 ( .A(\I_cache/cache[7][104] ), .B(n9861), .S0(n5846), .Y(
        n12006) );
  CLKMX2X2 U11045 ( .A(\I_cache/cache[6][104] ), .B(n9861), .S0(n5888), .Y(
        n12007) );
  CLKMX2X2 U11046 ( .A(\I_cache/cache[5][104] ), .B(n9861), .S0(n5756), .Y(
        n12008) );
  CLKMX2X2 U11047 ( .A(\I_cache/cache[4][104] ), .B(n9861), .S0(n5802), .Y(
        n12009) );
  CLKMX2X2 U11048 ( .A(\I_cache/cache[3][104] ), .B(n9861), .S0(n5667), .Y(
        n12010) );
  CLKMX2X2 U11049 ( .A(\I_cache/cache[2][104] ), .B(n9861), .S0(n5712), .Y(
        n12011) );
  CLKMX2X2 U11050 ( .A(\I_cache/cache[1][104] ), .B(n9861), .S0(n5578), .Y(
        n12012) );
  CLKMX2X2 U11051 ( .A(\I_cache/cache[0][104] ), .B(n9861), .S0(n5621), .Y(
        n12013) );
  CLKMX2X2 U11052 ( .A(\I_cache/cache[7][103] ), .B(n9905), .S0(n5846), .Y(
        n12014) );
  CLKMX2X2 U11053 ( .A(\I_cache/cache[6][103] ), .B(n9905), .S0(n5886), .Y(
        n12015) );
  CLKMX2X2 U11054 ( .A(\I_cache/cache[5][103] ), .B(n9905), .S0(n5756), .Y(
        n12016) );
  CLKMX2X2 U11055 ( .A(\I_cache/cache[4][103] ), .B(n9905), .S0(n5802), .Y(
        n12017) );
  CLKMX2X2 U11056 ( .A(\I_cache/cache[3][103] ), .B(n9905), .S0(n5667), .Y(
        n12018) );
  CLKMX2X2 U11057 ( .A(\I_cache/cache[2][103] ), .B(n9905), .S0(n5712), .Y(
        n12019) );
  CLKMX2X2 U11058 ( .A(\I_cache/cache[1][103] ), .B(n9905), .S0(n5577), .Y(
        n12020) );
  CLKMX2X2 U11059 ( .A(\I_cache/cache[0][103] ), .B(n9905), .S0(n5622), .Y(
        n12021) );
  CLKMX2X2 U11060 ( .A(\I_cache/cache[7][102] ), .B(n9927), .S0(n5847), .Y(
        n12022) );
  CLKMX2X2 U11061 ( .A(\I_cache/cache[6][102] ), .B(n9927), .S0(n5890), .Y(
        n12023) );
  CLKMX2X2 U11062 ( .A(\I_cache/cache[5][102] ), .B(n9927), .S0(n5757), .Y(
        n12024) );
  CLKMX2X2 U11063 ( .A(\I_cache/cache[4][102] ), .B(n9927), .S0(n5803), .Y(
        n12025) );
  CLKMX2X2 U11064 ( .A(\I_cache/cache[3][102] ), .B(n9927), .S0(n5668), .Y(
        n12026) );
  CLKMX2X2 U11065 ( .A(\I_cache/cache[2][102] ), .B(n9927), .S0(n5713), .Y(
        n12027) );
  CLKMX2X2 U11066 ( .A(\I_cache/cache[1][102] ), .B(n9927), .S0(n5579), .Y(
        n12028) );
  CLKMX2X2 U11067 ( .A(\I_cache/cache[0][102] ), .B(n9927), .S0(n5622), .Y(
        n12029) );
  CLKMX2X2 U11068 ( .A(\I_cache/cache[7][101] ), .B(n9720), .S0(n5842), .Y(
        n12030) );
  CLKMX2X2 U11069 ( .A(\I_cache/cache[6][101] ), .B(n9720), .S0(n5885), .Y(
        n12031) );
  CLKMX2X2 U11070 ( .A(\I_cache/cache[5][101] ), .B(n9720), .S0(n5757), .Y(
        n12032) );
  CLKMX2X2 U11071 ( .A(\I_cache/cache[4][101] ), .B(n9720), .S0(n5798), .Y(
        n12033) );
  CLKMX2X2 U11072 ( .A(\I_cache/cache[3][101] ), .B(n9720), .S0(n5663), .Y(
        n12034) );
  CLKMX2X2 U11073 ( .A(\I_cache/cache[2][101] ), .B(n9720), .S0(n5708), .Y(
        n12035) );
  CLKMX2X2 U11074 ( .A(\I_cache/cache[1][101] ), .B(n9720), .S0(n5574), .Y(
        n12036) );
  CLKMX2X2 U11075 ( .A(\I_cache/cache[0][101] ), .B(n9720), .S0(n5617), .Y(
        n12037) );
  CLKMX2X2 U11076 ( .A(\I_cache/cache[7][100] ), .B(n10860), .S0(n5850), .Y(
        n12038) );
  CLKMX2X2 U11077 ( .A(\I_cache/cache[6][100] ), .B(n10860), .S0(n5893), .Y(
        n12039) );
  CLKMX2X2 U11078 ( .A(\I_cache/cache[5][100] ), .B(n10860), .S0(n5759), .Y(
        n12040) );
  CLKMX2X2 U11079 ( .A(\I_cache/cache[4][100] ), .B(n10860), .S0(n5806), .Y(
        n12041) );
  CLKMX2X2 U11080 ( .A(\I_cache/cache[3][100] ), .B(n10860), .S0(n5671), .Y(
        n12042) );
  CLKMX2X2 U11081 ( .A(\I_cache/cache[2][100] ), .B(n10860), .S0(n5716), .Y(
        n12043) );
  CLKMX2X2 U11082 ( .A(\I_cache/cache[1][100] ), .B(n10860), .S0(n5582), .Y(
        n12044) );
  CLKMX2X2 U11083 ( .A(\I_cache/cache[0][100] ), .B(n10860), .S0(n5625), .Y(
        n12045) );
  CLKMX2X2 U11084 ( .A(\I_cache/cache[7][99] ), .B(n10954), .S0(n5842), .Y(
        n12046) );
  CLKMX2X2 U11085 ( .A(\I_cache/cache[6][99] ), .B(n10954), .S0(n5890), .Y(
        n12047) );
  CLKMX2X2 U11086 ( .A(\I_cache/cache[5][99] ), .B(n10954), .S0(n4831), .Y(
        n12048) );
  CLKMX2X2 U11087 ( .A(\I_cache/cache[4][99] ), .B(n10954), .S0(n5803), .Y(
        n12049) );
  CLKMX2X2 U11088 ( .A(\I_cache/cache[3][99] ), .B(n10954), .S0(n5668), .Y(
        n12050) );
  CLKMX2X2 U11089 ( .A(\I_cache/cache[2][99] ), .B(n10954), .S0(n5712), .Y(
        n12051) );
  CLKMX2X2 U11090 ( .A(\I_cache/cache[1][99] ), .B(n10954), .S0(n5582), .Y(
        n12052) );
  CLKMX2X2 U11091 ( .A(\I_cache/cache[0][99] ), .B(n10954), .S0(n5624), .Y(
        n12053) );
  CLKMX2X2 U11092 ( .A(\I_cache/cache[7][98] ), .B(n10925), .S0(n5843), .Y(
        n12054) );
  CLKMX2X2 U11093 ( .A(\I_cache/cache[6][98] ), .B(n10925), .S0(n5889), .Y(
        n12055) );
  CLKMX2X2 U11094 ( .A(\I_cache/cache[5][98] ), .B(n10925), .S0(n4830), .Y(
        n12056) );
  CLKMX2X2 U11095 ( .A(\I_cache/cache[4][98] ), .B(n10925), .S0(n5801), .Y(
        n12057) );
  CLKMX2X2 U11096 ( .A(\I_cache/cache[3][98] ), .B(n10925), .S0(n5665), .Y(
        n12058) );
  CLKMX2X2 U11097 ( .A(\I_cache/cache[2][98] ), .B(n10925), .S0(n5713), .Y(
        n12059) );
  CLKMX2X2 U11098 ( .A(\I_cache/cache[1][98] ), .B(n10925), .S0(n5576), .Y(
        n12060) );
  CLKMX2X2 U11099 ( .A(\I_cache/cache[0][98] ), .B(n10925), .S0(n5625), .Y(
        n12061) );
  CLKMX2X2 U11100 ( .A(\I_cache/cache[6][97] ), .B(n10883), .S0(n5892), .Y(
        n12063) );
  CLKMX2X2 U11101 ( .A(\I_cache/cache[5][97] ), .B(n10883), .S0(n5757), .Y(
        n12064) );
  CLKMX2X2 U11102 ( .A(\I_cache/cache[4][97] ), .B(n10883), .S0(n5805), .Y(
        n12065) );
  CLKMX2X2 U11103 ( .A(\I_cache/cache[3][97] ), .B(n10883), .S0(n5670), .Y(
        n12066) );
  CLKMX2X2 U11104 ( .A(\I_cache/cache[2][97] ), .B(n10883), .S0(n5715), .Y(
        n12067) );
  CLKMX2X2 U11105 ( .A(\I_cache/cache[1][97] ), .B(n10883), .S0(n5581), .Y(
        n12068) );
  CLKMX2X2 U11106 ( .A(\I_cache/cache[0][97] ), .B(n10883), .S0(n5617), .Y(
        n12069) );
  CLKMX2X2 U11107 ( .A(\I_cache/cache[7][96] ), .B(n10817), .S0(n5850), .Y(
        n12070) );
  CLKMX2X2 U11108 ( .A(\I_cache/cache[6][96] ), .B(n10817), .S0(n5893), .Y(
        n12071) );
  CLKMX2X2 U11109 ( .A(\I_cache/cache[5][96] ), .B(n10817), .S0(n5759), .Y(
        n12072) );
  CLKMX2X2 U11110 ( .A(\I_cache/cache[4][96] ), .B(n10817), .S0(n5806), .Y(
        n12073) );
  CLKMX2X2 U11111 ( .A(\I_cache/cache[3][96] ), .B(n10817), .S0(n5671), .Y(
        n12074) );
  CLKMX2X2 U11112 ( .A(\I_cache/cache[2][96] ), .B(n10817), .S0(n5716), .Y(
        n12075) );
  CLKMX2X2 U11113 ( .A(\I_cache/cache[1][96] ), .B(n10817), .S0(n5582), .Y(
        n12076) );
  CLKMX2X2 U11114 ( .A(\I_cache/cache[0][96] ), .B(n10817), .S0(n5625), .Y(
        n12077) );
  CLKMX2X2 U11115 ( .A(\I_cache/cache[7][31] ), .B(n9659), .S0(n5848), .Y(
        n12590) );
  CLKMX2X2 U11116 ( .A(\I_cache/cache[6][31] ), .B(n9659), .S0(n5887), .Y(
        n12591) );
  CLKMX2X2 U11117 ( .A(\I_cache/cache[5][31] ), .B(n9659), .S0(n5753), .Y(
        n12592) );
  CLKMX2X2 U11118 ( .A(\I_cache/cache[4][31] ), .B(n9659), .S0(n5798), .Y(
        n12593) );
  CLKMX2X2 U11119 ( .A(\I_cache/cache[3][31] ), .B(n9659), .S0(n5668), .Y(
        n12594) );
  CLKMX2X2 U11120 ( .A(\I_cache/cache[2][31] ), .B(n9659), .S0(n5709), .Y(
        n12595) );
  CLKMX2X2 U11121 ( .A(\I_cache/cache[1][31] ), .B(n9659), .S0(n5575), .Y(
        n12596) );
  CLKMX2X2 U11122 ( .A(\I_cache/cache[0][31] ), .B(n9659), .S0(n5619), .Y(
        n12597) );
  CLKMX2X2 U11123 ( .A(\I_cache/cache[7][30] ), .B(n9681), .S0(n5842), .Y(
        n12598) );
  CLKMX2X2 U11124 ( .A(\I_cache/cache[6][30] ), .B(n9681), .S0(n5885), .Y(
        n12599) );
  CLKMX2X2 U11125 ( .A(\I_cache/cache[5][30] ), .B(n9681), .S0(n5752), .Y(
        n12600) );
  CLKMX2X2 U11126 ( .A(\I_cache/cache[4][30] ), .B(n9681), .S0(n5798), .Y(
        n12601) );
  CLKMX2X2 U11127 ( .A(\I_cache/cache[3][30] ), .B(n9681), .S0(n5663), .Y(
        n12602) );
  CLKMX2X2 U11128 ( .A(\I_cache/cache[2][30] ), .B(n9681), .S0(n5708), .Y(
        n12603) );
  CLKMX2X2 U11129 ( .A(\I_cache/cache[1][30] ), .B(n9681), .S0(n5574), .Y(
        n12604) );
  CLKMX2X2 U11130 ( .A(\I_cache/cache[0][30] ), .B(n9681), .S0(n5617), .Y(
        n12605) );
  CLKMX2X2 U11131 ( .A(\I_cache/cache[7][29] ), .B(n9703), .S0(n5842), .Y(
        n12606) );
  CLKMX2X2 U11132 ( .A(\I_cache/cache[6][29] ), .B(n9703), .S0(n5885), .Y(
        n12607) );
  CLKMX2X2 U11133 ( .A(\I_cache/cache[5][29] ), .B(n9703), .S0(n5753), .Y(
        n12608) );
  CLKMX2X2 U11134 ( .A(\I_cache/cache[4][29] ), .B(n9703), .S0(n5798), .Y(
        n12609) );
  CLKMX2X2 U11135 ( .A(\I_cache/cache[3][29] ), .B(n9703), .S0(n5663), .Y(
        n12610) );
  CLKMX2X2 U11136 ( .A(\I_cache/cache[2][29] ), .B(n9703), .S0(n5708), .Y(
        n12611) );
  CLKMX2X2 U11137 ( .A(\I_cache/cache[1][29] ), .B(n9703), .S0(n5574), .Y(
        n12612) );
  CLKMX2X2 U11138 ( .A(\I_cache/cache[0][29] ), .B(n9703), .S0(n5617), .Y(
        n12613) );
  CLKMX2X2 U11139 ( .A(\I_cache/cache[7][28] ), .B(n9651), .S0(n5845), .Y(
        n12614) );
  CLKMX2X2 U11140 ( .A(\I_cache/cache[6][28] ), .B(n9651), .S0(n5887), .Y(
        n12615) );
  CLKMX2X2 U11141 ( .A(\I_cache/cache[5][28] ), .B(n9651), .S0(n5753), .Y(
        n12616) );
  CLKMX2X2 U11142 ( .A(\I_cache/cache[4][28] ), .B(n9651), .S0(n5803), .Y(
        n12617) );
  CLKMX2X2 U11143 ( .A(\I_cache/cache[3][28] ), .B(n9651), .S0(n5664), .Y(
        n12618) );
  CLKMX2X2 U11144 ( .A(\I_cache/cache[2][28] ), .B(n9651), .S0(n5709), .Y(
        n12619) );
  CLKMX2X2 U11145 ( .A(\I_cache/cache[1][28] ), .B(n9651), .S0(n5575), .Y(
        n12620) );
  CLKMX2X2 U11146 ( .A(\I_cache/cache[0][28] ), .B(n9651), .S0(n5622), .Y(
        n12621) );
  CLKMX2X2 U11147 ( .A(\I_cache/cache[7][27] ), .B(n9629), .S0(n5844), .Y(
        n12622) );
  CLKMX2X2 U11148 ( .A(\I_cache/cache[6][27] ), .B(n9629), .S0(n5887), .Y(
        n12623) );
  CLKMX2X2 U11149 ( .A(\I_cache/cache[5][27] ), .B(n9629), .S0(n5753), .Y(
        n12624) );
  CLKMX2X2 U11150 ( .A(\I_cache/cache[4][27] ), .B(n9629), .S0(n5801), .Y(
        n12625) );
  CLKMX2X2 U11151 ( .A(\I_cache/cache[3][27] ), .B(n9629), .S0(n5666), .Y(
        n12626) );
  CLKMX2X2 U11152 ( .A(\I_cache/cache[2][27] ), .B(n9629), .S0(n5709), .Y(
        n12627) );
  CLKMX2X2 U11153 ( .A(\I_cache/cache[1][27] ), .B(n9629), .S0(n5575), .Y(
        n12628) );
  CLKMX2X2 U11154 ( .A(\I_cache/cache[0][27] ), .B(n9629), .S0(n5617), .Y(
        n12629) );
  CLKMX2X2 U11155 ( .A(\I_cache/cache[7][26] ), .B(n6607), .S0(n5846), .Y(
        n12630) );
  CLKMX2X2 U11156 ( .A(\I_cache/cache[6][26] ), .B(n6607), .S0(n5886), .Y(
        n12631) );
  CLKMX2X2 U11157 ( .A(\I_cache/cache[5][26] ), .B(n6607), .S0(n5757), .Y(
        n12632) );
  CLKMX2X2 U11158 ( .A(\I_cache/cache[4][26] ), .B(n6607), .S0(n5802), .Y(
        n12633) );
  CLKMX2X2 U11159 ( .A(\I_cache/cache[3][26] ), .B(n6607), .S0(n5668), .Y(
        n12634) );
  CLKMX2X2 U11160 ( .A(\I_cache/cache[2][26] ), .B(n6607), .S0(n5708), .Y(
        n12635) );
  CLKMX2X2 U11161 ( .A(\I_cache/cache[1][26] ), .B(n6607), .S0(n5575), .Y(
        n12636) );
  CLKMX2X2 U11162 ( .A(\I_cache/cache[0][26] ), .B(n6607), .S0(n5618), .Y(
        n12637) );
  CLKMX2X2 U11163 ( .A(\I_cache/cache[7][25] ), .B(n10048), .S0(n5844), .Y(
        n12638) );
  CLKMX2X2 U11164 ( .A(\I_cache/cache[6][25] ), .B(n10048), .S0(n5888), .Y(
        n12639) );
  CLKMX2X2 U11165 ( .A(\I_cache/cache[5][25] ), .B(n10048), .S0(n5754), .Y(
        n12640) );
  CLKMX2X2 U11166 ( .A(\I_cache/cache[4][25] ), .B(n10048), .S0(n5800), .Y(
        n12641) );
  CLKMX2X2 U11167 ( .A(\I_cache/cache[3][25] ), .B(n10048), .S0(n5665), .Y(
        n12642) );
  CLKMX2X2 U11168 ( .A(\I_cache/cache[2][25] ), .B(n10048), .S0(n5710), .Y(
        n12643) );
  CLKMX2X2 U11169 ( .A(\I_cache/cache[1][25] ), .B(n10048), .S0(n5576), .Y(
        n12644) );
  CLKMX2X2 U11170 ( .A(\I_cache/cache[0][25] ), .B(n10048), .S0(n5619), .Y(
        n12645) );
  CLKMX2X2 U11171 ( .A(\I_cache/cache[7][24] ), .B(n10843), .S0(n5850), .Y(
        n12646) );
  CLKMX2X2 U11172 ( .A(\I_cache/cache[6][24] ), .B(n10843), .S0(n5893), .Y(
        n12647) );
  CLKMX2X2 U11173 ( .A(\I_cache/cache[5][24] ), .B(n10843), .S0(n5759), .Y(
        n12648) );
  CLKMX2X2 U11174 ( .A(\I_cache/cache[4][24] ), .B(n10843), .S0(n5806), .Y(
        n12649) );
  CLKMX2X2 U11175 ( .A(\I_cache/cache[3][24] ), .B(n10843), .S0(n5671), .Y(
        n12650) );
  CLKMX2X2 U11176 ( .A(\I_cache/cache[2][24] ), .B(n10843), .S0(n5716), .Y(
        n12651) );
  CLKMX2X2 U11177 ( .A(\I_cache/cache[1][24] ), .B(n10843), .S0(n5582), .Y(
        n12652) );
  CLKMX2X2 U11178 ( .A(\I_cache/cache[0][24] ), .B(n10843), .S0(n5625), .Y(
        n12653) );
  CLKMX2X2 U11179 ( .A(\I_cache/cache[7][23] ), .B(n10026), .S0(n5844), .Y(
        n12654) );
  CLKMX2X2 U11180 ( .A(\I_cache/cache[6][23] ), .B(n10026), .S0(n5888), .Y(
        n12655) );
  CLKMX2X2 U11181 ( .A(\I_cache/cache[5][23] ), .B(n10026), .S0(n5754), .Y(
        n12656) );
  CLKMX2X2 U11182 ( .A(\I_cache/cache[4][23] ), .B(n10026), .S0(n5800), .Y(
        n12657) );
  CLKMX2X2 U11183 ( .A(\I_cache/cache[3][23] ), .B(n10026), .S0(n5665), .Y(
        n12658) );
  CLKMX2X2 U11184 ( .A(\I_cache/cache[2][23] ), .B(n10026), .S0(n5710), .Y(
        n12659) );
  CLKMX2X2 U11185 ( .A(\I_cache/cache[1][23] ), .B(n10026), .S0(n5576), .Y(
        n12660) );
  CLKMX2X2 U11186 ( .A(\I_cache/cache[0][23] ), .B(n10026), .S0(n5619), .Y(
        n12661) );
  CLKMX2X2 U11187 ( .A(\I_cache/cache[7][22] ), .B(n9982), .S0(n5847), .Y(
        n12662) );
  CLKMX2X2 U11188 ( .A(\I_cache/cache[6][22] ), .B(n9982), .S0(n5890), .Y(
        n12663) );
  CLKMX2X2 U11189 ( .A(\I_cache/cache[5][22] ), .B(n9982), .S0(n5757), .Y(
        n12664) );
  CLKMX2X2 U11190 ( .A(\I_cache/cache[4][22] ), .B(n9982), .S0(n5803), .Y(
        n12665) );
  CLKMX2X2 U11191 ( .A(\I_cache/cache[3][22] ), .B(n9982), .S0(n5668), .Y(
        n12666) );
  CLKMX2X2 U11192 ( .A(\I_cache/cache[2][22] ), .B(n9982), .S0(n5713), .Y(
        n12667) );
  CLKMX2X2 U11193 ( .A(\I_cache/cache[1][22] ), .B(n9982), .S0(n5579), .Y(
        n12668) );
  CLKMX2X2 U11194 ( .A(\I_cache/cache[0][22] ), .B(n9982), .S0(n5622), .Y(
        n12669) );
  CLKMX2X2 U11195 ( .A(\I_cache/cache[7][21] ), .B(n10004), .S0(n5847), .Y(
        n12670) );
  CLKMX2X2 U11196 ( .A(\I_cache/cache[6][21] ), .B(n10004), .S0(n5890), .Y(
        n12671) );
  CLKMX2X2 U11197 ( .A(\I_cache/cache[5][21] ), .B(n10004), .S0(n5757), .Y(
        n12672) );
  CLKMX2X2 U11198 ( .A(\I_cache/cache[4][21] ), .B(n10004), .S0(n5803), .Y(
        n12673) );
  CLKMX2X2 U11199 ( .A(\I_cache/cache[3][21] ), .B(n10004), .S0(n5668), .Y(
        n12674) );
  CLKMX2X2 U11200 ( .A(\I_cache/cache[2][21] ), .B(n10004), .S0(n5713), .Y(
        n12675) );
  CLKMX2X2 U11201 ( .A(\I_cache/cache[1][21] ), .B(n10004), .S0(n5578), .Y(
        n12676) );
  CLKMX2X2 U11202 ( .A(\I_cache/cache[0][21] ), .B(n10004), .S0(n5619), .Y(
        n12677) );
  CLKMX2X2 U11203 ( .A(\I_cache/cache[7][20] ), .B(n9793), .S0(n5843), .Y(
        n12678) );
  CLKMX2X2 U11204 ( .A(\I_cache/cache[6][20] ), .B(n9793), .S0(n5886), .Y(
        n12679) );
  CLKMX2X2 U11205 ( .A(\I_cache/cache[5][20] ), .B(n9793), .S0(n5752), .Y(
        n12680) );
  CLKMX2X2 U11206 ( .A(\I_cache/cache[4][20] ), .B(n9793), .S0(n5799), .Y(
        n12681) );
  CLKMX2X2 U11207 ( .A(\I_cache/cache[3][20] ), .B(n9793), .S0(n5664), .Y(
        n12682) );
  CLKMX2X2 U11208 ( .A(\I_cache/cache[2][20] ), .B(n9793), .S0(n5713), .Y(
        n12683) );
  CLKMX2X2 U11209 ( .A(\I_cache/cache[1][20] ), .B(n9793), .S0(n5579), .Y(
        n12684) );
  CLKMX2X2 U11210 ( .A(\I_cache/cache[0][20] ), .B(n9793), .S0(n5618), .Y(
        n12685) );
  CLKMX2X2 U11211 ( .A(\I_cache/cache[7][19] ), .B(n11092), .S0(n5848), .Y(
        n12686) );
  CLKMX2X2 U11212 ( .A(\I_cache/cache[6][19] ), .B(n11092), .S0(n5891), .Y(
        n12687) );
  CLKMX2X2 U11213 ( .A(\I_cache/cache[5][19] ), .B(n11092), .S0(n5758), .Y(
        n12688) );
  CLKMX2X2 U11214 ( .A(\I_cache/cache[4][19] ), .B(n11092), .S0(n5804), .Y(
        n12689) );
  CLKMX2X2 U11215 ( .A(\I_cache/cache[3][19] ), .B(n11092), .S0(n5669), .Y(
        n12690) );
  CLKMX2X2 U11216 ( .A(\I_cache/cache[2][19] ), .B(n11092), .S0(n5714), .Y(
        n12691) );
  CLKMX2X2 U11217 ( .A(\I_cache/cache[1][19] ), .B(n11092), .S0(n5580), .Y(
        n12692) );
  CLKMX2X2 U11218 ( .A(\I_cache/cache[0][19] ), .B(n11092), .S0(n5623), .Y(
        n12693) );
  CLKMX2X2 U11219 ( .A(\I_cache/cache[7][18] ), .B(n9773), .S0(n5843), .Y(
        n12694) );
  CLKMX2X2 U11220 ( .A(\I_cache/cache[6][18] ), .B(n9773), .S0(n5886), .Y(
        n12695) );
  CLKMX2X2 U11221 ( .A(\I_cache/cache[5][18] ), .B(n9773), .S0(n5752), .Y(
        n12696) );
  CLKMX2X2 U11222 ( .A(\I_cache/cache[4][18] ), .B(n9773), .S0(n5799), .Y(
        n12697) );
  CLKMX2X2 U11223 ( .A(\I_cache/cache[3][18] ), .B(n9773), .S0(n5664), .Y(
        n12698) );
  CLKMX2X2 U11224 ( .A(\I_cache/cache[2][18] ), .B(n9773), .S0(n5711), .Y(
        n12699) );
  CLKMX2X2 U11225 ( .A(\I_cache/cache[1][18] ), .B(n9773), .S0(n5582), .Y(
        n12700) );
  CLKMX2X2 U11226 ( .A(\I_cache/cache[0][18] ), .B(n9773), .S0(n5618), .Y(
        n12701) );
  CLKMX2X2 U11227 ( .A(\I_cache/cache[7][17] ), .B(n9745), .S0(n5842), .Y(
        n12702) );
  CLKMX2X2 U11228 ( .A(\I_cache/cache[6][17] ), .B(n9745), .S0(n5885), .Y(
        n12703) );
  CLKMX2X2 U11229 ( .A(\I_cache/cache[5][17] ), .B(n9745), .S0(n5754), .Y(
        n12704) );
  CLKMX2X2 U11230 ( .A(\I_cache/cache[4][17] ), .B(n9745), .S0(n5798), .Y(
        n12705) );
  CLKMX2X2 U11231 ( .A(\I_cache/cache[3][17] ), .B(n9745), .S0(n5663), .Y(
        n12706) );
  CLKMX2X2 U11232 ( .A(\I_cache/cache[2][17] ), .B(n9745), .S0(n5708), .Y(
        n12707) );
  CLKMX2X2 U11233 ( .A(\I_cache/cache[1][17] ), .B(n9745), .S0(n5574), .Y(
        n12708) );
  CLKMX2X2 U11234 ( .A(\I_cache/cache[0][17] ), .B(n9745), .S0(n5620), .Y(
        n12709) );
  CLKMX2X2 U11235 ( .A(\I_cache/cache[7][16] ), .B(n9767), .S0(n5843), .Y(
        n12710) );
  CLKMX2X2 U11236 ( .A(\I_cache/cache[6][16] ), .B(n9767), .S0(n5886), .Y(
        n12711) );
  CLKMX2X2 U11237 ( .A(\I_cache/cache[5][16] ), .B(n9767), .S0(n5752), .Y(
        n12712) );
  CLKMX2X2 U11238 ( .A(\I_cache/cache[4][16] ), .B(n9767), .S0(n5799), .Y(
        n12713) );
  CLKMX2X2 U11239 ( .A(\I_cache/cache[3][16] ), .B(n9767), .S0(n5664), .Y(
        n12714) );
  CLKMX2X2 U11240 ( .A(\I_cache/cache[2][16] ), .B(n9767), .S0(n5709), .Y(
        n12715) );
  CLKMX2X2 U11241 ( .A(\I_cache/cache[1][16] ), .B(n9767), .S0(n5575), .Y(
        n12716) );
  CLKMX2X2 U11242 ( .A(\I_cache/cache[0][16] ), .B(n9767), .S0(n5618), .Y(
        n12717) );
  CLKMX2X2 U11243 ( .A(\I_cache/cache[7][15] ), .B(n10072), .S0(n5846), .Y(
        n12718) );
  CLKMX2X2 U11244 ( .A(\I_cache/cache[6][15] ), .B(n10072), .S0(n5887), .Y(
        n12719) );
  CLKMX2X2 U11245 ( .A(\I_cache/cache[5][15] ), .B(n10072), .S0(n5753), .Y(
        n12720) );
  CLKMX2X2 U11246 ( .A(\I_cache/cache[4][15] ), .B(n10072), .S0(n5799), .Y(
        n12721) );
  CLKMX2X2 U11247 ( .A(\I_cache/cache[3][15] ), .B(n10072), .S0(n5663), .Y(
        n12722) );
  CLKMX2X2 U11248 ( .A(\I_cache/cache[2][15] ), .B(n10072), .S0(n5709), .Y(
        n12723) );
  CLKMX2X2 U11249 ( .A(\I_cache/cache[1][15] ), .B(n10072), .S0(n5575), .Y(
        n12724) );
  CLKMX2X2 U11250 ( .A(\I_cache/cache[0][15] ), .B(n10072), .S0(n5620), .Y(
        n12725) );
  CLKMX2X2 U11251 ( .A(\I_cache/cache[7][14] ), .B(n10251), .S0(n5850), .Y(
        n12726) );
  CLKMX2X2 U11252 ( .A(\I_cache/cache[6][14] ), .B(n10251), .S0(n5893), .Y(
        n12727) );
  CLKMX2X2 U11253 ( .A(\I_cache/cache[5][14] ), .B(n10251), .S0(n5759), .Y(
        n12728) );
  CLKMX2X2 U11254 ( .A(\I_cache/cache[4][14] ), .B(n10251), .S0(n5806), .Y(
        n12729) );
  CLKMX2X2 U11255 ( .A(\I_cache/cache[3][14] ), .B(n10251), .S0(n5671), .Y(
        n12730) );
  CLKMX2X2 U11256 ( .A(\I_cache/cache[2][14] ), .B(n10251), .S0(n5716), .Y(
        n12731) );
  CLKMX2X2 U11257 ( .A(\I_cache/cache[1][14] ), .B(n10251), .S0(n5582), .Y(
        n12732) );
  CLKMX2X2 U11258 ( .A(\I_cache/cache[0][14] ), .B(n10251), .S0(n5625), .Y(
        n12733) );
  CLKMX2X2 U11259 ( .A(\I_cache/cache[7][13] ), .B(n10229), .S0(n5845), .Y(
        n12734) );
  CLKMX2X2 U11260 ( .A(\I_cache/cache[6][13] ), .B(n10229), .S0(n5889), .Y(
        n12735) );
  CLKMX2X2 U11261 ( .A(\I_cache/cache[5][13] ), .B(n10229), .S0(n5755), .Y(
        n12736) );
  CLKMX2X2 U11262 ( .A(\I_cache/cache[4][13] ), .B(n10229), .S0(n5801), .Y(
        n12737) );
  CLKMX2X2 U11263 ( .A(\I_cache/cache[3][13] ), .B(n10229), .S0(n5666), .Y(
        n12738) );
  CLKMX2X2 U11264 ( .A(\I_cache/cache[2][13] ), .B(n10229), .S0(n5711), .Y(
        n12739) );
  CLKMX2X2 U11265 ( .A(\I_cache/cache[1][13] ), .B(n10229), .S0(n5576), .Y(
        n12740) );
  CLKMX2X2 U11266 ( .A(\I_cache/cache[0][13] ), .B(n10229), .S0(n5619), .Y(
        n12741) );
  CLKMX2X2 U11267 ( .A(\I_cache/cache[7][12] ), .B(n10131), .S0(n5845), .Y(
        n12742) );
  CLKMX2X2 U11268 ( .A(\I_cache/cache[6][12] ), .B(n10131), .S0(n5889), .Y(
        n12743) );
  CLKMX2X2 U11269 ( .A(\I_cache/cache[5][12] ), .B(n10131), .S0(n5755), .Y(
        n12744) );
  CLKMX2X2 U11270 ( .A(\I_cache/cache[4][12] ), .B(n10131), .S0(n5801), .Y(
        n12745) );
  CLKMX2X2 U11271 ( .A(\I_cache/cache[3][12] ), .B(n10131), .S0(n5666), .Y(
        n12746) );
  CLKMX2X2 U11272 ( .A(\I_cache/cache[2][12] ), .B(n10131), .S0(n5711), .Y(
        n12747) );
  CLKMX2X2 U11273 ( .A(\I_cache/cache[1][12] ), .B(n10131), .S0(n5577), .Y(
        n12748) );
  CLKMX2X2 U11274 ( .A(\I_cache/cache[0][12] ), .B(n10131), .S0(n5620), .Y(
        n12749) );
  CLKMX2X2 U11275 ( .A(\I_cache/cache[7][11] ), .B(n10095), .S0(n5845), .Y(
        n12750) );
  CLKMX2X2 U11276 ( .A(\I_cache/cache[6][11] ), .B(n10095), .S0(n5889), .Y(
        n12751) );
  CLKMX2X2 U11277 ( .A(\I_cache/cache[5][11] ), .B(n10095), .S0(n5755), .Y(
        n12752) );
  CLKMX2X2 U11278 ( .A(\I_cache/cache[4][11] ), .B(n10095), .S0(n5801), .Y(
        n12753) );
  CLKMX2X2 U11279 ( .A(\I_cache/cache[3][11] ), .B(n10095), .S0(n5666), .Y(
        n12754) );
  CLKMX2X2 U11280 ( .A(\I_cache/cache[2][11] ), .B(n10095), .S0(n5711), .Y(
        n12755) );
  CLKMX2X2 U11281 ( .A(\I_cache/cache[1][11] ), .B(n10095), .S0(n5577), .Y(
        n12756) );
  CLKMX2X2 U11282 ( .A(\I_cache/cache[0][11] ), .B(n10095), .S0(n5620), .Y(
        n12757) );
  CLKMX2X2 U11283 ( .A(\I_cache/cache[7][10] ), .B(n9844), .S0(n5846), .Y(
        n12758) );
  CLKMX2X2 U11284 ( .A(\I_cache/cache[6][10] ), .B(n9844), .S0(n5887), .Y(
        n12759) );
  CLKMX2X2 U11285 ( .A(\I_cache/cache[5][10] ), .B(n9844), .S0(n5756), .Y(
        n12760) );
  CLKMX2X2 U11286 ( .A(\I_cache/cache[4][10] ), .B(n9844), .S0(n5802), .Y(
        n12761) );
  CLKMX2X2 U11287 ( .A(\I_cache/cache[3][10] ), .B(n9844), .S0(n5667), .Y(
        n12762) );
  CLKMX2X2 U11288 ( .A(\I_cache/cache[2][10] ), .B(n9844), .S0(n5712), .Y(
        n12763) );
  CLKMX2X2 U11289 ( .A(\I_cache/cache[1][10] ), .B(n9844), .S0(n5578), .Y(
        n12764) );
  CLKMX2X2 U11290 ( .A(\I_cache/cache[0][10] ), .B(n9844), .S0(n5621), .Y(
        n12765) );
  CLKMX2X2 U11291 ( .A(\I_cache/cache[7][9] ), .B(n9888), .S0(n5846), .Y(
        n12766) );
  CLKMX2X2 U11292 ( .A(\I_cache/cache[6][9] ), .B(n9888), .S0(n5889), .Y(
        n12767) );
  CLKMX2X2 U11293 ( .A(\I_cache/cache[5][9] ), .B(n9888), .S0(n5756), .Y(
        n12768) );
  CLKMX2X2 U11294 ( .A(\I_cache/cache[4][9] ), .B(n9888), .S0(n5802), .Y(
        n12769) );
  CLKMX2X2 U11295 ( .A(\I_cache/cache[3][9] ), .B(n9888), .S0(n5667), .Y(
        n12770) );
  CLKMX2X2 U11296 ( .A(\I_cache/cache[2][9] ), .B(n9888), .S0(n5712), .Y(
        n12771) );
  CLKMX2X2 U11297 ( .A(\I_cache/cache[1][9] ), .B(n9888), .S0(n5578), .Y(
        n12772) );
  CLKMX2X2 U11298 ( .A(\I_cache/cache[0][9] ), .B(n9888), .S0(n5621), .Y(
        n12773) );
  CLKMX2X2 U11299 ( .A(\I_cache/cache[7][8] ), .B(n9866), .S0(n5846), .Y(
        n12774) );
  CLKMX2X2 U11300 ( .A(\I_cache/cache[6][8] ), .B(n9866), .S0(n5885), .Y(
        n12775) );
  CLKMX2X2 U11301 ( .A(\I_cache/cache[5][8] ), .B(n9866), .S0(n5756), .Y(
        n12776) );
  CLKMX2X2 U11302 ( .A(\I_cache/cache[4][8] ), .B(n9866), .S0(n5802), .Y(
        n12777) );
  CLKMX2X2 U11303 ( .A(\I_cache/cache[3][8] ), .B(n9866), .S0(n5667), .Y(
        n12778) );
  CLKMX2X2 U11304 ( .A(\I_cache/cache[2][8] ), .B(n9866), .S0(n5712), .Y(
        n12779) );
  CLKMX2X2 U11305 ( .A(\I_cache/cache[1][8] ), .B(n9866), .S0(n5578), .Y(
        n12780) );
  CLKMX2X2 U11306 ( .A(\I_cache/cache[0][8] ), .B(n9866), .S0(n5621), .Y(
        n12781) );
  CLKMX2X2 U11307 ( .A(\I_cache/cache[7][7] ), .B(n9910), .S0(n5845), .Y(
        n12782) );
  CLKMX2X2 U11308 ( .A(\I_cache/cache[6][7] ), .B(n9910), .S0(n5889), .Y(
        n12783) );
  CLKMX2X2 U11309 ( .A(\I_cache/cache[5][7] ), .B(n9910), .S0(n5755), .Y(
        n12784) );
  CLKMX2X2 U11310 ( .A(\I_cache/cache[4][7] ), .B(n9910), .S0(n5801), .Y(
        n12785) );
  CLKMX2X2 U11311 ( .A(\I_cache/cache[3][7] ), .B(n9910), .S0(n5666), .Y(
        n12786) );
  CLKMX2X2 U11312 ( .A(\I_cache/cache[2][7] ), .B(n9910), .S0(n5711), .Y(
        n12787) );
  CLKMX2X2 U11313 ( .A(\I_cache/cache[1][7] ), .B(n9910), .S0(n5579), .Y(
        n12788) );
  CLKMX2X2 U11314 ( .A(\I_cache/cache[0][7] ), .B(n9910), .S0(n5622), .Y(
        n12789) );
  CLKMX2X2 U11315 ( .A(\I_cache/cache[7][6] ), .B(n9932), .S0(n5847), .Y(
        n12790) );
  CLKMX2X2 U11316 ( .A(\I_cache/cache[6][6] ), .B(n9932), .S0(n5890), .Y(
        n12791) );
  CLKMX2X2 U11317 ( .A(\I_cache/cache[5][6] ), .B(n9932), .S0(n5757), .Y(
        n12792) );
  CLKMX2X2 U11318 ( .A(\I_cache/cache[4][6] ), .B(n9932), .S0(n5803), .Y(
        n12793) );
  CLKMX2X2 U11319 ( .A(\I_cache/cache[3][6] ), .B(n9932), .S0(n5668), .Y(
        n12794) );
  CLKMX2X2 U11320 ( .A(\I_cache/cache[2][6] ), .B(n9932), .S0(n5713), .Y(
        n12795) );
  CLKMX2X2 U11321 ( .A(\I_cache/cache[1][6] ), .B(n9932), .S0(n5579), .Y(
        n12796) );
  CLKMX2X2 U11322 ( .A(\I_cache/cache[0][6] ), .B(n9932), .S0(n5622), .Y(
        n12797) );
  CLKMX2X2 U11323 ( .A(\I_cache/cache[7][5] ), .B(n9725), .S0(n5842), .Y(
        n12798) );
  CLKMX2X2 U11324 ( .A(\I_cache/cache[6][5] ), .B(n9725), .S0(n5885), .Y(
        n12799) );
  CLKMX2X2 U11325 ( .A(\I_cache/cache[5][5] ), .B(n9725), .S0(n5752), .Y(
        n12800) );
  CLKMX2X2 U11326 ( .A(\I_cache/cache[4][5] ), .B(n9725), .S0(n5798), .Y(
        n12801) );
  CLKMX2X2 U11327 ( .A(\I_cache/cache[3][5] ), .B(n9725), .S0(n5663), .Y(
        n12802) );
  CLKMX2X2 U11328 ( .A(\I_cache/cache[2][5] ), .B(n9725), .S0(n5708), .Y(
        n12803) );
  CLKMX2X2 U11329 ( .A(\I_cache/cache[1][5] ), .B(n9725), .S0(n5574), .Y(
        n12804) );
  CLKMX2X2 U11330 ( .A(\I_cache/cache[0][5] ), .B(n9725), .S0(n5617), .Y(
        n12805) );
  CLKMX2X2 U11331 ( .A(\I_cache/cache[7][4] ), .B(n10865), .S0(n5850), .Y(
        n12806) );
  CLKMX2X2 U11332 ( .A(\I_cache/cache[6][4] ), .B(n10865), .S0(n5893), .Y(
        n12807) );
  CLKMX2X2 U11333 ( .A(\I_cache/cache[5][4] ), .B(n10865), .S0(n5759), .Y(
        n12808) );
  CLKMX2X2 U11334 ( .A(\I_cache/cache[4][4] ), .B(n10865), .S0(n5806), .Y(
        n12809) );
  CLKMX2X2 U11335 ( .A(\I_cache/cache[3][4] ), .B(n10865), .S0(n5671), .Y(
        n12810) );
  CLKMX2X2 U11336 ( .A(\I_cache/cache[2][4] ), .B(n10865), .S0(n5716), .Y(
        n12811) );
  CLKMX2X2 U11337 ( .A(\I_cache/cache[1][4] ), .B(n10865), .S0(n5582), .Y(
        n12812) );
  CLKMX2X2 U11338 ( .A(\I_cache/cache[0][4] ), .B(n10865), .S0(n5625), .Y(
        n12813) );
  CLKMX2X2 U11339 ( .A(\I_cache/cache[7][3] ), .B(n10959), .S0(n5842), .Y(
        n12814) );
  CLKMX2X2 U11340 ( .A(\I_cache/cache[6][3] ), .B(n10959), .S0(n5887), .Y(
        n12815) );
  CLKMX2X2 U11341 ( .A(\I_cache/cache[5][3] ), .B(n10959), .S0(n4828), .Y(
        n12816) );
  CLKMX2X2 U11342 ( .A(\I_cache/cache[4][3] ), .B(n10959), .S0(n5799), .Y(
        n12817) );
  CLKMX2X2 U11343 ( .A(\I_cache/cache[3][3] ), .B(n10959), .S0(n5664), .Y(
        n12818) );
  CLKMX2X2 U11344 ( .A(\I_cache/cache[2][3] ), .B(n10959), .S0(n5711), .Y(
        n12819) );
  CLKMX2X2 U11345 ( .A(\I_cache/cache[1][3] ), .B(n10959), .S0(n5581), .Y(
        n12820) );
  CLKMX2X2 U11346 ( .A(\I_cache/cache[0][3] ), .B(n10959), .S0(n5620), .Y(
        n12821) );
  CLKMX2X2 U11347 ( .A(\I_cache/cache[7][2] ), .B(n10930), .S0(n5843), .Y(
        n12822) );
  CLKMX2X2 U11348 ( .A(\I_cache/cache[6][2] ), .B(n10930), .S0(n5888), .Y(
        n12823) );
  CLKMX2X2 U11349 ( .A(\I_cache/cache[5][2] ), .B(n10930), .S0(n4829), .Y(
        n12824) );
  CLKMX2X2 U11350 ( .A(\I_cache/cache[4][2] ), .B(n10930), .S0(n5800), .Y(
        n12825) );
  CLKMX2X2 U11351 ( .A(\I_cache/cache[3][2] ), .B(n10930), .S0(n5666), .Y(
        n12826) );
  CLKMX2X2 U11352 ( .A(\I_cache/cache[2][2] ), .B(n10930), .S0(n5710), .Y(
        n12827) );
  CLKMX2X2 U11353 ( .A(\I_cache/cache[1][2] ), .B(n10930), .S0(n5580), .Y(
        n12828) );
  CLKMX2X2 U11354 ( .A(\I_cache/cache[0][2] ), .B(n10930), .S0(n5622), .Y(
        n12829) );
  CLKMX2X2 U11355 ( .A(\I_cache/cache[7][1] ), .B(n10888), .S0(n5842), .Y(
        n12830) );
  CLKMX2X2 U11356 ( .A(\I_cache/cache[6][1] ), .B(n10888), .S0(n5885), .Y(
        n12831) );
  CLKMX2X2 U11357 ( .A(\I_cache/cache[5][1] ), .B(n10888), .S0(n5753), .Y(
        n12832) );
  CLKMX2X2 U11358 ( .A(\I_cache/cache[4][1] ), .B(n10888), .S0(n5798), .Y(
        n12833) );
  CLKMX2X2 U11359 ( .A(\I_cache/cache[3][1] ), .B(n10888), .S0(n5663), .Y(
        n12834) );
  CLKMX2X2 U11360 ( .A(\I_cache/cache[2][1] ), .B(n10888), .S0(n5708), .Y(
        n12835) );
  CLKMX2X2 U11361 ( .A(\I_cache/cache[1][1] ), .B(n10888), .S0(n5574), .Y(
        n12836) );
  CLKMX2X2 U11362 ( .A(\I_cache/cache[0][1] ), .B(n10888), .S0(n5619), .Y(
        n12837) );
  CLKMX2X2 U11363 ( .A(\I_cache/cache[7][0] ), .B(n10822), .S0(n5850), .Y(
        n12845) );
  CLKMX2X2 U11364 ( .A(\I_cache/cache[6][0] ), .B(n10822), .S0(n5893), .Y(
        n12838) );
  CLKMX2X2 U11365 ( .A(\I_cache/cache[5][0] ), .B(n10822), .S0(n5759), .Y(
        n12839) );
  CLKMX2X2 U11366 ( .A(\I_cache/cache[4][0] ), .B(n10822), .S0(n5806), .Y(
        n12840) );
  CLKMX2X2 U11367 ( .A(\I_cache/cache[3][0] ), .B(n10822), .S0(n5671), .Y(
        n12841) );
  CLKMX2X2 U11368 ( .A(\I_cache/cache[2][0] ), .B(n10822), .S0(n5716), .Y(
        n12842) );
  CLKMX2X2 U11369 ( .A(\I_cache/cache[1][0] ), .B(n10822), .S0(n5582), .Y(
        n12843) );
  CLKMX2X2 U11370 ( .A(\I_cache/cache[0][0] ), .B(n10822), .S0(n5625), .Y(
        n12844) );
  MX2XL U11371 ( .A(\D_cache/cache[7][142] ), .B(n11051), .S0(n3561), .Y(
        \D_cache/n653 ) );
  MX2XL U11372 ( .A(\D_cache/cache[6][142] ), .B(n11051), .S0(n5368), .Y(
        \D_cache/n654 ) );
  MX2XL U11373 ( .A(\D_cache/cache[5][142] ), .B(n11051), .S0(n5344), .Y(
        \D_cache/n655 ) );
  MX2XL U11374 ( .A(\D_cache/cache[4][142] ), .B(n11051), .S0(n5317), .Y(
        \D_cache/n656 ) );
  MX2XL U11375 ( .A(\D_cache/cache[3][142] ), .B(n11051), .S0(n5272), .Y(
        \D_cache/n657 ) );
  MX2XL U11376 ( .A(\D_cache/cache[2][142] ), .B(n11051), .S0(n5230), .Y(
        \D_cache/n658 ) );
  MX2XL U11377 ( .A(\D_cache/cache[1][142] ), .B(n11051), .S0(n5202), .Y(
        \D_cache/n659 ) );
  MX2XL U11378 ( .A(\D_cache/cache[0][142] ), .B(n11051), .S0(n5162), .Y(
        \D_cache/n660 ) );
  MX2XL U11379 ( .A(\I_cache/cache[6][95] ), .B(n6577), .S0(n5891), .Y(n12079)
         );
  MX2XL U11380 ( .A(\I_cache/cache[5][95] ), .B(n6577), .S0(n5755), .Y(n12080)
         );
  MX2XL U11381 ( .A(\I_cache/cache[4][95] ), .B(n6577), .S0(n5804), .Y(n12081)
         );
  MX2XL U11382 ( .A(\I_cache/cache[3][95] ), .B(n6577), .S0(n5669), .Y(n12082)
         );
  MX2XL U11383 ( .A(\I_cache/cache[2][95] ), .B(n6577), .S0(n5714), .Y(n12083)
         );
  MX2XL U11384 ( .A(\I_cache/cache[1][95] ), .B(n6577), .S0(n5577), .Y(n12084)
         );
  MX2XL U11385 ( .A(\I_cache/cache[0][95] ), .B(n6577), .S0(n5621), .Y(n12085)
         );
  MX2XL U11386 ( .A(\I_cache/cache[6][94] ), .B(n9666), .S0(n5887), .Y(n12087)
         );
  MX2XL U11387 ( .A(\I_cache/cache[5][94] ), .B(n9666), .S0(n5753), .Y(n12088)
         );
  MX2XL U11388 ( .A(\I_cache/cache[4][94] ), .B(n9666), .S0(n5799), .Y(n12089)
         );
  MX2XL U11389 ( .A(\I_cache/cache[3][94] ), .B(n9666), .S0(n5671), .Y(n12090)
         );
  MX2XL U11390 ( .A(\I_cache/cache[2][94] ), .B(n9666), .S0(n5709), .Y(n12091)
         );
  MX2XL U11391 ( .A(\I_cache/cache[1][94] ), .B(n9666), .S0(n5579), .Y(n12092)
         );
  MX2XL U11392 ( .A(\I_cache/cache[0][94] ), .B(n9666), .S0(n5621), .Y(n12093)
         );
  MX2XL U11393 ( .A(\I_cache/cache[6][93] ), .B(n9688), .S0(n5885), .Y(n12095)
         );
  MX2XL U11394 ( .A(\I_cache/cache[5][93] ), .B(n9688), .S0(n5754), .Y(n12096)
         );
  MX2XL U11395 ( .A(\I_cache/cache[4][93] ), .B(n9688), .S0(n5798), .Y(n12097)
         );
  MX2XL U11396 ( .A(\I_cache/cache[3][93] ), .B(n9688), .S0(n5663), .Y(n12098)
         );
  MX2XL U11397 ( .A(\I_cache/cache[2][93] ), .B(n9688), .S0(n5708), .Y(n12099)
         );
  MX2XL U11398 ( .A(\I_cache/cache[1][93] ), .B(n9688), .S0(n5574), .Y(n12100)
         );
  MX2XL U11399 ( .A(\I_cache/cache[0][93] ), .B(n9688), .S0(n5617), .Y(n12101)
         );
  MX2XL U11400 ( .A(\I_cache/cache[6][92] ), .B(n9636), .S0(n5887), .Y(n12103)
         );
  MX2XL U11401 ( .A(\I_cache/cache[5][92] ), .B(n9636), .S0(n5753), .Y(n12104)
         );
  MX2XL U11402 ( .A(\I_cache/cache[4][92] ), .B(n9636), .S0(n5802), .Y(n12105)
         );
  MX2XL U11403 ( .A(\I_cache/cache[3][92] ), .B(n9636), .S0(n5664), .Y(n12106)
         );
  MX2XL U11404 ( .A(\I_cache/cache[2][92] ), .B(n9636), .S0(n5709), .Y(n12107)
         );
  MX2XL U11405 ( .A(\I_cache/cache[1][92] ), .B(n9636), .S0(n5575), .Y(n12108)
         );
  MX2XL U11406 ( .A(\I_cache/cache[0][92] ), .B(n9636), .S0(n5625), .Y(n12109)
         );
  MX2XL U11407 ( .A(\I_cache/cache[6][91] ), .B(n9614), .S0(n5887), .Y(n12111)
         );
  MX2XL U11408 ( .A(\I_cache/cache[5][91] ), .B(n9614), .S0(n5753), .Y(n12112)
         );
  MX2XL U11409 ( .A(\I_cache/cache[4][91] ), .B(n9614), .S0(n5800), .Y(n12113)
         );
  MX2XL U11410 ( .A(\I_cache/cache[3][91] ), .B(n9614), .S0(n5666), .Y(n12114)
         );
  MX2XL U11411 ( .A(\I_cache/cache[2][91] ), .B(n9614), .S0(n5709), .Y(n12115)
         );
  MX2XL U11412 ( .A(\I_cache/cache[1][91] ), .B(n9614), .S0(n5575), .Y(n12116)
         );
  MX2XL U11413 ( .A(\I_cache/cache[0][91] ), .B(n9614), .S0(n5624), .Y(n12117)
         );
  MX2XL U11414 ( .A(\I_cache/cache[6][90] ), .B(n6592), .S0(n5891), .Y(n12119)
         );
  MX2XL U11415 ( .A(\I_cache/cache[5][90] ), .B(n6592), .S0(n5756), .Y(n12120)
         );
  MX2XL U11416 ( .A(\I_cache/cache[4][90] ), .B(n6592), .S0(n5804), .Y(n12121)
         );
  MX2XL U11417 ( .A(\I_cache/cache[3][90] ), .B(n6592), .S0(n5669), .Y(n12122)
         );
  MX2XL U11418 ( .A(\I_cache/cache[2][90] ), .B(n6592), .S0(n5714), .Y(n12123)
         );
  MX2XL U11419 ( .A(\I_cache/cache[1][90] ), .B(n6592), .S0(n5578), .Y(n12124)
         );
  MX2XL U11420 ( .A(\I_cache/cache[0][90] ), .B(n6592), .S0(n5625), .Y(n12125)
         );
  MX2XL U11421 ( .A(\I_cache/cache[1][88] ), .B(n6547), .S0(n5582), .Y(n12140)
         );
  MX2XL U11422 ( .A(\I_cache/cache[6][87] ), .B(n10011), .S0(n5887), .Y(n12143) );
  MX2XL U11423 ( .A(\I_cache/cache[5][87] ), .B(n10011), .S0(n5756), .Y(n12144) );
  MX2XL U11424 ( .A(\I_cache/cache[4][87] ), .B(n10011), .S0(n5802), .Y(n12145) );
  MX2XL U11425 ( .A(\I_cache/cache[3][87] ), .B(n10011), .S0(n5667), .Y(n12146) );
  MX2XL U11426 ( .A(\I_cache/cache[2][87] ), .B(n10011), .S0(n5712), .Y(n12147) );
  MX2XL U11427 ( .A(\I_cache/cache[1][87] ), .B(n10011), .S0(n5576), .Y(n12148) );
  MX2XL U11428 ( .A(\I_cache/cache[0][87] ), .B(n10011), .S0(n5619), .Y(n12149) );
  MX2XL U11429 ( .A(\I_cache/cache[6][86] ), .B(n9967), .S0(n5890), .Y(n12151)
         );
  MX2XL U11430 ( .A(\I_cache/cache[5][86] ), .B(n9967), .S0(n5757), .Y(n12152)
         );
  MX2XL U11431 ( .A(\I_cache/cache[4][86] ), .B(n9967), .S0(n5803), .Y(n12153)
         );
  MX2XL U11432 ( .A(\I_cache/cache[3][86] ), .B(n9967), .S0(n5668), .Y(n12154)
         );
  MX2XL U11433 ( .A(\I_cache/cache[2][86] ), .B(n9967), .S0(n5713), .Y(n12155)
         );
  MX2XL U11434 ( .A(\I_cache/cache[1][86] ), .B(n9967), .S0(n5579), .Y(n12156)
         );
  MX2XL U11435 ( .A(\I_cache/cache[0][86] ), .B(n9967), .S0(n5622), .Y(n12157)
         );
  MX2XL U11436 ( .A(\I_cache/cache[6][84] ), .B(n9778), .S0(n5886), .Y(n12167)
         );
  MX2XL U11437 ( .A(\I_cache/cache[5][84] ), .B(n9778), .S0(n5752), .Y(n12168)
         );
  MX2XL U11438 ( .A(\I_cache/cache[4][84] ), .B(n9778), .S0(n5799), .Y(n12169)
         );
  MX2XL U11439 ( .A(\I_cache/cache[3][84] ), .B(n9778), .S0(n5664), .Y(n12170)
         );
  MX2XL U11440 ( .A(\I_cache/cache[2][84] ), .B(n9778), .S0(n5709), .Y(n12171)
         );
  MX2XL U11441 ( .A(\I_cache/cache[1][84] ), .B(n9778), .S0(n5576), .Y(n12172)
         );
  MX2XL U11442 ( .A(\I_cache/cache[0][84] ), .B(n9778), .S0(n5618), .Y(n12173)
         );
  MX2XL U11443 ( .A(\I_cache/cache[5][82] ), .B(n9770), .S0(n5752), .Y(n12184)
         );
  MX2XL U11444 ( .A(\I_cache/cache[2][82] ), .B(n9770), .S0(n5708), .Y(n12187)
         );
  MX2XL U11445 ( .A(\I_cache/cache[6][81] ), .B(n6567), .S0(n5891), .Y(n12191)
         );
  MX2XL U11446 ( .A(\I_cache/cache[5][81] ), .B(n6567), .S0(n5757), .Y(n12192)
         );
  MX2XL U11447 ( .A(\I_cache/cache[4][81] ), .B(n6567), .S0(n5804), .Y(n12193)
         );
  MX2XL U11448 ( .A(\I_cache/cache[3][81] ), .B(n6567), .S0(n5669), .Y(n12194)
         );
  MX2XL U11449 ( .A(\I_cache/cache[2][81] ), .B(n6567), .S0(n5714), .Y(n12195)
         );
  MX2XL U11450 ( .A(\I_cache/cache[1][81] ), .B(n6567), .S0(n5577), .Y(n12196)
         );
  MX2XL U11451 ( .A(\I_cache/cache[0][81] ), .B(n6567), .S0(n5622), .Y(n12197)
         );
  MX2XL U11452 ( .A(\I_cache/cache[2][80] ), .B(n9752), .S0(n5708), .Y(n12203)
         );
  MX2XL U11453 ( .A(\I_cache/cache[6][74] ), .B(n9829), .S0(n5886), .Y(n12247)
         );
  MX2XL U11454 ( .A(\I_cache/cache[5][74] ), .B(n9829), .S0(n5752), .Y(n12248)
         );
  MX2XL U11455 ( .A(\I_cache/cache[4][74] ), .B(n9829), .S0(n5799), .Y(n12249)
         );
  MX2XL U11456 ( .A(\I_cache/cache[3][74] ), .B(n9829), .S0(n5664), .Y(n12250)
         );
  MX2XL U11457 ( .A(\I_cache/cache[2][74] ), .B(n9829), .S0(n5710), .Y(n12251)
         );
  MX2XL U11458 ( .A(\I_cache/cache[1][74] ), .B(n9829), .S0(n5578), .Y(n12252)
         );
  MX2XL U11459 ( .A(\I_cache/cache[0][74] ), .B(n9829), .S0(n5618), .Y(n12253)
         );
  MX2XL U11460 ( .A(\I_cache/cache[6][73] ), .B(n9873), .S0(n5885), .Y(n12255)
         );
  MX2XL U11461 ( .A(\I_cache/cache[5][73] ), .B(n9873), .S0(n5756), .Y(n12256)
         );
  MX2XL U11462 ( .A(\I_cache/cache[4][73] ), .B(n9873), .S0(n5802), .Y(n12257)
         );
  MX2XL U11463 ( .A(\I_cache/cache[3][73] ), .B(n9873), .S0(n5667), .Y(n12258)
         );
  MX2XL U11464 ( .A(\I_cache/cache[2][73] ), .B(n9873), .S0(n5712), .Y(n12259)
         );
  MX2XL U11465 ( .A(\I_cache/cache[1][73] ), .B(n9873), .S0(n5578), .Y(n12260)
         );
  MX2XL U11466 ( .A(\I_cache/cache[0][73] ), .B(n9873), .S0(n5621), .Y(n12261)
         );
  MX2XL U11467 ( .A(\I_cache/cache[6][72] ), .B(n9851), .S0(n5889), .Y(n12263)
         );
  MX2XL U11468 ( .A(\I_cache/cache[5][72] ), .B(n9851), .S0(n5756), .Y(n12264)
         );
  MX2XL U11469 ( .A(\I_cache/cache[4][72] ), .B(n9851), .S0(n5802), .Y(n12265)
         );
  MX2XL U11470 ( .A(\I_cache/cache[3][72] ), .B(n9851), .S0(n5667), .Y(n12266)
         );
  MX2XL U11471 ( .A(\I_cache/cache[2][72] ), .B(n9851), .S0(n5712), .Y(n12267)
         );
  MX2XL U11472 ( .A(\I_cache/cache[1][72] ), .B(n9851), .S0(n5578), .Y(n12268)
         );
  MX2XL U11473 ( .A(\I_cache/cache[0][72] ), .B(n9851), .S0(n5621), .Y(n12269)
         );
  MX2XL U11474 ( .A(\I_cache/cache[6][71] ), .B(n9895), .S0(n5890), .Y(n12271)
         );
  MX2XL U11475 ( .A(\I_cache/cache[5][71] ), .B(n9895), .S0(n5756), .Y(n12272)
         );
  MX2XL U11476 ( .A(\I_cache/cache[4][71] ), .B(n9895), .S0(n5802), .Y(n12273)
         );
  MX2XL U11477 ( .A(\I_cache/cache[3][71] ), .B(n9895), .S0(n5667), .Y(n12274)
         );
  MX2XL U11478 ( .A(\I_cache/cache[2][71] ), .B(n9895), .S0(n5712), .Y(n12275)
         );
  MX2XL U11479 ( .A(\I_cache/cache[1][71] ), .B(n9895), .S0(n5578), .Y(n12276)
         );
  MX2XL U11480 ( .A(\I_cache/cache[0][71] ), .B(n9895), .S0(n5621), .Y(n12277)
         );
  MX2XL U11481 ( .A(\I_cache/cache[6][70] ), .B(n9917), .S0(n5890), .Y(n12279)
         );
  MX2XL U11482 ( .A(\I_cache/cache[5][70] ), .B(n9917), .S0(n5757), .Y(n12280)
         );
  MX2XL U11483 ( .A(\I_cache/cache[4][70] ), .B(n9917), .S0(n5803), .Y(n12281)
         );
  MX2XL U11484 ( .A(\I_cache/cache[3][70] ), .B(n9917), .S0(n5668), .Y(n12282)
         );
  MX2XL U11485 ( .A(\I_cache/cache[2][70] ), .B(n9917), .S0(n5713), .Y(n12283)
         );
  MX2XL U11486 ( .A(\I_cache/cache[1][70] ), .B(n9917), .S0(n5579), .Y(n12284)
         );
  MX2XL U11487 ( .A(\I_cache/cache[0][70] ), .B(n9917), .S0(n5622), .Y(n12285)
         );
  MX2XL U11488 ( .A(\I_cache/cache[6][69] ), .B(n9710), .S0(n5885), .Y(n12287)
         );
  MX2XL U11489 ( .A(\I_cache/cache[5][69] ), .B(n9710), .S0(n5752), .Y(n12288)
         );
  MX2XL U11490 ( .A(\I_cache/cache[4][69] ), .B(n9710), .S0(n5798), .Y(n12289)
         );
  MX2XL U11491 ( .A(\I_cache/cache[3][69] ), .B(n9710), .S0(n5663), .Y(n12290)
         );
  MX2XL U11492 ( .A(\I_cache/cache[2][69] ), .B(n9710), .S0(n5708), .Y(n12291)
         );
  MX2XL U11493 ( .A(\I_cache/cache[1][69] ), .B(n9710), .S0(n5574), .Y(n12292)
         );
  MX2XL U11494 ( .A(\I_cache/cache[0][69] ), .B(n9710), .S0(n5617), .Y(n12293)
         );
  MX2XL U11495 ( .A(\I_cache/cache[6][68] ), .B(n6542), .S0(n5891), .Y(n12295)
         );
  MX2XL U11496 ( .A(\I_cache/cache[5][68] ), .B(n6542), .S0(n5758), .Y(n12296)
         );
  MX2XL U11497 ( .A(\I_cache/cache[4][68] ), .B(n6542), .S0(n5804), .Y(n12297)
         );
  MX2XL U11498 ( .A(\I_cache/cache[3][68] ), .B(n6542), .S0(n5669), .Y(n12298)
         );
  MX2XL U11499 ( .A(\I_cache/cache[2][68] ), .B(n6542), .S0(n5714), .Y(n12299)
         );
  MX2XL U11500 ( .A(\I_cache/cache[1][68] ), .B(n6542), .S0(n5579), .Y(n12300)
         );
  MX2XL U11501 ( .A(\I_cache/cache[0][68] ), .B(n6542), .S0(n5623), .Y(n12301)
         );
  MX2XL U11502 ( .A(\I_cache/cache[6][63] ), .B(n6582), .S0(n5891), .Y(n12335)
         );
  MX2XL U11503 ( .A(\I_cache/cache[5][63] ), .B(n6582), .S0(n5756), .Y(n12336)
         );
  MX2XL U11504 ( .A(\I_cache/cache[4][63] ), .B(n6582), .S0(n5804), .Y(n12337)
         );
  MX2XL U11505 ( .A(\I_cache/cache[3][63] ), .B(n6582), .S0(n5669), .Y(n12338)
         );
  MX2XL U11506 ( .A(\I_cache/cache[2][63] ), .B(n6582), .S0(n5714), .Y(n12339)
         );
  MX2XL U11507 ( .A(\I_cache/cache[1][63] ), .B(n6582), .S0(n5578), .Y(n12340)
         );
  MX2XL U11508 ( .A(\I_cache/cache[0][63] ), .B(n6582), .S0(n5621), .Y(n12341)
         );
  MX2XL U11509 ( .A(\I_cache/cache[6][62] ), .B(n9671), .S0(n5893), .Y(n12343)
         );
  MX2XL U11510 ( .A(\I_cache/cache[5][62] ), .B(n9671), .S0(n5754), .Y(n12344)
         );
  MX2XL U11511 ( .A(\I_cache/cache[4][62] ), .B(n9671), .S0(n5806), .Y(n12345)
         );
  MX2XL U11512 ( .A(\I_cache/cache[3][62] ), .B(n9671), .S0(n5671), .Y(n12346)
         );
  MX2XL U11513 ( .A(\I_cache/cache[2][62] ), .B(n9671), .S0(n5716), .Y(n12347)
         );
  MX2XL U11514 ( .A(\I_cache/cache[1][62] ), .B(n9671), .S0(n5582), .Y(n12348)
         );
  MX2XL U11515 ( .A(\I_cache/cache[0][62] ), .B(n9671), .S0(n5617), .Y(n12349)
         );
  MX2XL U11516 ( .A(\I_cache/cache[6][61] ), .B(n3610), .S0(n5885), .Y(n12351)
         );
  MX2XL U11517 ( .A(\I_cache/cache[5][61] ), .B(n3610), .S0(n5753), .Y(n12352)
         );
  MX2XL U11518 ( .A(\I_cache/cache[4][61] ), .B(n3610), .S0(n5798), .Y(n12353)
         );
  MX2XL U11519 ( .A(\I_cache/cache[3][61] ), .B(n3610), .S0(n5663), .Y(n12354)
         );
  MX2XL U11520 ( .A(\I_cache/cache[2][61] ), .B(n3610), .S0(n5708), .Y(n12355)
         );
  MX2XL U11521 ( .A(\I_cache/cache[1][61] ), .B(n3610), .S0(n5574), .Y(n12356)
         );
  MX2XL U11522 ( .A(\I_cache/cache[0][61] ), .B(n3610), .S0(n5617), .Y(n12357)
         );
  MX2XL U11523 ( .A(\I_cache/cache[6][60] ), .B(n9641), .S0(n5887), .Y(n12359)
         );
  MX2XL U11524 ( .A(\I_cache/cache[5][60] ), .B(n9641), .S0(n5753), .Y(n12360)
         );
  MX2XL U11525 ( .A(\I_cache/cache[4][60] ), .B(n9641), .S0(n5798), .Y(n12361)
         );
  MX2XL U11526 ( .A(\I_cache/cache[3][60] ), .B(n9641), .S0(n5663), .Y(n12362)
         );
  MX2XL U11527 ( .A(\I_cache/cache[2][60] ), .B(n9641), .S0(n5709), .Y(n12363)
         );
  MX2XL U11528 ( .A(\I_cache/cache[1][60] ), .B(n9641), .S0(n5575), .Y(n12364)
         );
  MX2XL U11529 ( .A(\I_cache/cache[0][60] ), .B(n9641), .S0(n5620), .Y(n12365)
         );
  MX2XL U11530 ( .A(\I_cache/cache[6][59] ), .B(n9619), .S0(n5887), .Y(n12367)
         );
  MX2XL U11531 ( .A(\I_cache/cache[5][59] ), .B(n9619), .S0(n5753), .Y(n12368)
         );
  MX2XL U11532 ( .A(\I_cache/cache[4][59] ), .B(n9619), .S0(n5803), .Y(n12369)
         );
  MX2XL U11533 ( .A(\I_cache/cache[3][59] ), .B(n9619), .S0(n5664), .Y(n12370)
         );
  MX2XL U11534 ( .A(\I_cache/cache[2][59] ), .B(n9619), .S0(n5709), .Y(n12371)
         );
  MX2XL U11535 ( .A(\I_cache/cache[1][59] ), .B(n9619), .S0(n5575), .Y(n12372)
         );
  MX2XL U11536 ( .A(\I_cache/cache[0][59] ), .B(n9619), .S0(n5621), .Y(n12373)
         );
  MX2XL U11537 ( .A(\I_cache/cache[6][58] ), .B(n6597), .S0(n5891), .Y(n12375)
         );
  MX2XL U11538 ( .A(\I_cache/cache[5][58] ), .B(n6597), .S0(n5757), .Y(n12376)
         );
  MX2XL U11539 ( .A(\I_cache/cache[4][58] ), .B(n6597), .S0(n5804), .Y(n12377)
         );
  MX2XL U11540 ( .A(\I_cache/cache[3][58] ), .B(n6597), .S0(n5669), .Y(n12378)
         );
  MX2XL U11541 ( .A(\I_cache/cache[2][58] ), .B(n6597), .S0(n5714), .Y(n12379)
         );
  MX2XL U11542 ( .A(\I_cache/cache[1][58] ), .B(n6597), .S0(n5575), .Y(n12380)
         );
  MX2XL U11543 ( .A(\I_cache/cache[0][58] ), .B(n6597), .S0(n5624), .Y(n12381)
         );
  MX2XL U11544 ( .A(\I_cache/cache[6][57] ), .B(n10038), .S0(n5888), .Y(n12383) );
  MX2XL U11545 ( .A(\I_cache/cache[5][57] ), .B(n10038), .S0(n5754), .Y(n12384) );
  MX2XL U11546 ( .A(\I_cache/cache[4][57] ), .B(n10038), .S0(n5800), .Y(n12385) );
  MX2XL U11547 ( .A(\I_cache/cache[3][57] ), .B(n10038), .S0(n5665), .Y(n12386) );
  MX2XL U11548 ( .A(\I_cache/cache[2][57] ), .B(n10038), .S0(n5710), .Y(n12387) );
  MX2XL U11549 ( .A(\I_cache/cache[1][57] ), .B(n10038), .S0(n5576), .Y(n12388) );
  MX2XL U11550 ( .A(\I_cache/cache[0][57] ), .B(n10038), .S0(n5619), .Y(n12389) );
  MX2XL U11551 ( .A(\I_cache/cache[6][55] ), .B(n10016), .S0(n5888), .Y(n12399) );
  MX2XL U11552 ( .A(\I_cache/cache[5][55] ), .B(n10016), .S0(n5754), .Y(n12400) );
  MX2XL U11553 ( .A(\I_cache/cache[4][55] ), .B(n10016), .S0(n5800), .Y(n12401) );
  MX2XL U11554 ( .A(\I_cache/cache[3][55] ), .B(n10016), .S0(n5665), .Y(n12402) );
  MX2XL U11555 ( .A(\I_cache/cache[2][55] ), .B(n10016), .S0(n5710), .Y(n12403) );
  MX2XL U11556 ( .A(\I_cache/cache[1][55] ), .B(n10016), .S0(n5576), .Y(n12404) );
  MX2XL U11557 ( .A(\I_cache/cache[0][55] ), .B(n10016), .S0(n5619), .Y(n12405) );
  MX2XL U11558 ( .A(\I_cache/cache[6][54] ), .B(n9972), .S0(n5890), .Y(n12407)
         );
  MX2XL U11559 ( .A(\I_cache/cache[5][54] ), .B(n9972), .S0(n5757), .Y(n12408)
         );
  MX2XL U11560 ( .A(\I_cache/cache[4][54] ), .B(n9972), .S0(n5803), .Y(n12409)
         );
  MX2XL U11561 ( .A(\I_cache/cache[3][54] ), .B(n9972), .S0(n5668), .Y(n12410)
         );
  MX2XL U11562 ( .A(\I_cache/cache[2][54] ), .B(n9972), .S0(n5713), .Y(n12411)
         );
  MX2XL U11563 ( .A(\I_cache/cache[1][54] ), .B(n9972), .S0(n5579), .Y(n12412)
         );
  MX2XL U11564 ( .A(\I_cache/cache[0][54] ), .B(n9972), .S0(n5622), .Y(n12413)
         );
  MX2XL U11565 ( .A(\I_cache/cache[6][53] ), .B(n9994), .S0(n5890), .Y(n12415)
         );
  MX2XL U11566 ( .A(\I_cache/cache[5][53] ), .B(n9994), .S0(n5757), .Y(n12416)
         );
  MX2XL U11567 ( .A(\I_cache/cache[4][53] ), .B(n9994), .S0(n5803), .Y(n12417)
         );
  MX2XL U11568 ( .A(\I_cache/cache[3][53] ), .B(n9994), .S0(n5668), .Y(n12418)
         );
  MX2XL U11569 ( .A(\I_cache/cache[2][53] ), .B(n9994), .S0(n5713), .Y(n12419)
         );
  MX2XL U11570 ( .A(\I_cache/cache[1][53] ), .B(n9994), .S0(n5579), .Y(n12420)
         );
  MX2XL U11571 ( .A(\I_cache/cache[0][53] ), .B(n9994), .S0(n5622), .Y(n12421)
         );
  MX2XL U11572 ( .A(\I_cache/cache[6][52] ), .B(n9783), .S0(n5886), .Y(n12423)
         );
  MX2XL U11573 ( .A(\I_cache/cache[5][52] ), .B(n9783), .S0(n5752), .Y(n12424)
         );
  MX2XL U11574 ( .A(\I_cache/cache[4][52] ), .B(n9783), .S0(n5799), .Y(n12425)
         );
  MX2XL U11575 ( .A(\I_cache/cache[3][52] ), .B(n9783), .S0(n5664), .Y(n12426)
         );
  MX2XL U11576 ( .A(\I_cache/cache[2][52] ), .B(n9783), .S0(n5712), .Y(n12427)
         );
  MX2XL U11577 ( .A(\I_cache/cache[1][52] ), .B(n9783), .S0(n5580), .Y(n12428)
         );
  MX2XL U11578 ( .A(\I_cache/cache[0][52] ), .B(n9783), .S0(n5618), .Y(n12429)
         );
  MX2XL U11579 ( .A(\I_cache/cache[6][50] ), .B(n3615), .S0(n5886), .Y(n12439)
         );
  MX2XL U11580 ( .A(\I_cache/cache[5][50] ), .B(n3615), .S0(n5752), .Y(n12440)
         );
  MX2XL U11581 ( .A(\I_cache/cache[4][50] ), .B(n3615), .S0(n5799), .Y(n12441)
         );
  MX2XL U11582 ( .A(\I_cache/cache[3][50] ), .B(n3615), .S0(n5664), .Y(n12442)
         );
  MX2XL U11583 ( .A(\I_cache/cache[2][50] ), .B(n3615), .S0(n5713), .Y(n12443)
         );
  MX2XL U11584 ( .A(\I_cache/cache[1][50] ), .B(n3615), .S0(n5582), .Y(n12444)
         );
  MX2XL U11585 ( .A(\I_cache/cache[0][50] ), .B(n3615), .S0(n5618), .Y(n12445)
         );
  MX2XL U11586 ( .A(\I_cache/cache[6][49] ), .B(n6572), .S0(n5893), .Y(n12447)
         );
  MX2XL U11587 ( .A(\I_cache/cache[5][49] ), .B(n6572), .S0(n5755), .Y(n12448)
         );
  MX2XL U11588 ( .A(\I_cache/cache[4][49] ), .B(n6572), .S0(n5806), .Y(n12449)
         );
  MX2XL U11589 ( .A(\I_cache/cache[3][49] ), .B(n6572), .S0(n5671), .Y(n12450)
         );
  MX2XL U11590 ( .A(\I_cache/cache[2][49] ), .B(n6572), .S0(n5716), .Y(n12451)
         );
  MX2XL U11591 ( .A(\I_cache/cache[1][49] ), .B(n6572), .S0(n5581), .Y(n12452)
         );
  MX2XL U11592 ( .A(\I_cache/cache[0][49] ), .B(n6572), .S0(n5620), .Y(n12453)
         );
  MX2XL U11593 ( .A(\I_cache/cache[6][48] ), .B(n3611), .S0(n5889), .Y(n12455)
         );
  MX2XL U11594 ( .A(\I_cache/cache[5][48] ), .B(n3611), .S0(n5755), .Y(n12456)
         );
  MX2XL U11595 ( .A(\I_cache/cache[4][48] ), .B(n3611), .S0(n5801), .Y(n12457)
         );
  MX2XL U11596 ( .A(\I_cache/cache[3][48] ), .B(n3611), .S0(n5666), .Y(n12458)
         );
  MX2XL U11597 ( .A(\I_cache/cache[2][48] ), .B(n3611), .S0(n5711), .Y(n12459)
         );
  MX2XL U11598 ( .A(\I_cache/cache[1][48] ), .B(n3611), .S0(n5576), .Y(n12460)
         );
  MX2XL U11599 ( .A(\I_cache/cache[0][48] ), .B(n3611), .S0(n5618), .Y(n12461)
         );
  MX2XL U11600 ( .A(\I_cache/cache[6][47] ), .B(n10062), .S0(n5888), .Y(n12463) );
  MX2XL U11601 ( .A(\I_cache/cache[5][47] ), .B(n10062), .S0(n5754), .Y(n12464) );
  MX2XL U11602 ( .A(\I_cache/cache[4][47] ), .B(n10062), .S0(n5800), .Y(n12465) );
  MX2XL U11603 ( .A(\I_cache/cache[3][47] ), .B(n10062), .S0(n5665), .Y(n12466) );
  MX2XL U11604 ( .A(\I_cache/cache[2][47] ), .B(n10062), .S0(n5710), .Y(n12467) );
  MX2XL U11605 ( .A(\I_cache/cache[1][47] ), .B(n10062), .S0(n5576), .Y(n12468) );
  MX2XL U11606 ( .A(\I_cache/cache[0][47] ), .B(n10062), .S0(n5622), .Y(n12469) );
  MX2XL U11607 ( .A(\I_cache/cache[6][44] ), .B(n10121), .S0(n5889), .Y(n12487) );
  MX2XL U11608 ( .A(\I_cache/cache[5][44] ), .B(n10121), .S0(n5755), .Y(n12488) );
  MX2XL U11609 ( .A(\I_cache/cache[4][44] ), .B(n10121), .S0(n5801), .Y(n12489) );
  MX2XL U11610 ( .A(\I_cache/cache[3][44] ), .B(n10121), .S0(n5666), .Y(n12490) );
  MX2XL U11611 ( .A(\I_cache/cache[2][44] ), .B(n10121), .S0(n5711), .Y(n12491) );
  MX2XL U11612 ( .A(\I_cache/cache[1][44] ), .B(n10121), .S0(n5577), .Y(n12492) );
  MX2XL U11613 ( .A(\I_cache/cache[0][44] ), .B(n10121), .S0(n5620), .Y(n12493) );
  MX2XL U11614 ( .A(\I_cache/cache[6][43] ), .B(n10085), .S0(n5889), .Y(n12495) );
  MX2XL U11615 ( .A(\I_cache/cache[5][43] ), .B(n10085), .S0(n5755), .Y(n12496) );
  MX2XL U11616 ( .A(\I_cache/cache[4][43] ), .B(n10085), .S0(n5801), .Y(n12497) );
  MX2XL U11617 ( .A(\I_cache/cache[3][43] ), .B(n10085), .S0(n5666), .Y(n12498) );
  MX2XL U11618 ( .A(\I_cache/cache[2][43] ), .B(n10085), .S0(n5711), .Y(n12499) );
  MX2XL U11619 ( .A(\I_cache/cache[1][43] ), .B(n10085), .S0(n5577), .Y(n12500) );
  MX2XL U11620 ( .A(\I_cache/cache[0][43] ), .B(n10085), .S0(n5620), .Y(n12501) );
  MX2XL U11621 ( .A(\I_cache/cache[6][42] ), .B(n9834), .S0(n5886), .Y(n12503)
         );
  MX2XL U11622 ( .A(\I_cache/cache[5][42] ), .B(n9834), .S0(n5752), .Y(n12504)
         );
  MX2XL U11623 ( .A(\I_cache/cache[4][42] ), .B(n9834), .S0(n5799), .Y(n12505)
         );
  MX2XL U11624 ( .A(\I_cache/cache[3][42] ), .B(n9834), .S0(n5664), .Y(n12506)
         );
  MX2XL U11625 ( .A(\I_cache/cache[2][42] ), .B(n9834), .S0(n5711), .Y(n12507)
         );
  MX2XL U11626 ( .A(\I_cache/cache[1][42] ), .B(n9834), .S0(n5581), .Y(n12508)
         );
  MX2XL U11627 ( .A(\I_cache/cache[0][42] ), .B(n9834), .S0(n5621), .Y(n12509)
         );
  MX2XL U11628 ( .A(\I_cache/cache[6][41] ), .B(n9878), .S0(n5887), .Y(n12511)
         );
  MX2XL U11629 ( .A(\I_cache/cache[5][41] ), .B(n9878), .S0(n5756), .Y(n12512)
         );
  MX2XL U11630 ( .A(\I_cache/cache[4][41] ), .B(n9878), .S0(n5802), .Y(n12513)
         );
  MX2XL U11631 ( .A(\I_cache/cache[3][41] ), .B(n9878), .S0(n5667), .Y(n12514)
         );
  MX2XL U11632 ( .A(\I_cache/cache[2][41] ), .B(n9878), .S0(n5712), .Y(n12515)
         );
  MX2XL U11633 ( .A(\I_cache/cache[1][41] ), .B(n9878), .S0(n5578), .Y(n12516)
         );
  MX2XL U11634 ( .A(\I_cache/cache[0][41] ), .B(n9878), .S0(n5621), .Y(n12517)
         );
  MX2XL U11635 ( .A(\I_cache/cache[6][40] ), .B(n9856), .S0(n5889), .Y(n12519)
         );
  MX2XL U11636 ( .A(\I_cache/cache[5][40] ), .B(n9856), .S0(n5756), .Y(n12520)
         );
  MX2XL U11637 ( .A(\I_cache/cache[4][40] ), .B(n9856), .S0(n5802), .Y(n12521)
         );
  MX2XL U11638 ( .A(\I_cache/cache[3][40] ), .B(n9856), .S0(n5667), .Y(n12522)
         );
  MX2XL U11639 ( .A(\I_cache/cache[2][40] ), .B(n9856), .S0(n5712), .Y(n12523)
         );
  MX2XL U11640 ( .A(\I_cache/cache[1][40] ), .B(n9856), .S0(n5578), .Y(n12524)
         );
  MX2XL U11641 ( .A(\I_cache/cache[0][40] ), .B(n9856), .S0(n5621), .Y(n12525)
         );
  MX2XL U11642 ( .A(\I_cache/cache[6][39] ), .B(n9900), .S0(n5885), .Y(n12527)
         );
  MX2XL U11643 ( .A(\I_cache/cache[5][39] ), .B(n9900), .S0(n5756), .Y(n12528)
         );
  MX2XL U11644 ( .A(\I_cache/cache[4][39] ), .B(n9900), .S0(n5802), .Y(n12529)
         );
  MX2XL U11645 ( .A(\I_cache/cache[3][39] ), .B(n9900), .S0(n5667), .Y(n12530)
         );
  MX2XL U11646 ( .A(\I_cache/cache[2][39] ), .B(n9900), .S0(n5712), .Y(n12531)
         );
  MX2XL U11647 ( .A(\I_cache/cache[1][39] ), .B(n9900), .S0(n5578), .Y(n12532)
         );
  MX2XL U11648 ( .A(\I_cache/cache[0][39] ), .B(n9900), .S0(n5620), .Y(n12533)
         );
  MX2XL U11649 ( .A(\I_cache/cache[6][38] ), .B(n9922), .S0(n5890), .Y(n12535)
         );
  MX2XL U11650 ( .A(\I_cache/cache[5][38] ), .B(n9922), .S0(n5757), .Y(n12536)
         );
  MX2XL U11651 ( .A(\I_cache/cache[4][38] ), .B(n9922), .S0(n5803), .Y(n12537)
         );
  MX2XL U11652 ( .A(\I_cache/cache[3][38] ), .B(n9922), .S0(n5668), .Y(n12538)
         );
  MX2XL U11653 ( .A(\I_cache/cache[2][38] ), .B(n9922), .S0(n5713), .Y(n12539)
         );
  MX2XL U11654 ( .A(\I_cache/cache[1][38] ), .B(n9922), .S0(n5579), .Y(n12540)
         );
  MX2XL U11655 ( .A(\I_cache/cache[0][38] ), .B(n9922), .S0(n5622), .Y(n12541)
         );
  MX2XL U11656 ( .A(\I_cache/cache[6][37] ), .B(n3607), .S0(n5885), .Y(n12543)
         );
  MX2XL U11657 ( .A(\I_cache/cache[5][37] ), .B(n3607), .S0(n5756), .Y(n12544)
         );
  MX2XL U11658 ( .A(\I_cache/cache[4][37] ), .B(n3607), .S0(n5798), .Y(n12545)
         );
  MX2XL U11659 ( .A(\I_cache/cache[3][37] ), .B(n3607), .S0(n5663), .Y(n12546)
         );
  MX2XL U11660 ( .A(\I_cache/cache[2][37] ), .B(n3607), .S0(n5708), .Y(n12547)
         );
  MX2XL U11661 ( .A(\I_cache/cache[1][37] ), .B(n3607), .S0(n5574), .Y(n12548)
         );
  MX2XL U11662 ( .A(\I_cache/cache[0][37] ), .B(n3607), .S0(n5617), .Y(n12549)
         );
  MX2XL U11663 ( .A(\I_cache/cache[6][32] ), .B(n6557), .S0(n5891), .Y(n12583)
         );
  MX2XL U11664 ( .A(\I_cache/cache[5][32] ), .B(n6557), .S0(n5756), .Y(n12584)
         );
  MX2XL U11665 ( .A(\I_cache/cache[4][32] ), .B(n6557), .S0(n5804), .Y(n12585)
         );
  MX2XL U11666 ( .A(\I_cache/cache[3][32] ), .B(n6557), .S0(n5669), .Y(n12586)
         );
  MX2XL U11667 ( .A(\I_cache/cache[2][32] ), .B(n6557), .S0(n5714), .Y(n12587)
         );
  MX2XL U11668 ( .A(\I_cache/cache[1][32] ), .B(n6557), .S0(n5580), .Y(n12588)
         );
  MX2XL U11669 ( .A(\I_cache/cache[0][32] ), .B(n6557), .S0(n5622), .Y(n12589)
         );
  MX2XL U11670 ( .A(\I_cache/cache[6][89] ), .B(n10033), .S0(n5888), .Y(n12127) );
  MX2XL U11671 ( .A(\I_cache/cache[5][89] ), .B(n10033), .S0(n5754), .Y(n12128) );
  MX2XL U11672 ( .A(\I_cache/cache[4][89] ), .B(n10033), .S0(n5800), .Y(n12129) );
  MX2XL U11673 ( .A(\I_cache/cache[3][89] ), .B(n10033), .S0(n5665), .Y(n12130) );
  MX2XL U11674 ( .A(\I_cache/cache[2][89] ), .B(n10033), .S0(n5710), .Y(n12131) );
  MX2XL U11675 ( .A(\I_cache/cache[1][89] ), .B(n10033), .S0(n5576), .Y(n12132) );
  MX2XL U11676 ( .A(\I_cache/cache[0][89] ), .B(n10033), .S0(n5619), .Y(n12133) );
  MX2XL U11677 ( .A(\I_cache/cache[6][83] ), .B(n11074), .S0(n5891), .Y(n12175) );
  MX2XL U11678 ( .A(\I_cache/cache[5][83] ), .B(n11074), .S0(n5758), .Y(n12176) );
  MX2XL U11679 ( .A(\I_cache/cache[4][83] ), .B(n11074), .S0(n5804), .Y(n12177) );
  MX2XL U11680 ( .A(\I_cache/cache[3][83] ), .B(n11074), .S0(n5669), .Y(n12178) );
  MX2XL U11681 ( .A(\I_cache/cache[2][83] ), .B(n11074), .S0(n5714), .Y(n12179) );
  MX2XL U11682 ( .A(\I_cache/cache[1][83] ), .B(n11074), .S0(n5580), .Y(n12180) );
  MX2XL U11683 ( .A(\I_cache/cache[0][83] ), .B(n11074), .S0(n5623), .Y(n12181) );
  MX2XL U11684 ( .A(\I_cache/cache[6][78] ), .B(n10236), .S0(n5888), .Y(n12215) );
  MX2XL U11685 ( .A(\I_cache/cache[5][78] ), .B(n10236), .S0(n5754), .Y(n12216) );
  MX2XL U11686 ( .A(\I_cache/cache[4][78] ), .B(n10236), .S0(n5800), .Y(n12217) );
  MX2XL U11687 ( .A(\I_cache/cache[3][78] ), .B(n10236), .S0(n5665), .Y(n12218) );
  MX2XL U11688 ( .A(\I_cache/cache[2][78] ), .B(n10236), .S0(n5710), .Y(n12219) );
  MX2XL U11689 ( .A(\I_cache/cache[1][78] ), .B(n10236), .S0(n5576), .Y(n12220) );
  MX2XL U11690 ( .A(\I_cache/cache[0][78] ), .B(n10236), .S0(n5625), .Y(n12221) );
  MX2XL U11691 ( .A(\I_cache/cache[6][77] ), .B(n10214), .S0(n5889), .Y(n12223) );
  MX2XL U11692 ( .A(\I_cache/cache[5][77] ), .B(n10214), .S0(n5755), .Y(n12224) );
  MX2XL U11693 ( .A(\I_cache/cache[4][77] ), .B(n10214), .S0(n5801), .Y(n12225) );
  MX2XL U11694 ( .A(\I_cache/cache[3][77] ), .B(n10214), .S0(n5666), .Y(n12226) );
  MX2XL U11695 ( .A(\I_cache/cache[2][77] ), .B(n10214), .S0(n5711), .Y(n12227) );
  MX2XL U11696 ( .A(\I_cache/cache[1][77] ), .B(n10214), .S0(n5577), .Y(n12228) );
  MX2XL U11697 ( .A(\I_cache/cache[0][77] ), .B(n10214), .S0(n5620), .Y(n12229) );
  MX2XL U11698 ( .A(\I_cache/cache[6][76] ), .B(n10116), .S0(n5889), .Y(n12231) );
  MX2XL U11699 ( .A(\I_cache/cache[5][76] ), .B(n10116), .S0(n5755), .Y(n12232) );
  MX2XL U11700 ( .A(\I_cache/cache[4][76] ), .B(n10116), .S0(n5801), .Y(n12233) );
  MX2XL U11701 ( .A(\I_cache/cache[3][76] ), .B(n10116), .S0(n5666), .Y(n12234) );
  MX2XL U11702 ( .A(\I_cache/cache[2][76] ), .B(n10116), .S0(n5711), .Y(n12235) );
  MX2XL U11703 ( .A(\I_cache/cache[1][76] ), .B(n10116), .S0(n5577), .Y(n12236) );
  MX2XL U11704 ( .A(\I_cache/cache[0][76] ), .B(n10116), .S0(n5620), .Y(n12237) );
  MX2XL U11705 ( .A(\I_cache/cache[6][75] ), .B(n10080), .S0(n5887), .Y(n12239) );
  MX2XL U11706 ( .A(\I_cache/cache[5][75] ), .B(n10080), .S0(n5753), .Y(n12240) );
  MX2XL U11707 ( .A(\I_cache/cache[4][75] ), .B(n10080), .S0(n5801), .Y(n12241) );
  MX2XL U11708 ( .A(\I_cache/cache[3][75] ), .B(n10080), .S0(n5666), .Y(n12242) );
  MX2XL U11709 ( .A(\I_cache/cache[2][75] ), .B(n10080), .S0(n5709), .Y(n12243) );
  MX2XL U11710 ( .A(\I_cache/cache[1][75] ), .B(n10080), .S0(n5577), .Y(n12244) );
  MX2XL U11711 ( .A(\I_cache/cache[0][75] ), .B(n10080), .S0(n5620), .Y(n12245) );
  MX2XL U11712 ( .A(\I_cache/cache[6][67] ), .B(n10944), .S0(n5887), .Y(n12303) );
  MX2XL U11713 ( .A(\I_cache/cache[5][67] ), .B(n10944), .S0(n4831), .Y(n12304) );
  MX2XL U11714 ( .A(\I_cache/cache[4][67] ), .B(n10944), .S0(n5803), .Y(n12305) );
  MX2XL U11715 ( .A(\I_cache/cache[3][67] ), .B(n10944), .S0(n5665), .Y(n12306) );
  MX2XL U11716 ( .A(\I_cache/cache[2][67] ), .B(n10944), .S0(n5713), .Y(n12307) );
  MX2XL U11717 ( .A(\I_cache/cache[1][67] ), .B(n10944), .S0(n5581), .Y(n12308) );
  MX2XL U11718 ( .A(\I_cache/cache[0][67] ), .B(n10944), .S0(n5624), .Y(n12309) );
  MX2XL U11719 ( .A(\I_cache/cache[6][56] ), .B(n10833), .S0(n5893), .Y(n12391) );
  MX2XL U11720 ( .A(\I_cache/cache[5][56] ), .B(n10833), .S0(n5759), .Y(n12392) );
  MX2XL U11721 ( .A(\I_cache/cache[4][56] ), .B(n10833), .S0(n5806), .Y(n12393) );
  MX2XL U11722 ( .A(\I_cache/cache[3][56] ), .B(n10833), .S0(n5671), .Y(n12394) );
  MX2XL U11723 ( .A(\I_cache/cache[2][56] ), .B(n10833), .S0(n5716), .Y(n12395) );
  MX2XL U11724 ( .A(\I_cache/cache[1][56] ), .B(n10833), .S0(n5582), .Y(n12396) );
  MX2XL U11725 ( .A(\I_cache/cache[0][56] ), .B(n10833), .S0(n5625), .Y(n12397) );
  MX2XL U11726 ( .A(\I_cache/cache[6][51] ), .B(n3614), .S0(n5891), .Y(n12431)
         );
  MX2XL U11727 ( .A(\I_cache/cache[5][51] ), .B(n3614), .S0(n5758), .Y(n12432)
         );
  MX2XL U11728 ( .A(\I_cache/cache[4][51] ), .B(n3614), .S0(n5804), .Y(n12433)
         );
  MX2XL U11729 ( .A(\I_cache/cache[3][51] ), .B(n3614), .S0(n5669), .Y(n12434)
         );
  MX2XL U11730 ( .A(\I_cache/cache[2][51] ), .B(n3614), .S0(n5714), .Y(n12435)
         );
  MX2XL U11731 ( .A(\I_cache/cache[1][51] ), .B(n3614), .S0(n5580), .Y(n12436)
         );
  MX2XL U11732 ( .A(\I_cache/cache[0][51] ), .B(n3614), .S0(n5623), .Y(n12437)
         );
  MX2XL U11733 ( .A(\I_cache/cache[6][46] ), .B(n10241), .S0(n5888), .Y(n12471) );
  MX2XL U11734 ( .A(\I_cache/cache[5][46] ), .B(n10241), .S0(n5754), .Y(n12472) );
  MX2XL U11735 ( .A(\I_cache/cache[4][46] ), .B(n10241), .S0(n5800), .Y(n12473) );
  MX2XL U11736 ( .A(\I_cache/cache[3][46] ), .B(n10241), .S0(n5665), .Y(n12474) );
  MX2XL U11737 ( .A(\I_cache/cache[2][46] ), .B(n10241), .S0(n5710), .Y(n12475) );
  MX2XL U11738 ( .A(\I_cache/cache[1][46] ), .B(n10241), .S0(n5582), .Y(n12476) );
  MX2XL U11739 ( .A(\I_cache/cache[0][46] ), .B(n10241), .S0(n5625), .Y(n12477) );
  MX2XL U11740 ( .A(\I_cache/cache[6][45] ), .B(n10219), .S0(n5889), .Y(n12479) );
  MX2XL U11741 ( .A(\I_cache/cache[5][45] ), .B(n10219), .S0(n5755), .Y(n12480) );
  MX2XL U11742 ( .A(\I_cache/cache[4][45] ), .B(n10219), .S0(n5801), .Y(n12481) );
  MX2XL U11743 ( .A(\I_cache/cache[3][45] ), .B(n10219), .S0(n5666), .Y(n12482) );
  MX2XL U11744 ( .A(\I_cache/cache[2][45] ), .B(n10219), .S0(n5711), .Y(n12483) );
  MX2XL U11745 ( .A(\I_cache/cache[1][45] ), .B(n10219), .S0(n5577), .Y(n12484) );
  MX2XL U11746 ( .A(\I_cache/cache[0][45] ), .B(n10219), .S0(n5620), .Y(n12485) );
  MX2XL U11747 ( .A(\I_cache/cache[6][36] ), .B(n10855), .S0(n5893), .Y(n12551) );
  MX2XL U11748 ( .A(\I_cache/cache[5][36] ), .B(n10855), .S0(n5759), .Y(n12552) );
  MX2XL U11749 ( .A(\I_cache/cache[4][36] ), .B(n10855), .S0(n5806), .Y(n12553) );
  MX2XL U11750 ( .A(\I_cache/cache[3][36] ), .B(n10855), .S0(n5671), .Y(n12554) );
  MX2XL U11751 ( .A(\I_cache/cache[2][36] ), .B(n10855), .S0(n5716), .Y(n12555) );
  MX2XL U11752 ( .A(\I_cache/cache[1][36] ), .B(n10855), .S0(n5582), .Y(n12556) );
  MX2XL U11753 ( .A(\I_cache/cache[0][36] ), .B(n10855), .S0(n5625), .Y(n12557) );
  MX2XL U11754 ( .A(\I_cache/cache[6][35] ), .B(n3618), .S0(n5888), .Y(n12559)
         );
  MX2XL U11755 ( .A(\I_cache/cache[5][35] ), .B(n3618), .S0(n4831), .Y(n12560)
         );
  MX2XL U11756 ( .A(\I_cache/cache[4][35] ), .B(n3618), .S0(n5801), .Y(n12561)
         );
  MX2XL U11757 ( .A(\I_cache/cache[3][35] ), .B(n3618), .S0(n5664), .Y(n12562)
         );
  MX2XL U11758 ( .A(\I_cache/cache[2][35] ), .B(n3618), .S0(n5711), .Y(n12563)
         );
  MX2XL U11759 ( .A(\I_cache/cache[1][35] ), .B(n3618), .S0(n5577), .Y(n12564)
         );
  MX2XL U11760 ( .A(\I_cache/cache[0][35] ), .B(n3618), .S0(n5623), .Y(n12565)
         );
  MX2XL U11761 ( .A(\I_cache/cache[6][34] ), .B(n3619), .S0(n5886), .Y(n12567)
         );
  MX2XL U11762 ( .A(\I_cache/cache[5][34] ), .B(n3619), .S0(n4831), .Y(n12568)
         );
  MX2XL U11763 ( .A(\I_cache/cache[4][34] ), .B(n3619), .S0(n5800), .Y(n12569)
         );
  MX2XL U11764 ( .A(\I_cache/cache[3][34] ), .B(n3619), .S0(n5666), .Y(n12570)
         );
  MX2XL U11765 ( .A(\I_cache/cache[2][34] ), .B(n3619), .S0(n5708), .Y(n12571)
         );
  MX2XL U11766 ( .A(\I_cache/cache[1][34] ), .B(n3619), .S0(n5579), .Y(n12572)
         );
  MX2XL U11767 ( .A(\I_cache/cache[0][34] ), .B(n3619), .S0(n5625), .Y(n12573)
         );
  MX2XL U11768 ( .A(\I_cache/cache[6][33] ), .B(n10878), .S0(n5893), .Y(n12575) );
  MX2XL U11769 ( .A(\I_cache/cache[5][33] ), .B(n10878), .S0(n5759), .Y(n12576) );
  MX2XL U11770 ( .A(\I_cache/cache[4][33] ), .B(n10878), .S0(n5806), .Y(n12577) );
  MX2XL U11771 ( .A(\I_cache/cache[3][33] ), .B(n10878), .S0(n5671), .Y(n12578) );
  MX2XL U11772 ( .A(\I_cache/cache[2][33] ), .B(n10878), .S0(n5716), .Y(n12579) );
  MX2XL U11773 ( .A(\I_cache/cache[1][33] ), .B(n10878), .S0(n5582), .Y(n12580) );
  MX2XL U11774 ( .A(\I_cache/cache[0][33] ), .B(n10878), .S0(n5624), .Y(n12581) );
  MX2XL U11775 ( .A(n3554), .B(n3630), .S0(n3588), .Y(\i_MIPS/n331 ) );
  MX2XL U11776 ( .A(n3550), .B(net105250), .S0(n3597), .Y(\i_MIPS/n337 ) );
  MX2XL U11777 ( .A(n10673), .B(net104884), .S0(n3593), .Y(\i_MIPS/n353 ) );
  CLKINVX1 U11778 ( .A(\i_MIPS/n230 ), .Y(n10673) );
  CLKINVX1 U11779 ( .A(\i_MIPS/n240 ), .Y(n10185) );
  MX2XL U11780 ( .A(n9939), .B(net106290), .S0(n3601), .Y(\i_MIPS/n355 ) );
  CLKINVX1 U11781 ( .A(\i_MIPS/n232 ), .Y(n9939) );
  MX2XL U11782 ( .A(n3551), .B(n4078), .S0(n3590), .Y(\i_MIPS/n343 ) );
  MX2XL U11783 ( .A(\i_MIPS/ID_EX[78] ), .B(\i_MIPS/Sign_Extend[5] ), .S0(
        n3603), .Y(\i_MIPS/n443 ) );
  CLKMX2X2 U11784 ( .A(n5520), .B(\i_MIPS/Register/register[0][31] ), .S0(
        n6015), .Y(\i_MIPS/Register/n1139 ) );
  CLKMX2X2 U11785 ( .A(n5518), .B(\i_MIPS/Register/register[0][23] ), .S0(
        n6015), .Y(\i_MIPS/Register/n1131 ) );
  CLKMX2X2 U11786 ( .A(n5526), .B(\i_MIPS/Register/register[0][13] ), .S0(
        n6015), .Y(\i_MIPS/Register/n1121 ) );
  CLKMX2X2 U11787 ( .A(n5524), .B(\i_MIPS/Register/register[0][11] ), .S0(
        n6014), .Y(\i_MIPS/Register/n1119 ) );
  CLKMX2X2 U11788 ( .A(n5516), .B(\i_MIPS/Register/register[0][7] ), .S0(n6014), .Y(\i_MIPS/Register/n1115 ) );
  CLKMX2X2 U11789 ( .A(n5522), .B(\i_MIPS/Register/register[0][0] ), .S0(
        \i_MIPS/Register/n147 ), .Y(\i_MIPS/Register/n1108 ) );
  CLKMX2X2 U11790 ( .A(n5520), .B(\i_MIPS/Register/register[1][31] ), .S0(
        n6013), .Y(\i_MIPS/Register/n1107 ) );
  CLKMX2X2 U11791 ( .A(n5518), .B(\i_MIPS/Register/register[1][23] ), .S0(
        n6013), .Y(\i_MIPS/Register/n1099 ) );
  CLKMX2X2 U11792 ( .A(n5526), .B(\i_MIPS/Register/register[1][13] ), .S0(
        n6013), .Y(\i_MIPS/Register/n1089 ) );
  CLKMX2X2 U11793 ( .A(n5524), .B(\i_MIPS/Register/register[1][11] ), .S0(
        n6012), .Y(\i_MIPS/Register/n1087 ) );
  CLKMX2X2 U11794 ( .A(n5516), .B(\i_MIPS/Register/register[1][7] ), .S0(n6012), .Y(\i_MIPS/Register/n1083 ) );
  CLKMX2X2 U11795 ( .A(n5522), .B(\i_MIPS/Register/register[1][0] ), .S0(
        \i_MIPS/Register/n146 ), .Y(\i_MIPS/Register/n1076 ) );
  CLKMX2X2 U11796 ( .A(n5520), .B(\i_MIPS/Register/register[2][31] ), .S0(
        n6011), .Y(\i_MIPS/Register/n1075 ) );
  CLKMX2X2 U11797 ( .A(n5518), .B(\i_MIPS/Register/register[2][23] ), .S0(
        n6011), .Y(\i_MIPS/Register/n1067 ) );
  CLKMX2X2 U11798 ( .A(n5526), .B(\i_MIPS/Register/register[2][13] ), .S0(
        n6011), .Y(\i_MIPS/Register/n1057 ) );
  CLKMX2X2 U11799 ( .A(n5524), .B(\i_MIPS/Register/register[2][11] ), .S0(
        n6010), .Y(\i_MIPS/Register/n1055 ) );
  CLKMX2X2 U11800 ( .A(n5516), .B(\i_MIPS/Register/register[2][7] ), .S0(n6010), .Y(\i_MIPS/Register/n1051 ) );
  CLKMX2X2 U11801 ( .A(n5522), .B(\i_MIPS/Register/register[2][0] ), .S0(
        \i_MIPS/Register/n145 ), .Y(\i_MIPS/Register/n1044 ) );
  CLKMX2X2 U11802 ( .A(n5520), .B(\i_MIPS/Register/register[3][31] ), .S0(
        n6009), .Y(\i_MIPS/Register/n1043 ) );
  CLKMX2X2 U11803 ( .A(n5518), .B(\i_MIPS/Register/register[3][23] ), .S0(
        n6009), .Y(\i_MIPS/Register/n1035 ) );
  CLKMX2X2 U11804 ( .A(n5526), .B(\i_MIPS/Register/register[3][13] ), .S0(
        n6009), .Y(\i_MIPS/Register/n1025 ) );
  CLKMX2X2 U11805 ( .A(n5524), .B(\i_MIPS/Register/register[3][11] ), .S0(
        n6008), .Y(\i_MIPS/Register/n1023 ) );
  CLKMX2X2 U11806 ( .A(n5516), .B(\i_MIPS/Register/register[3][7] ), .S0(n6008), .Y(\i_MIPS/Register/n1019 ) );
  CLKMX2X2 U11807 ( .A(n5522), .B(\i_MIPS/Register/register[3][0] ), .S0(
        \i_MIPS/Register/n144 ), .Y(\i_MIPS/Register/n1012 ) );
  CLKMX2X2 U11808 ( .A(n5520), .B(\i_MIPS/Register/register[4][31] ), .S0(
        n6007), .Y(\i_MIPS/Register/n1011 ) );
  CLKMX2X2 U11809 ( .A(n5518), .B(\i_MIPS/Register/register[4][23] ), .S0(
        n6007), .Y(\i_MIPS/Register/n1003 ) );
  CLKMX2X2 U11810 ( .A(n5526), .B(\i_MIPS/Register/register[4][13] ), .S0(
        n6007), .Y(\i_MIPS/Register/n993 ) );
  CLKMX2X2 U11811 ( .A(n5524), .B(\i_MIPS/Register/register[4][11] ), .S0(
        n6006), .Y(\i_MIPS/Register/n991 ) );
  CLKMX2X2 U11812 ( .A(n5516), .B(\i_MIPS/Register/register[4][7] ), .S0(n6006), .Y(\i_MIPS/Register/n987 ) );
  CLKMX2X2 U11813 ( .A(n5522), .B(\i_MIPS/Register/register[4][0] ), .S0(
        \i_MIPS/Register/n143 ), .Y(\i_MIPS/Register/n980 ) );
  CLKMX2X2 U11814 ( .A(n5520), .B(\i_MIPS/Register/register[5][31] ), .S0(
        n6005), .Y(\i_MIPS/Register/n979 ) );
  CLKMX2X2 U11815 ( .A(n5518), .B(\i_MIPS/Register/register[5][23] ), .S0(
        n6005), .Y(\i_MIPS/Register/n971 ) );
  CLKMX2X2 U11816 ( .A(n5526), .B(\i_MIPS/Register/register[5][13] ), .S0(
        n6005), .Y(\i_MIPS/Register/n961 ) );
  CLKMX2X2 U11817 ( .A(n5524), .B(\i_MIPS/Register/register[5][11] ), .S0(
        n6004), .Y(\i_MIPS/Register/n959 ) );
  CLKMX2X2 U11818 ( .A(n5516), .B(\i_MIPS/Register/register[5][7] ), .S0(n6004), .Y(\i_MIPS/Register/n955 ) );
  CLKMX2X2 U11819 ( .A(n5522), .B(\i_MIPS/Register/register[5][0] ), .S0(
        \i_MIPS/Register/n142 ), .Y(\i_MIPS/Register/n948 ) );
  CLKMX2X2 U11820 ( .A(n5520), .B(\i_MIPS/Register/register[6][31] ), .S0(
        n6003), .Y(\i_MIPS/Register/n947 ) );
  CLKMX2X2 U11821 ( .A(n5518), .B(\i_MIPS/Register/register[6][23] ), .S0(
        n6003), .Y(\i_MIPS/Register/n939 ) );
  CLKMX2X2 U11822 ( .A(n5526), .B(\i_MIPS/Register/register[6][13] ), .S0(
        n6003), .Y(\i_MIPS/Register/n929 ) );
  CLKMX2X2 U11823 ( .A(n5524), .B(\i_MIPS/Register/register[6][11] ), .S0(
        n6002), .Y(\i_MIPS/Register/n927 ) );
  CLKMX2X2 U11824 ( .A(n5516), .B(\i_MIPS/Register/register[6][7] ), .S0(n6002), .Y(\i_MIPS/Register/n923 ) );
  CLKMX2X2 U11825 ( .A(n5522), .B(\i_MIPS/Register/register[6][0] ), .S0(
        \i_MIPS/Register/n141 ), .Y(\i_MIPS/Register/n916 ) );
  CLKMX2X2 U11826 ( .A(n5521), .B(\i_MIPS/Register/register[7][31] ), .S0(
        n6001), .Y(\i_MIPS/Register/n915 ) );
  CLKMX2X2 U11827 ( .A(n5519), .B(\i_MIPS/Register/register[7][23] ), .S0(
        n6001), .Y(\i_MIPS/Register/n907 ) );
  CLKMX2X2 U11828 ( .A(n5527), .B(\i_MIPS/Register/register[7][13] ), .S0(
        n6001), .Y(\i_MIPS/Register/n897 ) );
  CLKMX2X2 U11829 ( .A(n5525), .B(\i_MIPS/Register/register[7][11] ), .S0(
        n6000), .Y(\i_MIPS/Register/n895 ) );
  CLKMX2X2 U11830 ( .A(n5517), .B(\i_MIPS/Register/register[7][7] ), .S0(n6000), .Y(\i_MIPS/Register/n891 ) );
  CLKMX2X2 U11831 ( .A(n5523), .B(\i_MIPS/Register/register[7][0] ), .S0(
        \i_MIPS/Register/n139 ), .Y(\i_MIPS/Register/n884 ) );
  CLKMX2X2 U11832 ( .A(n5520), .B(\i_MIPS/Register/register[8][31] ), .S0(
        n5999), .Y(\i_MIPS/Register/n883 ) );
  CLKMX2X2 U11833 ( .A(n5518), .B(\i_MIPS/Register/register[8][23] ), .S0(
        n5999), .Y(\i_MIPS/Register/n875 ) );
  CLKMX2X2 U11834 ( .A(n5526), .B(\i_MIPS/Register/register[8][13] ), .S0(
        n5999), .Y(\i_MIPS/Register/n865 ) );
  CLKMX2X2 U11835 ( .A(n5524), .B(\i_MIPS/Register/register[8][11] ), .S0(
        n5998), .Y(\i_MIPS/Register/n863 ) );
  CLKMX2X2 U11836 ( .A(n5516), .B(\i_MIPS/Register/register[8][7] ), .S0(n5998), .Y(\i_MIPS/Register/n859 ) );
  CLKMX2X2 U11837 ( .A(n5522), .B(\i_MIPS/Register/register[8][0] ), .S0(
        \i_MIPS/Register/n138 ), .Y(\i_MIPS/Register/n852 ) );
  CLKMX2X2 U11838 ( .A(n5520), .B(\i_MIPS/Register/register[9][31] ), .S0(
        n5997), .Y(\i_MIPS/Register/n851 ) );
  CLKMX2X2 U11839 ( .A(n5518), .B(\i_MIPS/Register/register[9][23] ), .S0(
        n5997), .Y(\i_MIPS/Register/n843 ) );
  CLKMX2X2 U11840 ( .A(n5526), .B(\i_MIPS/Register/register[9][13] ), .S0(
        n5997), .Y(\i_MIPS/Register/n833 ) );
  CLKMX2X2 U11841 ( .A(n5524), .B(\i_MIPS/Register/register[9][11] ), .S0(
        n5996), .Y(\i_MIPS/Register/n831 ) );
  CLKMX2X2 U11842 ( .A(n5516), .B(\i_MIPS/Register/register[9][7] ), .S0(n5996), .Y(\i_MIPS/Register/n827 ) );
  CLKMX2X2 U11843 ( .A(n5522), .B(\i_MIPS/Register/register[9][0] ), .S0(
        \i_MIPS/Register/n137 ), .Y(\i_MIPS/Register/n820 ) );
  CLKMX2X2 U11844 ( .A(n5520), .B(\i_MIPS/Register/register[10][31] ), .S0(
        n5995), .Y(\i_MIPS/Register/n819 ) );
  CLKMX2X2 U11845 ( .A(n5518), .B(\i_MIPS/Register/register[10][23] ), .S0(
        n5995), .Y(\i_MIPS/Register/n811 ) );
  CLKMX2X2 U11846 ( .A(n5526), .B(\i_MIPS/Register/register[10][13] ), .S0(
        n5995), .Y(\i_MIPS/Register/n801 ) );
  CLKMX2X2 U11847 ( .A(n5524), .B(\i_MIPS/Register/register[10][11] ), .S0(
        n5994), .Y(\i_MIPS/Register/n799 ) );
  CLKMX2X2 U11848 ( .A(n5516), .B(\i_MIPS/Register/register[10][7] ), .S0(
        n5994), .Y(\i_MIPS/Register/n795 ) );
  CLKMX2X2 U11849 ( .A(n5522), .B(\i_MIPS/Register/register[10][0] ), .S0(
        \i_MIPS/Register/n136 ), .Y(\i_MIPS/Register/n788 ) );
  CLKMX2X2 U11850 ( .A(n5521), .B(\i_MIPS/Register/register[11][31] ), .S0(
        n5993), .Y(\i_MIPS/Register/n787 ) );
  CLKMX2X2 U11851 ( .A(n5519), .B(\i_MIPS/Register/register[11][23] ), .S0(
        n5993), .Y(\i_MIPS/Register/n779 ) );
  CLKMX2X2 U11852 ( .A(n5527), .B(\i_MIPS/Register/register[11][13] ), .S0(
        n5993), .Y(\i_MIPS/Register/n769 ) );
  CLKMX2X2 U11853 ( .A(n5525), .B(\i_MIPS/Register/register[11][11] ), .S0(
        n5992), .Y(\i_MIPS/Register/n767 ) );
  CLKMX2X2 U11854 ( .A(n5517), .B(\i_MIPS/Register/register[11][7] ), .S0(
        n5992), .Y(\i_MIPS/Register/n763 ) );
  CLKMX2X2 U11855 ( .A(n5523), .B(\i_MIPS/Register/register[11][0] ), .S0(
        \i_MIPS/Register/n135 ), .Y(\i_MIPS/Register/n756 ) );
  CLKMX2X2 U11856 ( .A(n5520), .B(\i_MIPS/Register/register[12][31] ), .S0(
        n5991), .Y(\i_MIPS/Register/n755 ) );
  CLKMX2X2 U11857 ( .A(n5518), .B(\i_MIPS/Register/register[12][23] ), .S0(
        n5991), .Y(\i_MIPS/Register/n747 ) );
  CLKMX2X2 U11858 ( .A(n5526), .B(\i_MIPS/Register/register[12][13] ), .S0(
        n5991), .Y(\i_MIPS/Register/n737 ) );
  CLKMX2X2 U11859 ( .A(n5524), .B(\i_MIPS/Register/register[12][11] ), .S0(
        n5990), .Y(\i_MIPS/Register/n735 ) );
  CLKMX2X2 U11860 ( .A(n5516), .B(\i_MIPS/Register/register[12][7] ), .S0(
        n5990), .Y(\i_MIPS/Register/n731 ) );
  CLKMX2X2 U11861 ( .A(n5522), .B(\i_MIPS/Register/register[12][0] ), .S0(
        \i_MIPS/Register/n134 ), .Y(\i_MIPS/Register/n724 ) );
  CLKMX2X2 U11862 ( .A(n5520), .B(\i_MIPS/Register/register[13][31] ), .S0(
        n5989), .Y(\i_MIPS/Register/n723 ) );
  CLKMX2X2 U11863 ( .A(n5518), .B(\i_MIPS/Register/register[13][23] ), .S0(
        n5989), .Y(\i_MIPS/Register/n715 ) );
  CLKMX2X2 U11864 ( .A(n5526), .B(\i_MIPS/Register/register[13][13] ), .S0(
        n5989), .Y(\i_MIPS/Register/n705 ) );
  CLKMX2X2 U11865 ( .A(n5524), .B(\i_MIPS/Register/register[13][11] ), .S0(
        n5988), .Y(\i_MIPS/Register/n703 ) );
  CLKMX2X2 U11866 ( .A(n5516), .B(\i_MIPS/Register/register[13][7] ), .S0(
        n5988), .Y(\i_MIPS/Register/n699 ) );
  CLKMX2X2 U11867 ( .A(n5522), .B(\i_MIPS/Register/register[13][0] ), .S0(
        \i_MIPS/Register/n133 ), .Y(\i_MIPS/Register/n692 ) );
  CLKMX2X2 U11868 ( .A(n5520), .B(\i_MIPS/Register/register[14][31] ), .S0(
        n5987), .Y(\i_MIPS/Register/n691 ) );
  CLKMX2X2 U11869 ( .A(n5518), .B(\i_MIPS/Register/register[14][23] ), .S0(
        n5987), .Y(\i_MIPS/Register/n683 ) );
  CLKMX2X2 U11870 ( .A(n5526), .B(\i_MIPS/Register/register[14][13] ), .S0(
        n5987), .Y(\i_MIPS/Register/n673 ) );
  CLKMX2X2 U11871 ( .A(n5524), .B(\i_MIPS/Register/register[14][11] ), .S0(
        n5986), .Y(\i_MIPS/Register/n671 ) );
  CLKMX2X2 U11872 ( .A(n5516), .B(\i_MIPS/Register/register[14][7] ), .S0(
        n5986), .Y(\i_MIPS/Register/n667 ) );
  CLKMX2X2 U11873 ( .A(n5522), .B(\i_MIPS/Register/register[14][0] ), .S0(
        \i_MIPS/Register/n132 ), .Y(\i_MIPS/Register/n660 ) );
  CLKMX2X2 U11874 ( .A(n5521), .B(\i_MIPS/Register/register[15][31] ), .S0(
        n5985), .Y(\i_MIPS/Register/n659 ) );
  CLKMX2X2 U11875 ( .A(n5519), .B(\i_MIPS/Register/register[15][23] ), .S0(
        n5985), .Y(\i_MIPS/Register/n651 ) );
  CLKMX2X2 U11876 ( .A(n5527), .B(\i_MIPS/Register/register[15][13] ), .S0(
        n5985), .Y(\i_MIPS/Register/n641 ) );
  CLKMX2X2 U11877 ( .A(n5525), .B(\i_MIPS/Register/register[15][11] ), .S0(
        n5984), .Y(\i_MIPS/Register/n639 ) );
  CLKMX2X2 U11878 ( .A(n5517), .B(\i_MIPS/Register/register[15][7] ), .S0(
        n5984), .Y(\i_MIPS/Register/n635 ) );
  CLKMX2X2 U11879 ( .A(n5523), .B(\i_MIPS/Register/register[15][0] ), .S0(
        \i_MIPS/Register/n130 ), .Y(\i_MIPS/Register/n628 ) );
  CLKMX2X2 U11880 ( .A(n5521), .B(\i_MIPS/Register/register[16][31] ), .S0(
        n5983), .Y(\i_MIPS/Register/n627 ) );
  CLKMX2X2 U11881 ( .A(n5519), .B(\i_MIPS/Register/register[16][23] ), .S0(
        n5983), .Y(\i_MIPS/Register/n619 ) );
  CLKMX2X2 U11882 ( .A(n5527), .B(\i_MIPS/Register/register[16][13] ), .S0(
        n5983), .Y(\i_MIPS/Register/n609 ) );
  CLKMX2X2 U11883 ( .A(n5525), .B(\i_MIPS/Register/register[16][11] ), .S0(
        n5982), .Y(\i_MIPS/Register/n607 ) );
  CLKMX2X2 U11884 ( .A(n5517), .B(\i_MIPS/Register/register[16][7] ), .S0(
        n5982), .Y(\i_MIPS/Register/n603 ) );
  CLKMX2X2 U11885 ( .A(n5523), .B(\i_MIPS/Register/register[16][0] ), .S0(
        \i_MIPS/Register/n129 ), .Y(\i_MIPS/Register/n596 ) );
  CLKMX2X2 U11886 ( .A(n5521), .B(\i_MIPS/Register/register[17][31] ), .S0(
        n5981), .Y(\i_MIPS/Register/n595 ) );
  CLKMX2X2 U11887 ( .A(n5519), .B(\i_MIPS/Register/register[17][23] ), .S0(
        n5981), .Y(\i_MIPS/Register/n587 ) );
  CLKMX2X2 U11888 ( .A(n5527), .B(\i_MIPS/Register/register[17][13] ), .S0(
        n5981), .Y(\i_MIPS/Register/n577 ) );
  CLKMX2X2 U11889 ( .A(n5525), .B(\i_MIPS/Register/register[17][11] ), .S0(
        n5980), .Y(\i_MIPS/Register/n575 ) );
  CLKMX2X2 U11890 ( .A(n5517), .B(\i_MIPS/Register/register[17][7] ), .S0(
        n5980), .Y(\i_MIPS/Register/n571 ) );
  CLKMX2X2 U11891 ( .A(n5523), .B(\i_MIPS/Register/register[17][0] ), .S0(
        \i_MIPS/Register/n128 ), .Y(\i_MIPS/Register/n564 ) );
  CLKMX2X2 U11892 ( .A(n5521), .B(\i_MIPS/Register/register[18][31] ), .S0(
        n5979), .Y(\i_MIPS/Register/n563 ) );
  CLKMX2X2 U11893 ( .A(n5519), .B(\i_MIPS/Register/register[18][23] ), .S0(
        n5979), .Y(\i_MIPS/Register/n555 ) );
  CLKMX2X2 U11894 ( .A(n5527), .B(\i_MIPS/Register/register[18][13] ), .S0(
        n5979), .Y(\i_MIPS/Register/n545 ) );
  CLKMX2X2 U11895 ( .A(n5525), .B(\i_MIPS/Register/register[18][11] ), .S0(
        n5978), .Y(\i_MIPS/Register/n543 ) );
  CLKMX2X2 U11896 ( .A(n5517), .B(\i_MIPS/Register/register[18][7] ), .S0(
        n5978), .Y(\i_MIPS/Register/n539 ) );
  CLKMX2X2 U11897 ( .A(n5523), .B(\i_MIPS/Register/register[18][0] ), .S0(
        \i_MIPS/Register/n127 ), .Y(\i_MIPS/Register/n532 ) );
  CLKMX2X2 U11898 ( .A(n5520), .B(\i_MIPS/Register/register[19][31] ), .S0(
        n5976), .Y(\i_MIPS/Register/n531 ) );
  CLKMX2X2 U11899 ( .A(n5518), .B(\i_MIPS/Register/register[19][23] ), .S0(
        n5977), .Y(\i_MIPS/Register/n523 ) );
  CLKMX2X2 U11900 ( .A(n5527), .B(\i_MIPS/Register/register[19][13] ), .S0(
        n5976), .Y(\i_MIPS/Register/n513 ) );
  CLKMX2X2 U11901 ( .A(n5516), .B(\i_MIPS/Register/register[19][7] ), .S0(
        n5977), .Y(\i_MIPS/Register/n507 ) );
  CLKMX2X2 U11902 ( .A(n5522), .B(\i_MIPS/Register/register[19][0] ), .S0(
        \i_MIPS/Register/n126 ), .Y(\i_MIPS/Register/n500 ) );
  CLKMX2X2 U11903 ( .A(n5521), .B(\i_MIPS/Register/register[20][31] ), .S0(
        n5975), .Y(\i_MIPS/Register/n499 ) );
  CLKMX2X2 U11904 ( .A(n5519), .B(\i_MIPS/Register/register[20][23] ), .S0(
        n5975), .Y(\i_MIPS/Register/n491 ) );
  CLKMX2X2 U11905 ( .A(n5527), .B(\i_MIPS/Register/register[20][13] ), .S0(
        n5975), .Y(\i_MIPS/Register/n481 ) );
  CLKMX2X2 U11906 ( .A(n5525), .B(\i_MIPS/Register/register[20][11] ), .S0(
        n5974), .Y(\i_MIPS/Register/n479 ) );
  CLKMX2X2 U11907 ( .A(n5517), .B(\i_MIPS/Register/register[20][7] ), .S0(
        n5974), .Y(\i_MIPS/Register/n475 ) );
  CLKMX2X2 U11908 ( .A(n5523), .B(\i_MIPS/Register/register[20][0] ), .S0(
        \i_MIPS/Register/n125 ), .Y(\i_MIPS/Register/n468 ) );
  CLKMX2X2 U11909 ( .A(n5521), .B(\i_MIPS/Register/register[21][31] ), .S0(
        n5972), .Y(\i_MIPS/Register/n467 ) );
  CLKMX2X2 U11910 ( .A(n5519), .B(\i_MIPS/Register/register[21][23] ), .S0(
        n5973), .Y(\i_MIPS/Register/n459 ) );
  CLKMX2X2 U11911 ( .A(n5526), .B(\i_MIPS/Register/register[21][13] ), .S0(
        n5972), .Y(\i_MIPS/Register/n449 ) );
  CLKMX2X2 U11912 ( .A(n5517), .B(\i_MIPS/Register/register[21][7] ), .S0(
        n5973), .Y(\i_MIPS/Register/n443 ) );
  CLKMX2X2 U11913 ( .A(n5523), .B(\i_MIPS/Register/register[21][0] ), .S0(
        \i_MIPS/Register/n124 ), .Y(\i_MIPS/Register/n436 ) );
  CLKMX2X2 U11914 ( .A(n5521), .B(\i_MIPS/Register/register[22][31] ), .S0(
        n5971), .Y(\i_MIPS/Register/n435 ) );
  CLKMX2X2 U11915 ( .A(n5519), .B(\i_MIPS/Register/register[22][23] ), .S0(
        n5971), .Y(\i_MIPS/Register/n427 ) );
  CLKMX2X2 U11916 ( .A(n5527), .B(\i_MIPS/Register/register[22][13] ), .S0(
        n5971), .Y(\i_MIPS/Register/n417 ) );
  CLKMX2X2 U11917 ( .A(n5525), .B(\i_MIPS/Register/register[22][11] ), .S0(
        n5970), .Y(\i_MIPS/Register/n415 ) );
  CLKMX2X2 U11918 ( .A(n5517), .B(\i_MIPS/Register/register[22][7] ), .S0(
        n5970), .Y(\i_MIPS/Register/n411 ) );
  CLKMX2X2 U11919 ( .A(n5523), .B(\i_MIPS/Register/register[22][0] ), .S0(
        \i_MIPS/Register/n123 ), .Y(\i_MIPS/Register/n404 ) );
  CLKMX2X2 U11920 ( .A(n5520), .B(\i_MIPS/Register/register[23][31] ), .S0(
        n5968), .Y(\i_MIPS/Register/n403 ) );
  CLKMX2X2 U11921 ( .A(n5518), .B(\i_MIPS/Register/register[23][23] ), .S0(
        n5969), .Y(\i_MIPS/Register/n395 ) );
  CLKMX2X2 U11922 ( .A(n5527), .B(\i_MIPS/Register/register[23][13] ), .S0(
        n5968), .Y(\i_MIPS/Register/n385 ) );
  CLKMX2X2 U11923 ( .A(n5516), .B(\i_MIPS/Register/register[23][7] ), .S0(
        n5969), .Y(\i_MIPS/Register/n379 ) );
  CLKMX2X2 U11924 ( .A(n5522), .B(\i_MIPS/Register/register[23][0] ), .S0(
        \i_MIPS/Register/n121 ), .Y(\i_MIPS/Register/n372 ) );
  MXI2XL U11925 ( .A(\i_MIPS/n202 ), .B(net108323), .S0(n3597), .Y(
        \i_MIPS/n325 ) );
  MXI2XL U11926 ( .A(\i_MIPS/n236 ), .B(net108012), .S0(n3589), .Y(
        \i_MIPS/n359 ) );
  CLKMX2X2 U11927 ( .A(n5517), .B(\i_MIPS/Register/register[24][7] ), .S0(
        n5967), .Y(\i_MIPS/Register/n347 ) );
  CLKMX2X2 U11928 ( .A(n5521), .B(\i_MIPS/Register/register[25][31] ), .S0(
        n5965), .Y(\i_MIPS/Register/n339 ) );
  CLKMX2X2 U11929 ( .A(n5519), .B(\i_MIPS/Register/register[25][23] ), .S0(
        n5965), .Y(\i_MIPS/Register/n331 ) );
  CLKMX2X2 U11930 ( .A(n5527), .B(\i_MIPS/Register/register[25][13] ), .S0(
        n5965), .Y(\i_MIPS/Register/n321 ) );
  CLKMX2X2 U11931 ( .A(n5525), .B(\i_MIPS/Register/register[25][11] ), .S0(
        n5964), .Y(\i_MIPS/Register/n319 ) );
  CLKMX2X2 U11932 ( .A(n5517), .B(\i_MIPS/Register/register[25][7] ), .S0(
        n5964), .Y(\i_MIPS/Register/n315 ) );
  CLKMX2X2 U11933 ( .A(n5523), .B(\i_MIPS/Register/register[25][0] ), .S0(
        \i_MIPS/Register/n116 ), .Y(\i_MIPS/Register/n308 ) );
  CLKMX2X2 U11934 ( .A(n5527), .B(\i_MIPS/Register/register[26][13] ), .S0(
        n5963), .Y(\i_MIPS/Register/n289 ) );
  CLKMX2X2 U11935 ( .A(n5517), .B(\i_MIPS/Register/register[26][7] ), .S0(
        n5963), .Y(\i_MIPS/Register/n283 ) );
  CLKMX2X2 U11936 ( .A(n5523), .B(\i_MIPS/Register/register[26][0] ), .S0(
        n5963), .Y(\i_MIPS/Register/n276 ) );
  CLKMX2X2 U11937 ( .A(n5521), .B(\i_MIPS/Register/register[27][31] ), .S0(
        n5960), .Y(\i_MIPS/Register/n275 ) );
  CLKMX2X2 U11938 ( .A(n5519), .B(\i_MIPS/Register/register[27][23] ), .S0(
        n5961), .Y(\i_MIPS/Register/n267 ) );
  CLKMX2X2 U11939 ( .A(n5526), .B(\i_MIPS/Register/register[27][13] ), .S0(
        n5960), .Y(\i_MIPS/Register/n257 ) );
  CLKMX2X2 U11940 ( .A(n5517), .B(\i_MIPS/Register/register[27][7] ), .S0(
        n5961), .Y(\i_MIPS/Register/n251 ) );
  CLKMX2X2 U11941 ( .A(n5523), .B(\i_MIPS/Register/register[27][0] ), .S0(
        \i_MIPS/Register/n112 ), .Y(\i_MIPS/Register/n244 ) );
  CLKMX2X2 U11942 ( .A(n5519), .B(\i_MIPS/Register/register[28][23] ), .S0(
        n5959), .Y(\i_MIPS/Register/n235 ) );
  CLKMX2X2 U11943 ( .A(n5527), .B(\i_MIPS/Register/register[28][13] ), .S0(
        n5959), .Y(\i_MIPS/Register/n225 ) );
  CLKMX2X2 U11944 ( .A(n5525), .B(\i_MIPS/Register/register[28][11] ), .S0(
        n5959), .Y(\i_MIPS/Register/n223 ) );
  CLKMX2X2 U11945 ( .A(n5517), .B(\i_MIPS/Register/register[28][7] ), .S0(
        n5958), .Y(\i_MIPS/Register/n219 ) );
  CLKMX2X2 U11946 ( .A(n5523), .B(\i_MIPS/Register/register[28][0] ), .S0(
        n5958), .Y(\i_MIPS/Register/n212 ) );
  CLKMX2X2 U11947 ( .A(n5520), .B(\i_MIPS/Register/register[29][31] ), .S0(
        n5956), .Y(\i_MIPS/Register/n211 ) );
  CLKMX2X2 U11948 ( .A(n5518), .B(\i_MIPS/Register/register[29][23] ), .S0(
        n5957), .Y(\i_MIPS/Register/n203 ) );
  CLKMX2X2 U11949 ( .A(n5527), .B(\i_MIPS/Register/register[29][13] ), .S0(
        n5956), .Y(\i_MIPS/Register/n193 ) );
  CLKMX2X2 U11950 ( .A(n5516), .B(\i_MIPS/Register/register[29][7] ), .S0(
        n5957), .Y(\i_MIPS/Register/n187 ) );
  CLKMX2X2 U11951 ( .A(n5522), .B(\i_MIPS/Register/register[29][0] ), .S0(
        \i_MIPS/Register/n108 ), .Y(\i_MIPS/Register/n180 ) );
  CLKMX2X2 U11952 ( .A(n5521), .B(\i_MIPS/Register/register[30][31] ), .S0(
        n5955), .Y(\i_MIPS/Register/n179 ) );
  CLKMX2X2 U11953 ( .A(n5519), .B(\i_MIPS/Register/register[30][23] ), .S0(
        n5955), .Y(\i_MIPS/Register/n171 ) );
  CLKMX2X2 U11954 ( .A(n5527), .B(\i_MIPS/Register/register[30][13] ), .S0(
        n5955), .Y(\i_MIPS/Register/n161 ) );
  CLKMX2X2 U11955 ( .A(n5525), .B(\i_MIPS/Register/register[30][11] ), .S0(
        n5954), .Y(\i_MIPS/Register/n159 ) );
  CLKMX2X2 U11956 ( .A(n5517), .B(\i_MIPS/Register/register[30][7] ), .S0(
        n5954), .Y(\i_MIPS/Register/n155 ) );
  CLKMX2X2 U11957 ( .A(n5523), .B(\i_MIPS/Register/register[30][0] ), .S0(
        \i_MIPS/Register/n106 ), .Y(\i_MIPS/Register/n148 ) );
  CLKMX2X2 U11958 ( .A(n5525), .B(\i_MIPS/Register/register[19][11] ), .S0(
        \i_MIPS/Register/n126 ), .Y(\i_MIPS/Register/n511 ) );
  CLKMX2X2 U11959 ( .A(n5524), .B(\i_MIPS/Register/register[21][11] ), .S0(
        \i_MIPS/Register/n124 ), .Y(\i_MIPS/Register/n447 ) );
  CLKMX2X2 U11960 ( .A(n5525), .B(\i_MIPS/Register/register[23][11] ), .S0(
        \i_MIPS/Register/n121 ), .Y(\i_MIPS/Register/n383 ) );
  CLKMX2X2 U11961 ( .A(n5521), .B(\i_MIPS/Register/register[24][31] ), .S0(
        n5967), .Y(\i_MIPS/Register/n371 ) );
  CLKMX2X2 U11962 ( .A(n5519), .B(\i_MIPS/Register/register[24][23] ), .S0(
        n5967), .Y(\i_MIPS/Register/n363 ) );
  CLKMX2X2 U11963 ( .A(n5527), .B(\i_MIPS/Register/register[24][13] ), .S0(
        n5966), .Y(\i_MIPS/Register/n353 ) );
  CLKMX2X2 U11964 ( .A(n5525), .B(\i_MIPS/Register/register[24][11] ), .S0(
        n5966), .Y(\i_MIPS/Register/n351 ) );
  CLKMX2X2 U11965 ( .A(n5523), .B(\i_MIPS/Register/register[24][0] ), .S0(
        \i_MIPS/Register/n118 ), .Y(\i_MIPS/Register/n340 ) );
  CLKMX2X2 U11966 ( .A(n5521), .B(\i_MIPS/Register/register[26][31] ), .S0(
        n5962), .Y(\i_MIPS/Register/n307 ) );
  CLKMX2X2 U11967 ( .A(n5519), .B(\i_MIPS/Register/register[26][23] ), .S0(
        n5962), .Y(\i_MIPS/Register/n299 ) );
  CLKMX2X2 U11968 ( .A(n5525), .B(\i_MIPS/Register/register[26][11] ), .S0(
        \i_MIPS/Register/n114 ), .Y(\i_MIPS/Register/n287 ) );
  CLKMX2X2 U11969 ( .A(n5521), .B(\i_MIPS/Register/register[28][31] ), .S0(
        \i_MIPS/Register/n110 ), .Y(\i_MIPS/Register/n243 ) );
  CLKMX2X2 U11970 ( .A(n5524), .B(\i_MIPS/Register/register[27][11] ), .S0(
        \i_MIPS/Register/n112 ), .Y(\i_MIPS/Register/n255 ) );
  CLKMX2X2 U11971 ( .A(n5524), .B(\i_MIPS/Register/register[29][11] ), .S0(
        \i_MIPS/Register/n108 ), .Y(\i_MIPS/Register/n191 ) );
  MX2XL U11972 ( .A(n5051), .B(n1287), .S0(n3590), .Y(\i_MIPS/n441 ) );
  MX2XL U11973 ( .A(n3682), .B(n168), .S0(n3605), .Y(\i_MIPS/n444 ) );
  MX2XL U11974 ( .A(\i_MIPS/ID_EX[81] ), .B(\i_MIPS/Sign_Extend[8] ), .S0(
        n3590), .Y(\i_MIPS/n440 ) );
  MX2XL U11975 ( .A(\i_MIPS/ID_EX[84] ), .B(\i_MIPS/Sign_Extend[11] ), .S0(
        n3601), .Y(\i_MIPS/n437 ) );
  MX2XL U11976 ( .A(\i_MIPS/ID_EX[86] ), .B(\i_MIPS/Sign_Extend[13] ), .S0(
        n3597), .Y(\i_MIPS/n435 ) );
  CLKMX2X2 U11977 ( .A(n5500), .B(\i_MIPS/Register/register[0][29] ), .S0(
        n6015), .Y(\i_MIPS/Register/n1137 ) );
  CLKMX2X2 U11978 ( .A(n5497), .B(\i_MIPS/Register/register[0][28] ), .S0(
        n6015), .Y(\i_MIPS/Register/n1136 ) );
  CLKMX2X2 U11979 ( .A(n5471), .B(\i_MIPS/Register/register[0][27] ), .S0(
        n6014), .Y(\i_MIPS/Register/n1135 ) );
  CLKMX2X2 U11980 ( .A(n5480), .B(\i_MIPS/Register/register[0][26] ), .S0(
        n6015), .Y(\i_MIPS/Register/n1134 ) );
  CLKMX2X2 U11981 ( .A(n5469), .B(\i_MIPS/Register/register[0][22] ), .S0(
        n6014), .Y(\i_MIPS/Register/n1130 ) );
  CLKMX2X2 U11982 ( .A(n5492), .B(\i_MIPS/Register/register[0][21] ), .S0(
        n6015), .Y(\i_MIPS/Register/n1129 ) );
  CLKMX2X2 U11983 ( .A(n5473), .B(\i_MIPS/Register/register[0][20] ), .S0(
        n6014), .Y(\i_MIPS/Register/n1128 ) );
  CLKMX2X2 U11984 ( .A(n5466), .B(\i_MIPS/Register/register[0][19] ), .S0(
        n6014), .Y(\i_MIPS/Register/n1127 ) );
  CLKMX2X2 U11985 ( .A(n5508), .B(\i_MIPS/Register/register[0][18] ), .S0(
        n6015), .Y(\i_MIPS/Register/n1126 ) );
  CLKMX2X2 U11986 ( .A(n5505), .B(\i_MIPS/Register/register[0][17] ), .S0(
        n6015), .Y(\i_MIPS/Register/n1125 ) );
  CLKMX2X2 U11987 ( .A(n5489), .B(\i_MIPS/Register/register[0][16] ), .S0(
        n6015), .Y(\i_MIPS/Register/n1124 ) );
  CLKMX2X2 U11988 ( .A(n5482), .B(\i_MIPS/Register/register[0][15] ), .S0(
        n6015), .Y(\i_MIPS/Register/n1123 ) );
  CLKMX2X2 U11989 ( .A(n5487), .B(\i_MIPS/Register/register[0][14] ), .S0(
        n6014), .Y(\i_MIPS/Register/n1122 ) );
  CLKMX2X2 U11990 ( .A(n5484), .B(\i_MIPS/Register/register[0][12] ), .S0(
        n6015), .Y(\i_MIPS/Register/n1120 ) );
  CLKMX2X2 U11991 ( .A(n5494), .B(\i_MIPS/Register/register[0][10] ), .S0(
        n6015), .Y(\i_MIPS/Register/n1118 ) );
  CLKMX2X2 U11992 ( .A(n5502), .B(\i_MIPS/Register/register[0][9] ), .S0(n6015), .Y(\i_MIPS/Register/n1117 ) );
  CLKMX2X2 U11993 ( .A(n5511), .B(\i_MIPS/Register/register[0][8] ), .S0(n6015), .Y(\i_MIPS/Register/n1116 ) );
  CLKMX2X2 U11994 ( .A(n5455), .B(\i_MIPS/Register/register[0][6] ), .S0(n6014), .Y(\i_MIPS/Register/n1114 ) );
  CLKMX2X2 U11995 ( .A(n5226), .B(\i_MIPS/Register/register[0][4] ), .S0(n6014), .Y(\i_MIPS/Register/n1112 ) );
  CLKMX2X2 U11996 ( .A(n5195), .B(\i_MIPS/Register/register[0][3] ), .S0(n6014), .Y(\i_MIPS/Register/n1111 ) );
  CLKMX2X2 U11997 ( .A(n5463), .B(\i_MIPS/Register/register[0][2] ), .S0(n6014), .Y(\i_MIPS/Register/n1110 ) );
  CLKMX2X2 U11998 ( .A(n5513), .B(\i_MIPS/Register/register[0][1] ), .S0(n6015), .Y(\i_MIPS/Register/n1109 ) );
  CLKMX2X2 U11999 ( .A(n5500), .B(\i_MIPS/Register/register[1][29] ), .S0(
        n6013), .Y(\i_MIPS/Register/n1105 ) );
  CLKMX2X2 U12000 ( .A(n5497), .B(\i_MIPS/Register/register[1][28] ), .S0(
        n6013), .Y(\i_MIPS/Register/n1104 ) );
  CLKMX2X2 U12001 ( .A(n5471), .B(\i_MIPS/Register/register[1][27] ), .S0(
        n6012), .Y(\i_MIPS/Register/n1103 ) );
  CLKMX2X2 U12002 ( .A(n5480), .B(\i_MIPS/Register/register[1][26] ), .S0(
        n6013), .Y(\i_MIPS/Register/n1102 ) );
  CLKMX2X2 U12003 ( .A(n5469), .B(\i_MIPS/Register/register[1][22] ), .S0(
        n6012), .Y(\i_MIPS/Register/n1098 ) );
  CLKMX2X2 U12004 ( .A(n5492), .B(\i_MIPS/Register/register[1][21] ), .S0(
        n6013), .Y(\i_MIPS/Register/n1097 ) );
  CLKMX2X2 U12005 ( .A(n5473), .B(\i_MIPS/Register/register[1][20] ), .S0(
        n6012), .Y(\i_MIPS/Register/n1096 ) );
  CLKMX2X2 U12006 ( .A(n5466), .B(\i_MIPS/Register/register[1][19] ), .S0(
        n6012), .Y(\i_MIPS/Register/n1095 ) );
  CLKMX2X2 U12007 ( .A(n5508), .B(\i_MIPS/Register/register[1][18] ), .S0(
        n6013), .Y(\i_MIPS/Register/n1094 ) );
  CLKMX2X2 U12008 ( .A(n5505), .B(\i_MIPS/Register/register[1][17] ), .S0(
        n6013), .Y(\i_MIPS/Register/n1093 ) );
  CLKMX2X2 U12009 ( .A(n5489), .B(\i_MIPS/Register/register[1][16] ), .S0(
        n6013), .Y(\i_MIPS/Register/n1092 ) );
  CLKMX2X2 U12010 ( .A(n5482), .B(\i_MIPS/Register/register[1][15] ), .S0(
        n6013), .Y(\i_MIPS/Register/n1091 ) );
  CLKMX2X2 U12011 ( .A(n5487), .B(\i_MIPS/Register/register[1][14] ), .S0(
        n6012), .Y(\i_MIPS/Register/n1090 ) );
  CLKMX2X2 U12012 ( .A(n5484), .B(\i_MIPS/Register/register[1][12] ), .S0(
        n6013), .Y(\i_MIPS/Register/n1088 ) );
  CLKMX2X2 U12013 ( .A(n5494), .B(\i_MIPS/Register/register[1][10] ), .S0(
        n6013), .Y(\i_MIPS/Register/n1086 ) );
  CLKMX2X2 U12014 ( .A(n5502), .B(\i_MIPS/Register/register[1][9] ), .S0(n6013), .Y(\i_MIPS/Register/n1085 ) );
  CLKMX2X2 U12015 ( .A(n5511), .B(\i_MIPS/Register/register[1][8] ), .S0(n6013), .Y(\i_MIPS/Register/n1084 ) );
  CLKMX2X2 U12016 ( .A(n5455), .B(\i_MIPS/Register/register[1][6] ), .S0(n6012), .Y(\i_MIPS/Register/n1082 ) );
  CLKMX2X2 U12017 ( .A(n5226), .B(\i_MIPS/Register/register[1][4] ), .S0(n6012), .Y(\i_MIPS/Register/n1080 ) );
  CLKMX2X2 U12018 ( .A(n5195), .B(\i_MIPS/Register/register[1][3] ), .S0(n6012), .Y(\i_MIPS/Register/n1079 ) );
  CLKMX2X2 U12019 ( .A(n5463), .B(\i_MIPS/Register/register[1][2] ), .S0(n6012), .Y(\i_MIPS/Register/n1078 ) );
  CLKMX2X2 U12020 ( .A(n5513), .B(\i_MIPS/Register/register[1][1] ), .S0(n6013), .Y(\i_MIPS/Register/n1077 ) );
  CLKMX2X2 U12021 ( .A(n5500), .B(\i_MIPS/Register/register[2][29] ), .S0(
        n6011), .Y(\i_MIPS/Register/n1073 ) );
  CLKMX2X2 U12022 ( .A(n5497), .B(\i_MIPS/Register/register[2][28] ), .S0(
        n6011), .Y(\i_MIPS/Register/n1072 ) );
  CLKMX2X2 U12023 ( .A(n5471), .B(\i_MIPS/Register/register[2][27] ), .S0(
        n6010), .Y(\i_MIPS/Register/n1071 ) );
  CLKMX2X2 U12024 ( .A(n5480), .B(\i_MIPS/Register/register[2][26] ), .S0(
        n6011), .Y(\i_MIPS/Register/n1070 ) );
  CLKMX2X2 U12025 ( .A(n5469), .B(\i_MIPS/Register/register[2][22] ), .S0(
        n6010), .Y(\i_MIPS/Register/n1066 ) );
  CLKMX2X2 U12026 ( .A(n5492), .B(\i_MIPS/Register/register[2][21] ), .S0(
        n6011), .Y(\i_MIPS/Register/n1065 ) );
  CLKMX2X2 U12027 ( .A(n5473), .B(\i_MIPS/Register/register[2][20] ), .S0(
        n6010), .Y(\i_MIPS/Register/n1064 ) );
  CLKMX2X2 U12028 ( .A(n5466), .B(\i_MIPS/Register/register[2][19] ), .S0(
        n6010), .Y(\i_MIPS/Register/n1063 ) );
  CLKMX2X2 U12029 ( .A(n5508), .B(\i_MIPS/Register/register[2][18] ), .S0(
        n6011), .Y(\i_MIPS/Register/n1062 ) );
  CLKMX2X2 U12030 ( .A(n5505), .B(\i_MIPS/Register/register[2][17] ), .S0(
        n6011), .Y(\i_MIPS/Register/n1061 ) );
  CLKMX2X2 U12031 ( .A(n5489), .B(\i_MIPS/Register/register[2][16] ), .S0(
        n6011), .Y(\i_MIPS/Register/n1060 ) );
  CLKMX2X2 U12032 ( .A(n5482), .B(\i_MIPS/Register/register[2][15] ), .S0(
        n6011), .Y(\i_MIPS/Register/n1059 ) );
  CLKMX2X2 U12033 ( .A(n5487), .B(\i_MIPS/Register/register[2][14] ), .S0(
        n6010), .Y(\i_MIPS/Register/n1058 ) );
  CLKMX2X2 U12034 ( .A(n5484), .B(\i_MIPS/Register/register[2][12] ), .S0(
        n6011), .Y(\i_MIPS/Register/n1056 ) );
  CLKMX2X2 U12035 ( .A(n5494), .B(\i_MIPS/Register/register[2][10] ), .S0(
        n6011), .Y(\i_MIPS/Register/n1054 ) );
  CLKMX2X2 U12036 ( .A(n5502), .B(\i_MIPS/Register/register[2][9] ), .S0(n6011), .Y(\i_MIPS/Register/n1053 ) );
  CLKMX2X2 U12037 ( .A(n5511), .B(\i_MIPS/Register/register[2][8] ), .S0(n6011), .Y(\i_MIPS/Register/n1052 ) );
  CLKMX2X2 U12038 ( .A(n5455), .B(\i_MIPS/Register/register[2][6] ), .S0(n6010), .Y(\i_MIPS/Register/n1050 ) );
  CLKMX2X2 U12039 ( .A(n5226), .B(\i_MIPS/Register/register[2][4] ), .S0(n6010), .Y(\i_MIPS/Register/n1048 ) );
  CLKMX2X2 U12040 ( .A(n5195), .B(\i_MIPS/Register/register[2][3] ), .S0(n6010), .Y(\i_MIPS/Register/n1047 ) );
  CLKMX2X2 U12041 ( .A(n5463), .B(\i_MIPS/Register/register[2][2] ), .S0(n6010), .Y(\i_MIPS/Register/n1046 ) );
  CLKMX2X2 U12042 ( .A(n5513), .B(\i_MIPS/Register/register[2][1] ), .S0(n6011), .Y(\i_MIPS/Register/n1045 ) );
  CLKMX2X2 U12043 ( .A(n5500), .B(\i_MIPS/Register/register[3][29] ), .S0(
        n6009), .Y(\i_MIPS/Register/n1041 ) );
  CLKMX2X2 U12044 ( .A(n5497), .B(\i_MIPS/Register/register[3][28] ), .S0(
        n6009), .Y(\i_MIPS/Register/n1040 ) );
  CLKMX2X2 U12045 ( .A(n5471), .B(\i_MIPS/Register/register[3][27] ), .S0(
        n6008), .Y(\i_MIPS/Register/n1039 ) );
  CLKMX2X2 U12046 ( .A(n5480), .B(\i_MIPS/Register/register[3][26] ), .S0(
        n6009), .Y(\i_MIPS/Register/n1038 ) );
  CLKMX2X2 U12047 ( .A(n5469), .B(\i_MIPS/Register/register[3][22] ), .S0(
        n6008), .Y(\i_MIPS/Register/n1034 ) );
  CLKMX2X2 U12048 ( .A(n5492), .B(\i_MIPS/Register/register[3][21] ), .S0(
        n6009), .Y(\i_MIPS/Register/n1033 ) );
  CLKMX2X2 U12049 ( .A(n5473), .B(\i_MIPS/Register/register[3][20] ), .S0(
        n6008), .Y(\i_MIPS/Register/n1032 ) );
  CLKMX2X2 U12050 ( .A(n5466), .B(\i_MIPS/Register/register[3][19] ), .S0(
        n6008), .Y(\i_MIPS/Register/n1031 ) );
  CLKMX2X2 U12051 ( .A(n5508), .B(\i_MIPS/Register/register[3][18] ), .S0(
        n6009), .Y(\i_MIPS/Register/n1030 ) );
  CLKMX2X2 U12052 ( .A(n5505), .B(\i_MIPS/Register/register[3][17] ), .S0(
        n6009), .Y(\i_MIPS/Register/n1029 ) );
  CLKMX2X2 U12053 ( .A(n5489), .B(\i_MIPS/Register/register[3][16] ), .S0(
        n6009), .Y(\i_MIPS/Register/n1028 ) );
  CLKMX2X2 U12054 ( .A(n5482), .B(\i_MIPS/Register/register[3][15] ), .S0(
        n6009), .Y(\i_MIPS/Register/n1027 ) );
  CLKMX2X2 U12055 ( .A(n5487), .B(\i_MIPS/Register/register[3][14] ), .S0(
        n6008), .Y(\i_MIPS/Register/n1026 ) );
  CLKMX2X2 U12056 ( .A(n5484), .B(\i_MIPS/Register/register[3][12] ), .S0(
        n6009), .Y(\i_MIPS/Register/n1024 ) );
  CLKMX2X2 U12057 ( .A(n5494), .B(\i_MIPS/Register/register[3][10] ), .S0(
        n6009), .Y(\i_MIPS/Register/n1022 ) );
  CLKMX2X2 U12058 ( .A(n5502), .B(\i_MIPS/Register/register[3][9] ), .S0(n6009), .Y(\i_MIPS/Register/n1021 ) );
  CLKMX2X2 U12059 ( .A(n5511), .B(\i_MIPS/Register/register[3][8] ), .S0(n6009), .Y(\i_MIPS/Register/n1020 ) );
  CLKMX2X2 U12060 ( .A(n5455), .B(\i_MIPS/Register/register[3][6] ), .S0(n6008), .Y(\i_MIPS/Register/n1018 ) );
  CLKMX2X2 U12061 ( .A(n5226), .B(\i_MIPS/Register/register[3][4] ), .S0(n6008), .Y(\i_MIPS/Register/n1016 ) );
  CLKMX2X2 U12062 ( .A(n5195), .B(\i_MIPS/Register/register[3][3] ), .S0(n6008), .Y(\i_MIPS/Register/n1015 ) );
  CLKMX2X2 U12063 ( .A(n5463), .B(\i_MIPS/Register/register[3][2] ), .S0(n6008), .Y(\i_MIPS/Register/n1014 ) );
  CLKMX2X2 U12064 ( .A(n5513), .B(\i_MIPS/Register/register[3][1] ), .S0(n6009), .Y(\i_MIPS/Register/n1013 ) );
  CLKMX2X2 U12065 ( .A(n5500), .B(\i_MIPS/Register/register[4][29] ), .S0(
        n6007), .Y(\i_MIPS/Register/n1009 ) );
  CLKMX2X2 U12066 ( .A(n5497), .B(\i_MIPS/Register/register[4][28] ), .S0(
        n6007), .Y(\i_MIPS/Register/n1008 ) );
  CLKMX2X2 U12067 ( .A(n5471), .B(\i_MIPS/Register/register[4][27] ), .S0(
        n6006), .Y(\i_MIPS/Register/n1007 ) );
  CLKMX2X2 U12068 ( .A(n5480), .B(\i_MIPS/Register/register[4][26] ), .S0(
        n6007), .Y(\i_MIPS/Register/n1006 ) );
  CLKMX2X2 U12069 ( .A(n5469), .B(\i_MIPS/Register/register[4][22] ), .S0(
        n6006), .Y(\i_MIPS/Register/n1002 ) );
  CLKMX2X2 U12070 ( .A(n5492), .B(\i_MIPS/Register/register[4][21] ), .S0(
        n6007), .Y(\i_MIPS/Register/n1001 ) );
  CLKMX2X2 U12071 ( .A(n5473), .B(\i_MIPS/Register/register[4][20] ), .S0(
        n6006), .Y(\i_MIPS/Register/n1000 ) );
  CLKMX2X2 U12072 ( .A(n5466), .B(\i_MIPS/Register/register[4][19] ), .S0(
        n6006), .Y(\i_MIPS/Register/n999 ) );
  CLKMX2X2 U12073 ( .A(n5508), .B(\i_MIPS/Register/register[4][18] ), .S0(
        n6007), .Y(\i_MIPS/Register/n998 ) );
  CLKMX2X2 U12074 ( .A(n5505), .B(\i_MIPS/Register/register[4][17] ), .S0(
        n6007), .Y(\i_MIPS/Register/n997 ) );
  CLKMX2X2 U12075 ( .A(n5489), .B(\i_MIPS/Register/register[4][16] ), .S0(
        n6007), .Y(\i_MIPS/Register/n996 ) );
  CLKMX2X2 U12076 ( .A(n5482), .B(\i_MIPS/Register/register[4][15] ), .S0(
        n6007), .Y(\i_MIPS/Register/n995 ) );
  CLKMX2X2 U12077 ( .A(n5487), .B(\i_MIPS/Register/register[4][14] ), .S0(
        n6006), .Y(\i_MIPS/Register/n994 ) );
  CLKMX2X2 U12078 ( .A(n5484), .B(\i_MIPS/Register/register[4][12] ), .S0(
        n6007), .Y(\i_MIPS/Register/n992 ) );
  CLKMX2X2 U12079 ( .A(n5494), .B(\i_MIPS/Register/register[4][10] ), .S0(
        n6007), .Y(\i_MIPS/Register/n990 ) );
  CLKMX2X2 U12080 ( .A(n5502), .B(\i_MIPS/Register/register[4][9] ), .S0(n6007), .Y(\i_MIPS/Register/n989 ) );
  CLKMX2X2 U12081 ( .A(n5511), .B(\i_MIPS/Register/register[4][8] ), .S0(n6007), .Y(\i_MIPS/Register/n988 ) );
  CLKMX2X2 U12082 ( .A(n5455), .B(\i_MIPS/Register/register[4][6] ), .S0(n6006), .Y(\i_MIPS/Register/n986 ) );
  CLKMX2X2 U12083 ( .A(n5226), .B(\i_MIPS/Register/register[4][4] ), .S0(n6006), .Y(\i_MIPS/Register/n984 ) );
  CLKMX2X2 U12084 ( .A(n5195), .B(\i_MIPS/Register/register[4][3] ), .S0(n6006), .Y(\i_MIPS/Register/n983 ) );
  CLKMX2X2 U12085 ( .A(n5463), .B(\i_MIPS/Register/register[4][2] ), .S0(n6006), .Y(\i_MIPS/Register/n982 ) );
  CLKMX2X2 U12086 ( .A(n5513), .B(\i_MIPS/Register/register[4][1] ), .S0(n6007), .Y(\i_MIPS/Register/n981 ) );
  CLKMX2X2 U12087 ( .A(n5500), .B(\i_MIPS/Register/register[5][29] ), .S0(
        n6005), .Y(\i_MIPS/Register/n977 ) );
  CLKMX2X2 U12088 ( .A(n5497), .B(\i_MIPS/Register/register[5][28] ), .S0(
        n6005), .Y(\i_MIPS/Register/n976 ) );
  CLKMX2X2 U12089 ( .A(n5471), .B(\i_MIPS/Register/register[5][27] ), .S0(
        n6004), .Y(\i_MIPS/Register/n975 ) );
  CLKMX2X2 U12090 ( .A(n5480), .B(\i_MIPS/Register/register[5][26] ), .S0(
        n6005), .Y(\i_MIPS/Register/n974 ) );
  CLKMX2X2 U12091 ( .A(n5469), .B(\i_MIPS/Register/register[5][22] ), .S0(
        n6004), .Y(\i_MIPS/Register/n970 ) );
  CLKMX2X2 U12092 ( .A(n5492), .B(\i_MIPS/Register/register[5][21] ), .S0(
        n6005), .Y(\i_MIPS/Register/n969 ) );
  CLKMX2X2 U12093 ( .A(n5473), .B(\i_MIPS/Register/register[5][20] ), .S0(
        n6004), .Y(\i_MIPS/Register/n968 ) );
  CLKMX2X2 U12094 ( .A(n5466), .B(\i_MIPS/Register/register[5][19] ), .S0(
        n6004), .Y(\i_MIPS/Register/n967 ) );
  CLKMX2X2 U12095 ( .A(n5508), .B(\i_MIPS/Register/register[5][18] ), .S0(
        n6005), .Y(\i_MIPS/Register/n966 ) );
  CLKMX2X2 U12096 ( .A(n5505), .B(\i_MIPS/Register/register[5][17] ), .S0(
        n6005), .Y(\i_MIPS/Register/n965 ) );
  CLKMX2X2 U12097 ( .A(n5489), .B(\i_MIPS/Register/register[5][16] ), .S0(
        n6005), .Y(\i_MIPS/Register/n964 ) );
  CLKMX2X2 U12098 ( .A(n5482), .B(\i_MIPS/Register/register[5][15] ), .S0(
        n6005), .Y(\i_MIPS/Register/n963 ) );
  CLKMX2X2 U12099 ( .A(n5487), .B(\i_MIPS/Register/register[5][14] ), .S0(
        n6004), .Y(\i_MIPS/Register/n962 ) );
  CLKMX2X2 U12100 ( .A(n5484), .B(\i_MIPS/Register/register[5][12] ), .S0(
        n6005), .Y(\i_MIPS/Register/n960 ) );
  CLKMX2X2 U12101 ( .A(n5494), .B(\i_MIPS/Register/register[5][10] ), .S0(
        n6005), .Y(\i_MIPS/Register/n958 ) );
  CLKMX2X2 U12102 ( .A(n5502), .B(\i_MIPS/Register/register[5][9] ), .S0(n6005), .Y(\i_MIPS/Register/n957 ) );
  CLKMX2X2 U12103 ( .A(n5511), .B(\i_MIPS/Register/register[5][8] ), .S0(n6005), .Y(\i_MIPS/Register/n956 ) );
  CLKMX2X2 U12104 ( .A(n5455), .B(\i_MIPS/Register/register[5][6] ), .S0(n6004), .Y(\i_MIPS/Register/n954 ) );
  CLKMX2X2 U12105 ( .A(n5226), .B(\i_MIPS/Register/register[5][4] ), .S0(n6004), .Y(\i_MIPS/Register/n952 ) );
  CLKMX2X2 U12106 ( .A(n5195), .B(\i_MIPS/Register/register[5][3] ), .S0(n6004), .Y(\i_MIPS/Register/n951 ) );
  CLKMX2X2 U12107 ( .A(n5463), .B(\i_MIPS/Register/register[5][2] ), .S0(n6004), .Y(\i_MIPS/Register/n950 ) );
  CLKMX2X2 U12108 ( .A(n5513), .B(\i_MIPS/Register/register[5][1] ), .S0(n6005), .Y(\i_MIPS/Register/n949 ) );
  CLKMX2X2 U12109 ( .A(n5500), .B(\i_MIPS/Register/register[6][29] ), .S0(
        n6003), .Y(\i_MIPS/Register/n945 ) );
  CLKMX2X2 U12110 ( .A(n5497), .B(\i_MIPS/Register/register[6][28] ), .S0(
        n6003), .Y(\i_MIPS/Register/n944 ) );
  CLKMX2X2 U12111 ( .A(n5471), .B(\i_MIPS/Register/register[6][27] ), .S0(
        n6002), .Y(\i_MIPS/Register/n943 ) );
  CLKMX2X2 U12112 ( .A(n5480), .B(\i_MIPS/Register/register[6][26] ), .S0(
        n6003), .Y(\i_MIPS/Register/n942 ) );
  CLKMX2X2 U12113 ( .A(n5469), .B(\i_MIPS/Register/register[6][22] ), .S0(
        n6002), .Y(\i_MIPS/Register/n938 ) );
  CLKMX2X2 U12114 ( .A(n5492), .B(\i_MIPS/Register/register[6][21] ), .S0(
        n6003), .Y(\i_MIPS/Register/n937 ) );
  CLKMX2X2 U12115 ( .A(n5473), .B(\i_MIPS/Register/register[6][20] ), .S0(
        n6002), .Y(\i_MIPS/Register/n936 ) );
  CLKMX2X2 U12116 ( .A(n5466), .B(\i_MIPS/Register/register[6][19] ), .S0(
        n6002), .Y(\i_MIPS/Register/n935 ) );
  CLKMX2X2 U12117 ( .A(n5508), .B(\i_MIPS/Register/register[6][18] ), .S0(
        n6003), .Y(\i_MIPS/Register/n934 ) );
  CLKMX2X2 U12118 ( .A(n5505), .B(\i_MIPS/Register/register[6][17] ), .S0(
        n6003), .Y(\i_MIPS/Register/n933 ) );
  CLKMX2X2 U12119 ( .A(n5489), .B(\i_MIPS/Register/register[6][16] ), .S0(
        n6003), .Y(\i_MIPS/Register/n932 ) );
  CLKMX2X2 U12120 ( .A(n5482), .B(\i_MIPS/Register/register[6][15] ), .S0(
        n6003), .Y(\i_MIPS/Register/n931 ) );
  CLKMX2X2 U12121 ( .A(n5487), .B(\i_MIPS/Register/register[6][14] ), .S0(
        n6002), .Y(\i_MIPS/Register/n930 ) );
  CLKMX2X2 U12122 ( .A(n5484), .B(\i_MIPS/Register/register[6][12] ), .S0(
        n6003), .Y(\i_MIPS/Register/n928 ) );
  CLKMX2X2 U12123 ( .A(n5494), .B(\i_MIPS/Register/register[6][10] ), .S0(
        n6003), .Y(\i_MIPS/Register/n926 ) );
  CLKMX2X2 U12124 ( .A(n5502), .B(\i_MIPS/Register/register[6][9] ), .S0(n6003), .Y(\i_MIPS/Register/n925 ) );
  CLKMX2X2 U12125 ( .A(n5511), .B(\i_MIPS/Register/register[6][8] ), .S0(n6003), .Y(\i_MIPS/Register/n924 ) );
  CLKMX2X2 U12126 ( .A(n5455), .B(\i_MIPS/Register/register[6][6] ), .S0(n6002), .Y(\i_MIPS/Register/n922 ) );
  CLKMX2X2 U12127 ( .A(n5226), .B(\i_MIPS/Register/register[6][4] ), .S0(n6002), .Y(\i_MIPS/Register/n920 ) );
  CLKMX2X2 U12128 ( .A(n5195), .B(\i_MIPS/Register/register[6][3] ), .S0(n6002), .Y(\i_MIPS/Register/n919 ) );
  CLKMX2X2 U12129 ( .A(n5463), .B(\i_MIPS/Register/register[6][2] ), .S0(n6002), .Y(\i_MIPS/Register/n918 ) );
  CLKMX2X2 U12130 ( .A(n5513), .B(\i_MIPS/Register/register[6][1] ), .S0(n6003), .Y(\i_MIPS/Register/n917 ) );
  CLKMX2X2 U12131 ( .A(n5501), .B(\i_MIPS/Register/register[7][29] ), .S0(
        n6001), .Y(\i_MIPS/Register/n913 ) );
  CLKMX2X2 U12132 ( .A(n5498), .B(\i_MIPS/Register/register[7][28] ), .S0(
        n6001), .Y(\i_MIPS/Register/n912 ) );
  CLKMX2X2 U12133 ( .A(n5472), .B(\i_MIPS/Register/register[7][27] ), .S0(
        n6000), .Y(\i_MIPS/Register/n911 ) );
  CLKMX2X2 U12134 ( .A(n5481), .B(\i_MIPS/Register/register[7][26] ), .S0(
        n6001), .Y(\i_MIPS/Register/n910 ) );
  CLKMX2X2 U12135 ( .A(n5470), .B(\i_MIPS/Register/register[7][22] ), .S0(
        n6000), .Y(\i_MIPS/Register/n906 ) );
  CLKMX2X2 U12136 ( .A(n5493), .B(\i_MIPS/Register/register[7][21] ), .S0(
        n6001), .Y(\i_MIPS/Register/n905 ) );
  CLKMX2X2 U12137 ( .A(n5474), .B(\i_MIPS/Register/register[7][20] ), .S0(
        n6000), .Y(\i_MIPS/Register/n904 ) );
  CLKMX2X2 U12138 ( .A(n5467), .B(\i_MIPS/Register/register[7][19] ), .S0(
        n6000), .Y(\i_MIPS/Register/n903 ) );
  CLKMX2X2 U12139 ( .A(n5509), .B(\i_MIPS/Register/register[7][18] ), .S0(
        n6001), .Y(\i_MIPS/Register/n902 ) );
  CLKMX2X2 U12140 ( .A(n5506), .B(\i_MIPS/Register/register[7][17] ), .S0(
        n6001), .Y(\i_MIPS/Register/n901 ) );
  CLKMX2X2 U12141 ( .A(n5490), .B(\i_MIPS/Register/register[7][16] ), .S0(
        n6001), .Y(\i_MIPS/Register/n900 ) );
  CLKMX2X2 U12142 ( .A(n5483), .B(\i_MIPS/Register/register[7][15] ), .S0(
        n6001), .Y(\i_MIPS/Register/n899 ) );
  CLKMX2X2 U12143 ( .A(n5488), .B(\i_MIPS/Register/register[7][14] ), .S0(
        n6000), .Y(\i_MIPS/Register/n898 ) );
  CLKMX2X2 U12144 ( .A(n5485), .B(\i_MIPS/Register/register[7][12] ), .S0(
        n6001), .Y(\i_MIPS/Register/n896 ) );
  CLKMX2X2 U12145 ( .A(n5495), .B(\i_MIPS/Register/register[7][10] ), .S0(
        n6001), .Y(\i_MIPS/Register/n894 ) );
  CLKMX2X2 U12146 ( .A(n5503), .B(\i_MIPS/Register/register[7][9] ), .S0(n6001), .Y(\i_MIPS/Register/n893 ) );
  CLKMX2X2 U12147 ( .A(n5512), .B(\i_MIPS/Register/register[7][8] ), .S0(n6001), .Y(\i_MIPS/Register/n892 ) );
  CLKMX2X2 U12148 ( .A(n5456), .B(\i_MIPS/Register/register[7][6] ), .S0(n6000), .Y(\i_MIPS/Register/n890 ) );
  CLKMX2X2 U12149 ( .A(n5227), .B(\i_MIPS/Register/register[7][4] ), .S0(n6000), .Y(\i_MIPS/Register/n888 ) );
  CLKMX2X2 U12150 ( .A(n5196), .B(\i_MIPS/Register/register[7][3] ), .S0(n6000), .Y(\i_MIPS/Register/n887 ) );
  CLKMX2X2 U12151 ( .A(n5464), .B(\i_MIPS/Register/register[7][2] ), .S0(n6000), .Y(\i_MIPS/Register/n886 ) );
  CLKMX2X2 U12152 ( .A(n5514), .B(\i_MIPS/Register/register[7][1] ), .S0(n6001), .Y(\i_MIPS/Register/n885 ) );
  CLKMX2X2 U12153 ( .A(n5500), .B(\i_MIPS/Register/register[8][29] ), .S0(
        n5999), .Y(\i_MIPS/Register/n881 ) );
  CLKMX2X2 U12154 ( .A(n5497), .B(\i_MIPS/Register/register[8][28] ), .S0(
        n5999), .Y(\i_MIPS/Register/n880 ) );
  CLKMX2X2 U12155 ( .A(n5471), .B(\i_MIPS/Register/register[8][27] ), .S0(
        n5998), .Y(\i_MIPS/Register/n879 ) );
  CLKMX2X2 U12156 ( .A(n5480), .B(\i_MIPS/Register/register[8][26] ), .S0(
        n5999), .Y(\i_MIPS/Register/n878 ) );
  CLKMX2X2 U12157 ( .A(n5469), .B(\i_MIPS/Register/register[8][22] ), .S0(
        n5998), .Y(\i_MIPS/Register/n874 ) );
  CLKMX2X2 U12158 ( .A(n5492), .B(\i_MIPS/Register/register[8][21] ), .S0(
        n5999), .Y(\i_MIPS/Register/n873 ) );
  CLKMX2X2 U12159 ( .A(n5473), .B(\i_MIPS/Register/register[8][20] ), .S0(
        n5998), .Y(\i_MIPS/Register/n872 ) );
  CLKMX2X2 U12160 ( .A(n5466), .B(\i_MIPS/Register/register[8][19] ), .S0(
        n5998), .Y(\i_MIPS/Register/n871 ) );
  CLKMX2X2 U12161 ( .A(n5508), .B(\i_MIPS/Register/register[8][18] ), .S0(
        n5999), .Y(\i_MIPS/Register/n870 ) );
  CLKMX2X2 U12162 ( .A(n5505), .B(\i_MIPS/Register/register[8][17] ), .S0(
        n5999), .Y(\i_MIPS/Register/n869 ) );
  CLKMX2X2 U12163 ( .A(n5489), .B(\i_MIPS/Register/register[8][16] ), .S0(
        n5999), .Y(\i_MIPS/Register/n868 ) );
  CLKMX2X2 U12164 ( .A(n5482), .B(\i_MIPS/Register/register[8][15] ), .S0(
        n5999), .Y(\i_MIPS/Register/n867 ) );
  CLKMX2X2 U12165 ( .A(n5487), .B(\i_MIPS/Register/register[8][14] ), .S0(
        n5998), .Y(\i_MIPS/Register/n866 ) );
  CLKMX2X2 U12166 ( .A(n5484), .B(\i_MIPS/Register/register[8][12] ), .S0(
        n5999), .Y(\i_MIPS/Register/n864 ) );
  CLKMX2X2 U12167 ( .A(n5494), .B(\i_MIPS/Register/register[8][10] ), .S0(
        n5999), .Y(\i_MIPS/Register/n862 ) );
  CLKMX2X2 U12168 ( .A(n5502), .B(\i_MIPS/Register/register[8][9] ), .S0(n5999), .Y(\i_MIPS/Register/n861 ) );
  CLKMX2X2 U12169 ( .A(n5511), .B(\i_MIPS/Register/register[8][8] ), .S0(n5999), .Y(\i_MIPS/Register/n860 ) );
  CLKMX2X2 U12170 ( .A(n5455), .B(\i_MIPS/Register/register[8][6] ), .S0(n5998), .Y(\i_MIPS/Register/n858 ) );
  CLKMX2X2 U12171 ( .A(n5226), .B(\i_MIPS/Register/register[8][4] ), .S0(n5998), .Y(\i_MIPS/Register/n856 ) );
  CLKMX2X2 U12172 ( .A(n5195), .B(\i_MIPS/Register/register[8][3] ), .S0(n5998), .Y(\i_MIPS/Register/n855 ) );
  CLKMX2X2 U12173 ( .A(n5463), .B(\i_MIPS/Register/register[8][2] ), .S0(n5998), .Y(\i_MIPS/Register/n854 ) );
  CLKMX2X2 U12174 ( .A(n5513), .B(\i_MIPS/Register/register[8][1] ), .S0(n5999), .Y(\i_MIPS/Register/n853 ) );
  CLKMX2X2 U12175 ( .A(n5500), .B(\i_MIPS/Register/register[9][29] ), .S0(
        n5997), .Y(\i_MIPS/Register/n849 ) );
  CLKMX2X2 U12176 ( .A(n5497), .B(\i_MIPS/Register/register[9][28] ), .S0(
        n5997), .Y(\i_MIPS/Register/n848 ) );
  CLKMX2X2 U12177 ( .A(n5471), .B(\i_MIPS/Register/register[9][27] ), .S0(
        n5996), .Y(\i_MIPS/Register/n847 ) );
  CLKMX2X2 U12178 ( .A(n5480), .B(\i_MIPS/Register/register[9][26] ), .S0(
        n5997), .Y(\i_MIPS/Register/n846 ) );
  CLKMX2X2 U12179 ( .A(n5469), .B(\i_MIPS/Register/register[9][22] ), .S0(
        n5996), .Y(\i_MIPS/Register/n842 ) );
  CLKMX2X2 U12180 ( .A(n5492), .B(\i_MIPS/Register/register[9][21] ), .S0(
        n5997), .Y(\i_MIPS/Register/n841 ) );
  CLKMX2X2 U12181 ( .A(n5473), .B(\i_MIPS/Register/register[9][20] ), .S0(
        n5996), .Y(\i_MIPS/Register/n840 ) );
  CLKMX2X2 U12182 ( .A(n5466), .B(\i_MIPS/Register/register[9][19] ), .S0(
        n5996), .Y(\i_MIPS/Register/n839 ) );
  CLKMX2X2 U12183 ( .A(n5508), .B(\i_MIPS/Register/register[9][18] ), .S0(
        n5997), .Y(\i_MIPS/Register/n838 ) );
  CLKMX2X2 U12184 ( .A(n5505), .B(\i_MIPS/Register/register[9][17] ), .S0(
        n5997), .Y(\i_MIPS/Register/n837 ) );
  CLKMX2X2 U12185 ( .A(n5489), .B(\i_MIPS/Register/register[9][16] ), .S0(
        n5997), .Y(\i_MIPS/Register/n836 ) );
  CLKMX2X2 U12186 ( .A(n5482), .B(\i_MIPS/Register/register[9][15] ), .S0(
        n5997), .Y(\i_MIPS/Register/n835 ) );
  CLKMX2X2 U12187 ( .A(n5487), .B(\i_MIPS/Register/register[9][14] ), .S0(
        n5996), .Y(\i_MIPS/Register/n834 ) );
  CLKMX2X2 U12188 ( .A(n5484), .B(\i_MIPS/Register/register[9][12] ), .S0(
        n5997), .Y(\i_MIPS/Register/n832 ) );
  CLKMX2X2 U12189 ( .A(n5494), .B(\i_MIPS/Register/register[9][10] ), .S0(
        n5997), .Y(\i_MIPS/Register/n830 ) );
  CLKMX2X2 U12190 ( .A(n5502), .B(\i_MIPS/Register/register[9][9] ), .S0(n5997), .Y(\i_MIPS/Register/n829 ) );
  CLKMX2X2 U12191 ( .A(n5511), .B(\i_MIPS/Register/register[9][8] ), .S0(n5997), .Y(\i_MIPS/Register/n828 ) );
  CLKMX2X2 U12192 ( .A(n5455), .B(\i_MIPS/Register/register[9][6] ), .S0(n5996), .Y(\i_MIPS/Register/n826 ) );
  CLKMX2X2 U12193 ( .A(n5226), .B(\i_MIPS/Register/register[9][4] ), .S0(n5996), .Y(\i_MIPS/Register/n824 ) );
  CLKMX2X2 U12194 ( .A(n5195), .B(\i_MIPS/Register/register[9][3] ), .S0(n5996), .Y(\i_MIPS/Register/n823 ) );
  CLKMX2X2 U12195 ( .A(n5463), .B(\i_MIPS/Register/register[9][2] ), .S0(n5996), .Y(\i_MIPS/Register/n822 ) );
  CLKMX2X2 U12196 ( .A(n5513), .B(\i_MIPS/Register/register[9][1] ), .S0(n5997), .Y(\i_MIPS/Register/n821 ) );
  CLKMX2X2 U12197 ( .A(n5500), .B(\i_MIPS/Register/register[10][29] ), .S0(
        n5995), .Y(\i_MIPS/Register/n817 ) );
  CLKMX2X2 U12198 ( .A(n5497), .B(\i_MIPS/Register/register[10][28] ), .S0(
        n5995), .Y(\i_MIPS/Register/n816 ) );
  CLKMX2X2 U12199 ( .A(n5471), .B(\i_MIPS/Register/register[10][27] ), .S0(
        n5994), .Y(\i_MIPS/Register/n815 ) );
  CLKMX2X2 U12200 ( .A(n5480), .B(\i_MIPS/Register/register[10][26] ), .S0(
        n5995), .Y(\i_MIPS/Register/n814 ) );
  CLKMX2X2 U12201 ( .A(n5469), .B(\i_MIPS/Register/register[10][22] ), .S0(
        n5994), .Y(\i_MIPS/Register/n810 ) );
  CLKMX2X2 U12202 ( .A(n5492), .B(\i_MIPS/Register/register[10][21] ), .S0(
        n5995), .Y(\i_MIPS/Register/n809 ) );
  CLKMX2X2 U12203 ( .A(n5473), .B(\i_MIPS/Register/register[10][20] ), .S0(
        n5994), .Y(\i_MIPS/Register/n808 ) );
  CLKMX2X2 U12204 ( .A(n5466), .B(\i_MIPS/Register/register[10][19] ), .S0(
        n5994), .Y(\i_MIPS/Register/n807 ) );
  CLKMX2X2 U12205 ( .A(n5508), .B(\i_MIPS/Register/register[10][18] ), .S0(
        n5995), .Y(\i_MIPS/Register/n806 ) );
  CLKMX2X2 U12206 ( .A(n5505), .B(\i_MIPS/Register/register[10][17] ), .S0(
        n5995), .Y(\i_MIPS/Register/n805 ) );
  CLKMX2X2 U12207 ( .A(n5489), .B(\i_MIPS/Register/register[10][16] ), .S0(
        n5995), .Y(\i_MIPS/Register/n804 ) );
  CLKMX2X2 U12208 ( .A(n5482), .B(\i_MIPS/Register/register[10][15] ), .S0(
        n5995), .Y(\i_MIPS/Register/n803 ) );
  CLKMX2X2 U12209 ( .A(n5487), .B(\i_MIPS/Register/register[10][14] ), .S0(
        n5994), .Y(\i_MIPS/Register/n802 ) );
  CLKMX2X2 U12210 ( .A(n5484), .B(\i_MIPS/Register/register[10][12] ), .S0(
        n5995), .Y(\i_MIPS/Register/n800 ) );
  CLKMX2X2 U12211 ( .A(n5494), .B(\i_MIPS/Register/register[10][10] ), .S0(
        n5995), .Y(\i_MIPS/Register/n798 ) );
  CLKMX2X2 U12212 ( .A(n5502), .B(\i_MIPS/Register/register[10][9] ), .S0(
        n5995), .Y(\i_MIPS/Register/n797 ) );
  CLKMX2X2 U12213 ( .A(n5511), .B(\i_MIPS/Register/register[10][8] ), .S0(
        n5995), .Y(\i_MIPS/Register/n796 ) );
  CLKMX2X2 U12214 ( .A(n5455), .B(\i_MIPS/Register/register[10][6] ), .S0(
        n5994), .Y(\i_MIPS/Register/n794 ) );
  CLKMX2X2 U12215 ( .A(n5226), .B(\i_MIPS/Register/register[10][4] ), .S0(
        n5994), .Y(\i_MIPS/Register/n792 ) );
  CLKMX2X2 U12216 ( .A(n5195), .B(\i_MIPS/Register/register[10][3] ), .S0(
        n5994), .Y(\i_MIPS/Register/n791 ) );
  CLKMX2X2 U12217 ( .A(n5463), .B(\i_MIPS/Register/register[10][2] ), .S0(
        n5994), .Y(\i_MIPS/Register/n790 ) );
  CLKMX2X2 U12218 ( .A(n5513), .B(\i_MIPS/Register/register[10][1] ), .S0(
        n5995), .Y(\i_MIPS/Register/n789 ) );
  CLKMX2X2 U12219 ( .A(n5501), .B(\i_MIPS/Register/register[11][29] ), .S0(
        n5993), .Y(\i_MIPS/Register/n785 ) );
  CLKMX2X2 U12220 ( .A(n5498), .B(\i_MIPS/Register/register[11][28] ), .S0(
        n5993), .Y(\i_MIPS/Register/n784 ) );
  CLKMX2X2 U12221 ( .A(n5472), .B(\i_MIPS/Register/register[11][27] ), .S0(
        n5992), .Y(\i_MIPS/Register/n783 ) );
  CLKMX2X2 U12222 ( .A(n5481), .B(\i_MIPS/Register/register[11][26] ), .S0(
        n5993), .Y(\i_MIPS/Register/n782 ) );
  CLKMX2X2 U12223 ( .A(n5470), .B(\i_MIPS/Register/register[11][22] ), .S0(
        n5992), .Y(\i_MIPS/Register/n778 ) );
  CLKMX2X2 U12224 ( .A(n5493), .B(\i_MIPS/Register/register[11][21] ), .S0(
        n5993), .Y(\i_MIPS/Register/n777 ) );
  CLKMX2X2 U12225 ( .A(n5474), .B(\i_MIPS/Register/register[11][20] ), .S0(
        n5992), .Y(\i_MIPS/Register/n776 ) );
  CLKMX2X2 U12226 ( .A(n5467), .B(\i_MIPS/Register/register[11][19] ), .S0(
        n5992), .Y(\i_MIPS/Register/n775 ) );
  CLKMX2X2 U12227 ( .A(n5509), .B(\i_MIPS/Register/register[11][18] ), .S0(
        n5993), .Y(\i_MIPS/Register/n774 ) );
  CLKMX2X2 U12228 ( .A(n5506), .B(\i_MIPS/Register/register[11][17] ), .S0(
        n5993), .Y(\i_MIPS/Register/n773 ) );
  CLKMX2X2 U12229 ( .A(n5490), .B(\i_MIPS/Register/register[11][16] ), .S0(
        n5993), .Y(\i_MIPS/Register/n772 ) );
  CLKMX2X2 U12230 ( .A(n5483), .B(\i_MIPS/Register/register[11][15] ), .S0(
        n5993), .Y(\i_MIPS/Register/n771 ) );
  CLKMX2X2 U12231 ( .A(n5488), .B(\i_MIPS/Register/register[11][14] ), .S0(
        n5992), .Y(\i_MIPS/Register/n770 ) );
  CLKMX2X2 U12232 ( .A(n5485), .B(\i_MIPS/Register/register[11][12] ), .S0(
        n5993), .Y(\i_MIPS/Register/n768 ) );
  CLKMX2X2 U12233 ( .A(n5495), .B(\i_MIPS/Register/register[11][10] ), .S0(
        n5993), .Y(\i_MIPS/Register/n766 ) );
  CLKMX2X2 U12234 ( .A(n5503), .B(\i_MIPS/Register/register[11][9] ), .S0(
        n5993), .Y(\i_MIPS/Register/n765 ) );
  CLKMX2X2 U12235 ( .A(n5512), .B(\i_MIPS/Register/register[11][8] ), .S0(
        n5993), .Y(\i_MIPS/Register/n764 ) );
  CLKMX2X2 U12236 ( .A(n5456), .B(\i_MIPS/Register/register[11][6] ), .S0(
        n5992), .Y(\i_MIPS/Register/n762 ) );
  CLKMX2X2 U12237 ( .A(n5227), .B(\i_MIPS/Register/register[11][4] ), .S0(
        n5992), .Y(\i_MIPS/Register/n760 ) );
  CLKMX2X2 U12238 ( .A(n5196), .B(\i_MIPS/Register/register[11][3] ), .S0(
        n5992), .Y(\i_MIPS/Register/n759 ) );
  CLKMX2X2 U12239 ( .A(n5464), .B(\i_MIPS/Register/register[11][2] ), .S0(
        n5992), .Y(\i_MIPS/Register/n758 ) );
  CLKMX2X2 U12240 ( .A(n5514), .B(\i_MIPS/Register/register[11][1] ), .S0(
        n5993), .Y(\i_MIPS/Register/n757 ) );
  CLKMX2X2 U12241 ( .A(n5500), .B(\i_MIPS/Register/register[12][29] ), .S0(
        n5991), .Y(\i_MIPS/Register/n753 ) );
  CLKMX2X2 U12242 ( .A(n5497), .B(\i_MIPS/Register/register[12][28] ), .S0(
        n5991), .Y(\i_MIPS/Register/n752 ) );
  CLKMX2X2 U12243 ( .A(n5471), .B(\i_MIPS/Register/register[12][27] ), .S0(
        n5990), .Y(\i_MIPS/Register/n751 ) );
  CLKMX2X2 U12244 ( .A(n5480), .B(\i_MIPS/Register/register[12][26] ), .S0(
        n5991), .Y(\i_MIPS/Register/n750 ) );
  CLKMX2X2 U12245 ( .A(n5469), .B(\i_MIPS/Register/register[12][22] ), .S0(
        n5990), .Y(\i_MIPS/Register/n746 ) );
  CLKMX2X2 U12246 ( .A(n5492), .B(\i_MIPS/Register/register[12][21] ), .S0(
        n5991), .Y(\i_MIPS/Register/n745 ) );
  CLKMX2X2 U12247 ( .A(n5473), .B(\i_MIPS/Register/register[12][20] ), .S0(
        n5990), .Y(\i_MIPS/Register/n744 ) );
  CLKMX2X2 U12248 ( .A(n5466), .B(\i_MIPS/Register/register[12][19] ), .S0(
        n5990), .Y(\i_MIPS/Register/n743 ) );
  CLKMX2X2 U12249 ( .A(n5508), .B(\i_MIPS/Register/register[12][18] ), .S0(
        n5991), .Y(\i_MIPS/Register/n742 ) );
  CLKMX2X2 U12250 ( .A(n5505), .B(\i_MIPS/Register/register[12][17] ), .S0(
        n5991), .Y(\i_MIPS/Register/n741 ) );
  CLKMX2X2 U12251 ( .A(n5489), .B(\i_MIPS/Register/register[12][16] ), .S0(
        n5991), .Y(\i_MIPS/Register/n740 ) );
  CLKMX2X2 U12252 ( .A(n5482), .B(\i_MIPS/Register/register[12][15] ), .S0(
        n5991), .Y(\i_MIPS/Register/n739 ) );
  CLKMX2X2 U12253 ( .A(n5487), .B(\i_MIPS/Register/register[12][14] ), .S0(
        n5990), .Y(\i_MIPS/Register/n738 ) );
  CLKMX2X2 U12254 ( .A(n5484), .B(\i_MIPS/Register/register[12][12] ), .S0(
        n5991), .Y(\i_MIPS/Register/n736 ) );
  CLKMX2X2 U12255 ( .A(n5494), .B(\i_MIPS/Register/register[12][10] ), .S0(
        n5991), .Y(\i_MIPS/Register/n734 ) );
  CLKMX2X2 U12256 ( .A(n5502), .B(\i_MIPS/Register/register[12][9] ), .S0(
        n5991), .Y(\i_MIPS/Register/n733 ) );
  CLKMX2X2 U12257 ( .A(n5511), .B(\i_MIPS/Register/register[12][8] ), .S0(
        n5991), .Y(\i_MIPS/Register/n732 ) );
  CLKMX2X2 U12258 ( .A(n5455), .B(\i_MIPS/Register/register[12][6] ), .S0(
        n5990), .Y(\i_MIPS/Register/n730 ) );
  CLKMX2X2 U12259 ( .A(n5226), .B(\i_MIPS/Register/register[12][4] ), .S0(
        n5990), .Y(\i_MIPS/Register/n728 ) );
  CLKMX2X2 U12260 ( .A(n5195), .B(\i_MIPS/Register/register[12][3] ), .S0(
        n5990), .Y(\i_MIPS/Register/n727 ) );
  CLKMX2X2 U12261 ( .A(n5463), .B(\i_MIPS/Register/register[12][2] ), .S0(
        n5990), .Y(\i_MIPS/Register/n726 ) );
  CLKMX2X2 U12262 ( .A(n5513), .B(\i_MIPS/Register/register[12][1] ), .S0(
        n5991), .Y(\i_MIPS/Register/n725 ) );
  CLKMX2X2 U12263 ( .A(n5500), .B(\i_MIPS/Register/register[13][29] ), .S0(
        n5989), .Y(\i_MIPS/Register/n721 ) );
  CLKMX2X2 U12264 ( .A(n5497), .B(\i_MIPS/Register/register[13][28] ), .S0(
        n5989), .Y(\i_MIPS/Register/n720 ) );
  CLKMX2X2 U12265 ( .A(n5471), .B(\i_MIPS/Register/register[13][27] ), .S0(
        n5988), .Y(\i_MIPS/Register/n719 ) );
  CLKMX2X2 U12266 ( .A(n5480), .B(\i_MIPS/Register/register[13][26] ), .S0(
        n5989), .Y(\i_MIPS/Register/n718 ) );
  CLKMX2X2 U12267 ( .A(n5469), .B(\i_MIPS/Register/register[13][22] ), .S0(
        n5988), .Y(\i_MIPS/Register/n714 ) );
  CLKMX2X2 U12268 ( .A(n5492), .B(\i_MIPS/Register/register[13][21] ), .S0(
        n5989), .Y(\i_MIPS/Register/n713 ) );
  CLKMX2X2 U12269 ( .A(n5473), .B(\i_MIPS/Register/register[13][20] ), .S0(
        n5988), .Y(\i_MIPS/Register/n712 ) );
  CLKMX2X2 U12270 ( .A(n5466), .B(\i_MIPS/Register/register[13][19] ), .S0(
        n5988), .Y(\i_MIPS/Register/n711 ) );
  CLKMX2X2 U12271 ( .A(n5508), .B(\i_MIPS/Register/register[13][18] ), .S0(
        n5989), .Y(\i_MIPS/Register/n710 ) );
  CLKMX2X2 U12272 ( .A(n5505), .B(\i_MIPS/Register/register[13][17] ), .S0(
        n5989), .Y(\i_MIPS/Register/n709 ) );
  CLKMX2X2 U12273 ( .A(n5489), .B(\i_MIPS/Register/register[13][16] ), .S0(
        n5989), .Y(\i_MIPS/Register/n708 ) );
  CLKMX2X2 U12274 ( .A(n5482), .B(\i_MIPS/Register/register[13][15] ), .S0(
        n5989), .Y(\i_MIPS/Register/n707 ) );
  CLKMX2X2 U12275 ( .A(n5487), .B(\i_MIPS/Register/register[13][14] ), .S0(
        n5988), .Y(\i_MIPS/Register/n706 ) );
  CLKMX2X2 U12276 ( .A(n5484), .B(\i_MIPS/Register/register[13][12] ), .S0(
        n5989), .Y(\i_MIPS/Register/n704 ) );
  CLKMX2X2 U12277 ( .A(n5494), .B(\i_MIPS/Register/register[13][10] ), .S0(
        n5989), .Y(\i_MIPS/Register/n702 ) );
  CLKMX2X2 U12278 ( .A(n5502), .B(\i_MIPS/Register/register[13][9] ), .S0(
        n5989), .Y(\i_MIPS/Register/n701 ) );
  CLKMX2X2 U12279 ( .A(n5511), .B(\i_MIPS/Register/register[13][8] ), .S0(
        n5989), .Y(\i_MIPS/Register/n700 ) );
  CLKMX2X2 U12280 ( .A(n5455), .B(\i_MIPS/Register/register[13][6] ), .S0(
        n5988), .Y(\i_MIPS/Register/n698 ) );
  CLKMX2X2 U12281 ( .A(n5226), .B(\i_MIPS/Register/register[13][4] ), .S0(
        n5988), .Y(\i_MIPS/Register/n696 ) );
  CLKMX2X2 U12282 ( .A(n5195), .B(\i_MIPS/Register/register[13][3] ), .S0(
        n5988), .Y(\i_MIPS/Register/n695 ) );
  CLKMX2X2 U12283 ( .A(n5463), .B(\i_MIPS/Register/register[13][2] ), .S0(
        n5988), .Y(\i_MIPS/Register/n694 ) );
  CLKMX2X2 U12284 ( .A(n5513), .B(\i_MIPS/Register/register[13][1] ), .S0(
        n5989), .Y(\i_MIPS/Register/n693 ) );
  CLKMX2X2 U12285 ( .A(n5500), .B(\i_MIPS/Register/register[14][29] ), .S0(
        n5987), .Y(\i_MIPS/Register/n689 ) );
  CLKMX2X2 U12286 ( .A(n5497), .B(\i_MIPS/Register/register[14][28] ), .S0(
        n5987), .Y(\i_MIPS/Register/n688 ) );
  CLKMX2X2 U12287 ( .A(n5471), .B(\i_MIPS/Register/register[14][27] ), .S0(
        n5986), .Y(\i_MIPS/Register/n687 ) );
  CLKMX2X2 U12288 ( .A(n5480), .B(\i_MIPS/Register/register[14][26] ), .S0(
        n5987), .Y(\i_MIPS/Register/n686 ) );
  CLKMX2X2 U12289 ( .A(n5469), .B(\i_MIPS/Register/register[14][22] ), .S0(
        n5986), .Y(\i_MIPS/Register/n682 ) );
  CLKMX2X2 U12290 ( .A(n5492), .B(\i_MIPS/Register/register[14][21] ), .S0(
        n5987), .Y(\i_MIPS/Register/n681 ) );
  CLKMX2X2 U12291 ( .A(n5473), .B(\i_MIPS/Register/register[14][20] ), .S0(
        n5986), .Y(\i_MIPS/Register/n680 ) );
  CLKMX2X2 U12292 ( .A(n5466), .B(\i_MIPS/Register/register[14][19] ), .S0(
        n5986), .Y(\i_MIPS/Register/n679 ) );
  CLKMX2X2 U12293 ( .A(n5508), .B(\i_MIPS/Register/register[14][18] ), .S0(
        n5987), .Y(\i_MIPS/Register/n678 ) );
  CLKMX2X2 U12294 ( .A(n5505), .B(\i_MIPS/Register/register[14][17] ), .S0(
        n5987), .Y(\i_MIPS/Register/n677 ) );
  CLKMX2X2 U12295 ( .A(n5489), .B(\i_MIPS/Register/register[14][16] ), .S0(
        n5987), .Y(\i_MIPS/Register/n676 ) );
  CLKMX2X2 U12296 ( .A(n5482), .B(\i_MIPS/Register/register[14][15] ), .S0(
        n5987), .Y(\i_MIPS/Register/n675 ) );
  CLKMX2X2 U12297 ( .A(n5487), .B(\i_MIPS/Register/register[14][14] ), .S0(
        n5986), .Y(\i_MIPS/Register/n674 ) );
  CLKMX2X2 U12298 ( .A(n5484), .B(\i_MIPS/Register/register[14][12] ), .S0(
        n5987), .Y(\i_MIPS/Register/n672 ) );
  CLKMX2X2 U12299 ( .A(n5494), .B(\i_MIPS/Register/register[14][10] ), .S0(
        n5987), .Y(\i_MIPS/Register/n670 ) );
  CLKMX2X2 U12300 ( .A(n5502), .B(\i_MIPS/Register/register[14][9] ), .S0(
        n5987), .Y(\i_MIPS/Register/n669 ) );
  CLKMX2X2 U12301 ( .A(n5511), .B(\i_MIPS/Register/register[14][8] ), .S0(
        n5987), .Y(\i_MIPS/Register/n668 ) );
  CLKMX2X2 U12302 ( .A(n5455), .B(\i_MIPS/Register/register[14][6] ), .S0(
        n5986), .Y(\i_MIPS/Register/n666 ) );
  CLKMX2X2 U12303 ( .A(n5226), .B(\i_MIPS/Register/register[14][4] ), .S0(
        n5986), .Y(\i_MIPS/Register/n664 ) );
  CLKMX2X2 U12304 ( .A(n5195), .B(\i_MIPS/Register/register[14][3] ), .S0(
        n5986), .Y(\i_MIPS/Register/n663 ) );
  CLKMX2X2 U12305 ( .A(n5463), .B(\i_MIPS/Register/register[14][2] ), .S0(
        n5986), .Y(\i_MIPS/Register/n662 ) );
  CLKMX2X2 U12306 ( .A(n5513), .B(\i_MIPS/Register/register[14][1] ), .S0(
        n5987), .Y(\i_MIPS/Register/n661 ) );
  CLKMX2X2 U12307 ( .A(n5501), .B(\i_MIPS/Register/register[15][29] ), .S0(
        n5985), .Y(\i_MIPS/Register/n657 ) );
  CLKMX2X2 U12308 ( .A(n5498), .B(\i_MIPS/Register/register[15][28] ), .S0(
        n5985), .Y(\i_MIPS/Register/n656 ) );
  CLKMX2X2 U12309 ( .A(n5472), .B(\i_MIPS/Register/register[15][27] ), .S0(
        n5984), .Y(\i_MIPS/Register/n655 ) );
  CLKMX2X2 U12310 ( .A(n5481), .B(\i_MIPS/Register/register[15][26] ), .S0(
        n5985), .Y(\i_MIPS/Register/n654 ) );
  CLKMX2X2 U12311 ( .A(n5470), .B(\i_MIPS/Register/register[15][22] ), .S0(
        n5984), .Y(\i_MIPS/Register/n650 ) );
  CLKMX2X2 U12312 ( .A(n5493), .B(\i_MIPS/Register/register[15][21] ), .S0(
        n5985), .Y(\i_MIPS/Register/n649 ) );
  CLKMX2X2 U12313 ( .A(n5474), .B(\i_MIPS/Register/register[15][20] ), .S0(
        n5984), .Y(\i_MIPS/Register/n648 ) );
  CLKMX2X2 U12314 ( .A(n5467), .B(\i_MIPS/Register/register[15][19] ), .S0(
        n5984), .Y(\i_MIPS/Register/n647 ) );
  CLKMX2X2 U12315 ( .A(n5509), .B(\i_MIPS/Register/register[15][18] ), .S0(
        n5985), .Y(\i_MIPS/Register/n646 ) );
  CLKMX2X2 U12316 ( .A(n5506), .B(\i_MIPS/Register/register[15][17] ), .S0(
        n5985), .Y(\i_MIPS/Register/n645 ) );
  CLKMX2X2 U12317 ( .A(n5490), .B(\i_MIPS/Register/register[15][16] ), .S0(
        n5985), .Y(\i_MIPS/Register/n644 ) );
  CLKMX2X2 U12318 ( .A(n5483), .B(\i_MIPS/Register/register[15][15] ), .S0(
        n5985), .Y(\i_MIPS/Register/n643 ) );
  CLKMX2X2 U12319 ( .A(n5488), .B(\i_MIPS/Register/register[15][14] ), .S0(
        n5984), .Y(\i_MIPS/Register/n642 ) );
  CLKMX2X2 U12320 ( .A(n5485), .B(\i_MIPS/Register/register[15][12] ), .S0(
        n5985), .Y(\i_MIPS/Register/n640 ) );
  CLKMX2X2 U12321 ( .A(n5495), .B(\i_MIPS/Register/register[15][10] ), .S0(
        n5985), .Y(\i_MIPS/Register/n638 ) );
  CLKMX2X2 U12322 ( .A(n5503), .B(\i_MIPS/Register/register[15][9] ), .S0(
        n5985), .Y(\i_MIPS/Register/n637 ) );
  CLKMX2X2 U12323 ( .A(n5512), .B(\i_MIPS/Register/register[15][8] ), .S0(
        n5985), .Y(\i_MIPS/Register/n636 ) );
  CLKMX2X2 U12324 ( .A(n5456), .B(\i_MIPS/Register/register[15][6] ), .S0(
        n5984), .Y(\i_MIPS/Register/n634 ) );
  CLKMX2X2 U12325 ( .A(n5227), .B(\i_MIPS/Register/register[15][4] ), .S0(
        n5984), .Y(\i_MIPS/Register/n632 ) );
  CLKMX2X2 U12326 ( .A(n5196), .B(\i_MIPS/Register/register[15][3] ), .S0(
        n5984), .Y(\i_MIPS/Register/n631 ) );
  CLKMX2X2 U12327 ( .A(n5464), .B(\i_MIPS/Register/register[15][2] ), .S0(
        n5984), .Y(\i_MIPS/Register/n630 ) );
  CLKMX2X2 U12328 ( .A(n5514), .B(\i_MIPS/Register/register[15][1] ), .S0(
        n5985), .Y(\i_MIPS/Register/n629 ) );
  CLKMX2X2 U12329 ( .A(n5501), .B(\i_MIPS/Register/register[16][29] ), .S0(
        n5983), .Y(\i_MIPS/Register/n625 ) );
  CLKMX2X2 U12330 ( .A(n5498), .B(\i_MIPS/Register/register[16][28] ), .S0(
        n5983), .Y(\i_MIPS/Register/n624 ) );
  CLKMX2X2 U12331 ( .A(n5472), .B(\i_MIPS/Register/register[16][27] ), .S0(
        n5982), .Y(\i_MIPS/Register/n623 ) );
  CLKMX2X2 U12332 ( .A(n5481), .B(\i_MIPS/Register/register[16][26] ), .S0(
        n5983), .Y(\i_MIPS/Register/n622 ) );
  CLKMX2X2 U12333 ( .A(n5470), .B(\i_MIPS/Register/register[16][22] ), .S0(
        n5982), .Y(\i_MIPS/Register/n618 ) );
  CLKMX2X2 U12334 ( .A(n5493), .B(\i_MIPS/Register/register[16][21] ), .S0(
        n5983), .Y(\i_MIPS/Register/n617 ) );
  CLKMX2X2 U12335 ( .A(n5474), .B(\i_MIPS/Register/register[16][20] ), .S0(
        n5982), .Y(\i_MIPS/Register/n616 ) );
  CLKMX2X2 U12336 ( .A(n5467), .B(\i_MIPS/Register/register[16][19] ), .S0(
        n5982), .Y(\i_MIPS/Register/n615 ) );
  CLKMX2X2 U12337 ( .A(n5509), .B(\i_MIPS/Register/register[16][18] ), .S0(
        n5983), .Y(\i_MIPS/Register/n614 ) );
  CLKMX2X2 U12338 ( .A(n5506), .B(\i_MIPS/Register/register[16][17] ), .S0(
        n5983), .Y(\i_MIPS/Register/n613 ) );
  CLKMX2X2 U12339 ( .A(n5490), .B(\i_MIPS/Register/register[16][16] ), .S0(
        n5983), .Y(\i_MIPS/Register/n612 ) );
  CLKMX2X2 U12340 ( .A(n5483), .B(\i_MIPS/Register/register[16][15] ), .S0(
        n5983), .Y(\i_MIPS/Register/n611 ) );
  CLKMX2X2 U12341 ( .A(n5488), .B(\i_MIPS/Register/register[16][14] ), .S0(
        n5982), .Y(\i_MIPS/Register/n610 ) );
  CLKMX2X2 U12342 ( .A(n5485), .B(\i_MIPS/Register/register[16][12] ), .S0(
        n5983), .Y(\i_MIPS/Register/n608 ) );
  CLKMX2X2 U12343 ( .A(n5495), .B(\i_MIPS/Register/register[16][10] ), .S0(
        n5983), .Y(\i_MIPS/Register/n606 ) );
  CLKMX2X2 U12344 ( .A(n5503), .B(\i_MIPS/Register/register[16][9] ), .S0(
        n5983), .Y(\i_MIPS/Register/n605 ) );
  CLKMX2X2 U12345 ( .A(n5512), .B(\i_MIPS/Register/register[16][8] ), .S0(
        n5983), .Y(\i_MIPS/Register/n604 ) );
  CLKMX2X2 U12346 ( .A(n5456), .B(\i_MIPS/Register/register[16][6] ), .S0(
        n5982), .Y(\i_MIPS/Register/n602 ) );
  CLKMX2X2 U12347 ( .A(n5227), .B(\i_MIPS/Register/register[16][4] ), .S0(
        n5982), .Y(\i_MIPS/Register/n600 ) );
  CLKMX2X2 U12348 ( .A(n5196), .B(\i_MIPS/Register/register[16][3] ), .S0(
        n5982), .Y(\i_MIPS/Register/n599 ) );
  CLKMX2X2 U12349 ( .A(n5464), .B(\i_MIPS/Register/register[16][2] ), .S0(
        n5982), .Y(\i_MIPS/Register/n598 ) );
  CLKMX2X2 U12350 ( .A(n5514), .B(\i_MIPS/Register/register[16][1] ), .S0(
        n5983), .Y(\i_MIPS/Register/n597 ) );
  CLKMX2X2 U12351 ( .A(n5501), .B(\i_MIPS/Register/register[17][29] ), .S0(
        n5981), .Y(\i_MIPS/Register/n593 ) );
  CLKMX2X2 U12352 ( .A(n5498), .B(\i_MIPS/Register/register[17][28] ), .S0(
        n5981), .Y(\i_MIPS/Register/n592 ) );
  CLKMX2X2 U12353 ( .A(n5472), .B(\i_MIPS/Register/register[17][27] ), .S0(
        n5980), .Y(\i_MIPS/Register/n591 ) );
  CLKMX2X2 U12354 ( .A(n5481), .B(\i_MIPS/Register/register[17][26] ), .S0(
        n5981), .Y(\i_MIPS/Register/n590 ) );
  CLKMX2X2 U12355 ( .A(n5470), .B(\i_MIPS/Register/register[17][22] ), .S0(
        n5980), .Y(\i_MIPS/Register/n586 ) );
  CLKMX2X2 U12356 ( .A(n5493), .B(\i_MIPS/Register/register[17][21] ), .S0(
        n5981), .Y(\i_MIPS/Register/n585 ) );
  CLKMX2X2 U12357 ( .A(n5474), .B(\i_MIPS/Register/register[17][20] ), .S0(
        n5980), .Y(\i_MIPS/Register/n584 ) );
  CLKMX2X2 U12358 ( .A(n5467), .B(\i_MIPS/Register/register[17][19] ), .S0(
        n5980), .Y(\i_MIPS/Register/n583 ) );
  CLKMX2X2 U12359 ( .A(n5509), .B(\i_MIPS/Register/register[17][18] ), .S0(
        n5981), .Y(\i_MIPS/Register/n582 ) );
  CLKMX2X2 U12360 ( .A(n5506), .B(\i_MIPS/Register/register[17][17] ), .S0(
        n5981), .Y(\i_MIPS/Register/n581 ) );
  CLKMX2X2 U12361 ( .A(n5490), .B(\i_MIPS/Register/register[17][16] ), .S0(
        n5981), .Y(\i_MIPS/Register/n580 ) );
  CLKMX2X2 U12362 ( .A(n5483), .B(\i_MIPS/Register/register[17][15] ), .S0(
        n5981), .Y(\i_MIPS/Register/n579 ) );
  CLKMX2X2 U12363 ( .A(n5488), .B(\i_MIPS/Register/register[17][14] ), .S0(
        n5980), .Y(\i_MIPS/Register/n578 ) );
  CLKMX2X2 U12364 ( .A(n5485), .B(\i_MIPS/Register/register[17][12] ), .S0(
        n5981), .Y(\i_MIPS/Register/n576 ) );
  CLKMX2X2 U12365 ( .A(n5495), .B(\i_MIPS/Register/register[17][10] ), .S0(
        n5981), .Y(\i_MIPS/Register/n574 ) );
  CLKMX2X2 U12366 ( .A(n5503), .B(\i_MIPS/Register/register[17][9] ), .S0(
        n5981), .Y(\i_MIPS/Register/n573 ) );
  CLKMX2X2 U12367 ( .A(n5512), .B(\i_MIPS/Register/register[17][8] ), .S0(
        n5981), .Y(\i_MIPS/Register/n572 ) );
  CLKMX2X2 U12368 ( .A(n5456), .B(\i_MIPS/Register/register[17][6] ), .S0(
        n5980), .Y(\i_MIPS/Register/n570 ) );
  CLKMX2X2 U12369 ( .A(n5227), .B(\i_MIPS/Register/register[17][4] ), .S0(
        n5980), .Y(\i_MIPS/Register/n568 ) );
  CLKMX2X2 U12370 ( .A(n5196), .B(\i_MIPS/Register/register[17][3] ), .S0(
        n5980), .Y(\i_MIPS/Register/n567 ) );
  CLKMX2X2 U12371 ( .A(n5464), .B(\i_MIPS/Register/register[17][2] ), .S0(
        n5980), .Y(\i_MIPS/Register/n566 ) );
  CLKMX2X2 U12372 ( .A(n5514), .B(\i_MIPS/Register/register[17][1] ), .S0(
        n5981), .Y(\i_MIPS/Register/n565 ) );
  CLKMX2X2 U12373 ( .A(n5501), .B(\i_MIPS/Register/register[18][29] ), .S0(
        n5979), .Y(\i_MIPS/Register/n561 ) );
  CLKMX2X2 U12374 ( .A(n5498), .B(\i_MIPS/Register/register[18][28] ), .S0(
        n5979), .Y(\i_MIPS/Register/n560 ) );
  CLKMX2X2 U12375 ( .A(n5472), .B(\i_MIPS/Register/register[18][27] ), .S0(
        n5978), .Y(\i_MIPS/Register/n559 ) );
  CLKMX2X2 U12376 ( .A(n5481), .B(\i_MIPS/Register/register[18][26] ), .S0(
        n5979), .Y(\i_MIPS/Register/n558 ) );
  CLKMX2X2 U12377 ( .A(n5470), .B(\i_MIPS/Register/register[18][22] ), .S0(
        n5978), .Y(\i_MIPS/Register/n554 ) );
  CLKMX2X2 U12378 ( .A(n5493), .B(\i_MIPS/Register/register[18][21] ), .S0(
        n5979), .Y(\i_MIPS/Register/n553 ) );
  CLKMX2X2 U12379 ( .A(n5474), .B(\i_MIPS/Register/register[18][20] ), .S0(
        n5978), .Y(\i_MIPS/Register/n552 ) );
  CLKMX2X2 U12380 ( .A(n5467), .B(\i_MIPS/Register/register[18][19] ), .S0(
        n5978), .Y(\i_MIPS/Register/n551 ) );
  CLKMX2X2 U12381 ( .A(n5509), .B(\i_MIPS/Register/register[18][18] ), .S0(
        n5979), .Y(\i_MIPS/Register/n550 ) );
  CLKMX2X2 U12382 ( .A(n5506), .B(\i_MIPS/Register/register[18][17] ), .S0(
        n5979), .Y(\i_MIPS/Register/n549 ) );
  CLKMX2X2 U12383 ( .A(n5490), .B(\i_MIPS/Register/register[18][16] ), .S0(
        n5979), .Y(\i_MIPS/Register/n548 ) );
  CLKMX2X2 U12384 ( .A(n5483), .B(\i_MIPS/Register/register[18][15] ), .S0(
        n5979), .Y(\i_MIPS/Register/n547 ) );
  CLKMX2X2 U12385 ( .A(n5488), .B(\i_MIPS/Register/register[18][14] ), .S0(
        n5978), .Y(\i_MIPS/Register/n546 ) );
  CLKMX2X2 U12386 ( .A(n5485), .B(\i_MIPS/Register/register[18][12] ), .S0(
        n5979), .Y(\i_MIPS/Register/n544 ) );
  CLKMX2X2 U12387 ( .A(n5495), .B(\i_MIPS/Register/register[18][10] ), .S0(
        n5979), .Y(\i_MIPS/Register/n542 ) );
  CLKMX2X2 U12388 ( .A(n5503), .B(\i_MIPS/Register/register[18][9] ), .S0(
        n5979), .Y(\i_MIPS/Register/n541 ) );
  CLKMX2X2 U12389 ( .A(n5512), .B(\i_MIPS/Register/register[18][8] ), .S0(
        n5979), .Y(\i_MIPS/Register/n540 ) );
  CLKMX2X2 U12390 ( .A(n5456), .B(\i_MIPS/Register/register[18][6] ), .S0(
        n5978), .Y(\i_MIPS/Register/n538 ) );
  CLKMX2X2 U12391 ( .A(n5227), .B(\i_MIPS/Register/register[18][4] ), .S0(
        n5978), .Y(\i_MIPS/Register/n536 ) );
  CLKMX2X2 U12392 ( .A(n5196), .B(\i_MIPS/Register/register[18][3] ), .S0(
        n5978), .Y(\i_MIPS/Register/n535 ) );
  CLKMX2X2 U12393 ( .A(n5464), .B(\i_MIPS/Register/register[18][2] ), .S0(
        n5978), .Y(\i_MIPS/Register/n534 ) );
  CLKMX2X2 U12394 ( .A(n5514), .B(\i_MIPS/Register/register[18][1] ), .S0(
        n5979), .Y(\i_MIPS/Register/n533 ) );
  CLKMX2X2 U12395 ( .A(n5501), .B(\i_MIPS/Register/register[19][29] ), .S0(
        n5977), .Y(\i_MIPS/Register/n529 ) );
  CLKMX2X2 U12396 ( .A(n10539), .B(\i_MIPS/Register/register[19][28] ), .S0(
        n5977), .Y(\i_MIPS/Register/n528 ) );
  CLKMX2X2 U12397 ( .A(n5471), .B(\i_MIPS/Register/register[19][27] ), .S0(
        n5976), .Y(\i_MIPS/Register/n527 ) );
  CLKMX2X2 U12398 ( .A(n5481), .B(\i_MIPS/Register/register[19][26] ), .S0(
        n5977), .Y(\i_MIPS/Register/n526 ) );
  CLKMX2X2 U12399 ( .A(n5478), .B(\i_MIPS/Register/register[19][25] ), .S0(
        n5976), .Y(\i_MIPS/Register/n525 ) );
  CLKMX2X2 U12400 ( .A(n5476), .B(\i_MIPS/Register/register[19][24] ), .S0(
        n5976), .Y(\i_MIPS/Register/n524 ) );
  CLKMX2X2 U12401 ( .A(n5469), .B(\i_MIPS/Register/register[19][22] ), .S0(
        n5976), .Y(\i_MIPS/Register/n522 ) );
  CLKMX2X2 U12402 ( .A(n5493), .B(\i_MIPS/Register/register[19][21] ), .S0(
        n5977), .Y(\i_MIPS/Register/n521 ) );
  CLKMX2X2 U12403 ( .A(n5474), .B(\i_MIPS/Register/register[19][20] ), .S0(
        n5976), .Y(\i_MIPS/Register/n520 ) );
  CLKMX2X2 U12404 ( .A(n5467), .B(\i_MIPS/Register/register[19][19] ), .S0(
        n5976), .Y(\i_MIPS/Register/n519 ) );
  CLKMX2X2 U12405 ( .A(n5509), .B(\i_MIPS/Register/register[19][18] ), .S0(
        n5977), .Y(\i_MIPS/Register/n518 ) );
  CLKMX2X2 U12406 ( .A(n5506), .B(\i_MIPS/Register/register[19][17] ), .S0(
        n5977), .Y(\i_MIPS/Register/n517 ) );
  CLKMX2X2 U12407 ( .A(n5490), .B(\i_MIPS/Register/register[19][16] ), .S0(
        n5977), .Y(\i_MIPS/Register/n516 ) );
  CLKMX2X2 U12408 ( .A(n5483), .B(\i_MIPS/Register/register[19][15] ), .S0(
        n5977), .Y(\i_MIPS/Register/n515 ) );
  CLKMX2X2 U12409 ( .A(n5487), .B(\i_MIPS/Register/register[19][14] ), .S0(
        n5976), .Y(\i_MIPS/Register/n514 ) );
  CLKMX2X2 U12410 ( .A(n5485), .B(\i_MIPS/Register/register[19][12] ), .S0(
        n5977), .Y(\i_MIPS/Register/n512 ) );
  CLKMX2X2 U12411 ( .A(n5495), .B(\i_MIPS/Register/register[19][10] ), .S0(
        n5977), .Y(\i_MIPS/Register/n510 ) );
  CLKMX2X2 U12412 ( .A(n5503), .B(\i_MIPS/Register/register[19][9] ), .S0(
        n5977), .Y(\i_MIPS/Register/n509 ) );
  CLKMX2X2 U12413 ( .A(n5512), .B(\i_MIPS/Register/register[19][8] ), .S0(
        n5977), .Y(\i_MIPS/Register/n508 ) );
  CLKMX2X2 U12414 ( .A(n5456), .B(\i_MIPS/Register/register[19][6] ), .S0(
        n5976), .Y(\i_MIPS/Register/n506 ) );
  CLKMX2X2 U12415 ( .A(n5227), .B(\i_MIPS/Register/register[19][4] ), .S0(
        n5976), .Y(\i_MIPS/Register/n504 ) );
  CLKMX2X2 U12416 ( .A(n5195), .B(\i_MIPS/Register/register[19][3] ), .S0(
        n5976), .Y(\i_MIPS/Register/n503 ) );
  CLKMX2X2 U12417 ( .A(n5463), .B(\i_MIPS/Register/register[19][2] ), .S0(
        n5976), .Y(\i_MIPS/Register/n502 ) );
  CLKMX2X2 U12418 ( .A(n5513), .B(\i_MIPS/Register/register[19][1] ), .S0(
        n5977), .Y(\i_MIPS/Register/n501 ) );
  CLKMX2X2 U12419 ( .A(n5501), .B(\i_MIPS/Register/register[20][29] ), .S0(
        n5975), .Y(\i_MIPS/Register/n497 ) );
  CLKMX2X2 U12420 ( .A(n5498), .B(\i_MIPS/Register/register[20][28] ), .S0(
        n5975), .Y(\i_MIPS/Register/n496 ) );
  CLKMX2X2 U12421 ( .A(n5472), .B(\i_MIPS/Register/register[20][27] ), .S0(
        n5974), .Y(\i_MIPS/Register/n495 ) );
  CLKMX2X2 U12422 ( .A(n5481), .B(\i_MIPS/Register/register[20][26] ), .S0(
        n5975), .Y(\i_MIPS/Register/n494 ) );
  CLKMX2X2 U12423 ( .A(n5470), .B(\i_MIPS/Register/register[20][22] ), .S0(
        n5974), .Y(\i_MIPS/Register/n490 ) );
  CLKMX2X2 U12424 ( .A(n5493), .B(\i_MIPS/Register/register[20][21] ), .S0(
        n5975), .Y(\i_MIPS/Register/n489 ) );
  CLKMX2X2 U12425 ( .A(n5474), .B(\i_MIPS/Register/register[20][20] ), .S0(
        n5974), .Y(\i_MIPS/Register/n488 ) );
  CLKMX2X2 U12426 ( .A(n5467), .B(\i_MIPS/Register/register[20][19] ), .S0(
        n5974), .Y(\i_MIPS/Register/n487 ) );
  CLKMX2X2 U12427 ( .A(n5509), .B(\i_MIPS/Register/register[20][18] ), .S0(
        n5975), .Y(\i_MIPS/Register/n486 ) );
  CLKMX2X2 U12428 ( .A(n5506), .B(\i_MIPS/Register/register[20][17] ), .S0(
        n5975), .Y(\i_MIPS/Register/n485 ) );
  CLKMX2X2 U12429 ( .A(n5490), .B(\i_MIPS/Register/register[20][16] ), .S0(
        n5975), .Y(\i_MIPS/Register/n484 ) );
  CLKMX2X2 U12430 ( .A(n5483), .B(\i_MIPS/Register/register[20][15] ), .S0(
        n5975), .Y(\i_MIPS/Register/n483 ) );
  CLKMX2X2 U12431 ( .A(n5488), .B(\i_MIPS/Register/register[20][14] ), .S0(
        n5974), .Y(\i_MIPS/Register/n482 ) );
  CLKMX2X2 U12432 ( .A(n5485), .B(\i_MIPS/Register/register[20][12] ), .S0(
        n5975), .Y(\i_MIPS/Register/n480 ) );
  CLKMX2X2 U12433 ( .A(n5495), .B(\i_MIPS/Register/register[20][10] ), .S0(
        n5975), .Y(\i_MIPS/Register/n478 ) );
  CLKMX2X2 U12434 ( .A(n5503), .B(\i_MIPS/Register/register[20][9] ), .S0(
        n5975), .Y(\i_MIPS/Register/n477 ) );
  CLKMX2X2 U12435 ( .A(n5512), .B(\i_MIPS/Register/register[20][8] ), .S0(
        n5975), .Y(\i_MIPS/Register/n476 ) );
  CLKMX2X2 U12436 ( .A(n5456), .B(\i_MIPS/Register/register[20][6] ), .S0(
        n5974), .Y(\i_MIPS/Register/n474 ) );
  CLKMX2X2 U12437 ( .A(n5227), .B(\i_MIPS/Register/register[20][4] ), .S0(
        n5974), .Y(\i_MIPS/Register/n472 ) );
  CLKMX2X2 U12438 ( .A(n5196), .B(\i_MIPS/Register/register[20][3] ), .S0(
        n5974), .Y(\i_MIPS/Register/n471 ) );
  CLKMX2X2 U12439 ( .A(n5464), .B(\i_MIPS/Register/register[20][2] ), .S0(
        n5974), .Y(\i_MIPS/Register/n470 ) );
  CLKMX2X2 U12440 ( .A(n5514), .B(\i_MIPS/Register/register[20][1] ), .S0(
        n5975), .Y(\i_MIPS/Register/n469 ) );
  CLKMX2X2 U12441 ( .A(n5500), .B(\i_MIPS/Register/register[21][29] ), .S0(
        n5973), .Y(\i_MIPS/Register/n465 ) );
  CLKMX2X2 U12442 ( .A(n10539), .B(\i_MIPS/Register/register[21][28] ), .S0(
        n5973), .Y(\i_MIPS/Register/n464 ) );
  CLKMX2X2 U12443 ( .A(n5472), .B(\i_MIPS/Register/register[21][27] ), .S0(
        n5972), .Y(\i_MIPS/Register/n463 ) );
  CLKMX2X2 U12444 ( .A(n5480), .B(\i_MIPS/Register/register[21][26] ), .S0(
        n5973), .Y(\i_MIPS/Register/n462 ) );
  CLKMX2X2 U12445 ( .A(n5479), .B(\i_MIPS/Register/register[21][25] ), .S0(
        n5972), .Y(\i_MIPS/Register/n461 ) );
  CLKMX2X2 U12446 ( .A(n5477), .B(\i_MIPS/Register/register[21][24] ), .S0(
        n5972), .Y(\i_MIPS/Register/n460 ) );
  CLKMX2X2 U12447 ( .A(n5470), .B(\i_MIPS/Register/register[21][22] ), .S0(
        n5972), .Y(\i_MIPS/Register/n458 ) );
  CLKMX2X2 U12448 ( .A(n5492), .B(\i_MIPS/Register/register[21][21] ), .S0(
        n5973), .Y(\i_MIPS/Register/n457 ) );
  CLKMX2X2 U12449 ( .A(n5473), .B(\i_MIPS/Register/register[21][20] ), .S0(
        n5972), .Y(\i_MIPS/Register/n456 ) );
  CLKMX2X2 U12450 ( .A(n5466), .B(\i_MIPS/Register/register[21][19] ), .S0(
        n5972), .Y(\i_MIPS/Register/n455 ) );
  CLKMX2X2 U12451 ( .A(n5508), .B(\i_MIPS/Register/register[21][18] ), .S0(
        n5973), .Y(\i_MIPS/Register/n454 ) );
  CLKMX2X2 U12452 ( .A(n5505), .B(\i_MIPS/Register/register[21][17] ), .S0(
        n5973), .Y(\i_MIPS/Register/n453 ) );
  CLKMX2X2 U12453 ( .A(n5489), .B(\i_MIPS/Register/register[21][16] ), .S0(
        n5973), .Y(\i_MIPS/Register/n452 ) );
  CLKMX2X2 U12454 ( .A(n5482), .B(\i_MIPS/Register/register[21][15] ), .S0(
        n5973), .Y(\i_MIPS/Register/n451 ) );
  CLKMX2X2 U12455 ( .A(n5488), .B(\i_MIPS/Register/register[21][14] ), .S0(
        n5972), .Y(\i_MIPS/Register/n450 ) );
  CLKMX2X2 U12456 ( .A(n5484), .B(\i_MIPS/Register/register[21][12] ), .S0(
        n5973), .Y(\i_MIPS/Register/n448 ) );
  CLKMX2X2 U12457 ( .A(n5494), .B(\i_MIPS/Register/register[21][10] ), .S0(
        n5973), .Y(\i_MIPS/Register/n446 ) );
  CLKMX2X2 U12458 ( .A(n5502), .B(\i_MIPS/Register/register[21][9] ), .S0(
        n5973), .Y(\i_MIPS/Register/n445 ) );
  CLKMX2X2 U12459 ( .A(n5511), .B(\i_MIPS/Register/register[21][8] ), .S0(
        n5973), .Y(\i_MIPS/Register/n444 ) );
  CLKMX2X2 U12460 ( .A(n5455), .B(\i_MIPS/Register/register[21][6] ), .S0(
        n5972), .Y(\i_MIPS/Register/n442 ) );
  CLKMX2X2 U12461 ( .A(n5226), .B(\i_MIPS/Register/register[21][4] ), .S0(
        n5972), .Y(\i_MIPS/Register/n440 ) );
  CLKMX2X2 U12462 ( .A(n5196), .B(\i_MIPS/Register/register[21][3] ), .S0(
        n5972), .Y(\i_MIPS/Register/n439 ) );
  CLKMX2X2 U12463 ( .A(n5464), .B(\i_MIPS/Register/register[21][2] ), .S0(
        n5972), .Y(\i_MIPS/Register/n438 ) );
  CLKMX2X2 U12464 ( .A(n5514), .B(\i_MIPS/Register/register[21][1] ), .S0(
        n5973), .Y(\i_MIPS/Register/n437 ) );
  CLKMX2X2 U12465 ( .A(n5501), .B(\i_MIPS/Register/register[22][29] ), .S0(
        n5971), .Y(\i_MIPS/Register/n433 ) );
  CLKMX2X2 U12466 ( .A(n5498), .B(\i_MIPS/Register/register[22][28] ), .S0(
        n5971), .Y(\i_MIPS/Register/n432 ) );
  CLKMX2X2 U12467 ( .A(n5472), .B(\i_MIPS/Register/register[22][27] ), .S0(
        n5970), .Y(\i_MIPS/Register/n431 ) );
  CLKMX2X2 U12468 ( .A(n5481), .B(\i_MIPS/Register/register[22][26] ), .S0(
        n5971), .Y(\i_MIPS/Register/n430 ) );
  CLKMX2X2 U12469 ( .A(n5470), .B(\i_MIPS/Register/register[22][22] ), .S0(
        n5970), .Y(\i_MIPS/Register/n426 ) );
  CLKMX2X2 U12470 ( .A(n5493), .B(\i_MIPS/Register/register[22][21] ), .S0(
        n5971), .Y(\i_MIPS/Register/n425 ) );
  CLKMX2X2 U12471 ( .A(n5474), .B(\i_MIPS/Register/register[22][20] ), .S0(
        n5970), .Y(\i_MIPS/Register/n424 ) );
  CLKMX2X2 U12472 ( .A(n5467), .B(\i_MIPS/Register/register[22][19] ), .S0(
        n5970), .Y(\i_MIPS/Register/n423 ) );
  CLKMX2X2 U12473 ( .A(n5509), .B(\i_MIPS/Register/register[22][18] ), .S0(
        n5971), .Y(\i_MIPS/Register/n422 ) );
  CLKMX2X2 U12474 ( .A(n5506), .B(\i_MIPS/Register/register[22][17] ), .S0(
        n5971), .Y(\i_MIPS/Register/n421 ) );
  CLKMX2X2 U12475 ( .A(n5490), .B(\i_MIPS/Register/register[22][16] ), .S0(
        n5971), .Y(\i_MIPS/Register/n420 ) );
  CLKMX2X2 U12476 ( .A(n5483), .B(\i_MIPS/Register/register[22][15] ), .S0(
        n5971), .Y(\i_MIPS/Register/n419 ) );
  CLKMX2X2 U12477 ( .A(n5488), .B(\i_MIPS/Register/register[22][14] ), .S0(
        n5970), .Y(\i_MIPS/Register/n418 ) );
  CLKMX2X2 U12478 ( .A(n5485), .B(\i_MIPS/Register/register[22][12] ), .S0(
        n5971), .Y(\i_MIPS/Register/n416 ) );
  CLKMX2X2 U12479 ( .A(n5495), .B(\i_MIPS/Register/register[22][10] ), .S0(
        n5971), .Y(\i_MIPS/Register/n414 ) );
  CLKMX2X2 U12480 ( .A(n5503), .B(\i_MIPS/Register/register[22][9] ), .S0(
        n5971), .Y(\i_MIPS/Register/n413 ) );
  CLKMX2X2 U12481 ( .A(n5512), .B(\i_MIPS/Register/register[22][8] ), .S0(
        n5971), .Y(\i_MIPS/Register/n412 ) );
  CLKMX2X2 U12482 ( .A(n5456), .B(\i_MIPS/Register/register[22][6] ), .S0(
        n5970), .Y(\i_MIPS/Register/n410 ) );
  CLKMX2X2 U12483 ( .A(n5227), .B(\i_MIPS/Register/register[22][4] ), .S0(
        n5970), .Y(\i_MIPS/Register/n408 ) );
  CLKMX2X2 U12484 ( .A(n5196), .B(\i_MIPS/Register/register[22][3] ), .S0(
        n5970), .Y(\i_MIPS/Register/n407 ) );
  CLKMX2X2 U12485 ( .A(n5464), .B(\i_MIPS/Register/register[22][2] ), .S0(
        n5970), .Y(\i_MIPS/Register/n406 ) );
  CLKMX2X2 U12486 ( .A(n5514), .B(\i_MIPS/Register/register[22][1] ), .S0(
        n5971), .Y(\i_MIPS/Register/n405 ) );
  CLKMX2X2 U12487 ( .A(n5501), .B(\i_MIPS/Register/register[23][29] ), .S0(
        n5969), .Y(\i_MIPS/Register/n401 ) );
  CLKMX2X2 U12488 ( .A(n10539), .B(\i_MIPS/Register/register[23][28] ), .S0(
        n5969), .Y(\i_MIPS/Register/n400 ) );
  CLKMX2X2 U12489 ( .A(n5471), .B(\i_MIPS/Register/register[23][27] ), .S0(
        n5968), .Y(\i_MIPS/Register/n399 ) );
  CLKMX2X2 U12490 ( .A(n5481), .B(\i_MIPS/Register/register[23][26] ), .S0(
        n5969), .Y(\i_MIPS/Register/n398 ) );
  CLKMX2X2 U12491 ( .A(n5478), .B(\i_MIPS/Register/register[23][25] ), .S0(
        n5968), .Y(\i_MIPS/Register/n397 ) );
  CLKMX2X2 U12492 ( .A(n5476), .B(\i_MIPS/Register/register[23][24] ), .S0(
        n5968), .Y(\i_MIPS/Register/n396 ) );
  CLKMX2X2 U12493 ( .A(n5469), .B(\i_MIPS/Register/register[23][22] ), .S0(
        n5968), .Y(\i_MIPS/Register/n394 ) );
  CLKMX2X2 U12494 ( .A(n5493), .B(\i_MIPS/Register/register[23][21] ), .S0(
        n5969), .Y(\i_MIPS/Register/n393 ) );
  CLKMX2X2 U12495 ( .A(n5474), .B(\i_MIPS/Register/register[23][20] ), .S0(
        n5968), .Y(\i_MIPS/Register/n392 ) );
  CLKMX2X2 U12496 ( .A(n5467), .B(\i_MIPS/Register/register[23][19] ), .S0(
        n5968), .Y(\i_MIPS/Register/n391 ) );
  CLKMX2X2 U12497 ( .A(n5509), .B(\i_MIPS/Register/register[23][18] ), .S0(
        n5969), .Y(\i_MIPS/Register/n390 ) );
  CLKMX2X2 U12498 ( .A(n5506), .B(\i_MIPS/Register/register[23][17] ), .S0(
        n5969), .Y(\i_MIPS/Register/n389 ) );
  CLKMX2X2 U12499 ( .A(n5490), .B(\i_MIPS/Register/register[23][16] ), .S0(
        n5969), .Y(\i_MIPS/Register/n388 ) );
  CLKMX2X2 U12500 ( .A(n5483), .B(\i_MIPS/Register/register[23][15] ), .S0(
        n5969), .Y(\i_MIPS/Register/n387 ) );
  CLKMX2X2 U12501 ( .A(n5487), .B(\i_MIPS/Register/register[23][14] ), .S0(
        n5968), .Y(\i_MIPS/Register/n386 ) );
  CLKMX2X2 U12502 ( .A(n5485), .B(\i_MIPS/Register/register[23][12] ), .S0(
        n5969), .Y(\i_MIPS/Register/n384 ) );
  CLKMX2X2 U12503 ( .A(n5495), .B(\i_MIPS/Register/register[23][10] ), .S0(
        n5969), .Y(\i_MIPS/Register/n382 ) );
  CLKMX2X2 U12504 ( .A(n5503), .B(\i_MIPS/Register/register[23][9] ), .S0(
        n5969), .Y(\i_MIPS/Register/n381 ) );
  CLKMX2X2 U12505 ( .A(n5512), .B(\i_MIPS/Register/register[23][8] ), .S0(
        n5969), .Y(\i_MIPS/Register/n380 ) );
  CLKMX2X2 U12506 ( .A(n5456), .B(\i_MIPS/Register/register[23][6] ), .S0(
        n5968), .Y(\i_MIPS/Register/n378 ) );
  CLKMX2X2 U12507 ( .A(n5227), .B(\i_MIPS/Register/register[23][4] ), .S0(
        n5968), .Y(\i_MIPS/Register/n376 ) );
  CLKMX2X2 U12508 ( .A(n5195), .B(\i_MIPS/Register/register[23][3] ), .S0(
        n5968), .Y(\i_MIPS/Register/n375 ) );
  CLKMX2X2 U12509 ( .A(n5463), .B(\i_MIPS/Register/register[23][2] ), .S0(
        n5968), .Y(\i_MIPS/Register/n374 ) );
  CLKMX2X2 U12510 ( .A(n5513), .B(\i_MIPS/Register/register[23][1] ), .S0(
        n5969), .Y(\i_MIPS/Register/n373 ) );
  CLKMX2X2 U12511 ( .A(n5501), .B(\i_MIPS/Register/register[24][29] ), .S0(
        n5967), .Y(\i_MIPS/Register/n369 ) );
  CLKMX2X2 U12512 ( .A(n5498), .B(\i_MIPS/Register/register[24][28] ), .S0(
        n5967), .Y(\i_MIPS/Register/n368 ) );
  CLKMX2X2 U12513 ( .A(n5472), .B(\i_MIPS/Register/register[24][27] ), .S0(
        n5966), .Y(\i_MIPS/Register/n367 ) );
  CLKMX2X2 U12514 ( .A(n5481), .B(\i_MIPS/Register/register[24][26] ), .S0(
        n5967), .Y(\i_MIPS/Register/n366 ) );
  CLKMX2X2 U12515 ( .A(n5470), .B(\i_MIPS/Register/register[24][22] ), .S0(
        n5966), .Y(\i_MIPS/Register/n362 ) );
  CLKMX2X2 U12516 ( .A(n5493), .B(\i_MIPS/Register/register[24][21] ), .S0(
        n5967), .Y(\i_MIPS/Register/n361 ) );
  CLKMX2X2 U12517 ( .A(n5474), .B(\i_MIPS/Register/register[24][20] ), .S0(
        n5966), .Y(\i_MIPS/Register/n360 ) );
  CLKMX2X2 U12518 ( .A(n5467), .B(\i_MIPS/Register/register[24][19] ), .S0(
        n5966), .Y(\i_MIPS/Register/n359 ) );
  CLKMX2X2 U12519 ( .A(n5509), .B(\i_MIPS/Register/register[24][18] ), .S0(
        n5967), .Y(\i_MIPS/Register/n358 ) );
  CLKMX2X2 U12520 ( .A(n5506), .B(\i_MIPS/Register/register[24][17] ), .S0(
        n5967), .Y(\i_MIPS/Register/n357 ) );
  CLKMX2X2 U12521 ( .A(n5490), .B(\i_MIPS/Register/register[24][16] ), .S0(
        n5967), .Y(\i_MIPS/Register/n356 ) );
  CLKMX2X2 U12522 ( .A(n5483), .B(\i_MIPS/Register/register[24][15] ), .S0(
        n5967), .Y(\i_MIPS/Register/n355 ) );
  CLKMX2X2 U12523 ( .A(n5488), .B(\i_MIPS/Register/register[24][14] ), .S0(
        n5966), .Y(\i_MIPS/Register/n354 ) );
  CLKMX2X2 U12524 ( .A(n5485), .B(\i_MIPS/Register/register[24][12] ), .S0(
        n5967), .Y(\i_MIPS/Register/n352 ) );
  CLKMX2X2 U12525 ( .A(n5495), .B(\i_MIPS/Register/register[24][10] ), .S0(
        n5967), .Y(\i_MIPS/Register/n350 ) );
  CLKMX2X2 U12526 ( .A(n5503), .B(\i_MIPS/Register/register[24][9] ), .S0(
        n5967), .Y(\i_MIPS/Register/n349 ) );
  CLKMX2X2 U12527 ( .A(n5512), .B(\i_MIPS/Register/register[24][8] ), .S0(
        n5967), .Y(\i_MIPS/Register/n348 ) );
  CLKMX2X2 U12528 ( .A(n5456), .B(\i_MIPS/Register/register[24][6] ), .S0(
        n5966), .Y(\i_MIPS/Register/n346 ) );
  CLKMX2X2 U12529 ( .A(n5227), .B(\i_MIPS/Register/register[24][4] ), .S0(
        n5966), .Y(\i_MIPS/Register/n344 ) );
  CLKMX2X2 U12530 ( .A(n5196), .B(\i_MIPS/Register/register[24][3] ), .S0(
        n5966), .Y(\i_MIPS/Register/n343 ) );
  CLKMX2X2 U12531 ( .A(n5464), .B(\i_MIPS/Register/register[24][2] ), .S0(
        n5966), .Y(\i_MIPS/Register/n342 ) );
  CLKMX2X2 U12532 ( .A(n5514), .B(\i_MIPS/Register/register[24][1] ), .S0(
        n5967), .Y(\i_MIPS/Register/n341 ) );
  CLKMX2X2 U12533 ( .A(n5501), .B(\i_MIPS/Register/register[25][29] ), .S0(
        n5965), .Y(\i_MIPS/Register/n337 ) );
  CLKMX2X2 U12534 ( .A(n5498), .B(\i_MIPS/Register/register[25][28] ), .S0(
        n5965), .Y(\i_MIPS/Register/n336 ) );
  CLKMX2X2 U12535 ( .A(n5472), .B(\i_MIPS/Register/register[25][27] ), .S0(
        n5964), .Y(\i_MIPS/Register/n335 ) );
  CLKMX2X2 U12536 ( .A(n5481), .B(\i_MIPS/Register/register[25][26] ), .S0(
        n5965), .Y(\i_MIPS/Register/n334 ) );
  CLKMX2X2 U12537 ( .A(n5470), .B(\i_MIPS/Register/register[25][22] ), .S0(
        n5964), .Y(\i_MIPS/Register/n330 ) );
  CLKMX2X2 U12538 ( .A(n5493), .B(\i_MIPS/Register/register[25][21] ), .S0(
        n5965), .Y(\i_MIPS/Register/n329 ) );
  CLKMX2X2 U12539 ( .A(n5474), .B(\i_MIPS/Register/register[25][20] ), .S0(
        n5964), .Y(\i_MIPS/Register/n328 ) );
  CLKMX2X2 U12540 ( .A(n5467), .B(\i_MIPS/Register/register[25][19] ), .S0(
        n5964), .Y(\i_MIPS/Register/n327 ) );
  CLKMX2X2 U12541 ( .A(n5509), .B(\i_MIPS/Register/register[25][18] ), .S0(
        n5965), .Y(\i_MIPS/Register/n326 ) );
  CLKMX2X2 U12542 ( .A(n5506), .B(\i_MIPS/Register/register[25][17] ), .S0(
        n5965), .Y(\i_MIPS/Register/n325 ) );
  CLKMX2X2 U12543 ( .A(n5490), .B(\i_MIPS/Register/register[25][16] ), .S0(
        n5965), .Y(\i_MIPS/Register/n324 ) );
  CLKMX2X2 U12544 ( .A(n5483), .B(\i_MIPS/Register/register[25][15] ), .S0(
        n5965), .Y(\i_MIPS/Register/n323 ) );
  CLKMX2X2 U12545 ( .A(n5488), .B(\i_MIPS/Register/register[25][14] ), .S0(
        n5964), .Y(\i_MIPS/Register/n322 ) );
  CLKMX2X2 U12546 ( .A(n5485), .B(\i_MIPS/Register/register[25][12] ), .S0(
        n5965), .Y(\i_MIPS/Register/n320 ) );
  CLKMX2X2 U12547 ( .A(n5495), .B(\i_MIPS/Register/register[25][10] ), .S0(
        n5965), .Y(\i_MIPS/Register/n318 ) );
  CLKMX2X2 U12548 ( .A(n5503), .B(\i_MIPS/Register/register[25][9] ), .S0(
        n5965), .Y(\i_MIPS/Register/n317 ) );
  CLKMX2X2 U12549 ( .A(n5512), .B(\i_MIPS/Register/register[25][8] ), .S0(
        n5965), .Y(\i_MIPS/Register/n316 ) );
  CLKMX2X2 U12550 ( .A(n5456), .B(\i_MIPS/Register/register[25][6] ), .S0(
        n5964), .Y(\i_MIPS/Register/n314 ) );
  CLKMX2X2 U12551 ( .A(n5227), .B(\i_MIPS/Register/register[25][4] ), .S0(
        n5964), .Y(\i_MIPS/Register/n312 ) );
  CLKMX2X2 U12552 ( .A(n5196), .B(\i_MIPS/Register/register[25][3] ), .S0(
        n5964), .Y(\i_MIPS/Register/n311 ) );
  CLKMX2X2 U12553 ( .A(n5464), .B(\i_MIPS/Register/register[25][2] ), .S0(
        n5964), .Y(\i_MIPS/Register/n310 ) );
  CLKMX2X2 U12554 ( .A(n5514), .B(\i_MIPS/Register/register[25][1] ), .S0(
        n5965), .Y(\i_MIPS/Register/n309 ) );
  CLKMX2X2 U12555 ( .A(n5501), .B(\i_MIPS/Register/register[26][29] ), .S0(
        n5963), .Y(\i_MIPS/Register/n305 ) );
  CLKMX2X2 U12556 ( .A(n5498), .B(\i_MIPS/Register/register[26][28] ), .S0(
        n5963), .Y(\i_MIPS/Register/n304 ) );
  CLKMX2X2 U12557 ( .A(n5472), .B(\i_MIPS/Register/register[26][27] ), .S0(
        n5962), .Y(\i_MIPS/Register/n303 ) );
  CLKMX2X2 U12558 ( .A(n5481), .B(\i_MIPS/Register/register[26][26] ), .S0(
        n5963), .Y(\i_MIPS/Register/n302 ) );
  CLKMX2X2 U12559 ( .A(n5470), .B(\i_MIPS/Register/register[26][22] ), .S0(
        n5962), .Y(\i_MIPS/Register/n298 ) );
  CLKMX2X2 U12560 ( .A(n5493), .B(\i_MIPS/Register/register[26][21] ), .S0(
        n5963), .Y(\i_MIPS/Register/n297 ) );
  CLKMX2X2 U12561 ( .A(n5474), .B(\i_MIPS/Register/register[26][20] ), .S0(
        n5962), .Y(\i_MIPS/Register/n296 ) );
  CLKMX2X2 U12562 ( .A(n5467), .B(\i_MIPS/Register/register[26][19] ), .S0(
        n5962), .Y(\i_MIPS/Register/n295 ) );
  CLKMX2X2 U12563 ( .A(n5509), .B(\i_MIPS/Register/register[26][18] ), .S0(
        n5963), .Y(\i_MIPS/Register/n294 ) );
  CLKMX2X2 U12564 ( .A(n5506), .B(\i_MIPS/Register/register[26][17] ), .S0(
        n5963), .Y(\i_MIPS/Register/n293 ) );
  CLKMX2X2 U12565 ( .A(n5490), .B(\i_MIPS/Register/register[26][16] ), .S0(
        n5963), .Y(\i_MIPS/Register/n292 ) );
  CLKMX2X2 U12566 ( .A(n5483), .B(\i_MIPS/Register/register[26][15] ), .S0(
        n5963), .Y(\i_MIPS/Register/n291 ) );
  CLKMX2X2 U12567 ( .A(n5488), .B(\i_MIPS/Register/register[26][14] ), .S0(
        n5962), .Y(\i_MIPS/Register/n290 ) );
  CLKMX2X2 U12568 ( .A(n5485), .B(\i_MIPS/Register/register[26][12] ), .S0(
        n5963), .Y(\i_MIPS/Register/n288 ) );
  CLKMX2X2 U12569 ( .A(n5495), .B(\i_MIPS/Register/register[26][10] ), .S0(
        n5963), .Y(\i_MIPS/Register/n286 ) );
  CLKMX2X2 U12570 ( .A(n5503), .B(\i_MIPS/Register/register[26][9] ), .S0(
        n5963), .Y(\i_MIPS/Register/n285 ) );
  CLKMX2X2 U12571 ( .A(n5512), .B(\i_MIPS/Register/register[26][8] ), .S0(
        n5963), .Y(\i_MIPS/Register/n284 ) );
  CLKMX2X2 U12572 ( .A(n5456), .B(\i_MIPS/Register/register[26][6] ), .S0(
        n5962), .Y(\i_MIPS/Register/n282 ) );
  CLKMX2X2 U12573 ( .A(n5227), .B(\i_MIPS/Register/register[26][4] ), .S0(
        n5962), .Y(\i_MIPS/Register/n280 ) );
  CLKMX2X2 U12574 ( .A(n5196), .B(\i_MIPS/Register/register[26][3] ), .S0(
        n5962), .Y(\i_MIPS/Register/n279 ) );
  CLKMX2X2 U12575 ( .A(n5464), .B(\i_MIPS/Register/register[26][2] ), .S0(
        n5962), .Y(\i_MIPS/Register/n278 ) );
  CLKMX2X2 U12576 ( .A(n5514), .B(\i_MIPS/Register/register[26][1] ), .S0(
        n5963), .Y(\i_MIPS/Register/n277 ) );
  CLKMX2X2 U12577 ( .A(n5500), .B(\i_MIPS/Register/register[27][29] ), .S0(
        n5961), .Y(\i_MIPS/Register/n273 ) );
  CLKMX2X2 U12578 ( .A(n10539), .B(\i_MIPS/Register/register[27][28] ), .S0(
        n5961), .Y(\i_MIPS/Register/n272 ) );
  CLKMX2X2 U12579 ( .A(n5472), .B(\i_MIPS/Register/register[27][27] ), .S0(
        n5960), .Y(\i_MIPS/Register/n271 ) );
  CLKMX2X2 U12580 ( .A(n5480), .B(\i_MIPS/Register/register[27][26] ), .S0(
        n5961), .Y(\i_MIPS/Register/n270 ) );
  CLKMX2X2 U12581 ( .A(n5479), .B(\i_MIPS/Register/register[27][25] ), .S0(
        n5960), .Y(\i_MIPS/Register/n269 ) );
  CLKMX2X2 U12582 ( .A(n5477), .B(\i_MIPS/Register/register[27][24] ), .S0(
        n5960), .Y(\i_MIPS/Register/n268 ) );
  CLKMX2X2 U12583 ( .A(n5470), .B(\i_MIPS/Register/register[27][22] ), .S0(
        n5960), .Y(\i_MIPS/Register/n266 ) );
  CLKMX2X2 U12584 ( .A(n5492), .B(\i_MIPS/Register/register[27][21] ), .S0(
        n5961), .Y(\i_MIPS/Register/n265 ) );
  CLKMX2X2 U12585 ( .A(n5473), .B(\i_MIPS/Register/register[27][20] ), .S0(
        n5960), .Y(\i_MIPS/Register/n264 ) );
  CLKMX2X2 U12586 ( .A(n5466), .B(\i_MIPS/Register/register[27][19] ), .S0(
        n5960), .Y(\i_MIPS/Register/n263 ) );
  CLKMX2X2 U12587 ( .A(n5508), .B(\i_MIPS/Register/register[27][18] ), .S0(
        n5961), .Y(\i_MIPS/Register/n262 ) );
  CLKMX2X2 U12588 ( .A(n5505), .B(\i_MIPS/Register/register[27][17] ), .S0(
        n5961), .Y(\i_MIPS/Register/n261 ) );
  CLKMX2X2 U12589 ( .A(n5489), .B(\i_MIPS/Register/register[27][16] ), .S0(
        n5961), .Y(\i_MIPS/Register/n260 ) );
  CLKMX2X2 U12590 ( .A(n5482), .B(\i_MIPS/Register/register[27][15] ), .S0(
        n5961), .Y(\i_MIPS/Register/n259 ) );
  CLKMX2X2 U12591 ( .A(n5488), .B(\i_MIPS/Register/register[27][14] ), .S0(
        n5960), .Y(\i_MIPS/Register/n258 ) );
  CLKMX2X2 U12592 ( .A(n5484), .B(\i_MIPS/Register/register[27][12] ), .S0(
        n5961), .Y(\i_MIPS/Register/n256 ) );
  CLKMX2X2 U12593 ( .A(n5494), .B(\i_MIPS/Register/register[27][10] ), .S0(
        n5961), .Y(\i_MIPS/Register/n254 ) );
  CLKMX2X2 U12594 ( .A(n5502), .B(\i_MIPS/Register/register[27][9] ), .S0(
        n5961), .Y(\i_MIPS/Register/n253 ) );
  CLKMX2X2 U12595 ( .A(n5511), .B(\i_MIPS/Register/register[27][8] ), .S0(
        n5961), .Y(\i_MIPS/Register/n252 ) );
  CLKMX2X2 U12596 ( .A(n5455), .B(\i_MIPS/Register/register[27][6] ), .S0(
        n5960), .Y(\i_MIPS/Register/n250 ) );
  CLKMX2X2 U12597 ( .A(n5226), .B(\i_MIPS/Register/register[27][4] ), .S0(
        n5960), .Y(\i_MIPS/Register/n248 ) );
  CLKMX2X2 U12598 ( .A(n5196), .B(\i_MIPS/Register/register[27][3] ), .S0(
        n5960), .Y(\i_MIPS/Register/n247 ) );
  CLKMX2X2 U12599 ( .A(n5464), .B(\i_MIPS/Register/register[27][2] ), .S0(
        n5960), .Y(\i_MIPS/Register/n246 ) );
  CLKMX2X2 U12600 ( .A(n5514), .B(\i_MIPS/Register/register[27][1] ), .S0(
        n5961), .Y(\i_MIPS/Register/n245 ) );
  CLKMX2X2 U12601 ( .A(n5501), .B(\i_MIPS/Register/register[28][29] ), .S0(
        n5959), .Y(\i_MIPS/Register/n241 ) );
  CLKMX2X2 U12602 ( .A(n5498), .B(\i_MIPS/Register/register[28][28] ), .S0(
        n5959), .Y(\i_MIPS/Register/n240 ) );
  CLKMX2X2 U12603 ( .A(n5472), .B(\i_MIPS/Register/register[28][27] ), .S0(
        n5958), .Y(\i_MIPS/Register/n239 ) );
  CLKMX2X2 U12604 ( .A(n5481), .B(\i_MIPS/Register/register[28][26] ), .S0(
        n5959), .Y(\i_MIPS/Register/n238 ) );
  CLKMX2X2 U12605 ( .A(n5470), .B(\i_MIPS/Register/register[28][22] ), .S0(
        n5958), .Y(\i_MIPS/Register/n234 ) );
  CLKMX2X2 U12606 ( .A(n5493), .B(\i_MIPS/Register/register[28][21] ), .S0(
        n5959), .Y(\i_MIPS/Register/n233 ) );
  CLKMX2X2 U12607 ( .A(n5474), .B(\i_MIPS/Register/register[28][20] ), .S0(
        n5958), .Y(\i_MIPS/Register/n232 ) );
  CLKMX2X2 U12608 ( .A(n5467), .B(\i_MIPS/Register/register[28][19] ), .S0(
        n5958), .Y(\i_MIPS/Register/n231 ) );
  CLKMX2X2 U12609 ( .A(n5509), .B(\i_MIPS/Register/register[28][18] ), .S0(
        n5959), .Y(\i_MIPS/Register/n230 ) );
  CLKMX2X2 U12610 ( .A(n5506), .B(\i_MIPS/Register/register[28][17] ), .S0(
        n5959), .Y(\i_MIPS/Register/n229 ) );
  CLKMX2X2 U12611 ( .A(n5490), .B(\i_MIPS/Register/register[28][16] ), .S0(
        n5959), .Y(\i_MIPS/Register/n228 ) );
  CLKMX2X2 U12612 ( .A(n5483), .B(\i_MIPS/Register/register[28][15] ), .S0(
        n5959), .Y(\i_MIPS/Register/n227 ) );
  CLKMX2X2 U12613 ( .A(n5488), .B(\i_MIPS/Register/register[28][14] ), .S0(
        n5958), .Y(\i_MIPS/Register/n226 ) );
  CLKMX2X2 U12614 ( .A(n5485), .B(\i_MIPS/Register/register[28][12] ), .S0(
        n5959), .Y(\i_MIPS/Register/n224 ) );
  CLKMX2X2 U12615 ( .A(n5495), .B(\i_MIPS/Register/register[28][10] ), .S0(
        n5959), .Y(\i_MIPS/Register/n222 ) );
  CLKMX2X2 U12616 ( .A(n5503), .B(\i_MIPS/Register/register[28][9] ), .S0(
        n5959), .Y(\i_MIPS/Register/n221 ) );
  CLKMX2X2 U12617 ( .A(n5512), .B(\i_MIPS/Register/register[28][8] ), .S0(
        n5959), .Y(\i_MIPS/Register/n220 ) );
  CLKMX2X2 U12618 ( .A(n5456), .B(\i_MIPS/Register/register[28][6] ), .S0(
        n5958), .Y(\i_MIPS/Register/n218 ) );
  CLKMX2X2 U12619 ( .A(n5227), .B(\i_MIPS/Register/register[28][4] ), .S0(
        n5958), .Y(\i_MIPS/Register/n216 ) );
  CLKMX2X2 U12620 ( .A(n5196), .B(\i_MIPS/Register/register[28][3] ), .S0(
        n5958), .Y(\i_MIPS/Register/n215 ) );
  CLKMX2X2 U12621 ( .A(n5464), .B(\i_MIPS/Register/register[28][2] ), .S0(
        n5958), .Y(\i_MIPS/Register/n214 ) );
  CLKMX2X2 U12622 ( .A(n5514), .B(\i_MIPS/Register/register[28][1] ), .S0(
        n5959), .Y(\i_MIPS/Register/n213 ) );
  CLKMX2X2 U12623 ( .A(n5501), .B(\i_MIPS/Register/register[29][29] ), .S0(
        n5957), .Y(\i_MIPS/Register/n209 ) );
  CLKMX2X2 U12624 ( .A(n10539), .B(\i_MIPS/Register/register[29][28] ), .S0(
        n5957), .Y(\i_MIPS/Register/n208 ) );
  CLKMX2X2 U12625 ( .A(n5471), .B(\i_MIPS/Register/register[29][27] ), .S0(
        n5956), .Y(\i_MIPS/Register/n207 ) );
  CLKMX2X2 U12626 ( .A(n5481), .B(\i_MIPS/Register/register[29][26] ), .S0(
        n5957), .Y(\i_MIPS/Register/n206 ) );
  CLKMX2X2 U12627 ( .A(n5478), .B(\i_MIPS/Register/register[29][25] ), .S0(
        n5956), .Y(\i_MIPS/Register/n205 ) );
  CLKMX2X2 U12628 ( .A(n5476), .B(\i_MIPS/Register/register[29][24] ), .S0(
        n5956), .Y(\i_MIPS/Register/n204 ) );
  CLKMX2X2 U12629 ( .A(n5469), .B(\i_MIPS/Register/register[29][22] ), .S0(
        n5956), .Y(\i_MIPS/Register/n202 ) );
  CLKMX2X2 U12630 ( .A(n5493), .B(\i_MIPS/Register/register[29][21] ), .S0(
        n5957), .Y(\i_MIPS/Register/n201 ) );
  CLKMX2X2 U12631 ( .A(n5474), .B(\i_MIPS/Register/register[29][20] ), .S0(
        n5956), .Y(\i_MIPS/Register/n200 ) );
  CLKMX2X2 U12632 ( .A(n5467), .B(\i_MIPS/Register/register[29][19] ), .S0(
        n5956), .Y(\i_MIPS/Register/n199 ) );
  CLKMX2X2 U12633 ( .A(n5509), .B(\i_MIPS/Register/register[29][18] ), .S0(
        n5957), .Y(\i_MIPS/Register/n198 ) );
  CLKMX2X2 U12634 ( .A(n5506), .B(\i_MIPS/Register/register[29][17] ), .S0(
        n5957), .Y(\i_MIPS/Register/n197 ) );
  CLKMX2X2 U12635 ( .A(n5490), .B(\i_MIPS/Register/register[29][16] ), .S0(
        n5957), .Y(\i_MIPS/Register/n196 ) );
  CLKMX2X2 U12636 ( .A(n5483), .B(\i_MIPS/Register/register[29][15] ), .S0(
        n5957), .Y(\i_MIPS/Register/n195 ) );
  CLKMX2X2 U12637 ( .A(n5487), .B(\i_MIPS/Register/register[29][14] ), .S0(
        n5956), .Y(\i_MIPS/Register/n194 ) );
  CLKMX2X2 U12638 ( .A(n5485), .B(\i_MIPS/Register/register[29][12] ), .S0(
        n5957), .Y(\i_MIPS/Register/n192 ) );
  CLKMX2X2 U12639 ( .A(n5495), .B(\i_MIPS/Register/register[29][10] ), .S0(
        n5957), .Y(\i_MIPS/Register/n190 ) );
  CLKMX2X2 U12640 ( .A(n5503), .B(\i_MIPS/Register/register[29][9] ), .S0(
        n5957), .Y(\i_MIPS/Register/n189 ) );
  CLKMX2X2 U12641 ( .A(n5512), .B(\i_MIPS/Register/register[29][8] ), .S0(
        n5957), .Y(\i_MIPS/Register/n188 ) );
  CLKMX2X2 U12642 ( .A(n9938), .B(\i_MIPS/Register/register[29][6] ), .S0(
        n5956), .Y(\i_MIPS/Register/n186 ) );
  CLKMX2X2 U12643 ( .A(n5227), .B(\i_MIPS/Register/register[29][4] ), .S0(
        n5956), .Y(\i_MIPS/Register/n184 ) );
  CLKMX2X2 U12644 ( .A(n5195), .B(\i_MIPS/Register/register[29][3] ), .S0(
        n5956), .Y(\i_MIPS/Register/n183 ) );
  CLKMX2X2 U12645 ( .A(n5463), .B(\i_MIPS/Register/register[29][2] ), .S0(
        n5956), .Y(\i_MIPS/Register/n182 ) );
  CLKMX2X2 U12646 ( .A(n5513), .B(\i_MIPS/Register/register[29][1] ), .S0(
        n5957), .Y(\i_MIPS/Register/n181 ) );
  CLKMX2X2 U12647 ( .A(n5501), .B(\i_MIPS/Register/register[30][29] ), .S0(
        n5955), .Y(\i_MIPS/Register/n177 ) );
  CLKMX2X2 U12648 ( .A(n5498), .B(\i_MIPS/Register/register[30][28] ), .S0(
        n5955), .Y(\i_MIPS/Register/n176 ) );
  CLKMX2X2 U12649 ( .A(n5472), .B(\i_MIPS/Register/register[30][27] ), .S0(
        n5954), .Y(\i_MIPS/Register/n175 ) );
  CLKMX2X2 U12650 ( .A(n5481), .B(\i_MIPS/Register/register[30][26] ), .S0(
        n5955), .Y(\i_MIPS/Register/n174 ) );
  CLKMX2X2 U12651 ( .A(n5470), .B(\i_MIPS/Register/register[30][22] ), .S0(
        n5954), .Y(\i_MIPS/Register/n170 ) );
  CLKMX2X2 U12652 ( .A(n5493), .B(\i_MIPS/Register/register[30][21] ), .S0(
        n5955), .Y(\i_MIPS/Register/n169 ) );
  CLKMX2X2 U12653 ( .A(n5474), .B(\i_MIPS/Register/register[30][20] ), .S0(
        n5954), .Y(\i_MIPS/Register/n168 ) );
  CLKMX2X2 U12654 ( .A(n5467), .B(\i_MIPS/Register/register[30][19] ), .S0(
        n5954), .Y(\i_MIPS/Register/n167 ) );
  CLKMX2X2 U12655 ( .A(n5509), .B(\i_MIPS/Register/register[30][18] ), .S0(
        n5955), .Y(\i_MIPS/Register/n166 ) );
  CLKMX2X2 U12656 ( .A(n5506), .B(\i_MIPS/Register/register[30][17] ), .S0(
        n5955), .Y(\i_MIPS/Register/n165 ) );
  CLKMX2X2 U12657 ( .A(n5490), .B(\i_MIPS/Register/register[30][16] ), .S0(
        n5955), .Y(\i_MIPS/Register/n164 ) );
  CLKMX2X2 U12658 ( .A(n5483), .B(\i_MIPS/Register/register[30][15] ), .S0(
        n5955), .Y(\i_MIPS/Register/n163 ) );
  CLKMX2X2 U12659 ( .A(n5488), .B(\i_MIPS/Register/register[30][14] ), .S0(
        n5954), .Y(\i_MIPS/Register/n162 ) );
  CLKMX2X2 U12660 ( .A(n5485), .B(\i_MIPS/Register/register[30][12] ), .S0(
        n5955), .Y(\i_MIPS/Register/n160 ) );
  CLKMX2X2 U12661 ( .A(n5495), .B(\i_MIPS/Register/register[30][10] ), .S0(
        n5955), .Y(\i_MIPS/Register/n158 ) );
  CLKMX2X2 U12662 ( .A(n5503), .B(\i_MIPS/Register/register[30][9] ), .S0(
        n5955), .Y(\i_MIPS/Register/n157 ) );
  CLKMX2X2 U12663 ( .A(n5512), .B(\i_MIPS/Register/register[30][8] ), .S0(
        n5955), .Y(\i_MIPS/Register/n156 ) );
  CLKMX2X2 U12664 ( .A(n5456), .B(\i_MIPS/Register/register[30][6] ), .S0(
        n5954), .Y(\i_MIPS/Register/n154 ) );
  CLKMX2X2 U12665 ( .A(n5227), .B(\i_MIPS/Register/register[30][4] ), .S0(
        n5954), .Y(\i_MIPS/Register/n152 ) );
  CLKMX2X2 U12666 ( .A(n5196), .B(\i_MIPS/Register/register[30][3] ), .S0(
        n5954), .Y(\i_MIPS/Register/n151 ) );
  CLKMX2X2 U12667 ( .A(n5464), .B(\i_MIPS/Register/register[30][2] ), .S0(
        n5954), .Y(\i_MIPS/Register/n150 ) );
  CLKMX2X2 U12668 ( .A(n5514), .B(\i_MIPS/Register/register[30][1] ), .S0(
        n5955), .Y(\i_MIPS/Register/n149 ) );
  MX2XL U12669 ( .A(n5050), .B(n2948), .S0(n3591), .Y(\i_MIPS/n442 ) );
  MXI2X1 U12670 ( .A(n3674), .B(\i_MIPS/n512 ), .S0(n3591), .Y(\i_MIPS/n439 )
         );
  MX2XL U12671 ( .A(n5478), .B(\i_MIPS/Register/register[1][25] ), .S0(n6012), 
        .Y(\i_MIPS/Register/n1101 ) );
  MX2XL U12672 ( .A(n5476), .B(\i_MIPS/Register/register[1][24] ), .S0(n6012), 
        .Y(\i_MIPS/Register/n1100 ) );
  MX2XL U12673 ( .A(n5478), .B(\i_MIPS/Register/register[2][25] ), .S0(n6010), 
        .Y(\i_MIPS/Register/n1069 ) );
  MX2XL U12674 ( .A(n5476), .B(\i_MIPS/Register/register[2][24] ), .S0(n6010), 
        .Y(\i_MIPS/Register/n1068 ) );
  MX2XL U12675 ( .A(n5478), .B(\i_MIPS/Register/register[3][25] ), .S0(n6008), 
        .Y(\i_MIPS/Register/n1037 ) );
  MX2XL U12676 ( .A(n5476), .B(\i_MIPS/Register/register[3][24] ), .S0(n6008), 
        .Y(\i_MIPS/Register/n1036 ) );
  MX2XL U12677 ( .A(n5478), .B(\i_MIPS/Register/register[4][25] ), .S0(n6006), 
        .Y(\i_MIPS/Register/n1005 ) );
  MX2XL U12678 ( .A(n5476), .B(\i_MIPS/Register/register[4][24] ), .S0(n6006), 
        .Y(\i_MIPS/Register/n1004 ) );
  MX2XL U12679 ( .A(n5478), .B(\i_MIPS/Register/register[5][25] ), .S0(n6004), 
        .Y(\i_MIPS/Register/n973 ) );
  MX2XL U12680 ( .A(n5476), .B(\i_MIPS/Register/register[5][24] ), .S0(n6004), 
        .Y(\i_MIPS/Register/n972 ) );
  MX2XL U12681 ( .A(n5478), .B(\i_MIPS/Register/register[6][25] ), .S0(n6002), 
        .Y(\i_MIPS/Register/n941 ) );
  MX2XL U12682 ( .A(n5476), .B(\i_MIPS/Register/register[6][24] ), .S0(n6002), 
        .Y(\i_MIPS/Register/n940 ) );
  MX2XL U12683 ( .A(n5478), .B(\i_MIPS/Register/register[8][25] ), .S0(n5998), 
        .Y(\i_MIPS/Register/n877 ) );
  MX2XL U12684 ( .A(n5476), .B(\i_MIPS/Register/register[8][24] ), .S0(n5998), 
        .Y(\i_MIPS/Register/n876 ) );
  MX2XL U12685 ( .A(n5478), .B(\i_MIPS/Register/register[9][25] ), .S0(n5996), 
        .Y(\i_MIPS/Register/n845 ) );
  MX2XL U12686 ( .A(n5476), .B(\i_MIPS/Register/register[9][24] ), .S0(n5996), 
        .Y(\i_MIPS/Register/n844 ) );
  MX2XL U12687 ( .A(n5478), .B(\i_MIPS/Register/register[10][25] ), .S0(n5994), 
        .Y(\i_MIPS/Register/n813 ) );
  MX2XL U12688 ( .A(n5476), .B(\i_MIPS/Register/register[10][24] ), .S0(n5994), 
        .Y(\i_MIPS/Register/n812 ) );
  MX2XL U12689 ( .A(n5479), .B(\i_MIPS/Register/register[11][25] ), .S0(n5992), 
        .Y(\i_MIPS/Register/n781 ) );
  MX2XL U12690 ( .A(n5477), .B(\i_MIPS/Register/register[11][24] ), .S0(n5992), 
        .Y(\i_MIPS/Register/n780 ) );
  MX2XL U12691 ( .A(n5478), .B(\i_MIPS/Register/register[12][25] ), .S0(n5990), 
        .Y(\i_MIPS/Register/n749 ) );
  MX2XL U12692 ( .A(n5476), .B(\i_MIPS/Register/register[12][24] ), .S0(n5990), 
        .Y(\i_MIPS/Register/n748 ) );
  MX2XL U12693 ( .A(n5478), .B(\i_MIPS/Register/register[13][25] ), .S0(n5988), 
        .Y(\i_MIPS/Register/n717 ) );
  MX2XL U12694 ( .A(n5476), .B(\i_MIPS/Register/register[13][24] ), .S0(n5988), 
        .Y(\i_MIPS/Register/n716 ) );
  MX2XL U12695 ( .A(n5478), .B(\i_MIPS/Register/register[14][25] ), .S0(n5986), 
        .Y(\i_MIPS/Register/n685 ) );
  MX2XL U12696 ( .A(n5476), .B(\i_MIPS/Register/register[14][24] ), .S0(n5986), 
        .Y(\i_MIPS/Register/n684 ) );
  MX2XL U12697 ( .A(n5479), .B(\i_MIPS/Register/register[15][25] ), .S0(n5984), 
        .Y(\i_MIPS/Register/n653 ) );
  MX2XL U12698 ( .A(n5477), .B(\i_MIPS/Register/register[15][24] ), .S0(n5984), 
        .Y(\i_MIPS/Register/n652 ) );
  MX2XL U12699 ( .A(n5479), .B(\i_MIPS/Register/register[16][25] ), .S0(n5982), 
        .Y(\i_MIPS/Register/n621 ) );
  MX2XL U12700 ( .A(n5477), .B(\i_MIPS/Register/register[16][24] ), .S0(n5982), 
        .Y(\i_MIPS/Register/n620 ) );
  MX2XL U12701 ( .A(n5479), .B(\i_MIPS/Register/register[17][25] ), .S0(n5980), 
        .Y(\i_MIPS/Register/n589 ) );
  MX2XL U12702 ( .A(n5477), .B(\i_MIPS/Register/register[17][24] ), .S0(n5980), 
        .Y(\i_MIPS/Register/n588 ) );
  MX2XL U12703 ( .A(n5479), .B(\i_MIPS/Register/register[18][25] ), .S0(n5978), 
        .Y(\i_MIPS/Register/n557 ) );
  MX2XL U12704 ( .A(n5477), .B(\i_MIPS/Register/register[18][24] ), .S0(n5978), 
        .Y(\i_MIPS/Register/n556 ) );
  MX2XL U12705 ( .A(n5479), .B(\i_MIPS/Register/register[20][25] ), .S0(n5974), 
        .Y(\i_MIPS/Register/n493 ) );
  MX2XL U12706 ( .A(n5477), .B(\i_MIPS/Register/register[20][24] ), .S0(n5974), 
        .Y(\i_MIPS/Register/n492 ) );
  MX2XL U12707 ( .A(n5479), .B(\i_MIPS/Register/register[22][25] ), .S0(n5970), 
        .Y(\i_MIPS/Register/n429 ) );
  MX2XL U12708 ( .A(n5477), .B(\i_MIPS/Register/register[22][24] ), .S0(n5970), 
        .Y(\i_MIPS/Register/n428 ) );
  MX2XL U12709 ( .A(n5479), .B(\i_MIPS/Register/register[24][25] ), .S0(n5966), 
        .Y(\i_MIPS/Register/n365 ) );
  MX2XL U12710 ( .A(n5477), .B(\i_MIPS/Register/register[24][24] ), .S0(n5966), 
        .Y(\i_MIPS/Register/n364 ) );
  MX2XL U12711 ( .A(n5479), .B(\i_MIPS/Register/register[25][25] ), .S0(n5964), 
        .Y(\i_MIPS/Register/n333 ) );
  MX2XL U12712 ( .A(n5477), .B(\i_MIPS/Register/register[25][24] ), .S0(n5964), 
        .Y(\i_MIPS/Register/n332 ) );
  MX2XL U12713 ( .A(n5479), .B(\i_MIPS/Register/register[26][25] ), .S0(n5962), 
        .Y(\i_MIPS/Register/n301 ) );
  MX2XL U12714 ( .A(n5477), .B(\i_MIPS/Register/register[26][24] ), .S0(n5962), 
        .Y(\i_MIPS/Register/n300 ) );
  MX2XL U12715 ( .A(n5479), .B(\i_MIPS/Register/register[28][25] ), .S0(n5958), 
        .Y(\i_MIPS/Register/n237 ) );
  MX2XL U12716 ( .A(n5477), .B(\i_MIPS/Register/register[28][24] ), .S0(n5958), 
        .Y(\i_MIPS/Register/n236 ) );
  MX2XL U12717 ( .A(n5479), .B(\i_MIPS/Register/register[30][25] ), .S0(n5954), 
        .Y(\i_MIPS/Register/n173 ) );
  MX2XL U12718 ( .A(n5477), .B(\i_MIPS/Register/register[30][24] ), .S0(n5954), 
        .Y(\i_MIPS/Register/n172 ) );
  CLKMX2X2 U12719 ( .A(n5460), .B(\i_MIPS/Register/register[0][30] ), .S0(
        n6014), .Y(\i_MIPS/Register/n1138 ) );
  CLKMX2X2 U12720 ( .A(n5458), .B(\i_MIPS/Register/register[0][5] ), .S0(n6014), .Y(\i_MIPS/Register/n1113 ) );
  CLKMX2X2 U12721 ( .A(n5460), .B(\i_MIPS/Register/register[1][30] ), .S0(
        n6012), .Y(\i_MIPS/Register/n1106 ) );
  CLKMX2X2 U12722 ( .A(n5458), .B(\i_MIPS/Register/register[1][5] ), .S0(n6012), .Y(\i_MIPS/Register/n1081 ) );
  CLKMX2X2 U12723 ( .A(n5460), .B(\i_MIPS/Register/register[2][30] ), .S0(
        n6010), .Y(\i_MIPS/Register/n1074 ) );
  CLKMX2X2 U12724 ( .A(n5458), .B(\i_MIPS/Register/register[2][5] ), .S0(n6010), .Y(\i_MIPS/Register/n1049 ) );
  CLKMX2X2 U12725 ( .A(n5460), .B(\i_MIPS/Register/register[3][30] ), .S0(
        n6008), .Y(\i_MIPS/Register/n1042 ) );
  CLKMX2X2 U12726 ( .A(n5458), .B(\i_MIPS/Register/register[3][5] ), .S0(n6008), .Y(\i_MIPS/Register/n1017 ) );
  CLKMX2X2 U12727 ( .A(n5460), .B(\i_MIPS/Register/register[4][30] ), .S0(
        n6006), .Y(\i_MIPS/Register/n1010 ) );
  CLKMX2X2 U12728 ( .A(n5458), .B(\i_MIPS/Register/register[4][5] ), .S0(n6006), .Y(\i_MIPS/Register/n985 ) );
  CLKMX2X2 U12729 ( .A(n5460), .B(\i_MIPS/Register/register[5][30] ), .S0(
        n6004), .Y(\i_MIPS/Register/n978 ) );
  CLKMX2X2 U12730 ( .A(n5458), .B(\i_MIPS/Register/register[5][5] ), .S0(n6004), .Y(\i_MIPS/Register/n953 ) );
  CLKMX2X2 U12731 ( .A(n5460), .B(\i_MIPS/Register/register[6][30] ), .S0(
        n6002), .Y(\i_MIPS/Register/n946 ) );
  CLKMX2X2 U12732 ( .A(n5458), .B(\i_MIPS/Register/register[6][5] ), .S0(n6002), .Y(\i_MIPS/Register/n921 ) );
  CLKMX2X2 U12733 ( .A(n5461), .B(\i_MIPS/Register/register[7][30] ), .S0(
        n6000), .Y(\i_MIPS/Register/n914 ) );
  CLKMX2X2 U12734 ( .A(n5459), .B(\i_MIPS/Register/register[7][5] ), .S0(n6000), .Y(\i_MIPS/Register/n889 ) );
  CLKMX2X2 U12735 ( .A(n5460), .B(\i_MIPS/Register/register[8][30] ), .S0(
        n5998), .Y(\i_MIPS/Register/n882 ) );
  CLKMX2X2 U12736 ( .A(n5458), .B(\i_MIPS/Register/register[8][5] ), .S0(n5998), .Y(\i_MIPS/Register/n857 ) );
  CLKMX2X2 U12737 ( .A(n5460), .B(\i_MIPS/Register/register[9][30] ), .S0(
        n5996), .Y(\i_MIPS/Register/n850 ) );
  CLKMX2X2 U12738 ( .A(n5458), .B(\i_MIPS/Register/register[9][5] ), .S0(n5996), .Y(\i_MIPS/Register/n825 ) );
  CLKMX2X2 U12739 ( .A(n5460), .B(\i_MIPS/Register/register[10][30] ), .S0(
        n5994), .Y(\i_MIPS/Register/n818 ) );
  CLKMX2X2 U12740 ( .A(n5458), .B(\i_MIPS/Register/register[10][5] ), .S0(
        n5994), .Y(\i_MIPS/Register/n793 ) );
  CLKMX2X2 U12741 ( .A(n5461), .B(\i_MIPS/Register/register[11][30] ), .S0(
        n5992), .Y(\i_MIPS/Register/n786 ) );
  CLKMX2X2 U12742 ( .A(n5459), .B(\i_MIPS/Register/register[11][5] ), .S0(
        n5992), .Y(\i_MIPS/Register/n761 ) );
  CLKMX2X2 U12743 ( .A(n5460), .B(\i_MIPS/Register/register[12][30] ), .S0(
        n5990), .Y(\i_MIPS/Register/n754 ) );
  CLKMX2X2 U12744 ( .A(n5458), .B(\i_MIPS/Register/register[12][5] ), .S0(
        n5990), .Y(\i_MIPS/Register/n729 ) );
  CLKMX2X2 U12745 ( .A(n5460), .B(\i_MIPS/Register/register[13][30] ), .S0(
        n5988), .Y(\i_MIPS/Register/n722 ) );
  CLKMX2X2 U12746 ( .A(n5458), .B(\i_MIPS/Register/register[13][5] ), .S0(
        n5988), .Y(\i_MIPS/Register/n697 ) );
  CLKMX2X2 U12747 ( .A(n5460), .B(\i_MIPS/Register/register[14][30] ), .S0(
        n5986), .Y(\i_MIPS/Register/n690 ) );
  CLKMX2X2 U12748 ( .A(n5458), .B(\i_MIPS/Register/register[14][5] ), .S0(
        n5986), .Y(\i_MIPS/Register/n665 ) );
  CLKMX2X2 U12749 ( .A(n5461), .B(\i_MIPS/Register/register[15][30] ), .S0(
        n5984), .Y(\i_MIPS/Register/n658 ) );
  CLKMX2X2 U12750 ( .A(n5459), .B(\i_MIPS/Register/register[15][5] ), .S0(
        n5984), .Y(\i_MIPS/Register/n633 ) );
  CLKMX2X2 U12751 ( .A(n5461), .B(\i_MIPS/Register/register[16][30] ), .S0(
        n5982), .Y(\i_MIPS/Register/n626 ) );
  CLKMX2X2 U12752 ( .A(n5459), .B(\i_MIPS/Register/register[16][5] ), .S0(
        n5982), .Y(\i_MIPS/Register/n601 ) );
  CLKMX2X2 U12753 ( .A(n5461), .B(\i_MIPS/Register/register[17][30] ), .S0(
        n5980), .Y(\i_MIPS/Register/n594 ) );
  CLKMX2X2 U12754 ( .A(n5459), .B(\i_MIPS/Register/register[17][5] ), .S0(
        n5980), .Y(\i_MIPS/Register/n569 ) );
  CLKMX2X2 U12755 ( .A(n5461), .B(\i_MIPS/Register/register[18][30] ), .S0(
        n5978), .Y(\i_MIPS/Register/n562 ) );
  CLKMX2X2 U12756 ( .A(n5459), .B(\i_MIPS/Register/register[18][5] ), .S0(
        n5978), .Y(\i_MIPS/Register/n537 ) );
  CLKMX2X2 U12757 ( .A(n5460), .B(\i_MIPS/Register/register[19][30] ), .S0(
        n5976), .Y(\i_MIPS/Register/n530 ) );
  CLKMX2X2 U12758 ( .A(n5459), .B(\i_MIPS/Register/register[19][5] ), .S0(
        n5976), .Y(\i_MIPS/Register/n505 ) );
  CLKMX2X2 U12759 ( .A(n5461), .B(\i_MIPS/Register/register[20][30] ), .S0(
        n5974), .Y(\i_MIPS/Register/n498 ) );
  CLKMX2X2 U12760 ( .A(n5459), .B(\i_MIPS/Register/register[20][5] ), .S0(
        n5974), .Y(\i_MIPS/Register/n473 ) );
  CLKMX2X2 U12761 ( .A(n5460), .B(\i_MIPS/Register/register[21][30] ), .S0(
        n5972), .Y(\i_MIPS/Register/n466 ) );
  CLKMX2X2 U12762 ( .A(n5458), .B(\i_MIPS/Register/register[21][5] ), .S0(
        n5972), .Y(\i_MIPS/Register/n441 ) );
  CLKMX2X2 U12763 ( .A(n5461), .B(\i_MIPS/Register/register[22][30] ), .S0(
        n5970), .Y(\i_MIPS/Register/n434 ) );
  CLKMX2X2 U12764 ( .A(n5459), .B(\i_MIPS/Register/register[22][5] ), .S0(
        n5970), .Y(\i_MIPS/Register/n409 ) );
  CLKMX2X2 U12765 ( .A(n5461), .B(\i_MIPS/Register/register[23][30] ), .S0(
        n5968), .Y(\i_MIPS/Register/n402 ) );
  CLKMX2X2 U12766 ( .A(n5459), .B(\i_MIPS/Register/register[23][5] ), .S0(
        n5968), .Y(\i_MIPS/Register/n377 ) );
  CLKMX2X2 U12767 ( .A(n5461), .B(\i_MIPS/Register/register[24][30] ), .S0(
        n5966), .Y(\i_MIPS/Register/n370 ) );
  CLKMX2X2 U12768 ( .A(n5459), .B(\i_MIPS/Register/register[24][5] ), .S0(
        n5966), .Y(\i_MIPS/Register/n345 ) );
  CLKMX2X2 U12769 ( .A(n5461), .B(\i_MIPS/Register/register[25][30] ), .S0(
        n5964), .Y(\i_MIPS/Register/n338 ) );
  CLKMX2X2 U12770 ( .A(n5459), .B(\i_MIPS/Register/register[25][5] ), .S0(
        n5964), .Y(\i_MIPS/Register/n313 ) );
  CLKMX2X2 U12771 ( .A(n5461), .B(\i_MIPS/Register/register[26][30] ), .S0(
        n5962), .Y(\i_MIPS/Register/n306 ) );
  CLKMX2X2 U12772 ( .A(n5459), .B(\i_MIPS/Register/register[26][5] ), .S0(
        n5962), .Y(\i_MIPS/Register/n281 ) );
  CLKMX2X2 U12773 ( .A(n5461), .B(\i_MIPS/Register/register[27][30] ), .S0(
        n5960), .Y(\i_MIPS/Register/n274 ) );
  CLKMX2X2 U12774 ( .A(n5458), .B(\i_MIPS/Register/register[27][5] ), .S0(
        n5960), .Y(\i_MIPS/Register/n249 ) );
  CLKMX2X2 U12775 ( .A(n5461), .B(\i_MIPS/Register/register[28][30] ), .S0(
        n5958), .Y(\i_MIPS/Register/n242 ) );
  CLKMX2X2 U12776 ( .A(n5459), .B(\i_MIPS/Register/register[28][5] ), .S0(
        n5958), .Y(\i_MIPS/Register/n217 ) );
  CLKMX2X2 U12777 ( .A(n5460), .B(\i_MIPS/Register/register[29][30] ), .S0(
        n5956), .Y(\i_MIPS/Register/n210 ) );
  CLKMX2X2 U12778 ( .A(n5459), .B(\i_MIPS/Register/register[29][5] ), .S0(
        n5956), .Y(\i_MIPS/Register/n185 ) );
  CLKMX2X2 U12779 ( .A(n5461), .B(\i_MIPS/Register/register[30][30] ), .S0(
        n5954), .Y(\i_MIPS/Register/n178 ) );
  CLKMX2X2 U12780 ( .A(n5459), .B(\i_MIPS/Register/register[30][5] ), .S0(
        n5954), .Y(\i_MIPS/Register/n153 ) );
  MX2XL U12781 ( .A(n11), .B(\i_MIPS/Sign_Extend[0] ), .S0(n3588), .Y(
        \i_MIPS/n448 ) );
  MX2XL U12782 ( .A(n10430), .B(n3907), .S0(n3589), .Y(\i_MIPS/n317 ) );
  CLKINVX1 U12783 ( .A(\i_MIPS/n194 ), .Y(n10430) );
  MX2XL U12784 ( .A(\i_MIPS/ID_EX[85] ), .B(\i_MIPS/Sign_Extend[12] ), .S0(
        n3595), .Y(\i_MIPS/n436 ) );
  NAND3BXL U12785 ( .AN(net105433), .B(net105434), .C(net105435), .Y(n10348)
         );
  INVXL U12786 ( .A(net105436), .Y(net105433) );
  XOR3XL U12787 ( .A(\i_MIPS/IF_ID[4] ), .B(\i_MIPS/Sign_Extend[2] ), .C(n4768), .Y(n10937) );
  XOR3XL U12788 ( .A(\i_MIPS/IF_ID[3] ), .B(\i_MIPS/Sign_Extend[1] ), .C(
        n10134), .Y(n9735) );
  AOI2BB1XL U12789 ( .A0N(\i_MIPS/PC/n5 ), .A1N(net115789), .B0(n9732), .Y(
        n9733) );
  AO22X1 U12790 ( .A0(n5555), .A1(n10768), .B0(n11054), .B1(
        \i_MIPS/Sign_Extend[1] ), .Y(n9732) );
  AO22X1 U12791 ( .A0(n5556), .A1(n10811), .B0(n11054), .B1(
        \i_MIPS/Sign_Extend[11] ), .Y(n10482) );
  XOR3XL U12792 ( .A(\i_MIPS/IF_ID[9] ), .B(n1287), .C(n4767), .Y(n10161) );
  AO22X1 U12793 ( .A0(n5555), .A1(n10618), .B0(n11054), .B1(n1287), .Y(n10159)
         );
  AO22X1 U12794 ( .A0(n5556), .A1(n10698), .B0(n11054), .B1(n10355), .Y(n10356) );
  CLKINVX1 U12795 ( .A(\i_MIPS/n500 ), .Y(n10355) );
  XOR3XL U12796 ( .A(\i_MIPS/IF_ID[27] ), .B(n6016), .C(n10529), .Y(n10388) );
  AO22X1 U12797 ( .A0(n5556), .A1(n3888), .B0(n11054), .B1(n3001), .Y(n10386)
         );
  AO22X1 U12798 ( .A0(n5555), .A1(n10528), .B0(n11054), .B1(
        \i_MIPS/Sign_Extend[8] ), .Y(n10169) );
  AO22X1 U12799 ( .A0(n5555), .A1(n10659), .B0(n11054), .B1(n2948), .Y(n10148)
         );
  XOR3XL U12800 ( .A(\i_MIPS/IF_ID[12] ), .B(\i_MIPS/Sign_Extend[10] ), .C(
        n4770), .Y(n10476) );
  AO22X1 U12801 ( .A0(n5556), .A1(n10473), .B0(n11054), .B1(
        \i_MIPS/Sign_Extend[10] ), .Y(n10474) );
  AO22X1 U12802 ( .A0(n5555), .A1(n10511), .B0(n11054), .B1(
        \i_MIPS/Sign_Extend[14] ), .Y(n10274) );
  XOR3XL U12803 ( .A(\i_MIPS/IF_ID[26] ), .B(n6016), .C(n4808), .Y(n10381) );
  AOI2BB1XL U12804 ( .A0N(\i_MIPS/PC/n28 ), .A1N(net115799), .B0(n10379), .Y(
        n10380) );
  AO22X1 U12805 ( .A0(n5556), .A1(n10443), .B0(n11054), .B1(n10378), .Y(n10379) );
  AO22X1 U12806 ( .A0(n5556), .A1(n10429), .B0(n11054), .B1(n254), .Y(n10366)
         );
  AO22X1 U12807 ( .A0(n5556), .A1(n10825), .B0(n11054), .B1(
        \i_MIPS/Sign_Extend[0] ), .Y(n10826) );
  XOR3XL U12808 ( .A(\i_MIPS/IF_ID[6] ), .B(n168), .C(n4766), .Y(n10872) );
  AO22X1 U12809 ( .A0(n5555), .A1(n11055), .B0(n11054), .B1(n11053), .Y(n11057) );
  AO22X1 U12810 ( .A0(n5556), .A1(n10349), .B0(n11054), .B1(net114081), .Y(
        n10343) );
  AO22X1 U12811 ( .A0(n5555), .A1(n10416), .B0(n11054), .B1(net105477), .Y(
        n10325) );
  MX2XL U12812 ( .A(n12971), .B(n3956), .S0(n3597), .Y(\i_MIPS/n385 ) );
  MX2XL U12813 ( .A(n12956), .B(n4053), .S0(n3599), .Y(\i_MIPS/n370 ) );
  MX2XL U12814 ( .A(n12969), .B(net105167), .S0(n3601), .Y(\i_MIPS/n383 ) );
  MX2XL U12815 ( .A(n12973), .B(n3980), .S0(n3599), .Y(\i_MIPS/n387 ) );
  MX2XL U12816 ( .A(n12961), .B(net105313), .S0(n3591), .Y(\i_MIPS/n375 ) );
  NAND2BX1 U12817 ( .AN(n7744), .B(\i_MIPS/ID_EX_3 ), .Y(net36639) );
  AOI33X1 U12818 ( .A0(\i_MIPS/Hazard_detection/n7 ), .A1(n7743), .A2(n7742), 
        .B0(\i_MIPS/Hazard_detection/n4 ), .B1(n7741), .B2(n7740), .Y(n7744)
         );
  XOR2XL U12819 ( .A(\i_MIPS/n500 ), .B(\i_MIPS/ID_EX[111] ), .Y(n7742) );
  AO22XL U12820 ( .A0(n3032), .A1(n3589), .B0(n3586), .B1(\i_MIPS/ALUOp[1] ), 
        .Y(\i_MIPS/n401 ) );
  AO22XL U12821 ( .A0(n11575), .A1(n3595), .B0(n3586), .B1(\i_MIPS/ID_EX_5 ), 
        .Y(\i_MIPS/n408 ) );
  CLKINVX1 U12822 ( .A(n11588), .Y(n11575) );
  BUFX20 U12823 ( .A(n3976), .Y(n5051) );
  AO21XL U12824 ( .A0(\i_MIPS/ID_EX[93] ), .A1(n3586), .B0(n4642), .Y(
        \i_MIPS/n428 ) );
  AO21XL U12825 ( .A0(\i_MIPS/ID_EX[95] ), .A1(n3586), .B0(n4642), .Y(
        \i_MIPS/n426 ) );
  AO21XL U12826 ( .A0(\i_MIPS/ID_EX[96] ), .A1(n3586), .B0(n4642), .Y(
        \i_MIPS/n425 ) );
  AO21XL U12827 ( .A0(\i_MIPS/ID_EX[98] ), .A1(n3586), .B0(n4642), .Y(
        \i_MIPS/n423 ) );
  AO21XL U12828 ( .A0(\i_MIPS/ID_EX[100] ), .A1(n3586), .B0(n4642), .Y(
        \i_MIPS/n421 ) );
  AO21XL U12829 ( .A0(\i_MIPS/ID_EX[94] ), .A1(n3586), .B0(n4642), .Y(
        \i_MIPS/n427 ) );
  AO21XL U12830 ( .A0(\i_MIPS/ID_EX[97] ), .A1(n3586), .B0(n4642), .Y(
        \i_MIPS/n424 ) );
  AO21XL U12831 ( .A0(\i_MIPS/ID_EX[99] ), .A1(n3586), .B0(n4642), .Y(
        \i_MIPS/n422 ) );
  AO21XL U12832 ( .A0(\i_MIPS/ID_EX[101] ), .A1(n3586), .B0(n4642), .Y(
        \i_MIPS/n420 ) );
  AO21XL U12833 ( .A0(\i_MIPS/ID_EX[102] ), .A1(n3586), .B0(n4642), .Y(
        \i_MIPS/n419 ) );
  AO21XL U12834 ( .A0(\i_MIPS/ID_EX[103] ), .A1(n3586), .B0(n4642), .Y(
        \i_MIPS/n418 ) );
  AO21XL U12835 ( .A0(\i_MIPS/ID_EX[104] ), .A1(n3586), .B0(n4642), .Y(
        \i_MIPS/n417 ) );
  AND2X2 U12836 ( .A(n9731), .B(\i_MIPS/IR[26] ), .Y(n4837) );
  AND3X2 U12837 ( .A(\i_MIPS/Register/n120 ), .B(\i_MIPS/Reg_W[3] ), .C(
        \i_MIPS/Reg_W[4] ), .Y(\i_MIPS/Register/n104 ) );
  NAND3BX1 U12838 ( .AN(n9819), .B(\i_MIPS/IR[29] ), .C(n9818), .Y(
        \i_MIPS/Control/n14 ) );
  AOI2BB1X1 U12839 ( .A0N(n9817), .A1N(n9816), .B0(\i_MIPS/IR[30] ), .Y(n9818)
         );
  XOR2X1 U12840 ( .A(n9815), .B(n9814), .Y(n9819) );
  NAND2X1 U12841 ( .A(n9817), .B(n9816), .Y(n9815) );
  NAND2XL U12842 ( .A(n10138), .B(ICACHE_addr[3]), .Y(n9936) );
  NAND2XL U12843 ( .A(n10179), .B(ICACHE_addr[7]), .Y(n10168) );
  NAND2XL U12844 ( .A(n10471), .B(ICACHE_addr[9]), .Y(n10472) );
  NAND2XL U12845 ( .A(n10158), .B(ICACHE_addr[5]), .Y(n10147) );
  NAND2XL U12846 ( .A(n10491), .B(ICACHE_addr[11]), .Y(n10492) );
  NOR2BX1 U12847 ( .AN(\i_MIPS/EX_MEM_0 ), .B(\i_MIPS/EX_MEM_74 ), .Y(
        \i_MIPS/Register/n120 ) );
  CLKINVX1 U12848 ( .A(\i_MIPS/IR[28] ), .Y(n9820) );
  NAND3BX1 U12849 ( .AN(n9603), .B(\i_MIPS/IR[27] ), .C(n9820), .Y(n9654) );
  CLKINVX1 U12850 ( .A(\i_MIPS/IR[26] ), .Y(n9817) );
  CLKINVX1 U12851 ( .A(\i_MIPS/IR[27] ), .Y(n9600) );
  CLKINVX1 U12852 ( .A(mem_ready_D), .Y(n11539) );
  CLKINVX1 U12853 ( .A(mem_ready_I), .Y(n11540) );
  CLKBUFX3 U12854 ( .A(\i_MIPS/jump_addr[22] ), .Y(net114081) );
  XOR2X1 U12855 ( .A(\i_MIPS/n506 ), .B(\i_MIPS/jump_addr[30] ), .Y(n10582) );
  CLKINVX1 U12856 ( .A(\i_MIPS/jump_addr[29] ), .Y(n10577) );
  NOR2X1 U12857 ( .A(n9823), .B(n9822), .Y(n11574) );
  CLKINVX1 U12858 ( .A(\i_MIPS/jump_addr[30] ), .Y(n10723) );
  CLKINVX1 U12859 ( .A(\i_MIPS/n524 ), .Y(n10574) );
  CLKINVX1 U12860 ( .A(\i_MIPS/n525 ), .Y(n10537) );
  CLKINVX1 U12861 ( .A(\i_MIPS/n505 ), .Y(n10294) );
  CLKINVX6 U12862 ( .A(n12865), .Y(n4838) );
  INVX20 U12863 ( .A(n4838), .Y(mem_addr_I[21]) );
  AO22X1 U12864 ( .A0(ICACHE_addr[20]), .A1(mem_read_I), .B0(mem_write_I), 
        .B1(n11362), .Y(n12864) );
  INVX20 U12865 ( .A(n4842), .Y(mem_addr_I[23]) );
  AO22X1 U12866 ( .A0(ICACHE_addr[22]), .A1(mem_read_I), .B0(mem_write_I), 
        .B1(n11364), .Y(n12862) );
  AO22X1 U12867 ( .A0(ICACHE_addr[23]), .A1(mem_read_I), .B0(mem_write_I), 
        .B1(n11365), .Y(n12861) );
  AO22X1 U12868 ( .A0(ICACHE_addr[24]), .A1(mem_read_I), .B0(mem_write_I), 
        .B1(n11366), .Y(n12860) );
  CLKINVX6 U12869 ( .A(n12858), .Y(n4852) );
  INVX20 U12870 ( .A(n4852), .Y(mem_addr_I[28]) );
  AO22X1 U12871 ( .A0(ICACHE_addr[27]), .A1(mem_read_I), .B0(mem_write_I), 
        .B1(n11369), .Y(n12857) );
  AO22X1 U12872 ( .A0(ICACHE_addr[28]), .A1(mem_read_I), .B0(mem_write_I), 
        .B1(n11370), .Y(n12856) );
  AO22X1 U12873 ( .A0(ICACHE_addr[29]), .A1(mem_read_I), .B0(mem_write_I), 
        .B1(n11371), .Y(n12855) );
  MX2XL U12874 ( .A(n3608), .B(n4100), .S0(n3597), .Y(\i_MIPS/n347 ) );
  MX2XL U12875 ( .A(DCACHE_addr[21]), .B(n4101), .S0(n3599), .Y(\i_MIPS/n376 )
         );
  AND2XL U12876 ( .A(DCACHE_addr[3]), .B(n11507), .Y(n12849) );
  OAI211X2 U12877 ( .A0(n6648), .A1(n6647), .B0(n4835), .C0(net112544), .Y(
        n8698) );
  MX2XL U12878 ( .A(n10541), .B(n3706), .S0(n3603), .Y(\i_MIPS/n311 ) );
  AO22X1 U12879 ( .A0(DCACHE_addr[18]), .A1(n11534), .B0(n5042), .B1(n11522), 
        .Y(n12847) );
  AND2XL U12880 ( .A(n5044), .B(n11443), .Y(n12853) );
  AND2XL U12881 ( .A(n5042), .B(n11444), .Y(n12852) );
  AND2XL U12882 ( .A(n5043), .B(n11466), .Y(n12851) );
  INVX12 U12883 ( .A(n4920), .Y(DCACHE_addr[17]) );
  AO22X1 U12884 ( .A0(DCACHE_addr[16]), .A1(n11534), .B0(n5042), .B1(n11520), 
        .Y(n12848) );
  OAI221XL U12885 ( .A0(net107854), .A1(net117709), .B0(net107855), .B1(
        net117731), .C0(n3949), .Y(n4937) );
  AND2XL U12886 ( .A(n5043), .B(n11493), .Y(n12850) );
  NAND2X8 U12887 ( .A(\i_MIPS/n264 ), .B(\i_MIPS/n245 ), .Y(n10979) );
  OAI221XL U12888 ( .A0(net112328), .A1(net117713), .B0(net112329), .B1(
        net117733), .C0(net112330), .Y(n4987) );
  OA22X2 U12889 ( .A0(n5918), .A1(n1330), .B0(n5876), .B1(n2983), .Y(n11123)
         );
  XOR2X4 U12890 ( .A(ICACHE_addr[19]), .B(n11202), .Y(n11603) );
  CLKAND2X12 U12891 ( .A(n5048), .B(n11342), .Y(mem_wdata_I[127]) );
  INVX12 U12892 ( .A(net118925), .Y(net118926) );
  INVX12 U12893 ( .A(n5006), .Y(DCACHE_addr[9]) );
  INVX12 U12894 ( .A(n5008), .Y(DCACHE_addr[27]) );
  NAND2X1 U12895 ( .A(DCACHE_addr[1]), .B(n5190), .Y(net106674) );
  NAND2X1 U12896 ( .A(n11034), .B(n3718), .Y(n11524) );
  AO22X1 U12897 ( .A0(DCACHE_addr[21]), .A1(mem_read_D), .B0(mem_write_D), 
        .B1(n11525), .Y(n5011) );
  AO22X1 U12898 ( .A0(n12961), .A1(mem_read_D), .B0(mem_write_D), .B1(n11526), 
        .Y(n5012) );
  NAND2X1 U12899 ( .A(n11018), .B(n11017), .Y(n11526) );
  AO22X1 U12900 ( .A0(DCACHE_addr[23]), .A1(mem_read_D), .B0(mem_write_D), 
        .B1(n11527), .Y(n5013) );
  NAND2X1 U12901 ( .A(n11032), .B(n11031), .Y(n11527) );
  AO22X1 U12902 ( .A0(n12959), .A1(mem_read_D), .B0(mem_write_D), .B1(n11528), 
        .Y(n5014) );
  AO22X1 U12903 ( .A0(DCACHE_addr[25]), .A1(mem_read_D), .B0(mem_write_D), 
        .B1(n11529), .Y(n5015) );
  AO22X1 U12904 ( .A0(n12956), .A1(mem_read_D), .B0(mem_write_D), .B1(n11531), 
        .Y(n5017) );
  NAND2X1 U12905 ( .A(n11000), .B(n10999), .Y(n11532) );
  NAND2X1 U12906 ( .A(n10991), .B(n10990), .Y(n11533) );
  INVX12 U12907 ( .A(n5021), .Y(DCACHE_addr[24]) );
  INVX12 U12908 ( .A(n5024), .Y(DCACHE_addr[22]) );
  NAND2X1 U12909 ( .A(DCACHE_addr[23]), .B(n5190), .Y(net105288) );
  CLKAND2X12 U12910 ( .A(n5044), .B(n11494), .Y(mem_wdata_D[118]) );
  NAND2X1 U12911 ( .A(DCACHE_addr[25]), .B(n5190), .Y(net105423) );
  NAND2X8 U12912 ( .A(n11218), .B(n6528), .Y(net36572) );
  XOR2X4 U12913 ( .A(ICACHE_addr[20]), .B(n11216), .Y(n11605) );
  NAND3BXL U12914 ( .AN(n3648), .B(n10713), .C(net104830), .Y(n10719) );
  CLKAND2X12 U12915 ( .A(n5044), .B(n11503), .Y(mem_wdata_D[127]) );
  NAND2X8 U12916 ( .A(\i_MIPS/ID_EX[83] ), .B(n6675), .Y(n9316) );
  CLKBUFX20 U12917 ( .A(n11536), .Y(mem_read_I) );
  OA22X4 U12918 ( .A0(n5743), .A1(n2884), .B0(n5672), .B1(n1266), .Y(n6361) );
  OA22X4 U12919 ( .A0(n5838), .A1(n2885), .B0(n5763), .B1(n1267), .Y(n6360) );
  OA22X4 U12920 ( .A0(n138), .A1(n2941), .B0(n5704), .B1(n1290), .Y(n6364) );
  OA22X4 U12921 ( .A0(n5917), .A1(n2942), .B0(n5851), .B1(n1291), .Y(n6362) );
  OA22X4 U12922 ( .A0(n5741), .A1(n2943), .B0(n5672), .B1(n1292), .Y(n6368) );
  OA22X4 U12923 ( .A0(n5928), .A1(n2932), .B0(n5851), .B1(n1293), .Y(n6366) );
  OA22X4 U12924 ( .A0(n5743), .A1(n1299), .B0(n5698), .B1(n3009), .Y(n6372) );
  XOR2X2 U12925 ( .A(n11371), .B(ICACHE_addr[29]), .Y(n6385) );
  OA22X4 U12926 ( .A0(n5895), .A1(n1300), .B0(n5880), .B1(n2966), .Y(n6376) );
  OA22X4 U12927 ( .A0(n5719), .A1(n2973), .B0(n5702), .B1(n1295), .Y(n6381) );
  OA22X4 U12928 ( .A0(n5920), .A1(n1301), .B0(n5853), .B1(n2967), .Y(n6379) );
  OA22X4 U12929 ( .A0(n5401), .A1(n434), .B0(n5444), .B1(n2060), .Y(n6496) );
  CLKINVX3 U12930 ( .A(n6499), .Y(n11003) );
  NAND2BX4 U12931 ( .AN(n5406), .B(\D_cache/cache[6][154] ), .Y(n6517) );
  NAND2BX4 U12932 ( .AN(n5219), .B(\D_cache/cache[1][154] ), .Y(n6521) );
  NAND2BX4 U12933 ( .AN(n5303), .B(\D_cache/cache[3][154] ), .Y(n6519) );
  OR2X8 U12934 ( .A(n6524), .B(n6523), .Y(n11374) );
  OA22X4 U12935 ( .A0(n5746), .A1(n2583), .B0(n5697), .B1(n1077), .Y(n6527) );
  OA22X4 U12936 ( .A0(n5834), .A1(n2584), .B0(n5763), .B1(n1078), .Y(n6526) );
  OA22X4 U12937 ( .A0(n5895), .A1(n1286), .B0(n5880), .B1(n2935), .Y(n6525) );
  NAND2X2 U12938 ( .A(n4738), .B(n9606), .Y(n11079) );
  NAND4X2 U12939 ( .A(n6641), .B(n6640), .C(n6639), .D(n6638), .Y(net107196)
         );
  CLKINVX6 U12940 ( .A(\i_MIPS/forward_unit/n10 ), .Y(n6643) );
  OAI2BB1X4 U12941 ( .A0N(n6651), .A1N(n6650), .B0(n6649), .Y(n6669) );
  NAND2X2 U12942 ( .A(\i_MIPS/ALUin1[14] ), .B(n6696), .Y(net110406) );
  NAND2X2 U12943 ( .A(n6691), .B(n300), .Y(net109179) );
  NAND2X2 U12944 ( .A(\i_MIPS/ALUin1[25] ), .B(n144), .Y(n11103) );
  OAI31X2 U12945 ( .A0(n6925), .A1(n6924), .A2(n6923), .B0(n6922), .Y(n7592)
         );
  OAI31X2 U12946 ( .A0(n7060), .A1(n7059), .A2(n7058), .B0(n7057), .Y(
        net104868) );
  OAI221X2 U12947 ( .A0(n7815), .A1(net107138), .B0(n7838), .B1(net107141), 
        .C0(n7814), .Y(net105179) );
  NAND3BX2 U12948 ( .AN(n7866), .B(net117745), .C(n7865), .Y(n7872) );
  AOI2BB1X2 U12949 ( .A0N(net108290), .A1N(n8978), .B0(n8977), .Y(n8981) );
  AO22X4 U12950 ( .A0(n10769), .A1(net118215), .B0(net118225), .B1(n9079), .Y(
        net108101) );
  OA22X4 U12951 ( .A0(n3979), .A1(n3878), .B0(n10755), .B1(n4495), .Y(n9096)
         );
  CLKINVX3 U12952 ( .A(n9305), .Y(n9307) );
  AO22X4 U12953 ( .A0(DCACHE_addr[28]), .A1(n5190), .B0(n4407), .B1(n9421), 
        .Y(n10075) );
  OAI222X2 U12954 ( .A0(n9466), .A1(net117709), .B0(n5462), .B1(net117723), 
        .C0(n9487), .C1(net117731), .Y(n10590) );
  NAND2X2 U12955 ( .A(n9945), .B(n4689), .Y(n9956) );
  NAND2X2 U12956 ( .A(n4737), .B(n9958), .Y(n10970) );
  CLKINVX3 U12957 ( .A(n10164), .Y(n10176) );
  CLKINVX3 U12958 ( .A(n10938), .Y(n10939) );
  OA22X4 U12959 ( .A0(n5830), .A1(n2974), .B0(n5785), .B1(n1322), .Y(n11115)
         );
  OA22X4 U12960 ( .A0(n5830), .A1(n2975), .B0(n5785), .B1(n1323), .Y(n11120)
         );
  OA22X4 U12961 ( .A0(n5832), .A1(n2976), .B0(n5786), .B1(n1324), .Y(n11157)
         );
  OA22X4 U12962 ( .A0(n5832), .A1(n2977), .B0(n5796), .B1(n1325), .Y(n11169)
         );
  OA22X4 U12963 ( .A0(n5832), .A1(n2978), .B0(n5796), .B1(n1326), .Y(n11174)
         );
  OA22X4 U12964 ( .A0(n5832), .A1(n2979), .B0(n5762), .B1(n1327), .Y(n11179)
         );
  OA22X4 U12965 ( .A0(n138), .A1(n2933), .B0(n5696), .B1(n1296), .Y(n11200) );
  OA22X4 U12966 ( .A0(n5838), .A1(n2980), .B0(n5787), .B1(n1328), .Y(n11199)
         );
  OA22X4 U12967 ( .A0(n138), .A1(n3013), .B0(n5696), .B1(n1343), .Y(n11205) );
  OA22X4 U12968 ( .A0(n5807), .A1(n2155), .B0(n5787), .B1(n531), .Y(n11212) );
  AO22X4 U12969 ( .A0(ICACHE_addr[5]), .A1(mem_read_I), .B0(n5046), .B1(n11347), .Y(n12878) );
endmodule

